module basic_5000_50000_5000_5_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
nor U0 (N_0,In_3993,In_4250);
and U1 (N_1,In_2023,In_4190);
and U2 (N_2,In_2305,In_4483);
nand U3 (N_3,In_3727,In_3797);
or U4 (N_4,In_286,In_833);
nor U5 (N_5,In_4602,In_2848);
or U6 (N_6,In_3218,In_2304);
or U7 (N_7,In_490,In_4967);
and U8 (N_8,In_4732,In_4287);
and U9 (N_9,In_814,In_1092);
and U10 (N_10,In_3068,In_1831);
or U11 (N_11,In_4750,In_158);
and U12 (N_12,In_3953,In_119);
and U13 (N_13,In_4315,In_3470);
nor U14 (N_14,In_2863,In_2051);
or U15 (N_15,In_848,In_830);
and U16 (N_16,In_3633,In_128);
or U17 (N_17,In_4715,In_4993);
nand U18 (N_18,In_690,In_2237);
or U19 (N_19,In_4301,In_2829);
nor U20 (N_20,In_265,In_4857);
and U21 (N_21,In_4242,In_1738);
xnor U22 (N_22,In_577,In_4837);
and U23 (N_23,In_3612,In_1191);
nor U24 (N_24,In_221,In_1624);
nor U25 (N_25,In_1618,In_750);
or U26 (N_26,In_4720,In_4839);
nand U27 (N_27,In_988,In_2668);
xnor U28 (N_28,In_596,In_4832);
and U29 (N_29,In_3145,In_3021);
and U30 (N_30,In_2802,In_4812);
nand U31 (N_31,In_3559,In_2257);
and U32 (N_32,In_2739,In_1921);
and U33 (N_33,In_3093,In_2590);
nand U34 (N_34,In_3434,In_1175);
or U35 (N_35,In_2118,In_923);
or U36 (N_36,In_650,In_3188);
nor U37 (N_37,In_2797,In_1623);
nor U38 (N_38,In_374,In_3087);
xnor U39 (N_39,In_4643,In_1833);
nor U40 (N_40,In_3579,In_124);
and U41 (N_41,In_2277,In_4788);
and U42 (N_42,In_2620,In_1080);
nand U43 (N_43,In_4476,In_795);
or U44 (N_44,In_1221,In_288);
or U45 (N_45,In_2775,In_3252);
or U46 (N_46,In_4859,In_1401);
nor U47 (N_47,In_4659,In_4655);
nor U48 (N_48,In_1448,In_4161);
or U49 (N_49,In_416,In_1453);
and U50 (N_50,In_2597,In_60);
nand U51 (N_51,In_2883,In_1415);
or U52 (N_52,In_1145,In_1419);
and U53 (N_53,In_3983,In_2140);
xnor U54 (N_54,In_3221,In_4464);
nor U55 (N_55,In_501,In_2814);
xor U56 (N_56,In_1678,In_2933);
nor U57 (N_57,In_3994,In_2199);
xor U58 (N_58,In_3508,In_4105);
and U59 (N_59,In_3687,In_1369);
or U60 (N_60,In_3195,In_3905);
nor U61 (N_61,In_572,In_2343);
or U62 (N_62,In_4463,In_3943);
nand U63 (N_63,In_406,In_3113);
xnor U64 (N_64,In_4961,In_1484);
nor U65 (N_65,In_1840,In_3928);
and U66 (N_66,In_4754,In_2423);
or U67 (N_67,In_4546,In_3914);
xor U68 (N_68,In_3705,In_3151);
and U69 (N_69,In_3133,In_2669);
nand U70 (N_70,In_1841,In_4906);
nand U71 (N_71,In_4776,In_1333);
nor U72 (N_72,In_3383,In_4639);
nand U73 (N_73,In_963,In_4415);
nor U74 (N_74,In_4699,In_195);
xor U75 (N_75,In_277,In_4321);
and U76 (N_76,In_4127,In_4605);
or U77 (N_77,In_560,In_4890);
nor U78 (N_78,In_2674,In_620);
and U79 (N_79,In_805,In_1220);
nor U80 (N_80,In_2671,In_700);
or U81 (N_81,In_3898,In_956);
xnor U82 (N_82,In_737,In_1542);
nor U83 (N_83,In_4418,In_1797);
nor U84 (N_84,In_2654,In_1003);
and U85 (N_85,In_3251,In_2230);
or U86 (N_86,In_2033,In_66);
and U87 (N_87,In_4998,In_3351);
nor U88 (N_88,In_2129,In_4196);
or U89 (N_89,In_1929,In_1256);
and U90 (N_90,In_3591,In_1262);
nand U91 (N_91,In_1413,In_4638);
nor U92 (N_92,In_2449,In_2910);
or U93 (N_93,In_4099,In_2354);
nor U94 (N_94,In_3032,In_4133);
or U95 (N_95,In_4852,In_685);
or U96 (N_96,In_3833,In_2349);
nand U97 (N_97,In_3426,In_1231);
and U98 (N_98,In_1507,In_3749);
nor U99 (N_99,In_3874,In_4875);
and U100 (N_100,In_4063,In_3134);
and U101 (N_101,In_3842,In_426);
or U102 (N_102,In_2563,In_2397);
and U103 (N_103,In_2228,In_4809);
nor U104 (N_104,In_952,In_1423);
nand U105 (N_105,In_3205,In_1988);
nor U106 (N_106,In_1025,In_3788);
and U107 (N_107,In_1596,In_4888);
or U108 (N_108,In_2582,In_1053);
nor U109 (N_109,In_4,In_1059);
nand U110 (N_110,In_2243,In_4977);
and U111 (N_111,In_2715,In_624);
or U112 (N_112,In_4747,In_3206);
nor U113 (N_113,In_1064,In_2725);
and U114 (N_114,In_954,In_2793);
nor U115 (N_115,In_4798,In_3040);
nand U116 (N_116,In_3014,In_3051);
nand U117 (N_117,In_1837,In_4182);
nor U118 (N_118,In_4647,In_1719);
and U119 (N_119,In_2889,In_4762);
and U120 (N_120,In_3223,In_4223);
or U121 (N_121,In_3499,In_3318);
xor U122 (N_122,In_161,In_2955);
nor U123 (N_123,In_1216,In_144);
and U124 (N_124,In_2536,In_4261);
or U125 (N_125,In_215,In_4529);
and U126 (N_126,In_3599,In_3438);
or U127 (N_127,In_4227,In_3873);
nand U128 (N_128,In_216,In_1628);
or U129 (N_129,In_1155,In_205);
xnor U130 (N_130,In_1888,In_3100);
or U131 (N_131,In_2637,In_4279);
xor U132 (N_132,In_2088,In_99);
or U133 (N_133,In_1965,In_2247);
xor U134 (N_134,In_682,In_2111);
nand U135 (N_135,In_4936,In_666);
xnor U136 (N_136,In_4629,In_1827);
nor U137 (N_137,In_2570,In_4158);
or U138 (N_138,In_3877,In_3474);
nand U139 (N_139,In_1537,In_1244);
or U140 (N_140,In_38,In_2571);
or U141 (N_141,In_1062,In_1088);
nor U142 (N_142,In_4586,In_2854);
nor U143 (N_143,In_3148,In_2296);
and U144 (N_144,In_3534,In_3922);
nor U145 (N_145,In_2884,In_3598);
nor U146 (N_146,In_4368,In_969);
nand U147 (N_147,In_2587,In_424);
or U148 (N_148,In_2638,In_3626);
nand U149 (N_149,In_2787,In_1141);
and U150 (N_150,In_2436,In_270);
nand U151 (N_151,In_2031,In_3333);
or U152 (N_152,In_1403,In_3125);
or U153 (N_153,In_2204,In_3791);
or U154 (N_154,In_4517,In_2123);
or U155 (N_155,In_1248,In_3005);
nor U156 (N_156,In_4098,In_537);
or U157 (N_157,In_3452,In_3752);
or U158 (N_158,In_2653,In_1920);
nand U159 (N_159,In_4610,In_2085);
xor U160 (N_160,In_4978,In_2252);
and U161 (N_161,In_2134,In_3819);
nor U162 (N_162,In_2192,In_467);
or U163 (N_163,In_2321,In_291);
xor U164 (N_164,In_4912,In_3437);
nand U165 (N_165,In_932,In_2075);
nor U166 (N_166,In_2487,In_4024);
nand U167 (N_167,In_2062,In_1915);
nand U168 (N_168,In_2401,In_4328);
and U169 (N_169,In_4675,In_1202);
nand U170 (N_170,In_4150,In_422);
and U171 (N_171,In_930,In_2726);
or U172 (N_172,In_3763,In_1967);
nand U173 (N_173,In_759,In_3957);
nand U174 (N_174,In_4664,In_3972);
nand U175 (N_175,In_1309,In_3121);
or U176 (N_176,In_3412,In_3140);
and U177 (N_177,In_2265,In_1326);
xor U178 (N_178,In_4472,In_19);
or U179 (N_179,In_2159,In_2368);
xnor U180 (N_180,In_4646,In_3616);
nor U181 (N_181,In_2960,In_2675);
and U182 (N_182,In_357,In_944);
or U183 (N_183,In_2639,In_2818);
nor U184 (N_184,In_2189,In_4248);
or U185 (N_185,In_3492,In_1568);
xnor U186 (N_186,In_3240,In_4139);
nand U187 (N_187,In_3865,In_2843);
and U188 (N_188,In_3137,In_4892);
nor U189 (N_189,In_533,In_1702);
or U190 (N_190,In_3702,In_3774);
nor U191 (N_191,In_1767,In_3436);
nor U192 (N_192,In_3780,In_959);
or U193 (N_193,In_1363,In_354);
nand U194 (N_194,In_2248,In_2412);
nand U195 (N_195,In_2161,In_2498);
nand U196 (N_196,In_414,In_4184);
or U197 (N_197,In_462,In_2385);
and U198 (N_198,In_278,In_1676);
nand U199 (N_199,In_4830,In_3025);
or U200 (N_200,In_4534,In_1447);
nor U201 (N_201,In_2615,In_1913);
nor U202 (N_202,In_3464,In_4727);
xor U203 (N_203,In_1972,In_768);
or U204 (N_204,In_4652,In_1501);
and U205 (N_205,In_309,In_106);
or U206 (N_206,In_4550,In_3662);
or U207 (N_207,In_2378,In_1261);
and U208 (N_208,In_4760,In_4642);
and U209 (N_209,In_1692,In_1475);
nor U210 (N_210,In_342,In_3544);
nand U211 (N_211,In_1630,In_3408);
xor U212 (N_212,In_3673,In_298);
nor U213 (N_213,In_3253,In_4612);
xnor U214 (N_214,In_2196,In_194);
or U215 (N_215,In_4120,In_3523);
or U216 (N_216,In_731,In_2728);
or U217 (N_217,In_780,In_1928);
nand U218 (N_218,In_2180,In_672);
nand U219 (N_219,In_3688,In_3704);
nor U220 (N_220,In_621,In_246);
or U221 (N_221,In_2408,In_1651);
nand U222 (N_222,In_4613,In_3536);
and U223 (N_223,In_476,In_3399);
nand U224 (N_224,In_1685,In_3476);
or U225 (N_225,In_4866,In_3096);
xor U226 (N_226,In_2493,In_2270);
and U227 (N_227,In_450,In_2737);
nor U228 (N_228,In_4896,In_3185);
nor U229 (N_229,In_2631,In_352);
xor U230 (N_230,In_3389,In_581);
nand U231 (N_231,In_917,In_1566);
nor U232 (N_232,In_4990,In_1587);
nand U233 (N_233,In_989,In_500);
or U234 (N_234,In_1954,In_2393);
or U235 (N_235,In_515,In_1437);
nand U236 (N_236,In_3292,In_2081);
nand U237 (N_237,In_1951,In_3305);
or U238 (N_238,In_4649,In_874);
nor U239 (N_239,In_2577,In_3674);
and U240 (N_240,In_4351,In_4653);
xnor U241 (N_241,In_4902,In_1170);
nand U242 (N_242,In_3012,In_4855);
or U243 (N_243,In_364,In_2014);
or U244 (N_244,In_4778,In_1891);
nor U245 (N_245,In_871,In_2238);
and U246 (N_246,In_4460,In_3696);
nand U247 (N_247,In_4164,In_2913);
xor U248 (N_248,In_3301,In_2741);
and U249 (N_249,In_3933,In_1663);
nand U250 (N_250,In_3855,In_2053);
nand U251 (N_251,In_3467,In_1481);
nand U252 (N_252,In_867,In_4304);
or U253 (N_253,In_182,In_1458);
nand U254 (N_254,In_4174,In_3118);
nand U255 (N_255,In_3701,In_2927);
nand U256 (N_256,In_896,In_1902);
nand U257 (N_257,In_1776,In_3104);
or U258 (N_258,In_4871,In_2488);
nand U259 (N_259,In_3091,In_573);
nand U260 (N_260,In_137,In_2792);
nand U261 (N_261,In_17,In_2137);
nand U262 (N_262,In_3821,In_1657);
or U263 (N_263,In_4543,In_2670);
nand U264 (N_264,In_2037,In_891);
nand U265 (N_265,In_1372,In_3655);
nor U266 (N_266,In_3267,In_4124);
or U267 (N_267,In_1510,In_1107);
or U268 (N_268,In_4052,In_3463);
and U269 (N_269,In_1368,In_1182);
and U270 (N_270,In_769,In_2678);
and U271 (N_271,In_3075,In_2875);
nand U272 (N_272,In_4109,In_3656);
or U273 (N_273,In_746,In_3083);
or U274 (N_274,In_4791,In_1995);
and U275 (N_275,In_2198,In_3827);
and U276 (N_276,In_3281,In_906);
xnor U277 (N_277,In_4309,In_1726);
nand U278 (N_278,In_4393,In_4909);
nor U279 (N_279,In_224,In_3226);
and U280 (N_280,In_98,In_171);
and U281 (N_281,In_1686,In_4352);
or U282 (N_282,In_2092,In_4381);
and U283 (N_283,In_2731,In_4818);
and U284 (N_284,In_1733,In_2372);
or U285 (N_285,In_4341,In_1468);
or U286 (N_286,In_4836,In_1519);
or U287 (N_287,In_4983,In_2322);
and U288 (N_288,In_1117,In_1895);
nor U289 (N_289,In_3472,In_2736);
and U290 (N_290,In_658,In_4195);
nor U291 (N_291,In_2988,In_1304);
and U292 (N_292,In_1658,In_1775);
nand U293 (N_293,In_55,In_3527);
and U294 (N_294,In_3249,In_3047);
nand U295 (N_295,In_2759,In_84);
and U296 (N_296,In_1756,In_4011);
or U297 (N_297,In_2535,In_3154);
and U298 (N_298,In_1329,In_845);
nor U299 (N_299,In_402,In_4380);
or U300 (N_300,In_4660,In_4826);
and U301 (N_301,In_3478,In_4320);
and U302 (N_302,In_860,In_1000);
or U303 (N_303,In_3684,In_745);
or U304 (N_304,In_3921,In_2402);
or U305 (N_305,In_425,In_2026);
and U306 (N_306,In_346,In_1856);
and U307 (N_307,In_720,In_2290);
nor U308 (N_308,In_1177,In_3268);
nor U309 (N_309,In_4975,In_3454);
xnor U310 (N_310,In_126,In_4867);
nand U311 (N_311,In_2478,In_753);
nor U312 (N_312,In_928,In_32);
or U313 (N_313,In_2060,In_1135);
and U314 (N_314,In_1600,In_1858);
or U315 (N_315,In_114,In_1367);
or U316 (N_316,In_3066,In_1901);
and U317 (N_317,In_4670,In_3966);
and U318 (N_318,In_4154,In_242);
nor U319 (N_319,In_3179,In_1905);
nor U320 (N_320,In_1266,In_1161);
and U321 (N_321,In_1679,In_3331);
and U322 (N_322,In_2989,In_4879);
nor U323 (N_323,In_680,In_3120);
and U324 (N_324,In_3988,In_1996);
or U325 (N_325,In_4807,In_2015);
or U326 (N_326,In_3681,In_2516);
and U327 (N_327,In_3679,In_4526);
xor U328 (N_328,In_1994,In_1142);
nand U329 (N_329,In_4014,In_2454);
nor U330 (N_330,In_202,In_1524);
nor U331 (N_331,In_3385,In_1520);
nand U332 (N_332,In_2216,In_262);
nor U333 (N_333,In_2581,In_2844);
nand U334 (N_334,In_1290,In_1680);
or U335 (N_335,In_2229,In_222);
nor U336 (N_336,In_1287,In_1825);
nor U337 (N_337,In_4118,In_825);
nor U338 (N_338,In_3609,In_2356);
nand U339 (N_339,In_1506,In_484);
nand U340 (N_340,In_4581,In_3009);
or U341 (N_341,In_3288,In_4359);
and U342 (N_342,In_2254,In_1004);
or U343 (N_343,In_1260,In_3347);
nor U344 (N_344,In_4492,In_3123);
nand U345 (N_345,In_2086,In_3882);
and U346 (N_346,In_391,In_506);
and U347 (N_347,In_3242,In_1946);
and U348 (N_348,In_4413,In_3329);
nor U349 (N_349,In_1698,In_3871);
or U350 (N_350,In_1695,In_2628);
and U351 (N_351,In_865,In_4443);
or U352 (N_352,In_2207,In_4721);
nand U353 (N_353,In_118,In_3708);
or U354 (N_354,In_1787,In_2016);
or U355 (N_355,In_2231,In_148);
and U356 (N_356,In_4205,In_2179);
nor U357 (N_357,In_4259,In_1527);
and U358 (N_358,In_469,In_2302);
xnor U359 (N_359,In_1662,In_4173);
and U360 (N_360,In_210,In_2365);
or U361 (N_361,In_1132,In_4910);
nor U362 (N_362,In_2333,In_49);
nand U363 (N_363,In_1500,In_1130);
and U364 (N_364,In_3246,In_1075);
or U365 (N_365,In_2028,In_2939);
and U366 (N_366,In_2337,In_2586);
nor U367 (N_367,In_2937,In_1395);
or U368 (N_368,In_4827,In_1265);
or U369 (N_369,In_4204,In_566);
or U370 (N_370,In_1496,In_3175);
nand U371 (N_371,In_3157,In_2840);
and U372 (N_372,In_4237,In_604);
and U373 (N_373,In_2867,In_4152);
nand U374 (N_374,In_1974,In_439);
xnor U375 (N_375,In_2407,In_4022);
xor U376 (N_376,In_1953,In_993);
and U377 (N_377,In_3308,In_1364);
or U378 (N_378,In_372,In_3278);
nor U379 (N_379,In_550,In_2469);
or U380 (N_380,In_2197,In_2981);
or U381 (N_381,In_4712,In_1433);
or U382 (N_382,In_597,In_3208);
nor U383 (N_383,In_2915,In_3564);
and U384 (N_384,In_1674,In_63);
or U385 (N_385,In_3884,In_308);
and U386 (N_386,In_1466,In_3703);
and U387 (N_387,In_1782,In_4696);
and U388 (N_388,In_1343,In_3896);
xnor U389 (N_389,In_735,In_2830);
nor U390 (N_390,In_4191,In_82);
nand U391 (N_391,In_3306,In_2657);
or U392 (N_392,In_376,In_494);
or U393 (N_393,In_1682,In_3386);
nor U394 (N_394,In_1892,In_1997);
nor U395 (N_395,In_3273,In_3166);
or U396 (N_396,In_1404,In_4614);
nor U397 (N_397,In_4693,In_4201);
or U398 (N_398,In_3152,In_390);
nand U399 (N_399,In_3038,In_1198);
xor U400 (N_400,In_1412,In_1313);
nand U401 (N_401,In_42,In_1950);
and U402 (N_402,In_2706,In_1811);
nand U403 (N_403,In_1370,In_1887);
or U404 (N_404,In_3477,In_2271);
or U405 (N_405,In_4789,In_96);
nand U406 (N_406,In_1633,In_4437);
or U407 (N_407,In_329,In_2439);
nand U408 (N_408,In_2819,In_1110);
and U409 (N_409,In_3839,In_420);
and U410 (N_410,In_1780,In_832);
nor U411 (N_411,In_233,In_4078);
or U412 (N_412,In_355,In_4245);
and U413 (N_413,In_503,In_1882);
or U414 (N_414,In_115,In_4900);
xnor U415 (N_415,In_1529,In_2431);
or U416 (N_416,In_2719,In_122);
nor U417 (N_417,In_2643,In_2705);
and U418 (N_418,In_1073,In_838);
and U419 (N_419,In_2774,In_1761);
or U420 (N_420,In_4264,In_2853);
nor U421 (N_421,In_1989,In_3284);
nand U422 (N_422,In_2442,In_131);
nand U423 (N_423,In_4107,In_1234);
nor U424 (N_424,In_3165,In_3772);
nor U425 (N_425,In_272,In_3343);
and U426 (N_426,In_2148,In_1955);
or U427 (N_427,In_2095,In_456);
or U428 (N_428,In_147,In_1610);
and U429 (N_429,In_489,In_570);
or U430 (N_430,In_1101,In_4356);
and U431 (N_431,In_4311,In_677);
nand U432 (N_432,In_3738,In_4369);
nand U433 (N_433,In_2400,In_4119);
or U434 (N_434,In_1085,In_884);
and U435 (N_435,In_567,In_4383);
nand U436 (N_436,In_670,In_2603);
nand U437 (N_437,In_4992,In_2240);
nand U438 (N_438,In_4084,In_3321);
nor U439 (N_439,In_2396,In_4718);
xnor U440 (N_440,In_4451,In_399);
nand U441 (N_441,In_970,In_2785);
xnor U442 (N_442,In_2951,In_444);
or U443 (N_443,In_3504,In_3101);
or U444 (N_444,In_4669,In_626);
and U445 (N_445,In_1802,In_2532);
nor U446 (N_446,In_3806,In_1183);
and U447 (N_447,In_1576,In_2384);
or U448 (N_448,In_4056,In_1308);
nand U449 (N_449,In_831,In_856);
xnor U450 (N_450,In_2859,In_3995);
nor U451 (N_451,In_2851,In_2714);
nand U452 (N_452,In_2403,In_4845);
nand U453 (N_453,In_2846,In_727);
nand U454 (N_454,In_4467,In_892);
nand U455 (N_455,In_2505,In_1476);
or U456 (N_456,In_2044,In_301);
and U457 (N_457,In_3132,In_3868);
xnor U458 (N_458,In_3954,In_1207);
nand U459 (N_459,In_542,In_1);
nand U460 (N_460,In_590,In_130);
nor U461 (N_461,In_3356,In_3519);
xor U462 (N_462,In_2489,In_556);
xor U463 (N_463,In_4177,In_3430);
nand U464 (N_464,In_3238,In_229);
or U465 (N_465,In_1579,In_473);
nand U466 (N_466,In_2330,In_4880);
nand U467 (N_467,In_1286,In_145);
nor U468 (N_468,In_1327,In_2663);
xor U469 (N_469,In_25,In_2443);
xnor U470 (N_470,In_2214,In_1543);
nor U471 (N_471,In_1931,In_1646);
or U472 (N_472,In_326,In_3232);
or U473 (N_473,In_1580,In_4407);
nand U474 (N_474,In_3310,In_3875);
and U475 (N_475,In_1452,In_78);
and U476 (N_476,In_2146,In_3088);
or U477 (N_477,In_1553,In_2256);
or U478 (N_478,In_152,In_4016);
nand U479 (N_479,In_1082,In_2080);
nand U480 (N_480,In_2924,In_1631);
or U481 (N_481,In_2624,In_267);
nor U482 (N_482,In_4314,In_3072);
or U483 (N_483,In_1836,In_1795);
or U484 (N_484,In_4230,In_3737);
and U485 (N_485,In_3001,In_3835);
and U486 (N_486,In_875,In_529);
or U487 (N_487,In_3759,In_2143);
nor U488 (N_488,In_393,In_3501);
and U489 (N_489,In_1104,In_1328);
or U490 (N_490,In_2782,In_3851);
nor U491 (N_491,In_3927,In_4829);
nand U492 (N_492,In_1667,In_787);
nor U493 (N_493,In_2528,In_4797);
and U494 (N_494,In_3946,In_1539);
nand U495 (N_495,In_61,In_26);
nand U496 (N_496,In_4724,In_495);
or U497 (N_497,In_3158,In_4673);
nand U498 (N_498,In_1607,In_4536);
nand U499 (N_499,In_4601,In_771);
and U500 (N_500,In_1925,In_3515);
nor U501 (N_501,In_1463,In_4037);
nor U502 (N_502,In_1139,In_990);
or U503 (N_503,In_2602,In_2126);
nor U504 (N_504,In_1502,In_3909);
nor U505 (N_505,In_2894,In_2429);
nand U506 (N_506,In_2310,In_4917);
or U507 (N_507,In_3776,In_68);
or U508 (N_508,In_4121,In_1190);
nand U509 (N_509,In_4233,In_4633);
and U510 (N_510,In_4001,In_3406);
nand U511 (N_511,In_1681,In_3554);
and U512 (N_512,In_654,In_674);
nor U513 (N_513,In_721,In_3244);
xor U514 (N_514,In_2722,In_3258);
and U515 (N_515,In_4503,In_3722);
and U516 (N_516,In_2005,In_4471);
xnor U517 (N_517,In_3611,In_4360);
and U518 (N_518,In_2038,In_4104);
nor U519 (N_519,In_2917,In_562);
nand U520 (N_520,In_2022,In_103);
nand U521 (N_521,In_3675,In_2856);
nand U522 (N_522,In_211,In_2780);
nand U523 (N_523,In_692,In_883);
nor U524 (N_524,In_4183,In_3449);
or U525 (N_525,In_3074,In_1647);
or U526 (N_526,In_1509,In_4528);
nand U527 (N_527,In_125,In_3643);
xor U528 (N_528,In_1753,In_4462);
and U529 (N_529,In_4582,In_4566);
nand U530 (N_530,In_3736,In_518);
nand U531 (N_531,In_179,In_1969);
nand U532 (N_532,In_2178,In_3904);
nor U533 (N_533,In_3561,In_1919);
nand U534 (N_534,In_3056,In_1393);
or U535 (N_535,In_1058,In_2965);
or U536 (N_536,In_2500,In_2327);
nor U537 (N_537,In_2762,In_4275);
or U538 (N_538,In_477,In_852);
nor U539 (N_539,In_281,In_2236);
nor U540 (N_540,In_593,In_2648);
xor U541 (N_541,In_1334,In_3588);
and U542 (N_542,In_3431,In_18);
or U543 (N_543,In_4247,In_2210);
or U544 (N_544,In_189,In_3220);
nor U545 (N_545,In_3639,In_4456);
and U546 (N_546,In_3992,In_3229);
and U547 (N_547,In_3298,In_1962);
xnor U548 (N_548,In_686,In_1410);
nand U549 (N_549,In_1922,In_1602);
and U550 (N_550,In_4843,In_3231);
nor U551 (N_551,In_302,In_3000);
nor U552 (N_552,In_1293,In_931);
nand U553 (N_553,In_4335,In_3592);
nor U554 (N_554,In_2942,In_1977);
or U555 (N_555,In_3027,In_4446);
xnor U556 (N_556,In_2078,In_2559);
nand U557 (N_557,In_1627,In_4132);
nor U558 (N_558,In_2331,In_808);
nand U559 (N_559,In_1439,In_108);
and U560 (N_560,In_4804,In_1823);
and U561 (N_561,In_2869,In_4215);
and U562 (N_562,In_4111,In_4046);
nor U563 (N_563,In_3586,In_4650);
or U564 (N_564,In_684,In_2376);
nor U565 (N_565,In_509,In_1298);
and U566 (N_566,In_1586,In_1522);
nand U567 (N_567,In_2712,In_2635);
nor U568 (N_568,In_3934,In_635);
nor U569 (N_569,In_3621,In_3161);
and U570 (N_570,In_4608,In_3828);
xor U571 (N_571,In_2905,In_3413);
or U572 (N_572,In_3234,In_3345);
nor U573 (N_573,In_3969,In_3307);
or U574 (N_574,In_675,In_2097);
and U575 (N_575,In_1555,In_3439);
or U576 (N_576,In_1813,In_649);
nor U577 (N_577,In_208,In_4606);
nand U578 (N_578,In_764,In_4085);
and U579 (N_579,In_4216,In_1855);
xnor U580 (N_580,In_2115,In_2119);
or U581 (N_581,In_2166,In_2490);
nor U582 (N_582,In_3911,In_1794);
or U583 (N_583,In_676,In_2084);
and U584 (N_584,In_2906,In_2650);
nand U585 (N_585,In_4420,In_3542);
xor U586 (N_586,In_1380,In_3060);
nand U587 (N_587,In_3571,In_2717);
nand U588 (N_588,In_755,In_3017);
nor U589 (N_589,In_615,In_3395);
and U590 (N_590,In_4524,In_2833);
nand U591 (N_591,In_4716,In_1514);
and U592 (N_592,In_1982,In_56);
and U593 (N_593,In_4522,In_2515);
xnor U594 (N_594,In_1200,In_2926);
or U595 (N_595,In_257,In_2177);
and U596 (N_596,In_2632,In_2480);
xor U597 (N_597,In_1356,In_2441);
and U598 (N_598,In_1083,In_4895);
and U599 (N_599,In_3334,In_3631);
nand U600 (N_600,In_4726,In_3979);
nor U601 (N_601,In_950,In_2172);
xnor U602 (N_602,In_2877,In_4219);
or U603 (N_603,In_3974,In_3065);
and U604 (N_604,In_4021,In_4624);
or U605 (N_605,In_1129,In_2646);
and U606 (N_606,In_2056,In_585);
nand U607 (N_607,In_3615,In_488);
nor U608 (N_608,In_110,In_2213);
nand U609 (N_609,In_1081,In_1728);
and U610 (N_610,In_977,In_1319);
nand U611 (N_611,In_696,In_4539);
or U612 (N_612,In_3907,In_2580);
and U613 (N_613,In_1005,In_2584);
nor U614 (N_614,In_1821,In_1634);
nand U615 (N_615,In_910,In_306);
or U616 (N_616,In_3685,In_1020);
or U617 (N_617,In_3381,In_1284);
and U618 (N_618,In_4165,In_3617);
nand U619 (N_619,In_2522,In_457);
xnor U620 (N_620,In_287,In_259);
or U621 (N_621,In_1077,In_586);
or U622 (N_622,In_3115,In_4562);
nand U623 (N_623,In_3566,In_4153);
or U624 (N_624,In_849,In_3396);
or U625 (N_625,In_2220,In_2768);
or U626 (N_626,In_384,In_2556);
nor U627 (N_627,In_3192,In_2755);
nand U628 (N_628,In_722,In_653);
nor U629 (N_629,In_4143,In_843);
or U630 (N_630,In_2217,In_4209);
nor U631 (N_631,In_3644,In_668);
nand U632 (N_632,In_1548,In_978);
nand U633 (N_633,In_2735,In_3779);
nand U634 (N_634,In_4925,In_3716);
and U635 (N_635,In_1362,In_138);
or U636 (N_636,In_4591,In_3751);
nand U637 (N_637,In_3136,In_2908);
nand U638 (N_638,In_1731,In_2982);
nor U639 (N_639,In_2693,In_3276);
and U640 (N_640,In_3372,In_3533);
nand U641 (N_641,In_3540,In_667);
and U642 (N_642,In_2325,In_1722);
nor U643 (N_643,In_3186,In_2190);
nand U644 (N_644,In_3235,In_3071);
and U645 (N_645,In_2687,In_1860);
nor U646 (N_646,In_4956,In_4554);
or U647 (N_647,In_293,In_4815);
or U648 (N_648,In_3930,In_1167);
nand U649 (N_649,In_2279,In_4980);
or U650 (N_650,In_313,In_3895);
nor U651 (N_651,In_4623,In_2465);
or U652 (N_652,In_411,In_4891);
and U653 (N_653,In_1148,In_3119);
or U654 (N_654,In_574,In_3785);
or U655 (N_655,In_1069,In_1545);
and U656 (N_656,In_563,In_172);
nor U657 (N_657,In_2404,In_4565);
nor U658 (N_658,In_4346,In_594);
and U659 (N_659,In_2120,In_4512);
nand U660 (N_660,In_4478,In_117);
nor U661 (N_661,In_3479,In_4276);
or U662 (N_662,In_4445,In_2614);
and U663 (N_663,In_1559,In_4357);
nand U664 (N_664,In_3709,In_2673);
nand U665 (N_665,In_4881,In_961);
nand U666 (N_666,In_1512,In_4518);
and U667 (N_667,In_2233,In_255);
nand U668 (N_668,In_3581,In_855);
and U669 (N_669,In_1684,In_2452);
or U670 (N_670,In_3666,In_4440);
or U671 (N_671,In_1461,In_2339);
or U672 (N_672,In_1639,In_3786);
nand U673 (N_673,In_1869,In_4596);
xnor U674 (N_674,In_294,In_3980);
nor U675 (N_675,In_3332,In_895);
or U676 (N_676,In_2692,In_2171);
and U677 (N_677,In_2608,In_785);
nor U678 (N_678,In_4738,In_4563);
and U679 (N_679,In_4469,In_3078);
nor U680 (N_680,In_3913,In_35);
and U681 (N_681,In_4665,In_3102);
nand U682 (N_682,In_798,In_368);
nand U683 (N_683,In_2125,In_3991);
or U684 (N_684,In_4619,In_3899);
nand U685 (N_685,In_206,In_2679);
or U686 (N_686,In_70,In_4162);
nor U687 (N_687,In_1636,In_1123);
nor U688 (N_688,In_2681,In_2251);
xnor U689 (N_689,In_4286,In_2764);
and U690 (N_690,In_27,In_3750);
and U691 (N_691,In_223,In_4382);
nand U692 (N_692,In_4841,In_4294);
or U693 (N_693,In_2460,In_1133);
xnor U694 (N_694,In_836,In_271);
nand U695 (N_695,In_3063,In_522);
nor U696 (N_696,In_1716,In_2286);
and U697 (N_697,In_3572,In_3646);
or U698 (N_698,In_2285,In_1001);
and U699 (N_699,In_784,In_664);
nand U700 (N_700,In_4801,In_525);
xnor U701 (N_701,In_4773,In_3171);
nand U702 (N_702,In_2549,In_4805);
nand U703 (N_703,In_1357,In_1617);
nor U704 (N_704,In_3442,In_4885);
nand U705 (N_705,In_4074,In_4695);
and U706 (N_706,In_1443,In_1268);
nor U707 (N_707,In_359,In_751);
or U708 (N_708,In_3176,In_1884);
nand U709 (N_709,In_2502,In_1759);
or U710 (N_710,In_2223,In_4533);
nand U711 (N_711,In_3049,In_2440);
nand U712 (N_712,In_1832,In_4081);
nand U713 (N_713,In_3550,In_2758);
and U714 (N_714,In_1948,In_502);
nand U715 (N_715,In_3309,In_4987);
or U716 (N_716,In_2021,In_421);
and U717 (N_717,In_3694,In_4680);
nand U718 (N_718,In_592,In_901);
nand U719 (N_719,In_409,In_1567);
nor U720 (N_720,In_907,In_3975);
nand U721 (N_721,In_1923,In_2868);
nand U722 (N_722,In_3022,In_1006);
nand U723 (N_723,In_607,In_4535);
nor U724 (N_724,In_1347,In_1583);
nor U725 (N_725,In_1034,In_3444);
and U726 (N_726,In_1295,In_2633);
nand U727 (N_727,In_219,In_3451);
nand U728 (N_728,In_4803,In_3816);
nand U729 (N_729,In_2373,In_4934);
xnor U730 (N_730,In_3368,In_3058);
nor U731 (N_731,In_289,In_2071);
nand U732 (N_732,In_436,In_446);
nor U733 (N_733,In_552,In_1973);
and U734 (N_734,In_3224,In_2389);
nor U735 (N_735,In_2655,In_282);
nand U736 (N_736,In_1978,In_2520);
or U737 (N_737,In_94,In_4927);
and U738 (N_738,In_74,In_3023);
or U739 (N_739,In_4995,In_2328);
nand U740 (N_740,In_2861,In_4299);
nor U741 (N_741,In_3010,In_1483);
and U742 (N_742,In_4459,In_3624);
nand U743 (N_743,In_2383,In_2032);
nand U744 (N_744,In_1100,In_2623);
and U745 (N_745,In_538,In_3424);
and U746 (N_746,In_603,In_1247);
or U747 (N_747,In_1714,In_1774);
or U748 (N_748,In_4397,In_1382);
or U749 (N_749,In_1863,In_4792);
or U750 (N_750,In_4268,In_4960);
nand U751 (N_751,In_3950,In_1879);
and U752 (N_752,In_4938,In_1523);
nor U753 (N_753,In_2723,In_4666);
and U754 (N_754,In_3141,In_2471);
nor U755 (N_755,In_4225,In_4971);
nand U756 (N_756,In_3496,In_2609);
and U757 (N_757,In_1344,In_2893);
or U758 (N_758,In_3362,In_97);
nand U759 (N_759,In_303,In_1505);
or U760 (N_760,In_640,In_3062);
and U761 (N_761,In_2361,In_4061);
nand U762 (N_762,In_4603,In_2020);
nor U763 (N_763,In_4100,In_2769);
nor U764 (N_764,In_23,In_3723);
or U765 (N_765,In_2250,In_1442);
nand U766 (N_766,In_3574,In_2476);
xor U767 (N_767,In_1531,In_2734);
or U768 (N_768,In_4151,In_929);
or U769 (N_769,In_924,In_3124);
xor U770 (N_770,In_718,In_3792);
xnor U771 (N_771,In_1157,In_767);
nor U772 (N_772,In_1669,In_1930);
nand U773 (N_773,In_1280,In_3417);
nand U774 (N_774,In_4387,In_1424);
or U775 (N_775,In_2694,In_1622);
and U776 (N_776,In_2826,In_4854);
nor U777 (N_777,In_1388,In_2461);
and U778 (N_778,In_2752,In_3122);
nor U779 (N_779,In_4968,In_2353);
xnor U780 (N_780,In_3019,In_4943);
or U781 (N_781,In_1611,In_3374);
nand U782 (N_782,In_3985,In_2747);
and U783 (N_783,In_212,In_1993);
or U784 (N_784,In_1801,In_4873);
nor U785 (N_785,In_3589,In_1398);
and U786 (N_786,In_4322,In_241);
xnor U787 (N_787,In_1185,In_1427);
or U788 (N_788,In_2922,In_319);
xor U789 (N_789,In_167,In_3050);
nand U790 (N_790,In_3414,In_2409);
or U791 (N_791,In_898,In_3551);
xor U792 (N_792,In_3303,In_2950);
nand U793 (N_793,In_3590,In_1546);
or U794 (N_794,In_320,In_510);
and U795 (N_795,In_4023,In_3652);
nor U796 (N_796,In_3742,In_1914);
or U797 (N_797,In_4192,In_2149);
or U798 (N_798,In_3300,In_2292);
xor U799 (N_799,In_2929,In_3767);
and U800 (N_800,In_2904,In_2727);
or U801 (N_801,In_4681,In_4972);
and U802 (N_802,In_1834,In_3164);
or U803 (N_803,In_4265,In_4210);
nor U804 (N_804,In_479,In_392);
nand U805 (N_805,In_4865,In_4730);
nand U806 (N_806,In_3834,In_4714);
nand U807 (N_807,In_3850,In_4682);
nand U808 (N_808,In_1871,In_1561);
or U809 (N_809,In_3582,In_1346);
nor U810 (N_810,In_2181,In_1517);
or U811 (N_811,In_191,In_4238);
nand U812 (N_812,In_736,In_1605);
or U813 (N_813,In_3447,In_4054);
and U814 (N_814,In_1222,In_2850);
nand U815 (N_815,In_3784,In_325);
or U816 (N_816,In_351,In_3924);
and U817 (N_817,In_4057,In_459);
nor U818 (N_818,In_4932,In_2317);
nand U819 (N_819,In_2718,In_2923);
nand U820 (N_820,In_2195,In_3813);
nor U821 (N_821,In_3156,In_4366);
nand U822 (N_822,In_960,In_3926);
nor U823 (N_823,In_4783,In_4771);
nor U824 (N_824,In_3790,In_4436);
nand U825 (N_825,In_4169,In_1169);
nand U826 (N_826,In_3082,In_3848);
nand U827 (N_827,In_3888,In_2043);
or U828 (N_828,In_539,In_4757);
and U829 (N_829,In_2479,In_3843);
nand U830 (N_830,In_1480,In_766);
nor U831 (N_831,In_4491,In_73);
or U832 (N_832,In_4018,In_1643);
nor U833 (N_833,In_4684,In_3446);
or U834 (N_834,In_2649,In_1397);
nand U835 (N_835,In_4755,In_3538);
nor U836 (N_836,In_2636,In_362);
and U837 (N_837,In_4043,In_2130);
nand U838 (N_838,In_669,In_285);
and U839 (N_839,In_2919,In_4574);
nand U840 (N_840,In_3502,In_2540);
xor U841 (N_841,In_879,In_1336);
or U842 (N_842,In_622,In_3094);
nor U843 (N_843,In_744,In_276);
xnor U844 (N_844,In_2059,In_2364);
nor U845 (N_845,In_3729,In_3885);
nand U846 (N_846,In_1551,In_1224);
or U847 (N_847,In_4235,In_1785);
or U848 (N_848,In_3734,In_2221);
or U849 (N_849,In_127,In_197);
xnor U850 (N_850,In_4945,In_4371);
xor U851 (N_851,In_2259,In_4683);
xor U852 (N_852,In_2139,In_3728);
nand U853 (N_853,In_3730,In_2147);
nor U854 (N_854,In_2219,In_4398);
nor U855 (N_855,In_1365,In_1140);
nor U856 (N_856,In_2641,In_4587);
or U857 (N_857,In_279,In_1031);
xor U858 (N_858,In_2824,In_660);
nor U859 (N_859,In_370,In_3775);
or U860 (N_860,In_1575,In_327);
nand U861 (N_861,In_1493,In_1338);
xnor U862 (N_862,In_4542,In_50);
or U863 (N_863,In_3583,In_16);
and U864 (N_864,In_3401,In_844);
and U865 (N_865,In_979,In_1573);
or U866 (N_866,In_2416,In_1768);
nor U867 (N_867,In_236,In_1668);
or U868 (N_868,In_629,In_398);
and U869 (N_869,In_2552,In_2072);
or U870 (N_870,In_703,In_3200);
and U871 (N_871,In_4567,In_905);
nand U872 (N_872,In_1099,In_1238);
xnor U873 (N_873,In_3739,In_4030);
or U874 (N_874,In_4853,In_1459);
and U875 (N_875,In_2618,In_2011);
nor U876 (N_876,In_2589,In_2314);
and U877 (N_877,In_3573,In_3002);
nand U878 (N_878,In_1784,In_602);
nor U879 (N_879,In_4414,In_1886);
and U880 (N_880,In_1482,In_2959);
nand U881 (N_881,In_4310,In_3798);
nor U882 (N_882,In_725,In_102);
xnor U883 (N_883,In_4020,In_3879);
nor U884 (N_884,In_1911,In_383);
or U885 (N_885,In_4188,In_129);
or U886 (N_886,In_4708,In_269);
nor U887 (N_887,In_80,In_2415);
and U888 (N_888,In_2352,In_3741);
nand U889 (N_889,In_4808,In_4847);
or U890 (N_890,In_4551,In_343);
or U891 (N_891,In_433,In_4146);
or U892 (N_892,In_1477,In_528);
nand U893 (N_893,In_2459,In_1525);
and U894 (N_894,In_2617,In_3055);
and U895 (N_895,In_774,In_2063);
and U896 (N_896,In_4913,In_1940);
xnor U897 (N_897,In_2665,In_3971);
or U898 (N_898,In_3127,In_4347);
nand U899 (N_899,In_3256,In_1127);
xor U900 (N_900,In_4203,In_4448);
nor U901 (N_901,In_1120,In_2647);
and U902 (N_902,In_2878,In_4628);
or U903 (N_903,In_4864,In_3789);
nand U904 (N_904,In_2299,In_464);
nand U905 (N_905,In_1783,In_2222);
or U906 (N_906,In_955,In_4434);
nand U907 (N_907,In_968,In_1422);
or U908 (N_908,In_2173,In_1411);
xor U909 (N_909,In_1859,In_792);
nor U910 (N_910,In_519,In_4140);
and U911 (N_911,In_4431,In_280);
nor U912 (N_912,In_3322,In_4849);
nor U913 (N_913,In_2897,In_1359);
nor U914 (N_914,In_3388,In_4234);
and U915 (N_915,In_3944,In_4433);
and U916 (N_916,In_4079,In_3883);
or U917 (N_917,In_4484,In_3422);
nand U918 (N_918,In_840,In_2823);
nor U919 (N_919,In_1032,In_1051);
and U920 (N_920,In_2876,In_739);
or U921 (N_921,In_2503,In_3111);
nand U922 (N_922,In_783,In_4131);
xnor U923 (N_923,In_3912,In_4821);
or U924 (N_924,In_2799,In_2273);
nand U925 (N_925,In_3272,In_4123);
or U926 (N_926,In_3364,In_405);
nor U927 (N_927,In_1418,In_2307);
nand U928 (N_928,In_3948,In_1675);
nor U929 (N_929,In_4441,In_2426);
or U930 (N_930,In_1163,In_2804);
xor U931 (N_931,In_4135,In_3854);
nand U932 (N_932,In_1924,In_356);
xor U933 (N_933,In_1040,In_2235);
and U934 (N_934,In_1824,In_4810);
nand U935 (N_935,In_1067,In_1445);
nand U936 (N_936,In_2899,In_4363);
nor U937 (N_937,In_1820,In_4819);
xor U938 (N_938,In_1288,In_4134);
nor U939 (N_939,In_3608,In_316);
and U940 (N_940,In_4694,In_36);
or U941 (N_941,In_3257,In_3320);
or U942 (N_942,In_353,In_3657);
nor U943 (N_943,In_1570,In_1998);
nor U944 (N_944,In_857,In_2076);
xnor U945 (N_945,In_1975,In_2474);
nor U946 (N_946,In_3026,In_4728);
and U947 (N_947,In_625,In_2165);
or U948 (N_948,In_1211,In_415);
nor U949 (N_949,In_557,In_1371);
or U950 (N_950,In_863,In_1043);
and U951 (N_951,In_1942,In_192);
nor U952 (N_952,In_2382,In_2338);
and U953 (N_953,In_1376,In_4733);
xnor U954 (N_954,In_3663,In_4071);
or U955 (N_955,In_3938,In_3596);
nand U956 (N_956,In_3487,In_3760);
xor U957 (N_957,In_1375,In_1518);
xor U958 (N_958,In_1242,In_634);
nor U959 (N_959,In_3822,In_1846);
nand U960 (N_960,In_20,In_1556);
nor U961 (N_961,In_1981,In_4661);
nand U962 (N_962,In_1342,In_4922);
nand U963 (N_963,In_151,In_86);
and U964 (N_964,In_3497,In_166);
xor U965 (N_965,In_3720,In_2838);
xor U966 (N_966,In_2141,In_4058);
nand U967 (N_967,In_251,In_3937);
or U968 (N_968,In_644,In_2380);
nor U969 (N_969,In_449,In_709);
nand U970 (N_970,In_3664,In_3443);
nor U971 (N_971,In_3044,In_12);
nor U972 (N_972,In_2242,In_1569);
and U973 (N_973,In_4800,In_806);
nor U974 (N_974,In_3525,In_4156);
nand U975 (N_975,In_1660,In_4218);
nand U976 (N_976,In_1296,In_3569);
or U977 (N_977,In_4970,In_3211);
or U978 (N_978,In_4035,In_812);
and U979 (N_979,In_2627,In_3015);
nand U980 (N_980,In_2558,In_1853);
and U981 (N_981,In_890,In_1434);
and U982 (N_982,In_3159,In_1958);
and U983 (N_983,In_3823,In_601);
nor U984 (N_984,In_4632,In_2091);
and U985 (N_985,In_804,In_1354);
and U986 (N_986,In_1102,In_3841);
and U987 (N_987,In_217,In_1330);
nor U988 (N_988,In_4122,In_2275);
nand U989 (N_989,In_1274,In_1604);
nand U990 (N_990,In_4658,In_321);
or U991 (N_991,In_2659,In_4636);
and U992 (N_992,In_3304,In_2598);
and U993 (N_993,In_1699,In_4045);
nor U994 (N_994,In_296,In_2102);
and U995 (N_995,In_800,In_2684);
nand U996 (N_996,In_1849,In_2969);
nor U997 (N_997,In_4041,In_4736);
nand U998 (N_998,In_2967,In_3602);
or U999 (N_999,In_2902,In_4860);
nor U1000 (N_1000,In_2034,In_1881);
and U1001 (N_1001,In_1150,In_1828);
nand U1002 (N_1002,In_2131,In_46);
or U1003 (N_1003,In_4531,In_3567);
nand U1004 (N_1004,In_911,In_2484);
or U1005 (N_1005,In_3144,In_3295);
or U1006 (N_1006,In_4000,In_2232);
nand U1007 (N_1007,In_1430,In_1349);
nor U1008 (N_1008,In_4408,In_142);
or U1009 (N_1009,In_4176,In_3942);
and U1010 (N_1010,In_4944,In_4272);
and U1011 (N_1011,In_4115,In_646);
or U1012 (N_1012,In_2433,In_3455);
or U1013 (N_1013,In_645,In_712);
xnor U1014 (N_1014,In_4180,In_3064);
or U1015 (N_1015,In_1273,In_3658);
and U1016 (N_1016,In_2776,In_816);
and U1017 (N_1017,In_51,In_4498);
and U1018 (N_1018,In_2550,In_157);
or U1019 (N_1019,In_338,In_862);
nand U1020 (N_1020,In_4395,In_2990);
nor U1021 (N_1021,In_803,In_935);
or U1022 (N_1022,In_4868,In_1745);
or U1023 (N_1023,In_4772,In_2770);
or U1024 (N_1024,In_4555,In_3375);
nor U1025 (N_1025,In_2521,In_765);
or U1026 (N_1026,In_2744,In_2791);
nand U1027 (N_1027,In_1018,In_2492);
or U1028 (N_1028,In_1291,In_3291);
nor U1029 (N_1029,In_3518,In_4003);
or U1030 (N_1030,In_3236,In_1460);
nand U1031 (N_1031,In_1976,In_159);
or U1032 (N_1032,In_2227,In_921);
or U1033 (N_1033,In_4211,In_3367);
xnor U1034 (N_1034,In_3667,In_2507);
nand U1035 (N_1035,In_4502,In_140);
or U1036 (N_1036,In_3625,In_2870);
or U1037 (N_1037,In_4969,In_2326);
nor U1038 (N_1038,In_3138,In_1339);
and U1039 (N_1039,In_2301,In_4050);
or U1040 (N_1040,In_4883,In_1626);
or U1041 (N_1041,In_482,In_1332);
nand U1042 (N_1042,In_339,In_1944);
nand U1043 (N_1043,In_1184,In_3593);
xnor U1044 (N_1044,In_3647,In_468);
nand U1045 (N_1045,In_841,In_3201);
nand U1046 (N_1046,In_1078,In_3194);
and U1047 (N_1047,In_548,In_1990);
nor U1048 (N_1048,In_2255,In_4055);
nor U1049 (N_1049,In_1079,In_1848);
or U1050 (N_1050,In_916,In_1935);
or U1051 (N_1051,In_4034,In_4952);
nor U1052 (N_1052,In_3098,In_1513);
and U1053 (N_1053,In_4470,In_3706);
nor U1054 (N_1054,In_2975,In_2079);
xnor U1055 (N_1055,In_4051,In_3963);
xnor U1056 (N_1056,In_2891,In_2266);
or U1057 (N_1057,In_551,In_350);
or U1058 (N_1058,In_926,In_1350);
or U1059 (N_1059,In_4213,In_4262);
or U1060 (N_1060,In_4690,In_3858);
nand U1061 (N_1061,In_881,In_2316);
and U1062 (N_1062,In_4168,In_2760);
xor U1063 (N_1063,In_3804,In_1593);
nor U1064 (N_1064,In_465,In_4454);
and U1065 (N_1065,In_656,In_1770);
or U1066 (N_1066,In_1454,In_4076);
xnor U1067 (N_1067,In_4325,In_2320);
nor U1068 (N_1068,In_3067,In_2815);
nor U1069 (N_1069,In_1677,In_2527);
nand U1070 (N_1070,In_2472,In_4548);
and U1071 (N_1071,In_4044,In_239);
xnor U1072 (N_1072,In_2012,In_2837);
or U1073 (N_1073,In_2002,In_2977);
nand U1074 (N_1074,In_1947,In_4271);
nand U1075 (N_1075,In_1166,In_1540);
and U1076 (N_1076,In_3869,In_2142);
or U1077 (N_1077,In_4403,In_2546);
nor U1078 (N_1078,In_1090,In_4377);
nand U1079 (N_1079,In_2644,In_1599);
and U1080 (N_1080,In_4597,In_4010);
and U1081 (N_1081,In_4384,In_437);
nand U1082 (N_1082,In_367,In_4160);
and U1083 (N_1083,In_4015,In_1276);
nand U1084 (N_1084,In_3986,In_3030);
or U1085 (N_1085,In_3549,In_1515);
nand U1086 (N_1086,In_47,In_1275);
or U1087 (N_1087,In_4406,In_671);
and U1088 (N_1088,In_4179,In_1949);
or U1089 (N_1089,In_2121,In_4609);
xor U1090 (N_1090,In_4541,In_4466);
or U1091 (N_1091,In_2406,In_1812);
nor U1092 (N_1092,In_3109,In_1927);
and U1093 (N_1093,In_4965,In_918);
nand U1094 (N_1094,In_4698,In_4662);
or U1095 (N_1095,In_4222,In_2616);
and U1096 (N_1096,In_2446,In_2077);
or U1097 (N_1097,In_2280,In_1991);
nor U1098 (N_1098,In_4362,In_160);
nand U1099 (N_1099,In_949,In_1444);
and U1100 (N_1100,In_113,In_2788);
nand U1101 (N_1101,In_188,In_4423);
and U1102 (N_1102,In_2583,In_920);
xor U1103 (N_1103,In_4511,In_1214);
nand U1104 (N_1104,In_3654,In_3346);
or U1105 (N_1105,In_980,In_1503);
nor U1106 (N_1106,In_4096,In_2934);
or U1107 (N_1107,In_747,In_250);
or U1108 (N_1108,In_3910,In_1642);
and U1109 (N_1109,In_4297,In_4333);
and U1110 (N_1110,In_3390,In_1377);
xor U1111 (N_1111,In_3354,In_169);
nand U1112 (N_1112,In_2163,In_4419);
nand U1113 (N_1113,In_3204,In_3978);
or U1114 (N_1114,In_2003,In_4741);
nand U1115 (N_1115,In_2154,In_1724);
nand U1116 (N_1116,In_2392,In_648);
or U1117 (N_1117,In_2388,In_1180);
nor U1118 (N_1118,In_3503,In_253);
xor U1119 (N_1119,In_3614,In_1489);
and U1120 (N_1120,In_2212,In_7);
nor U1121 (N_1121,In_2313,In_1735);
xor U1122 (N_1122,In_4473,In_1883);
or U1123 (N_1123,In_22,In_1387);
and U1124 (N_1124,In_2530,In_1134);
or U1125 (N_1125,In_3488,In_4825);
xor U1126 (N_1126,In_4729,In_3348);
nor U1127 (N_1127,In_4735,In_3665);
nor U1128 (N_1128,In_4878,In_4025);
or U1129 (N_1129,In_1650,In_4480);
or U1130 (N_1130,In_2662,In_1992);
or U1131 (N_1131,In_4206,In_1652);
nand U1132 (N_1132,In_1315,In_1010);
nand U1133 (N_1133,In_4386,In_3584);
nand U1134 (N_1134,In_4640,In_1353);
and U1135 (N_1135,In_1670,In_1449);
nand U1136 (N_1136,In_1049,In_4313);
and U1137 (N_1137,In_3465,In_4572);
nand U1138 (N_1138,In_4510,In_143);
nand U1139 (N_1139,In_358,In_1890);
or U1140 (N_1140,In_336,In_547);
or U1141 (N_1141,In_4507,In_3178);
or U1142 (N_1142,In_4108,In_569);
nand U1143 (N_1143,In_3837,In_4038);
nand U1144 (N_1144,In_1159,In_3241);
and U1145 (N_1145,In_155,In_1406);
and U1146 (N_1146,In_2329,In_3483);
nor U1147 (N_1147,In_1904,In_2612);
or U1148 (N_1148,In_1804,In_3289);
and U1149 (N_1149,In_605,In_1864);
and U1150 (N_1150,In_69,In_423);
nor U1151 (N_1151,In_1653,In_3740);
nor U1152 (N_1152,In_1282,In_1778);
nor U1153 (N_1153,In_2444,In_317);
and U1154 (N_1154,In_3041,In_1564);
xor U1155 (N_1155,In_1378,In_2524);
and U1156 (N_1156,In_829,In_2430);
or U1157 (N_1157,In_121,In_2999);
nand U1158 (N_1158,In_2847,In_332);
nand U1159 (N_1159,In_983,In_1544);
nand U1160 (N_1160,In_3147,In_1693);
nand U1161 (N_1161,In_2007,In_3725);
and U1162 (N_1162,In_438,In_1968);
and U1163 (N_1163,In_434,In_3903);
nor U1164 (N_1164,In_3939,In_4877);
and U1165 (N_1165,In_2370,In_2786);
nand U1166 (N_1166,In_204,In_2835);
and U1167 (N_1167,In_3970,In_1210);
nor U1168 (N_1168,In_2117,In_3277);
xor U1169 (N_1169,In_1664,In_1179);
nand U1170 (N_1170,In_1259,In_2529);
or U1171 (N_1171,In_4790,In_900);
nand U1172 (N_1172,In_1771,In_1227);
nand U1173 (N_1173,In_3428,In_2475);
xnor U1174 (N_1174,In_1945,In_1880);
or U1175 (N_1175,In_2457,In_4985);
or U1176 (N_1176,In_796,In_775);
xnor U1177 (N_1177,In_401,In_1066);
and U1178 (N_1178,In_4200,In_2434);
and U1179 (N_1179,In_3415,In_4385);
or U1180 (N_1180,In_3576,In_3990);
and U1181 (N_1181,In_2993,In_1154);
or U1182 (N_1182,In_4040,In_1659);
xnor U1183 (N_1183,In_714,In_478);
nand U1184 (N_1184,In_4953,In_595);
nor U1185 (N_1185,In_2268,In_1932);
and U1186 (N_1186,In_4318,In_3239);
nand U1187 (N_1187,In_2685,In_3035);
nand U1188 (N_1188,In_1612,In_3274);
nor U1189 (N_1189,In_4779,In_2347);
nand U1190 (N_1190,In_3416,In_3327);
or U1191 (N_1191,In_4752,In_3977);
or U1192 (N_1192,In_4246,In_663);
or U1193 (N_1193,In_1637,In_1748);
and U1194 (N_1194,In_3660,In_4430);
nor U1195 (N_1195,In_2511,In_3747);
and U1196 (N_1196,In_4257,In_2218);
and U1197 (N_1197,In_4997,In_2074);
or U1198 (N_1198,In_1479,In_3849);
or U1199 (N_1199,In_1253,In_4465);
or U1200 (N_1200,In_4584,In_992);
and U1201 (N_1201,In_1562,In_2896);
nor U1202 (N_1202,In_1186,In_925);
and U1203 (N_1203,In_3642,In_1526);
or U1204 (N_1204,In_2864,In_2289);
nand U1205 (N_1205,In_3678,In_4786);
and U1206 (N_1206,In_3766,In_1436);
or U1207 (N_1207,In_3955,In_4186);
nor U1208 (N_1208,In_3468,In_1399);
xor U1209 (N_1209,In_1011,In_4592);
nand U1210 (N_1210,In_1467,In_2374);
and U1211 (N_1211,In_2112,In_1470);
or U1212 (N_1212,In_1462,In_1013);
and U1213 (N_1213,In_951,In_380);
and U1214 (N_1214,In_1277,In_3537);
and U1215 (N_1215,In_1126,In_3036);
nand U1216 (N_1216,In_187,In_1086);
and U1217 (N_1217,In_4091,In_4876);
nand U1218 (N_1218,In_564,In_1045);
nor U1219 (N_1219,In_536,In_1383);
and U1220 (N_1220,In_249,In_54);
or U1221 (N_1221,In_91,In_1755);
or U1222 (N_1222,In_2903,In_4688);
nor U1223 (N_1223,In_749,In_227);
nand U1224 (N_1224,In_2626,In_3462);
nor U1225 (N_1225,In_1690,In_1817);
nand U1226 (N_1226,In_4671,In_2946);
nor U1227 (N_1227,In_3546,In_2187);
nor U1228 (N_1228,In_1144,In_3481);
nand U1229 (N_1229,In_4277,In_3698);
and U1230 (N_1230,In_4838,In_65);
and U1231 (N_1231,In_1861,In_2508);
nor U1232 (N_1232,In_1306,In_3193);
nor U1233 (N_1233,In_2607,In_3380);
or U1234 (N_1234,In_799,In_2300);
or U1235 (N_1235,In_3831,In_2701);
and U1236 (N_1236,In_116,In_957);
or U1237 (N_1237,In_3929,In_850);
and U1238 (N_1238,In_4710,In_1016);
nand U1239 (N_1239,In_1152,In_4319);
and U1240 (N_1240,In_3618,In_2984);
and U1241 (N_1241,In_1806,In_3311);
or U1242 (N_1242,In_4626,In_2174);
or U1243 (N_1243,In_429,In_3486);
nand U1244 (N_1244,In_777,In_3817);
nor U1245 (N_1245,In_2652,In_1289);
nand U1246 (N_1246,In_4617,In_4713);
and U1247 (N_1247,In_4094,In_4080);
and U1248 (N_1248,In_3787,In_965);
nand U1249 (N_1249,In_1711,In_48);
nor U1250 (N_1250,In_1044,In_1125);
nand U1251 (N_1251,In_4101,In_168);
or U1252 (N_1252,In_4557,In_4898);
or U1253 (N_1253,In_4709,In_4068);
nand U1254 (N_1254,In_3243,In_2209);
and U1255 (N_1255,In_2101,In_591);
and U1256 (N_1256,In_3744,In_3524);
xor U1257 (N_1257,In_2150,In_2357);
nor U1258 (N_1258,In_3105,In_1903);
or U1259 (N_1259,In_1438,In_3445);
nor U1260 (N_1260,In_1715,In_2050);
or U1261 (N_1261,In_4958,In_4254);
nand U1262 (N_1262,In_4138,In_1158);
and U1263 (N_1263,In_162,In_1536);
xnor U1264 (N_1264,In_1068,In_1429);
and U1265 (N_1265,In_3006,In_4060);
nand U1266 (N_1266,In_442,In_4167);
and U1267 (N_1267,In_1807,In_1803);
nand U1268 (N_1268,In_3799,In_375);
nand U1269 (N_1269,In_846,In_133);
or U1270 (N_1270,In_261,In_2470);
and U1271 (N_1271,In_2485,In_4178);
and U1272 (N_1272,In_3466,In_2765);
and U1273 (N_1273,In_4580,In_1193);
xor U1274 (N_1274,In_4117,In_33);
or U1275 (N_1275,In_10,In_3107);
or U1276 (N_1276,In_1019,In_3410);
or U1277 (N_1277,In_4692,In_3448);
and U1278 (N_1278,In_2569,In_3506);
nor U1279 (N_1279,In_3764,In_2772);
and U1280 (N_1280,In_2288,In_3941);
or U1281 (N_1281,In_1389,In_3580);
nand U1282 (N_1282,In_2363,In_4870);
nand U1283 (N_1283,In_379,In_4342);
nor U1284 (N_1284,In_652,In_3230);
and U1285 (N_1285,In_4648,In_1379);
nor U1286 (N_1286,In_1294,In_532);
nand U1287 (N_1287,In_3285,In_878);
or U1288 (N_1288,In_4402,In_4349);
or U1289 (N_1289,In_4147,In_4831);
or U1290 (N_1290,In_2008,In_1229);
nor U1291 (N_1291,In_1096,In_642);
nand U1292 (N_1292,In_4722,In_4485);
xnor U1293 (N_1293,In_4781,In_4047);
nand U1294 (N_1294,In_304,In_4495);
and U1295 (N_1295,In_4083,In_1318);
and U1296 (N_1296,In_2754,In_1056);
nand U1297 (N_1297,In_1360,In_2183);
xor U1298 (N_1298,In_2811,In_4370);
nand U1299 (N_1299,In_4645,In_4281);
and U1300 (N_1300,In_4862,In_1898);
and U1301 (N_1301,In_1021,In_2514);
nand U1302 (N_1302,In_3712,In_4266);
nor U1303 (N_1303,In_4391,In_582);
nand U1304 (N_1304,In_2405,In_561);
nor U1305 (N_1305,In_4006,In_3641);
and U1306 (N_1306,In_4421,In_2986);
nor U1307 (N_1307,In_3283,In_4761);
and U1308 (N_1308,In_1899,In_2039);
nand U1309 (N_1309,In_150,In_4544);
and U1310 (N_1310,In_3080,In_3510);
nor U1311 (N_1311,In_135,In_3150);
nand U1312 (N_1312,In_4175,In_2494);
or U1313 (N_1313,In_2239,In_912);
nor U1314 (N_1314,In_410,In_1048);
nor U1315 (N_1315,In_4858,In_1766);
nor U1316 (N_1316,In_454,In_2371);
or U1317 (N_1317,In_263,In_2857);
nand U1318 (N_1318,In_3824,In_2783);
nor U1319 (N_1319,In_453,In_2249);
nand U1320 (N_1320,In_3004,In_1769);
nor U1321 (N_1321,In_3552,In_2909);
nor U1322 (N_1322,In_4239,In_4795);
nand U1323 (N_1323,In_4258,In_3961);
nand U1324 (N_1324,In_4793,In_480);
or U1325 (N_1325,In_3323,In_3782);
nor U1326 (N_1326,In_688,In_4630);
or U1327 (N_1327,In_2944,In_3494);
xor U1328 (N_1328,In_4785,In_655);
nand U1329 (N_1329,In_4907,In_199);
or U1330 (N_1330,In_497,In_4514);
or U1331 (N_1331,In_2281,In_4412);
nand U1332 (N_1332,In_4949,In_4942);
or U1333 (N_1333,In_4486,In_2453);
nand U1334 (N_1334,In_3965,In_3003);
nor U1335 (N_1335,In_1204,In_4558);
or U1336 (N_1336,In_2324,In_4269);
and U1337 (N_1337,In_3352,In_2746);
or U1338 (N_1338,In_4703,In_3212);
nand U1339 (N_1339,In_794,In_1035);
nor U1340 (N_1340,In_876,In_4114);
nand U1341 (N_1341,In_934,In_2901);
nand U1342 (N_1342,In_3650,In_4595);
or U1343 (N_1343,In_1114,In_1322);
or U1344 (N_1344,In_3653,In_435);
nand U1345 (N_1345,In_1877,In_4753);
or U1346 (N_1346,In_1941,In_2880);
and U1347 (N_1347,In_1143,In_4705);
nand U1348 (N_1348,In_839,In_163);
nor U1349 (N_1349,In_820,In_2761);
nor U1350 (N_1350,In_797,In_348);
and U1351 (N_1351,In_967,In_575);
or U1352 (N_1352,In_2194,In_2284);
nor U1353 (N_1353,In_1961,In_2998);
nor U1354 (N_1354,In_1980,In_471);
nor U1355 (N_1355,In_1414,In_3844);
nand U1356 (N_1356,In_4093,In_4493);
xor U1357 (N_1357,In_470,In_1494);
or U1358 (N_1358,In_3604,In_3595);
nor U1359 (N_1359,In_2987,In_71);
nand U1360 (N_1360,In_2613,In_4479);
or U1361 (N_1361,In_4823,In_193);
or U1362 (N_1362,In_1852,In_1595);
or U1363 (N_1363,In_1581,In_3427);
nor U1364 (N_1364,In_2144,In_2778);
and U1365 (N_1365,In_226,In_617);
and U1366 (N_1366,In_3801,In_2832);
nor U1367 (N_1367,In_0,In_3997);
nand U1368 (N_1368,In_3459,In_4802);
and U1369 (N_1369,In_2745,In_710);
and U1370 (N_1370,In_3715,In_156);
or U1371 (N_1371,In_1516,In_3172);
or U1372 (N_1372,In_283,In_3139);
and U1373 (N_1373,In_2017,In_3563);
nor U1374 (N_1374,In_3690,In_717);
and U1375 (N_1375,In_228,In_3275);
xor U1376 (N_1376,In_3037,In_4026);
nor U1377 (N_1377,In_4064,In_3480);
nor U1378 (N_1378,In_2971,In_3964);
or U1379 (N_1379,In_2451,In_149);
xnor U1380 (N_1380,In_183,In_4157);
nor U1381 (N_1381,In_492,In_3471);
and U1382 (N_1382,In_3371,In_136);
and U1383 (N_1383,In_2845,In_2188);
nor U1384 (N_1384,In_3967,In_2566);
and U1385 (N_1385,In_3981,In_4288);
nand U1386 (N_1386,In_4128,In_1936);
and U1387 (N_1387,In_2100,In_2182);
and U1388 (N_1388,In_310,In_4964);
xor U1389 (N_1389,In_3893,In_3126);
and U1390 (N_1390,In_3250,In_2061);
xor U1391 (N_1391,In_3881,In_1885);
or U1392 (N_1392,In_2773,In_4303);
and U1393 (N_1393,In_2211,In_2336);
nand U1394 (N_1394,In_3337,In_4053);
and U1395 (N_1395,In_4243,In_4348);
nand U1396 (N_1396,In_3473,In_394);
nand U1397 (N_1397,In_1741,In_3227);
nor U1398 (N_1398,In_1235,In_4130);
and U1399 (N_1399,In_1300,In_1417);
and U1400 (N_1400,In_1839,In_1425);
nor U1401 (N_1401,In_4404,In_1033);
or U1402 (N_1402,In_4401,In_4373);
and U1403 (N_1403,In_1830,In_1323);
xor U1404 (N_1404,In_1028,In_4400);
nand U1405 (N_1405,In_1223,In_1199);
nand U1406 (N_1406,In_483,In_2702);
or U1407 (N_1407,In_2816,In_3418);
nand U1408 (N_1408,In_1251,In_1499);
nand U1409 (N_1409,In_2708,In_1615);
and U1410 (N_1410,In_1878,In_4350);
or U1411 (N_1411,In_2342,In_3770);
nand U1412 (N_1412,In_4181,In_1938);
nand U1413 (N_1413,In_2976,In_1845);
or U1414 (N_1414,In_1022,In_1606);
or U1415 (N_1415,In_3475,In_1269);
nand U1416 (N_1416,In_3160,In_2463);
or U1417 (N_1417,In_295,In_4822);
and U1418 (N_1418,In_1857,In_1751);
and U1419 (N_1419,In_1189,In_3531);
nor U1420 (N_1420,In_1638,In_5);
nor U1421 (N_1421,In_4700,In_1616);
or U1422 (N_1422,In_1687,In_4884);
and U1423 (N_1423,In_3271,In_535);
and U1424 (N_1424,In_3735,In_4644);
nand U1425 (N_1425,In_154,In_3721);
nand U1426 (N_1426,In_752,In_3918);
xnor U1427 (N_1427,In_2496,In_2035);
or U1428 (N_1428,In_3557,In_4765);
and U1429 (N_1429,In_3695,In_880);
and U1430 (N_1430,In_4499,In_1151);
or U1431 (N_1431,In_1122,In_400);
and U1432 (N_1432,In_2027,In_4283);
nand U1433 (N_1433,In_526,In_3509);
and U1434 (N_1434,In_1723,In_4291);
and U1435 (N_1435,In_1218,In_4125);
or U1436 (N_1436,In_385,In_1721);
or U1437 (N_1437,In_2625,In_2104);
nor U1438 (N_1438,In_1390,In_4679);
nor U1439 (N_1439,In_2928,In_1405);
nand U1440 (N_1440,In_1729,In_4453);
xor U1441 (N_1441,In_1391,In_4559);
or U1442 (N_1442,In_2047,In_2158);
nand U1443 (N_1443,In_4894,In_3532);
nor U1444 (N_1444,In_1272,In_2167);
nor U1445 (N_1445,In_1578,In_1805);
or U1446 (N_1446,In_2246,In_4488);
nor U1447 (N_1447,In_861,In_2046);
and U1448 (N_1448,In_4439,In_4828);
xor U1449 (N_1449,In_939,In_2004);
and U1450 (N_1450,In_201,In_3651);
nor U1451 (N_1451,In_2355,In_1552);
nor U1452 (N_1452,In_589,In_1565);
nand U1453 (N_1453,In_3420,In_4145);
or U1454 (N_1454,In_3800,In_886);
xor U1455 (N_1455,In_2069,In_691);
nor U1456 (N_1456,In_4748,In_943);
nand U1457 (N_1457,In_4545,In_1838);
and U1458 (N_1458,In_971,In_3069);
nand U1459 (N_1459,In_3325,In_3155);
nor U1460 (N_1460,In_4339,In_1894);
or U1461 (N_1461,In_4009,In_4749);
and U1462 (N_1462,In_609,In_2151);
nand U1463 (N_1463,In_2680,In_2193);
xor U1464 (N_1464,In_3316,In_4948);
or U1465 (N_1465,In_2348,In_2138);
and U1466 (N_1466,In_1742,In_3810);
nand U1467 (N_1467,In_1239,In_2170);
xnor U1468 (N_1468,In_530,In_1366);
and U1469 (N_1469,In_1874,In_689);
nor U1470 (N_1470,In_1900,In_499);
nor U1471 (N_1471,In_730,In_4782);
or U1472 (N_1472,In_2592,In_4532);
nand U1473 (N_1473,In_4926,In_2018);
or U1474 (N_1474,In_2340,In_4012);
nand U1475 (N_1475,In_3645,In_3042);
and U1476 (N_1476,In_3699,In_4527);
or U1477 (N_1477,In_3114,In_3225);
or U1478 (N_1478,In_3976,In_2185);
and U1479 (N_1479,In_1822,In_4678);
nor U1480 (N_1480,In_34,In_360);
and U1481 (N_1481,In_361,In_3680);
or U1482 (N_1482,In_568,In_762);
nand U1483 (N_1483,In_4504,In_268);
or U1484 (N_1484,In_2629,In_2160);
nand U1485 (N_1485,In_3575,In_2661);
nor U1486 (N_1486,In_3606,In_673);
nor U1487 (N_1487,In_284,In_2557);
nor U1488 (N_1488,In_3543,In_3457);
or U1489 (N_1489,In_2481,In_4144);
xnor U1490 (N_1490,In_4540,In_4489);
or U1491 (N_1491,In_3866,In_2114);
and U1492 (N_1492,In_2730,In_2895);
and U1493 (N_1493,In_888,In_763);
or U1494 (N_1494,In_498,In_4240);
nand U1495 (N_1495,In_2096,In_2567);
or U1496 (N_1496,In_2852,In_3923);
nand U1497 (N_1497,In_3409,In_3084);
nor U1498 (N_1498,In_2561,In_1408);
nand U1499 (N_1499,In_3919,In_1147);
nor U1500 (N_1500,In_1549,In_827);
and U1501 (N_1501,In_8,In_59);
or U1502 (N_1502,In_3290,In_810);
nand U1503 (N_1503,In_1426,In_4163);
nor U1504 (N_1504,In_2601,In_3659);
nor U1505 (N_1505,In_3209,In_146);
xor U1506 (N_1506,In_1541,In_3339);
nor U1507 (N_1507,In_4811,In_2945);
nand U1508 (N_1508,In_4077,In_4955);
xor U1509 (N_1509,In_580,In_3585);
and U1510 (N_1510,In_639,In_4396);
nor U1511 (N_1511,In_1635,In_3753);
and U1512 (N_1512,In_1194,In_3432);
and U1513 (N_1513,In_1036,In_3048);
and U1514 (N_1514,In_3959,In_3732);
and U1515 (N_1515,In_2425,In_4340);
xnor U1516 (N_1516,In_4901,In_3106);
nor U1517 (N_1517,In_1054,In_3920);
xnor U1518 (N_1518,In_181,In_2067);
nor U1519 (N_1519,In_2790,In_904);
nand U1520 (N_1520,In_3485,In_2447);
nor U1521 (N_1521,In_1119,In_3489);
xnor U1522 (N_1522,In_728,In_2640);
and U1523 (N_1523,In_2936,In_4330);
or U1524 (N_1524,In_3906,In_3335);
and U1525 (N_1525,In_1008,In_2358);
and U1526 (N_1526,In_314,In_1285);
or U1527 (N_1527,In_4090,In_3517);
and U1528 (N_1528,In_4744,In_4806);
nor U1529 (N_1529,In_948,In_240);
nand U1530 (N_1530,In_164,In_565);
or U1531 (N_1531,In_2676,In_2953);
nor U1532 (N_1532,In_3931,In_599);
nor U1533 (N_1533,In_4893,In_3932);
and U1534 (N_1534,In_2282,In_549);
and U1535 (N_1535,In_2767,In_341);
nand U1536 (N_1536,In_683,In_417);
and U1537 (N_1537,In_3149,In_4092);
or U1538 (N_1538,In_2495,In_1297);
or U1539 (N_1539,In_1917,In_4979);
and U1540 (N_1540,In_2438,In_1026);
nand U1541 (N_1541,In_299,In_4607);
and U1542 (N_1542,In_2834,In_3423);
nor U1543 (N_1543,In_4332,In_964);
nor U1544 (N_1544,In_662,In_1601);
nor U1545 (N_1545,In_4775,In_369);
xor U1546 (N_1546,In_2066,In_2539);
nor U1547 (N_1547,In_1791,In_2387);
and U1548 (N_1548,In_1620,In_4229);
and U1549 (N_1549,In_922,In_2686);
nor U1550 (N_1550,In_826,In_1381);
or U1551 (N_1551,In_1717,In_3677);
or U1552 (N_1552,In_4635,In_4625);
nand U1553 (N_1553,In_4013,In_2604);
nand U1554 (N_1554,In_1705,In_1588);
or U1555 (N_1555,In_2346,In_4916);
nor U1556 (N_1556,In_2113,In_2585);
and U1557 (N_1557,In_1173,In_1810);
nand U1558 (N_1558,In_773,In_4075);
or U1559 (N_1559,In_377,In_28);
nor U1560 (N_1560,In_3130,In_1340);
xnor U1561 (N_1561,In_41,In_3686);
and U1562 (N_1562,In_3378,In_3756);
or U1563 (N_1563,In_1321,In_4477);
or U1564 (N_1564,In_1374,In_460);
and U1565 (N_1565,In_4723,In_1009);
nor U1566 (N_1566,In_2992,In_973);
and U1567 (N_1567,In_687,In_4874);
and U1568 (N_1568,In_2622,In_903);
nand U1569 (N_1569,In_2591,In_3450);
nand U1570 (N_1570,In_1174,In_1491);
and U1571 (N_1571,In_933,In_4199);
or U1572 (N_1572,In_311,In_809);
xor U1573 (N_1573,In_3996,In_2537);
nor U1574 (N_1574,In_92,In_1706);
nor U1575 (N_1575,In_2094,In_4840);
nand U1576 (N_1576,In_3630,In_4920);
or U1577 (N_1577,In_1146,In_3099);
and U1578 (N_1578,In_2428,In_1305);
or U1579 (N_1579,In_2245,In_2972);
and U1580 (N_1580,In_1851,In_4166);
xnor U1581 (N_1581,In_868,In_2961);
or U1582 (N_1582,In_2297,In_2122);
nor U1583 (N_1583,In_44,In_3670);
xor U1584 (N_1584,In_2882,In_3802);
and U1585 (N_1585,In_3892,In_4982);
nor U1586 (N_1586,In_1603,In_4685);
nor U1587 (N_1587,In_2691,In_3435);
nand U1588 (N_1588,In_913,In_4734);
nor U1589 (N_1589,In_2128,In_4253);
or U1590 (N_1590,In_776,In_1560);
or U1591 (N_1591,In_4141,In_1230);
and U1592 (N_1592,In_4438,In_4835);
xnor U1593 (N_1593,In_2394,In_1237);
or U1594 (N_1594,In_2424,In_2874);
xnor U1595 (N_1595,In_4549,In_1208);
nor U1596 (N_1596,In_2024,In_3116);
nand U1597 (N_1597,In_3982,In_4148);
or U1598 (N_1598,In_521,In_1012);
and U1599 (N_1599,In_1311,In_2985);
xor U1600 (N_1600,In_4290,In_822);
or U1601 (N_1601,In_1472,In_2544);
or U1602 (N_1602,In_915,In_3013);
and U1603 (N_1603,In_1407,In_1691);
and U1604 (N_1604,In_4784,In_1105);
and U1605 (N_1605,In_3135,In_2045);
nand U1606 (N_1606,In_4583,In_3915);
nand U1607 (N_1607,In_4863,In_2526);
nand U1608 (N_1608,In_134,In_2907);
and U1609 (N_1609,In_1263,In_3743);
nand U1610 (N_1610,In_4842,In_2911);
or U1611 (N_1611,In_178,In_1351);
nand U1612 (N_1612,In_4447,In_430);
nor U1613 (N_1613,In_3668,In_4497);
nand U1614 (N_1614,In_463,In_3818);
nand U1615 (N_1615,In_3925,In_4005);
nand U1616 (N_1616,In_1862,In_1786);
nand U1617 (N_1617,In_2427,In_1165);
and U1618 (N_1618,In_2954,In_2156);
nor U1619 (N_1619,In_947,In_3421);
or U1620 (N_1620,In_637,In_3086);
nor U1621 (N_1621,In_1217,In_893);
nor U1622 (N_1622,In_4442,In_3522);
or U1623 (N_1623,In_3973,In_3097);
and U1624 (N_1624,In_4746,In_4355);
nand U1625 (N_1625,In_1598,In_4631);
and U1626 (N_1626,In_1450,In_165);
nor U1627 (N_1627,In_458,In_2707);
nand U1628 (N_1628,In_1708,In_2464);
xnor U1629 (N_1629,In_4244,In_2842);
or U1630 (N_1630,In_4193,In_1547);
or U1631 (N_1631,In_505,In_3627);
nand U1632 (N_1632,In_3197,In_3493);
nand U1633 (N_1633,In_345,In_2881);
and U1634 (N_1634,In_29,In_2466);
nor U1635 (N_1635,In_4149,In_909);
and U1636 (N_1636,In_786,In_1076);
nand U1637 (N_1637,In_4560,In_4280);
nand U1638 (N_1638,In_1113,In_1416);
nor U1639 (N_1639,In_995,In_4256);
nor U1640 (N_1640,In_541,In_986);
or U1641 (N_1641,In_1192,In_15);
and U1642 (N_1642,In_3163,In_2462);
nor U1643 (N_1643,In_1212,In_3620);
nand U1644 (N_1644,In_3162,In_4308);
or U1645 (N_1645,In_2013,In_1710);
and U1646 (N_1646,In_1245,In_2554);
and U1647 (N_1647,In_4604,In_4392);
nor U1648 (N_1648,In_1727,In_322);
and U1649 (N_1649,In_1337,In_2226);
nand U1650 (N_1650,In_1314,In_1550);
or U1651 (N_1651,In_2860,In_3011);
nand U1652 (N_1652,In_2572,In_2202);
nor U1653 (N_1653,In_3248,In_4725);
nor U1654 (N_1654,In_3795,In_4365);
and U1655 (N_1655,In_3632,In_1435);
or U1656 (N_1656,In_4704,In_859);
xnor U1657 (N_1657,In_1352,In_2672);
xnor U1658 (N_1658,In_2135,In_30);
or U1659 (N_1659,In_4088,In_1709);
nand U1660 (N_1660,In_3520,In_3733);
or U1661 (N_1661,In_2600,In_3807);
and U1662 (N_1662,In_2740,In_3031);
nor U1663 (N_1663,In_3342,In_3189);
or U1664 (N_1664,In_708,In_4255);
nor U1665 (N_1665,In_1661,In_4375);
nor U1666 (N_1666,In_4260,In_87);
nand U1667 (N_1667,In_4226,In_887);
and U1668 (N_1668,In_748,In_3958);
nor U1669 (N_1669,In_2795,In_738);
and U1670 (N_1670,In_186,In_3328);
or U1671 (N_1671,In_2010,In_2287);
nand U1672 (N_1672,In_3177,In_3783);
nand U1673 (N_1673,In_659,In_2873);
or U1674 (N_1674,In_1267,In_858);
nor U1675 (N_1675,In_2720,In_4519);
or U1676 (N_1676,In_1999,In_2525);
or U1677 (N_1677,In_1292,In_3358);
nand U1678 (N_1678,In_4657,In_333);
xnor U1679 (N_1679,In_2105,In_4903);
or U1680 (N_1680,In_3280,In_702);
xor U1681 (N_1681,In_2334,In_3491);
nor U1682 (N_1682,In_3046,In_811);
nand U1683 (N_1683,In_2234,In_13);
nor U1684 (N_1684,In_4425,In_2456);
nor U1685 (N_1685,In_347,In_3535);
or U1686 (N_1686,In_2291,In_1153);
nor U1687 (N_1687,In_4487,In_174);
nor U1688 (N_1688,In_1641,In_3202);
nand U1689 (N_1689,In_1747,In_2145);
nor U1690 (N_1690,In_1814,In_4676);
or U1691 (N_1691,In_4197,In_3369);
xor U1692 (N_1692,In_4994,In_2831);
and U1693 (N_1693,In_4974,In_4112);
nor U1694 (N_1694,In_2350,In_3382);
and U1695 (N_1695,In_440,In_4185);
or U1696 (N_1696,In_3692,In_2898);
xnor U1697 (N_1697,In_4929,In_2634);
nand U1698 (N_1698,In_3397,In_2395);
xor U1699 (N_1699,In_31,In_1168);
or U1700 (N_1700,In_4697,In_1243);
nor U1701 (N_1701,In_3247,In_4298);
nand U1702 (N_1702,In_2311,In_4991);
nor U1703 (N_1703,In_11,In_647);
or U1704 (N_1704,In_3805,In_1264);
nand U1705 (N_1705,In_3902,In_2057);
xor U1706 (N_1706,In_4428,In_578);
nand U1707 (N_1707,In_3634,In_2332);
nor U1708 (N_1708,In_994,In_1730);
and U1709 (N_1709,In_3024,In_3207);
nor U1710 (N_1710,In_4561,In_1024);
nand U1711 (N_1711,In_4252,In_4872);
nor U1712 (N_1712,In_2048,In_2551);
nand U1713 (N_1713,In_2055,In_4717);
or U1714 (N_1714,In_247,In_2082);
nor U1715 (N_1715,In_4817,In_2938);
xor U1716 (N_1716,In_3956,In_4756);
nand U1717 (N_1717,In_835,In_523);
nor U1718 (N_1718,In_305,In_3638);
and U1719 (N_1719,In_2606,In_779);
xnor U1720 (N_1720,In_4505,In_1488);
xnor U1721 (N_1721,In_598,In_4769);
nand U1722 (N_1722,In_1872,In_337);
nor U1723 (N_1723,In_485,In_1331);
or U1724 (N_1724,In_1409,In_2827);
and U1725 (N_1725,In_2420,In_2312);
nor U1726 (N_1726,In_2742,In_4848);
or U1727 (N_1727,In_2749,In_3210);
or U1728 (N_1728,In_1943,In_2366);
or U1729 (N_1729,In_4766,In_512);
nor U1730 (N_1730,In_2359,In_517);
and U1731 (N_1731,In_2315,In_1181);
or U1732 (N_1732,In_981,In_2467);
nor U1733 (N_1733,In_2191,In_1440);
nand U1734 (N_1734,In_2958,In_4416);
nor U1735 (N_1735,In_2225,In_2124);
or U1736 (N_1736,In_3293,In_2);
and U1737 (N_1737,In_1655,In_1465);
or U1738 (N_1738,In_559,In_2390);
or U1739 (N_1739,In_3324,In_1250);
and U1740 (N_1740,In_3945,In_4996);
nor U1741 (N_1741,In_619,In_2886);
xnor U1742 (N_1742,In_546,In_1057);
or U1743 (N_1743,In_4263,In_695);
nor U1744 (N_1744,In_681,In_2176);
or U1745 (N_1745,In_2399,In_2711);
xnor U1746 (N_1746,In_1195,In_2200);
or U1747 (N_1747,In_3771,In_4481);
and U1748 (N_1748,In_4751,In_75);
or U1749 (N_1749,In_312,In_2777);
xor U1750 (N_1750,In_2421,In_610);
xor U1751 (N_1751,In_4458,In_870);
and U1752 (N_1752,In_3370,In_4126);
nand U1753 (N_1753,In_4988,In_2611);
xor U1754 (N_1754,In_2836,In_4249);
or U1755 (N_1755,In_3460,In_2224);
nand U1756 (N_1756,In_1725,In_2704);
nand U1757 (N_1757,In_3622,In_3402);
nor U1758 (N_1758,In_3603,In_3355);
or U1759 (N_1759,In_1765,In_2784);
or U1760 (N_1760,In_1172,In_889);
or U1761 (N_1761,In_2319,In_3594);
nand U1762 (N_1762,In_962,In_3829);
and U1763 (N_1763,In_2716,In_4089);
or U1764 (N_1764,In_3636,In_4137);
or U1765 (N_1765,In_1052,In_2538);
xor U1766 (N_1766,In_3085,In_213);
nand U1767 (N_1767,In_2733,In_1739);
or U1768 (N_1768,In_3294,In_1219);
nand U1769 (N_1769,In_418,In_3314);
or U1770 (N_1770,In_3516,In_139);
and U1771 (N_1771,In_3498,In_1469);
nor U1772 (N_1772,In_828,In_83);
and U1773 (N_1773,In_2619,In_3117);
and U1774 (N_1774,In_2789,In_4689);
or U1775 (N_1775,In_238,In_611);
nor U1776 (N_1776,In_4816,In_37);
nor U1777 (N_1777,In_4207,In_4899);
and U1778 (N_1778,In_4711,In_3769);
nand U1779 (N_1779,In_2916,In_1983);
and U1780 (N_1780,In_3691,In_1619);
or U1781 (N_1781,In_3748,In_3340);
or U1782 (N_1782,In_231,In_4589);
nand U1783 (N_1783,In_576,In_2757);
nor U1784 (N_1784,In_2419,In_987);
nand U1785 (N_1785,In_4966,In_984);
xnor U1786 (N_1786,In_3754,In_1065);
nor U1787 (N_1787,In_2696,In_2957);
and U1788 (N_1788,In_1116,In_627);
nor U1789 (N_1789,In_3400,In_104);
nand U1790 (N_1790,In_3054,In_2381);
nand U1791 (N_1791,In_4691,In_2019);
nand U1792 (N_1792,In_938,In_2560);
and U1793 (N_1793,In_4490,In_2369);
or U1794 (N_1794,In_2900,In_3146);
and U1795 (N_1795,In_1358,In_1758);
nand U1796 (N_1796,In_3184,In_2794);
and U1797 (N_1797,In_1649,In_2817);
nor U1798 (N_1798,In_1176,In_4946);
nor U1799 (N_1799,In_2501,In_1492);
or U1800 (N_1800,In_1964,In_1609);
nor U1801 (N_1801,In_1301,In_4701);
and U1802 (N_1802,In_2947,In_2645);
nand U1803 (N_1803,In_742,In_2367);
xor U1804 (N_1804,In_1441,In_1590);
and U1805 (N_1805,In_3845,In_4042);
nor U1806 (N_1806,In_2049,In_3908);
nand U1807 (N_1807,In_3170,In_4516);
nand U1808 (N_1808,In_2341,In_3629);
nor U1809 (N_1809,In_3713,In_382);
and U1810 (N_1810,In_209,In_2510);
xnor U1811 (N_1811,In_791,In_1672);
nand U1812 (N_1812,In_3846,In_4976);
xor U1813 (N_1813,In_4067,In_2839);
and U1814 (N_1814,In_2807,In_1589);
and U1815 (N_1815,In_1039,In_2351);
and U1816 (N_1816,In_1178,In_3357);
and U1817 (N_1817,In_3076,In_2241);
nor U1818 (N_1818,In_1455,In_1534);
nand U1819 (N_1819,In_4097,In_4455);
nand U1820 (N_1820,In_1528,In_618);
and U1821 (N_1821,In_2344,In_4353);
or U1822 (N_1822,In_2805,In_2682);
nand U1823 (N_1823,In_2962,In_3838);
or U1824 (N_1824,In_958,In_741);
or U1825 (N_1825,In_3456,In_2206);
or U1826 (N_1826,In_4082,In_4521);
nand U1827 (N_1827,In_2000,In_4579);
and U1828 (N_1828,In_2473,In_4813);
or U1829 (N_1829,In_3530,In_914);
or U1830 (N_1830,In_4273,In_3891);
xor U1831 (N_1831,In_1648,In_2855);
and U1832 (N_1832,In_4004,In_2593);
nand U1833 (N_1833,In_3034,In_3830);
nand U1834 (N_1834,In_1233,In_3312);
nor U1835 (N_1835,In_4508,In_1071);
nor U1836 (N_1836,In_290,In_292);
nor U1837 (N_1837,In_4228,In_4129);
xor U1838 (N_1838,In_802,In_180);
nor U1839 (N_1839,In_4594,In_4777);
xnor U1840 (N_1840,In_1640,In_3640);
nor U1841 (N_1841,In_4095,In_4833);
xor U1842 (N_1842,In_4897,In_1746);
nand U1843 (N_1843,In_4236,In_4599);
nand U1844 (N_1844,In_1149,In_3876);
xnor U1845 (N_1845,In_2041,In_4672);
nand U1846 (N_1846,In_2887,In_3073);
nor U1847 (N_1847,In_3577,In_4429);
nand U1848 (N_1848,In_1696,In_1896);
nor U1849 (N_1849,In_3317,In_2813);
xnor U1850 (N_1850,In_461,In_3366);
or U1851 (N_1851,In_1736,In_3886);
nand U1852 (N_1852,In_2621,In_2642);
nand U1853 (N_1853,In_3490,In_373);
or U1854 (N_1854,In_2700,In_1341);
nor U1855 (N_1855,In_1498,In_4731);
xnor U1856 (N_1856,In_3648,In_514);
nor U1857 (N_1857,In_3719,In_2748);
or U1858 (N_1858,In_4036,In_1816);
or U1859 (N_1859,In_4221,In_1431);
xor U1860 (N_1860,In_1937,In_614);
nand U1861 (N_1861,In_3526,In_3862);
or U1862 (N_1862,In_3297,In_2963);
and U1863 (N_1863,In_207,In_754);
or U1864 (N_1864,In_2106,In_872);
nor U1865 (N_1865,In_697,In_3825);
xnor U1866 (N_1866,In_3384,In_2244);
and U1867 (N_1867,In_4285,In_723);
or U1868 (N_1868,In_2729,In_2298);
xnor U1869 (N_1869,In_854,In_4306);
nor U1870 (N_1870,In_2862,In_3077);
and U1871 (N_1871,In_1868,In_4367);
or U1872 (N_1872,In_3859,In_4435);
nand U1873 (N_1873,In_1843,In_2698);
nand U1874 (N_1874,In_679,In_3215);
nand U1875 (N_1875,In_1278,In_3635);
and U1876 (N_1876,In_4305,In_3270);
and U1877 (N_1877,In_203,In_4170);
or U1878 (N_1878,In_704,In_919);
or U1879 (N_1879,In_3214,In_4008);
nor U1880 (N_1880,In_4986,In_3778);
nand U1881 (N_1881,In_3610,In_4354);
and U1882 (N_1882,In_1303,In_2574);
or U1883 (N_1883,In_4914,In_4951);
and U1884 (N_1884,In_248,In_3199);
nor U1885 (N_1885,In_328,In_3710);
and U1886 (N_1886,In_4588,In_1763);
xnor U1887 (N_1887,In_335,In_4073);
and U1888 (N_1888,In_4032,In_3555);
nor U1889 (N_1889,In_3968,In_3809);
xor U1890 (N_1890,In_1070,In_451);
nand U1891 (N_1891,In_4547,In_274);
and U1892 (N_1892,In_2518,In_3359);
nor U1893 (N_1893,In_2377,In_1490);
and U1894 (N_1894,In_2925,In_220);
xor U1895 (N_1895,In_3870,In_4208);
and U1896 (N_1896,In_2578,In_2750);
nand U1897 (N_1897,In_1038,In_4846);
nand U1898 (N_1898,In_1255,In_4358);
or U1899 (N_1899,In_1554,In_1757);
nor U1900 (N_1900,In_612,In_3279);
nor U1901 (N_1901,In_1656,In_945);
and U1902 (N_1902,In_2483,In_4663);
or U1903 (N_1903,In_1027,In_807);
nor U1904 (N_1904,In_175,In_1281);
nand U1905 (N_1905,In_4768,In_3405);
xor U1906 (N_1906,In_3182,In_2362);
nand U1907 (N_1907,In_3265,In_4344);
xnor U1908 (N_1908,In_2455,In_185);
nor U1909 (N_1909,In_2258,In_4525);
or U1910 (N_1910,In_466,In_1091);
nor U1911 (N_1911,In_2743,In_2253);
and U1912 (N_1912,In_2803,In_3761);
xor U1913 (N_1913,In_2688,In_1015);
and U1914 (N_1914,In_1918,In_782);
or U1915 (N_1915,In_1645,In_3880);
nand U1916 (N_1916,In_1283,In_4962);
nand U1917 (N_1917,In_1310,In_2871);
and U1918 (N_1918,In_4739,In_4924);
nor U1919 (N_1919,In_1654,In_4552);
nand U1920 (N_1920,In_441,In_1906);
nor U1921 (N_1921,In_4590,In_4027);
or U1922 (N_1922,In_531,In_743);
nor U1923 (N_1923,In_524,In_1345);
and U1924 (N_1924,In_3057,In_2738);
and U1925 (N_1925,In_999,In_4116);
or U1926 (N_1926,In_4702,In_2952);
nor U1927 (N_1927,In_2303,In_4086);
nand U1928 (N_1928,In_3600,In_1307);
nor U1929 (N_1929,In_937,In_4621);
nor U1930 (N_1930,In_79,In_3407);
or U1931 (N_1931,In_3425,In_2509);
nor U1932 (N_1932,In_975,In_1793);
and U1933 (N_1933,In_1781,In_4834);
xnor U1934 (N_1934,In_2562,In_927);
or U1935 (N_1935,In_1196,In_4070);
and U1936 (N_1936,In_3020,In_2610);
and U1937 (N_1937,In_1632,In_4921);
nor U1938 (N_1938,In_4820,In_3363);
and U1939 (N_1939,In_2709,In_447);
and U1940 (N_1940,In_631,In_705);
nand U1941 (N_1941,In_4379,In_1713);
xnor U1942 (N_1942,In_3112,In_711);
nor U1943 (N_1943,In_2186,In_2849);
and U1944 (N_1944,In_1876,In_4394);
and U1945 (N_1945,In_3693,In_4142);
or U1946 (N_1946,In_651,In_4989);
and U1947 (N_1947,In_584,In_2205);
and U1948 (N_1948,In_3689,In_4059);
nor U1949 (N_1949,In_2810,In_76);
nor U1950 (N_1950,In_2555,In_2579);
nand U1951 (N_1951,In_2099,In_2162);
and U1952 (N_1952,In_4758,In_408);
xor U1953 (N_1953,In_544,In_3404);
xnor U1954 (N_1954,In_3815,In_4930);
nor U1955 (N_1955,In_558,In_1762);
or U1956 (N_1956,In_1574,In_2930);
nor U1957 (N_1957,In_793,In_3768);
nor U1958 (N_1958,In_3453,In_1136);
nand U1959 (N_1959,In_2090,In_244);
or U1960 (N_1960,In_2274,In_4399);
nor U1961 (N_1961,In_2931,In_72);
nand U1962 (N_1962,In_976,In_297);
or U1963 (N_1963,In_4327,In_1960);
nor U1964 (N_1964,In_200,In_2116);
nor U1965 (N_1965,In_2573,In_2272);
or U1966 (N_1966,In_4941,In_527);
nand U1967 (N_1967,In_2435,In_3196);
nor U1968 (N_1968,In_1815,In_3377);
or U1969 (N_1969,In_1471,In_2534);
xor U1970 (N_1970,In_2267,In_2683);
and U1971 (N_1971,In_4787,In_3864);
and U1972 (N_1972,In_972,In_761);
nand U1973 (N_1973,In_2030,In_3039);
or U1974 (N_1974,In_2806,In_1097);
nand U1975 (N_1975,In_475,In_235);
nor U1976 (N_1976,In_2801,In_1007);
xnor U1977 (N_1977,In_4049,In_3262);
xor U1978 (N_1978,In_1254,In_2605);
or U1979 (N_1979,In_4110,In_4615);
nand U1980 (N_1980,In_4282,In_1671);
xnor U1981 (N_1981,In_3142,In_1348);
or U1982 (N_1982,In_3853,In_214);
nor U1983 (N_1983,In_1798,In_3952);
nand U1984 (N_1984,In_1373,In_1809);
and U1985 (N_1985,In_713,In_3500);
nor U1986 (N_1986,In_2073,In_2261);
nand U1987 (N_1987,In_3187,In_3376);
and U1988 (N_1988,In_1112,In_1279);
nand U1989 (N_1989,In_623,In_4515);
or U1990 (N_1990,In_1456,In_1701);
and U1991 (N_1991,In_2935,In_3043);
nand U1992 (N_1992,In_851,In_4919);
or U1993 (N_1993,In_1160,In_3353);
and U1994 (N_1994,In_504,In_2699);
or U1995 (N_1995,In_3326,In_4939);
nand U1996 (N_1996,In_1779,In_496);
or U1997 (N_1997,In_2599,In_1037);
nor U1998 (N_1998,In_1258,In_1055);
or U1999 (N_1999,In_3245,In_2531);
or U2000 (N_2000,In_4908,In_698);
or U2001 (N_2001,In_1108,In_2697);
nor U2002 (N_2002,In_1959,In_1385);
or U2003 (N_2003,In_882,In_3558);
xor U2004 (N_2004,In_4861,In_2422);
or U2005 (N_2005,In_3836,In_2006);
and U2006 (N_2006,In_724,In_1270);
and U2007 (N_2007,In_2064,In_184);
or U2008 (N_2008,In_636,In_894);
nand U2009 (N_2009,In_2753,In_2065);
or U2010 (N_2010,In_4389,In_3495);
or U2011 (N_2011,In_3601,In_3403);
and U2012 (N_2012,In_2677,In_772);
and U2013 (N_2013,In_3649,In_3180);
or U2014 (N_2014,In_2001,In_3016);
nand U2015 (N_2015,In_1625,In_1047);
nand U2016 (N_2016,In_2994,In_853);
nor U2017 (N_2017,In_756,In_4707);
nor U2018 (N_2018,In_1451,In_4331);
or U2019 (N_2019,In_64,In_2417);
nand U2020 (N_2020,In_2009,In_4062);
nor U2021 (N_2021,In_3847,In_2276);
and U2022 (N_2022,In_330,In_3373);
and U2023 (N_2023,In_3260,In_2800);
nand U2024 (N_2024,In_817,In_3962);
and U2025 (N_2025,In_789,In_511);
and U2026 (N_2026,In_974,In_3315);
nand U2027 (N_2027,In_3560,In_1749);
nor U2028 (N_2028,In_455,In_2070);
xnor U2029 (N_2029,In_4904,In_701);
nand U2030 (N_2030,In_4494,In_1093);
and U2031 (N_2031,In_4598,In_4564);
nand U2032 (N_2032,In_1910,In_2656);
nor U2033 (N_2033,In_815,In_3514);
or U2034 (N_2034,In_513,In_4267);
or U2035 (N_2035,In_4618,In_3714);
or U2036 (N_2036,In_2763,In_3894);
nand U2037 (N_2037,In_3777,In_3313);
and U2038 (N_2038,In_661,In_493);
xor U2039 (N_2039,In_4361,In_53);
or U2040 (N_2040,In_1084,In_4007);
and U2041 (N_2041,In_3671,In_3266);
xor U2042 (N_2042,In_388,In_4667);
nand U2043 (N_2043,In_3984,In_4295);
nand U2044 (N_2044,In_4887,In_323);
or U2045 (N_2045,In_1608,In_1796);
or U2046 (N_2046,In_1171,In_90);
and U2047 (N_2047,In_4937,In_403);
or U2048 (N_2048,In_3613,In_4743);
xnor U2049 (N_2049,In_4576,In_2576);
nor U2050 (N_2050,In_324,In_1228);
nor U2051 (N_2051,In_1106,In_14);
or U2052 (N_2052,In_600,In_757);
nor U2053 (N_2053,In_3061,In_4317);
nor U2054 (N_2054,In_3867,In_4770);
and U2055 (N_2055,In_3008,In_821);
nor U2056 (N_2056,In_4364,In_2974);
nand U2057 (N_2057,In_4019,In_3623);
and U2058 (N_2058,In_2970,In_4422);
nor U2059 (N_2059,In_413,In_1594);
and U2060 (N_2060,In_1970,In_1826);
nand U2061 (N_2061,In_432,In_365);
and U2062 (N_2062,In_4620,In_1629);
nor U2063 (N_2063,In_40,In_1206);
nor U2064 (N_2064,In_2689,In_170);
nand U2065 (N_2065,In_1030,In_2109);
nand U2066 (N_2066,In_89,In_4923);
and U2067 (N_2067,In_4424,In_1209);
nor U2068 (N_2068,In_1909,In_4869);
xor U2069 (N_2069,In_4300,In_2858);
nor U2070 (N_2070,In_4251,In_3429);
or U2071 (N_2071,In_2036,In_2912);
or U2072 (N_2072,In_3897,In_123);
nand U2073 (N_2073,In_1752,In_2208);
nor U2074 (N_2074,In_4796,In_57);
nor U2075 (N_2075,In_3628,In_1889);
nor U2076 (N_2076,In_258,In_2517);
xor U2077 (N_2077,In_1421,In_4954);
nand U2078 (N_2078,In_2309,In_2477);
nand U2079 (N_2079,In_1355,In_632);
or U2080 (N_2080,In_3553,In_4065);
xnor U2081 (N_2081,In_1597,In_396);
or U2082 (N_2082,In_902,In_3219);
or U2083 (N_2083,In_4889,In_719);
nor U2084 (N_2084,In_3440,In_2458);
or U2085 (N_2085,In_3469,In_4641);
and U2086 (N_2086,In_2152,In_1754);
nand U2087 (N_2087,In_4324,In_331);
and U2088 (N_2088,In_3556,In_1939);
and U2089 (N_2089,In_4187,In_1246);
nor U2090 (N_2090,In_1557,In_3419);
and U2091 (N_2091,In_412,In_275);
nand U2092 (N_2092,In_1866,In_1014);
nand U2093 (N_2093,In_344,In_985);
or U2094 (N_2094,In_4814,In_4378);
nor U2095 (N_2095,In_4706,In_21);
nor U2096 (N_2096,In_4172,In_3263);
and U2097 (N_2097,In_3597,In_4217);
or U2098 (N_2098,In_1023,In_3758);
and U2099 (N_2099,In_897,In_4556);
nand U2100 (N_2100,In_2110,In_1835);
and U2101 (N_2101,In_4759,In_834);
nand U2102 (N_2102,In_3878,In_3213);
or U2103 (N_2103,In_62,In_633);
or U2104 (N_2104,In_4851,In_2948);
or U2105 (N_2105,In_1072,In_2991);
or U2106 (N_2106,In_3174,In_3261);
nand U2107 (N_2107,In_1621,In_1788);
nor U2108 (N_2108,In_6,In_1299);
or U2109 (N_2109,In_4212,In_2262);
nor U2110 (N_2110,In_4882,In_1673);
nor U2111 (N_2111,In_3887,In_1854);
xnor U2112 (N_2112,In_4915,In_2885);
nand U2113 (N_2113,In_3724,In_3167);
and U2114 (N_2114,In_4571,In_4296);
nor U2115 (N_2115,In_1188,In_3394);
and U2116 (N_2116,In_899,In_2568);
or U2117 (N_2117,In_378,In_1215);
xnor U2118 (N_2118,In_4202,In_2588);
and U2119 (N_2119,In_3143,In_4637);
or U2120 (N_2120,In_2630,In_4410);
nor U2121 (N_2121,In_3299,In_847);
or U2122 (N_2122,In_340,In_2918);
and U2123 (N_2123,In_112,In_3059);
and U2124 (N_2124,In_3296,In_1850);
nand U2125 (N_2125,In_665,In_491);
nand U2126 (N_2126,In_4523,In_678);
and U2127 (N_2127,In_4302,In_4651);
nor U2128 (N_2128,In_1870,In_1187);
and U2129 (N_2129,In_4585,In_2973);
and U2130 (N_2130,In_996,In_2413);
and U2131 (N_2131,In_3287,In_2108);
nor U2132 (N_2132,In_3365,In_397);
or U2133 (N_2133,In_2410,In_3826);
nand U2134 (N_2134,In_230,In_3998);
or U2135 (N_2135,In_4336,In_3700);
nand U2136 (N_2136,In_936,In_4764);
xor U2137 (N_2137,In_141,In_3755);
xor U2138 (N_2138,In_3338,In_1446);
and U2139 (N_2139,In_1789,In_3336);
nand U2140 (N_2140,In_1203,In_3361);
and U2141 (N_2141,In_67,In_9);
or U2142 (N_2142,In_1325,In_4002);
xor U2143 (N_2143,In_2828,In_1061);
nand U2144 (N_2144,In_3081,In_3391);
nand U2145 (N_2145,In_2822,In_2796);
and U2146 (N_2146,In_363,In_1703);
nand U2147 (N_2147,In_3089,In_4029);
or U2148 (N_2148,In_2133,In_1063);
nor U2149 (N_2149,In_1335,In_1985);
and U2150 (N_2150,In_3935,In_1613);
xor U2151 (N_2151,In_1571,In_1164);
xnor U2152 (N_2152,In_3173,In_1875);
nor U2153 (N_2153,In_1432,In_801);
nand U2154 (N_2154,In_4578,In_4284);
xor U2155 (N_2155,In_3198,In_543);
nor U2156 (N_2156,In_1732,In_2025);
nor U2157 (N_2157,In_4674,In_4278);
and U2158 (N_2158,In_1487,In_1386);
nand U2159 (N_2159,In_2594,In_1103);
nor U2160 (N_2160,In_1760,In_2921);
and U2161 (N_2161,In_3028,In_1396);
or U2162 (N_2162,In_2411,In_3661);
and U2163 (N_2163,In_734,In_4017);
xor U2164 (N_2164,In_4774,In_657);
or U2165 (N_2165,In_4928,In_2164);
or U2166 (N_2166,In_4066,In_196);
and U2167 (N_2167,In_266,In_4856);
and U2168 (N_2168,In_2323,In_3441);
xor U2169 (N_2169,In_1829,In_1420);
nand U2170 (N_2170,In_2506,In_4656);
or U2171 (N_2171,In_2448,In_3570);
or U2172 (N_2172,In_908,In_4911);
nor U2173 (N_2173,In_2548,In_3547);
and U2174 (N_2174,In_2943,In_2721);
nor U2175 (N_2175,In_587,In_4220);
nor U2176 (N_2176,In_3773,In_4388);
nand U2177 (N_2177,In_3108,In_1966);
nand U2178 (N_2178,In_2107,In_4963);
or U2179 (N_2179,In_4905,In_1865);
nor U2180 (N_2180,In_2058,In_395);
or U2181 (N_2181,In_4627,In_3254);
xor U2182 (N_2182,In_1041,In_2932);
and U2183 (N_2183,In_1777,In_153);
or U2184 (N_2184,In_1400,In_2450);
or U2185 (N_2185,In_2308,In_3900);
nor U2186 (N_2186,In_1457,In_4452);
nand U2187 (N_2187,In_4530,In_1240);
nor U2188 (N_2188,In_781,In_2414);
and U2189 (N_2189,In_2996,In_2201);
nand U2190 (N_2190,In_2968,In_1402);
nor U2191 (N_2191,In_2360,In_4390);
or U2192 (N_2192,In_4072,In_2879);
nor U2193 (N_2193,In_1530,In_2978);
and U2194 (N_2194,In_1474,In_443);
nor U2195 (N_2195,In_1986,In_3718);
nand U2196 (N_2196,In_3746,In_448);
nand U2197 (N_2197,In_4323,In_3350);
or U2198 (N_2198,In_2595,In_3757);
nor U2199 (N_2199,In_3987,In_111);
or U2200 (N_2200,In_4337,In_1844);
nand U2201 (N_2201,In_3282,In_2997);
nand U2202 (N_2202,In_4039,In_2052);
or U2203 (N_2203,In_760,In_1074);
nor U2204 (N_2204,In_778,In_1744);
nand U2205 (N_2205,In_3947,In_1109);
nand U2206 (N_2206,In_1743,In_173);
or U2207 (N_2207,In_4444,In_707);
xnor U2208 (N_2208,In_4194,In_579);
or U2209 (N_2209,In_93,In_4940);
xor U2210 (N_2210,In_2418,In_2513);
xnor U2211 (N_2211,In_991,In_1773);
or U2212 (N_2212,In_4316,In_3745);
xnor U2213 (N_2213,In_3433,In_1320);
nor U2214 (N_2214,In_2132,In_4468);
nor U2215 (N_2215,In_1764,In_3528);
nand U2216 (N_2216,In_3860,In_4155);
nand U2217 (N_2217,In_520,In_334);
nand U2218 (N_2218,In_4159,In_1392);
nand U2219 (N_2219,In_4616,In_24);
or U2220 (N_2220,In_3812,In_4417);
nor U2221 (N_2221,In_554,In_4136);
nand U2222 (N_2222,In_2949,In_3392);
nor U2223 (N_2223,In_1584,In_1979);
and U2224 (N_2224,In_3861,In_2519);
and U2225 (N_2225,In_2398,In_2812);
nand U2226 (N_2226,In_3548,In_1511);
or U2227 (N_2227,In_100,In_487);
xnor U2228 (N_2228,In_2345,In_3901);
nand U2229 (N_2229,In_4329,In_3090);
nand U2230 (N_2230,In_4984,In_1087);
nand U2231 (N_2231,In_234,In_3794);
nor U2232 (N_2232,In_740,In_1572);
or U2233 (N_2233,In_2914,In_4933);
nand U2234 (N_2234,In_3319,In_819);
nor U2235 (N_2235,In_4293,In_2318);
nor U2236 (N_2236,In_4241,In_1933);
nor U2237 (N_2237,In_3562,In_3029);
xor U2238 (N_2238,In_873,In_2575);
nor U2239 (N_2239,In_1712,In_3949);
and U2240 (N_2240,In_2264,In_2651);
nor U2241 (N_2241,In_4409,In_2533);
and U2242 (N_2242,In_2713,In_481);
nand U2243 (N_2243,In_2596,In_371);
and U2244 (N_2244,In_3936,In_758);
nand U2245 (N_2245,In_2890,In_4372);
xnor U2246 (N_2246,In_4677,In_3183);
nor U2247 (N_2247,In_2866,In_2295);
xnor U2248 (N_2248,In_1704,In_982);
and U2249 (N_2249,In_2920,In_218);
nand U2250 (N_2250,In_3676,In_2445);
or U2251 (N_2251,In_729,In_4687);
or U2252 (N_2252,In_1384,In_3216);
nor U2253 (N_2253,In_4577,In_1029);
and U2254 (N_2254,In_3578,In_4931);
nand U2255 (N_2255,In_4103,In_4031);
nand U2256 (N_2256,In_3762,In_1094);
or U2257 (N_2257,In_953,In_486);
or U2258 (N_2258,In_77,In_3568);
or U2259 (N_2259,In_1718,In_694);
nand U2260 (N_2260,In_4411,In_638);
nor U2261 (N_2261,In_1252,In_2504);
and U2262 (N_2262,In_1138,In_1847);
or U2263 (N_2263,In_1302,In_3110);
or U2264 (N_2264,In_1111,In_4611);
xor U2265 (N_2265,In_516,In_3153);
nand U2266 (N_2266,In_2512,In_1236);
nand U2267 (N_2267,In_273,In_788);
xnor U2268 (N_2268,In_4622,In_534);
and U2269 (N_2269,In_630,In_1971);
or U2270 (N_2270,In_39,In_431);
xnor U2271 (N_2271,In_4767,In_452);
nand U2272 (N_2272,In_1582,In_4376);
and U2273 (N_2273,In_2964,In_3484);
nand U2274 (N_2274,In_2995,In_1867);
and U2275 (N_2275,In_2491,In_3387);
nand U2276 (N_2276,In_389,In_699);
nand U2277 (N_2277,In_198,In_1934);
nand U2278 (N_2278,In_2089,In_1098);
and U2279 (N_2279,In_1495,In_3360);
nand U2280 (N_2280,In_427,In_4189);
and U2281 (N_2281,In_1800,In_3960);
and U2282 (N_2282,In_264,In_2724);
nor U2283 (N_2283,In_2695,In_1893);
nand U2284 (N_2284,In_1819,In_4496);
nor U2285 (N_2285,In_2136,In_2168);
and U2286 (N_2286,In_3808,In_1089);
nor U2287 (N_2287,In_2068,In_1508);
or U2288 (N_2288,In_4345,In_3168);
nand U2289 (N_2289,In_3683,In_1665);
and U2290 (N_2290,In_1464,In_3889);
or U2291 (N_2291,In_318,In_1042);
nor U2292 (N_2292,In_4935,In_81);
nand U2293 (N_2293,In_2966,In_1734);
and U2294 (N_2294,In_4509,In_641);
xnor U2295 (N_2295,In_3222,In_4343);
nor U2296 (N_2296,In_3513,In_583);
nand U2297 (N_2297,In_4231,In_4850);
nor U2298 (N_2298,In_2808,In_4450);
nand U2299 (N_2299,In_1060,In_1614);
nor U2300 (N_2300,In_997,In_3033);
or U2301 (N_2301,In_381,In_864);
nand U2302 (N_2302,In_1987,In_1808);
nor U2303 (N_2303,In_942,In_2184);
nand U2304 (N_2304,In_2565,In_1577);
or U2305 (N_2305,In_4214,In_2667);
and U2306 (N_2306,In_2157,In_4570);
or U2307 (N_2307,In_1118,In_4737);
xnor U2308 (N_2308,In_2841,In_3711);
nor U2309 (N_2309,In_419,In_1226);
nand U2310 (N_2310,In_3203,In_2771);
and U2311 (N_2311,In_2054,In_1394);
and U2312 (N_2312,In_1591,In_1952);
and U2313 (N_2313,In_2820,In_3169);
nand U2314 (N_2314,In_3330,In_2892);
and U2315 (N_2315,In_2203,In_1535);
nor U2316 (N_2316,In_3379,In_3070);
nand U2317 (N_2317,In_2821,In_4745);
and U2318 (N_2318,In_2153,In_3872);
nor U2319 (N_2319,In_2391,In_2888);
and U2320 (N_2320,In_1897,In_2098);
nor U2321 (N_2321,In_1121,In_1497);
and U2322 (N_2322,In_540,In_4374);
xor U2323 (N_2323,In_2175,In_4033);
nand U2324 (N_2324,In_715,In_3917);
nor U2325 (N_2325,In_88,In_109);
nor U2326 (N_2326,In_2703,In_1317);
nor U2327 (N_2327,In_1241,In_3482);
nor U2328 (N_2328,In_1485,In_732);
and U2329 (N_2329,In_2294,In_693);
nand U2330 (N_2330,In_1694,In_245);
and U2331 (N_2331,In_1792,In_1046);
nor U2332 (N_2332,In_4959,In_1478);
and U2333 (N_2333,In_3505,In_2278);
nand U2334 (N_2334,In_616,In_4087);
nor U2335 (N_2335,In_4461,In_4326);
nand U2336 (N_2336,In_2497,In_4501);
nor U2337 (N_2337,In_2293,In_349);
nor U2338 (N_2338,In_2666,In_1700);
nor U2339 (N_2339,In_2553,In_3951);
and U2340 (N_2340,In_4573,In_1772);
and U2341 (N_2341,In_966,In_2732);
xnor U2342 (N_2342,In_1271,In_2375);
or U2343 (N_2343,In_4427,In_52);
or U2344 (N_2344,In_643,In_2751);
nor U2345 (N_2345,In_4270,In_4232);
and U2346 (N_2346,In_3545,In_3);
xor U2347 (N_2347,In_1916,In_3840);
nor U2348 (N_2348,In_1017,In_3587);
xor U2349 (N_2349,In_1697,In_2779);
nor U2350 (N_2350,In_101,In_2543);
nand U2351 (N_2351,In_2523,In_3007);
nor U2352 (N_2352,In_4048,In_866);
or U2353 (N_2353,In_2283,In_2940);
nand U2354 (N_2354,In_3697,In_366);
and U2355 (N_2355,In_1324,In_4405);
or U2356 (N_2356,In_4575,In_4426);
nor U2357 (N_2357,In_3539,In_1131);
xor U2358 (N_2358,In_3619,In_3233);
nand U2359 (N_2359,In_386,In_606);
nand U2360 (N_2360,In_4799,In_4794);
and U2361 (N_2361,In_3916,In_3092);
and U2362 (N_2362,In_445,In_3707);
and U2363 (N_2363,In_3565,In_508);
and U2364 (N_2364,In_2093,In_4028);
nand U2365 (N_2365,In_1486,In_2798);
and U2366 (N_2366,In_824,In_3393);
nor U2367 (N_2367,In_2269,In_3672);
or U2368 (N_2368,In_4432,In_4654);
and U2369 (N_2369,In_1720,In_3128);
nor U2370 (N_2370,In_3731,In_225);
nor U2371 (N_2371,In_252,In_1137);
and U2372 (N_2372,In_1750,In_877);
and U2373 (N_2373,In_3302,In_1644);
nor U2374 (N_2374,In_1873,In_3103);
nor U2375 (N_2375,In_813,In_555);
nor U2376 (N_2376,In_3999,In_613);
xor U2377 (N_2377,In_474,In_1156);
nor U2378 (N_2378,In_3511,In_3052);
and U2379 (N_2379,In_2756,In_1197);
or U2380 (N_2380,In_2542,In_2983);
nor U2381 (N_2381,In_4292,In_190);
and U2382 (N_2382,In_2825,In_4947);
nand U2383 (N_2383,In_733,In_3255);
nand U2384 (N_2384,In_4334,In_3191);
or U2385 (N_2385,In_4553,In_3793);
or U2386 (N_2386,In_842,In_3940);
nand U2387 (N_2387,In_3890,In_1532);
or U2388 (N_2388,In_1907,In_120);
and U2389 (N_2389,In_2545,In_3286);
nor U2390 (N_2390,In_3989,In_3717);
or U2391 (N_2391,In_1558,In_3018);
nor U2392 (N_2392,In_3796,In_4844);
nand U2393 (N_2393,In_4538,In_2486);
nand U2394 (N_2394,In_472,In_1316);
or U2395 (N_2395,In_2386,In_232);
nand U2396 (N_2396,In_2155,In_2980);
xor U2397 (N_2397,In_2664,In_4482);
nor U2398 (N_2398,In_3803,In_105);
and U2399 (N_2399,In_4886,In_3832);
nor U2400 (N_2400,In_387,In_1740);
nand U2401 (N_2401,In_3259,In_2103);
nand U2402 (N_2402,In_3857,In_4224);
nor U2403 (N_2403,In_4740,In_2215);
nor U2404 (N_2404,In_2083,In_1128);
or U2405 (N_2405,In_4634,In_2040);
or U2406 (N_2406,In_176,In_4449);
or U2407 (N_2407,In_1504,In_300);
nand U2408 (N_2408,In_4520,In_3129);
nor U2409 (N_2409,In_1737,In_1963);
or U2410 (N_2410,In_3814,In_2127);
nor U2411 (N_2411,In_260,In_1984);
nor U2412 (N_2412,In_1249,In_2865);
nand U2413 (N_2413,In_4973,In_45);
or U2414 (N_2414,In_1926,In_2169);
or U2415 (N_2415,In_2979,In_1473);
and U2416 (N_2416,In_2766,In_3458);
nand U2417 (N_2417,In_3461,In_4198);
xor U2418 (N_2418,In_85,In_3217);
and U2419 (N_2419,In_3820,In_4457);
nor U2420 (N_2420,In_4106,In_4999);
nor U2421 (N_2421,In_4568,In_3607);
nand U2422 (N_2422,In_4742,In_1095);
xor U2423 (N_2423,In_254,In_588);
nand U2424 (N_2424,In_2335,In_4780);
nor U2425 (N_2425,In_1666,In_4918);
or U2426 (N_2426,In_4307,In_2437);
xnor U2427 (N_2427,In_941,In_4289);
nand U2428 (N_2428,In_95,In_3181);
and U2429 (N_2429,In_1956,In_507);
and U2430 (N_2430,In_3344,In_2468);
xnor U2431 (N_2431,In_2029,In_243);
nor U2432 (N_2432,In_770,In_885);
and U2433 (N_2433,In_407,In_1707);
xnor U2434 (N_2434,In_177,In_1790);
and U2435 (N_2435,In_3269,In_998);
and U2436 (N_2436,In_837,In_3682);
nor U2437 (N_2437,In_608,In_571);
nor U2438 (N_2438,In_706,In_1050);
and U2439 (N_2439,In_2690,In_3237);
nand U2440 (N_2440,In_3781,In_4312);
or U2441 (N_2441,In_4981,In_1818);
and U2442 (N_2442,In_2956,In_3529);
and U2443 (N_2443,In_1002,In_3228);
nor U2444 (N_2444,In_3507,In_3521);
nor U2445 (N_2445,In_1799,In_3637);
nand U2446 (N_2446,In_2710,In_2482);
nor U2447 (N_2447,In_1683,In_869);
nand U2448 (N_2448,In_3190,In_404);
or U2449 (N_2449,In_4824,In_4474);
nor U2450 (N_2450,In_315,In_2809);
nand U2451 (N_2451,In_4069,In_237);
nand U2452 (N_2452,In_428,In_1225);
nor U2453 (N_2453,In_3264,In_4537);
and U2454 (N_2454,In_818,In_553);
or U2455 (N_2455,In_3411,In_4569);
and U2456 (N_2456,In_4113,In_1201);
or U2457 (N_2457,In_1257,In_2872);
and U2458 (N_2458,In_2499,In_1585);
or U2459 (N_2459,In_3131,In_1689);
nand U2460 (N_2460,In_4513,In_1912);
nor U2461 (N_2461,In_1361,In_2260);
nor U2462 (N_2462,In_2379,In_716);
or U2463 (N_2463,In_256,In_2781);
nand U2464 (N_2464,In_4668,In_1124);
and U2465 (N_2465,In_3398,In_1213);
and U2466 (N_2466,In_2547,In_3053);
and U2467 (N_2467,In_1533,In_4957);
and U2468 (N_2468,In_2042,In_4338);
or U2469 (N_2469,In_2564,In_4274);
and U2470 (N_2470,In_3045,In_1428);
xnor U2471 (N_2471,In_307,In_3726);
or U2472 (N_2472,In_43,In_940);
and U2473 (N_2473,In_4600,In_4171);
xor U2474 (N_2474,In_790,In_1688);
and U2475 (N_2475,In_3341,In_3541);
nor U2476 (N_2476,In_3669,In_2541);
or U2477 (N_2477,In_2941,In_2432);
and U2478 (N_2478,In_726,In_1908);
nand U2479 (N_2479,In_3512,In_4719);
and U2480 (N_2480,In_107,In_946);
nand U2481 (N_2481,In_3856,In_3852);
xnor U2482 (N_2482,In_1205,In_4593);
nor U2483 (N_2483,In_2658,In_4475);
nand U2484 (N_2484,In_2263,In_1312);
nand U2485 (N_2485,In_132,In_2306);
nand U2486 (N_2486,In_4500,In_3811);
nor U2487 (N_2487,In_4686,In_1592);
or U2488 (N_2488,In_4763,In_1842);
and U2489 (N_2489,In_1232,In_1162);
nand U2490 (N_2490,In_1957,In_4102);
nor U2491 (N_2491,In_3079,In_3349);
nor U2492 (N_2492,In_3605,In_628);
and U2493 (N_2493,In_823,In_58);
nor U2494 (N_2494,In_3095,In_3863);
or U2495 (N_2495,In_1538,In_4950);
or U2496 (N_2496,In_1521,In_1115);
nor U2497 (N_2497,In_1563,In_4506);
nand U2498 (N_2498,In_2660,In_545);
and U2499 (N_2499,In_3765,In_2087);
nand U2500 (N_2500,In_1143,In_1835);
and U2501 (N_2501,In_4444,In_2990);
and U2502 (N_2502,In_113,In_4911);
or U2503 (N_2503,In_4550,In_1924);
nand U2504 (N_2504,In_873,In_756);
nor U2505 (N_2505,In_1905,In_2578);
xnor U2506 (N_2506,In_2227,In_4926);
nand U2507 (N_2507,In_4142,In_4919);
xnor U2508 (N_2508,In_1170,In_1239);
nor U2509 (N_2509,In_1061,In_2177);
nor U2510 (N_2510,In_2717,In_971);
nor U2511 (N_2511,In_499,In_3825);
nor U2512 (N_2512,In_3461,In_882);
and U2513 (N_2513,In_3062,In_4942);
nand U2514 (N_2514,In_3215,In_4014);
nor U2515 (N_2515,In_3547,In_2804);
and U2516 (N_2516,In_4228,In_134);
and U2517 (N_2517,In_3423,In_4421);
and U2518 (N_2518,In_4963,In_436);
nor U2519 (N_2519,In_1372,In_310);
nor U2520 (N_2520,In_2894,In_2496);
and U2521 (N_2521,In_4685,In_2439);
or U2522 (N_2522,In_1066,In_4194);
nor U2523 (N_2523,In_2876,In_2630);
or U2524 (N_2524,In_2354,In_411);
nor U2525 (N_2525,In_1007,In_3880);
and U2526 (N_2526,In_2765,In_3382);
nor U2527 (N_2527,In_2551,In_3625);
nor U2528 (N_2528,In_2165,In_3106);
nor U2529 (N_2529,In_2258,In_3895);
nor U2530 (N_2530,In_2471,In_247);
and U2531 (N_2531,In_3517,In_4678);
nor U2532 (N_2532,In_164,In_351);
and U2533 (N_2533,In_628,In_4107);
and U2534 (N_2534,In_1138,In_855);
and U2535 (N_2535,In_3262,In_2297);
nor U2536 (N_2536,In_147,In_742);
or U2537 (N_2537,In_231,In_308);
xnor U2538 (N_2538,In_3768,In_4351);
and U2539 (N_2539,In_414,In_1860);
nor U2540 (N_2540,In_2860,In_3770);
or U2541 (N_2541,In_1508,In_4289);
and U2542 (N_2542,In_3224,In_618);
and U2543 (N_2543,In_226,In_3615);
nand U2544 (N_2544,In_2144,In_1433);
and U2545 (N_2545,In_4203,In_1105);
nand U2546 (N_2546,In_1210,In_2303);
and U2547 (N_2547,In_2249,In_2526);
and U2548 (N_2548,In_4553,In_2779);
xnor U2549 (N_2549,In_1764,In_2998);
nand U2550 (N_2550,In_506,In_175);
and U2551 (N_2551,In_433,In_1860);
or U2552 (N_2552,In_1491,In_2824);
nor U2553 (N_2553,In_4743,In_4720);
and U2554 (N_2554,In_1870,In_1645);
and U2555 (N_2555,In_2663,In_1544);
xnor U2556 (N_2556,In_3367,In_749);
nor U2557 (N_2557,In_669,In_4581);
xnor U2558 (N_2558,In_3028,In_1732);
xnor U2559 (N_2559,In_2582,In_1367);
xor U2560 (N_2560,In_2102,In_4593);
nor U2561 (N_2561,In_4142,In_3627);
and U2562 (N_2562,In_1423,In_1817);
nor U2563 (N_2563,In_3385,In_1122);
or U2564 (N_2564,In_943,In_4498);
nor U2565 (N_2565,In_994,In_2722);
nor U2566 (N_2566,In_3127,In_1191);
nand U2567 (N_2567,In_2409,In_1951);
or U2568 (N_2568,In_4698,In_1891);
or U2569 (N_2569,In_3095,In_4548);
nor U2570 (N_2570,In_2900,In_3203);
nand U2571 (N_2571,In_2787,In_265);
nand U2572 (N_2572,In_3850,In_2499);
nand U2573 (N_2573,In_4282,In_954);
xor U2574 (N_2574,In_4841,In_347);
and U2575 (N_2575,In_1417,In_2339);
nand U2576 (N_2576,In_1400,In_4982);
and U2577 (N_2577,In_1327,In_2494);
or U2578 (N_2578,In_1070,In_4619);
and U2579 (N_2579,In_60,In_160);
or U2580 (N_2580,In_1995,In_495);
nor U2581 (N_2581,In_4658,In_1792);
nor U2582 (N_2582,In_4312,In_3052);
nor U2583 (N_2583,In_295,In_100);
xnor U2584 (N_2584,In_215,In_3492);
nor U2585 (N_2585,In_2173,In_1581);
or U2586 (N_2586,In_3243,In_3461);
and U2587 (N_2587,In_120,In_1249);
or U2588 (N_2588,In_2604,In_4712);
nor U2589 (N_2589,In_104,In_313);
xor U2590 (N_2590,In_4830,In_3674);
and U2591 (N_2591,In_3648,In_3093);
nand U2592 (N_2592,In_306,In_3688);
or U2593 (N_2593,In_4016,In_2657);
nand U2594 (N_2594,In_335,In_1715);
nor U2595 (N_2595,In_2302,In_3861);
or U2596 (N_2596,In_2117,In_3664);
nor U2597 (N_2597,In_2090,In_1468);
or U2598 (N_2598,In_1823,In_1532);
or U2599 (N_2599,In_1274,In_2892);
nor U2600 (N_2600,In_2547,In_1305);
or U2601 (N_2601,In_601,In_2572);
nor U2602 (N_2602,In_1135,In_1555);
or U2603 (N_2603,In_1945,In_2174);
and U2604 (N_2604,In_4672,In_3191);
nand U2605 (N_2605,In_132,In_4176);
and U2606 (N_2606,In_2735,In_4799);
or U2607 (N_2607,In_1144,In_3659);
or U2608 (N_2608,In_3660,In_4903);
nor U2609 (N_2609,In_1027,In_1989);
nand U2610 (N_2610,In_3167,In_4200);
nand U2611 (N_2611,In_3294,In_2778);
and U2612 (N_2612,In_4459,In_2798);
nor U2613 (N_2613,In_3742,In_2482);
or U2614 (N_2614,In_72,In_1793);
nand U2615 (N_2615,In_1225,In_4982);
or U2616 (N_2616,In_2952,In_1448);
or U2617 (N_2617,In_1953,In_1107);
and U2618 (N_2618,In_3937,In_4747);
nand U2619 (N_2619,In_2371,In_2991);
nor U2620 (N_2620,In_3811,In_3384);
and U2621 (N_2621,In_2673,In_1387);
and U2622 (N_2622,In_3105,In_3286);
and U2623 (N_2623,In_1722,In_1152);
nand U2624 (N_2624,In_2821,In_1606);
and U2625 (N_2625,In_4580,In_2277);
and U2626 (N_2626,In_4294,In_832);
or U2627 (N_2627,In_1920,In_1294);
or U2628 (N_2628,In_4921,In_4736);
or U2629 (N_2629,In_3942,In_1687);
xnor U2630 (N_2630,In_3275,In_2808);
nand U2631 (N_2631,In_3911,In_3660);
or U2632 (N_2632,In_2567,In_754);
nor U2633 (N_2633,In_1458,In_789);
xnor U2634 (N_2634,In_110,In_714);
nand U2635 (N_2635,In_4924,In_4783);
or U2636 (N_2636,In_4006,In_1207);
nor U2637 (N_2637,In_3226,In_4038);
or U2638 (N_2638,In_4965,In_118);
nor U2639 (N_2639,In_3400,In_2113);
nand U2640 (N_2640,In_3814,In_3119);
nor U2641 (N_2641,In_1811,In_1050);
or U2642 (N_2642,In_3171,In_4787);
nand U2643 (N_2643,In_3299,In_2691);
nor U2644 (N_2644,In_3264,In_741);
and U2645 (N_2645,In_1975,In_274);
nand U2646 (N_2646,In_166,In_1598);
and U2647 (N_2647,In_2063,In_2350);
nand U2648 (N_2648,In_3972,In_3309);
and U2649 (N_2649,In_3992,In_2588);
and U2650 (N_2650,In_131,In_4919);
and U2651 (N_2651,In_2567,In_4822);
or U2652 (N_2652,In_4083,In_147);
and U2653 (N_2653,In_315,In_3608);
nor U2654 (N_2654,In_954,In_4649);
or U2655 (N_2655,In_1502,In_2919);
nand U2656 (N_2656,In_411,In_3160);
and U2657 (N_2657,In_2349,In_2197);
nor U2658 (N_2658,In_850,In_4740);
xnor U2659 (N_2659,In_2196,In_8);
nor U2660 (N_2660,In_958,In_2894);
and U2661 (N_2661,In_2691,In_3748);
nand U2662 (N_2662,In_1568,In_2671);
nor U2663 (N_2663,In_894,In_4541);
nand U2664 (N_2664,In_2051,In_3012);
nand U2665 (N_2665,In_1579,In_910);
xor U2666 (N_2666,In_3731,In_1094);
xnor U2667 (N_2667,In_4317,In_2439);
or U2668 (N_2668,In_178,In_4209);
or U2669 (N_2669,In_3143,In_4926);
or U2670 (N_2670,In_235,In_909);
and U2671 (N_2671,In_1672,In_2877);
and U2672 (N_2672,In_1315,In_3421);
or U2673 (N_2673,In_1299,In_4242);
xor U2674 (N_2674,In_4703,In_1408);
or U2675 (N_2675,In_1314,In_2840);
nand U2676 (N_2676,In_2969,In_2352);
nor U2677 (N_2677,In_396,In_2689);
or U2678 (N_2678,In_2804,In_3059);
nor U2679 (N_2679,In_4458,In_4784);
nor U2680 (N_2680,In_2177,In_535);
xnor U2681 (N_2681,In_2735,In_3148);
nand U2682 (N_2682,In_2007,In_4617);
and U2683 (N_2683,In_1360,In_2820);
nor U2684 (N_2684,In_3226,In_2295);
xor U2685 (N_2685,In_2054,In_3590);
or U2686 (N_2686,In_2276,In_2394);
nor U2687 (N_2687,In_71,In_718);
or U2688 (N_2688,In_4209,In_397);
or U2689 (N_2689,In_1449,In_721);
and U2690 (N_2690,In_133,In_1169);
and U2691 (N_2691,In_2128,In_2302);
xnor U2692 (N_2692,In_282,In_293);
nand U2693 (N_2693,In_4319,In_2777);
nand U2694 (N_2694,In_4922,In_1680);
and U2695 (N_2695,In_1858,In_617);
and U2696 (N_2696,In_1074,In_2956);
nor U2697 (N_2697,In_1847,In_2177);
or U2698 (N_2698,In_2841,In_669);
and U2699 (N_2699,In_2666,In_3902);
and U2700 (N_2700,In_4193,In_4149);
nand U2701 (N_2701,In_202,In_4126);
nand U2702 (N_2702,In_4820,In_1955);
and U2703 (N_2703,In_2169,In_1484);
nand U2704 (N_2704,In_3245,In_3264);
xnor U2705 (N_2705,In_4329,In_3014);
xor U2706 (N_2706,In_4448,In_3055);
and U2707 (N_2707,In_1531,In_1400);
nor U2708 (N_2708,In_641,In_3677);
and U2709 (N_2709,In_19,In_1303);
nand U2710 (N_2710,In_4572,In_2329);
nor U2711 (N_2711,In_3851,In_3550);
xor U2712 (N_2712,In_821,In_2076);
and U2713 (N_2713,In_1425,In_264);
and U2714 (N_2714,In_1495,In_818);
xnor U2715 (N_2715,In_4228,In_2032);
nand U2716 (N_2716,In_2134,In_3378);
or U2717 (N_2717,In_4536,In_4022);
xnor U2718 (N_2718,In_3780,In_7);
nand U2719 (N_2719,In_1378,In_3882);
nand U2720 (N_2720,In_667,In_3062);
or U2721 (N_2721,In_2601,In_300);
or U2722 (N_2722,In_389,In_4278);
xor U2723 (N_2723,In_630,In_1619);
or U2724 (N_2724,In_1603,In_77);
or U2725 (N_2725,In_947,In_1587);
nor U2726 (N_2726,In_2769,In_1620);
nand U2727 (N_2727,In_4848,In_4286);
or U2728 (N_2728,In_4184,In_4085);
xnor U2729 (N_2729,In_1879,In_797);
and U2730 (N_2730,In_4288,In_2699);
or U2731 (N_2731,In_2450,In_3821);
or U2732 (N_2732,In_2321,In_4153);
and U2733 (N_2733,In_1530,In_825);
and U2734 (N_2734,In_334,In_3188);
nand U2735 (N_2735,In_1636,In_4227);
nor U2736 (N_2736,In_889,In_325);
nor U2737 (N_2737,In_134,In_731);
nor U2738 (N_2738,In_439,In_2874);
and U2739 (N_2739,In_2015,In_4323);
nor U2740 (N_2740,In_937,In_1557);
xnor U2741 (N_2741,In_1831,In_2376);
nor U2742 (N_2742,In_3112,In_2520);
nor U2743 (N_2743,In_1359,In_3858);
nand U2744 (N_2744,In_647,In_3074);
nand U2745 (N_2745,In_1582,In_3104);
or U2746 (N_2746,In_3542,In_3884);
xor U2747 (N_2747,In_2626,In_1423);
nand U2748 (N_2748,In_1959,In_1350);
nor U2749 (N_2749,In_3267,In_4162);
nor U2750 (N_2750,In_830,In_4409);
and U2751 (N_2751,In_585,In_2453);
nand U2752 (N_2752,In_3813,In_3203);
or U2753 (N_2753,In_4486,In_568);
nand U2754 (N_2754,In_4841,In_3772);
and U2755 (N_2755,In_3466,In_2635);
nand U2756 (N_2756,In_2498,In_1767);
and U2757 (N_2757,In_3910,In_4416);
and U2758 (N_2758,In_1397,In_4183);
xor U2759 (N_2759,In_1223,In_1326);
and U2760 (N_2760,In_639,In_3153);
nand U2761 (N_2761,In_3481,In_2294);
nor U2762 (N_2762,In_1706,In_4419);
and U2763 (N_2763,In_1595,In_966);
nand U2764 (N_2764,In_3067,In_3383);
and U2765 (N_2765,In_3970,In_3919);
and U2766 (N_2766,In_92,In_212);
and U2767 (N_2767,In_3742,In_3693);
nor U2768 (N_2768,In_4760,In_1027);
or U2769 (N_2769,In_300,In_1323);
and U2770 (N_2770,In_4136,In_3614);
or U2771 (N_2771,In_1452,In_3393);
or U2772 (N_2772,In_1262,In_1992);
or U2773 (N_2773,In_3566,In_712);
xnor U2774 (N_2774,In_1203,In_3290);
nand U2775 (N_2775,In_1693,In_1743);
nand U2776 (N_2776,In_1435,In_3586);
or U2777 (N_2777,In_3371,In_475);
or U2778 (N_2778,In_731,In_2558);
and U2779 (N_2779,In_1665,In_3392);
nand U2780 (N_2780,In_4699,In_3242);
and U2781 (N_2781,In_4393,In_3551);
xor U2782 (N_2782,In_3704,In_4988);
and U2783 (N_2783,In_4887,In_2005);
nor U2784 (N_2784,In_411,In_3425);
nor U2785 (N_2785,In_1192,In_2568);
and U2786 (N_2786,In_2216,In_2431);
or U2787 (N_2787,In_2918,In_1743);
nor U2788 (N_2788,In_2721,In_1823);
xor U2789 (N_2789,In_2141,In_1519);
and U2790 (N_2790,In_4733,In_2872);
or U2791 (N_2791,In_4691,In_1170);
and U2792 (N_2792,In_3748,In_1293);
nand U2793 (N_2793,In_2912,In_432);
nor U2794 (N_2794,In_2275,In_1985);
nand U2795 (N_2795,In_3543,In_3996);
nand U2796 (N_2796,In_3570,In_327);
and U2797 (N_2797,In_4974,In_4072);
nand U2798 (N_2798,In_307,In_1972);
xnor U2799 (N_2799,In_1678,In_3434);
and U2800 (N_2800,In_100,In_4922);
nor U2801 (N_2801,In_3647,In_3839);
xor U2802 (N_2802,In_1794,In_472);
or U2803 (N_2803,In_3368,In_3327);
or U2804 (N_2804,In_2588,In_217);
and U2805 (N_2805,In_740,In_3011);
nand U2806 (N_2806,In_1523,In_2505);
and U2807 (N_2807,In_1040,In_2562);
nor U2808 (N_2808,In_734,In_2218);
nor U2809 (N_2809,In_2431,In_4029);
nand U2810 (N_2810,In_4651,In_3672);
or U2811 (N_2811,In_2158,In_4239);
xnor U2812 (N_2812,In_3210,In_1527);
or U2813 (N_2813,In_3749,In_2781);
or U2814 (N_2814,In_4736,In_4547);
or U2815 (N_2815,In_1104,In_14);
nand U2816 (N_2816,In_1645,In_1144);
and U2817 (N_2817,In_472,In_2538);
or U2818 (N_2818,In_712,In_815);
or U2819 (N_2819,In_4287,In_2209);
nand U2820 (N_2820,In_3200,In_304);
and U2821 (N_2821,In_908,In_4213);
or U2822 (N_2822,In_49,In_2581);
nand U2823 (N_2823,In_3320,In_4697);
or U2824 (N_2824,In_658,In_3456);
nand U2825 (N_2825,In_1558,In_2608);
or U2826 (N_2826,In_1912,In_3062);
xor U2827 (N_2827,In_80,In_1824);
xnor U2828 (N_2828,In_985,In_3914);
nor U2829 (N_2829,In_921,In_0);
xor U2830 (N_2830,In_1014,In_2485);
xnor U2831 (N_2831,In_4935,In_3115);
nand U2832 (N_2832,In_3618,In_3014);
nor U2833 (N_2833,In_523,In_3629);
or U2834 (N_2834,In_2929,In_1381);
nand U2835 (N_2835,In_4629,In_1814);
xor U2836 (N_2836,In_2456,In_4340);
and U2837 (N_2837,In_2032,In_1647);
xor U2838 (N_2838,In_4392,In_2253);
or U2839 (N_2839,In_578,In_1667);
nor U2840 (N_2840,In_3614,In_3960);
and U2841 (N_2841,In_573,In_4866);
nand U2842 (N_2842,In_4472,In_2684);
nand U2843 (N_2843,In_3485,In_2849);
and U2844 (N_2844,In_1933,In_3711);
and U2845 (N_2845,In_3072,In_4550);
and U2846 (N_2846,In_185,In_1040);
nand U2847 (N_2847,In_1933,In_2972);
xnor U2848 (N_2848,In_2299,In_1430);
and U2849 (N_2849,In_3392,In_2359);
or U2850 (N_2850,In_1730,In_49);
nor U2851 (N_2851,In_4932,In_4546);
nor U2852 (N_2852,In_4367,In_2142);
nand U2853 (N_2853,In_3537,In_405);
and U2854 (N_2854,In_2335,In_3871);
xnor U2855 (N_2855,In_2532,In_3919);
nor U2856 (N_2856,In_4230,In_2833);
and U2857 (N_2857,In_3525,In_1174);
nand U2858 (N_2858,In_2389,In_4171);
nor U2859 (N_2859,In_3320,In_4427);
nor U2860 (N_2860,In_2172,In_1827);
nor U2861 (N_2861,In_2259,In_1332);
and U2862 (N_2862,In_3176,In_2157);
or U2863 (N_2863,In_1119,In_2853);
nor U2864 (N_2864,In_2056,In_1385);
xor U2865 (N_2865,In_3853,In_1806);
nor U2866 (N_2866,In_86,In_2856);
nor U2867 (N_2867,In_2675,In_573);
and U2868 (N_2868,In_4818,In_4672);
xor U2869 (N_2869,In_2285,In_1210);
and U2870 (N_2870,In_3241,In_4880);
nor U2871 (N_2871,In_3934,In_441);
nand U2872 (N_2872,In_1160,In_988);
and U2873 (N_2873,In_2308,In_431);
nor U2874 (N_2874,In_468,In_1022);
nor U2875 (N_2875,In_1522,In_1470);
and U2876 (N_2876,In_4913,In_1357);
nand U2877 (N_2877,In_1245,In_2485);
or U2878 (N_2878,In_1061,In_312);
or U2879 (N_2879,In_1696,In_2099);
nor U2880 (N_2880,In_4333,In_2574);
nand U2881 (N_2881,In_4363,In_4);
nor U2882 (N_2882,In_2193,In_1878);
and U2883 (N_2883,In_3678,In_1072);
nor U2884 (N_2884,In_3388,In_1761);
nor U2885 (N_2885,In_55,In_540);
nor U2886 (N_2886,In_1626,In_4724);
nor U2887 (N_2887,In_2689,In_2292);
or U2888 (N_2888,In_1298,In_128);
nand U2889 (N_2889,In_27,In_2402);
or U2890 (N_2890,In_2408,In_1881);
nand U2891 (N_2891,In_2990,In_3927);
and U2892 (N_2892,In_4570,In_4272);
nor U2893 (N_2893,In_3412,In_1353);
nor U2894 (N_2894,In_2194,In_1876);
and U2895 (N_2895,In_2599,In_450);
or U2896 (N_2896,In_4616,In_1046);
and U2897 (N_2897,In_1298,In_2770);
nand U2898 (N_2898,In_809,In_1469);
nor U2899 (N_2899,In_215,In_1078);
or U2900 (N_2900,In_1666,In_3937);
nor U2901 (N_2901,In_949,In_3166);
or U2902 (N_2902,In_2683,In_4187);
nand U2903 (N_2903,In_3867,In_4643);
and U2904 (N_2904,In_3102,In_2183);
xnor U2905 (N_2905,In_3225,In_573);
nand U2906 (N_2906,In_2612,In_2001);
or U2907 (N_2907,In_3326,In_4879);
and U2908 (N_2908,In_273,In_4565);
nor U2909 (N_2909,In_2349,In_2462);
nor U2910 (N_2910,In_79,In_4141);
and U2911 (N_2911,In_390,In_4421);
nor U2912 (N_2912,In_4768,In_4537);
nor U2913 (N_2913,In_936,In_2225);
xnor U2914 (N_2914,In_2324,In_3554);
and U2915 (N_2915,In_1629,In_2407);
nor U2916 (N_2916,In_889,In_875);
xnor U2917 (N_2917,In_2963,In_3550);
or U2918 (N_2918,In_778,In_1994);
nor U2919 (N_2919,In_2746,In_2997);
and U2920 (N_2920,In_1261,In_4425);
nor U2921 (N_2921,In_228,In_3114);
nand U2922 (N_2922,In_4617,In_282);
or U2923 (N_2923,In_1483,In_44);
nor U2924 (N_2924,In_4648,In_4169);
nor U2925 (N_2925,In_3335,In_1493);
nand U2926 (N_2926,In_229,In_4630);
nor U2927 (N_2927,In_3817,In_1898);
or U2928 (N_2928,In_1107,In_2796);
nand U2929 (N_2929,In_1137,In_423);
and U2930 (N_2930,In_4559,In_4414);
xnor U2931 (N_2931,In_1690,In_3248);
nor U2932 (N_2932,In_2837,In_1601);
or U2933 (N_2933,In_3541,In_4322);
and U2934 (N_2934,In_1957,In_3023);
nand U2935 (N_2935,In_970,In_1299);
or U2936 (N_2936,In_3460,In_4714);
and U2937 (N_2937,In_3366,In_1811);
nand U2938 (N_2938,In_3723,In_4494);
xnor U2939 (N_2939,In_117,In_3148);
nor U2940 (N_2940,In_2147,In_181);
nand U2941 (N_2941,In_3842,In_632);
nand U2942 (N_2942,In_1128,In_4353);
xor U2943 (N_2943,In_4199,In_4603);
nor U2944 (N_2944,In_2895,In_3852);
or U2945 (N_2945,In_4383,In_3464);
or U2946 (N_2946,In_3311,In_373);
nand U2947 (N_2947,In_5,In_2279);
xor U2948 (N_2948,In_2027,In_2231);
nor U2949 (N_2949,In_3168,In_4049);
xnor U2950 (N_2950,In_3537,In_802);
or U2951 (N_2951,In_1508,In_1597);
and U2952 (N_2952,In_936,In_2387);
nor U2953 (N_2953,In_2078,In_2964);
nand U2954 (N_2954,In_209,In_3555);
nand U2955 (N_2955,In_2914,In_2815);
xor U2956 (N_2956,In_1327,In_2786);
or U2957 (N_2957,In_4411,In_1258);
nand U2958 (N_2958,In_2763,In_407);
or U2959 (N_2959,In_161,In_2783);
or U2960 (N_2960,In_2936,In_1857);
nor U2961 (N_2961,In_2709,In_1019);
nor U2962 (N_2962,In_1068,In_1274);
xnor U2963 (N_2963,In_63,In_1988);
and U2964 (N_2964,In_819,In_3327);
nand U2965 (N_2965,In_4008,In_478);
and U2966 (N_2966,In_250,In_4940);
nand U2967 (N_2967,In_152,In_4869);
or U2968 (N_2968,In_4674,In_2965);
nand U2969 (N_2969,In_4554,In_3313);
or U2970 (N_2970,In_2649,In_2198);
xnor U2971 (N_2971,In_1701,In_2635);
or U2972 (N_2972,In_1224,In_632);
nor U2973 (N_2973,In_2740,In_796);
xor U2974 (N_2974,In_4752,In_2820);
nor U2975 (N_2975,In_489,In_3340);
and U2976 (N_2976,In_447,In_2972);
nand U2977 (N_2977,In_1392,In_2541);
and U2978 (N_2978,In_4353,In_216);
nor U2979 (N_2979,In_2817,In_4051);
xor U2980 (N_2980,In_4086,In_2845);
nor U2981 (N_2981,In_644,In_2592);
nand U2982 (N_2982,In_438,In_3826);
or U2983 (N_2983,In_4707,In_4026);
or U2984 (N_2984,In_1569,In_2868);
or U2985 (N_2985,In_2170,In_2142);
and U2986 (N_2986,In_821,In_1972);
nor U2987 (N_2987,In_1734,In_2483);
xnor U2988 (N_2988,In_1844,In_499);
and U2989 (N_2989,In_1096,In_4081);
or U2990 (N_2990,In_3308,In_4642);
nand U2991 (N_2991,In_4100,In_44);
or U2992 (N_2992,In_4938,In_3651);
nor U2993 (N_2993,In_1829,In_1364);
nand U2994 (N_2994,In_244,In_804);
nor U2995 (N_2995,In_2702,In_1639);
nand U2996 (N_2996,In_2771,In_3187);
or U2997 (N_2997,In_455,In_3647);
or U2998 (N_2998,In_2514,In_586);
and U2999 (N_2999,In_1604,In_2181);
nand U3000 (N_3000,In_4427,In_4340);
and U3001 (N_3001,In_1203,In_4437);
nand U3002 (N_3002,In_330,In_791);
nor U3003 (N_3003,In_3024,In_207);
and U3004 (N_3004,In_4398,In_979);
or U3005 (N_3005,In_1827,In_2932);
nand U3006 (N_3006,In_599,In_2164);
and U3007 (N_3007,In_4553,In_505);
nor U3008 (N_3008,In_1433,In_2258);
or U3009 (N_3009,In_3846,In_2942);
and U3010 (N_3010,In_936,In_3585);
or U3011 (N_3011,In_3922,In_4480);
and U3012 (N_3012,In_4952,In_2340);
xor U3013 (N_3013,In_1417,In_2679);
xor U3014 (N_3014,In_331,In_4788);
nand U3015 (N_3015,In_4454,In_2188);
nor U3016 (N_3016,In_3554,In_4166);
nor U3017 (N_3017,In_877,In_3623);
and U3018 (N_3018,In_4922,In_3259);
or U3019 (N_3019,In_2686,In_4495);
nor U3020 (N_3020,In_3935,In_764);
nor U3021 (N_3021,In_3226,In_524);
nor U3022 (N_3022,In_2918,In_1202);
or U3023 (N_3023,In_3273,In_934);
and U3024 (N_3024,In_1868,In_2489);
nor U3025 (N_3025,In_4715,In_495);
xor U3026 (N_3026,In_1490,In_2455);
and U3027 (N_3027,In_3416,In_505);
nor U3028 (N_3028,In_139,In_2844);
and U3029 (N_3029,In_3148,In_651);
or U3030 (N_3030,In_3998,In_1519);
nand U3031 (N_3031,In_132,In_2328);
xor U3032 (N_3032,In_1831,In_1095);
nor U3033 (N_3033,In_3591,In_1817);
nor U3034 (N_3034,In_3311,In_965);
nand U3035 (N_3035,In_8,In_2662);
nand U3036 (N_3036,In_137,In_2209);
and U3037 (N_3037,In_2610,In_493);
and U3038 (N_3038,In_3281,In_1122);
and U3039 (N_3039,In_1286,In_4044);
nand U3040 (N_3040,In_3817,In_2681);
xnor U3041 (N_3041,In_865,In_1646);
nor U3042 (N_3042,In_4752,In_1782);
and U3043 (N_3043,In_4674,In_1053);
nand U3044 (N_3044,In_3592,In_3018);
and U3045 (N_3045,In_2418,In_88);
or U3046 (N_3046,In_4072,In_2857);
nand U3047 (N_3047,In_2805,In_1415);
xor U3048 (N_3048,In_3706,In_1161);
nand U3049 (N_3049,In_1121,In_310);
or U3050 (N_3050,In_4274,In_719);
and U3051 (N_3051,In_3935,In_1373);
nor U3052 (N_3052,In_32,In_3431);
nand U3053 (N_3053,In_2878,In_2244);
or U3054 (N_3054,In_4840,In_4895);
or U3055 (N_3055,In_4372,In_4291);
nand U3056 (N_3056,In_377,In_3638);
nand U3057 (N_3057,In_1983,In_3228);
or U3058 (N_3058,In_4554,In_3802);
or U3059 (N_3059,In_3169,In_4225);
nor U3060 (N_3060,In_3863,In_2348);
nor U3061 (N_3061,In_75,In_148);
or U3062 (N_3062,In_2631,In_522);
or U3063 (N_3063,In_833,In_601);
nor U3064 (N_3064,In_1071,In_2478);
or U3065 (N_3065,In_3119,In_1526);
and U3066 (N_3066,In_4896,In_4768);
nand U3067 (N_3067,In_1151,In_2616);
nand U3068 (N_3068,In_3844,In_424);
and U3069 (N_3069,In_3582,In_176);
nand U3070 (N_3070,In_3607,In_203);
and U3071 (N_3071,In_1847,In_3507);
or U3072 (N_3072,In_3199,In_4746);
or U3073 (N_3073,In_2849,In_4745);
or U3074 (N_3074,In_4258,In_157);
or U3075 (N_3075,In_1958,In_2863);
or U3076 (N_3076,In_2254,In_3569);
and U3077 (N_3077,In_3044,In_1200);
or U3078 (N_3078,In_2513,In_3294);
nor U3079 (N_3079,In_902,In_2766);
xor U3080 (N_3080,In_2871,In_2025);
or U3081 (N_3081,In_4147,In_940);
nand U3082 (N_3082,In_2564,In_2532);
and U3083 (N_3083,In_1695,In_2414);
nor U3084 (N_3084,In_3103,In_4559);
nor U3085 (N_3085,In_4555,In_4228);
and U3086 (N_3086,In_4608,In_3963);
nor U3087 (N_3087,In_138,In_1741);
nand U3088 (N_3088,In_3172,In_1123);
or U3089 (N_3089,In_205,In_4544);
or U3090 (N_3090,In_4456,In_4731);
or U3091 (N_3091,In_33,In_495);
nand U3092 (N_3092,In_1292,In_893);
nor U3093 (N_3093,In_1135,In_2428);
and U3094 (N_3094,In_4446,In_60);
nand U3095 (N_3095,In_4390,In_2344);
or U3096 (N_3096,In_4508,In_1873);
and U3097 (N_3097,In_1814,In_1367);
and U3098 (N_3098,In_1708,In_2863);
nand U3099 (N_3099,In_2699,In_2611);
and U3100 (N_3100,In_4895,In_3300);
and U3101 (N_3101,In_3447,In_3718);
and U3102 (N_3102,In_107,In_3607);
nand U3103 (N_3103,In_3171,In_2467);
nor U3104 (N_3104,In_3217,In_2652);
xnor U3105 (N_3105,In_2003,In_4670);
xor U3106 (N_3106,In_4835,In_189);
nand U3107 (N_3107,In_126,In_917);
xnor U3108 (N_3108,In_1541,In_4576);
xor U3109 (N_3109,In_1654,In_1768);
nor U3110 (N_3110,In_885,In_397);
xor U3111 (N_3111,In_3539,In_432);
or U3112 (N_3112,In_4017,In_1979);
nand U3113 (N_3113,In_4775,In_2356);
and U3114 (N_3114,In_3912,In_3072);
nor U3115 (N_3115,In_4242,In_4502);
and U3116 (N_3116,In_4487,In_2542);
nor U3117 (N_3117,In_646,In_1347);
or U3118 (N_3118,In_4647,In_3616);
nor U3119 (N_3119,In_3107,In_1402);
nand U3120 (N_3120,In_3473,In_2673);
and U3121 (N_3121,In_4988,In_2162);
nor U3122 (N_3122,In_4422,In_658);
or U3123 (N_3123,In_2225,In_1836);
and U3124 (N_3124,In_2935,In_822);
and U3125 (N_3125,In_4143,In_2328);
or U3126 (N_3126,In_4876,In_2283);
or U3127 (N_3127,In_396,In_4283);
xnor U3128 (N_3128,In_809,In_3282);
xor U3129 (N_3129,In_4855,In_4754);
and U3130 (N_3130,In_4226,In_2097);
or U3131 (N_3131,In_1095,In_3880);
xnor U3132 (N_3132,In_2901,In_1323);
or U3133 (N_3133,In_3564,In_1658);
and U3134 (N_3134,In_2086,In_3731);
nand U3135 (N_3135,In_3094,In_1957);
nor U3136 (N_3136,In_991,In_1301);
nor U3137 (N_3137,In_2232,In_681);
or U3138 (N_3138,In_1771,In_4591);
and U3139 (N_3139,In_2501,In_2428);
nand U3140 (N_3140,In_1914,In_1327);
and U3141 (N_3141,In_1648,In_4);
and U3142 (N_3142,In_2752,In_1411);
nand U3143 (N_3143,In_4275,In_2333);
or U3144 (N_3144,In_4211,In_3765);
or U3145 (N_3145,In_3920,In_1832);
or U3146 (N_3146,In_4372,In_2442);
or U3147 (N_3147,In_498,In_4796);
nor U3148 (N_3148,In_1376,In_1824);
nor U3149 (N_3149,In_2269,In_3979);
nor U3150 (N_3150,In_332,In_3040);
xnor U3151 (N_3151,In_3387,In_581);
or U3152 (N_3152,In_2474,In_1559);
nor U3153 (N_3153,In_1896,In_2633);
nand U3154 (N_3154,In_3596,In_624);
nand U3155 (N_3155,In_3365,In_801);
and U3156 (N_3156,In_484,In_4067);
xor U3157 (N_3157,In_3660,In_2844);
nand U3158 (N_3158,In_4459,In_252);
nand U3159 (N_3159,In_2304,In_1425);
nand U3160 (N_3160,In_1051,In_1880);
nand U3161 (N_3161,In_593,In_3308);
nor U3162 (N_3162,In_1601,In_180);
nand U3163 (N_3163,In_1143,In_2387);
nor U3164 (N_3164,In_292,In_4136);
xnor U3165 (N_3165,In_4924,In_3441);
and U3166 (N_3166,In_64,In_4972);
xnor U3167 (N_3167,In_214,In_1179);
nor U3168 (N_3168,In_2395,In_2904);
nand U3169 (N_3169,In_2943,In_1949);
nand U3170 (N_3170,In_4978,In_4151);
or U3171 (N_3171,In_2037,In_1775);
xor U3172 (N_3172,In_342,In_3985);
xnor U3173 (N_3173,In_3110,In_875);
nor U3174 (N_3174,In_4672,In_3904);
and U3175 (N_3175,In_341,In_4884);
nor U3176 (N_3176,In_1846,In_660);
nor U3177 (N_3177,In_2895,In_3791);
and U3178 (N_3178,In_1818,In_1159);
and U3179 (N_3179,In_1128,In_3887);
and U3180 (N_3180,In_3818,In_2793);
nor U3181 (N_3181,In_2886,In_302);
and U3182 (N_3182,In_4732,In_3492);
nand U3183 (N_3183,In_2486,In_414);
nand U3184 (N_3184,In_2305,In_4503);
and U3185 (N_3185,In_1870,In_1270);
nor U3186 (N_3186,In_4944,In_2765);
xnor U3187 (N_3187,In_2849,In_1714);
or U3188 (N_3188,In_548,In_3369);
nor U3189 (N_3189,In_2288,In_627);
nand U3190 (N_3190,In_1345,In_19);
xnor U3191 (N_3191,In_1721,In_1506);
xnor U3192 (N_3192,In_3118,In_3235);
and U3193 (N_3193,In_2747,In_931);
or U3194 (N_3194,In_4734,In_1422);
and U3195 (N_3195,In_3278,In_2518);
nand U3196 (N_3196,In_531,In_582);
or U3197 (N_3197,In_3579,In_2375);
and U3198 (N_3198,In_4871,In_4141);
and U3199 (N_3199,In_4288,In_394);
and U3200 (N_3200,In_1367,In_2958);
or U3201 (N_3201,In_3425,In_4066);
nor U3202 (N_3202,In_3009,In_23);
nor U3203 (N_3203,In_623,In_2751);
and U3204 (N_3204,In_4817,In_932);
nor U3205 (N_3205,In_1211,In_474);
nor U3206 (N_3206,In_1427,In_289);
or U3207 (N_3207,In_1675,In_3783);
or U3208 (N_3208,In_2610,In_2374);
nor U3209 (N_3209,In_3721,In_3239);
and U3210 (N_3210,In_1868,In_1893);
or U3211 (N_3211,In_651,In_1940);
xor U3212 (N_3212,In_1599,In_4258);
nor U3213 (N_3213,In_3310,In_3517);
nand U3214 (N_3214,In_3434,In_343);
nand U3215 (N_3215,In_4991,In_4667);
nor U3216 (N_3216,In_4583,In_2919);
nor U3217 (N_3217,In_243,In_694);
or U3218 (N_3218,In_3259,In_4224);
or U3219 (N_3219,In_4351,In_4683);
or U3220 (N_3220,In_3704,In_3213);
nand U3221 (N_3221,In_2884,In_1700);
nand U3222 (N_3222,In_2002,In_838);
and U3223 (N_3223,In_2494,In_4273);
and U3224 (N_3224,In_4087,In_2864);
nand U3225 (N_3225,In_2415,In_96);
nand U3226 (N_3226,In_124,In_4269);
xnor U3227 (N_3227,In_982,In_2955);
and U3228 (N_3228,In_94,In_3584);
or U3229 (N_3229,In_1661,In_4429);
or U3230 (N_3230,In_4470,In_4600);
nor U3231 (N_3231,In_3906,In_4414);
nand U3232 (N_3232,In_1165,In_819);
and U3233 (N_3233,In_3881,In_2305);
nor U3234 (N_3234,In_1877,In_731);
nand U3235 (N_3235,In_3801,In_557);
nand U3236 (N_3236,In_2582,In_2304);
nor U3237 (N_3237,In_4765,In_634);
xor U3238 (N_3238,In_3910,In_4690);
or U3239 (N_3239,In_4812,In_506);
or U3240 (N_3240,In_2022,In_2208);
and U3241 (N_3241,In_2054,In_1159);
nor U3242 (N_3242,In_439,In_2711);
nand U3243 (N_3243,In_1758,In_1470);
and U3244 (N_3244,In_3507,In_2196);
nand U3245 (N_3245,In_1140,In_14);
nor U3246 (N_3246,In_2570,In_86);
and U3247 (N_3247,In_4532,In_1254);
nand U3248 (N_3248,In_4187,In_395);
xor U3249 (N_3249,In_1005,In_4050);
nand U3250 (N_3250,In_1977,In_169);
and U3251 (N_3251,In_4474,In_1439);
nand U3252 (N_3252,In_4521,In_1334);
or U3253 (N_3253,In_565,In_3204);
and U3254 (N_3254,In_971,In_533);
nand U3255 (N_3255,In_10,In_4417);
or U3256 (N_3256,In_2540,In_170);
nor U3257 (N_3257,In_609,In_605);
nor U3258 (N_3258,In_194,In_2825);
nor U3259 (N_3259,In_2494,In_4651);
nand U3260 (N_3260,In_4643,In_1164);
nand U3261 (N_3261,In_696,In_1126);
and U3262 (N_3262,In_4970,In_259);
nand U3263 (N_3263,In_3559,In_3890);
or U3264 (N_3264,In_767,In_991);
nand U3265 (N_3265,In_4232,In_2859);
and U3266 (N_3266,In_758,In_2371);
or U3267 (N_3267,In_568,In_4290);
xor U3268 (N_3268,In_2166,In_2952);
and U3269 (N_3269,In_2463,In_4674);
xor U3270 (N_3270,In_4734,In_1516);
or U3271 (N_3271,In_2055,In_3070);
and U3272 (N_3272,In_3207,In_3674);
or U3273 (N_3273,In_1498,In_1205);
nor U3274 (N_3274,In_2625,In_2906);
nand U3275 (N_3275,In_3547,In_2363);
and U3276 (N_3276,In_4859,In_2715);
nor U3277 (N_3277,In_4886,In_2266);
nand U3278 (N_3278,In_1935,In_383);
xor U3279 (N_3279,In_3177,In_1438);
or U3280 (N_3280,In_914,In_438);
or U3281 (N_3281,In_1355,In_2727);
nand U3282 (N_3282,In_132,In_2397);
nand U3283 (N_3283,In_904,In_3840);
or U3284 (N_3284,In_4726,In_473);
xnor U3285 (N_3285,In_2499,In_399);
nor U3286 (N_3286,In_1679,In_47);
xnor U3287 (N_3287,In_3688,In_4524);
nand U3288 (N_3288,In_3865,In_3202);
and U3289 (N_3289,In_3915,In_1696);
nand U3290 (N_3290,In_2436,In_4794);
or U3291 (N_3291,In_3129,In_2550);
or U3292 (N_3292,In_1527,In_651);
nand U3293 (N_3293,In_1461,In_2784);
and U3294 (N_3294,In_826,In_564);
or U3295 (N_3295,In_3104,In_3176);
nor U3296 (N_3296,In_38,In_2750);
nor U3297 (N_3297,In_68,In_4475);
nand U3298 (N_3298,In_1562,In_4362);
nand U3299 (N_3299,In_4343,In_877);
xnor U3300 (N_3300,In_2534,In_1682);
xor U3301 (N_3301,In_4508,In_3100);
nor U3302 (N_3302,In_4168,In_2753);
nand U3303 (N_3303,In_4472,In_2563);
and U3304 (N_3304,In_2419,In_4917);
nand U3305 (N_3305,In_4000,In_77);
nand U3306 (N_3306,In_2872,In_4525);
or U3307 (N_3307,In_4248,In_4817);
xnor U3308 (N_3308,In_993,In_350);
or U3309 (N_3309,In_681,In_1336);
nor U3310 (N_3310,In_3402,In_411);
nand U3311 (N_3311,In_1387,In_2617);
or U3312 (N_3312,In_4214,In_69);
xnor U3313 (N_3313,In_1426,In_1231);
nand U3314 (N_3314,In_1015,In_655);
xor U3315 (N_3315,In_2236,In_2712);
or U3316 (N_3316,In_2825,In_4939);
or U3317 (N_3317,In_676,In_3969);
and U3318 (N_3318,In_1012,In_100);
nor U3319 (N_3319,In_3543,In_1937);
or U3320 (N_3320,In_1064,In_1825);
nand U3321 (N_3321,In_4071,In_1617);
xnor U3322 (N_3322,In_2144,In_2320);
or U3323 (N_3323,In_1744,In_4075);
and U3324 (N_3324,In_4259,In_3020);
or U3325 (N_3325,In_3069,In_1138);
nor U3326 (N_3326,In_3147,In_4164);
nand U3327 (N_3327,In_4887,In_1370);
nor U3328 (N_3328,In_569,In_1063);
xnor U3329 (N_3329,In_4469,In_252);
xor U3330 (N_3330,In_3191,In_2060);
nor U3331 (N_3331,In_365,In_4921);
nor U3332 (N_3332,In_1218,In_4546);
nand U3333 (N_3333,In_791,In_3284);
nor U3334 (N_3334,In_935,In_767);
and U3335 (N_3335,In_917,In_110);
or U3336 (N_3336,In_2623,In_3586);
nor U3337 (N_3337,In_2466,In_1092);
and U3338 (N_3338,In_2680,In_435);
nand U3339 (N_3339,In_566,In_4700);
and U3340 (N_3340,In_3538,In_328);
nand U3341 (N_3341,In_3230,In_3042);
nand U3342 (N_3342,In_2513,In_1945);
xnor U3343 (N_3343,In_1221,In_1047);
nand U3344 (N_3344,In_992,In_3917);
xor U3345 (N_3345,In_1594,In_571);
xnor U3346 (N_3346,In_4560,In_3603);
or U3347 (N_3347,In_4577,In_502);
and U3348 (N_3348,In_1171,In_3193);
and U3349 (N_3349,In_1997,In_4165);
nand U3350 (N_3350,In_3736,In_1336);
and U3351 (N_3351,In_140,In_4857);
nand U3352 (N_3352,In_1808,In_1703);
nand U3353 (N_3353,In_1271,In_3784);
nand U3354 (N_3354,In_939,In_3576);
nor U3355 (N_3355,In_77,In_3180);
nor U3356 (N_3356,In_2451,In_4785);
nand U3357 (N_3357,In_367,In_2185);
and U3358 (N_3358,In_1991,In_1134);
nor U3359 (N_3359,In_2863,In_2597);
xnor U3360 (N_3360,In_1582,In_4479);
and U3361 (N_3361,In_1962,In_2179);
nand U3362 (N_3362,In_4159,In_663);
and U3363 (N_3363,In_2671,In_3174);
nor U3364 (N_3364,In_4122,In_3970);
nand U3365 (N_3365,In_1370,In_4696);
nor U3366 (N_3366,In_4315,In_4359);
or U3367 (N_3367,In_3132,In_3790);
xor U3368 (N_3368,In_1238,In_4124);
xor U3369 (N_3369,In_1866,In_4131);
xnor U3370 (N_3370,In_4311,In_1202);
and U3371 (N_3371,In_4679,In_4717);
and U3372 (N_3372,In_4749,In_2122);
and U3373 (N_3373,In_4718,In_3302);
nor U3374 (N_3374,In_4385,In_343);
nand U3375 (N_3375,In_4870,In_2661);
nand U3376 (N_3376,In_2539,In_1969);
nor U3377 (N_3377,In_4447,In_2174);
nand U3378 (N_3378,In_3544,In_2572);
nand U3379 (N_3379,In_2197,In_4549);
and U3380 (N_3380,In_4580,In_749);
nor U3381 (N_3381,In_4750,In_1499);
or U3382 (N_3382,In_4246,In_1571);
nand U3383 (N_3383,In_3112,In_1218);
or U3384 (N_3384,In_2076,In_3799);
and U3385 (N_3385,In_129,In_586);
or U3386 (N_3386,In_1827,In_1962);
nand U3387 (N_3387,In_3132,In_4520);
nor U3388 (N_3388,In_2265,In_3570);
nor U3389 (N_3389,In_4972,In_4549);
nand U3390 (N_3390,In_3110,In_697);
nor U3391 (N_3391,In_1699,In_2201);
nor U3392 (N_3392,In_1214,In_2753);
and U3393 (N_3393,In_1118,In_1871);
nor U3394 (N_3394,In_4393,In_2675);
and U3395 (N_3395,In_4985,In_4063);
or U3396 (N_3396,In_912,In_294);
xor U3397 (N_3397,In_3479,In_4224);
or U3398 (N_3398,In_4367,In_2202);
and U3399 (N_3399,In_333,In_2408);
or U3400 (N_3400,In_569,In_3860);
nor U3401 (N_3401,In_2655,In_2442);
nand U3402 (N_3402,In_3765,In_3392);
and U3403 (N_3403,In_4661,In_4912);
nand U3404 (N_3404,In_2571,In_1634);
nand U3405 (N_3405,In_2190,In_4952);
nor U3406 (N_3406,In_2322,In_1650);
nand U3407 (N_3407,In_976,In_3867);
nor U3408 (N_3408,In_4844,In_4850);
nor U3409 (N_3409,In_2241,In_1706);
or U3410 (N_3410,In_2087,In_617);
nor U3411 (N_3411,In_2361,In_4656);
xnor U3412 (N_3412,In_321,In_4847);
xor U3413 (N_3413,In_4984,In_2995);
nor U3414 (N_3414,In_2933,In_392);
and U3415 (N_3415,In_1377,In_1850);
and U3416 (N_3416,In_2504,In_1798);
nor U3417 (N_3417,In_1218,In_4572);
and U3418 (N_3418,In_2803,In_1762);
or U3419 (N_3419,In_2900,In_1708);
nand U3420 (N_3420,In_1934,In_4205);
nor U3421 (N_3421,In_4053,In_3673);
or U3422 (N_3422,In_1553,In_4641);
nand U3423 (N_3423,In_3292,In_3029);
and U3424 (N_3424,In_3433,In_2151);
or U3425 (N_3425,In_1037,In_2784);
nand U3426 (N_3426,In_260,In_564);
nor U3427 (N_3427,In_698,In_949);
nand U3428 (N_3428,In_1786,In_661);
nor U3429 (N_3429,In_894,In_1351);
xor U3430 (N_3430,In_56,In_1617);
or U3431 (N_3431,In_1578,In_3760);
nand U3432 (N_3432,In_3889,In_4339);
or U3433 (N_3433,In_2873,In_3526);
or U3434 (N_3434,In_2674,In_3934);
nor U3435 (N_3435,In_4016,In_1111);
xor U3436 (N_3436,In_1275,In_3397);
and U3437 (N_3437,In_1305,In_1330);
nor U3438 (N_3438,In_3012,In_3847);
nand U3439 (N_3439,In_4127,In_3835);
nand U3440 (N_3440,In_3009,In_1349);
nand U3441 (N_3441,In_558,In_1935);
nand U3442 (N_3442,In_863,In_3382);
nor U3443 (N_3443,In_179,In_4212);
nor U3444 (N_3444,In_2177,In_4717);
and U3445 (N_3445,In_2063,In_424);
nand U3446 (N_3446,In_1985,In_4769);
xor U3447 (N_3447,In_962,In_3275);
and U3448 (N_3448,In_3904,In_4226);
nor U3449 (N_3449,In_4508,In_3124);
nand U3450 (N_3450,In_3476,In_1099);
or U3451 (N_3451,In_2884,In_571);
nand U3452 (N_3452,In_4257,In_1339);
xor U3453 (N_3453,In_0,In_2440);
nand U3454 (N_3454,In_2729,In_3111);
and U3455 (N_3455,In_3330,In_597);
or U3456 (N_3456,In_2004,In_3444);
nand U3457 (N_3457,In_4211,In_2884);
and U3458 (N_3458,In_4284,In_875);
and U3459 (N_3459,In_2695,In_3895);
nor U3460 (N_3460,In_4673,In_3896);
nor U3461 (N_3461,In_4817,In_1122);
nand U3462 (N_3462,In_3592,In_197);
xor U3463 (N_3463,In_4473,In_298);
or U3464 (N_3464,In_3702,In_4374);
and U3465 (N_3465,In_2043,In_4853);
nor U3466 (N_3466,In_3012,In_4349);
or U3467 (N_3467,In_2651,In_2272);
or U3468 (N_3468,In_4059,In_3869);
and U3469 (N_3469,In_3156,In_4940);
nand U3470 (N_3470,In_4323,In_614);
and U3471 (N_3471,In_3439,In_499);
nor U3472 (N_3472,In_457,In_2543);
nand U3473 (N_3473,In_1400,In_1948);
nor U3474 (N_3474,In_436,In_4792);
or U3475 (N_3475,In_2514,In_348);
nand U3476 (N_3476,In_4344,In_3390);
or U3477 (N_3477,In_1516,In_4844);
nor U3478 (N_3478,In_315,In_2236);
or U3479 (N_3479,In_2950,In_3042);
and U3480 (N_3480,In_3362,In_4447);
and U3481 (N_3481,In_71,In_1772);
nor U3482 (N_3482,In_1598,In_960);
and U3483 (N_3483,In_1638,In_4538);
and U3484 (N_3484,In_4998,In_4209);
and U3485 (N_3485,In_4038,In_4328);
nor U3486 (N_3486,In_4131,In_3724);
nor U3487 (N_3487,In_1133,In_144);
or U3488 (N_3488,In_824,In_2016);
and U3489 (N_3489,In_2354,In_1907);
xor U3490 (N_3490,In_4693,In_3767);
nand U3491 (N_3491,In_827,In_646);
nand U3492 (N_3492,In_4801,In_4557);
or U3493 (N_3493,In_3050,In_497);
nor U3494 (N_3494,In_1270,In_1086);
nor U3495 (N_3495,In_3069,In_2408);
or U3496 (N_3496,In_20,In_288);
or U3497 (N_3497,In_3175,In_4221);
or U3498 (N_3498,In_3166,In_775);
nand U3499 (N_3499,In_171,In_79);
nor U3500 (N_3500,In_2549,In_2667);
or U3501 (N_3501,In_4107,In_3975);
or U3502 (N_3502,In_3685,In_4994);
nand U3503 (N_3503,In_3539,In_4542);
nand U3504 (N_3504,In_3843,In_2854);
xnor U3505 (N_3505,In_2629,In_2146);
and U3506 (N_3506,In_1200,In_4655);
nand U3507 (N_3507,In_1323,In_3909);
nand U3508 (N_3508,In_2454,In_2788);
and U3509 (N_3509,In_690,In_2981);
nand U3510 (N_3510,In_1153,In_2416);
nor U3511 (N_3511,In_987,In_3705);
and U3512 (N_3512,In_3460,In_3431);
nand U3513 (N_3513,In_3808,In_15);
nand U3514 (N_3514,In_4727,In_4944);
nand U3515 (N_3515,In_712,In_1596);
nor U3516 (N_3516,In_2843,In_947);
nor U3517 (N_3517,In_4828,In_1885);
nor U3518 (N_3518,In_631,In_1143);
nand U3519 (N_3519,In_4422,In_3125);
xnor U3520 (N_3520,In_1392,In_4808);
nand U3521 (N_3521,In_81,In_3143);
nand U3522 (N_3522,In_1850,In_1317);
nor U3523 (N_3523,In_2789,In_1148);
nand U3524 (N_3524,In_2319,In_4715);
or U3525 (N_3525,In_2392,In_3956);
nor U3526 (N_3526,In_4853,In_3096);
nor U3527 (N_3527,In_1053,In_3843);
nand U3528 (N_3528,In_1672,In_1867);
and U3529 (N_3529,In_2021,In_4838);
xnor U3530 (N_3530,In_199,In_4448);
nor U3531 (N_3531,In_2824,In_4522);
or U3532 (N_3532,In_404,In_1668);
nand U3533 (N_3533,In_1118,In_3570);
and U3534 (N_3534,In_4879,In_4818);
nor U3535 (N_3535,In_2895,In_4213);
and U3536 (N_3536,In_4088,In_2993);
nand U3537 (N_3537,In_2634,In_1696);
nor U3538 (N_3538,In_4309,In_3329);
and U3539 (N_3539,In_3951,In_587);
nor U3540 (N_3540,In_2622,In_4957);
nor U3541 (N_3541,In_30,In_2156);
nand U3542 (N_3542,In_4692,In_4464);
or U3543 (N_3543,In_413,In_1408);
nand U3544 (N_3544,In_787,In_3703);
or U3545 (N_3545,In_4952,In_2349);
nand U3546 (N_3546,In_2512,In_3938);
nor U3547 (N_3547,In_3435,In_460);
and U3548 (N_3548,In_1385,In_4952);
or U3549 (N_3549,In_4392,In_2593);
nor U3550 (N_3550,In_1612,In_3209);
nand U3551 (N_3551,In_4147,In_461);
or U3552 (N_3552,In_4338,In_3420);
nand U3553 (N_3553,In_3104,In_883);
nand U3554 (N_3554,In_1438,In_4170);
nand U3555 (N_3555,In_2437,In_3565);
or U3556 (N_3556,In_4223,In_4053);
or U3557 (N_3557,In_4979,In_4429);
and U3558 (N_3558,In_2360,In_4999);
nand U3559 (N_3559,In_3652,In_4921);
xnor U3560 (N_3560,In_1694,In_685);
or U3561 (N_3561,In_424,In_2521);
or U3562 (N_3562,In_528,In_420);
and U3563 (N_3563,In_3142,In_1083);
nor U3564 (N_3564,In_4135,In_914);
xnor U3565 (N_3565,In_1611,In_2185);
nand U3566 (N_3566,In_3866,In_1645);
nand U3567 (N_3567,In_2666,In_463);
nor U3568 (N_3568,In_3210,In_2442);
nand U3569 (N_3569,In_4785,In_4491);
and U3570 (N_3570,In_3780,In_1376);
and U3571 (N_3571,In_1353,In_2806);
and U3572 (N_3572,In_1214,In_2725);
or U3573 (N_3573,In_3548,In_364);
or U3574 (N_3574,In_680,In_2685);
nand U3575 (N_3575,In_4392,In_4000);
nand U3576 (N_3576,In_2863,In_4199);
nor U3577 (N_3577,In_3980,In_4027);
xor U3578 (N_3578,In_3859,In_1766);
nand U3579 (N_3579,In_1266,In_344);
and U3580 (N_3580,In_3183,In_1121);
nand U3581 (N_3581,In_4390,In_2850);
and U3582 (N_3582,In_1572,In_4453);
and U3583 (N_3583,In_3202,In_1261);
nor U3584 (N_3584,In_532,In_341);
nor U3585 (N_3585,In_3017,In_4597);
nor U3586 (N_3586,In_397,In_3031);
or U3587 (N_3587,In_4164,In_4967);
and U3588 (N_3588,In_1084,In_2039);
or U3589 (N_3589,In_3545,In_2416);
nand U3590 (N_3590,In_3255,In_4375);
nor U3591 (N_3591,In_911,In_4067);
nor U3592 (N_3592,In_1229,In_4409);
and U3593 (N_3593,In_4340,In_1118);
nand U3594 (N_3594,In_3582,In_4488);
or U3595 (N_3595,In_743,In_4035);
and U3596 (N_3596,In_1151,In_2592);
and U3597 (N_3597,In_2668,In_4040);
nand U3598 (N_3598,In_1689,In_4535);
or U3599 (N_3599,In_3714,In_3479);
and U3600 (N_3600,In_982,In_279);
nor U3601 (N_3601,In_4576,In_1611);
nor U3602 (N_3602,In_3735,In_691);
nand U3603 (N_3603,In_4150,In_1144);
nor U3604 (N_3604,In_2156,In_2923);
or U3605 (N_3605,In_498,In_470);
nor U3606 (N_3606,In_3060,In_1974);
nor U3607 (N_3607,In_3444,In_767);
nor U3608 (N_3608,In_974,In_4612);
or U3609 (N_3609,In_488,In_1439);
and U3610 (N_3610,In_4907,In_4497);
and U3611 (N_3611,In_712,In_4804);
or U3612 (N_3612,In_2319,In_4029);
and U3613 (N_3613,In_179,In_851);
and U3614 (N_3614,In_4511,In_4506);
nor U3615 (N_3615,In_783,In_1538);
and U3616 (N_3616,In_215,In_966);
and U3617 (N_3617,In_782,In_4020);
or U3618 (N_3618,In_2769,In_1806);
and U3619 (N_3619,In_3986,In_2835);
nor U3620 (N_3620,In_1465,In_2944);
and U3621 (N_3621,In_794,In_1101);
nor U3622 (N_3622,In_4611,In_1645);
xor U3623 (N_3623,In_1531,In_641);
and U3624 (N_3624,In_2588,In_2248);
nor U3625 (N_3625,In_2013,In_3284);
nand U3626 (N_3626,In_831,In_552);
and U3627 (N_3627,In_1090,In_236);
nand U3628 (N_3628,In_2190,In_2260);
and U3629 (N_3629,In_913,In_536);
nand U3630 (N_3630,In_1156,In_3782);
and U3631 (N_3631,In_1518,In_4260);
nand U3632 (N_3632,In_4505,In_4046);
or U3633 (N_3633,In_1135,In_1203);
nand U3634 (N_3634,In_4380,In_4041);
nand U3635 (N_3635,In_3793,In_4965);
or U3636 (N_3636,In_4312,In_234);
nor U3637 (N_3637,In_3701,In_2031);
and U3638 (N_3638,In_4062,In_3108);
nor U3639 (N_3639,In_4478,In_3026);
xor U3640 (N_3640,In_388,In_4761);
and U3641 (N_3641,In_4104,In_2234);
or U3642 (N_3642,In_279,In_1655);
nor U3643 (N_3643,In_4931,In_3330);
or U3644 (N_3644,In_4156,In_3368);
nor U3645 (N_3645,In_4341,In_1093);
or U3646 (N_3646,In_4222,In_4593);
or U3647 (N_3647,In_3974,In_3223);
and U3648 (N_3648,In_674,In_3897);
nor U3649 (N_3649,In_802,In_1588);
and U3650 (N_3650,In_4873,In_1563);
or U3651 (N_3651,In_3353,In_1890);
nand U3652 (N_3652,In_1077,In_2232);
nand U3653 (N_3653,In_4886,In_1043);
nor U3654 (N_3654,In_4333,In_4808);
nor U3655 (N_3655,In_3467,In_4295);
nor U3656 (N_3656,In_4356,In_1212);
or U3657 (N_3657,In_4878,In_2006);
nor U3658 (N_3658,In_3923,In_3484);
and U3659 (N_3659,In_3859,In_1146);
and U3660 (N_3660,In_2753,In_2370);
nand U3661 (N_3661,In_498,In_3137);
or U3662 (N_3662,In_4777,In_4540);
xnor U3663 (N_3663,In_913,In_1594);
nand U3664 (N_3664,In_3324,In_4425);
or U3665 (N_3665,In_3017,In_72);
and U3666 (N_3666,In_3578,In_2389);
nor U3667 (N_3667,In_2288,In_132);
nand U3668 (N_3668,In_2897,In_4132);
nand U3669 (N_3669,In_49,In_1070);
nor U3670 (N_3670,In_167,In_1408);
and U3671 (N_3671,In_1929,In_3388);
or U3672 (N_3672,In_4706,In_4143);
and U3673 (N_3673,In_4031,In_510);
nand U3674 (N_3674,In_1333,In_1471);
nor U3675 (N_3675,In_3425,In_928);
or U3676 (N_3676,In_3549,In_332);
nor U3677 (N_3677,In_4022,In_48);
or U3678 (N_3678,In_2034,In_1769);
or U3679 (N_3679,In_3280,In_4338);
and U3680 (N_3680,In_3486,In_1114);
nand U3681 (N_3681,In_3977,In_1139);
and U3682 (N_3682,In_2158,In_1627);
and U3683 (N_3683,In_1742,In_1784);
nand U3684 (N_3684,In_4023,In_996);
or U3685 (N_3685,In_2790,In_3397);
nor U3686 (N_3686,In_3787,In_2638);
and U3687 (N_3687,In_1241,In_3905);
or U3688 (N_3688,In_3777,In_525);
and U3689 (N_3689,In_2381,In_1491);
and U3690 (N_3690,In_4997,In_3288);
and U3691 (N_3691,In_4503,In_2949);
or U3692 (N_3692,In_2377,In_2794);
nand U3693 (N_3693,In_1389,In_4020);
nor U3694 (N_3694,In_3886,In_4753);
nand U3695 (N_3695,In_1284,In_4110);
and U3696 (N_3696,In_413,In_748);
nor U3697 (N_3697,In_2870,In_1182);
and U3698 (N_3698,In_4173,In_2286);
xnor U3699 (N_3699,In_4409,In_4264);
or U3700 (N_3700,In_48,In_4035);
xnor U3701 (N_3701,In_268,In_2694);
and U3702 (N_3702,In_4161,In_2908);
or U3703 (N_3703,In_3399,In_2630);
and U3704 (N_3704,In_3920,In_3191);
nand U3705 (N_3705,In_1790,In_685);
nand U3706 (N_3706,In_3802,In_3887);
and U3707 (N_3707,In_446,In_4338);
and U3708 (N_3708,In_1214,In_4593);
or U3709 (N_3709,In_1082,In_4931);
nor U3710 (N_3710,In_1357,In_1272);
nand U3711 (N_3711,In_984,In_3198);
or U3712 (N_3712,In_3240,In_1443);
nor U3713 (N_3713,In_2272,In_1924);
xnor U3714 (N_3714,In_4070,In_4294);
xnor U3715 (N_3715,In_4374,In_603);
nand U3716 (N_3716,In_4294,In_2011);
nand U3717 (N_3717,In_2358,In_105);
nand U3718 (N_3718,In_2564,In_3625);
and U3719 (N_3719,In_272,In_4154);
and U3720 (N_3720,In_4936,In_3928);
or U3721 (N_3721,In_1486,In_2613);
or U3722 (N_3722,In_559,In_695);
nand U3723 (N_3723,In_971,In_4362);
nand U3724 (N_3724,In_1195,In_3476);
nor U3725 (N_3725,In_1690,In_2107);
nor U3726 (N_3726,In_4089,In_1744);
nor U3727 (N_3727,In_2295,In_85);
nand U3728 (N_3728,In_4811,In_4489);
or U3729 (N_3729,In_2649,In_4241);
nand U3730 (N_3730,In_4743,In_1812);
or U3731 (N_3731,In_3332,In_1109);
nand U3732 (N_3732,In_2411,In_3242);
nor U3733 (N_3733,In_1115,In_2909);
and U3734 (N_3734,In_1978,In_4538);
nand U3735 (N_3735,In_2989,In_3693);
or U3736 (N_3736,In_2012,In_4288);
and U3737 (N_3737,In_235,In_1033);
xnor U3738 (N_3738,In_1790,In_1260);
xnor U3739 (N_3739,In_858,In_1177);
nand U3740 (N_3740,In_3169,In_2642);
nor U3741 (N_3741,In_2753,In_3817);
xor U3742 (N_3742,In_863,In_3122);
nor U3743 (N_3743,In_2792,In_1939);
nand U3744 (N_3744,In_2777,In_3663);
nor U3745 (N_3745,In_135,In_1425);
nand U3746 (N_3746,In_796,In_3486);
and U3747 (N_3747,In_2920,In_4279);
or U3748 (N_3748,In_4283,In_2698);
and U3749 (N_3749,In_3554,In_1656);
or U3750 (N_3750,In_1048,In_4995);
nand U3751 (N_3751,In_4876,In_851);
nand U3752 (N_3752,In_949,In_4424);
nor U3753 (N_3753,In_2363,In_4196);
xnor U3754 (N_3754,In_4868,In_863);
nor U3755 (N_3755,In_674,In_1437);
nor U3756 (N_3756,In_3539,In_796);
nor U3757 (N_3757,In_4295,In_1352);
or U3758 (N_3758,In_4004,In_2403);
nor U3759 (N_3759,In_4884,In_833);
and U3760 (N_3760,In_1512,In_2823);
and U3761 (N_3761,In_4761,In_3943);
or U3762 (N_3762,In_4935,In_2672);
and U3763 (N_3763,In_3224,In_2875);
or U3764 (N_3764,In_3554,In_4771);
nand U3765 (N_3765,In_321,In_3121);
xor U3766 (N_3766,In_770,In_2218);
or U3767 (N_3767,In_3203,In_1542);
xor U3768 (N_3768,In_3710,In_3782);
nor U3769 (N_3769,In_4132,In_2553);
and U3770 (N_3770,In_4673,In_4844);
and U3771 (N_3771,In_3947,In_2093);
nor U3772 (N_3772,In_3505,In_2143);
and U3773 (N_3773,In_9,In_1552);
nor U3774 (N_3774,In_393,In_4893);
nand U3775 (N_3775,In_4281,In_1681);
and U3776 (N_3776,In_4901,In_1131);
xor U3777 (N_3777,In_467,In_3654);
nor U3778 (N_3778,In_4474,In_4016);
nor U3779 (N_3779,In_4785,In_4181);
nand U3780 (N_3780,In_1953,In_839);
nor U3781 (N_3781,In_1027,In_4726);
or U3782 (N_3782,In_3134,In_889);
or U3783 (N_3783,In_4267,In_162);
xor U3784 (N_3784,In_2254,In_4111);
nor U3785 (N_3785,In_3813,In_4022);
xnor U3786 (N_3786,In_2466,In_2884);
nor U3787 (N_3787,In_1756,In_963);
nand U3788 (N_3788,In_4506,In_4510);
nand U3789 (N_3789,In_4984,In_2550);
and U3790 (N_3790,In_2287,In_1449);
nand U3791 (N_3791,In_2996,In_2007);
or U3792 (N_3792,In_1855,In_1598);
nor U3793 (N_3793,In_2242,In_4741);
nor U3794 (N_3794,In_3659,In_4592);
or U3795 (N_3795,In_1838,In_2299);
nor U3796 (N_3796,In_641,In_4526);
nand U3797 (N_3797,In_2489,In_4378);
and U3798 (N_3798,In_4176,In_1281);
and U3799 (N_3799,In_2067,In_336);
and U3800 (N_3800,In_1195,In_2867);
nand U3801 (N_3801,In_3184,In_4893);
or U3802 (N_3802,In_3946,In_4914);
nand U3803 (N_3803,In_2122,In_4326);
and U3804 (N_3804,In_1814,In_2567);
nor U3805 (N_3805,In_4948,In_1916);
nand U3806 (N_3806,In_3076,In_3884);
nor U3807 (N_3807,In_928,In_4987);
nor U3808 (N_3808,In_2505,In_3262);
nand U3809 (N_3809,In_4048,In_3343);
or U3810 (N_3810,In_3981,In_2540);
and U3811 (N_3811,In_1435,In_4044);
and U3812 (N_3812,In_3609,In_4369);
nor U3813 (N_3813,In_4537,In_1709);
or U3814 (N_3814,In_3168,In_870);
or U3815 (N_3815,In_1923,In_3583);
nor U3816 (N_3816,In_4749,In_1135);
nor U3817 (N_3817,In_652,In_2971);
nand U3818 (N_3818,In_780,In_3138);
or U3819 (N_3819,In_4493,In_860);
or U3820 (N_3820,In_3467,In_1662);
and U3821 (N_3821,In_4041,In_4846);
or U3822 (N_3822,In_4248,In_513);
and U3823 (N_3823,In_473,In_3527);
and U3824 (N_3824,In_26,In_1435);
nor U3825 (N_3825,In_4065,In_60);
nand U3826 (N_3826,In_3005,In_4364);
nor U3827 (N_3827,In_2302,In_2138);
nor U3828 (N_3828,In_4853,In_3972);
nand U3829 (N_3829,In_2888,In_3514);
nor U3830 (N_3830,In_1559,In_2055);
nand U3831 (N_3831,In_4215,In_1547);
nand U3832 (N_3832,In_1101,In_965);
or U3833 (N_3833,In_2801,In_101);
or U3834 (N_3834,In_4620,In_3488);
and U3835 (N_3835,In_4266,In_317);
nor U3836 (N_3836,In_3015,In_4189);
and U3837 (N_3837,In_685,In_1784);
nand U3838 (N_3838,In_1160,In_3200);
nand U3839 (N_3839,In_3658,In_4160);
nand U3840 (N_3840,In_2025,In_4001);
or U3841 (N_3841,In_624,In_150);
and U3842 (N_3842,In_604,In_2133);
or U3843 (N_3843,In_4308,In_2309);
nor U3844 (N_3844,In_1091,In_3110);
xnor U3845 (N_3845,In_1044,In_143);
nand U3846 (N_3846,In_1702,In_3605);
and U3847 (N_3847,In_711,In_2098);
xor U3848 (N_3848,In_546,In_3684);
nand U3849 (N_3849,In_376,In_3143);
nor U3850 (N_3850,In_348,In_1364);
xor U3851 (N_3851,In_2551,In_2049);
nor U3852 (N_3852,In_668,In_1982);
nor U3853 (N_3853,In_526,In_2641);
nand U3854 (N_3854,In_148,In_4945);
xnor U3855 (N_3855,In_3804,In_33);
and U3856 (N_3856,In_2660,In_1674);
and U3857 (N_3857,In_4560,In_2418);
or U3858 (N_3858,In_4513,In_1842);
and U3859 (N_3859,In_834,In_2730);
and U3860 (N_3860,In_3458,In_781);
and U3861 (N_3861,In_1862,In_2215);
nor U3862 (N_3862,In_2731,In_3193);
xnor U3863 (N_3863,In_242,In_3031);
nand U3864 (N_3864,In_3746,In_3404);
nor U3865 (N_3865,In_2880,In_4607);
xnor U3866 (N_3866,In_3339,In_394);
nor U3867 (N_3867,In_3644,In_4307);
xor U3868 (N_3868,In_1045,In_3713);
nand U3869 (N_3869,In_3202,In_1214);
nor U3870 (N_3870,In_757,In_4202);
and U3871 (N_3871,In_4440,In_4495);
and U3872 (N_3872,In_2492,In_4552);
nor U3873 (N_3873,In_288,In_2942);
and U3874 (N_3874,In_2660,In_3536);
nor U3875 (N_3875,In_2268,In_388);
nand U3876 (N_3876,In_4188,In_4954);
nand U3877 (N_3877,In_3695,In_1771);
nand U3878 (N_3878,In_3061,In_3638);
or U3879 (N_3879,In_824,In_1392);
and U3880 (N_3880,In_2341,In_1664);
nor U3881 (N_3881,In_4880,In_2005);
and U3882 (N_3882,In_1697,In_1686);
and U3883 (N_3883,In_2934,In_779);
and U3884 (N_3884,In_588,In_2413);
and U3885 (N_3885,In_1587,In_1386);
and U3886 (N_3886,In_3516,In_3459);
or U3887 (N_3887,In_2351,In_2935);
or U3888 (N_3888,In_236,In_2532);
nand U3889 (N_3889,In_3199,In_3203);
or U3890 (N_3890,In_2518,In_2667);
and U3891 (N_3891,In_289,In_551);
or U3892 (N_3892,In_2062,In_2939);
nor U3893 (N_3893,In_4100,In_1410);
nand U3894 (N_3894,In_421,In_922);
and U3895 (N_3895,In_2318,In_3711);
nand U3896 (N_3896,In_4595,In_1570);
nor U3897 (N_3897,In_1123,In_4788);
nor U3898 (N_3898,In_1164,In_3517);
and U3899 (N_3899,In_4642,In_2077);
nand U3900 (N_3900,In_2229,In_836);
nor U3901 (N_3901,In_2031,In_4489);
or U3902 (N_3902,In_3342,In_3423);
nor U3903 (N_3903,In_1137,In_2536);
or U3904 (N_3904,In_3665,In_3010);
nor U3905 (N_3905,In_3592,In_1670);
and U3906 (N_3906,In_3545,In_1332);
nand U3907 (N_3907,In_1203,In_1123);
nor U3908 (N_3908,In_1674,In_4663);
and U3909 (N_3909,In_1181,In_184);
or U3910 (N_3910,In_1715,In_8);
or U3911 (N_3911,In_90,In_2856);
nor U3912 (N_3912,In_1916,In_1855);
or U3913 (N_3913,In_248,In_2107);
nand U3914 (N_3914,In_4315,In_4695);
and U3915 (N_3915,In_3862,In_519);
and U3916 (N_3916,In_4105,In_4583);
nand U3917 (N_3917,In_3514,In_3745);
nand U3918 (N_3918,In_4312,In_2822);
or U3919 (N_3919,In_120,In_630);
or U3920 (N_3920,In_1448,In_823);
nand U3921 (N_3921,In_1650,In_4361);
nor U3922 (N_3922,In_2476,In_3939);
and U3923 (N_3923,In_3914,In_275);
or U3924 (N_3924,In_1598,In_864);
and U3925 (N_3925,In_3593,In_2117);
xnor U3926 (N_3926,In_1470,In_4590);
xnor U3927 (N_3927,In_1163,In_1341);
nand U3928 (N_3928,In_2475,In_3838);
nand U3929 (N_3929,In_3180,In_527);
nor U3930 (N_3930,In_1121,In_3232);
or U3931 (N_3931,In_4947,In_2493);
or U3932 (N_3932,In_3468,In_575);
nor U3933 (N_3933,In_1663,In_1863);
and U3934 (N_3934,In_2457,In_4474);
nor U3935 (N_3935,In_1208,In_1001);
and U3936 (N_3936,In_3634,In_354);
or U3937 (N_3937,In_785,In_1422);
nand U3938 (N_3938,In_3966,In_2737);
and U3939 (N_3939,In_4707,In_2572);
nor U3940 (N_3940,In_4171,In_180);
xnor U3941 (N_3941,In_1520,In_1738);
nor U3942 (N_3942,In_159,In_2586);
xnor U3943 (N_3943,In_188,In_4240);
nand U3944 (N_3944,In_4478,In_461);
nand U3945 (N_3945,In_3313,In_420);
and U3946 (N_3946,In_1434,In_3605);
nand U3947 (N_3947,In_2806,In_679);
nor U3948 (N_3948,In_3550,In_3217);
nand U3949 (N_3949,In_4486,In_845);
nand U3950 (N_3950,In_592,In_3121);
or U3951 (N_3951,In_666,In_2468);
and U3952 (N_3952,In_1893,In_988);
and U3953 (N_3953,In_839,In_223);
xor U3954 (N_3954,In_4147,In_2889);
nand U3955 (N_3955,In_2062,In_3574);
and U3956 (N_3956,In_3606,In_3388);
nand U3957 (N_3957,In_2818,In_1830);
and U3958 (N_3958,In_907,In_316);
nand U3959 (N_3959,In_4774,In_4748);
and U3960 (N_3960,In_352,In_972);
nor U3961 (N_3961,In_2038,In_3943);
nor U3962 (N_3962,In_3287,In_3802);
or U3963 (N_3963,In_3522,In_2499);
xor U3964 (N_3964,In_610,In_4391);
nand U3965 (N_3965,In_1180,In_4416);
and U3966 (N_3966,In_324,In_2909);
or U3967 (N_3967,In_1022,In_1871);
nor U3968 (N_3968,In_3210,In_854);
nand U3969 (N_3969,In_3525,In_1444);
and U3970 (N_3970,In_2583,In_4566);
nor U3971 (N_3971,In_1502,In_228);
nand U3972 (N_3972,In_300,In_3324);
nand U3973 (N_3973,In_4665,In_2783);
nor U3974 (N_3974,In_2751,In_2008);
and U3975 (N_3975,In_4576,In_3573);
nor U3976 (N_3976,In_3319,In_4117);
nand U3977 (N_3977,In_3632,In_738);
nor U3978 (N_3978,In_3840,In_3109);
nor U3979 (N_3979,In_3653,In_1914);
or U3980 (N_3980,In_628,In_4315);
nand U3981 (N_3981,In_1815,In_3201);
nand U3982 (N_3982,In_573,In_4274);
nor U3983 (N_3983,In_4253,In_3504);
xor U3984 (N_3984,In_1408,In_2666);
or U3985 (N_3985,In_1686,In_4389);
nand U3986 (N_3986,In_1524,In_941);
or U3987 (N_3987,In_1824,In_1470);
or U3988 (N_3988,In_650,In_4199);
or U3989 (N_3989,In_4334,In_1241);
nor U3990 (N_3990,In_3613,In_1361);
xor U3991 (N_3991,In_4928,In_2393);
or U3992 (N_3992,In_1722,In_2298);
nand U3993 (N_3993,In_2749,In_539);
and U3994 (N_3994,In_966,In_2772);
or U3995 (N_3995,In_3232,In_2426);
nand U3996 (N_3996,In_3017,In_3522);
and U3997 (N_3997,In_4386,In_1082);
nand U3998 (N_3998,In_1653,In_1093);
nor U3999 (N_3999,In_3105,In_1358);
nor U4000 (N_4000,In_31,In_706);
nor U4001 (N_4001,In_2379,In_2685);
nand U4002 (N_4002,In_198,In_4699);
or U4003 (N_4003,In_2566,In_1665);
and U4004 (N_4004,In_2661,In_1025);
xnor U4005 (N_4005,In_4792,In_2288);
nor U4006 (N_4006,In_1785,In_2216);
or U4007 (N_4007,In_2236,In_3418);
or U4008 (N_4008,In_2592,In_2478);
and U4009 (N_4009,In_3305,In_1716);
and U4010 (N_4010,In_4078,In_1241);
and U4011 (N_4011,In_4458,In_442);
nand U4012 (N_4012,In_2786,In_1600);
or U4013 (N_4013,In_920,In_2972);
or U4014 (N_4014,In_827,In_4077);
nor U4015 (N_4015,In_2392,In_1519);
and U4016 (N_4016,In_2557,In_3540);
and U4017 (N_4017,In_567,In_2336);
xnor U4018 (N_4018,In_932,In_1341);
and U4019 (N_4019,In_4030,In_3938);
nor U4020 (N_4020,In_1694,In_239);
nor U4021 (N_4021,In_1200,In_2751);
nor U4022 (N_4022,In_2407,In_439);
and U4023 (N_4023,In_4306,In_1316);
nand U4024 (N_4024,In_4058,In_4999);
or U4025 (N_4025,In_4088,In_1356);
nor U4026 (N_4026,In_1506,In_504);
xnor U4027 (N_4027,In_639,In_2435);
xnor U4028 (N_4028,In_4892,In_1278);
xnor U4029 (N_4029,In_998,In_3282);
xnor U4030 (N_4030,In_1515,In_1944);
nand U4031 (N_4031,In_1172,In_1828);
or U4032 (N_4032,In_2485,In_1396);
nor U4033 (N_4033,In_1902,In_3845);
nand U4034 (N_4034,In_720,In_1205);
or U4035 (N_4035,In_4853,In_4794);
nand U4036 (N_4036,In_4310,In_790);
xor U4037 (N_4037,In_1385,In_4823);
nand U4038 (N_4038,In_3022,In_66);
nand U4039 (N_4039,In_1445,In_3642);
or U4040 (N_4040,In_2782,In_2160);
or U4041 (N_4041,In_3544,In_3892);
and U4042 (N_4042,In_3184,In_817);
xnor U4043 (N_4043,In_1164,In_1803);
nand U4044 (N_4044,In_3667,In_265);
nor U4045 (N_4045,In_3844,In_108);
and U4046 (N_4046,In_1499,In_893);
and U4047 (N_4047,In_3661,In_589);
xnor U4048 (N_4048,In_1976,In_2719);
nor U4049 (N_4049,In_240,In_3666);
or U4050 (N_4050,In_1565,In_2206);
nand U4051 (N_4051,In_4066,In_578);
nor U4052 (N_4052,In_3719,In_343);
and U4053 (N_4053,In_131,In_4347);
and U4054 (N_4054,In_1551,In_3941);
nand U4055 (N_4055,In_1892,In_2720);
and U4056 (N_4056,In_3669,In_4974);
nor U4057 (N_4057,In_2161,In_3116);
xnor U4058 (N_4058,In_4328,In_4270);
nor U4059 (N_4059,In_755,In_909);
nor U4060 (N_4060,In_3164,In_4839);
or U4061 (N_4061,In_645,In_483);
and U4062 (N_4062,In_49,In_4170);
xor U4063 (N_4063,In_2673,In_2199);
or U4064 (N_4064,In_4554,In_924);
xor U4065 (N_4065,In_1804,In_4191);
and U4066 (N_4066,In_1840,In_3884);
nand U4067 (N_4067,In_893,In_1972);
nand U4068 (N_4068,In_258,In_2104);
or U4069 (N_4069,In_3160,In_3766);
nor U4070 (N_4070,In_517,In_3859);
nor U4071 (N_4071,In_4923,In_2079);
nand U4072 (N_4072,In_1172,In_4314);
and U4073 (N_4073,In_2886,In_667);
nand U4074 (N_4074,In_2464,In_4353);
or U4075 (N_4075,In_4770,In_2480);
nor U4076 (N_4076,In_604,In_1798);
or U4077 (N_4077,In_1282,In_4566);
or U4078 (N_4078,In_1212,In_4420);
or U4079 (N_4079,In_446,In_95);
and U4080 (N_4080,In_690,In_2582);
nand U4081 (N_4081,In_1351,In_4227);
nor U4082 (N_4082,In_3669,In_2367);
or U4083 (N_4083,In_2282,In_3800);
and U4084 (N_4084,In_655,In_3571);
nor U4085 (N_4085,In_4607,In_4343);
or U4086 (N_4086,In_4240,In_4082);
nand U4087 (N_4087,In_3130,In_3618);
nor U4088 (N_4088,In_2746,In_1679);
nor U4089 (N_4089,In_3936,In_2889);
and U4090 (N_4090,In_1785,In_4549);
or U4091 (N_4091,In_4023,In_1761);
nor U4092 (N_4092,In_145,In_290);
or U4093 (N_4093,In_1402,In_1366);
nor U4094 (N_4094,In_3303,In_4899);
and U4095 (N_4095,In_4628,In_76);
and U4096 (N_4096,In_887,In_1187);
nor U4097 (N_4097,In_1303,In_2700);
or U4098 (N_4098,In_3858,In_4694);
nand U4099 (N_4099,In_3632,In_4693);
nand U4100 (N_4100,In_4654,In_2515);
xor U4101 (N_4101,In_4403,In_531);
and U4102 (N_4102,In_4802,In_1757);
nand U4103 (N_4103,In_77,In_2702);
nand U4104 (N_4104,In_700,In_284);
nor U4105 (N_4105,In_1965,In_4922);
or U4106 (N_4106,In_2720,In_1837);
nand U4107 (N_4107,In_2310,In_4756);
and U4108 (N_4108,In_4722,In_2718);
or U4109 (N_4109,In_2068,In_4604);
nor U4110 (N_4110,In_4068,In_3298);
nand U4111 (N_4111,In_62,In_841);
xnor U4112 (N_4112,In_1989,In_2669);
or U4113 (N_4113,In_70,In_4838);
and U4114 (N_4114,In_4329,In_3896);
nor U4115 (N_4115,In_4770,In_1069);
nand U4116 (N_4116,In_892,In_1418);
or U4117 (N_4117,In_1597,In_3466);
and U4118 (N_4118,In_2305,In_3836);
nand U4119 (N_4119,In_4902,In_2406);
or U4120 (N_4120,In_639,In_2632);
nand U4121 (N_4121,In_1244,In_1184);
nand U4122 (N_4122,In_2751,In_3474);
or U4123 (N_4123,In_4346,In_2552);
or U4124 (N_4124,In_4640,In_3318);
or U4125 (N_4125,In_1875,In_2770);
nand U4126 (N_4126,In_1603,In_4532);
xor U4127 (N_4127,In_3349,In_4083);
and U4128 (N_4128,In_4900,In_925);
nor U4129 (N_4129,In_2690,In_2328);
or U4130 (N_4130,In_3231,In_975);
and U4131 (N_4131,In_3816,In_2816);
nor U4132 (N_4132,In_4135,In_766);
nor U4133 (N_4133,In_2494,In_2496);
nor U4134 (N_4134,In_2520,In_844);
nor U4135 (N_4135,In_15,In_2853);
or U4136 (N_4136,In_1020,In_2251);
and U4137 (N_4137,In_3777,In_4818);
and U4138 (N_4138,In_381,In_4237);
nand U4139 (N_4139,In_1647,In_4271);
nand U4140 (N_4140,In_3525,In_2034);
nor U4141 (N_4141,In_729,In_118);
nor U4142 (N_4142,In_2824,In_3155);
nor U4143 (N_4143,In_4019,In_4929);
nor U4144 (N_4144,In_4527,In_1886);
or U4145 (N_4145,In_4211,In_2842);
or U4146 (N_4146,In_649,In_3005);
xor U4147 (N_4147,In_3807,In_3661);
or U4148 (N_4148,In_667,In_3349);
nor U4149 (N_4149,In_3126,In_4072);
or U4150 (N_4150,In_4646,In_3072);
nand U4151 (N_4151,In_1290,In_2079);
nand U4152 (N_4152,In_2990,In_2873);
nand U4153 (N_4153,In_1082,In_1387);
and U4154 (N_4154,In_4629,In_2833);
nand U4155 (N_4155,In_4172,In_2166);
or U4156 (N_4156,In_614,In_747);
nand U4157 (N_4157,In_1808,In_2801);
and U4158 (N_4158,In_377,In_633);
and U4159 (N_4159,In_1964,In_3758);
or U4160 (N_4160,In_4439,In_3807);
and U4161 (N_4161,In_4973,In_4113);
xor U4162 (N_4162,In_2255,In_3573);
and U4163 (N_4163,In_9,In_3333);
and U4164 (N_4164,In_1954,In_4389);
nand U4165 (N_4165,In_811,In_3098);
or U4166 (N_4166,In_792,In_4506);
nor U4167 (N_4167,In_4734,In_2395);
nor U4168 (N_4168,In_4298,In_4605);
nand U4169 (N_4169,In_4313,In_2210);
or U4170 (N_4170,In_3367,In_76);
nor U4171 (N_4171,In_4762,In_3917);
or U4172 (N_4172,In_1678,In_4377);
or U4173 (N_4173,In_2431,In_1399);
nor U4174 (N_4174,In_3898,In_2219);
or U4175 (N_4175,In_1424,In_326);
nor U4176 (N_4176,In_1689,In_3492);
nand U4177 (N_4177,In_4340,In_1391);
or U4178 (N_4178,In_4522,In_892);
nor U4179 (N_4179,In_2306,In_4583);
nor U4180 (N_4180,In_663,In_4196);
nor U4181 (N_4181,In_481,In_3558);
nand U4182 (N_4182,In_2837,In_290);
nand U4183 (N_4183,In_787,In_3169);
nand U4184 (N_4184,In_3957,In_906);
or U4185 (N_4185,In_3747,In_3091);
xnor U4186 (N_4186,In_1734,In_1221);
nor U4187 (N_4187,In_2318,In_504);
or U4188 (N_4188,In_532,In_3974);
nand U4189 (N_4189,In_2786,In_2319);
nand U4190 (N_4190,In_1394,In_2661);
and U4191 (N_4191,In_4206,In_673);
and U4192 (N_4192,In_4793,In_3240);
nor U4193 (N_4193,In_1352,In_1292);
and U4194 (N_4194,In_2358,In_4843);
or U4195 (N_4195,In_661,In_2541);
or U4196 (N_4196,In_4280,In_4090);
nor U4197 (N_4197,In_4632,In_2720);
nand U4198 (N_4198,In_2895,In_2224);
or U4199 (N_4199,In_2413,In_4456);
and U4200 (N_4200,In_3404,In_3674);
nor U4201 (N_4201,In_3004,In_4606);
or U4202 (N_4202,In_449,In_1144);
nor U4203 (N_4203,In_1071,In_3767);
or U4204 (N_4204,In_4272,In_2538);
and U4205 (N_4205,In_4386,In_2860);
nand U4206 (N_4206,In_641,In_246);
and U4207 (N_4207,In_3232,In_1825);
nand U4208 (N_4208,In_4636,In_2041);
or U4209 (N_4209,In_1563,In_3301);
xor U4210 (N_4210,In_1572,In_2186);
or U4211 (N_4211,In_4916,In_1452);
nor U4212 (N_4212,In_1343,In_3502);
and U4213 (N_4213,In_854,In_211);
nand U4214 (N_4214,In_87,In_2580);
and U4215 (N_4215,In_1510,In_808);
xnor U4216 (N_4216,In_2441,In_4024);
nor U4217 (N_4217,In_2655,In_679);
and U4218 (N_4218,In_3951,In_2756);
xor U4219 (N_4219,In_1820,In_1171);
nand U4220 (N_4220,In_2232,In_46);
nor U4221 (N_4221,In_1646,In_4569);
nand U4222 (N_4222,In_3356,In_1029);
and U4223 (N_4223,In_819,In_2632);
nor U4224 (N_4224,In_3942,In_4918);
nor U4225 (N_4225,In_4242,In_4018);
or U4226 (N_4226,In_1310,In_1426);
nor U4227 (N_4227,In_4152,In_4348);
nand U4228 (N_4228,In_437,In_3976);
or U4229 (N_4229,In_4395,In_124);
nand U4230 (N_4230,In_2897,In_4591);
nand U4231 (N_4231,In_2103,In_3442);
nand U4232 (N_4232,In_1041,In_1181);
and U4233 (N_4233,In_4695,In_2846);
or U4234 (N_4234,In_238,In_22);
or U4235 (N_4235,In_2638,In_4510);
and U4236 (N_4236,In_1693,In_1304);
nand U4237 (N_4237,In_1836,In_4461);
nor U4238 (N_4238,In_713,In_2483);
or U4239 (N_4239,In_4173,In_185);
and U4240 (N_4240,In_4469,In_2147);
nand U4241 (N_4241,In_377,In_1585);
xnor U4242 (N_4242,In_98,In_1326);
xor U4243 (N_4243,In_4562,In_2081);
and U4244 (N_4244,In_1198,In_3050);
nor U4245 (N_4245,In_1617,In_3722);
or U4246 (N_4246,In_4363,In_1071);
nand U4247 (N_4247,In_837,In_3063);
or U4248 (N_4248,In_3462,In_2299);
nand U4249 (N_4249,In_1182,In_2100);
nand U4250 (N_4250,In_4278,In_3323);
xnor U4251 (N_4251,In_4067,In_2000);
or U4252 (N_4252,In_2747,In_1214);
or U4253 (N_4253,In_4433,In_1888);
nor U4254 (N_4254,In_1535,In_3414);
or U4255 (N_4255,In_1551,In_235);
or U4256 (N_4256,In_3949,In_1868);
nand U4257 (N_4257,In_2137,In_4467);
or U4258 (N_4258,In_2918,In_3079);
nor U4259 (N_4259,In_82,In_2470);
nor U4260 (N_4260,In_4421,In_4845);
nor U4261 (N_4261,In_113,In_2632);
nand U4262 (N_4262,In_1043,In_800);
and U4263 (N_4263,In_2818,In_2557);
nor U4264 (N_4264,In_1817,In_144);
nor U4265 (N_4265,In_332,In_4354);
or U4266 (N_4266,In_2201,In_92);
nand U4267 (N_4267,In_2358,In_177);
and U4268 (N_4268,In_1878,In_1);
and U4269 (N_4269,In_884,In_2936);
nor U4270 (N_4270,In_1943,In_1986);
nor U4271 (N_4271,In_3627,In_230);
or U4272 (N_4272,In_1344,In_3135);
nor U4273 (N_4273,In_4804,In_4262);
and U4274 (N_4274,In_1087,In_1351);
xnor U4275 (N_4275,In_98,In_1051);
and U4276 (N_4276,In_3736,In_1503);
xor U4277 (N_4277,In_535,In_2203);
nand U4278 (N_4278,In_2136,In_886);
xor U4279 (N_4279,In_2171,In_499);
or U4280 (N_4280,In_3636,In_909);
or U4281 (N_4281,In_1513,In_2404);
or U4282 (N_4282,In_1232,In_112);
xnor U4283 (N_4283,In_4885,In_58);
nand U4284 (N_4284,In_896,In_4748);
and U4285 (N_4285,In_3972,In_853);
nand U4286 (N_4286,In_3868,In_4712);
xor U4287 (N_4287,In_2747,In_1781);
or U4288 (N_4288,In_84,In_1070);
xor U4289 (N_4289,In_2358,In_2735);
or U4290 (N_4290,In_2901,In_805);
nor U4291 (N_4291,In_1349,In_4370);
nand U4292 (N_4292,In_790,In_2514);
nor U4293 (N_4293,In_3462,In_4600);
xnor U4294 (N_4294,In_2046,In_3219);
or U4295 (N_4295,In_3386,In_2404);
nand U4296 (N_4296,In_3655,In_1043);
or U4297 (N_4297,In_4186,In_571);
nor U4298 (N_4298,In_1122,In_1665);
or U4299 (N_4299,In_3786,In_636);
xnor U4300 (N_4300,In_2196,In_1126);
and U4301 (N_4301,In_719,In_2541);
nor U4302 (N_4302,In_907,In_4856);
or U4303 (N_4303,In_3554,In_3033);
nand U4304 (N_4304,In_1488,In_458);
nor U4305 (N_4305,In_4701,In_977);
xnor U4306 (N_4306,In_3644,In_2827);
nor U4307 (N_4307,In_3299,In_4476);
nor U4308 (N_4308,In_4049,In_1340);
and U4309 (N_4309,In_1334,In_3188);
or U4310 (N_4310,In_4962,In_2857);
xor U4311 (N_4311,In_1252,In_4185);
xnor U4312 (N_4312,In_1369,In_4353);
and U4313 (N_4313,In_3209,In_2258);
or U4314 (N_4314,In_2610,In_759);
and U4315 (N_4315,In_1618,In_1648);
or U4316 (N_4316,In_3469,In_2748);
nand U4317 (N_4317,In_3648,In_4110);
and U4318 (N_4318,In_3842,In_1458);
and U4319 (N_4319,In_984,In_1519);
nor U4320 (N_4320,In_1312,In_1691);
nor U4321 (N_4321,In_2273,In_4490);
nand U4322 (N_4322,In_635,In_3600);
nand U4323 (N_4323,In_3005,In_817);
nand U4324 (N_4324,In_865,In_228);
nand U4325 (N_4325,In_4044,In_1713);
or U4326 (N_4326,In_322,In_4500);
nor U4327 (N_4327,In_1302,In_3349);
or U4328 (N_4328,In_1395,In_3085);
and U4329 (N_4329,In_4850,In_4073);
and U4330 (N_4330,In_1742,In_3340);
nand U4331 (N_4331,In_871,In_2716);
and U4332 (N_4332,In_2363,In_4215);
and U4333 (N_4333,In_4784,In_3761);
and U4334 (N_4334,In_3240,In_2640);
and U4335 (N_4335,In_4097,In_704);
nand U4336 (N_4336,In_2714,In_2012);
nor U4337 (N_4337,In_22,In_3875);
nor U4338 (N_4338,In_3167,In_741);
and U4339 (N_4339,In_2876,In_3915);
nor U4340 (N_4340,In_2258,In_3336);
and U4341 (N_4341,In_2957,In_3915);
nor U4342 (N_4342,In_1659,In_4395);
and U4343 (N_4343,In_2849,In_2987);
nand U4344 (N_4344,In_2790,In_998);
and U4345 (N_4345,In_975,In_99);
or U4346 (N_4346,In_2329,In_579);
or U4347 (N_4347,In_2508,In_2327);
xnor U4348 (N_4348,In_3458,In_2161);
nor U4349 (N_4349,In_2197,In_3851);
and U4350 (N_4350,In_4376,In_3914);
nand U4351 (N_4351,In_1690,In_1985);
or U4352 (N_4352,In_2368,In_794);
nand U4353 (N_4353,In_2758,In_2441);
and U4354 (N_4354,In_382,In_490);
nand U4355 (N_4355,In_2871,In_3898);
or U4356 (N_4356,In_3388,In_4913);
nand U4357 (N_4357,In_1091,In_3182);
nor U4358 (N_4358,In_2800,In_4142);
or U4359 (N_4359,In_2167,In_777);
nand U4360 (N_4360,In_1506,In_3215);
or U4361 (N_4361,In_1187,In_2721);
or U4362 (N_4362,In_2568,In_1568);
nand U4363 (N_4363,In_2656,In_2725);
nor U4364 (N_4364,In_1342,In_2604);
and U4365 (N_4365,In_936,In_3768);
or U4366 (N_4366,In_2430,In_705);
nand U4367 (N_4367,In_1655,In_2384);
nor U4368 (N_4368,In_2273,In_3603);
nand U4369 (N_4369,In_1548,In_1878);
nor U4370 (N_4370,In_3826,In_3922);
and U4371 (N_4371,In_1121,In_1652);
nand U4372 (N_4372,In_302,In_652);
nand U4373 (N_4373,In_3925,In_4765);
or U4374 (N_4374,In_2268,In_1834);
xor U4375 (N_4375,In_4403,In_811);
and U4376 (N_4376,In_4313,In_2340);
xor U4377 (N_4377,In_2019,In_2159);
or U4378 (N_4378,In_3486,In_3715);
nand U4379 (N_4379,In_1281,In_2468);
and U4380 (N_4380,In_2581,In_4904);
or U4381 (N_4381,In_4334,In_2341);
nor U4382 (N_4382,In_1211,In_2040);
and U4383 (N_4383,In_2143,In_916);
and U4384 (N_4384,In_4137,In_855);
nor U4385 (N_4385,In_437,In_1614);
and U4386 (N_4386,In_4354,In_4716);
or U4387 (N_4387,In_4769,In_4529);
nor U4388 (N_4388,In_3987,In_3247);
nand U4389 (N_4389,In_1295,In_695);
and U4390 (N_4390,In_3694,In_883);
nor U4391 (N_4391,In_1544,In_3654);
nand U4392 (N_4392,In_3092,In_1991);
and U4393 (N_4393,In_2936,In_4528);
and U4394 (N_4394,In_2706,In_848);
xor U4395 (N_4395,In_4380,In_4462);
or U4396 (N_4396,In_1739,In_3748);
nor U4397 (N_4397,In_4506,In_4673);
and U4398 (N_4398,In_4650,In_3573);
or U4399 (N_4399,In_557,In_3418);
nor U4400 (N_4400,In_4281,In_3220);
nor U4401 (N_4401,In_4209,In_2921);
xnor U4402 (N_4402,In_1660,In_2089);
and U4403 (N_4403,In_1531,In_4652);
and U4404 (N_4404,In_2514,In_1479);
and U4405 (N_4405,In_4295,In_3820);
and U4406 (N_4406,In_2376,In_2983);
nand U4407 (N_4407,In_3219,In_1960);
nand U4408 (N_4408,In_1729,In_4800);
or U4409 (N_4409,In_2381,In_4396);
and U4410 (N_4410,In_583,In_4281);
nand U4411 (N_4411,In_3687,In_4517);
and U4412 (N_4412,In_3993,In_646);
nand U4413 (N_4413,In_1407,In_528);
and U4414 (N_4414,In_4186,In_3082);
nand U4415 (N_4415,In_131,In_2602);
and U4416 (N_4416,In_3955,In_108);
nand U4417 (N_4417,In_2459,In_2852);
nor U4418 (N_4418,In_668,In_851);
nor U4419 (N_4419,In_3611,In_1386);
or U4420 (N_4420,In_3080,In_4572);
and U4421 (N_4421,In_2305,In_3169);
and U4422 (N_4422,In_200,In_1186);
xor U4423 (N_4423,In_788,In_4878);
nor U4424 (N_4424,In_271,In_2262);
or U4425 (N_4425,In_1726,In_341);
nand U4426 (N_4426,In_896,In_720);
or U4427 (N_4427,In_1634,In_3032);
or U4428 (N_4428,In_689,In_1179);
nand U4429 (N_4429,In_1826,In_4084);
or U4430 (N_4430,In_4005,In_2893);
xor U4431 (N_4431,In_461,In_4673);
nor U4432 (N_4432,In_2854,In_4479);
nand U4433 (N_4433,In_425,In_4786);
or U4434 (N_4434,In_671,In_4535);
nand U4435 (N_4435,In_3772,In_2734);
and U4436 (N_4436,In_3756,In_948);
nand U4437 (N_4437,In_2010,In_390);
and U4438 (N_4438,In_2184,In_1954);
nand U4439 (N_4439,In_3214,In_916);
or U4440 (N_4440,In_4684,In_2945);
nand U4441 (N_4441,In_347,In_611);
nor U4442 (N_4442,In_266,In_2794);
nor U4443 (N_4443,In_1423,In_3840);
nand U4444 (N_4444,In_1498,In_4203);
nor U4445 (N_4445,In_2360,In_4227);
or U4446 (N_4446,In_3432,In_4515);
nand U4447 (N_4447,In_3996,In_3803);
or U4448 (N_4448,In_1688,In_3363);
nand U4449 (N_4449,In_4436,In_1985);
xnor U4450 (N_4450,In_1071,In_4968);
or U4451 (N_4451,In_2571,In_1282);
nor U4452 (N_4452,In_3727,In_1098);
nor U4453 (N_4453,In_4485,In_3158);
and U4454 (N_4454,In_904,In_2362);
or U4455 (N_4455,In_4649,In_4724);
and U4456 (N_4456,In_934,In_4505);
xor U4457 (N_4457,In_2618,In_2611);
nand U4458 (N_4458,In_1406,In_2637);
nand U4459 (N_4459,In_1587,In_1373);
nor U4460 (N_4460,In_4227,In_3685);
or U4461 (N_4461,In_1907,In_4749);
nand U4462 (N_4462,In_3404,In_422);
nand U4463 (N_4463,In_2814,In_639);
and U4464 (N_4464,In_4290,In_725);
nor U4465 (N_4465,In_2883,In_2284);
nor U4466 (N_4466,In_3069,In_4478);
nand U4467 (N_4467,In_4895,In_2085);
or U4468 (N_4468,In_2424,In_2525);
or U4469 (N_4469,In_1543,In_1103);
nand U4470 (N_4470,In_1894,In_2779);
or U4471 (N_4471,In_4415,In_3405);
nand U4472 (N_4472,In_608,In_547);
or U4473 (N_4473,In_4887,In_2767);
and U4474 (N_4474,In_4715,In_4644);
and U4475 (N_4475,In_2577,In_1097);
nand U4476 (N_4476,In_2345,In_1990);
nand U4477 (N_4477,In_2666,In_1384);
or U4478 (N_4478,In_4729,In_3284);
or U4479 (N_4479,In_143,In_2175);
nand U4480 (N_4480,In_1311,In_2084);
xnor U4481 (N_4481,In_1177,In_1610);
or U4482 (N_4482,In_2667,In_4178);
nand U4483 (N_4483,In_4294,In_3850);
nand U4484 (N_4484,In_2973,In_3394);
nand U4485 (N_4485,In_33,In_1503);
and U4486 (N_4486,In_961,In_2465);
nor U4487 (N_4487,In_266,In_2578);
nand U4488 (N_4488,In_3687,In_2990);
and U4489 (N_4489,In_2141,In_1702);
and U4490 (N_4490,In_1014,In_2326);
and U4491 (N_4491,In_1201,In_3681);
and U4492 (N_4492,In_3121,In_1029);
and U4493 (N_4493,In_2637,In_167);
xnor U4494 (N_4494,In_955,In_143);
or U4495 (N_4495,In_879,In_3997);
or U4496 (N_4496,In_1132,In_3165);
nor U4497 (N_4497,In_1480,In_4869);
or U4498 (N_4498,In_2525,In_3);
or U4499 (N_4499,In_2197,In_2500);
and U4500 (N_4500,In_3034,In_3536);
nand U4501 (N_4501,In_2596,In_4356);
and U4502 (N_4502,In_4562,In_3041);
and U4503 (N_4503,In_3300,In_952);
nor U4504 (N_4504,In_4871,In_3617);
or U4505 (N_4505,In_4521,In_4378);
and U4506 (N_4506,In_3760,In_1849);
nand U4507 (N_4507,In_2661,In_691);
nand U4508 (N_4508,In_859,In_1331);
and U4509 (N_4509,In_268,In_956);
nand U4510 (N_4510,In_4652,In_4507);
and U4511 (N_4511,In_967,In_1391);
or U4512 (N_4512,In_3930,In_1640);
and U4513 (N_4513,In_4470,In_1370);
or U4514 (N_4514,In_2647,In_1325);
nand U4515 (N_4515,In_4903,In_1654);
or U4516 (N_4516,In_1077,In_2820);
and U4517 (N_4517,In_2627,In_2111);
and U4518 (N_4518,In_2955,In_141);
nand U4519 (N_4519,In_53,In_744);
and U4520 (N_4520,In_820,In_4828);
xnor U4521 (N_4521,In_1111,In_3254);
nand U4522 (N_4522,In_1952,In_1088);
or U4523 (N_4523,In_1698,In_4887);
or U4524 (N_4524,In_67,In_4133);
or U4525 (N_4525,In_781,In_1069);
or U4526 (N_4526,In_1963,In_2768);
nor U4527 (N_4527,In_4373,In_3835);
nor U4528 (N_4528,In_431,In_4622);
nand U4529 (N_4529,In_3242,In_2203);
or U4530 (N_4530,In_2087,In_639);
nor U4531 (N_4531,In_4849,In_4896);
nand U4532 (N_4532,In_3359,In_2819);
nor U4533 (N_4533,In_4986,In_658);
xor U4534 (N_4534,In_1623,In_1603);
nor U4535 (N_4535,In_2334,In_881);
nand U4536 (N_4536,In_3244,In_3791);
nand U4537 (N_4537,In_2139,In_4919);
nor U4538 (N_4538,In_791,In_923);
or U4539 (N_4539,In_4737,In_3541);
nand U4540 (N_4540,In_398,In_2275);
nand U4541 (N_4541,In_3578,In_2125);
xor U4542 (N_4542,In_2991,In_4065);
or U4543 (N_4543,In_2343,In_606);
and U4544 (N_4544,In_3335,In_2201);
or U4545 (N_4545,In_3621,In_3472);
or U4546 (N_4546,In_4114,In_4697);
nor U4547 (N_4547,In_221,In_4778);
and U4548 (N_4548,In_1782,In_582);
nor U4549 (N_4549,In_1060,In_2242);
and U4550 (N_4550,In_1501,In_2782);
or U4551 (N_4551,In_1185,In_2314);
or U4552 (N_4552,In_2460,In_4048);
nor U4553 (N_4553,In_1842,In_2839);
nand U4554 (N_4554,In_3855,In_2027);
and U4555 (N_4555,In_4902,In_4332);
nor U4556 (N_4556,In_3952,In_3466);
or U4557 (N_4557,In_4798,In_1375);
nor U4558 (N_4558,In_3717,In_3120);
or U4559 (N_4559,In_896,In_2378);
xnor U4560 (N_4560,In_78,In_2062);
nand U4561 (N_4561,In_1371,In_4193);
or U4562 (N_4562,In_1349,In_1270);
or U4563 (N_4563,In_2986,In_3479);
nor U4564 (N_4564,In_2299,In_3358);
or U4565 (N_4565,In_3775,In_3186);
nand U4566 (N_4566,In_130,In_73);
nor U4567 (N_4567,In_4726,In_458);
nor U4568 (N_4568,In_339,In_2673);
and U4569 (N_4569,In_903,In_4494);
or U4570 (N_4570,In_3725,In_3702);
and U4571 (N_4571,In_4481,In_53);
nand U4572 (N_4572,In_3278,In_2784);
nor U4573 (N_4573,In_2572,In_471);
and U4574 (N_4574,In_4477,In_3978);
or U4575 (N_4575,In_1585,In_709);
and U4576 (N_4576,In_3986,In_2589);
nand U4577 (N_4577,In_2822,In_4099);
or U4578 (N_4578,In_4960,In_2503);
or U4579 (N_4579,In_2294,In_4736);
nor U4580 (N_4580,In_1771,In_4438);
nor U4581 (N_4581,In_1867,In_2787);
or U4582 (N_4582,In_4871,In_4433);
and U4583 (N_4583,In_614,In_1823);
or U4584 (N_4584,In_2341,In_2732);
nor U4585 (N_4585,In_209,In_1176);
nand U4586 (N_4586,In_4978,In_4400);
or U4587 (N_4587,In_4251,In_948);
nand U4588 (N_4588,In_2865,In_4870);
and U4589 (N_4589,In_881,In_804);
nor U4590 (N_4590,In_4178,In_2337);
nor U4591 (N_4591,In_3681,In_4571);
nand U4592 (N_4592,In_829,In_1740);
or U4593 (N_4593,In_4664,In_3606);
nor U4594 (N_4594,In_1887,In_1043);
xor U4595 (N_4595,In_2599,In_725);
or U4596 (N_4596,In_4600,In_4459);
and U4597 (N_4597,In_1858,In_2122);
or U4598 (N_4598,In_2728,In_1121);
xor U4599 (N_4599,In_4324,In_403);
or U4600 (N_4600,In_3787,In_2237);
nand U4601 (N_4601,In_2639,In_3176);
and U4602 (N_4602,In_4377,In_4983);
or U4603 (N_4603,In_4161,In_666);
nand U4604 (N_4604,In_167,In_403);
nand U4605 (N_4605,In_649,In_1165);
nand U4606 (N_4606,In_1882,In_4651);
nor U4607 (N_4607,In_2893,In_4356);
nor U4608 (N_4608,In_3435,In_2060);
xor U4609 (N_4609,In_4973,In_758);
or U4610 (N_4610,In_3852,In_880);
or U4611 (N_4611,In_921,In_4036);
or U4612 (N_4612,In_4936,In_1848);
nand U4613 (N_4613,In_3964,In_4735);
nor U4614 (N_4614,In_2041,In_3240);
nor U4615 (N_4615,In_4598,In_131);
and U4616 (N_4616,In_3711,In_4618);
nand U4617 (N_4617,In_974,In_2650);
nand U4618 (N_4618,In_1151,In_2647);
and U4619 (N_4619,In_3868,In_1574);
or U4620 (N_4620,In_3970,In_1051);
nor U4621 (N_4621,In_2831,In_3788);
nand U4622 (N_4622,In_4511,In_1919);
nand U4623 (N_4623,In_120,In_4777);
nand U4624 (N_4624,In_2635,In_4552);
and U4625 (N_4625,In_2172,In_905);
xnor U4626 (N_4626,In_403,In_4127);
and U4627 (N_4627,In_4058,In_353);
nand U4628 (N_4628,In_4018,In_2358);
xor U4629 (N_4629,In_4035,In_1208);
or U4630 (N_4630,In_22,In_3815);
nand U4631 (N_4631,In_4584,In_4289);
nand U4632 (N_4632,In_297,In_1676);
nor U4633 (N_4633,In_541,In_24);
and U4634 (N_4634,In_4573,In_189);
nor U4635 (N_4635,In_4083,In_1971);
or U4636 (N_4636,In_1969,In_1829);
or U4637 (N_4637,In_954,In_4183);
xor U4638 (N_4638,In_915,In_3063);
or U4639 (N_4639,In_1315,In_1956);
and U4640 (N_4640,In_2987,In_3388);
nor U4641 (N_4641,In_165,In_1794);
nor U4642 (N_4642,In_3428,In_2564);
or U4643 (N_4643,In_3111,In_3276);
or U4644 (N_4644,In_1944,In_1204);
and U4645 (N_4645,In_593,In_245);
nor U4646 (N_4646,In_769,In_1658);
and U4647 (N_4647,In_4945,In_3647);
or U4648 (N_4648,In_1130,In_3783);
nand U4649 (N_4649,In_618,In_1770);
nor U4650 (N_4650,In_3985,In_4407);
and U4651 (N_4651,In_2539,In_2265);
and U4652 (N_4652,In_2391,In_2392);
xnor U4653 (N_4653,In_986,In_4031);
or U4654 (N_4654,In_2984,In_3332);
and U4655 (N_4655,In_2708,In_2241);
xnor U4656 (N_4656,In_2480,In_1136);
or U4657 (N_4657,In_1009,In_578);
and U4658 (N_4658,In_1950,In_78);
or U4659 (N_4659,In_987,In_3948);
or U4660 (N_4660,In_1517,In_3999);
nand U4661 (N_4661,In_4618,In_1284);
nand U4662 (N_4662,In_1218,In_4405);
xor U4663 (N_4663,In_552,In_3272);
nor U4664 (N_4664,In_2408,In_3528);
nand U4665 (N_4665,In_2803,In_895);
nor U4666 (N_4666,In_4335,In_2666);
nand U4667 (N_4667,In_3338,In_3974);
xnor U4668 (N_4668,In_1756,In_2731);
xor U4669 (N_4669,In_4489,In_1857);
or U4670 (N_4670,In_1440,In_3804);
and U4671 (N_4671,In_2886,In_2127);
or U4672 (N_4672,In_1760,In_3215);
nor U4673 (N_4673,In_4808,In_64);
or U4674 (N_4674,In_4922,In_2043);
or U4675 (N_4675,In_4024,In_2024);
or U4676 (N_4676,In_197,In_1733);
xnor U4677 (N_4677,In_882,In_3771);
nor U4678 (N_4678,In_3901,In_4272);
nor U4679 (N_4679,In_3893,In_1794);
and U4680 (N_4680,In_1132,In_4746);
or U4681 (N_4681,In_444,In_2017);
nor U4682 (N_4682,In_4595,In_2298);
nor U4683 (N_4683,In_4781,In_4318);
nand U4684 (N_4684,In_2671,In_4635);
nand U4685 (N_4685,In_4705,In_2780);
xnor U4686 (N_4686,In_3432,In_3833);
nor U4687 (N_4687,In_1273,In_280);
nand U4688 (N_4688,In_2214,In_4410);
and U4689 (N_4689,In_4759,In_2494);
or U4690 (N_4690,In_3483,In_4545);
nand U4691 (N_4691,In_645,In_3527);
and U4692 (N_4692,In_3247,In_3740);
or U4693 (N_4693,In_3771,In_3292);
and U4694 (N_4694,In_4434,In_3638);
nand U4695 (N_4695,In_2512,In_3932);
xnor U4696 (N_4696,In_4571,In_1872);
and U4697 (N_4697,In_2370,In_4470);
or U4698 (N_4698,In_311,In_169);
and U4699 (N_4699,In_392,In_2380);
xnor U4700 (N_4700,In_913,In_556);
or U4701 (N_4701,In_2603,In_1360);
nor U4702 (N_4702,In_902,In_3957);
or U4703 (N_4703,In_3909,In_2353);
nor U4704 (N_4704,In_2530,In_848);
nor U4705 (N_4705,In_1638,In_2963);
or U4706 (N_4706,In_2733,In_3216);
xor U4707 (N_4707,In_2299,In_3838);
and U4708 (N_4708,In_1171,In_4945);
nor U4709 (N_4709,In_4271,In_1155);
nand U4710 (N_4710,In_362,In_2176);
or U4711 (N_4711,In_3227,In_233);
xor U4712 (N_4712,In_1155,In_3456);
nand U4713 (N_4713,In_3911,In_567);
nor U4714 (N_4714,In_2885,In_2824);
or U4715 (N_4715,In_57,In_3355);
and U4716 (N_4716,In_1312,In_704);
xnor U4717 (N_4717,In_4378,In_968);
and U4718 (N_4718,In_2117,In_534);
or U4719 (N_4719,In_2551,In_4097);
nor U4720 (N_4720,In_4433,In_517);
and U4721 (N_4721,In_3951,In_639);
or U4722 (N_4722,In_4238,In_4844);
nor U4723 (N_4723,In_2300,In_4054);
nor U4724 (N_4724,In_2964,In_3400);
nand U4725 (N_4725,In_2591,In_735);
nand U4726 (N_4726,In_3030,In_4591);
or U4727 (N_4727,In_1643,In_2487);
nor U4728 (N_4728,In_553,In_4520);
and U4729 (N_4729,In_4554,In_1988);
nand U4730 (N_4730,In_1919,In_3870);
nor U4731 (N_4731,In_4932,In_3810);
and U4732 (N_4732,In_1763,In_1318);
or U4733 (N_4733,In_4057,In_1907);
or U4734 (N_4734,In_4623,In_1223);
and U4735 (N_4735,In_1191,In_89);
nor U4736 (N_4736,In_4067,In_1788);
or U4737 (N_4737,In_4719,In_2406);
and U4738 (N_4738,In_505,In_899);
and U4739 (N_4739,In_3805,In_2244);
xor U4740 (N_4740,In_1834,In_4344);
or U4741 (N_4741,In_73,In_4202);
xnor U4742 (N_4742,In_4565,In_4449);
nor U4743 (N_4743,In_2961,In_891);
or U4744 (N_4744,In_4889,In_394);
nor U4745 (N_4745,In_3460,In_810);
and U4746 (N_4746,In_2713,In_3833);
nand U4747 (N_4747,In_905,In_3373);
and U4748 (N_4748,In_4092,In_1355);
nand U4749 (N_4749,In_511,In_189);
and U4750 (N_4750,In_4485,In_3760);
or U4751 (N_4751,In_2467,In_4236);
nor U4752 (N_4752,In_931,In_3723);
nand U4753 (N_4753,In_2564,In_652);
or U4754 (N_4754,In_1228,In_4919);
and U4755 (N_4755,In_3917,In_3378);
nand U4756 (N_4756,In_2265,In_4385);
nand U4757 (N_4757,In_3298,In_1883);
and U4758 (N_4758,In_1981,In_3108);
nor U4759 (N_4759,In_4147,In_414);
and U4760 (N_4760,In_213,In_1868);
and U4761 (N_4761,In_4501,In_1581);
nand U4762 (N_4762,In_741,In_1781);
nand U4763 (N_4763,In_2433,In_2010);
and U4764 (N_4764,In_3160,In_1957);
or U4765 (N_4765,In_2583,In_2608);
nor U4766 (N_4766,In_3691,In_1905);
xnor U4767 (N_4767,In_883,In_4412);
or U4768 (N_4768,In_1426,In_3890);
and U4769 (N_4769,In_35,In_3370);
nand U4770 (N_4770,In_4964,In_4493);
and U4771 (N_4771,In_3198,In_3533);
xor U4772 (N_4772,In_540,In_889);
nand U4773 (N_4773,In_1431,In_2350);
nor U4774 (N_4774,In_464,In_1680);
or U4775 (N_4775,In_1952,In_1991);
nand U4776 (N_4776,In_1445,In_3736);
and U4777 (N_4777,In_1093,In_4947);
nand U4778 (N_4778,In_1984,In_4688);
nand U4779 (N_4779,In_2450,In_4468);
or U4780 (N_4780,In_2394,In_3369);
nand U4781 (N_4781,In_4682,In_2092);
or U4782 (N_4782,In_3292,In_178);
or U4783 (N_4783,In_1095,In_3907);
nand U4784 (N_4784,In_4400,In_3136);
and U4785 (N_4785,In_4597,In_2535);
xor U4786 (N_4786,In_2284,In_3408);
nand U4787 (N_4787,In_2820,In_1381);
nor U4788 (N_4788,In_1121,In_2454);
or U4789 (N_4789,In_4212,In_3757);
or U4790 (N_4790,In_4580,In_4655);
and U4791 (N_4791,In_2935,In_4487);
or U4792 (N_4792,In_1930,In_926);
and U4793 (N_4793,In_4988,In_2468);
nand U4794 (N_4794,In_558,In_3242);
nor U4795 (N_4795,In_3880,In_1399);
nand U4796 (N_4796,In_30,In_1247);
nand U4797 (N_4797,In_4508,In_1957);
nand U4798 (N_4798,In_2983,In_1974);
nor U4799 (N_4799,In_383,In_1671);
xor U4800 (N_4800,In_3459,In_2876);
nor U4801 (N_4801,In_3014,In_131);
xor U4802 (N_4802,In_1884,In_4515);
and U4803 (N_4803,In_606,In_1002);
and U4804 (N_4804,In_13,In_1649);
or U4805 (N_4805,In_1124,In_2406);
nor U4806 (N_4806,In_65,In_4545);
and U4807 (N_4807,In_3382,In_2945);
nor U4808 (N_4808,In_1479,In_3711);
nand U4809 (N_4809,In_3271,In_1507);
and U4810 (N_4810,In_4736,In_607);
nor U4811 (N_4811,In_1572,In_1809);
and U4812 (N_4812,In_4568,In_1335);
or U4813 (N_4813,In_1247,In_2850);
or U4814 (N_4814,In_2090,In_574);
xor U4815 (N_4815,In_2439,In_3893);
and U4816 (N_4816,In_4547,In_4471);
nand U4817 (N_4817,In_88,In_588);
nand U4818 (N_4818,In_1489,In_1391);
nor U4819 (N_4819,In_4949,In_2959);
nand U4820 (N_4820,In_4144,In_4082);
and U4821 (N_4821,In_4413,In_3764);
nor U4822 (N_4822,In_4411,In_483);
nor U4823 (N_4823,In_43,In_3662);
or U4824 (N_4824,In_1589,In_32);
or U4825 (N_4825,In_4233,In_1563);
and U4826 (N_4826,In_2431,In_2174);
or U4827 (N_4827,In_4538,In_3258);
nand U4828 (N_4828,In_3062,In_4582);
nor U4829 (N_4829,In_2230,In_787);
and U4830 (N_4830,In_2573,In_469);
nor U4831 (N_4831,In_772,In_2629);
or U4832 (N_4832,In_1558,In_3974);
nand U4833 (N_4833,In_3428,In_238);
or U4834 (N_4834,In_3066,In_1068);
nand U4835 (N_4835,In_3457,In_963);
and U4836 (N_4836,In_4606,In_1509);
nor U4837 (N_4837,In_558,In_2920);
or U4838 (N_4838,In_231,In_3111);
and U4839 (N_4839,In_4142,In_1422);
nand U4840 (N_4840,In_185,In_3558);
nor U4841 (N_4841,In_133,In_574);
and U4842 (N_4842,In_3616,In_4949);
nor U4843 (N_4843,In_2248,In_1891);
nand U4844 (N_4844,In_1804,In_2064);
nor U4845 (N_4845,In_1790,In_3816);
nor U4846 (N_4846,In_1976,In_4178);
or U4847 (N_4847,In_280,In_4593);
nor U4848 (N_4848,In_1412,In_721);
or U4849 (N_4849,In_980,In_3355);
nor U4850 (N_4850,In_4362,In_15);
nand U4851 (N_4851,In_670,In_4358);
nor U4852 (N_4852,In_233,In_2471);
nor U4853 (N_4853,In_297,In_2925);
xnor U4854 (N_4854,In_1419,In_2678);
xnor U4855 (N_4855,In_551,In_4907);
nand U4856 (N_4856,In_2833,In_2072);
nor U4857 (N_4857,In_4782,In_3799);
nand U4858 (N_4858,In_2724,In_2710);
and U4859 (N_4859,In_4072,In_4446);
and U4860 (N_4860,In_2335,In_2414);
xor U4861 (N_4861,In_2772,In_4248);
and U4862 (N_4862,In_2003,In_1256);
or U4863 (N_4863,In_364,In_1833);
nand U4864 (N_4864,In_3848,In_3965);
xor U4865 (N_4865,In_1946,In_2180);
nor U4866 (N_4866,In_2178,In_1635);
nor U4867 (N_4867,In_2235,In_4848);
nor U4868 (N_4868,In_2098,In_2801);
xnor U4869 (N_4869,In_3979,In_3874);
and U4870 (N_4870,In_4685,In_2485);
nand U4871 (N_4871,In_4558,In_3270);
nand U4872 (N_4872,In_833,In_3067);
or U4873 (N_4873,In_4873,In_2575);
nand U4874 (N_4874,In_1985,In_120);
and U4875 (N_4875,In_919,In_2490);
nor U4876 (N_4876,In_4432,In_3647);
nor U4877 (N_4877,In_4829,In_1630);
nor U4878 (N_4878,In_4934,In_1937);
xor U4879 (N_4879,In_4650,In_299);
or U4880 (N_4880,In_4941,In_726);
nand U4881 (N_4881,In_4784,In_3080);
nor U4882 (N_4882,In_1854,In_4331);
or U4883 (N_4883,In_2958,In_2119);
or U4884 (N_4884,In_1942,In_1940);
nand U4885 (N_4885,In_2881,In_775);
nand U4886 (N_4886,In_2811,In_1644);
nand U4887 (N_4887,In_2844,In_4266);
and U4888 (N_4888,In_3312,In_4589);
and U4889 (N_4889,In_1395,In_302);
nand U4890 (N_4890,In_1745,In_3138);
xor U4891 (N_4891,In_167,In_2097);
nor U4892 (N_4892,In_4916,In_4193);
and U4893 (N_4893,In_3580,In_2174);
or U4894 (N_4894,In_4262,In_2838);
nor U4895 (N_4895,In_2217,In_3738);
or U4896 (N_4896,In_3341,In_4531);
and U4897 (N_4897,In_2425,In_4529);
and U4898 (N_4898,In_3409,In_616);
nor U4899 (N_4899,In_1171,In_3937);
and U4900 (N_4900,In_1892,In_827);
nor U4901 (N_4901,In_2975,In_3823);
nand U4902 (N_4902,In_592,In_1312);
or U4903 (N_4903,In_1690,In_4475);
xnor U4904 (N_4904,In_2053,In_4229);
or U4905 (N_4905,In_4866,In_3630);
nor U4906 (N_4906,In_3979,In_3176);
nand U4907 (N_4907,In_3283,In_3656);
or U4908 (N_4908,In_3560,In_4735);
or U4909 (N_4909,In_1583,In_12);
nand U4910 (N_4910,In_3289,In_4787);
nand U4911 (N_4911,In_4949,In_1289);
or U4912 (N_4912,In_1768,In_1680);
or U4913 (N_4913,In_4224,In_4046);
nor U4914 (N_4914,In_278,In_1246);
or U4915 (N_4915,In_4126,In_1774);
or U4916 (N_4916,In_412,In_447);
or U4917 (N_4917,In_1241,In_2948);
nand U4918 (N_4918,In_2447,In_87);
nand U4919 (N_4919,In_522,In_1135);
and U4920 (N_4920,In_4900,In_940);
or U4921 (N_4921,In_386,In_4008);
nor U4922 (N_4922,In_2198,In_4905);
and U4923 (N_4923,In_4596,In_2440);
or U4924 (N_4924,In_1752,In_2779);
or U4925 (N_4925,In_1003,In_1067);
and U4926 (N_4926,In_3657,In_403);
or U4927 (N_4927,In_4083,In_1537);
or U4928 (N_4928,In_81,In_4388);
and U4929 (N_4929,In_3741,In_2960);
xor U4930 (N_4930,In_3446,In_1801);
nor U4931 (N_4931,In_937,In_4578);
and U4932 (N_4932,In_3545,In_3697);
nand U4933 (N_4933,In_3218,In_2138);
and U4934 (N_4934,In_2031,In_4580);
nor U4935 (N_4935,In_4538,In_3199);
xor U4936 (N_4936,In_1392,In_1404);
or U4937 (N_4937,In_2389,In_716);
or U4938 (N_4938,In_320,In_2446);
or U4939 (N_4939,In_1605,In_46);
nor U4940 (N_4940,In_1185,In_1275);
and U4941 (N_4941,In_1917,In_2227);
and U4942 (N_4942,In_1042,In_494);
xnor U4943 (N_4943,In_1030,In_3568);
and U4944 (N_4944,In_1312,In_3962);
and U4945 (N_4945,In_2457,In_747);
or U4946 (N_4946,In_2058,In_4910);
or U4947 (N_4947,In_4223,In_1004);
or U4948 (N_4948,In_793,In_4838);
and U4949 (N_4949,In_1129,In_4188);
nand U4950 (N_4950,In_4427,In_873);
nor U4951 (N_4951,In_2418,In_3688);
or U4952 (N_4952,In_4925,In_4631);
nor U4953 (N_4953,In_4490,In_3910);
nor U4954 (N_4954,In_2451,In_4050);
nand U4955 (N_4955,In_4751,In_2761);
nand U4956 (N_4956,In_3218,In_2052);
nor U4957 (N_4957,In_2432,In_2745);
nor U4958 (N_4958,In_322,In_4753);
and U4959 (N_4959,In_2582,In_4409);
and U4960 (N_4960,In_2407,In_3949);
and U4961 (N_4961,In_891,In_666);
and U4962 (N_4962,In_615,In_604);
nor U4963 (N_4963,In_3412,In_4823);
or U4964 (N_4964,In_3067,In_4099);
or U4965 (N_4965,In_1170,In_1818);
nand U4966 (N_4966,In_589,In_1047);
xnor U4967 (N_4967,In_4757,In_1611);
xnor U4968 (N_4968,In_1558,In_611);
nor U4969 (N_4969,In_556,In_4068);
xor U4970 (N_4970,In_4061,In_1075);
xnor U4971 (N_4971,In_241,In_41);
or U4972 (N_4972,In_1622,In_724);
and U4973 (N_4973,In_289,In_1671);
and U4974 (N_4974,In_4383,In_3299);
or U4975 (N_4975,In_113,In_1660);
or U4976 (N_4976,In_80,In_4797);
and U4977 (N_4977,In_3391,In_2215);
or U4978 (N_4978,In_3672,In_3409);
nand U4979 (N_4979,In_2075,In_600);
or U4980 (N_4980,In_1023,In_1508);
nand U4981 (N_4981,In_4421,In_4367);
and U4982 (N_4982,In_2459,In_1636);
nand U4983 (N_4983,In_3103,In_3740);
xor U4984 (N_4984,In_3780,In_3806);
nor U4985 (N_4985,In_2833,In_2408);
nor U4986 (N_4986,In_1092,In_3813);
nor U4987 (N_4987,In_4594,In_2925);
nor U4988 (N_4988,In_4259,In_4590);
xor U4989 (N_4989,In_4735,In_2328);
or U4990 (N_4990,In_2977,In_2079);
nand U4991 (N_4991,In_4724,In_34);
or U4992 (N_4992,In_3323,In_490);
or U4993 (N_4993,In_1848,In_3715);
nand U4994 (N_4994,In_1462,In_3078);
nor U4995 (N_4995,In_359,In_4147);
nor U4996 (N_4996,In_4242,In_822);
or U4997 (N_4997,In_1602,In_1087);
or U4998 (N_4998,In_1434,In_625);
or U4999 (N_4999,In_162,In_4805);
and U5000 (N_5000,In_1076,In_2474);
nand U5001 (N_5001,In_2798,In_244);
and U5002 (N_5002,In_840,In_3961);
nand U5003 (N_5003,In_2965,In_1354);
or U5004 (N_5004,In_870,In_3848);
and U5005 (N_5005,In_4906,In_2304);
nor U5006 (N_5006,In_905,In_3962);
and U5007 (N_5007,In_2639,In_4945);
xor U5008 (N_5008,In_2408,In_1974);
xor U5009 (N_5009,In_4293,In_1563);
nor U5010 (N_5010,In_4048,In_4762);
or U5011 (N_5011,In_2737,In_974);
or U5012 (N_5012,In_1295,In_3267);
nand U5013 (N_5013,In_504,In_4393);
or U5014 (N_5014,In_635,In_1279);
and U5015 (N_5015,In_1231,In_4225);
nor U5016 (N_5016,In_1138,In_1387);
nor U5017 (N_5017,In_3388,In_2570);
and U5018 (N_5018,In_3220,In_1042);
nand U5019 (N_5019,In_1862,In_4125);
xor U5020 (N_5020,In_3889,In_2961);
nor U5021 (N_5021,In_4071,In_3712);
and U5022 (N_5022,In_201,In_2932);
nand U5023 (N_5023,In_2515,In_1749);
and U5024 (N_5024,In_1437,In_3432);
nor U5025 (N_5025,In_3670,In_3724);
nand U5026 (N_5026,In_371,In_253);
xnor U5027 (N_5027,In_3194,In_2198);
nor U5028 (N_5028,In_7,In_944);
xor U5029 (N_5029,In_2671,In_3046);
xor U5030 (N_5030,In_2916,In_4708);
and U5031 (N_5031,In_675,In_4966);
nand U5032 (N_5032,In_3083,In_66);
nand U5033 (N_5033,In_4578,In_1213);
or U5034 (N_5034,In_3072,In_4310);
or U5035 (N_5035,In_3830,In_4785);
nand U5036 (N_5036,In_2479,In_1692);
nor U5037 (N_5037,In_2567,In_1209);
or U5038 (N_5038,In_2497,In_716);
nand U5039 (N_5039,In_1158,In_1497);
nand U5040 (N_5040,In_4514,In_2544);
and U5041 (N_5041,In_1581,In_2321);
nor U5042 (N_5042,In_4874,In_4240);
or U5043 (N_5043,In_860,In_2281);
nand U5044 (N_5044,In_4178,In_4908);
or U5045 (N_5045,In_2232,In_1370);
or U5046 (N_5046,In_1929,In_1691);
nand U5047 (N_5047,In_2,In_2228);
and U5048 (N_5048,In_4796,In_1037);
or U5049 (N_5049,In_1595,In_1099);
nand U5050 (N_5050,In_113,In_4234);
or U5051 (N_5051,In_2612,In_4347);
and U5052 (N_5052,In_75,In_3023);
or U5053 (N_5053,In_4186,In_3932);
and U5054 (N_5054,In_4115,In_4717);
and U5055 (N_5055,In_2702,In_1519);
or U5056 (N_5056,In_3482,In_3274);
xnor U5057 (N_5057,In_814,In_2666);
and U5058 (N_5058,In_671,In_2376);
nand U5059 (N_5059,In_3081,In_980);
xnor U5060 (N_5060,In_3156,In_4966);
or U5061 (N_5061,In_1892,In_600);
nor U5062 (N_5062,In_3754,In_1015);
and U5063 (N_5063,In_1164,In_2169);
xor U5064 (N_5064,In_4110,In_4095);
and U5065 (N_5065,In_298,In_412);
nand U5066 (N_5066,In_1195,In_2536);
nand U5067 (N_5067,In_4451,In_4926);
or U5068 (N_5068,In_2615,In_65);
and U5069 (N_5069,In_100,In_2659);
or U5070 (N_5070,In_3840,In_285);
xor U5071 (N_5071,In_4375,In_289);
nor U5072 (N_5072,In_3962,In_4139);
nand U5073 (N_5073,In_2372,In_4940);
and U5074 (N_5074,In_841,In_74);
or U5075 (N_5075,In_26,In_1480);
and U5076 (N_5076,In_1322,In_3256);
xnor U5077 (N_5077,In_3233,In_296);
and U5078 (N_5078,In_2757,In_1168);
nand U5079 (N_5079,In_2168,In_2150);
and U5080 (N_5080,In_1488,In_3047);
and U5081 (N_5081,In_4563,In_2484);
or U5082 (N_5082,In_4117,In_4878);
and U5083 (N_5083,In_4505,In_2748);
or U5084 (N_5084,In_362,In_454);
nand U5085 (N_5085,In_2948,In_3239);
xnor U5086 (N_5086,In_2560,In_2003);
and U5087 (N_5087,In_1291,In_4246);
or U5088 (N_5088,In_1024,In_2824);
xnor U5089 (N_5089,In_4689,In_4780);
nor U5090 (N_5090,In_668,In_327);
or U5091 (N_5091,In_549,In_1621);
and U5092 (N_5092,In_3821,In_329);
or U5093 (N_5093,In_2614,In_4760);
or U5094 (N_5094,In_3661,In_2483);
or U5095 (N_5095,In_1387,In_923);
or U5096 (N_5096,In_4150,In_565);
nand U5097 (N_5097,In_1385,In_3108);
or U5098 (N_5098,In_854,In_3558);
and U5099 (N_5099,In_3082,In_4602);
and U5100 (N_5100,In_836,In_3508);
and U5101 (N_5101,In_1704,In_2511);
and U5102 (N_5102,In_541,In_1506);
or U5103 (N_5103,In_996,In_193);
or U5104 (N_5104,In_4297,In_4929);
nand U5105 (N_5105,In_3071,In_2681);
or U5106 (N_5106,In_3246,In_3222);
nor U5107 (N_5107,In_3543,In_1159);
and U5108 (N_5108,In_2853,In_2446);
or U5109 (N_5109,In_2787,In_1966);
nand U5110 (N_5110,In_4055,In_1800);
or U5111 (N_5111,In_117,In_1404);
and U5112 (N_5112,In_4037,In_3421);
and U5113 (N_5113,In_1439,In_794);
or U5114 (N_5114,In_3896,In_4393);
nand U5115 (N_5115,In_213,In_2661);
nor U5116 (N_5116,In_2605,In_696);
or U5117 (N_5117,In_3065,In_1339);
nand U5118 (N_5118,In_1322,In_4410);
nor U5119 (N_5119,In_4821,In_4792);
and U5120 (N_5120,In_4185,In_1376);
and U5121 (N_5121,In_4559,In_3789);
nand U5122 (N_5122,In_2408,In_1363);
nor U5123 (N_5123,In_2697,In_1869);
or U5124 (N_5124,In_2639,In_1740);
nor U5125 (N_5125,In_1865,In_4567);
or U5126 (N_5126,In_229,In_4973);
and U5127 (N_5127,In_310,In_3180);
xnor U5128 (N_5128,In_4501,In_1662);
or U5129 (N_5129,In_4606,In_1889);
nor U5130 (N_5130,In_235,In_2653);
nor U5131 (N_5131,In_3207,In_3809);
and U5132 (N_5132,In_4850,In_4662);
and U5133 (N_5133,In_968,In_129);
nand U5134 (N_5134,In_1642,In_1440);
nor U5135 (N_5135,In_2100,In_1956);
and U5136 (N_5136,In_4092,In_4332);
and U5137 (N_5137,In_4005,In_1635);
or U5138 (N_5138,In_3560,In_2281);
nand U5139 (N_5139,In_3037,In_1503);
nor U5140 (N_5140,In_1430,In_594);
or U5141 (N_5141,In_3852,In_2375);
xnor U5142 (N_5142,In_3219,In_4537);
or U5143 (N_5143,In_1047,In_957);
xnor U5144 (N_5144,In_3597,In_4972);
and U5145 (N_5145,In_3057,In_1061);
or U5146 (N_5146,In_4859,In_1529);
and U5147 (N_5147,In_4032,In_4214);
xor U5148 (N_5148,In_781,In_1732);
nand U5149 (N_5149,In_4621,In_647);
nor U5150 (N_5150,In_3625,In_4476);
nand U5151 (N_5151,In_4586,In_3788);
nor U5152 (N_5152,In_1421,In_2780);
nor U5153 (N_5153,In_4779,In_4451);
nor U5154 (N_5154,In_1656,In_625);
xor U5155 (N_5155,In_4700,In_4606);
nor U5156 (N_5156,In_3241,In_2727);
nor U5157 (N_5157,In_2771,In_397);
and U5158 (N_5158,In_4779,In_248);
and U5159 (N_5159,In_2600,In_1311);
and U5160 (N_5160,In_3635,In_3311);
nor U5161 (N_5161,In_1299,In_4472);
or U5162 (N_5162,In_4826,In_2644);
or U5163 (N_5163,In_2818,In_4241);
xnor U5164 (N_5164,In_4830,In_2088);
or U5165 (N_5165,In_4487,In_3845);
nor U5166 (N_5166,In_3038,In_4593);
and U5167 (N_5167,In_3931,In_1283);
nand U5168 (N_5168,In_4978,In_3546);
nand U5169 (N_5169,In_3664,In_2426);
or U5170 (N_5170,In_4605,In_1522);
or U5171 (N_5171,In_2381,In_3790);
xnor U5172 (N_5172,In_304,In_3512);
and U5173 (N_5173,In_6,In_2955);
nor U5174 (N_5174,In_2778,In_318);
nand U5175 (N_5175,In_4364,In_4995);
nor U5176 (N_5176,In_3503,In_4650);
nor U5177 (N_5177,In_525,In_3122);
xnor U5178 (N_5178,In_4563,In_912);
nand U5179 (N_5179,In_4770,In_41);
nand U5180 (N_5180,In_962,In_3096);
nand U5181 (N_5181,In_1197,In_1365);
and U5182 (N_5182,In_1813,In_2666);
and U5183 (N_5183,In_4687,In_2545);
xor U5184 (N_5184,In_3616,In_4466);
nand U5185 (N_5185,In_2011,In_4435);
nand U5186 (N_5186,In_1346,In_2803);
xnor U5187 (N_5187,In_4100,In_2984);
xnor U5188 (N_5188,In_4787,In_1565);
xor U5189 (N_5189,In_2051,In_2464);
or U5190 (N_5190,In_626,In_3841);
nand U5191 (N_5191,In_4577,In_2017);
or U5192 (N_5192,In_1873,In_4240);
or U5193 (N_5193,In_3847,In_1060);
and U5194 (N_5194,In_3415,In_99);
or U5195 (N_5195,In_1356,In_4964);
or U5196 (N_5196,In_3287,In_3704);
and U5197 (N_5197,In_4388,In_4639);
nor U5198 (N_5198,In_3361,In_4750);
nor U5199 (N_5199,In_591,In_779);
xnor U5200 (N_5200,In_4117,In_3741);
and U5201 (N_5201,In_2039,In_3022);
nor U5202 (N_5202,In_4148,In_3817);
nor U5203 (N_5203,In_4427,In_4148);
and U5204 (N_5204,In_3939,In_1786);
nand U5205 (N_5205,In_931,In_1967);
nand U5206 (N_5206,In_2122,In_4041);
nor U5207 (N_5207,In_1540,In_421);
and U5208 (N_5208,In_4940,In_377);
nand U5209 (N_5209,In_447,In_4982);
and U5210 (N_5210,In_2787,In_3572);
nor U5211 (N_5211,In_3386,In_2225);
and U5212 (N_5212,In_224,In_4387);
and U5213 (N_5213,In_1421,In_3276);
and U5214 (N_5214,In_3651,In_3775);
xnor U5215 (N_5215,In_1004,In_426);
nor U5216 (N_5216,In_3146,In_4882);
or U5217 (N_5217,In_415,In_183);
and U5218 (N_5218,In_2714,In_3307);
xnor U5219 (N_5219,In_154,In_1912);
and U5220 (N_5220,In_1151,In_3380);
nand U5221 (N_5221,In_2184,In_1201);
or U5222 (N_5222,In_2220,In_4064);
or U5223 (N_5223,In_690,In_4548);
nand U5224 (N_5224,In_4502,In_1251);
and U5225 (N_5225,In_130,In_3489);
nor U5226 (N_5226,In_1355,In_2508);
nand U5227 (N_5227,In_2548,In_185);
and U5228 (N_5228,In_1004,In_3614);
and U5229 (N_5229,In_3842,In_2400);
or U5230 (N_5230,In_759,In_4439);
nand U5231 (N_5231,In_3514,In_2622);
nor U5232 (N_5232,In_661,In_3270);
nor U5233 (N_5233,In_3257,In_4777);
and U5234 (N_5234,In_477,In_4600);
nand U5235 (N_5235,In_4806,In_416);
xnor U5236 (N_5236,In_4107,In_3182);
nand U5237 (N_5237,In_3876,In_2330);
nor U5238 (N_5238,In_47,In_2611);
or U5239 (N_5239,In_1089,In_3237);
and U5240 (N_5240,In_2491,In_1247);
or U5241 (N_5241,In_355,In_4330);
nand U5242 (N_5242,In_1573,In_2013);
nand U5243 (N_5243,In_824,In_2669);
nor U5244 (N_5244,In_2823,In_2586);
xor U5245 (N_5245,In_941,In_4959);
and U5246 (N_5246,In_1591,In_701);
or U5247 (N_5247,In_4263,In_3018);
nand U5248 (N_5248,In_1470,In_4446);
nor U5249 (N_5249,In_4112,In_71);
nand U5250 (N_5250,In_394,In_822);
xor U5251 (N_5251,In_2250,In_4833);
nor U5252 (N_5252,In_1913,In_4441);
nand U5253 (N_5253,In_4353,In_2743);
nor U5254 (N_5254,In_3318,In_648);
or U5255 (N_5255,In_1830,In_325);
or U5256 (N_5256,In_248,In_1297);
and U5257 (N_5257,In_1147,In_4603);
nand U5258 (N_5258,In_4534,In_746);
nand U5259 (N_5259,In_1442,In_3756);
nor U5260 (N_5260,In_3623,In_3630);
or U5261 (N_5261,In_3142,In_49);
and U5262 (N_5262,In_4210,In_2994);
or U5263 (N_5263,In_4703,In_3047);
nand U5264 (N_5264,In_75,In_1698);
nor U5265 (N_5265,In_1000,In_661);
and U5266 (N_5266,In_1613,In_189);
nor U5267 (N_5267,In_1641,In_160);
nand U5268 (N_5268,In_4072,In_1531);
or U5269 (N_5269,In_4684,In_4961);
or U5270 (N_5270,In_391,In_467);
nand U5271 (N_5271,In_2762,In_4905);
nor U5272 (N_5272,In_196,In_2175);
nand U5273 (N_5273,In_1307,In_1251);
or U5274 (N_5274,In_3844,In_2585);
or U5275 (N_5275,In_2558,In_2144);
nor U5276 (N_5276,In_512,In_3443);
nor U5277 (N_5277,In_1162,In_2746);
or U5278 (N_5278,In_286,In_284);
or U5279 (N_5279,In_4862,In_4860);
nor U5280 (N_5280,In_1994,In_3062);
xnor U5281 (N_5281,In_3168,In_3335);
nor U5282 (N_5282,In_674,In_137);
and U5283 (N_5283,In_3197,In_3467);
nand U5284 (N_5284,In_2538,In_2302);
and U5285 (N_5285,In_4792,In_918);
nor U5286 (N_5286,In_4268,In_3788);
nor U5287 (N_5287,In_2299,In_2437);
nor U5288 (N_5288,In_1647,In_2585);
and U5289 (N_5289,In_2660,In_929);
nand U5290 (N_5290,In_911,In_4082);
or U5291 (N_5291,In_2850,In_2088);
xnor U5292 (N_5292,In_1544,In_2336);
and U5293 (N_5293,In_1175,In_3968);
and U5294 (N_5294,In_2199,In_720);
and U5295 (N_5295,In_1047,In_721);
nand U5296 (N_5296,In_4489,In_892);
or U5297 (N_5297,In_1182,In_3759);
or U5298 (N_5298,In_3953,In_407);
or U5299 (N_5299,In_4002,In_2873);
nand U5300 (N_5300,In_4503,In_3860);
nand U5301 (N_5301,In_3816,In_2043);
xor U5302 (N_5302,In_3716,In_1035);
or U5303 (N_5303,In_2913,In_1095);
or U5304 (N_5304,In_4797,In_4950);
nor U5305 (N_5305,In_3100,In_4467);
and U5306 (N_5306,In_4421,In_2689);
nand U5307 (N_5307,In_1949,In_323);
nand U5308 (N_5308,In_4221,In_1384);
xnor U5309 (N_5309,In_1038,In_831);
nand U5310 (N_5310,In_4175,In_2991);
and U5311 (N_5311,In_3930,In_1879);
xor U5312 (N_5312,In_4042,In_2953);
nor U5313 (N_5313,In_522,In_3576);
and U5314 (N_5314,In_1792,In_1145);
and U5315 (N_5315,In_3291,In_1920);
xnor U5316 (N_5316,In_3653,In_3430);
or U5317 (N_5317,In_1320,In_1514);
nor U5318 (N_5318,In_1894,In_2432);
and U5319 (N_5319,In_744,In_3829);
or U5320 (N_5320,In_3939,In_893);
nor U5321 (N_5321,In_3347,In_4764);
and U5322 (N_5322,In_1757,In_3799);
nor U5323 (N_5323,In_1901,In_2307);
and U5324 (N_5324,In_1802,In_3859);
nor U5325 (N_5325,In_2933,In_1056);
and U5326 (N_5326,In_1003,In_1956);
or U5327 (N_5327,In_614,In_1566);
xor U5328 (N_5328,In_88,In_2606);
or U5329 (N_5329,In_3648,In_1319);
or U5330 (N_5330,In_2675,In_1372);
and U5331 (N_5331,In_1994,In_622);
nor U5332 (N_5332,In_2510,In_1949);
nor U5333 (N_5333,In_3815,In_3782);
and U5334 (N_5334,In_1463,In_3683);
nand U5335 (N_5335,In_2983,In_4094);
and U5336 (N_5336,In_4736,In_2536);
or U5337 (N_5337,In_4613,In_659);
or U5338 (N_5338,In_4994,In_3793);
or U5339 (N_5339,In_995,In_1905);
and U5340 (N_5340,In_4801,In_392);
nor U5341 (N_5341,In_2637,In_2368);
and U5342 (N_5342,In_4175,In_4493);
nand U5343 (N_5343,In_315,In_3598);
nand U5344 (N_5344,In_2874,In_4468);
nor U5345 (N_5345,In_1005,In_4850);
or U5346 (N_5346,In_4789,In_1781);
or U5347 (N_5347,In_284,In_2780);
and U5348 (N_5348,In_3232,In_4431);
nor U5349 (N_5349,In_667,In_3018);
or U5350 (N_5350,In_1127,In_4876);
nor U5351 (N_5351,In_566,In_2599);
nor U5352 (N_5352,In_3950,In_130);
or U5353 (N_5353,In_380,In_1184);
nand U5354 (N_5354,In_2893,In_3654);
nor U5355 (N_5355,In_1330,In_3057);
nand U5356 (N_5356,In_2807,In_2793);
nor U5357 (N_5357,In_1660,In_4549);
or U5358 (N_5358,In_4599,In_1383);
nand U5359 (N_5359,In_3792,In_3467);
nand U5360 (N_5360,In_4368,In_3391);
and U5361 (N_5361,In_2644,In_3280);
nor U5362 (N_5362,In_4360,In_1824);
xor U5363 (N_5363,In_344,In_4787);
and U5364 (N_5364,In_619,In_399);
nor U5365 (N_5365,In_4045,In_3604);
nor U5366 (N_5366,In_338,In_4923);
or U5367 (N_5367,In_2186,In_244);
nand U5368 (N_5368,In_4662,In_3288);
and U5369 (N_5369,In_539,In_3194);
nand U5370 (N_5370,In_2908,In_4125);
and U5371 (N_5371,In_4785,In_598);
nand U5372 (N_5372,In_2987,In_1763);
or U5373 (N_5373,In_2675,In_4251);
nor U5374 (N_5374,In_4089,In_3482);
nand U5375 (N_5375,In_368,In_4110);
and U5376 (N_5376,In_3583,In_4275);
nor U5377 (N_5377,In_2754,In_4150);
nand U5378 (N_5378,In_3831,In_2806);
nor U5379 (N_5379,In_3989,In_4316);
nand U5380 (N_5380,In_3729,In_4411);
nor U5381 (N_5381,In_4131,In_2666);
nand U5382 (N_5382,In_732,In_316);
nand U5383 (N_5383,In_155,In_597);
and U5384 (N_5384,In_229,In_4691);
xnor U5385 (N_5385,In_4381,In_3321);
nor U5386 (N_5386,In_34,In_2353);
and U5387 (N_5387,In_73,In_4811);
and U5388 (N_5388,In_541,In_2710);
nor U5389 (N_5389,In_1726,In_4134);
and U5390 (N_5390,In_2007,In_1149);
nor U5391 (N_5391,In_437,In_55);
nor U5392 (N_5392,In_3598,In_641);
or U5393 (N_5393,In_533,In_1996);
nor U5394 (N_5394,In_4533,In_967);
or U5395 (N_5395,In_4115,In_1617);
or U5396 (N_5396,In_3080,In_2485);
xnor U5397 (N_5397,In_4929,In_4355);
nand U5398 (N_5398,In_611,In_3327);
nor U5399 (N_5399,In_4892,In_1056);
nand U5400 (N_5400,In_4546,In_479);
nor U5401 (N_5401,In_2327,In_4792);
or U5402 (N_5402,In_3010,In_695);
nor U5403 (N_5403,In_2082,In_70);
or U5404 (N_5404,In_4116,In_3725);
nor U5405 (N_5405,In_4467,In_1566);
xnor U5406 (N_5406,In_880,In_2776);
nand U5407 (N_5407,In_1250,In_4186);
xor U5408 (N_5408,In_1599,In_1872);
nand U5409 (N_5409,In_3580,In_3085);
nand U5410 (N_5410,In_4536,In_3395);
and U5411 (N_5411,In_2432,In_4734);
nand U5412 (N_5412,In_4692,In_7);
and U5413 (N_5413,In_2389,In_1493);
nand U5414 (N_5414,In_2494,In_2705);
nand U5415 (N_5415,In_1499,In_2073);
nor U5416 (N_5416,In_555,In_790);
nor U5417 (N_5417,In_866,In_3243);
nor U5418 (N_5418,In_2577,In_2226);
xor U5419 (N_5419,In_2889,In_4227);
xor U5420 (N_5420,In_537,In_907);
or U5421 (N_5421,In_2548,In_191);
or U5422 (N_5422,In_3249,In_1292);
nand U5423 (N_5423,In_4030,In_880);
nor U5424 (N_5424,In_4097,In_1688);
xnor U5425 (N_5425,In_497,In_2368);
and U5426 (N_5426,In_4497,In_354);
nor U5427 (N_5427,In_965,In_2219);
nor U5428 (N_5428,In_686,In_3340);
or U5429 (N_5429,In_370,In_4510);
nor U5430 (N_5430,In_2748,In_4682);
and U5431 (N_5431,In_2285,In_4827);
and U5432 (N_5432,In_2560,In_2854);
nor U5433 (N_5433,In_2655,In_1445);
nor U5434 (N_5434,In_15,In_1086);
nand U5435 (N_5435,In_1246,In_212);
nand U5436 (N_5436,In_2324,In_286);
nor U5437 (N_5437,In_1913,In_1300);
nand U5438 (N_5438,In_2830,In_4643);
nor U5439 (N_5439,In_694,In_1525);
xor U5440 (N_5440,In_982,In_2396);
nand U5441 (N_5441,In_4478,In_2665);
nand U5442 (N_5442,In_3222,In_3482);
xnor U5443 (N_5443,In_2,In_3907);
nor U5444 (N_5444,In_683,In_3586);
and U5445 (N_5445,In_3048,In_975);
nor U5446 (N_5446,In_4366,In_4458);
and U5447 (N_5447,In_4161,In_2590);
and U5448 (N_5448,In_3504,In_2450);
and U5449 (N_5449,In_4581,In_1553);
nor U5450 (N_5450,In_1757,In_4357);
nor U5451 (N_5451,In_3959,In_174);
nor U5452 (N_5452,In_1347,In_1252);
or U5453 (N_5453,In_4813,In_4227);
or U5454 (N_5454,In_2741,In_4626);
nand U5455 (N_5455,In_2276,In_4968);
nor U5456 (N_5456,In_4073,In_1402);
and U5457 (N_5457,In_3498,In_4929);
nor U5458 (N_5458,In_880,In_4462);
nor U5459 (N_5459,In_84,In_1408);
or U5460 (N_5460,In_4906,In_1635);
nor U5461 (N_5461,In_532,In_475);
and U5462 (N_5462,In_355,In_3842);
nor U5463 (N_5463,In_352,In_4244);
nand U5464 (N_5464,In_1062,In_1044);
nand U5465 (N_5465,In_3759,In_117);
nor U5466 (N_5466,In_2243,In_3533);
nand U5467 (N_5467,In_1653,In_358);
and U5468 (N_5468,In_1742,In_510);
nor U5469 (N_5469,In_724,In_150);
nand U5470 (N_5470,In_3461,In_2936);
nor U5471 (N_5471,In_4064,In_4926);
and U5472 (N_5472,In_2818,In_2741);
nand U5473 (N_5473,In_1870,In_2253);
nand U5474 (N_5474,In_3453,In_2634);
xnor U5475 (N_5475,In_1629,In_1228);
nand U5476 (N_5476,In_2910,In_2739);
nor U5477 (N_5477,In_1479,In_4827);
nand U5478 (N_5478,In_485,In_2691);
and U5479 (N_5479,In_4453,In_4960);
and U5480 (N_5480,In_3125,In_4956);
nand U5481 (N_5481,In_4838,In_1479);
nand U5482 (N_5482,In_3129,In_2832);
or U5483 (N_5483,In_557,In_2315);
nor U5484 (N_5484,In_1572,In_3218);
nand U5485 (N_5485,In_3501,In_3359);
and U5486 (N_5486,In_4355,In_1534);
nor U5487 (N_5487,In_2692,In_3155);
and U5488 (N_5488,In_4557,In_188);
and U5489 (N_5489,In_4053,In_12);
nor U5490 (N_5490,In_1220,In_1033);
and U5491 (N_5491,In_1880,In_2586);
xor U5492 (N_5492,In_243,In_3247);
nor U5493 (N_5493,In_2446,In_3984);
or U5494 (N_5494,In_3469,In_2777);
and U5495 (N_5495,In_3591,In_4731);
or U5496 (N_5496,In_3208,In_3642);
and U5497 (N_5497,In_1867,In_3607);
and U5498 (N_5498,In_358,In_4252);
nor U5499 (N_5499,In_4941,In_2325);
or U5500 (N_5500,In_722,In_421);
and U5501 (N_5501,In_105,In_1388);
nor U5502 (N_5502,In_3510,In_2728);
and U5503 (N_5503,In_1135,In_1333);
nor U5504 (N_5504,In_1183,In_1971);
nor U5505 (N_5505,In_207,In_2062);
and U5506 (N_5506,In_3158,In_776);
nand U5507 (N_5507,In_2069,In_4096);
nand U5508 (N_5508,In_1047,In_3067);
or U5509 (N_5509,In_3762,In_855);
and U5510 (N_5510,In_2052,In_2265);
nor U5511 (N_5511,In_3541,In_765);
and U5512 (N_5512,In_2227,In_2484);
nand U5513 (N_5513,In_1128,In_3714);
nand U5514 (N_5514,In_3715,In_4511);
nor U5515 (N_5515,In_4591,In_4096);
nor U5516 (N_5516,In_4102,In_2126);
xnor U5517 (N_5517,In_4114,In_4257);
nand U5518 (N_5518,In_3417,In_2368);
or U5519 (N_5519,In_2856,In_758);
nor U5520 (N_5520,In_845,In_4104);
nand U5521 (N_5521,In_1057,In_2975);
xnor U5522 (N_5522,In_377,In_1336);
and U5523 (N_5523,In_3621,In_3888);
nand U5524 (N_5524,In_736,In_1976);
nor U5525 (N_5525,In_1812,In_2768);
nand U5526 (N_5526,In_2097,In_2821);
or U5527 (N_5527,In_1820,In_3987);
nand U5528 (N_5528,In_4805,In_613);
and U5529 (N_5529,In_145,In_1928);
nor U5530 (N_5530,In_1153,In_4712);
nor U5531 (N_5531,In_2731,In_3712);
nor U5532 (N_5532,In_3037,In_2929);
or U5533 (N_5533,In_1645,In_80);
nor U5534 (N_5534,In_4574,In_1280);
nand U5535 (N_5535,In_1950,In_3218);
nor U5536 (N_5536,In_3102,In_3387);
nor U5537 (N_5537,In_4516,In_1115);
nor U5538 (N_5538,In_531,In_2219);
nor U5539 (N_5539,In_2583,In_2889);
nand U5540 (N_5540,In_4531,In_1868);
nand U5541 (N_5541,In_2411,In_2870);
xor U5542 (N_5542,In_390,In_1437);
nand U5543 (N_5543,In_3925,In_1438);
nand U5544 (N_5544,In_1010,In_4673);
and U5545 (N_5545,In_850,In_1369);
and U5546 (N_5546,In_2900,In_568);
or U5547 (N_5547,In_1470,In_4943);
or U5548 (N_5548,In_3797,In_1001);
nand U5549 (N_5549,In_768,In_381);
nor U5550 (N_5550,In_1746,In_151);
and U5551 (N_5551,In_2416,In_2330);
nor U5552 (N_5552,In_3516,In_1655);
and U5553 (N_5553,In_2308,In_1744);
xnor U5554 (N_5554,In_1334,In_3042);
or U5555 (N_5555,In_4182,In_4348);
nor U5556 (N_5556,In_4738,In_4181);
xor U5557 (N_5557,In_17,In_3384);
nor U5558 (N_5558,In_513,In_4112);
and U5559 (N_5559,In_3577,In_2004);
nand U5560 (N_5560,In_2972,In_948);
nand U5561 (N_5561,In_3641,In_3595);
nand U5562 (N_5562,In_3316,In_4786);
or U5563 (N_5563,In_1260,In_4718);
or U5564 (N_5564,In_2693,In_2113);
and U5565 (N_5565,In_3932,In_981);
nand U5566 (N_5566,In_2130,In_2326);
nand U5567 (N_5567,In_4424,In_4560);
xnor U5568 (N_5568,In_773,In_3751);
and U5569 (N_5569,In_244,In_3592);
or U5570 (N_5570,In_1608,In_4100);
and U5571 (N_5571,In_1366,In_2347);
or U5572 (N_5572,In_85,In_3177);
or U5573 (N_5573,In_3114,In_1379);
nor U5574 (N_5574,In_3911,In_1661);
nor U5575 (N_5575,In_2181,In_2634);
nand U5576 (N_5576,In_296,In_3533);
and U5577 (N_5577,In_4115,In_2165);
or U5578 (N_5578,In_1245,In_2694);
or U5579 (N_5579,In_235,In_229);
nor U5580 (N_5580,In_4062,In_2444);
nor U5581 (N_5581,In_90,In_2561);
or U5582 (N_5582,In_4158,In_2116);
xnor U5583 (N_5583,In_53,In_4782);
nor U5584 (N_5584,In_1966,In_749);
nor U5585 (N_5585,In_1096,In_2544);
nor U5586 (N_5586,In_2432,In_1363);
nand U5587 (N_5587,In_3873,In_2146);
xnor U5588 (N_5588,In_4101,In_4354);
and U5589 (N_5589,In_2526,In_4439);
nand U5590 (N_5590,In_2509,In_1444);
nor U5591 (N_5591,In_55,In_244);
nor U5592 (N_5592,In_4878,In_2700);
and U5593 (N_5593,In_595,In_1371);
nor U5594 (N_5594,In_3483,In_2238);
or U5595 (N_5595,In_2377,In_2221);
and U5596 (N_5596,In_4990,In_4862);
nand U5597 (N_5597,In_1654,In_1299);
nor U5598 (N_5598,In_2273,In_3995);
and U5599 (N_5599,In_3582,In_2105);
xor U5600 (N_5600,In_4705,In_4982);
or U5601 (N_5601,In_1415,In_1809);
or U5602 (N_5602,In_668,In_3972);
nor U5603 (N_5603,In_2506,In_1983);
or U5604 (N_5604,In_1538,In_322);
nand U5605 (N_5605,In_977,In_4038);
xor U5606 (N_5606,In_3144,In_3705);
nand U5607 (N_5607,In_1780,In_2061);
and U5608 (N_5608,In_2694,In_3274);
nand U5609 (N_5609,In_760,In_3860);
or U5610 (N_5610,In_4449,In_3512);
nand U5611 (N_5611,In_203,In_1678);
and U5612 (N_5612,In_3946,In_588);
nand U5613 (N_5613,In_1446,In_534);
and U5614 (N_5614,In_2964,In_533);
nand U5615 (N_5615,In_3176,In_4374);
nor U5616 (N_5616,In_1116,In_4106);
nand U5617 (N_5617,In_3423,In_3421);
nand U5618 (N_5618,In_1985,In_2880);
or U5619 (N_5619,In_4565,In_3497);
xor U5620 (N_5620,In_3633,In_2043);
nand U5621 (N_5621,In_3152,In_1295);
nand U5622 (N_5622,In_2658,In_141);
and U5623 (N_5623,In_398,In_865);
and U5624 (N_5624,In_4302,In_1134);
nand U5625 (N_5625,In_3659,In_825);
nand U5626 (N_5626,In_3561,In_2165);
xnor U5627 (N_5627,In_3739,In_2549);
or U5628 (N_5628,In_3373,In_4070);
nor U5629 (N_5629,In_4124,In_935);
or U5630 (N_5630,In_1680,In_3332);
nor U5631 (N_5631,In_2071,In_35);
nor U5632 (N_5632,In_1348,In_1321);
nand U5633 (N_5633,In_3321,In_816);
nand U5634 (N_5634,In_1444,In_928);
nor U5635 (N_5635,In_1368,In_4124);
xor U5636 (N_5636,In_2048,In_353);
or U5637 (N_5637,In_3038,In_1808);
and U5638 (N_5638,In_981,In_4603);
nand U5639 (N_5639,In_237,In_4730);
nor U5640 (N_5640,In_4673,In_2158);
or U5641 (N_5641,In_1290,In_1375);
nor U5642 (N_5642,In_2779,In_2961);
and U5643 (N_5643,In_4696,In_3953);
or U5644 (N_5644,In_1794,In_4007);
or U5645 (N_5645,In_3899,In_3446);
xnor U5646 (N_5646,In_2852,In_4278);
and U5647 (N_5647,In_2232,In_941);
and U5648 (N_5648,In_685,In_4094);
and U5649 (N_5649,In_2538,In_3382);
xnor U5650 (N_5650,In_1018,In_1894);
xnor U5651 (N_5651,In_2439,In_96);
or U5652 (N_5652,In_1161,In_4683);
or U5653 (N_5653,In_2912,In_2678);
or U5654 (N_5654,In_878,In_3904);
or U5655 (N_5655,In_659,In_122);
and U5656 (N_5656,In_2786,In_4448);
xnor U5657 (N_5657,In_1646,In_2247);
xnor U5658 (N_5658,In_2698,In_3409);
xnor U5659 (N_5659,In_3347,In_578);
nor U5660 (N_5660,In_2304,In_64);
nor U5661 (N_5661,In_4062,In_4806);
nor U5662 (N_5662,In_3454,In_3549);
nor U5663 (N_5663,In_17,In_3064);
nor U5664 (N_5664,In_4421,In_3688);
xnor U5665 (N_5665,In_2325,In_2741);
and U5666 (N_5666,In_109,In_3871);
xor U5667 (N_5667,In_3029,In_236);
and U5668 (N_5668,In_494,In_3102);
nand U5669 (N_5669,In_1457,In_1342);
and U5670 (N_5670,In_2725,In_3326);
or U5671 (N_5671,In_317,In_3604);
nand U5672 (N_5672,In_1627,In_2622);
nand U5673 (N_5673,In_1524,In_711);
or U5674 (N_5674,In_3294,In_4836);
nor U5675 (N_5675,In_3079,In_1305);
nand U5676 (N_5676,In_2000,In_3835);
or U5677 (N_5677,In_4222,In_2073);
or U5678 (N_5678,In_2383,In_3974);
nand U5679 (N_5679,In_553,In_372);
and U5680 (N_5680,In_1982,In_565);
and U5681 (N_5681,In_86,In_4093);
nand U5682 (N_5682,In_2788,In_3490);
or U5683 (N_5683,In_4882,In_1891);
and U5684 (N_5684,In_3128,In_3005);
or U5685 (N_5685,In_4871,In_1709);
nor U5686 (N_5686,In_1139,In_1706);
and U5687 (N_5687,In_4802,In_4820);
and U5688 (N_5688,In_3507,In_1456);
nand U5689 (N_5689,In_4385,In_3195);
nand U5690 (N_5690,In_3489,In_1717);
or U5691 (N_5691,In_965,In_391);
xor U5692 (N_5692,In_1329,In_3907);
nand U5693 (N_5693,In_4919,In_4908);
and U5694 (N_5694,In_1812,In_3082);
or U5695 (N_5695,In_3586,In_1681);
and U5696 (N_5696,In_437,In_4784);
and U5697 (N_5697,In_2683,In_3759);
or U5698 (N_5698,In_4010,In_1907);
and U5699 (N_5699,In_1191,In_3438);
and U5700 (N_5700,In_2638,In_2722);
and U5701 (N_5701,In_3435,In_2305);
or U5702 (N_5702,In_1792,In_1025);
or U5703 (N_5703,In_3945,In_1407);
or U5704 (N_5704,In_2197,In_588);
nand U5705 (N_5705,In_1795,In_2052);
nor U5706 (N_5706,In_2476,In_673);
and U5707 (N_5707,In_2967,In_2329);
or U5708 (N_5708,In_4702,In_23);
and U5709 (N_5709,In_249,In_3730);
and U5710 (N_5710,In_4765,In_1685);
nand U5711 (N_5711,In_1920,In_3481);
or U5712 (N_5712,In_4186,In_1909);
nand U5713 (N_5713,In_447,In_3279);
xnor U5714 (N_5714,In_781,In_4791);
nor U5715 (N_5715,In_1191,In_4122);
nor U5716 (N_5716,In_1790,In_1924);
nor U5717 (N_5717,In_2797,In_2839);
nand U5718 (N_5718,In_92,In_363);
nor U5719 (N_5719,In_383,In_191);
and U5720 (N_5720,In_728,In_437);
nand U5721 (N_5721,In_3728,In_641);
or U5722 (N_5722,In_2988,In_2845);
and U5723 (N_5723,In_4952,In_212);
xor U5724 (N_5724,In_2097,In_3894);
nand U5725 (N_5725,In_4732,In_2058);
xnor U5726 (N_5726,In_4976,In_4245);
or U5727 (N_5727,In_68,In_2780);
nor U5728 (N_5728,In_4748,In_3367);
xor U5729 (N_5729,In_1128,In_584);
and U5730 (N_5730,In_549,In_3410);
and U5731 (N_5731,In_1307,In_3467);
and U5732 (N_5732,In_2423,In_723);
nand U5733 (N_5733,In_1853,In_3770);
or U5734 (N_5734,In_4253,In_570);
nor U5735 (N_5735,In_1735,In_1386);
or U5736 (N_5736,In_1327,In_4618);
nor U5737 (N_5737,In_4641,In_2954);
xnor U5738 (N_5738,In_1639,In_869);
nand U5739 (N_5739,In_1145,In_1695);
nor U5740 (N_5740,In_4120,In_1384);
nand U5741 (N_5741,In_353,In_2179);
nand U5742 (N_5742,In_3699,In_2190);
or U5743 (N_5743,In_3312,In_1616);
nor U5744 (N_5744,In_2523,In_2645);
nor U5745 (N_5745,In_1523,In_1291);
and U5746 (N_5746,In_146,In_816);
nor U5747 (N_5747,In_4118,In_414);
and U5748 (N_5748,In_3475,In_4746);
and U5749 (N_5749,In_4863,In_830);
or U5750 (N_5750,In_4397,In_2003);
nand U5751 (N_5751,In_3436,In_1159);
nor U5752 (N_5752,In_1677,In_2);
nand U5753 (N_5753,In_3352,In_1457);
nor U5754 (N_5754,In_3073,In_1596);
nand U5755 (N_5755,In_1272,In_996);
nand U5756 (N_5756,In_2860,In_2257);
nor U5757 (N_5757,In_2161,In_1106);
xnor U5758 (N_5758,In_1037,In_806);
or U5759 (N_5759,In_75,In_2056);
nand U5760 (N_5760,In_3639,In_4590);
and U5761 (N_5761,In_968,In_4915);
or U5762 (N_5762,In_3484,In_4597);
or U5763 (N_5763,In_1656,In_1561);
and U5764 (N_5764,In_1813,In_936);
nand U5765 (N_5765,In_4747,In_4807);
or U5766 (N_5766,In_1418,In_2054);
and U5767 (N_5767,In_4567,In_3066);
nand U5768 (N_5768,In_3489,In_3088);
or U5769 (N_5769,In_1137,In_4013);
nand U5770 (N_5770,In_1674,In_1178);
or U5771 (N_5771,In_3295,In_848);
nor U5772 (N_5772,In_1160,In_1005);
nand U5773 (N_5773,In_4548,In_4198);
and U5774 (N_5774,In_2016,In_722);
xor U5775 (N_5775,In_2516,In_3112);
or U5776 (N_5776,In_1422,In_2319);
nor U5777 (N_5777,In_4336,In_234);
nor U5778 (N_5778,In_1017,In_1009);
nand U5779 (N_5779,In_1646,In_4993);
or U5780 (N_5780,In_2572,In_2612);
and U5781 (N_5781,In_4565,In_4999);
nand U5782 (N_5782,In_2886,In_1207);
nor U5783 (N_5783,In_1315,In_906);
xor U5784 (N_5784,In_3363,In_1525);
nor U5785 (N_5785,In_4902,In_587);
nor U5786 (N_5786,In_3188,In_2879);
or U5787 (N_5787,In_4375,In_1625);
nor U5788 (N_5788,In_2160,In_2678);
and U5789 (N_5789,In_869,In_2604);
nor U5790 (N_5790,In_1882,In_891);
or U5791 (N_5791,In_4085,In_2192);
nor U5792 (N_5792,In_3981,In_1539);
xor U5793 (N_5793,In_3743,In_3662);
nor U5794 (N_5794,In_2584,In_4908);
or U5795 (N_5795,In_1454,In_4232);
nor U5796 (N_5796,In_335,In_2501);
nand U5797 (N_5797,In_3464,In_726);
or U5798 (N_5798,In_232,In_656);
nand U5799 (N_5799,In_551,In_2628);
nand U5800 (N_5800,In_19,In_4700);
nand U5801 (N_5801,In_2249,In_2509);
and U5802 (N_5802,In_615,In_3072);
xnor U5803 (N_5803,In_1574,In_2644);
or U5804 (N_5804,In_1725,In_2189);
nand U5805 (N_5805,In_2142,In_964);
xor U5806 (N_5806,In_416,In_4051);
xor U5807 (N_5807,In_2430,In_915);
nor U5808 (N_5808,In_3771,In_2797);
nor U5809 (N_5809,In_2440,In_3642);
and U5810 (N_5810,In_2574,In_522);
and U5811 (N_5811,In_2297,In_271);
and U5812 (N_5812,In_1192,In_3896);
nor U5813 (N_5813,In_3890,In_1091);
or U5814 (N_5814,In_3551,In_1627);
nor U5815 (N_5815,In_2247,In_1304);
and U5816 (N_5816,In_1311,In_154);
nand U5817 (N_5817,In_2941,In_708);
or U5818 (N_5818,In_851,In_2705);
xor U5819 (N_5819,In_3188,In_1887);
nor U5820 (N_5820,In_2877,In_1998);
nand U5821 (N_5821,In_2517,In_3082);
nand U5822 (N_5822,In_4515,In_4682);
and U5823 (N_5823,In_4066,In_2884);
nand U5824 (N_5824,In_4156,In_3254);
nor U5825 (N_5825,In_2045,In_1120);
and U5826 (N_5826,In_2063,In_1991);
or U5827 (N_5827,In_4044,In_4213);
nor U5828 (N_5828,In_1407,In_1383);
or U5829 (N_5829,In_4021,In_3883);
and U5830 (N_5830,In_4064,In_851);
nor U5831 (N_5831,In_4876,In_2811);
nand U5832 (N_5832,In_1997,In_3684);
and U5833 (N_5833,In_1049,In_3744);
nand U5834 (N_5834,In_3814,In_1013);
nor U5835 (N_5835,In_823,In_228);
nor U5836 (N_5836,In_4070,In_3411);
nand U5837 (N_5837,In_4632,In_1895);
and U5838 (N_5838,In_4724,In_4924);
nor U5839 (N_5839,In_298,In_2099);
or U5840 (N_5840,In_2383,In_2614);
nand U5841 (N_5841,In_4079,In_698);
or U5842 (N_5842,In_78,In_3667);
and U5843 (N_5843,In_2384,In_831);
or U5844 (N_5844,In_4127,In_1104);
nor U5845 (N_5845,In_3511,In_1160);
and U5846 (N_5846,In_1100,In_3346);
and U5847 (N_5847,In_3246,In_2376);
nand U5848 (N_5848,In_370,In_4882);
nor U5849 (N_5849,In_4621,In_4682);
nand U5850 (N_5850,In_2419,In_3003);
xor U5851 (N_5851,In_2251,In_2896);
and U5852 (N_5852,In_1230,In_1151);
xor U5853 (N_5853,In_1924,In_4442);
or U5854 (N_5854,In_1016,In_1150);
nand U5855 (N_5855,In_2660,In_265);
nand U5856 (N_5856,In_4498,In_3874);
nor U5857 (N_5857,In_2713,In_1336);
nor U5858 (N_5858,In_1204,In_887);
nand U5859 (N_5859,In_2548,In_2435);
or U5860 (N_5860,In_2800,In_1021);
and U5861 (N_5861,In_3603,In_3576);
or U5862 (N_5862,In_3050,In_300);
nor U5863 (N_5863,In_3970,In_3126);
xor U5864 (N_5864,In_3631,In_680);
nor U5865 (N_5865,In_4069,In_1046);
nor U5866 (N_5866,In_3521,In_3692);
nor U5867 (N_5867,In_2736,In_2231);
nand U5868 (N_5868,In_4283,In_2721);
xor U5869 (N_5869,In_4523,In_4009);
nor U5870 (N_5870,In_911,In_3113);
and U5871 (N_5871,In_1594,In_4108);
and U5872 (N_5872,In_2335,In_1547);
nor U5873 (N_5873,In_2605,In_4893);
nor U5874 (N_5874,In_1468,In_4219);
and U5875 (N_5875,In_2708,In_466);
and U5876 (N_5876,In_1901,In_2767);
or U5877 (N_5877,In_1186,In_1071);
xor U5878 (N_5878,In_4115,In_3375);
and U5879 (N_5879,In_2356,In_3528);
nand U5880 (N_5880,In_4448,In_4880);
nand U5881 (N_5881,In_1214,In_1510);
xor U5882 (N_5882,In_2926,In_3452);
and U5883 (N_5883,In_188,In_4472);
or U5884 (N_5884,In_4886,In_972);
nor U5885 (N_5885,In_4175,In_2712);
or U5886 (N_5886,In_855,In_570);
nand U5887 (N_5887,In_3224,In_1472);
nand U5888 (N_5888,In_3507,In_2613);
nor U5889 (N_5889,In_3608,In_2756);
nand U5890 (N_5890,In_2677,In_1347);
nor U5891 (N_5891,In_87,In_1994);
xor U5892 (N_5892,In_3921,In_4395);
or U5893 (N_5893,In_3780,In_2848);
nor U5894 (N_5894,In_3152,In_882);
or U5895 (N_5895,In_1332,In_4849);
nand U5896 (N_5896,In_3449,In_2175);
and U5897 (N_5897,In_2931,In_4137);
and U5898 (N_5898,In_3356,In_3939);
and U5899 (N_5899,In_4901,In_1456);
or U5900 (N_5900,In_2393,In_364);
xor U5901 (N_5901,In_2057,In_3862);
and U5902 (N_5902,In_178,In_2377);
and U5903 (N_5903,In_62,In_4534);
nor U5904 (N_5904,In_303,In_1695);
and U5905 (N_5905,In_1554,In_3079);
nor U5906 (N_5906,In_2731,In_1852);
or U5907 (N_5907,In_279,In_1014);
and U5908 (N_5908,In_304,In_1655);
and U5909 (N_5909,In_857,In_4273);
nor U5910 (N_5910,In_3207,In_1121);
nand U5911 (N_5911,In_3375,In_2074);
nor U5912 (N_5912,In_115,In_4779);
nand U5913 (N_5913,In_1824,In_881);
or U5914 (N_5914,In_2150,In_3637);
nor U5915 (N_5915,In_2201,In_3362);
xor U5916 (N_5916,In_2001,In_4693);
nor U5917 (N_5917,In_3968,In_331);
nand U5918 (N_5918,In_3167,In_609);
or U5919 (N_5919,In_2136,In_3569);
and U5920 (N_5920,In_3664,In_2194);
or U5921 (N_5921,In_165,In_327);
and U5922 (N_5922,In_2965,In_4385);
nor U5923 (N_5923,In_17,In_3621);
nand U5924 (N_5924,In_2557,In_2572);
or U5925 (N_5925,In_4211,In_290);
nand U5926 (N_5926,In_4981,In_672);
nor U5927 (N_5927,In_2355,In_5);
xor U5928 (N_5928,In_3739,In_2865);
and U5929 (N_5929,In_2267,In_4449);
or U5930 (N_5930,In_2859,In_1339);
or U5931 (N_5931,In_784,In_3149);
xor U5932 (N_5932,In_4948,In_4821);
nand U5933 (N_5933,In_4562,In_2664);
or U5934 (N_5934,In_2763,In_4024);
and U5935 (N_5935,In_1443,In_3523);
nand U5936 (N_5936,In_195,In_4740);
or U5937 (N_5937,In_4157,In_1984);
or U5938 (N_5938,In_2546,In_220);
xor U5939 (N_5939,In_642,In_1798);
and U5940 (N_5940,In_2998,In_2739);
nor U5941 (N_5941,In_1280,In_2246);
nand U5942 (N_5942,In_2595,In_3243);
nand U5943 (N_5943,In_1775,In_763);
and U5944 (N_5944,In_4073,In_3702);
xnor U5945 (N_5945,In_3930,In_2925);
or U5946 (N_5946,In_1071,In_2863);
nor U5947 (N_5947,In_1818,In_1539);
and U5948 (N_5948,In_3259,In_3069);
nand U5949 (N_5949,In_3971,In_2985);
nor U5950 (N_5950,In_4726,In_1564);
nand U5951 (N_5951,In_1169,In_1297);
nand U5952 (N_5952,In_997,In_1496);
nor U5953 (N_5953,In_2829,In_3812);
and U5954 (N_5954,In_3633,In_1557);
nand U5955 (N_5955,In_4276,In_2927);
nor U5956 (N_5956,In_338,In_2890);
and U5957 (N_5957,In_3311,In_427);
or U5958 (N_5958,In_94,In_1770);
and U5959 (N_5959,In_2038,In_3293);
and U5960 (N_5960,In_2779,In_1339);
nor U5961 (N_5961,In_1507,In_162);
or U5962 (N_5962,In_893,In_4781);
nand U5963 (N_5963,In_2309,In_664);
and U5964 (N_5964,In_2128,In_4625);
and U5965 (N_5965,In_218,In_3191);
or U5966 (N_5966,In_485,In_711);
nor U5967 (N_5967,In_4576,In_3575);
and U5968 (N_5968,In_3455,In_1136);
xor U5969 (N_5969,In_535,In_1794);
nor U5970 (N_5970,In_2094,In_2646);
or U5971 (N_5971,In_2,In_2534);
nand U5972 (N_5972,In_301,In_4871);
nor U5973 (N_5973,In_824,In_3785);
and U5974 (N_5974,In_4784,In_1560);
and U5975 (N_5975,In_2279,In_170);
nor U5976 (N_5976,In_414,In_3116);
and U5977 (N_5977,In_2803,In_2013);
or U5978 (N_5978,In_3699,In_438);
and U5979 (N_5979,In_3399,In_1219);
and U5980 (N_5980,In_1771,In_4753);
nor U5981 (N_5981,In_1713,In_787);
nor U5982 (N_5982,In_438,In_2606);
and U5983 (N_5983,In_2019,In_1961);
and U5984 (N_5984,In_4721,In_3516);
nand U5985 (N_5985,In_4729,In_3440);
and U5986 (N_5986,In_4895,In_2524);
or U5987 (N_5987,In_3357,In_484);
nand U5988 (N_5988,In_3871,In_2453);
xnor U5989 (N_5989,In_1608,In_4299);
nand U5990 (N_5990,In_636,In_1424);
and U5991 (N_5991,In_2603,In_3954);
nand U5992 (N_5992,In_704,In_4146);
and U5993 (N_5993,In_1042,In_2156);
nor U5994 (N_5994,In_839,In_2950);
and U5995 (N_5995,In_3582,In_1623);
nand U5996 (N_5996,In_2531,In_4056);
or U5997 (N_5997,In_3916,In_1258);
nand U5998 (N_5998,In_309,In_3561);
or U5999 (N_5999,In_4002,In_4663);
xnor U6000 (N_6000,In_78,In_3843);
xnor U6001 (N_6001,In_781,In_878);
nand U6002 (N_6002,In_2385,In_2283);
nand U6003 (N_6003,In_4038,In_3784);
nand U6004 (N_6004,In_2626,In_1250);
nor U6005 (N_6005,In_4421,In_4651);
nor U6006 (N_6006,In_4160,In_4998);
nand U6007 (N_6007,In_2917,In_1360);
or U6008 (N_6008,In_2448,In_1000);
nor U6009 (N_6009,In_4363,In_2528);
or U6010 (N_6010,In_788,In_1707);
nor U6011 (N_6011,In_2778,In_1108);
or U6012 (N_6012,In_3410,In_4030);
and U6013 (N_6013,In_588,In_3088);
nand U6014 (N_6014,In_707,In_79);
nor U6015 (N_6015,In_4827,In_3609);
nand U6016 (N_6016,In_3988,In_4908);
or U6017 (N_6017,In_4509,In_550);
or U6018 (N_6018,In_3541,In_1887);
nor U6019 (N_6019,In_4630,In_4479);
or U6020 (N_6020,In_4184,In_2492);
nand U6021 (N_6021,In_3225,In_1690);
nor U6022 (N_6022,In_4247,In_3053);
xor U6023 (N_6023,In_1379,In_751);
nand U6024 (N_6024,In_3586,In_2034);
or U6025 (N_6025,In_2483,In_3415);
and U6026 (N_6026,In_4991,In_3087);
xnor U6027 (N_6027,In_4001,In_3237);
nor U6028 (N_6028,In_1507,In_140);
and U6029 (N_6029,In_3752,In_3176);
nor U6030 (N_6030,In_1075,In_4089);
xnor U6031 (N_6031,In_2518,In_2397);
nand U6032 (N_6032,In_2576,In_819);
nor U6033 (N_6033,In_1105,In_2757);
nor U6034 (N_6034,In_3136,In_94);
and U6035 (N_6035,In_4202,In_3973);
and U6036 (N_6036,In_312,In_1780);
nor U6037 (N_6037,In_713,In_2105);
nor U6038 (N_6038,In_1400,In_887);
nor U6039 (N_6039,In_2139,In_4017);
nand U6040 (N_6040,In_1084,In_2308);
and U6041 (N_6041,In_4029,In_309);
nor U6042 (N_6042,In_1348,In_4074);
nor U6043 (N_6043,In_219,In_4970);
nor U6044 (N_6044,In_2976,In_1438);
xnor U6045 (N_6045,In_2567,In_2300);
xnor U6046 (N_6046,In_3876,In_1428);
xnor U6047 (N_6047,In_4040,In_3008);
or U6048 (N_6048,In_971,In_4439);
and U6049 (N_6049,In_1810,In_1177);
and U6050 (N_6050,In_536,In_1488);
nor U6051 (N_6051,In_1294,In_2104);
or U6052 (N_6052,In_857,In_2327);
or U6053 (N_6053,In_608,In_3918);
xor U6054 (N_6054,In_3066,In_2781);
or U6055 (N_6055,In_482,In_4165);
or U6056 (N_6056,In_3772,In_1090);
and U6057 (N_6057,In_68,In_909);
nand U6058 (N_6058,In_4685,In_1617);
nor U6059 (N_6059,In_4114,In_3184);
nor U6060 (N_6060,In_1651,In_1674);
or U6061 (N_6061,In_2984,In_2909);
xor U6062 (N_6062,In_1827,In_4661);
nand U6063 (N_6063,In_3302,In_221);
and U6064 (N_6064,In_4893,In_231);
nor U6065 (N_6065,In_961,In_3502);
nor U6066 (N_6066,In_4769,In_4023);
and U6067 (N_6067,In_2373,In_1584);
or U6068 (N_6068,In_3081,In_1256);
nand U6069 (N_6069,In_1047,In_107);
and U6070 (N_6070,In_4546,In_2567);
or U6071 (N_6071,In_2682,In_58);
xor U6072 (N_6072,In_3266,In_4625);
or U6073 (N_6073,In_2660,In_2495);
xnor U6074 (N_6074,In_2758,In_1611);
nor U6075 (N_6075,In_2624,In_2927);
nand U6076 (N_6076,In_2458,In_3782);
and U6077 (N_6077,In_4609,In_123);
nor U6078 (N_6078,In_1214,In_4991);
nand U6079 (N_6079,In_2534,In_34);
or U6080 (N_6080,In_4136,In_229);
nand U6081 (N_6081,In_4930,In_650);
and U6082 (N_6082,In_1350,In_1344);
nor U6083 (N_6083,In_1308,In_4674);
nand U6084 (N_6084,In_4414,In_591);
nor U6085 (N_6085,In_4446,In_1134);
or U6086 (N_6086,In_84,In_3382);
nor U6087 (N_6087,In_950,In_2220);
xnor U6088 (N_6088,In_2313,In_4087);
and U6089 (N_6089,In_4463,In_2501);
nand U6090 (N_6090,In_3307,In_1816);
and U6091 (N_6091,In_412,In_3524);
xnor U6092 (N_6092,In_3325,In_2806);
and U6093 (N_6093,In_3485,In_3184);
nor U6094 (N_6094,In_2811,In_4359);
and U6095 (N_6095,In_3583,In_3103);
xor U6096 (N_6096,In_3109,In_2123);
nor U6097 (N_6097,In_628,In_4609);
or U6098 (N_6098,In_4364,In_2190);
and U6099 (N_6099,In_223,In_1990);
or U6100 (N_6100,In_3491,In_560);
and U6101 (N_6101,In_4464,In_2538);
and U6102 (N_6102,In_4032,In_4154);
and U6103 (N_6103,In_2629,In_4524);
and U6104 (N_6104,In_370,In_2635);
and U6105 (N_6105,In_4352,In_1124);
or U6106 (N_6106,In_1499,In_4464);
and U6107 (N_6107,In_1098,In_2140);
and U6108 (N_6108,In_4826,In_4309);
and U6109 (N_6109,In_4348,In_1799);
and U6110 (N_6110,In_3194,In_1205);
or U6111 (N_6111,In_4012,In_911);
and U6112 (N_6112,In_2353,In_520);
or U6113 (N_6113,In_859,In_2083);
xnor U6114 (N_6114,In_2392,In_781);
and U6115 (N_6115,In_4329,In_4729);
nor U6116 (N_6116,In_3985,In_2110);
or U6117 (N_6117,In_24,In_97);
nand U6118 (N_6118,In_4476,In_1982);
or U6119 (N_6119,In_3009,In_1656);
or U6120 (N_6120,In_786,In_2146);
nor U6121 (N_6121,In_746,In_265);
nor U6122 (N_6122,In_858,In_394);
or U6123 (N_6123,In_3334,In_2778);
xor U6124 (N_6124,In_1576,In_3911);
or U6125 (N_6125,In_3186,In_1444);
nor U6126 (N_6126,In_2201,In_3332);
and U6127 (N_6127,In_3464,In_1498);
and U6128 (N_6128,In_549,In_4323);
nor U6129 (N_6129,In_1373,In_2648);
nand U6130 (N_6130,In_2439,In_753);
and U6131 (N_6131,In_2117,In_624);
nand U6132 (N_6132,In_3212,In_1388);
and U6133 (N_6133,In_1543,In_454);
and U6134 (N_6134,In_9,In_1567);
or U6135 (N_6135,In_1594,In_4073);
or U6136 (N_6136,In_2949,In_2456);
or U6137 (N_6137,In_2253,In_3471);
nor U6138 (N_6138,In_1015,In_4862);
and U6139 (N_6139,In_4889,In_554);
xnor U6140 (N_6140,In_2884,In_305);
xnor U6141 (N_6141,In_3648,In_2450);
nor U6142 (N_6142,In_488,In_3646);
or U6143 (N_6143,In_125,In_3209);
nand U6144 (N_6144,In_3329,In_418);
nand U6145 (N_6145,In_4418,In_2902);
xnor U6146 (N_6146,In_4351,In_576);
nand U6147 (N_6147,In_1060,In_4787);
nand U6148 (N_6148,In_4200,In_731);
and U6149 (N_6149,In_3853,In_4306);
and U6150 (N_6150,In_318,In_4354);
or U6151 (N_6151,In_1487,In_1106);
or U6152 (N_6152,In_4425,In_1835);
or U6153 (N_6153,In_2721,In_1412);
or U6154 (N_6154,In_3423,In_3963);
or U6155 (N_6155,In_3993,In_4151);
xor U6156 (N_6156,In_3316,In_3803);
or U6157 (N_6157,In_2799,In_755);
and U6158 (N_6158,In_2099,In_3113);
and U6159 (N_6159,In_1564,In_3109);
nand U6160 (N_6160,In_4999,In_1179);
nor U6161 (N_6161,In_4540,In_4066);
nor U6162 (N_6162,In_434,In_410);
or U6163 (N_6163,In_1789,In_361);
nor U6164 (N_6164,In_4305,In_960);
nand U6165 (N_6165,In_4543,In_2930);
xor U6166 (N_6166,In_1497,In_4160);
nor U6167 (N_6167,In_3958,In_2995);
nand U6168 (N_6168,In_2966,In_4555);
xor U6169 (N_6169,In_563,In_825);
nand U6170 (N_6170,In_4046,In_2757);
nor U6171 (N_6171,In_4507,In_2530);
and U6172 (N_6172,In_4088,In_4119);
nor U6173 (N_6173,In_4228,In_4906);
nand U6174 (N_6174,In_4964,In_3280);
xor U6175 (N_6175,In_3041,In_536);
or U6176 (N_6176,In_2119,In_2660);
nand U6177 (N_6177,In_283,In_4058);
nand U6178 (N_6178,In_3535,In_4954);
or U6179 (N_6179,In_3257,In_3815);
nor U6180 (N_6180,In_4706,In_2345);
nor U6181 (N_6181,In_2159,In_1083);
nand U6182 (N_6182,In_346,In_1776);
or U6183 (N_6183,In_3165,In_4735);
nand U6184 (N_6184,In_1770,In_590);
or U6185 (N_6185,In_1548,In_378);
and U6186 (N_6186,In_4106,In_2560);
nor U6187 (N_6187,In_3532,In_1403);
nor U6188 (N_6188,In_74,In_213);
and U6189 (N_6189,In_1276,In_2500);
or U6190 (N_6190,In_1361,In_2960);
or U6191 (N_6191,In_4952,In_412);
nor U6192 (N_6192,In_4683,In_1490);
xnor U6193 (N_6193,In_1839,In_3631);
or U6194 (N_6194,In_1686,In_507);
nand U6195 (N_6195,In_3446,In_1110);
and U6196 (N_6196,In_4189,In_3425);
or U6197 (N_6197,In_3429,In_4039);
or U6198 (N_6198,In_455,In_3431);
or U6199 (N_6199,In_1815,In_1970);
nor U6200 (N_6200,In_2376,In_1077);
or U6201 (N_6201,In_3063,In_3655);
nor U6202 (N_6202,In_2075,In_272);
xor U6203 (N_6203,In_2091,In_1501);
xnor U6204 (N_6204,In_1715,In_3828);
nor U6205 (N_6205,In_2234,In_4725);
and U6206 (N_6206,In_367,In_2015);
nand U6207 (N_6207,In_981,In_701);
nor U6208 (N_6208,In_3402,In_3499);
xor U6209 (N_6209,In_758,In_1518);
and U6210 (N_6210,In_1253,In_608);
or U6211 (N_6211,In_4513,In_2754);
and U6212 (N_6212,In_2002,In_2222);
nand U6213 (N_6213,In_3123,In_4438);
nand U6214 (N_6214,In_2031,In_2077);
and U6215 (N_6215,In_2803,In_2360);
and U6216 (N_6216,In_3788,In_16);
and U6217 (N_6217,In_3804,In_1354);
nand U6218 (N_6218,In_922,In_4773);
nand U6219 (N_6219,In_1926,In_4790);
nand U6220 (N_6220,In_758,In_1068);
or U6221 (N_6221,In_2378,In_91);
or U6222 (N_6222,In_3565,In_3733);
nand U6223 (N_6223,In_3189,In_3378);
nor U6224 (N_6224,In_4665,In_603);
or U6225 (N_6225,In_2861,In_4710);
nand U6226 (N_6226,In_2064,In_748);
nor U6227 (N_6227,In_329,In_1985);
nand U6228 (N_6228,In_234,In_3828);
nor U6229 (N_6229,In_1512,In_2147);
or U6230 (N_6230,In_2320,In_411);
and U6231 (N_6231,In_174,In_2489);
or U6232 (N_6232,In_117,In_2266);
nand U6233 (N_6233,In_2739,In_3900);
nor U6234 (N_6234,In_841,In_1143);
nand U6235 (N_6235,In_4438,In_3621);
nand U6236 (N_6236,In_3957,In_3785);
nand U6237 (N_6237,In_2301,In_960);
and U6238 (N_6238,In_1005,In_4304);
or U6239 (N_6239,In_1229,In_3297);
nor U6240 (N_6240,In_2806,In_408);
nor U6241 (N_6241,In_1481,In_2152);
or U6242 (N_6242,In_3538,In_3150);
or U6243 (N_6243,In_3041,In_4267);
and U6244 (N_6244,In_4907,In_736);
nor U6245 (N_6245,In_3959,In_2340);
nand U6246 (N_6246,In_2878,In_3270);
and U6247 (N_6247,In_1462,In_2188);
nand U6248 (N_6248,In_2565,In_4292);
xnor U6249 (N_6249,In_2144,In_2481);
nand U6250 (N_6250,In_754,In_4648);
nor U6251 (N_6251,In_2100,In_1436);
xor U6252 (N_6252,In_2033,In_1874);
nand U6253 (N_6253,In_2827,In_1253);
xor U6254 (N_6254,In_3114,In_255);
nand U6255 (N_6255,In_2032,In_4474);
nand U6256 (N_6256,In_62,In_3417);
nand U6257 (N_6257,In_135,In_1949);
and U6258 (N_6258,In_3172,In_3537);
nand U6259 (N_6259,In_164,In_2105);
nand U6260 (N_6260,In_2264,In_2430);
and U6261 (N_6261,In_4595,In_3065);
and U6262 (N_6262,In_4685,In_1053);
nor U6263 (N_6263,In_1146,In_3539);
nand U6264 (N_6264,In_1953,In_2327);
and U6265 (N_6265,In_3708,In_588);
xnor U6266 (N_6266,In_4601,In_3932);
or U6267 (N_6267,In_2286,In_4679);
and U6268 (N_6268,In_445,In_1655);
or U6269 (N_6269,In_1114,In_3441);
xnor U6270 (N_6270,In_2890,In_1580);
or U6271 (N_6271,In_1240,In_2439);
nand U6272 (N_6272,In_3498,In_726);
xor U6273 (N_6273,In_4802,In_1974);
nor U6274 (N_6274,In_4783,In_3224);
or U6275 (N_6275,In_2818,In_2680);
nand U6276 (N_6276,In_3077,In_2213);
or U6277 (N_6277,In_184,In_4137);
nor U6278 (N_6278,In_3752,In_2522);
xnor U6279 (N_6279,In_3705,In_4970);
nor U6280 (N_6280,In_4727,In_2050);
nor U6281 (N_6281,In_4047,In_296);
or U6282 (N_6282,In_952,In_2221);
or U6283 (N_6283,In_4945,In_1345);
nor U6284 (N_6284,In_1364,In_2940);
or U6285 (N_6285,In_2262,In_4237);
nand U6286 (N_6286,In_352,In_4267);
nor U6287 (N_6287,In_2950,In_870);
and U6288 (N_6288,In_2542,In_2397);
and U6289 (N_6289,In_1296,In_3479);
xnor U6290 (N_6290,In_3100,In_963);
or U6291 (N_6291,In_3794,In_1840);
xnor U6292 (N_6292,In_1958,In_233);
or U6293 (N_6293,In_2589,In_4700);
nand U6294 (N_6294,In_382,In_4163);
or U6295 (N_6295,In_682,In_2065);
xnor U6296 (N_6296,In_1780,In_659);
and U6297 (N_6297,In_1048,In_2007);
or U6298 (N_6298,In_817,In_4178);
or U6299 (N_6299,In_2653,In_3808);
or U6300 (N_6300,In_1934,In_4354);
nor U6301 (N_6301,In_3321,In_2308);
nand U6302 (N_6302,In_3743,In_3582);
nand U6303 (N_6303,In_4519,In_856);
nand U6304 (N_6304,In_2764,In_902);
nor U6305 (N_6305,In_4730,In_3186);
nor U6306 (N_6306,In_3689,In_3095);
or U6307 (N_6307,In_3337,In_2257);
or U6308 (N_6308,In_98,In_3096);
nand U6309 (N_6309,In_2676,In_4284);
xnor U6310 (N_6310,In_4674,In_1833);
nor U6311 (N_6311,In_3930,In_1807);
and U6312 (N_6312,In_2423,In_3859);
and U6313 (N_6313,In_213,In_1731);
or U6314 (N_6314,In_1557,In_3883);
and U6315 (N_6315,In_3893,In_2049);
and U6316 (N_6316,In_1426,In_4349);
or U6317 (N_6317,In_1041,In_561);
and U6318 (N_6318,In_1634,In_3743);
and U6319 (N_6319,In_1900,In_204);
nand U6320 (N_6320,In_1692,In_1988);
nand U6321 (N_6321,In_3809,In_1255);
xor U6322 (N_6322,In_2,In_715);
nand U6323 (N_6323,In_3169,In_575);
and U6324 (N_6324,In_3566,In_236);
or U6325 (N_6325,In_3037,In_456);
and U6326 (N_6326,In_131,In_787);
and U6327 (N_6327,In_4180,In_2467);
and U6328 (N_6328,In_877,In_229);
and U6329 (N_6329,In_1888,In_4589);
or U6330 (N_6330,In_1507,In_2004);
nand U6331 (N_6331,In_880,In_1663);
nand U6332 (N_6332,In_167,In_4692);
nand U6333 (N_6333,In_110,In_545);
nor U6334 (N_6334,In_2784,In_51);
nor U6335 (N_6335,In_739,In_205);
or U6336 (N_6336,In_2004,In_3144);
and U6337 (N_6337,In_3329,In_170);
nand U6338 (N_6338,In_2106,In_4116);
nor U6339 (N_6339,In_3222,In_4924);
nand U6340 (N_6340,In_1314,In_3485);
or U6341 (N_6341,In_1677,In_3084);
nor U6342 (N_6342,In_193,In_2033);
or U6343 (N_6343,In_3704,In_329);
nand U6344 (N_6344,In_46,In_3357);
or U6345 (N_6345,In_2081,In_4797);
or U6346 (N_6346,In_3002,In_2311);
xnor U6347 (N_6347,In_1373,In_1401);
or U6348 (N_6348,In_4690,In_950);
xor U6349 (N_6349,In_740,In_2576);
and U6350 (N_6350,In_3270,In_4419);
nor U6351 (N_6351,In_3284,In_2860);
nor U6352 (N_6352,In_678,In_2917);
xor U6353 (N_6353,In_4594,In_730);
xnor U6354 (N_6354,In_1286,In_627);
and U6355 (N_6355,In_4123,In_4919);
and U6356 (N_6356,In_943,In_3794);
or U6357 (N_6357,In_1762,In_1831);
nor U6358 (N_6358,In_2071,In_2698);
or U6359 (N_6359,In_4507,In_337);
nor U6360 (N_6360,In_1874,In_4454);
and U6361 (N_6361,In_2523,In_2426);
and U6362 (N_6362,In_4106,In_4227);
and U6363 (N_6363,In_914,In_3077);
nand U6364 (N_6364,In_2951,In_3228);
nor U6365 (N_6365,In_1386,In_2734);
nor U6366 (N_6366,In_2125,In_366);
nor U6367 (N_6367,In_3280,In_749);
nor U6368 (N_6368,In_1509,In_1789);
and U6369 (N_6369,In_4060,In_3961);
nor U6370 (N_6370,In_861,In_2022);
and U6371 (N_6371,In_3772,In_833);
nand U6372 (N_6372,In_705,In_1667);
nand U6373 (N_6373,In_1524,In_900);
nand U6374 (N_6374,In_3086,In_4468);
or U6375 (N_6375,In_1164,In_1384);
nor U6376 (N_6376,In_3349,In_4405);
nor U6377 (N_6377,In_2439,In_4828);
nand U6378 (N_6378,In_386,In_1015);
nor U6379 (N_6379,In_2031,In_3468);
and U6380 (N_6380,In_2513,In_1239);
and U6381 (N_6381,In_3124,In_3021);
or U6382 (N_6382,In_856,In_3579);
xor U6383 (N_6383,In_1420,In_1974);
and U6384 (N_6384,In_1519,In_831);
nand U6385 (N_6385,In_4883,In_4171);
xor U6386 (N_6386,In_168,In_2333);
or U6387 (N_6387,In_3478,In_938);
xnor U6388 (N_6388,In_402,In_668);
and U6389 (N_6389,In_2976,In_11);
nand U6390 (N_6390,In_4974,In_3346);
nor U6391 (N_6391,In_4951,In_2865);
nand U6392 (N_6392,In_4776,In_2978);
or U6393 (N_6393,In_3118,In_4555);
nor U6394 (N_6394,In_4254,In_1714);
or U6395 (N_6395,In_1712,In_3173);
and U6396 (N_6396,In_1459,In_1010);
xnor U6397 (N_6397,In_1147,In_2564);
or U6398 (N_6398,In_1428,In_4044);
and U6399 (N_6399,In_1044,In_3337);
nor U6400 (N_6400,In_2161,In_3818);
and U6401 (N_6401,In_4128,In_3517);
or U6402 (N_6402,In_3275,In_2019);
nand U6403 (N_6403,In_406,In_4876);
or U6404 (N_6404,In_4341,In_1121);
nand U6405 (N_6405,In_2093,In_3724);
or U6406 (N_6406,In_4242,In_2780);
nor U6407 (N_6407,In_1500,In_3015);
or U6408 (N_6408,In_169,In_338);
or U6409 (N_6409,In_1410,In_766);
nor U6410 (N_6410,In_2136,In_2418);
or U6411 (N_6411,In_1257,In_293);
or U6412 (N_6412,In_3003,In_1120);
or U6413 (N_6413,In_1705,In_653);
nor U6414 (N_6414,In_4248,In_4637);
nor U6415 (N_6415,In_2205,In_1361);
and U6416 (N_6416,In_1878,In_998);
nor U6417 (N_6417,In_2951,In_4896);
xor U6418 (N_6418,In_3839,In_4979);
and U6419 (N_6419,In_153,In_4874);
xor U6420 (N_6420,In_4280,In_3825);
and U6421 (N_6421,In_4844,In_2405);
or U6422 (N_6422,In_3692,In_2631);
nor U6423 (N_6423,In_4404,In_38);
or U6424 (N_6424,In_4620,In_3791);
nor U6425 (N_6425,In_3584,In_4780);
and U6426 (N_6426,In_141,In_3924);
nand U6427 (N_6427,In_292,In_2375);
or U6428 (N_6428,In_1694,In_651);
nor U6429 (N_6429,In_1400,In_458);
nor U6430 (N_6430,In_2783,In_1952);
nor U6431 (N_6431,In_761,In_4917);
nand U6432 (N_6432,In_206,In_1792);
or U6433 (N_6433,In_645,In_2797);
nand U6434 (N_6434,In_3627,In_943);
nor U6435 (N_6435,In_3868,In_1539);
nand U6436 (N_6436,In_4870,In_396);
and U6437 (N_6437,In_3481,In_1820);
nor U6438 (N_6438,In_4920,In_1868);
or U6439 (N_6439,In_2697,In_4412);
and U6440 (N_6440,In_2625,In_987);
and U6441 (N_6441,In_3994,In_2955);
nor U6442 (N_6442,In_895,In_2565);
and U6443 (N_6443,In_388,In_3852);
nor U6444 (N_6444,In_1894,In_539);
nand U6445 (N_6445,In_3024,In_4001);
nor U6446 (N_6446,In_1689,In_4659);
and U6447 (N_6447,In_636,In_3735);
nand U6448 (N_6448,In_4817,In_4644);
and U6449 (N_6449,In_4514,In_2999);
or U6450 (N_6450,In_2824,In_1188);
and U6451 (N_6451,In_2812,In_1692);
nor U6452 (N_6452,In_4979,In_2357);
nand U6453 (N_6453,In_3414,In_1604);
xnor U6454 (N_6454,In_4158,In_807);
or U6455 (N_6455,In_4199,In_1897);
nor U6456 (N_6456,In_3177,In_2822);
nor U6457 (N_6457,In_2597,In_2681);
or U6458 (N_6458,In_2400,In_20);
nand U6459 (N_6459,In_2175,In_4100);
nor U6460 (N_6460,In_2120,In_2600);
nand U6461 (N_6461,In_3741,In_3947);
or U6462 (N_6462,In_1858,In_2451);
and U6463 (N_6463,In_206,In_3254);
or U6464 (N_6464,In_1765,In_1520);
nand U6465 (N_6465,In_1692,In_3557);
and U6466 (N_6466,In_2273,In_2714);
xnor U6467 (N_6467,In_1375,In_701);
and U6468 (N_6468,In_3241,In_2923);
xor U6469 (N_6469,In_1855,In_3145);
and U6470 (N_6470,In_2740,In_902);
or U6471 (N_6471,In_3710,In_40);
nor U6472 (N_6472,In_134,In_1928);
nor U6473 (N_6473,In_4553,In_3298);
nor U6474 (N_6474,In_748,In_1117);
nand U6475 (N_6475,In_2935,In_2635);
or U6476 (N_6476,In_4120,In_3652);
and U6477 (N_6477,In_4373,In_288);
or U6478 (N_6478,In_993,In_684);
and U6479 (N_6479,In_2991,In_1999);
nor U6480 (N_6480,In_251,In_3902);
or U6481 (N_6481,In_396,In_1927);
or U6482 (N_6482,In_2653,In_1288);
nand U6483 (N_6483,In_1567,In_177);
or U6484 (N_6484,In_4513,In_2686);
nand U6485 (N_6485,In_2954,In_981);
nand U6486 (N_6486,In_4223,In_1618);
nor U6487 (N_6487,In_442,In_2894);
nor U6488 (N_6488,In_4967,In_1278);
nor U6489 (N_6489,In_577,In_3831);
nor U6490 (N_6490,In_1160,In_1492);
xor U6491 (N_6491,In_3901,In_2612);
nand U6492 (N_6492,In_1547,In_4681);
nor U6493 (N_6493,In_902,In_3291);
nor U6494 (N_6494,In_2960,In_2197);
nand U6495 (N_6495,In_1209,In_4739);
xnor U6496 (N_6496,In_81,In_3414);
nor U6497 (N_6497,In_4739,In_4667);
nor U6498 (N_6498,In_1930,In_313);
nor U6499 (N_6499,In_1376,In_405);
and U6500 (N_6500,In_4122,In_2796);
nand U6501 (N_6501,In_3340,In_2241);
nand U6502 (N_6502,In_1595,In_2698);
or U6503 (N_6503,In_829,In_584);
nand U6504 (N_6504,In_4146,In_824);
nand U6505 (N_6505,In_1953,In_3901);
xor U6506 (N_6506,In_4888,In_253);
and U6507 (N_6507,In_1482,In_4162);
nand U6508 (N_6508,In_1065,In_2325);
xnor U6509 (N_6509,In_2646,In_314);
or U6510 (N_6510,In_4220,In_4388);
nor U6511 (N_6511,In_1526,In_1576);
nand U6512 (N_6512,In_3944,In_1345);
nand U6513 (N_6513,In_2901,In_4213);
nand U6514 (N_6514,In_136,In_1868);
xor U6515 (N_6515,In_2903,In_630);
nand U6516 (N_6516,In_2030,In_3745);
nand U6517 (N_6517,In_4739,In_565);
and U6518 (N_6518,In_4358,In_3578);
or U6519 (N_6519,In_4551,In_2264);
nor U6520 (N_6520,In_4622,In_1240);
and U6521 (N_6521,In_3795,In_3801);
or U6522 (N_6522,In_3674,In_1953);
nor U6523 (N_6523,In_4241,In_1927);
nand U6524 (N_6524,In_3450,In_3070);
or U6525 (N_6525,In_3989,In_1047);
or U6526 (N_6526,In_4931,In_1734);
xnor U6527 (N_6527,In_4130,In_2925);
xor U6528 (N_6528,In_1433,In_2466);
and U6529 (N_6529,In_1443,In_3775);
and U6530 (N_6530,In_2280,In_4974);
nor U6531 (N_6531,In_4169,In_3577);
nand U6532 (N_6532,In_4230,In_1530);
or U6533 (N_6533,In_4813,In_4989);
nor U6534 (N_6534,In_886,In_1584);
nor U6535 (N_6535,In_505,In_103);
nand U6536 (N_6536,In_3779,In_4056);
and U6537 (N_6537,In_2928,In_3827);
and U6538 (N_6538,In_3322,In_4926);
and U6539 (N_6539,In_421,In_2424);
nand U6540 (N_6540,In_879,In_2333);
nor U6541 (N_6541,In_4464,In_2246);
or U6542 (N_6542,In_3439,In_4995);
or U6543 (N_6543,In_1212,In_3997);
and U6544 (N_6544,In_3202,In_33);
xnor U6545 (N_6545,In_3915,In_1634);
xnor U6546 (N_6546,In_3314,In_3618);
nor U6547 (N_6547,In_4572,In_1504);
or U6548 (N_6548,In_3014,In_1150);
and U6549 (N_6549,In_3488,In_2545);
nor U6550 (N_6550,In_4561,In_3333);
and U6551 (N_6551,In_1912,In_3473);
or U6552 (N_6552,In_3835,In_1694);
and U6553 (N_6553,In_858,In_4020);
or U6554 (N_6554,In_2458,In_2108);
or U6555 (N_6555,In_998,In_2766);
and U6556 (N_6556,In_1622,In_4903);
nor U6557 (N_6557,In_1206,In_1350);
and U6558 (N_6558,In_4482,In_4637);
nand U6559 (N_6559,In_2355,In_3029);
and U6560 (N_6560,In_4668,In_1939);
and U6561 (N_6561,In_2650,In_631);
or U6562 (N_6562,In_3159,In_4915);
nand U6563 (N_6563,In_2349,In_1248);
nand U6564 (N_6564,In_3094,In_2724);
or U6565 (N_6565,In_452,In_1360);
or U6566 (N_6566,In_1622,In_3037);
nand U6567 (N_6567,In_2107,In_3749);
nand U6568 (N_6568,In_3224,In_1269);
or U6569 (N_6569,In_1291,In_3990);
nand U6570 (N_6570,In_381,In_3890);
and U6571 (N_6571,In_1386,In_2237);
nand U6572 (N_6572,In_2920,In_1204);
xor U6573 (N_6573,In_2601,In_897);
nor U6574 (N_6574,In_3027,In_714);
or U6575 (N_6575,In_813,In_196);
nand U6576 (N_6576,In_2443,In_2619);
nand U6577 (N_6577,In_983,In_562);
nand U6578 (N_6578,In_4848,In_3885);
and U6579 (N_6579,In_2862,In_3283);
nand U6580 (N_6580,In_2354,In_1917);
xnor U6581 (N_6581,In_1067,In_2886);
or U6582 (N_6582,In_3404,In_4536);
and U6583 (N_6583,In_4371,In_2518);
nor U6584 (N_6584,In_200,In_2958);
nand U6585 (N_6585,In_2839,In_2622);
nand U6586 (N_6586,In_2187,In_20);
xor U6587 (N_6587,In_4037,In_1342);
xor U6588 (N_6588,In_3558,In_2768);
and U6589 (N_6589,In_3034,In_1028);
or U6590 (N_6590,In_3179,In_4070);
and U6591 (N_6591,In_2212,In_4624);
or U6592 (N_6592,In_2910,In_4316);
nor U6593 (N_6593,In_1008,In_2924);
and U6594 (N_6594,In_717,In_4349);
nand U6595 (N_6595,In_3144,In_2767);
xnor U6596 (N_6596,In_4472,In_2074);
or U6597 (N_6597,In_1485,In_3008);
and U6598 (N_6598,In_3981,In_371);
nand U6599 (N_6599,In_1063,In_4251);
and U6600 (N_6600,In_4074,In_3317);
nand U6601 (N_6601,In_138,In_146);
or U6602 (N_6602,In_2868,In_2929);
and U6603 (N_6603,In_454,In_2191);
nor U6604 (N_6604,In_722,In_730);
nor U6605 (N_6605,In_4515,In_4345);
or U6606 (N_6606,In_4045,In_3535);
or U6607 (N_6607,In_202,In_4705);
or U6608 (N_6608,In_3689,In_1831);
nand U6609 (N_6609,In_4564,In_4736);
nand U6610 (N_6610,In_1349,In_4343);
or U6611 (N_6611,In_1002,In_2017);
nor U6612 (N_6612,In_2457,In_2959);
xnor U6613 (N_6613,In_4834,In_4782);
xor U6614 (N_6614,In_1127,In_4888);
nor U6615 (N_6615,In_609,In_2026);
and U6616 (N_6616,In_4353,In_3452);
or U6617 (N_6617,In_3020,In_4372);
and U6618 (N_6618,In_4167,In_567);
nor U6619 (N_6619,In_2527,In_3084);
nor U6620 (N_6620,In_4507,In_566);
nor U6621 (N_6621,In_169,In_650);
and U6622 (N_6622,In_837,In_550);
or U6623 (N_6623,In_4346,In_144);
nor U6624 (N_6624,In_2993,In_3633);
nor U6625 (N_6625,In_284,In_2048);
nor U6626 (N_6626,In_4195,In_4292);
and U6627 (N_6627,In_4840,In_3882);
and U6628 (N_6628,In_3316,In_1943);
nand U6629 (N_6629,In_3869,In_3891);
nor U6630 (N_6630,In_2104,In_1208);
nor U6631 (N_6631,In_3944,In_2712);
or U6632 (N_6632,In_4798,In_178);
or U6633 (N_6633,In_2056,In_2477);
or U6634 (N_6634,In_956,In_4571);
xnor U6635 (N_6635,In_59,In_329);
or U6636 (N_6636,In_3978,In_4634);
or U6637 (N_6637,In_3427,In_2211);
and U6638 (N_6638,In_4942,In_2632);
nor U6639 (N_6639,In_3301,In_629);
nand U6640 (N_6640,In_3201,In_4878);
xnor U6641 (N_6641,In_3658,In_4497);
nand U6642 (N_6642,In_4100,In_1836);
nand U6643 (N_6643,In_2363,In_95);
or U6644 (N_6644,In_4791,In_2291);
or U6645 (N_6645,In_2556,In_4970);
nor U6646 (N_6646,In_3026,In_3257);
nand U6647 (N_6647,In_119,In_2413);
nor U6648 (N_6648,In_2669,In_2029);
and U6649 (N_6649,In_2748,In_1398);
or U6650 (N_6650,In_4652,In_4260);
xor U6651 (N_6651,In_945,In_4177);
or U6652 (N_6652,In_2116,In_1926);
nand U6653 (N_6653,In_2221,In_3028);
nand U6654 (N_6654,In_756,In_3212);
and U6655 (N_6655,In_3788,In_3910);
nor U6656 (N_6656,In_809,In_2142);
xnor U6657 (N_6657,In_1850,In_4818);
or U6658 (N_6658,In_463,In_4137);
or U6659 (N_6659,In_2625,In_4381);
nor U6660 (N_6660,In_938,In_1975);
or U6661 (N_6661,In_3981,In_3393);
and U6662 (N_6662,In_142,In_2775);
nor U6663 (N_6663,In_4910,In_4950);
nand U6664 (N_6664,In_1570,In_4047);
nor U6665 (N_6665,In_3613,In_3912);
xnor U6666 (N_6666,In_2133,In_2964);
nor U6667 (N_6667,In_585,In_2165);
or U6668 (N_6668,In_2362,In_2108);
and U6669 (N_6669,In_1237,In_972);
nand U6670 (N_6670,In_859,In_2972);
nand U6671 (N_6671,In_3254,In_3072);
or U6672 (N_6672,In_4401,In_2312);
or U6673 (N_6673,In_851,In_3531);
nor U6674 (N_6674,In_4227,In_1269);
nor U6675 (N_6675,In_4441,In_1836);
nand U6676 (N_6676,In_3377,In_3963);
nor U6677 (N_6677,In_217,In_2417);
nor U6678 (N_6678,In_4481,In_4160);
nand U6679 (N_6679,In_1677,In_1230);
nand U6680 (N_6680,In_3100,In_2629);
xor U6681 (N_6681,In_1974,In_30);
or U6682 (N_6682,In_920,In_4433);
nand U6683 (N_6683,In_106,In_2840);
nor U6684 (N_6684,In_3994,In_2612);
xor U6685 (N_6685,In_3121,In_567);
and U6686 (N_6686,In_2968,In_1484);
nand U6687 (N_6687,In_2094,In_2200);
nand U6688 (N_6688,In_2634,In_2985);
or U6689 (N_6689,In_3522,In_4387);
xnor U6690 (N_6690,In_1130,In_41);
and U6691 (N_6691,In_2488,In_2013);
or U6692 (N_6692,In_2012,In_3086);
xnor U6693 (N_6693,In_3034,In_2373);
or U6694 (N_6694,In_361,In_172);
nand U6695 (N_6695,In_838,In_1471);
or U6696 (N_6696,In_1470,In_2533);
and U6697 (N_6697,In_886,In_4734);
nor U6698 (N_6698,In_4899,In_829);
xnor U6699 (N_6699,In_1998,In_2160);
nor U6700 (N_6700,In_705,In_1588);
and U6701 (N_6701,In_2573,In_2388);
and U6702 (N_6702,In_3946,In_2825);
and U6703 (N_6703,In_2277,In_2104);
or U6704 (N_6704,In_559,In_2711);
nand U6705 (N_6705,In_3582,In_958);
or U6706 (N_6706,In_1041,In_3402);
and U6707 (N_6707,In_4532,In_1672);
and U6708 (N_6708,In_2918,In_4935);
and U6709 (N_6709,In_4841,In_1707);
nand U6710 (N_6710,In_3020,In_4224);
and U6711 (N_6711,In_660,In_945);
nand U6712 (N_6712,In_4570,In_2377);
nand U6713 (N_6713,In_1513,In_1349);
nor U6714 (N_6714,In_1608,In_4356);
nor U6715 (N_6715,In_3884,In_2047);
and U6716 (N_6716,In_3225,In_2286);
xor U6717 (N_6717,In_942,In_1444);
or U6718 (N_6718,In_1442,In_2132);
and U6719 (N_6719,In_1884,In_4863);
nor U6720 (N_6720,In_1024,In_2070);
nand U6721 (N_6721,In_2764,In_4608);
or U6722 (N_6722,In_1831,In_2879);
and U6723 (N_6723,In_1823,In_2131);
nor U6724 (N_6724,In_4919,In_2174);
or U6725 (N_6725,In_314,In_4487);
nand U6726 (N_6726,In_2288,In_4835);
xnor U6727 (N_6727,In_1871,In_1793);
or U6728 (N_6728,In_231,In_3052);
or U6729 (N_6729,In_1426,In_381);
nor U6730 (N_6730,In_1267,In_2100);
and U6731 (N_6731,In_1087,In_3354);
or U6732 (N_6732,In_273,In_643);
and U6733 (N_6733,In_1548,In_3553);
or U6734 (N_6734,In_1404,In_4952);
and U6735 (N_6735,In_4635,In_3354);
nand U6736 (N_6736,In_3266,In_2029);
nand U6737 (N_6737,In_1740,In_2990);
or U6738 (N_6738,In_4919,In_1821);
or U6739 (N_6739,In_1696,In_3384);
and U6740 (N_6740,In_3784,In_4241);
and U6741 (N_6741,In_1351,In_697);
nand U6742 (N_6742,In_3399,In_567);
or U6743 (N_6743,In_2262,In_574);
xnor U6744 (N_6744,In_4318,In_4540);
nor U6745 (N_6745,In_4354,In_856);
and U6746 (N_6746,In_774,In_4977);
and U6747 (N_6747,In_2682,In_1038);
nor U6748 (N_6748,In_969,In_61);
nor U6749 (N_6749,In_508,In_4871);
xor U6750 (N_6750,In_4998,In_1614);
xor U6751 (N_6751,In_419,In_266);
nand U6752 (N_6752,In_3878,In_2545);
nor U6753 (N_6753,In_3409,In_439);
xnor U6754 (N_6754,In_1812,In_4913);
nor U6755 (N_6755,In_3698,In_4045);
or U6756 (N_6756,In_2998,In_3934);
or U6757 (N_6757,In_4497,In_4316);
nand U6758 (N_6758,In_3250,In_1433);
nand U6759 (N_6759,In_1554,In_4176);
or U6760 (N_6760,In_124,In_2459);
nor U6761 (N_6761,In_4006,In_682);
or U6762 (N_6762,In_4421,In_502);
or U6763 (N_6763,In_3004,In_1046);
nor U6764 (N_6764,In_1038,In_1390);
and U6765 (N_6765,In_2098,In_3584);
and U6766 (N_6766,In_3654,In_529);
nand U6767 (N_6767,In_949,In_3104);
nor U6768 (N_6768,In_2921,In_3093);
or U6769 (N_6769,In_3631,In_353);
xnor U6770 (N_6770,In_4773,In_2078);
nor U6771 (N_6771,In_1923,In_1464);
nand U6772 (N_6772,In_3827,In_4908);
and U6773 (N_6773,In_4666,In_1332);
nand U6774 (N_6774,In_1744,In_950);
and U6775 (N_6775,In_706,In_982);
or U6776 (N_6776,In_1350,In_1128);
xor U6777 (N_6777,In_1383,In_2214);
nand U6778 (N_6778,In_4960,In_3942);
nor U6779 (N_6779,In_4572,In_1749);
nand U6780 (N_6780,In_4390,In_2505);
or U6781 (N_6781,In_4123,In_1137);
and U6782 (N_6782,In_2348,In_3807);
nor U6783 (N_6783,In_1473,In_1840);
nor U6784 (N_6784,In_3779,In_4035);
nor U6785 (N_6785,In_617,In_3150);
nor U6786 (N_6786,In_2853,In_1260);
and U6787 (N_6787,In_4502,In_3171);
or U6788 (N_6788,In_129,In_1447);
nor U6789 (N_6789,In_894,In_1241);
nand U6790 (N_6790,In_3512,In_3500);
xor U6791 (N_6791,In_1265,In_845);
nor U6792 (N_6792,In_1578,In_1644);
nand U6793 (N_6793,In_3302,In_2677);
xnor U6794 (N_6794,In_3821,In_4213);
and U6795 (N_6795,In_3810,In_3256);
nor U6796 (N_6796,In_4131,In_4311);
or U6797 (N_6797,In_954,In_4808);
or U6798 (N_6798,In_3127,In_1265);
xor U6799 (N_6799,In_3444,In_1432);
nand U6800 (N_6800,In_796,In_2747);
and U6801 (N_6801,In_4138,In_727);
xnor U6802 (N_6802,In_295,In_4634);
and U6803 (N_6803,In_1846,In_195);
nor U6804 (N_6804,In_1638,In_2224);
nor U6805 (N_6805,In_4550,In_2202);
and U6806 (N_6806,In_2923,In_1598);
xnor U6807 (N_6807,In_1385,In_402);
nand U6808 (N_6808,In_3795,In_2735);
or U6809 (N_6809,In_1765,In_1917);
or U6810 (N_6810,In_992,In_4631);
and U6811 (N_6811,In_2522,In_2145);
and U6812 (N_6812,In_655,In_2132);
or U6813 (N_6813,In_4299,In_465);
nor U6814 (N_6814,In_1625,In_4956);
nand U6815 (N_6815,In_2407,In_1521);
and U6816 (N_6816,In_4917,In_331);
nand U6817 (N_6817,In_630,In_2172);
nand U6818 (N_6818,In_3676,In_2720);
or U6819 (N_6819,In_1904,In_1180);
and U6820 (N_6820,In_4396,In_2897);
and U6821 (N_6821,In_4288,In_3346);
and U6822 (N_6822,In_1526,In_4015);
and U6823 (N_6823,In_1306,In_1231);
nor U6824 (N_6824,In_1814,In_4799);
or U6825 (N_6825,In_2590,In_4425);
nand U6826 (N_6826,In_1862,In_1642);
nor U6827 (N_6827,In_4428,In_352);
nand U6828 (N_6828,In_1060,In_2452);
nor U6829 (N_6829,In_2605,In_1542);
nand U6830 (N_6830,In_4685,In_3979);
nor U6831 (N_6831,In_2741,In_4425);
nor U6832 (N_6832,In_2824,In_4594);
nor U6833 (N_6833,In_220,In_1249);
and U6834 (N_6834,In_4388,In_257);
nand U6835 (N_6835,In_1375,In_1766);
nor U6836 (N_6836,In_2706,In_422);
and U6837 (N_6837,In_4428,In_2855);
nor U6838 (N_6838,In_1663,In_2617);
nand U6839 (N_6839,In_1919,In_3467);
or U6840 (N_6840,In_2224,In_175);
and U6841 (N_6841,In_2455,In_1048);
nand U6842 (N_6842,In_1212,In_4981);
nand U6843 (N_6843,In_3025,In_96);
nor U6844 (N_6844,In_3812,In_3760);
or U6845 (N_6845,In_1855,In_4208);
xor U6846 (N_6846,In_1903,In_377);
nand U6847 (N_6847,In_2277,In_4242);
xnor U6848 (N_6848,In_4551,In_3290);
and U6849 (N_6849,In_2733,In_3100);
nor U6850 (N_6850,In_2636,In_3404);
nand U6851 (N_6851,In_1394,In_1205);
and U6852 (N_6852,In_2726,In_679);
nor U6853 (N_6853,In_2220,In_1418);
nor U6854 (N_6854,In_1314,In_4333);
nand U6855 (N_6855,In_3111,In_3542);
xor U6856 (N_6856,In_2524,In_584);
and U6857 (N_6857,In_4477,In_656);
nor U6858 (N_6858,In_4169,In_3232);
or U6859 (N_6859,In_216,In_432);
and U6860 (N_6860,In_1824,In_2151);
and U6861 (N_6861,In_3132,In_2311);
nand U6862 (N_6862,In_985,In_2859);
or U6863 (N_6863,In_403,In_29);
nor U6864 (N_6864,In_4732,In_1330);
xnor U6865 (N_6865,In_2581,In_1064);
or U6866 (N_6866,In_1556,In_3080);
nor U6867 (N_6867,In_1214,In_4843);
or U6868 (N_6868,In_1522,In_2193);
or U6869 (N_6869,In_1687,In_4820);
nand U6870 (N_6870,In_17,In_3802);
xor U6871 (N_6871,In_3455,In_879);
xnor U6872 (N_6872,In_1407,In_260);
and U6873 (N_6873,In_1709,In_3894);
and U6874 (N_6874,In_4398,In_4776);
nor U6875 (N_6875,In_927,In_14);
or U6876 (N_6876,In_381,In_2492);
nand U6877 (N_6877,In_547,In_4676);
and U6878 (N_6878,In_2848,In_3733);
and U6879 (N_6879,In_884,In_3096);
nor U6880 (N_6880,In_1098,In_1800);
nor U6881 (N_6881,In_1181,In_1711);
and U6882 (N_6882,In_3768,In_2946);
nor U6883 (N_6883,In_2568,In_1423);
nand U6884 (N_6884,In_764,In_980);
or U6885 (N_6885,In_4276,In_1189);
nor U6886 (N_6886,In_4985,In_764);
or U6887 (N_6887,In_2046,In_4190);
nand U6888 (N_6888,In_3928,In_4117);
xnor U6889 (N_6889,In_4570,In_379);
and U6890 (N_6890,In_3500,In_1226);
or U6891 (N_6891,In_2530,In_3726);
or U6892 (N_6892,In_828,In_132);
and U6893 (N_6893,In_1151,In_220);
nand U6894 (N_6894,In_2437,In_4396);
nand U6895 (N_6895,In_310,In_3847);
and U6896 (N_6896,In_2199,In_54);
nand U6897 (N_6897,In_3661,In_574);
nand U6898 (N_6898,In_2728,In_3731);
and U6899 (N_6899,In_1862,In_374);
or U6900 (N_6900,In_1856,In_4920);
and U6901 (N_6901,In_680,In_820);
xnor U6902 (N_6902,In_1130,In_2598);
nor U6903 (N_6903,In_3020,In_3692);
nor U6904 (N_6904,In_3832,In_4789);
nor U6905 (N_6905,In_857,In_1071);
xnor U6906 (N_6906,In_127,In_1145);
or U6907 (N_6907,In_4407,In_4915);
nor U6908 (N_6908,In_839,In_2279);
nand U6909 (N_6909,In_3318,In_3693);
and U6910 (N_6910,In_2757,In_2389);
nor U6911 (N_6911,In_641,In_4686);
nor U6912 (N_6912,In_4569,In_3559);
and U6913 (N_6913,In_2734,In_3085);
or U6914 (N_6914,In_3148,In_1572);
nand U6915 (N_6915,In_536,In_4755);
nand U6916 (N_6916,In_4428,In_4054);
and U6917 (N_6917,In_3331,In_3767);
nor U6918 (N_6918,In_2276,In_2052);
nor U6919 (N_6919,In_3413,In_2880);
xor U6920 (N_6920,In_1954,In_1517);
nand U6921 (N_6921,In_3935,In_539);
nand U6922 (N_6922,In_1045,In_4500);
nand U6923 (N_6923,In_2265,In_1215);
nor U6924 (N_6924,In_2398,In_993);
nand U6925 (N_6925,In_1964,In_2066);
or U6926 (N_6926,In_1920,In_4531);
nor U6927 (N_6927,In_2172,In_628);
nor U6928 (N_6928,In_1592,In_3509);
xor U6929 (N_6929,In_3076,In_70);
or U6930 (N_6930,In_695,In_2428);
xor U6931 (N_6931,In_4069,In_2808);
nor U6932 (N_6932,In_1521,In_1889);
nand U6933 (N_6933,In_2736,In_4335);
nor U6934 (N_6934,In_3568,In_2213);
nor U6935 (N_6935,In_2057,In_830);
nor U6936 (N_6936,In_2486,In_2851);
or U6937 (N_6937,In_4980,In_3025);
and U6938 (N_6938,In_4888,In_2092);
xor U6939 (N_6939,In_603,In_111);
xnor U6940 (N_6940,In_580,In_3949);
nand U6941 (N_6941,In_3104,In_1509);
and U6942 (N_6942,In_4137,In_2224);
or U6943 (N_6943,In_2027,In_577);
nand U6944 (N_6944,In_4025,In_3125);
nand U6945 (N_6945,In_4554,In_4684);
and U6946 (N_6946,In_1624,In_387);
or U6947 (N_6947,In_1059,In_678);
nor U6948 (N_6948,In_3649,In_2941);
xor U6949 (N_6949,In_3820,In_4776);
and U6950 (N_6950,In_2365,In_6);
and U6951 (N_6951,In_4124,In_3647);
or U6952 (N_6952,In_609,In_4265);
nand U6953 (N_6953,In_4932,In_3329);
and U6954 (N_6954,In_4765,In_16);
and U6955 (N_6955,In_2916,In_925);
nor U6956 (N_6956,In_2905,In_852);
nand U6957 (N_6957,In_1186,In_1959);
and U6958 (N_6958,In_4481,In_2121);
or U6959 (N_6959,In_962,In_4526);
nand U6960 (N_6960,In_4787,In_1879);
nor U6961 (N_6961,In_4197,In_3094);
or U6962 (N_6962,In_2807,In_2507);
nand U6963 (N_6963,In_1077,In_2694);
or U6964 (N_6964,In_3981,In_2147);
and U6965 (N_6965,In_4928,In_4803);
and U6966 (N_6966,In_3708,In_2510);
and U6967 (N_6967,In_2215,In_3765);
nor U6968 (N_6968,In_2350,In_4833);
nor U6969 (N_6969,In_1728,In_836);
nor U6970 (N_6970,In_2176,In_3377);
and U6971 (N_6971,In_2842,In_1746);
nor U6972 (N_6972,In_3049,In_2181);
and U6973 (N_6973,In_392,In_2136);
or U6974 (N_6974,In_434,In_183);
nand U6975 (N_6975,In_2954,In_363);
nand U6976 (N_6976,In_888,In_4525);
and U6977 (N_6977,In_4747,In_4523);
or U6978 (N_6978,In_2815,In_3166);
and U6979 (N_6979,In_4088,In_1799);
xnor U6980 (N_6980,In_3446,In_430);
and U6981 (N_6981,In_1956,In_341);
or U6982 (N_6982,In_712,In_2028);
nor U6983 (N_6983,In_1469,In_798);
or U6984 (N_6984,In_1968,In_4322);
and U6985 (N_6985,In_2589,In_4347);
or U6986 (N_6986,In_2057,In_1332);
or U6987 (N_6987,In_750,In_32);
nand U6988 (N_6988,In_2588,In_3348);
or U6989 (N_6989,In_4741,In_57);
nand U6990 (N_6990,In_4302,In_2928);
nand U6991 (N_6991,In_4675,In_2119);
and U6992 (N_6992,In_2149,In_1855);
xnor U6993 (N_6993,In_3197,In_2992);
or U6994 (N_6994,In_3516,In_2293);
and U6995 (N_6995,In_1836,In_2474);
nor U6996 (N_6996,In_1722,In_4763);
nand U6997 (N_6997,In_2819,In_1781);
nand U6998 (N_6998,In_2469,In_3073);
xor U6999 (N_6999,In_3624,In_1973);
nor U7000 (N_7000,In_2244,In_3121);
xnor U7001 (N_7001,In_1081,In_1238);
xnor U7002 (N_7002,In_4001,In_4080);
or U7003 (N_7003,In_3649,In_3429);
nor U7004 (N_7004,In_3554,In_895);
xnor U7005 (N_7005,In_4567,In_1438);
nor U7006 (N_7006,In_95,In_3798);
xnor U7007 (N_7007,In_610,In_460);
nand U7008 (N_7008,In_1821,In_4001);
nand U7009 (N_7009,In_383,In_652);
nand U7010 (N_7010,In_2217,In_4518);
and U7011 (N_7011,In_3574,In_648);
or U7012 (N_7012,In_1217,In_3341);
nand U7013 (N_7013,In_3392,In_292);
or U7014 (N_7014,In_4451,In_2820);
nor U7015 (N_7015,In_2990,In_2062);
nor U7016 (N_7016,In_4596,In_3653);
nand U7017 (N_7017,In_2773,In_3287);
nand U7018 (N_7018,In_2682,In_2920);
nor U7019 (N_7019,In_3829,In_165);
or U7020 (N_7020,In_505,In_3435);
and U7021 (N_7021,In_620,In_3917);
nand U7022 (N_7022,In_2325,In_785);
or U7023 (N_7023,In_1820,In_782);
nand U7024 (N_7024,In_3522,In_4289);
nand U7025 (N_7025,In_4463,In_2721);
nor U7026 (N_7026,In_244,In_677);
nand U7027 (N_7027,In_733,In_4739);
or U7028 (N_7028,In_4229,In_4179);
nand U7029 (N_7029,In_3848,In_1190);
nand U7030 (N_7030,In_3207,In_4735);
or U7031 (N_7031,In_4995,In_3004);
nor U7032 (N_7032,In_700,In_761);
nand U7033 (N_7033,In_3410,In_1553);
and U7034 (N_7034,In_2230,In_4422);
nor U7035 (N_7035,In_3312,In_3982);
nor U7036 (N_7036,In_3925,In_662);
or U7037 (N_7037,In_414,In_3147);
nand U7038 (N_7038,In_1638,In_3719);
nand U7039 (N_7039,In_1342,In_2599);
nor U7040 (N_7040,In_2115,In_534);
and U7041 (N_7041,In_1718,In_3314);
and U7042 (N_7042,In_4972,In_3576);
or U7043 (N_7043,In_2665,In_1131);
or U7044 (N_7044,In_1984,In_745);
nand U7045 (N_7045,In_3358,In_549);
xnor U7046 (N_7046,In_377,In_853);
nand U7047 (N_7047,In_166,In_2062);
and U7048 (N_7048,In_1960,In_2908);
and U7049 (N_7049,In_116,In_2524);
nor U7050 (N_7050,In_2147,In_1634);
xor U7051 (N_7051,In_2765,In_1721);
xor U7052 (N_7052,In_399,In_3911);
or U7053 (N_7053,In_2874,In_4365);
or U7054 (N_7054,In_4214,In_305);
or U7055 (N_7055,In_1202,In_120);
nand U7056 (N_7056,In_806,In_2499);
nand U7057 (N_7057,In_1581,In_2211);
nor U7058 (N_7058,In_463,In_2709);
nor U7059 (N_7059,In_3980,In_2666);
xnor U7060 (N_7060,In_4588,In_3075);
nor U7061 (N_7061,In_4930,In_1315);
or U7062 (N_7062,In_3473,In_794);
nor U7063 (N_7063,In_2471,In_648);
nor U7064 (N_7064,In_4730,In_4582);
or U7065 (N_7065,In_1482,In_919);
and U7066 (N_7066,In_1340,In_3786);
and U7067 (N_7067,In_2295,In_4967);
nor U7068 (N_7068,In_2056,In_718);
nand U7069 (N_7069,In_3303,In_1942);
nand U7070 (N_7070,In_1396,In_4127);
nand U7071 (N_7071,In_2260,In_3229);
and U7072 (N_7072,In_2593,In_3092);
or U7073 (N_7073,In_222,In_4787);
and U7074 (N_7074,In_3706,In_3899);
nor U7075 (N_7075,In_2850,In_2744);
and U7076 (N_7076,In_1870,In_4231);
nor U7077 (N_7077,In_3236,In_2720);
or U7078 (N_7078,In_2199,In_1679);
nor U7079 (N_7079,In_2400,In_4661);
and U7080 (N_7080,In_2167,In_1964);
nand U7081 (N_7081,In_3083,In_4912);
and U7082 (N_7082,In_3843,In_616);
xor U7083 (N_7083,In_4730,In_1731);
nand U7084 (N_7084,In_2544,In_1452);
and U7085 (N_7085,In_3789,In_985);
and U7086 (N_7086,In_1280,In_2631);
nand U7087 (N_7087,In_2222,In_2883);
xor U7088 (N_7088,In_1142,In_988);
and U7089 (N_7089,In_209,In_4496);
xor U7090 (N_7090,In_4745,In_495);
and U7091 (N_7091,In_341,In_3278);
and U7092 (N_7092,In_1896,In_2228);
nor U7093 (N_7093,In_4209,In_3359);
nor U7094 (N_7094,In_2322,In_4419);
xnor U7095 (N_7095,In_2319,In_3271);
or U7096 (N_7096,In_323,In_1570);
nand U7097 (N_7097,In_4994,In_3033);
xor U7098 (N_7098,In_4927,In_3294);
and U7099 (N_7099,In_1787,In_2849);
nor U7100 (N_7100,In_608,In_784);
and U7101 (N_7101,In_3454,In_1585);
nand U7102 (N_7102,In_456,In_2829);
and U7103 (N_7103,In_4102,In_1504);
nand U7104 (N_7104,In_2543,In_1263);
or U7105 (N_7105,In_2461,In_1090);
and U7106 (N_7106,In_3625,In_1113);
and U7107 (N_7107,In_3563,In_3641);
and U7108 (N_7108,In_2830,In_3083);
nor U7109 (N_7109,In_354,In_3132);
or U7110 (N_7110,In_475,In_4324);
nor U7111 (N_7111,In_1558,In_3998);
nand U7112 (N_7112,In_3203,In_3671);
nor U7113 (N_7113,In_3943,In_802);
nand U7114 (N_7114,In_3519,In_1419);
xor U7115 (N_7115,In_576,In_266);
nand U7116 (N_7116,In_3934,In_2604);
nand U7117 (N_7117,In_2497,In_4676);
or U7118 (N_7118,In_1263,In_66);
nand U7119 (N_7119,In_3396,In_2162);
or U7120 (N_7120,In_4515,In_982);
nor U7121 (N_7121,In_4217,In_3560);
nor U7122 (N_7122,In_2756,In_617);
nand U7123 (N_7123,In_564,In_1743);
and U7124 (N_7124,In_1461,In_1119);
nor U7125 (N_7125,In_4663,In_2040);
and U7126 (N_7126,In_4531,In_471);
xnor U7127 (N_7127,In_674,In_185);
xnor U7128 (N_7128,In_1709,In_943);
nand U7129 (N_7129,In_963,In_3681);
xnor U7130 (N_7130,In_1690,In_405);
and U7131 (N_7131,In_468,In_2119);
or U7132 (N_7132,In_2661,In_1713);
nand U7133 (N_7133,In_1082,In_2605);
nand U7134 (N_7134,In_3238,In_4152);
nor U7135 (N_7135,In_4408,In_3529);
nor U7136 (N_7136,In_271,In_4520);
and U7137 (N_7137,In_4256,In_1639);
nor U7138 (N_7138,In_3338,In_2068);
nand U7139 (N_7139,In_2416,In_4625);
nor U7140 (N_7140,In_2720,In_4072);
and U7141 (N_7141,In_3443,In_2992);
or U7142 (N_7142,In_3292,In_400);
and U7143 (N_7143,In_2647,In_1957);
or U7144 (N_7144,In_1294,In_3010);
and U7145 (N_7145,In_179,In_2367);
or U7146 (N_7146,In_1860,In_1636);
nor U7147 (N_7147,In_2110,In_4668);
or U7148 (N_7148,In_1394,In_2405);
and U7149 (N_7149,In_289,In_641);
nor U7150 (N_7150,In_593,In_1176);
nand U7151 (N_7151,In_848,In_1583);
or U7152 (N_7152,In_1177,In_1277);
nor U7153 (N_7153,In_3346,In_4184);
or U7154 (N_7154,In_913,In_213);
xnor U7155 (N_7155,In_1459,In_2029);
nor U7156 (N_7156,In_2101,In_1517);
and U7157 (N_7157,In_133,In_4867);
nor U7158 (N_7158,In_374,In_362);
nand U7159 (N_7159,In_1167,In_3152);
and U7160 (N_7160,In_1529,In_418);
or U7161 (N_7161,In_3058,In_965);
nand U7162 (N_7162,In_2213,In_2410);
or U7163 (N_7163,In_4435,In_2935);
nor U7164 (N_7164,In_3108,In_1595);
and U7165 (N_7165,In_4353,In_1032);
nor U7166 (N_7166,In_2626,In_1958);
nor U7167 (N_7167,In_3777,In_2830);
nor U7168 (N_7168,In_416,In_4940);
nor U7169 (N_7169,In_2967,In_436);
or U7170 (N_7170,In_577,In_3493);
and U7171 (N_7171,In_3616,In_838);
nor U7172 (N_7172,In_4626,In_3016);
and U7173 (N_7173,In_4042,In_2103);
and U7174 (N_7174,In_4967,In_3399);
and U7175 (N_7175,In_352,In_2949);
and U7176 (N_7176,In_3669,In_1054);
nand U7177 (N_7177,In_4205,In_2875);
and U7178 (N_7178,In_3463,In_2792);
nor U7179 (N_7179,In_3635,In_149);
nor U7180 (N_7180,In_3045,In_4967);
or U7181 (N_7181,In_523,In_2541);
nor U7182 (N_7182,In_493,In_3132);
nor U7183 (N_7183,In_505,In_879);
or U7184 (N_7184,In_3893,In_4162);
or U7185 (N_7185,In_1010,In_2120);
or U7186 (N_7186,In_174,In_3352);
and U7187 (N_7187,In_1706,In_1893);
nand U7188 (N_7188,In_2016,In_3471);
nand U7189 (N_7189,In_4346,In_3167);
nor U7190 (N_7190,In_3208,In_1663);
nand U7191 (N_7191,In_970,In_3860);
and U7192 (N_7192,In_4151,In_4896);
and U7193 (N_7193,In_3079,In_3722);
nand U7194 (N_7194,In_2784,In_4344);
nand U7195 (N_7195,In_2894,In_3725);
and U7196 (N_7196,In_3875,In_1152);
nand U7197 (N_7197,In_2873,In_4881);
nand U7198 (N_7198,In_2820,In_3033);
or U7199 (N_7199,In_2018,In_3451);
or U7200 (N_7200,In_4763,In_4725);
xnor U7201 (N_7201,In_758,In_2965);
nor U7202 (N_7202,In_2790,In_4911);
and U7203 (N_7203,In_3063,In_4707);
xor U7204 (N_7204,In_1210,In_2777);
nand U7205 (N_7205,In_185,In_957);
nor U7206 (N_7206,In_3579,In_2182);
or U7207 (N_7207,In_4894,In_2597);
nor U7208 (N_7208,In_3130,In_1634);
or U7209 (N_7209,In_2753,In_988);
and U7210 (N_7210,In_1463,In_2022);
nor U7211 (N_7211,In_1171,In_3815);
nor U7212 (N_7212,In_1830,In_2852);
nand U7213 (N_7213,In_4742,In_4478);
or U7214 (N_7214,In_2215,In_4811);
nor U7215 (N_7215,In_2927,In_1186);
or U7216 (N_7216,In_1548,In_4147);
nand U7217 (N_7217,In_4599,In_559);
nor U7218 (N_7218,In_3136,In_3966);
xor U7219 (N_7219,In_1235,In_2442);
and U7220 (N_7220,In_637,In_1023);
and U7221 (N_7221,In_1273,In_4001);
or U7222 (N_7222,In_1630,In_938);
xor U7223 (N_7223,In_416,In_2592);
and U7224 (N_7224,In_3688,In_684);
and U7225 (N_7225,In_2200,In_1610);
or U7226 (N_7226,In_1544,In_882);
and U7227 (N_7227,In_1201,In_278);
nor U7228 (N_7228,In_3628,In_4431);
xnor U7229 (N_7229,In_1259,In_1733);
or U7230 (N_7230,In_4030,In_4432);
nand U7231 (N_7231,In_855,In_728);
xnor U7232 (N_7232,In_992,In_1487);
nand U7233 (N_7233,In_1159,In_3944);
or U7234 (N_7234,In_3009,In_3906);
or U7235 (N_7235,In_2958,In_4664);
and U7236 (N_7236,In_3136,In_3553);
xor U7237 (N_7237,In_4865,In_4804);
nor U7238 (N_7238,In_2089,In_4665);
nand U7239 (N_7239,In_2710,In_600);
and U7240 (N_7240,In_4759,In_543);
nand U7241 (N_7241,In_11,In_3170);
and U7242 (N_7242,In_4941,In_1482);
xor U7243 (N_7243,In_4861,In_3852);
or U7244 (N_7244,In_2806,In_36);
nor U7245 (N_7245,In_1208,In_225);
nor U7246 (N_7246,In_4829,In_1847);
and U7247 (N_7247,In_949,In_4662);
and U7248 (N_7248,In_2594,In_4970);
or U7249 (N_7249,In_3815,In_1997);
or U7250 (N_7250,In_4269,In_1794);
nand U7251 (N_7251,In_2473,In_4184);
nor U7252 (N_7252,In_3084,In_4535);
or U7253 (N_7253,In_989,In_1629);
and U7254 (N_7254,In_1738,In_2584);
or U7255 (N_7255,In_3649,In_4027);
or U7256 (N_7256,In_116,In_192);
nand U7257 (N_7257,In_371,In_2883);
or U7258 (N_7258,In_532,In_1040);
nor U7259 (N_7259,In_601,In_3264);
or U7260 (N_7260,In_1081,In_4513);
and U7261 (N_7261,In_3665,In_3382);
or U7262 (N_7262,In_4784,In_789);
or U7263 (N_7263,In_1069,In_1600);
or U7264 (N_7264,In_757,In_3469);
nand U7265 (N_7265,In_3569,In_4729);
or U7266 (N_7266,In_2145,In_4742);
and U7267 (N_7267,In_3802,In_3892);
xor U7268 (N_7268,In_3292,In_3662);
nor U7269 (N_7269,In_1293,In_593);
nand U7270 (N_7270,In_2441,In_782);
nor U7271 (N_7271,In_4780,In_4295);
nand U7272 (N_7272,In_3988,In_3493);
nor U7273 (N_7273,In_129,In_431);
and U7274 (N_7274,In_1630,In_4821);
and U7275 (N_7275,In_1347,In_1819);
nand U7276 (N_7276,In_2765,In_2820);
nor U7277 (N_7277,In_3098,In_914);
nor U7278 (N_7278,In_3146,In_1987);
and U7279 (N_7279,In_2313,In_4972);
xor U7280 (N_7280,In_3902,In_4257);
nor U7281 (N_7281,In_2325,In_1552);
nor U7282 (N_7282,In_4942,In_3319);
and U7283 (N_7283,In_4509,In_2014);
or U7284 (N_7284,In_2453,In_2953);
nor U7285 (N_7285,In_2217,In_16);
nor U7286 (N_7286,In_696,In_4172);
and U7287 (N_7287,In_2457,In_4666);
nor U7288 (N_7288,In_228,In_582);
xnor U7289 (N_7289,In_3873,In_2511);
or U7290 (N_7290,In_4326,In_1728);
nor U7291 (N_7291,In_990,In_3899);
nand U7292 (N_7292,In_3898,In_736);
or U7293 (N_7293,In_2731,In_3548);
or U7294 (N_7294,In_3403,In_3918);
nand U7295 (N_7295,In_3723,In_2152);
nor U7296 (N_7296,In_3302,In_4020);
or U7297 (N_7297,In_1492,In_2869);
xor U7298 (N_7298,In_1716,In_1854);
nor U7299 (N_7299,In_2778,In_2503);
nor U7300 (N_7300,In_2239,In_541);
nor U7301 (N_7301,In_4568,In_4864);
or U7302 (N_7302,In_394,In_2986);
or U7303 (N_7303,In_285,In_2250);
and U7304 (N_7304,In_2401,In_1363);
nor U7305 (N_7305,In_292,In_2050);
or U7306 (N_7306,In_89,In_4696);
and U7307 (N_7307,In_2671,In_2270);
nor U7308 (N_7308,In_3057,In_4198);
nor U7309 (N_7309,In_613,In_4259);
nand U7310 (N_7310,In_573,In_9);
nor U7311 (N_7311,In_4138,In_4858);
xnor U7312 (N_7312,In_1986,In_182);
and U7313 (N_7313,In_32,In_4827);
or U7314 (N_7314,In_763,In_3552);
nand U7315 (N_7315,In_3549,In_1476);
nand U7316 (N_7316,In_4779,In_4427);
nand U7317 (N_7317,In_226,In_4945);
and U7318 (N_7318,In_2465,In_4774);
and U7319 (N_7319,In_4254,In_3845);
and U7320 (N_7320,In_3203,In_1066);
or U7321 (N_7321,In_2820,In_3560);
or U7322 (N_7322,In_4968,In_132);
or U7323 (N_7323,In_256,In_1082);
nor U7324 (N_7324,In_2401,In_646);
and U7325 (N_7325,In_2313,In_1186);
and U7326 (N_7326,In_3203,In_4849);
nand U7327 (N_7327,In_1634,In_470);
and U7328 (N_7328,In_824,In_817);
nor U7329 (N_7329,In_2477,In_2673);
nor U7330 (N_7330,In_1254,In_1716);
and U7331 (N_7331,In_2461,In_4575);
nor U7332 (N_7332,In_2016,In_3801);
nor U7333 (N_7333,In_2863,In_454);
nor U7334 (N_7334,In_1285,In_3189);
xor U7335 (N_7335,In_2020,In_3784);
or U7336 (N_7336,In_2808,In_1909);
xnor U7337 (N_7337,In_414,In_3700);
nor U7338 (N_7338,In_3726,In_987);
nor U7339 (N_7339,In_3363,In_4220);
and U7340 (N_7340,In_3091,In_2698);
and U7341 (N_7341,In_3023,In_3191);
and U7342 (N_7342,In_798,In_4781);
or U7343 (N_7343,In_3523,In_2800);
or U7344 (N_7344,In_3456,In_180);
or U7345 (N_7345,In_4764,In_1251);
or U7346 (N_7346,In_602,In_2705);
nand U7347 (N_7347,In_3243,In_2534);
nand U7348 (N_7348,In_3302,In_133);
nand U7349 (N_7349,In_4318,In_3468);
nand U7350 (N_7350,In_79,In_2415);
nor U7351 (N_7351,In_549,In_4676);
nand U7352 (N_7352,In_3084,In_4198);
or U7353 (N_7353,In_1219,In_3610);
and U7354 (N_7354,In_626,In_2430);
nor U7355 (N_7355,In_4428,In_479);
nand U7356 (N_7356,In_1862,In_745);
or U7357 (N_7357,In_832,In_2283);
nand U7358 (N_7358,In_4409,In_155);
xor U7359 (N_7359,In_807,In_128);
nor U7360 (N_7360,In_4761,In_4391);
nand U7361 (N_7361,In_2563,In_3106);
nand U7362 (N_7362,In_1577,In_1351);
nor U7363 (N_7363,In_4126,In_4690);
and U7364 (N_7364,In_3072,In_525);
or U7365 (N_7365,In_2976,In_3679);
nand U7366 (N_7366,In_4700,In_2926);
and U7367 (N_7367,In_239,In_2985);
nor U7368 (N_7368,In_957,In_4322);
or U7369 (N_7369,In_1114,In_2855);
nor U7370 (N_7370,In_4151,In_47);
nor U7371 (N_7371,In_654,In_2954);
nand U7372 (N_7372,In_1618,In_3769);
and U7373 (N_7373,In_389,In_4105);
and U7374 (N_7374,In_1941,In_2388);
or U7375 (N_7375,In_1390,In_1857);
or U7376 (N_7376,In_2945,In_4825);
or U7377 (N_7377,In_4003,In_3112);
nor U7378 (N_7378,In_2111,In_778);
and U7379 (N_7379,In_3697,In_3753);
or U7380 (N_7380,In_3640,In_4630);
nand U7381 (N_7381,In_3295,In_3570);
or U7382 (N_7382,In_1516,In_4318);
nor U7383 (N_7383,In_4288,In_2521);
xor U7384 (N_7384,In_543,In_611);
and U7385 (N_7385,In_536,In_4012);
nand U7386 (N_7386,In_2387,In_4862);
or U7387 (N_7387,In_4625,In_1722);
nand U7388 (N_7388,In_4890,In_2097);
or U7389 (N_7389,In_2872,In_2941);
and U7390 (N_7390,In_4065,In_582);
or U7391 (N_7391,In_791,In_1107);
nand U7392 (N_7392,In_2193,In_3790);
or U7393 (N_7393,In_116,In_1041);
or U7394 (N_7394,In_2575,In_917);
nand U7395 (N_7395,In_1537,In_1571);
xor U7396 (N_7396,In_556,In_528);
or U7397 (N_7397,In_3634,In_4185);
xor U7398 (N_7398,In_28,In_4141);
or U7399 (N_7399,In_3020,In_2574);
nor U7400 (N_7400,In_4980,In_524);
and U7401 (N_7401,In_722,In_1479);
or U7402 (N_7402,In_594,In_2347);
and U7403 (N_7403,In_1941,In_1956);
nand U7404 (N_7404,In_3562,In_660);
and U7405 (N_7405,In_4696,In_4590);
nor U7406 (N_7406,In_2447,In_2099);
nand U7407 (N_7407,In_2161,In_1815);
nor U7408 (N_7408,In_3239,In_4393);
and U7409 (N_7409,In_2655,In_3638);
or U7410 (N_7410,In_1535,In_985);
or U7411 (N_7411,In_2280,In_4135);
nor U7412 (N_7412,In_4388,In_4497);
or U7413 (N_7413,In_1303,In_1279);
and U7414 (N_7414,In_4025,In_3965);
nand U7415 (N_7415,In_944,In_4922);
nor U7416 (N_7416,In_1238,In_14);
or U7417 (N_7417,In_711,In_377);
or U7418 (N_7418,In_404,In_1438);
and U7419 (N_7419,In_2756,In_4074);
nor U7420 (N_7420,In_773,In_1758);
nor U7421 (N_7421,In_472,In_54);
and U7422 (N_7422,In_3008,In_3645);
and U7423 (N_7423,In_327,In_4848);
nor U7424 (N_7424,In_3820,In_4825);
xnor U7425 (N_7425,In_1030,In_3698);
and U7426 (N_7426,In_122,In_4252);
nand U7427 (N_7427,In_4347,In_2961);
nor U7428 (N_7428,In_3230,In_4241);
nand U7429 (N_7429,In_2965,In_2320);
nor U7430 (N_7430,In_1011,In_2648);
xor U7431 (N_7431,In_2281,In_3623);
xor U7432 (N_7432,In_2942,In_976);
or U7433 (N_7433,In_2846,In_2820);
nor U7434 (N_7434,In_895,In_434);
and U7435 (N_7435,In_3006,In_1610);
or U7436 (N_7436,In_3788,In_3195);
xor U7437 (N_7437,In_2191,In_3526);
nor U7438 (N_7438,In_2783,In_1640);
nand U7439 (N_7439,In_4873,In_1232);
or U7440 (N_7440,In_4371,In_430);
nor U7441 (N_7441,In_1526,In_938);
xor U7442 (N_7442,In_1735,In_1890);
or U7443 (N_7443,In_1717,In_1952);
nand U7444 (N_7444,In_1257,In_792);
or U7445 (N_7445,In_2125,In_30);
nand U7446 (N_7446,In_435,In_3257);
nand U7447 (N_7447,In_3491,In_849);
or U7448 (N_7448,In_4507,In_1012);
or U7449 (N_7449,In_320,In_2571);
and U7450 (N_7450,In_383,In_2767);
xnor U7451 (N_7451,In_1557,In_1959);
nor U7452 (N_7452,In_55,In_2151);
xnor U7453 (N_7453,In_691,In_3353);
or U7454 (N_7454,In_3091,In_2485);
or U7455 (N_7455,In_3996,In_893);
xnor U7456 (N_7456,In_4505,In_3046);
nor U7457 (N_7457,In_4271,In_3303);
nor U7458 (N_7458,In_1540,In_2815);
and U7459 (N_7459,In_4134,In_2421);
and U7460 (N_7460,In_2636,In_122);
xor U7461 (N_7461,In_901,In_1050);
and U7462 (N_7462,In_2251,In_3209);
and U7463 (N_7463,In_2073,In_1877);
nand U7464 (N_7464,In_4600,In_607);
or U7465 (N_7465,In_4153,In_2511);
nor U7466 (N_7466,In_465,In_3855);
or U7467 (N_7467,In_36,In_1340);
xor U7468 (N_7468,In_1411,In_2502);
nand U7469 (N_7469,In_1269,In_902);
or U7470 (N_7470,In_2263,In_1718);
nand U7471 (N_7471,In_384,In_4371);
or U7472 (N_7472,In_1573,In_1926);
and U7473 (N_7473,In_1928,In_210);
nor U7474 (N_7474,In_3303,In_2935);
or U7475 (N_7475,In_2682,In_2132);
xnor U7476 (N_7476,In_249,In_2987);
nand U7477 (N_7477,In_1853,In_3982);
nor U7478 (N_7478,In_1452,In_4685);
xor U7479 (N_7479,In_4735,In_2818);
and U7480 (N_7480,In_2605,In_3332);
nor U7481 (N_7481,In_1784,In_4031);
and U7482 (N_7482,In_1494,In_1218);
and U7483 (N_7483,In_4574,In_4952);
nand U7484 (N_7484,In_4030,In_4317);
nand U7485 (N_7485,In_3500,In_2109);
nor U7486 (N_7486,In_4554,In_2625);
or U7487 (N_7487,In_3200,In_2884);
nor U7488 (N_7488,In_3220,In_2016);
and U7489 (N_7489,In_1619,In_4391);
and U7490 (N_7490,In_4274,In_923);
and U7491 (N_7491,In_4981,In_1316);
nor U7492 (N_7492,In_68,In_4314);
and U7493 (N_7493,In_2034,In_966);
or U7494 (N_7494,In_2635,In_1900);
nand U7495 (N_7495,In_37,In_690);
nand U7496 (N_7496,In_2413,In_4002);
or U7497 (N_7497,In_4323,In_19);
nor U7498 (N_7498,In_1222,In_4968);
nand U7499 (N_7499,In_3471,In_3959);
and U7500 (N_7500,In_1939,In_2017);
and U7501 (N_7501,In_3282,In_1936);
and U7502 (N_7502,In_989,In_2406);
xnor U7503 (N_7503,In_2703,In_4815);
and U7504 (N_7504,In_471,In_2449);
xnor U7505 (N_7505,In_1855,In_3931);
and U7506 (N_7506,In_3919,In_1585);
or U7507 (N_7507,In_4320,In_4429);
nand U7508 (N_7508,In_3741,In_235);
or U7509 (N_7509,In_4564,In_4375);
nand U7510 (N_7510,In_3468,In_2570);
xor U7511 (N_7511,In_389,In_3342);
nor U7512 (N_7512,In_4347,In_3850);
or U7513 (N_7513,In_3905,In_1584);
and U7514 (N_7514,In_3756,In_78);
or U7515 (N_7515,In_4230,In_3714);
nand U7516 (N_7516,In_1896,In_2794);
and U7517 (N_7517,In_2825,In_1660);
nor U7518 (N_7518,In_595,In_844);
nor U7519 (N_7519,In_2149,In_1803);
nand U7520 (N_7520,In_3582,In_620);
or U7521 (N_7521,In_4502,In_1777);
nor U7522 (N_7522,In_3009,In_2512);
or U7523 (N_7523,In_136,In_1927);
and U7524 (N_7524,In_434,In_1395);
and U7525 (N_7525,In_2578,In_4589);
nor U7526 (N_7526,In_2391,In_1111);
or U7527 (N_7527,In_4563,In_2886);
nor U7528 (N_7528,In_48,In_4119);
nor U7529 (N_7529,In_4978,In_2539);
nor U7530 (N_7530,In_506,In_925);
nand U7531 (N_7531,In_3685,In_878);
nor U7532 (N_7532,In_2083,In_1221);
nor U7533 (N_7533,In_1721,In_2766);
nor U7534 (N_7534,In_708,In_4545);
nand U7535 (N_7535,In_3727,In_3285);
and U7536 (N_7536,In_3799,In_1724);
nand U7537 (N_7537,In_4293,In_3700);
nand U7538 (N_7538,In_1157,In_1528);
and U7539 (N_7539,In_2977,In_1666);
nand U7540 (N_7540,In_562,In_3338);
nand U7541 (N_7541,In_426,In_1105);
or U7542 (N_7542,In_421,In_3213);
nor U7543 (N_7543,In_3775,In_1244);
nand U7544 (N_7544,In_3992,In_1557);
nand U7545 (N_7545,In_4147,In_4150);
xor U7546 (N_7546,In_4924,In_4383);
nand U7547 (N_7547,In_798,In_559);
or U7548 (N_7548,In_4355,In_398);
xnor U7549 (N_7549,In_4778,In_3688);
or U7550 (N_7550,In_711,In_2892);
or U7551 (N_7551,In_4813,In_37);
nor U7552 (N_7552,In_324,In_4376);
and U7553 (N_7553,In_2650,In_477);
and U7554 (N_7554,In_1612,In_2651);
or U7555 (N_7555,In_2101,In_4963);
nand U7556 (N_7556,In_1651,In_2528);
nor U7557 (N_7557,In_2149,In_2999);
or U7558 (N_7558,In_979,In_4879);
and U7559 (N_7559,In_1804,In_1329);
nand U7560 (N_7560,In_3491,In_3023);
and U7561 (N_7561,In_1275,In_2684);
nand U7562 (N_7562,In_1601,In_2191);
nor U7563 (N_7563,In_2740,In_3390);
or U7564 (N_7564,In_196,In_762);
nand U7565 (N_7565,In_3129,In_2840);
nand U7566 (N_7566,In_4846,In_2884);
or U7567 (N_7567,In_4730,In_1490);
nand U7568 (N_7568,In_3970,In_219);
or U7569 (N_7569,In_4360,In_4916);
and U7570 (N_7570,In_3975,In_4184);
nand U7571 (N_7571,In_4018,In_4922);
and U7572 (N_7572,In_4951,In_4885);
and U7573 (N_7573,In_577,In_2880);
or U7574 (N_7574,In_2821,In_1842);
and U7575 (N_7575,In_2971,In_1881);
and U7576 (N_7576,In_2680,In_7);
nand U7577 (N_7577,In_685,In_641);
nand U7578 (N_7578,In_251,In_1537);
nor U7579 (N_7579,In_3008,In_4889);
nor U7580 (N_7580,In_910,In_552);
nand U7581 (N_7581,In_4458,In_1244);
and U7582 (N_7582,In_1723,In_4534);
nand U7583 (N_7583,In_4616,In_3848);
nand U7584 (N_7584,In_2172,In_2780);
nor U7585 (N_7585,In_4571,In_2882);
and U7586 (N_7586,In_3057,In_1529);
xor U7587 (N_7587,In_2466,In_4407);
nand U7588 (N_7588,In_3763,In_723);
and U7589 (N_7589,In_2950,In_189);
and U7590 (N_7590,In_744,In_4528);
and U7591 (N_7591,In_1746,In_3285);
nor U7592 (N_7592,In_298,In_3336);
and U7593 (N_7593,In_352,In_857);
or U7594 (N_7594,In_1618,In_4326);
nor U7595 (N_7595,In_4115,In_802);
xnor U7596 (N_7596,In_493,In_4936);
nand U7597 (N_7597,In_4929,In_4266);
nor U7598 (N_7598,In_4323,In_3624);
nand U7599 (N_7599,In_1240,In_1605);
nand U7600 (N_7600,In_1459,In_4759);
and U7601 (N_7601,In_3886,In_4941);
and U7602 (N_7602,In_4991,In_4137);
xnor U7603 (N_7603,In_14,In_1585);
and U7604 (N_7604,In_2601,In_2172);
nand U7605 (N_7605,In_3091,In_4876);
or U7606 (N_7606,In_1482,In_725);
nand U7607 (N_7607,In_1367,In_3387);
nor U7608 (N_7608,In_1345,In_4543);
and U7609 (N_7609,In_200,In_4419);
nand U7610 (N_7610,In_4602,In_3476);
or U7611 (N_7611,In_2799,In_3401);
nor U7612 (N_7612,In_4349,In_695);
nand U7613 (N_7613,In_269,In_3738);
and U7614 (N_7614,In_4069,In_637);
nor U7615 (N_7615,In_4969,In_2724);
nand U7616 (N_7616,In_1152,In_1601);
nor U7617 (N_7617,In_909,In_2424);
or U7618 (N_7618,In_1503,In_112);
and U7619 (N_7619,In_2663,In_474);
and U7620 (N_7620,In_3686,In_602);
nand U7621 (N_7621,In_814,In_2680);
xnor U7622 (N_7622,In_3479,In_1227);
and U7623 (N_7623,In_891,In_4160);
or U7624 (N_7624,In_1838,In_4821);
nand U7625 (N_7625,In_1225,In_2938);
nand U7626 (N_7626,In_920,In_4412);
and U7627 (N_7627,In_1456,In_1192);
xnor U7628 (N_7628,In_1630,In_4775);
nand U7629 (N_7629,In_1009,In_1864);
nor U7630 (N_7630,In_2013,In_4293);
xor U7631 (N_7631,In_1652,In_1792);
and U7632 (N_7632,In_3376,In_3747);
or U7633 (N_7633,In_4908,In_194);
nand U7634 (N_7634,In_1349,In_597);
nand U7635 (N_7635,In_3850,In_3544);
nor U7636 (N_7636,In_1016,In_2685);
nand U7637 (N_7637,In_3213,In_2069);
nand U7638 (N_7638,In_4814,In_816);
nor U7639 (N_7639,In_1575,In_1808);
and U7640 (N_7640,In_2713,In_2537);
xor U7641 (N_7641,In_2219,In_2197);
or U7642 (N_7642,In_167,In_1608);
or U7643 (N_7643,In_1649,In_1968);
or U7644 (N_7644,In_3928,In_313);
nand U7645 (N_7645,In_1268,In_1946);
and U7646 (N_7646,In_1653,In_4649);
xnor U7647 (N_7647,In_4343,In_4453);
nand U7648 (N_7648,In_950,In_3287);
nor U7649 (N_7649,In_4246,In_350);
nand U7650 (N_7650,In_1031,In_622);
or U7651 (N_7651,In_415,In_3345);
nor U7652 (N_7652,In_249,In_1532);
or U7653 (N_7653,In_120,In_4600);
and U7654 (N_7654,In_1785,In_1134);
nor U7655 (N_7655,In_4970,In_2703);
nand U7656 (N_7656,In_4950,In_3270);
nor U7657 (N_7657,In_3505,In_3591);
and U7658 (N_7658,In_1389,In_3255);
nor U7659 (N_7659,In_922,In_4820);
and U7660 (N_7660,In_820,In_411);
or U7661 (N_7661,In_622,In_102);
nand U7662 (N_7662,In_2008,In_4960);
nand U7663 (N_7663,In_4218,In_3986);
nand U7664 (N_7664,In_4263,In_2363);
nand U7665 (N_7665,In_2946,In_939);
and U7666 (N_7666,In_4700,In_1325);
and U7667 (N_7667,In_1526,In_2748);
nor U7668 (N_7668,In_3753,In_1536);
or U7669 (N_7669,In_1543,In_4978);
nand U7670 (N_7670,In_4861,In_607);
nor U7671 (N_7671,In_2781,In_3931);
and U7672 (N_7672,In_4358,In_4779);
nand U7673 (N_7673,In_1580,In_951);
nor U7674 (N_7674,In_3419,In_3647);
nor U7675 (N_7675,In_2164,In_4484);
nand U7676 (N_7676,In_3817,In_534);
xnor U7677 (N_7677,In_4193,In_1413);
nand U7678 (N_7678,In_4281,In_520);
or U7679 (N_7679,In_3168,In_3867);
nor U7680 (N_7680,In_1362,In_4389);
xor U7681 (N_7681,In_935,In_2252);
or U7682 (N_7682,In_138,In_4720);
nor U7683 (N_7683,In_2123,In_3697);
or U7684 (N_7684,In_2352,In_1631);
or U7685 (N_7685,In_4790,In_4456);
nor U7686 (N_7686,In_381,In_469);
nand U7687 (N_7687,In_909,In_876);
nor U7688 (N_7688,In_4609,In_2811);
xnor U7689 (N_7689,In_1465,In_1918);
and U7690 (N_7690,In_4779,In_4746);
nor U7691 (N_7691,In_2896,In_4853);
nand U7692 (N_7692,In_77,In_2154);
nor U7693 (N_7693,In_3990,In_2536);
or U7694 (N_7694,In_4460,In_1067);
nand U7695 (N_7695,In_2964,In_2690);
and U7696 (N_7696,In_761,In_4596);
nand U7697 (N_7697,In_3431,In_294);
nand U7698 (N_7698,In_4540,In_1775);
nor U7699 (N_7699,In_3161,In_4102);
or U7700 (N_7700,In_859,In_2950);
nor U7701 (N_7701,In_496,In_1491);
and U7702 (N_7702,In_3203,In_318);
nor U7703 (N_7703,In_1607,In_3747);
and U7704 (N_7704,In_4230,In_2901);
nor U7705 (N_7705,In_4946,In_3564);
and U7706 (N_7706,In_1625,In_4898);
or U7707 (N_7707,In_4004,In_519);
and U7708 (N_7708,In_1788,In_3080);
nor U7709 (N_7709,In_3807,In_3879);
nor U7710 (N_7710,In_2636,In_414);
or U7711 (N_7711,In_4386,In_1717);
nand U7712 (N_7712,In_2552,In_1059);
nand U7713 (N_7713,In_1867,In_892);
or U7714 (N_7714,In_4535,In_4814);
nor U7715 (N_7715,In_227,In_978);
nor U7716 (N_7716,In_4798,In_1119);
nand U7717 (N_7717,In_3423,In_2103);
or U7718 (N_7718,In_1421,In_895);
nand U7719 (N_7719,In_4229,In_1220);
nand U7720 (N_7720,In_3422,In_3233);
and U7721 (N_7721,In_138,In_4999);
nand U7722 (N_7722,In_1616,In_4298);
nand U7723 (N_7723,In_1764,In_4533);
nand U7724 (N_7724,In_4205,In_3772);
nand U7725 (N_7725,In_4243,In_1565);
nand U7726 (N_7726,In_1792,In_1461);
and U7727 (N_7727,In_46,In_4025);
nor U7728 (N_7728,In_3704,In_58);
nand U7729 (N_7729,In_3729,In_3283);
or U7730 (N_7730,In_3762,In_3086);
and U7731 (N_7731,In_4344,In_2097);
nor U7732 (N_7732,In_729,In_790);
nor U7733 (N_7733,In_2855,In_3592);
or U7734 (N_7734,In_1208,In_3162);
and U7735 (N_7735,In_583,In_2637);
or U7736 (N_7736,In_3931,In_1661);
and U7737 (N_7737,In_1390,In_3987);
and U7738 (N_7738,In_2102,In_1977);
nand U7739 (N_7739,In_3034,In_945);
xnor U7740 (N_7740,In_1559,In_1727);
and U7741 (N_7741,In_1620,In_3395);
and U7742 (N_7742,In_4367,In_2931);
and U7743 (N_7743,In_2013,In_242);
and U7744 (N_7744,In_4053,In_3275);
nand U7745 (N_7745,In_1977,In_4543);
and U7746 (N_7746,In_2313,In_4871);
nand U7747 (N_7747,In_1711,In_150);
or U7748 (N_7748,In_4151,In_1174);
nor U7749 (N_7749,In_2259,In_615);
or U7750 (N_7750,In_2217,In_4924);
xor U7751 (N_7751,In_24,In_3415);
nand U7752 (N_7752,In_4793,In_4349);
and U7753 (N_7753,In_1446,In_4182);
nor U7754 (N_7754,In_4444,In_1249);
nor U7755 (N_7755,In_1362,In_1728);
nand U7756 (N_7756,In_4762,In_2935);
nand U7757 (N_7757,In_3998,In_1703);
nor U7758 (N_7758,In_3679,In_4629);
nor U7759 (N_7759,In_1608,In_2904);
and U7760 (N_7760,In_448,In_821);
nand U7761 (N_7761,In_3949,In_3619);
and U7762 (N_7762,In_4455,In_3946);
nor U7763 (N_7763,In_4618,In_3149);
or U7764 (N_7764,In_148,In_2395);
and U7765 (N_7765,In_3700,In_2934);
or U7766 (N_7766,In_1686,In_2893);
nor U7767 (N_7767,In_1099,In_4383);
nand U7768 (N_7768,In_4141,In_3847);
nor U7769 (N_7769,In_2143,In_216);
and U7770 (N_7770,In_1516,In_1129);
and U7771 (N_7771,In_4373,In_691);
and U7772 (N_7772,In_93,In_421);
nand U7773 (N_7773,In_2510,In_4359);
and U7774 (N_7774,In_1921,In_4256);
or U7775 (N_7775,In_2906,In_1291);
nand U7776 (N_7776,In_2975,In_1305);
nor U7777 (N_7777,In_1115,In_3492);
and U7778 (N_7778,In_251,In_3375);
nand U7779 (N_7779,In_2253,In_3665);
nand U7780 (N_7780,In_617,In_4849);
or U7781 (N_7781,In_4036,In_344);
and U7782 (N_7782,In_3935,In_227);
or U7783 (N_7783,In_522,In_4708);
nand U7784 (N_7784,In_784,In_2415);
or U7785 (N_7785,In_562,In_2273);
or U7786 (N_7786,In_542,In_4530);
and U7787 (N_7787,In_686,In_2590);
nor U7788 (N_7788,In_4825,In_3343);
or U7789 (N_7789,In_818,In_4794);
and U7790 (N_7790,In_4336,In_4296);
and U7791 (N_7791,In_3720,In_3637);
nand U7792 (N_7792,In_947,In_3256);
nand U7793 (N_7793,In_1052,In_3962);
or U7794 (N_7794,In_826,In_3930);
nand U7795 (N_7795,In_705,In_1534);
nor U7796 (N_7796,In_4262,In_660);
nand U7797 (N_7797,In_3306,In_1610);
and U7798 (N_7798,In_439,In_2512);
or U7799 (N_7799,In_4158,In_3275);
nand U7800 (N_7800,In_3191,In_3642);
and U7801 (N_7801,In_2252,In_3575);
nor U7802 (N_7802,In_4607,In_117);
and U7803 (N_7803,In_2483,In_4777);
nand U7804 (N_7804,In_2552,In_1203);
nor U7805 (N_7805,In_3532,In_2530);
and U7806 (N_7806,In_1598,In_3281);
or U7807 (N_7807,In_3610,In_3572);
and U7808 (N_7808,In_4256,In_3449);
nand U7809 (N_7809,In_4864,In_4589);
or U7810 (N_7810,In_1044,In_732);
and U7811 (N_7811,In_4066,In_3673);
nor U7812 (N_7812,In_1200,In_3410);
nor U7813 (N_7813,In_3788,In_1394);
or U7814 (N_7814,In_2113,In_2670);
or U7815 (N_7815,In_243,In_4170);
and U7816 (N_7816,In_2137,In_4840);
nor U7817 (N_7817,In_1532,In_2214);
xnor U7818 (N_7818,In_211,In_2523);
xor U7819 (N_7819,In_4958,In_4475);
or U7820 (N_7820,In_1755,In_693);
and U7821 (N_7821,In_3068,In_4446);
and U7822 (N_7822,In_3649,In_17);
xor U7823 (N_7823,In_4197,In_4523);
and U7824 (N_7824,In_1859,In_1369);
xor U7825 (N_7825,In_50,In_3457);
nand U7826 (N_7826,In_2823,In_45);
and U7827 (N_7827,In_2249,In_3248);
and U7828 (N_7828,In_2423,In_2683);
nand U7829 (N_7829,In_2474,In_560);
xnor U7830 (N_7830,In_1003,In_927);
or U7831 (N_7831,In_4282,In_3167);
nand U7832 (N_7832,In_3196,In_677);
nor U7833 (N_7833,In_2601,In_4634);
and U7834 (N_7834,In_4894,In_2863);
or U7835 (N_7835,In_4651,In_553);
or U7836 (N_7836,In_85,In_4642);
nor U7837 (N_7837,In_4694,In_1302);
or U7838 (N_7838,In_3529,In_2897);
or U7839 (N_7839,In_4075,In_3439);
or U7840 (N_7840,In_4736,In_4993);
or U7841 (N_7841,In_2413,In_666);
nand U7842 (N_7842,In_2380,In_4449);
nor U7843 (N_7843,In_1259,In_3290);
nand U7844 (N_7844,In_4182,In_2006);
and U7845 (N_7845,In_1417,In_732);
nand U7846 (N_7846,In_4881,In_844);
and U7847 (N_7847,In_4616,In_3113);
nand U7848 (N_7848,In_1860,In_4453);
and U7849 (N_7849,In_3456,In_945);
nor U7850 (N_7850,In_1255,In_4050);
and U7851 (N_7851,In_74,In_3837);
nor U7852 (N_7852,In_421,In_4622);
xor U7853 (N_7853,In_815,In_369);
and U7854 (N_7854,In_3651,In_3399);
nand U7855 (N_7855,In_4673,In_676);
nor U7856 (N_7856,In_3083,In_3585);
nor U7857 (N_7857,In_3982,In_2489);
and U7858 (N_7858,In_115,In_1862);
or U7859 (N_7859,In_3067,In_1501);
nor U7860 (N_7860,In_867,In_2375);
xnor U7861 (N_7861,In_3511,In_1289);
or U7862 (N_7862,In_4940,In_465);
nor U7863 (N_7863,In_4853,In_246);
nor U7864 (N_7864,In_2735,In_4061);
nor U7865 (N_7865,In_2440,In_2711);
and U7866 (N_7866,In_4274,In_2121);
nor U7867 (N_7867,In_1017,In_2829);
and U7868 (N_7868,In_3518,In_4934);
or U7869 (N_7869,In_4453,In_4977);
nor U7870 (N_7870,In_4774,In_3543);
and U7871 (N_7871,In_3891,In_3908);
and U7872 (N_7872,In_1703,In_4318);
and U7873 (N_7873,In_1647,In_1711);
nand U7874 (N_7874,In_3080,In_1638);
or U7875 (N_7875,In_1962,In_4409);
nor U7876 (N_7876,In_2760,In_3313);
and U7877 (N_7877,In_3179,In_1449);
nand U7878 (N_7878,In_1300,In_4333);
or U7879 (N_7879,In_4530,In_1370);
nand U7880 (N_7880,In_4281,In_104);
and U7881 (N_7881,In_4748,In_543);
nand U7882 (N_7882,In_994,In_1559);
and U7883 (N_7883,In_3761,In_2145);
nor U7884 (N_7884,In_145,In_2635);
nand U7885 (N_7885,In_151,In_3801);
nor U7886 (N_7886,In_2604,In_1633);
nand U7887 (N_7887,In_4231,In_1190);
nor U7888 (N_7888,In_3318,In_4945);
or U7889 (N_7889,In_223,In_733);
or U7890 (N_7890,In_1363,In_4278);
or U7891 (N_7891,In_4018,In_1200);
nor U7892 (N_7892,In_3651,In_2978);
nand U7893 (N_7893,In_749,In_3135);
or U7894 (N_7894,In_4936,In_1690);
nor U7895 (N_7895,In_647,In_1861);
nor U7896 (N_7896,In_90,In_3525);
and U7897 (N_7897,In_4802,In_2036);
nor U7898 (N_7898,In_977,In_1779);
or U7899 (N_7899,In_41,In_222);
and U7900 (N_7900,In_1160,In_2529);
nand U7901 (N_7901,In_1250,In_1027);
nand U7902 (N_7902,In_851,In_156);
or U7903 (N_7903,In_1985,In_2800);
nand U7904 (N_7904,In_2658,In_3511);
nor U7905 (N_7905,In_1660,In_1631);
or U7906 (N_7906,In_2335,In_2266);
nor U7907 (N_7907,In_2896,In_526);
nor U7908 (N_7908,In_4917,In_2280);
or U7909 (N_7909,In_2483,In_4355);
and U7910 (N_7910,In_4858,In_2400);
nor U7911 (N_7911,In_348,In_3637);
nand U7912 (N_7912,In_1516,In_3334);
and U7913 (N_7913,In_1510,In_3098);
xor U7914 (N_7914,In_2272,In_2017);
xor U7915 (N_7915,In_4186,In_4598);
nor U7916 (N_7916,In_490,In_2008);
or U7917 (N_7917,In_1060,In_477);
nand U7918 (N_7918,In_4110,In_3103);
nor U7919 (N_7919,In_1041,In_183);
nand U7920 (N_7920,In_3043,In_931);
nand U7921 (N_7921,In_2287,In_2493);
or U7922 (N_7922,In_4755,In_1165);
xnor U7923 (N_7923,In_327,In_4289);
or U7924 (N_7924,In_3184,In_1996);
xor U7925 (N_7925,In_4328,In_1939);
and U7926 (N_7926,In_2149,In_1224);
nor U7927 (N_7927,In_3744,In_2215);
and U7928 (N_7928,In_2741,In_136);
nand U7929 (N_7929,In_3344,In_4985);
nor U7930 (N_7930,In_668,In_2384);
nor U7931 (N_7931,In_1554,In_1901);
nor U7932 (N_7932,In_2456,In_3883);
and U7933 (N_7933,In_3991,In_3103);
nand U7934 (N_7934,In_2165,In_4444);
nand U7935 (N_7935,In_2147,In_1757);
or U7936 (N_7936,In_3844,In_2379);
nor U7937 (N_7937,In_2018,In_2795);
nor U7938 (N_7938,In_233,In_921);
nand U7939 (N_7939,In_458,In_1438);
nor U7940 (N_7940,In_1173,In_700);
xor U7941 (N_7941,In_3596,In_791);
nor U7942 (N_7942,In_2478,In_2439);
nand U7943 (N_7943,In_4921,In_2494);
nor U7944 (N_7944,In_2577,In_1505);
nor U7945 (N_7945,In_4710,In_1902);
nor U7946 (N_7946,In_2175,In_630);
nand U7947 (N_7947,In_2012,In_1021);
and U7948 (N_7948,In_3116,In_4879);
nor U7949 (N_7949,In_3642,In_1037);
nand U7950 (N_7950,In_582,In_1605);
nand U7951 (N_7951,In_3412,In_3275);
or U7952 (N_7952,In_3995,In_3583);
nand U7953 (N_7953,In_4321,In_3036);
nand U7954 (N_7954,In_961,In_3676);
and U7955 (N_7955,In_901,In_1152);
nor U7956 (N_7956,In_2298,In_4543);
nor U7957 (N_7957,In_3982,In_105);
and U7958 (N_7958,In_4101,In_2245);
nor U7959 (N_7959,In_1140,In_892);
or U7960 (N_7960,In_4536,In_2450);
or U7961 (N_7961,In_1388,In_4691);
or U7962 (N_7962,In_865,In_2241);
and U7963 (N_7963,In_1378,In_3056);
nor U7964 (N_7964,In_240,In_707);
or U7965 (N_7965,In_3459,In_3971);
and U7966 (N_7966,In_4524,In_3026);
or U7967 (N_7967,In_3944,In_62);
and U7968 (N_7968,In_590,In_4410);
nor U7969 (N_7969,In_560,In_412);
nand U7970 (N_7970,In_1060,In_3533);
nor U7971 (N_7971,In_3378,In_3781);
or U7972 (N_7972,In_4158,In_4431);
nand U7973 (N_7973,In_2381,In_3125);
nand U7974 (N_7974,In_4815,In_1215);
nor U7975 (N_7975,In_1503,In_3344);
and U7976 (N_7976,In_4987,In_4658);
nor U7977 (N_7977,In_1683,In_4299);
and U7978 (N_7978,In_4849,In_2548);
and U7979 (N_7979,In_4824,In_4238);
xnor U7980 (N_7980,In_2893,In_94);
or U7981 (N_7981,In_2470,In_1519);
and U7982 (N_7982,In_1659,In_4141);
nor U7983 (N_7983,In_2675,In_3837);
nor U7984 (N_7984,In_3945,In_4716);
nor U7985 (N_7985,In_3500,In_1439);
nand U7986 (N_7986,In_4768,In_3368);
or U7987 (N_7987,In_2547,In_4505);
xor U7988 (N_7988,In_3092,In_4069);
and U7989 (N_7989,In_3540,In_1146);
nand U7990 (N_7990,In_1312,In_1283);
nor U7991 (N_7991,In_1218,In_4191);
nor U7992 (N_7992,In_1107,In_2002);
nor U7993 (N_7993,In_2348,In_2546);
and U7994 (N_7994,In_1723,In_153);
nor U7995 (N_7995,In_4847,In_1056);
and U7996 (N_7996,In_1735,In_4999);
or U7997 (N_7997,In_4980,In_4323);
and U7998 (N_7998,In_1135,In_2663);
and U7999 (N_7999,In_136,In_4114);
xnor U8000 (N_8000,In_3541,In_2550);
or U8001 (N_8001,In_801,In_3336);
nor U8002 (N_8002,In_3750,In_1745);
nand U8003 (N_8003,In_3197,In_4846);
and U8004 (N_8004,In_1111,In_2867);
xor U8005 (N_8005,In_2522,In_819);
and U8006 (N_8006,In_1550,In_303);
nand U8007 (N_8007,In_3095,In_1197);
nand U8008 (N_8008,In_3561,In_2744);
nor U8009 (N_8009,In_2772,In_2404);
and U8010 (N_8010,In_3288,In_2957);
and U8011 (N_8011,In_3682,In_3342);
and U8012 (N_8012,In_309,In_4925);
nor U8013 (N_8013,In_2168,In_3425);
or U8014 (N_8014,In_1342,In_228);
or U8015 (N_8015,In_2861,In_832);
nand U8016 (N_8016,In_55,In_4796);
nand U8017 (N_8017,In_4832,In_2129);
and U8018 (N_8018,In_4913,In_4438);
nor U8019 (N_8019,In_3393,In_958);
nor U8020 (N_8020,In_4876,In_4705);
nor U8021 (N_8021,In_405,In_3499);
nand U8022 (N_8022,In_130,In_4429);
xor U8023 (N_8023,In_622,In_1605);
and U8024 (N_8024,In_4719,In_739);
nor U8025 (N_8025,In_4370,In_4987);
nand U8026 (N_8026,In_4971,In_1985);
or U8027 (N_8027,In_856,In_361);
nor U8028 (N_8028,In_1096,In_2445);
xnor U8029 (N_8029,In_1363,In_2095);
nor U8030 (N_8030,In_3118,In_1764);
or U8031 (N_8031,In_2412,In_1401);
nand U8032 (N_8032,In_3037,In_1876);
nor U8033 (N_8033,In_2690,In_993);
nand U8034 (N_8034,In_3172,In_4708);
and U8035 (N_8035,In_1850,In_3711);
xnor U8036 (N_8036,In_1768,In_3879);
nand U8037 (N_8037,In_4057,In_1720);
nand U8038 (N_8038,In_1130,In_561);
and U8039 (N_8039,In_4859,In_3186);
nand U8040 (N_8040,In_3334,In_4661);
and U8041 (N_8041,In_1889,In_4722);
xor U8042 (N_8042,In_3364,In_3406);
and U8043 (N_8043,In_568,In_3012);
or U8044 (N_8044,In_2829,In_3688);
and U8045 (N_8045,In_3735,In_2542);
and U8046 (N_8046,In_1250,In_957);
or U8047 (N_8047,In_1618,In_314);
xor U8048 (N_8048,In_3245,In_483);
or U8049 (N_8049,In_3442,In_3097);
nor U8050 (N_8050,In_548,In_4605);
or U8051 (N_8051,In_308,In_2733);
or U8052 (N_8052,In_3239,In_1224);
or U8053 (N_8053,In_412,In_461);
or U8054 (N_8054,In_4753,In_1276);
nor U8055 (N_8055,In_1555,In_3694);
nor U8056 (N_8056,In_1625,In_1851);
or U8057 (N_8057,In_2233,In_949);
nor U8058 (N_8058,In_3318,In_2546);
nand U8059 (N_8059,In_1888,In_2092);
and U8060 (N_8060,In_3133,In_4228);
nand U8061 (N_8061,In_1660,In_4965);
and U8062 (N_8062,In_1676,In_4455);
nand U8063 (N_8063,In_1180,In_1144);
nand U8064 (N_8064,In_1465,In_4082);
and U8065 (N_8065,In_3136,In_1288);
and U8066 (N_8066,In_4286,In_4415);
or U8067 (N_8067,In_306,In_1476);
or U8068 (N_8068,In_4886,In_1844);
or U8069 (N_8069,In_2249,In_3893);
and U8070 (N_8070,In_3285,In_3896);
nand U8071 (N_8071,In_1292,In_124);
nand U8072 (N_8072,In_187,In_4474);
nor U8073 (N_8073,In_2713,In_3498);
or U8074 (N_8074,In_34,In_3734);
or U8075 (N_8075,In_402,In_1849);
nor U8076 (N_8076,In_4666,In_762);
and U8077 (N_8077,In_2089,In_826);
nor U8078 (N_8078,In_4578,In_146);
nand U8079 (N_8079,In_11,In_2155);
or U8080 (N_8080,In_3140,In_1994);
or U8081 (N_8081,In_901,In_1375);
xor U8082 (N_8082,In_1440,In_3094);
nand U8083 (N_8083,In_1368,In_844);
and U8084 (N_8084,In_4807,In_1708);
and U8085 (N_8085,In_4252,In_2577);
and U8086 (N_8086,In_927,In_215);
xnor U8087 (N_8087,In_2433,In_2829);
and U8088 (N_8088,In_831,In_4881);
or U8089 (N_8089,In_1929,In_757);
or U8090 (N_8090,In_228,In_677);
or U8091 (N_8091,In_292,In_4302);
and U8092 (N_8092,In_884,In_4591);
or U8093 (N_8093,In_139,In_3033);
nor U8094 (N_8094,In_4171,In_3049);
or U8095 (N_8095,In_3403,In_3626);
nand U8096 (N_8096,In_615,In_4150);
nand U8097 (N_8097,In_2586,In_2666);
or U8098 (N_8098,In_745,In_3543);
nand U8099 (N_8099,In_4471,In_2020);
or U8100 (N_8100,In_4823,In_242);
and U8101 (N_8101,In_821,In_3227);
xor U8102 (N_8102,In_363,In_1229);
nand U8103 (N_8103,In_2941,In_4296);
and U8104 (N_8104,In_640,In_3847);
or U8105 (N_8105,In_1009,In_2885);
and U8106 (N_8106,In_1909,In_990);
xor U8107 (N_8107,In_187,In_4996);
nor U8108 (N_8108,In_2606,In_815);
and U8109 (N_8109,In_661,In_555);
xnor U8110 (N_8110,In_2704,In_653);
and U8111 (N_8111,In_754,In_513);
nor U8112 (N_8112,In_3754,In_1299);
nor U8113 (N_8113,In_4668,In_3866);
and U8114 (N_8114,In_4976,In_2416);
or U8115 (N_8115,In_2422,In_4842);
or U8116 (N_8116,In_4584,In_1631);
xnor U8117 (N_8117,In_2090,In_522);
nor U8118 (N_8118,In_205,In_421);
or U8119 (N_8119,In_4150,In_1920);
nand U8120 (N_8120,In_1480,In_387);
and U8121 (N_8121,In_3599,In_3424);
xor U8122 (N_8122,In_3230,In_900);
and U8123 (N_8123,In_980,In_2463);
and U8124 (N_8124,In_1576,In_4871);
and U8125 (N_8125,In_864,In_1588);
or U8126 (N_8126,In_3425,In_1763);
nand U8127 (N_8127,In_2269,In_2373);
nor U8128 (N_8128,In_1536,In_2840);
nor U8129 (N_8129,In_3381,In_2948);
or U8130 (N_8130,In_4993,In_2892);
nand U8131 (N_8131,In_22,In_2951);
nor U8132 (N_8132,In_2457,In_1534);
and U8133 (N_8133,In_863,In_921);
nor U8134 (N_8134,In_1929,In_167);
or U8135 (N_8135,In_4495,In_2402);
xnor U8136 (N_8136,In_4490,In_1663);
or U8137 (N_8137,In_4801,In_567);
nor U8138 (N_8138,In_4425,In_3405);
nor U8139 (N_8139,In_380,In_1131);
xnor U8140 (N_8140,In_671,In_3788);
nor U8141 (N_8141,In_263,In_3142);
or U8142 (N_8142,In_3314,In_1660);
nor U8143 (N_8143,In_4724,In_2383);
or U8144 (N_8144,In_2904,In_3447);
or U8145 (N_8145,In_3556,In_3873);
nand U8146 (N_8146,In_149,In_2676);
and U8147 (N_8147,In_189,In_3695);
xor U8148 (N_8148,In_979,In_2718);
xnor U8149 (N_8149,In_4135,In_231);
or U8150 (N_8150,In_4944,In_3781);
nand U8151 (N_8151,In_82,In_907);
xnor U8152 (N_8152,In_4051,In_2803);
and U8153 (N_8153,In_3003,In_4713);
or U8154 (N_8154,In_3230,In_4151);
and U8155 (N_8155,In_2869,In_3442);
nand U8156 (N_8156,In_3739,In_2285);
nor U8157 (N_8157,In_2584,In_4361);
nand U8158 (N_8158,In_1170,In_4723);
nand U8159 (N_8159,In_235,In_71);
and U8160 (N_8160,In_3785,In_809);
or U8161 (N_8161,In_4429,In_4467);
and U8162 (N_8162,In_4675,In_76);
nand U8163 (N_8163,In_2199,In_423);
nor U8164 (N_8164,In_614,In_3112);
or U8165 (N_8165,In_1165,In_2752);
nor U8166 (N_8166,In_1006,In_3367);
and U8167 (N_8167,In_4831,In_3491);
nor U8168 (N_8168,In_60,In_862);
and U8169 (N_8169,In_3629,In_1921);
or U8170 (N_8170,In_2092,In_4231);
or U8171 (N_8171,In_3904,In_602);
nand U8172 (N_8172,In_4470,In_2695);
or U8173 (N_8173,In_4325,In_1117);
nand U8174 (N_8174,In_3906,In_1975);
or U8175 (N_8175,In_972,In_2225);
nor U8176 (N_8176,In_4048,In_2015);
nand U8177 (N_8177,In_1402,In_3008);
nand U8178 (N_8178,In_978,In_3112);
and U8179 (N_8179,In_4969,In_3012);
or U8180 (N_8180,In_2171,In_4238);
or U8181 (N_8181,In_1617,In_1674);
xnor U8182 (N_8182,In_4842,In_1891);
or U8183 (N_8183,In_3701,In_3033);
and U8184 (N_8184,In_3193,In_3571);
nand U8185 (N_8185,In_1882,In_1390);
nor U8186 (N_8186,In_3558,In_3028);
nor U8187 (N_8187,In_1952,In_3178);
nand U8188 (N_8188,In_444,In_3747);
and U8189 (N_8189,In_4380,In_1286);
or U8190 (N_8190,In_1117,In_3934);
and U8191 (N_8191,In_452,In_4267);
nor U8192 (N_8192,In_836,In_1429);
and U8193 (N_8193,In_4320,In_4966);
nor U8194 (N_8194,In_4469,In_4396);
xor U8195 (N_8195,In_795,In_3801);
and U8196 (N_8196,In_3106,In_732);
nor U8197 (N_8197,In_4013,In_1668);
or U8198 (N_8198,In_4351,In_4084);
xor U8199 (N_8199,In_2808,In_2095);
nor U8200 (N_8200,In_3661,In_1982);
nor U8201 (N_8201,In_2961,In_3629);
nand U8202 (N_8202,In_1128,In_3699);
nor U8203 (N_8203,In_736,In_3616);
or U8204 (N_8204,In_2804,In_3350);
and U8205 (N_8205,In_3312,In_393);
and U8206 (N_8206,In_487,In_2909);
nand U8207 (N_8207,In_437,In_4215);
and U8208 (N_8208,In_1688,In_4936);
or U8209 (N_8209,In_4489,In_3161);
or U8210 (N_8210,In_4020,In_2731);
or U8211 (N_8211,In_4810,In_593);
nand U8212 (N_8212,In_4296,In_59);
and U8213 (N_8213,In_1396,In_157);
and U8214 (N_8214,In_1715,In_1791);
nand U8215 (N_8215,In_4192,In_554);
and U8216 (N_8216,In_3307,In_1130);
and U8217 (N_8217,In_2160,In_3604);
nand U8218 (N_8218,In_4126,In_42);
nand U8219 (N_8219,In_2051,In_3599);
nand U8220 (N_8220,In_2842,In_875);
or U8221 (N_8221,In_3252,In_1912);
nand U8222 (N_8222,In_3294,In_783);
or U8223 (N_8223,In_1525,In_854);
and U8224 (N_8224,In_3688,In_1554);
xor U8225 (N_8225,In_1757,In_798);
and U8226 (N_8226,In_3874,In_3474);
or U8227 (N_8227,In_4533,In_4983);
nand U8228 (N_8228,In_3881,In_4715);
nor U8229 (N_8229,In_2345,In_2983);
and U8230 (N_8230,In_1447,In_4276);
nor U8231 (N_8231,In_283,In_4627);
or U8232 (N_8232,In_4220,In_1115);
nor U8233 (N_8233,In_2497,In_1228);
or U8234 (N_8234,In_1685,In_1249);
xor U8235 (N_8235,In_1394,In_3308);
and U8236 (N_8236,In_3547,In_2439);
nor U8237 (N_8237,In_2945,In_597);
or U8238 (N_8238,In_4267,In_841);
nor U8239 (N_8239,In_2009,In_788);
or U8240 (N_8240,In_1438,In_847);
or U8241 (N_8241,In_2964,In_3424);
nor U8242 (N_8242,In_2146,In_583);
nor U8243 (N_8243,In_2902,In_1257);
nor U8244 (N_8244,In_387,In_2859);
nor U8245 (N_8245,In_1019,In_4051);
and U8246 (N_8246,In_4863,In_3222);
or U8247 (N_8247,In_402,In_4434);
nand U8248 (N_8248,In_3691,In_3156);
xor U8249 (N_8249,In_3473,In_315);
or U8250 (N_8250,In_1238,In_560);
nor U8251 (N_8251,In_3464,In_3082);
xnor U8252 (N_8252,In_3551,In_474);
or U8253 (N_8253,In_1981,In_2822);
xnor U8254 (N_8254,In_2745,In_2143);
nor U8255 (N_8255,In_4919,In_2129);
nor U8256 (N_8256,In_18,In_4338);
nor U8257 (N_8257,In_871,In_3841);
and U8258 (N_8258,In_1794,In_4915);
nand U8259 (N_8259,In_868,In_369);
nand U8260 (N_8260,In_4460,In_2168);
or U8261 (N_8261,In_2791,In_3820);
and U8262 (N_8262,In_4689,In_1147);
and U8263 (N_8263,In_2740,In_4425);
or U8264 (N_8264,In_2893,In_2669);
or U8265 (N_8265,In_676,In_4488);
or U8266 (N_8266,In_3821,In_2778);
or U8267 (N_8267,In_4421,In_1814);
and U8268 (N_8268,In_3525,In_314);
or U8269 (N_8269,In_1918,In_4934);
nor U8270 (N_8270,In_1770,In_922);
and U8271 (N_8271,In_4647,In_543);
or U8272 (N_8272,In_56,In_454);
and U8273 (N_8273,In_1151,In_2546);
nand U8274 (N_8274,In_1282,In_2646);
and U8275 (N_8275,In_4283,In_3659);
xnor U8276 (N_8276,In_2720,In_805);
nor U8277 (N_8277,In_3729,In_4464);
xnor U8278 (N_8278,In_4665,In_3216);
and U8279 (N_8279,In_2767,In_3427);
or U8280 (N_8280,In_2467,In_4564);
or U8281 (N_8281,In_1091,In_2815);
nor U8282 (N_8282,In_4963,In_4953);
nor U8283 (N_8283,In_905,In_2863);
nand U8284 (N_8284,In_4819,In_4665);
or U8285 (N_8285,In_946,In_2120);
nor U8286 (N_8286,In_4250,In_1200);
nand U8287 (N_8287,In_1465,In_4202);
nand U8288 (N_8288,In_2872,In_1082);
xnor U8289 (N_8289,In_498,In_3531);
and U8290 (N_8290,In_3422,In_2892);
or U8291 (N_8291,In_104,In_2783);
nand U8292 (N_8292,In_3726,In_2212);
nor U8293 (N_8293,In_2875,In_1506);
nand U8294 (N_8294,In_629,In_3367);
nand U8295 (N_8295,In_2287,In_2627);
xor U8296 (N_8296,In_994,In_4402);
and U8297 (N_8297,In_652,In_1542);
or U8298 (N_8298,In_3918,In_2574);
nor U8299 (N_8299,In_3909,In_244);
nor U8300 (N_8300,In_2566,In_1163);
and U8301 (N_8301,In_1236,In_3163);
xnor U8302 (N_8302,In_1162,In_4474);
and U8303 (N_8303,In_470,In_4961);
nor U8304 (N_8304,In_2404,In_1931);
or U8305 (N_8305,In_4056,In_4620);
and U8306 (N_8306,In_2503,In_3035);
xnor U8307 (N_8307,In_3548,In_4461);
or U8308 (N_8308,In_4653,In_4812);
xor U8309 (N_8309,In_4888,In_3831);
nand U8310 (N_8310,In_2101,In_3494);
or U8311 (N_8311,In_3715,In_4499);
nor U8312 (N_8312,In_671,In_4961);
or U8313 (N_8313,In_1290,In_1297);
nand U8314 (N_8314,In_1311,In_3894);
and U8315 (N_8315,In_724,In_4702);
nand U8316 (N_8316,In_4633,In_1393);
nor U8317 (N_8317,In_2231,In_590);
xor U8318 (N_8318,In_4226,In_1354);
xnor U8319 (N_8319,In_4951,In_368);
xnor U8320 (N_8320,In_537,In_284);
and U8321 (N_8321,In_1203,In_1146);
xnor U8322 (N_8322,In_1800,In_734);
nor U8323 (N_8323,In_2971,In_4269);
or U8324 (N_8324,In_3662,In_3857);
and U8325 (N_8325,In_563,In_3817);
and U8326 (N_8326,In_3235,In_4974);
and U8327 (N_8327,In_1364,In_574);
nand U8328 (N_8328,In_3699,In_843);
and U8329 (N_8329,In_2,In_1290);
or U8330 (N_8330,In_4460,In_1986);
or U8331 (N_8331,In_275,In_2896);
xor U8332 (N_8332,In_4487,In_1486);
or U8333 (N_8333,In_1052,In_1789);
nor U8334 (N_8334,In_265,In_1241);
and U8335 (N_8335,In_1004,In_1008);
or U8336 (N_8336,In_4881,In_3212);
nor U8337 (N_8337,In_3851,In_3183);
and U8338 (N_8338,In_4021,In_325);
nor U8339 (N_8339,In_3786,In_88);
and U8340 (N_8340,In_4899,In_4344);
nand U8341 (N_8341,In_2782,In_3098);
or U8342 (N_8342,In_2140,In_1128);
nor U8343 (N_8343,In_4865,In_4743);
nor U8344 (N_8344,In_2742,In_1450);
xnor U8345 (N_8345,In_3656,In_3822);
nand U8346 (N_8346,In_4372,In_2876);
xor U8347 (N_8347,In_3270,In_4863);
xnor U8348 (N_8348,In_2421,In_2093);
and U8349 (N_8349,In_2488,In_2755);
nand U8350 (N_8350,In_3835,In_40);
or U8351 (N_8351,In_3551,In_4949);
or U8352 (N_8352,In_3698,In_1462);
or U8353 (N_8353,In_2352,In_1437);
nand U8354 (N_8354,In_3322,In_3426);
and U8355 (N_8355,In_4822,In_186);
or U8356 (N_8356,In_1801,In_125);
nand U8357 (N_8357,In_2682,In_2098);
nand U8358 (N_8358,In_692,In_16);
nand U8359 (N_8359,In_4002,In_2874);
xor U8360 (N_8360,In_4720,In_3227);
xor U8361 (N_8361,In_1587,In_4711);
nand U8362 (N_8362,In_10,In_3358);
or U8363 (N_8363,In_4013,In_871);
nand U8364 (N_8364,In_2648,In_4259);
nand U8365 (N_8365,In_1735,In_354);
xor U8366 (N_8366,In_3299,In_1724);
nand U8367 (N_8367,In_1505,In_2809);
and U8368 (N_8368,In_4775,In_3841);
nand U8369 (N_8369,In_897,In_4024);
nor U8370 (N_8370,In_815,In_1436);
and U8371 (N_8371,In_946,In_2570);
nor U8372 (N_8372,In_1102,In_4225);
and U8373 (N_8373,In_4453,In_4020);
or U8374 (N_8374,In_1481,In_590);
and U8375 (N_8375,In_2715,In_1384);
nand U8376 (N_8376,In_716,In_2799);
or U8377 (N_8377,In_3463,In_1656);
nand U8378 (N_8378,In_1572,In_4741);
or U8379 (N_8379,In_759,In_440);
nor U8380 (N_8380,In_3048,In_2729);
nor U8381 (N_8381,In_3438,In_2758);
xnor U8382 (N_8382,In_3059,In_4282);
nor U8383 (N_8383,In_2384,In_4457);
nand U8384 (N_8384,In_4533,In_1540);
nor U8385 (N_8385,In_921,In_136);
and U8386 (N_8386,In_2742,In_2380);
and U8387 (N_8387,In_2706,In_4599);
xnor U8388 (N_8388,In_4189,In_3599);
nand U8389 (N_8389,In_2154,In_190);
nand U8390 (N_8390,In_4088,In_4316);
nor U8391 (N_8391,In_4330,In_758);
and U8392 (N_8392,In_1416,In_3468);
xor U8393 (N_8393,In_819,In_2610);
nand U8394 (N_8394,In_3264,In_238);
nor U8395 (N_8395,In_3752,In_2102);
or U8396 (N_8396,In_3947,In_1890);
and U8397 (N_8397,In_4668,In_3193);
or U8398 (N_8398,In_4117,In_2217);
or U8399 (N_8399,In_2707,In_2843);
or U8400 (N_8400,In_4208,In_2547);
and U8401 (N_8401,In_3645,In_2715);
nand U8402 (N_8402,In_148,In_4665);
and U8403 (N_8403,In_1117,In_422);
nand U8404 (N_8404,In_3860,In_2151);
nor U8405 (N_8405,In_411,In_1395);
nand U8406 (N_8406,In_3580,In_2295);
or U8407 (N_8407,In_2748,In_3618);
nand U8408 (N_8408,In_1308,In_2313);
nor U8409 (N_8409,In_4357,In_380);
nand U8410 (N_8410,In_939,In_687);
and U8411 (N_8411,In_814,In_635);
nor U8412 (N_8412,In_3415,In_4731);
and U8413 (N_8413,In_1239,In_2229);
xnor U8414 (N_8414,In_3420,In_931);
nand U8415 (N_8415,In_3716,In_1982);
nor U8416 (N_8416,In_3146,In_4568);
nor U8417 (N_8417,In_3541,In_99);
nand U8418 (N_8418,In_861,In_1672);
nand U8419 (N_8419,In_2792,In_4593);
or U8420 (N_8420,In_4768,In_1441);
or U8421 (N_8421,In_3054,In_3506);
nor U8422 (N_8422,In_4423,In_1525);
nand U8423 (N_8423,In_639,In_1215);
nand U8424 (N_8424,In_1505,In_2485);
nor U8425 (N_8425,In_1902,In_846);
nor U8426 (N_8426,In_4230,In_1517);
and U8427 (N_8427,In_3055,In_1114);
nor U8428 (N_8428,In_2261,In_497);
xnor U8429 (N_8429,In_4715,In_2482);
nor U8430 (N_8430,In_2243,In_1965);
or U8431 (N_8431,In_1884,In_4439);
nor U8432 (N_8432,In_804,In_849);
and U8433 (N_8433,In_2874,In_1798);
or U8434 (N_8434,In_140,In_3748);
or U8435 (N_8435,In_1768,In_2366);
and U8436 (N_8436,In_424,In_3966);
nand U8437 (N_8437,In_3847,In_1949);
nor U8438 (N_8438,In_1960,In_118);
nand U8439 (N_8439,In_1666,In_1754);
nor U8440 (N_8440,In_396,In_4672);
or U8441 (N_8441,In_1630,In_2708);
nor U8442 (N_8442,In_394,In_2087);
or U8443 (N_8443,In_3335,In_3664);
and U8444 (N_8444,In_192,In_2359);
nand U8445 (N_8445,In_1168,In_2211);
or U8446 (N_8446,In_1792,In_4283);
nand U8447 (N_8447,In_3251,In_3909);
or U8448 (N_8448,In_800,In_2614);
xnor U8449 (N_8449,In_1306,In_1304);
or U8450 (N_8450,In_735,In_1974);
nor U8451 (N_8451,In_4693,In_4839);
nor U8452 (N_8452,In_403,In_3253);
and U8453 (N_8453,In_4326,In_4878);
and U8454 (N_8454,In_3033,In_4048);
nor U8455 (N_8455,In_912,In_1119);
or U8456 (N_8456,In_3309,In_4363);
and U8457 (N_8457,In_4559,In_3345);
xor U8458 (N_8458,In_3184,In_4173);
xnor U8459 (N_8459,In_233,In_1565);
or U8460 (N_8460,In_2634,In_4972);
xnor U8461 (N_8461,In_539,In_3686);
or U8462 (N_8462,In_1922,In_3747);
or U8463 (N_8463,In_2269,In_2693);
or U8464 (N_8464,In_4044,In_3276);
and U8465 (N_8465,In_2465,In_839);
nand U8466 (N_8466,In_3143,In_1512);
or U8467 (N_8467,In_4081,In_3187);
nand U8468 (N_8468,In_193,In_154);
nand U8469 (N_8469,In_3074,In_2668);
or U8470 (N_8470,In_4529,In_1008);
or U8471 (N_8471,In_958,In_498);
or U8472 (N_8472,In_1247,In_619);
and U8473 (N_8473,In_1433,In_4145);
nand U8474 (N_8474,In_3511,In_1059);
nand U8475 (N_8475,In_1010,In_2187);
nor U8476 (N_8476,In_2058,In_1441);
or U8477 (N_8477,In_1614,In_1409);
nor U8478 (N_8478,In_4040,In_1626);
nand U8479 (N_8479,In_2921,In_3458);
and U8480 (N_8480,In_1947,In_4633);
and U8481 (N_8481,In_2074,In_1648);
nand U8482 (N_8482,In_4957,In_3218);
xnor U8483 (N_8483,In_3067,In_3872);
and U8484 (N_8484,In_3430,In_983);
and U8485 (N_8485,In_2064,In_1125);
and U8486 (N_8486,In_3369,In_2763);
nand U8487 (N_8487,In_4260,In_3628);
nand U8488 (N_8488,In_2388,In_220);
nand U8489 (N_8489,In_2995,In_1243);
xor U8490 (N_8490,In_3954,In_2577);
nand U8491 (N_8491,In_4969,In_1309);
and U8492 (N_8492,In_1578,In_3965);
and U8493 (N_8493,In_3223,In_2348);
nand U8494 (N_8494,In_464,In_2347);
and U8495 (N_8495,In_1612,In_3989);
nand U8496 (N_8496,In_993,In_3762);
nand U8497 (N_8497,In_2271,In_947);
xor U8498 (N_8498,In_2506,In_3896);
and U8499 (N_8499,In_496,In_1673);
and U8500 (N_8500,In_967,In_4511);
nand U8501 (N_8501,In_2572,In_3352);
or U8502 (N_8502,In_1338,In_4035);
nand U8503 (N_8503,In_1990,In_800);
xor U8504 (N_8504,In_921,In_4768);
nor U8505 (N_8505,In_1478,In_1499);
nand U8506 (N_8506,In_347,In_2243);
nor U8507 (N_8507,In_2163,In_205);
nand U8508 (N_8508,In_4223,In_3844);
or U8509 (N_8509,In_506,In_2228);
xnor U8510 (N_8510,In_4310,In_306);
and U8511 (N_8511,In_38,In_897);
or U8512 (N_8512,In_337,In_4380);
and U8513 (N_8513,In_2575,In_411);
nor U8514 (N_8514,In_2593,In_855);
and U8515 (N_8515,In_2016,In_4314);
and U8516 (N_8516,In_4126,In_4838);
and U8517 (N_8517,In_3674,In_3243);
nand U8518 (N_8518,In_4145,In_3317);
and U8519 (N_8519,In_1964,In_3835);
xnor U8520 (N_8520,In_3880,In_4587);
and U8521 (N_8521,In_4208,In_3842);
nor U8522 (N_8522,In_2421,In_2407);
nand U8523 (N_8523,In_3466,In_3507);
or U8524 (N_8524,In_228,In_2702);
nor U8525 (N_8525,In_917,In_4517);
and U8526 (N_8526,In_4743,In_425);
xor U8527 (N_8527,In_3819,In_2401);
or U8528 (N_8528,In_1327,In_3193);
nand U8529 (N_8529,In_2672,In_582);
xnor U8530 (N_8530,In_4642,In_4917);
nor U8531 (N_8531,In_1316,In_3001);
or U8532 (N_8532,In_2553,In_668);
nand U8533 (N_8533,In_2431,In_1405);
nand U8534 (N_8534,In_3331,In_1274);
nor U8535 (N_8535,In_1682,In_3368);
nand U8536 (N_8536,In_1138,In_2367);
and U8537 (N_8537,In_2947,In_744);
nand U8538 (N_8538,In_414,In_1619);
xor U8539 (N_8539,In_278,In_4138);
nand U8540 (N_8540,In_744,In_3499);
and U8541 (N_8541,In_433,In_4606);
and U8542 (N_8542,In_1125,In_3803);
or U8543 (N_8543,In_3204,In_3956);
nor U8544 (N_8544,In_3124,In_2546);
nand U8545 (N_8545,In_380,In_759);
nand U8546 (N_8546,In_4551,In_1156);
and U8547 (N_8547,In_287,In_1603);
and U8548 (N_8548,In_3505,In_1618);
or U8549 (N_8549,In_2189,In_2909);
nor U8550 (N_8550,In_2923,In_1636);
or U8551 (N_8551,In_3174,In_2695);
nor U8552 (N_8552,In_2883,In_2393);
or U8553 (N_8553,In_3267,In_1073);
or U8554 (N_8554,In_3962,In_4396);
nand U8555 (N_8555,In_2164,In_892);
or U8556 (N_8556,In_1426,In_2322);
nand U8557 (N_8557,In_2425,In_2842);
and U8558 (N_8558,In_7,In_1757);
and U8559 (N_8559,In_3039,In_3811);
nor U8560 (N_8560,In_755,In_3718);
or U8561 (N_8561,In_1032,In_791);
nor U8562 (N_8562,In_4437,In_3546);
xor U8563 (N_8563,In_2451,In_1366);
and U8564 (N_8564,In_1082,In_2613);
or U8565 (N_8565,In_3434,In_4770);
nor U8566 (N_8566,In_2895,In_518);
and U8567 (N_8567,In_3947,In_2998);
nor U8568 (N_8568,In_1825,In_1213);
and U8569 (N_8569,In_2662,In_4391);
and U8570 (N_8570,In_3079,In_1072);
and U8571 (N_8571,In_458,In_3981);
nand U8572 (N_8572,In_2890,In_1589);
or U8573 (N_8573,In_4516,In_1169);
or U8574 (N_8574,In_2113,In_172);
and U8575 (N_8575,In_2065,In_4840);
or U8576 (N_8576,In_622,In_3007);
and U8577 (N_8577,In_663,In_3578);
and U8578 (N_8578,In_3560,In_4438);
and U8579 (N_8579,In_4729,In_492);
or U8580 (N_8580,In_1597,In_3668);
nand U8581 (N_8581,In_2962,In_1033);
nand U8582 (N_8582,In_2395,In_626);
xnor U8583 (N_8583,In_3925,In_2210);
or U8584 (N_8584,In_1206,In_3326);
nand U8585 (N_8585,In_44,In_2232);
xor U8586 (N_8586,In_4411,In_1850);
nor U8587 (N_8587,In_4330,In_4725);
and U8588 (N_8588,In_847,In_3285);
and U8589 (N_8589,In_757,In_4382);
or U8590 (N_8590,In_1492,In_439);
and U8591 (N_8591,In_2273,In_3071);
and U8592 (N_8592,In_1897,In_3759);
nor U8593 (N_8593,In_3953,In_479);
and U8594 (N_8594,In_1803,In_4578);
nor U8595 (N_8595,In_971,In_262);
or U8596 (N_8596,In_756,In_1305);
nor U8597 (N_8597,In_4889,In_341);
and U8598 (N_8598,In_1043,In_2442);
and U8599 (N_8599,In_2939,In_1916);
or U8600 (N_8600,In_546,In_1362);
and U8601 (N_8601,In_4936,In_2262);
and U8602 (N_8602,In_65,In_816);
or U8603 (N_8603,In_4401,In_2140);
xnor U8604 (N_8604,In_2861,In_995);
or U8605 (N_8605,In_1164,In_1502);
and U8606 (N_8606,In_341,In_3172);
and U8607 (N_8607,In_2501,In_1783);
nor U8608 (N_8608,In_3262,In_2477);
or U8609 (N_8609,In_2149,In_4641);
nor U8610 (N_8610,In_4645,In_3015);
nor U8611 (N_8611,In_4505,In_706);
or U8612 (N_8612,In_1340,In_2909);
nor U8613 (N_8613,In_4622,In_2014);
nor U8614 (N_8614,In_2168,In_3467);
xnor U8615 (N_8615,In_775,In_2029);
or U8616 (N_8616,In_3387,In_258);
nand U8617 (N_8617,In_4638,In_1907);
and U8618 (N_8618,In_146,In_2400);
or U8619 (N_8619,In_704,In_1761);
or U8620 (N_8620,In_2163,In_478);
or U8621 (N_8621,In_268,In_2060);
nand U8622 (N_8622,In_1832,In_4004);
nor U8623 (N_8623,In_4461,In_1466);
and U8624 (N_8624,In_4681,In_3670);
xnor U8625 (N_8625,In_2731,In_4974);
and U8626 (N_8626,In_4745,In_420);
nor U8627 (N_8627,In_4251,In_3064);
nand U8628 (N_8628,In_1950,In_146);
xnor U8629 (N_8629,In_4801,In_1772);
and U8630 (N_8630,In_866,In_3409);
nor U8631 (N_8631,In_481,In_285);
nor U8632 (N_8632,In_1646,In_4861);
nor U8633 (N_8633,In_1700,In_3770);
or U8634 (N_8634,In_4157,In_2622);
nor U8635 (N_8635,In_732,In_1688);
nor U8636 (N_8636,In_3571,In_1665);
and U8637 (N_8637,In_1139,In_3991);
nor U8638 (N_8638,In_563,In_3896);
nand U8639 (N_8639,In_4113,In_900);
or U8640 (N_8640,In_1842,In_1944);
nand U8641 (N_8641,In_3926,In_3244);
or U8642 (N_8642,In_871,In_3184);
nand U8643 (N_8643,In_737,In_1184);
and U8644 (N_8644,In_2146,In_824);
and U8645 (N_8645,In_2202,In_4690);
nand U8646 (N_8646,In_1016,In_3503);
or U8647 (N_8647,In_4916,In_25);
nand U8648 (N_8648,In_988,In_4975);
or U8649 (N_8649,In_2567,In_714);
nor U8650 (N_8650,In_4583,In_3982);
nand U8651 (N_8651,In_4064,In_7);
nand U8652 (N_8652,In_4504,In_1540);
nor U8653 (N_8653,In_2907,In_1325);
or U8654 (N_8654,In_4050,In_567);
or U8655 (N_8655,In_224,In_3797);
nor U8656 (N_8656,In_3716,In_2604);
or U8657 (N_8657,In_541,In_4905);
xnor U8658 (N_8658,In_4420,In_4731);
nand U8659 (N_8659,In_1177,In_3201);
nor U8660 (N_8660,In_523,In_755);
or U8661 (N_8661,In_948,In_3826);
nor U8662 (N_8662,In_1173,In_1981);
nand U8663 (N_8663,In_4691,In_1702);
and U8664 (N_8664,In_2701,In_3640);
nor U8665 (N_8665,In_2615,In_1912);
nand U8666 (N_8666,In_4318,In_1285);
nor U8667 (N_8667,In_3916,In_2694);
nor U8668 (N_8668,In_1075,In_191);
xnor U8669 (N_8669,In_1072,In_4668);
nand U8670 (N_8670,In_2724,In_4421);
or U8671 (N_8671,In_4295,In_2701);
nor U8672 (N_8672,In_3741,In_2037);
and U8673 (N_8673,In_2337,In_3544);
and U8674 (N_8674,In_2033,In_886);
or U8675 (N_8675,In_1165,In_1753);
nand U8676 (N_8676,In_2087,In_2617);
and U8677 (N_8677,In_330,In_3649);
nand U8678 (N_8678,In_158,In_2710);
xor U8679 (N_8679,In_2355,In_2165);
nand U8680 (N_8680,In_2830,In_1316);
nand U8681 (N_8681,In_141,In_417);
or U8682 (N_8682,In_2307,In_4926);
or U8683 (N_8683,In_2912,In_1872);
nand U8684 (N_8684,In_2777,In_1192);
or U8685 (N_8685,In_1062,In_3111);
nand U8686 (N_8686,In_185,In_628);
xor U8687 (N_8687,In_4862,In_4998);
nor U8688 (N_8688,In_2136,In_2088);
or U8689 (N_8689,In_3229,In_4736);
nand U8690 (N_8690,In_256,In_3320);
nor U8691 (N_8691,In_4462,In_4735);
nand U8692 (N_8692,In_1001,In_931);
or U8693 (N_8693,In_1045,In_3006);
or U8694 (N_8694,In_2591,In_3823);
and U8695 (N_8695,In_91,In_1554);
and U8696 (N_8696,In_2649,In_287);
nor U8697 (N_8697,In_2250,In_2875);
and U8698 (N_8698,In_685,In_4979);
nor U8699 (N_8699,In_2118,In_4684);
or U8700 (N_8700,In_1779,In_4175);
or U8701 (N_8701,In_1398,In_609);
or U8702 (N_8702,In_3098,In_950);
and U8703 (N_8703,In_4602,In_1455);
xor U8704 (N_8704,In_2179,In_3323);
and U8705 (N_8705,In_4395,In_3815);
or U8706 (N_8706,In_4160,In_4570);
and U8707 (N_8707,In_4418,In_2525);
xnor U8708 (N_8708,In_1203,In_3907);
or U8709 (N_8709,In_833,In_2225);
and U8710 (N_8710,In_4067,In_4504);
nor U8711 (N_8711,In_1587,In_2742);
nand U8712 (N_8712,In_2645,In_264);
nor U8713 (N_8713,In_3848,In_2184);
nor U8714 (N_8714,In_1740,In_2218);
nor U8715 (N_8715,In_2674,In_3439);
and U8716 (N_8716,In_2432,In_3625);
nand U8717 (N_8717,In_555,In_4367);
nor U8718 (N_8718,In_812,In_1238);
xnor U8719 (N_8719,In_3099,In_4142);
nand U8720 (N_8720,In_3728,In_202);
nor U8721 (N_8721,In_1687,In_2514);
nor U8722 (N_8722,In_1949,In_1871);
nand U8723 (N_8723,In_4519,In_1339);
and U8724 (N_8724,In_3319,In_3899);
or U8725 (N_8725,In_1826,In_925);
xnor U8726 (N_8726,In_3749,In_1538);
or U8727 (N_8727,In_1151,In_3737);
and U8728 (N_8728,In_3540,In_150);
or U8729 (N_8729,In_3422,In_1064);
nand U8730 (N_8730,In_4503,In_3561);
nand U8731 (N_8731,In_3608,In_1361);
nand U8732 (N_8732,In_3509,In_4682);
or U8733 (N_8733,In_2924,In_4623);
or U8734 (N_8734,In_1701,In_3700);
nor U8735 (N_8735,In_3823,In_4064);
nand U8736 (N_8736,In_3252,In_1562);
nand U8737 (N_8737,In_4930,In_4409);
nand U8738 (N_8738,In_4436,In_4449);
nand U8739 (N_8739,In_355,In_1902);
nand U8740 (N_8740,In_3874,In_2348);
xnor U8741 (N_8741,In_2222,In_940);
nor U8742 (N_8742,In_4292,In_2644);
nand U8743 (N_8743,In_3991,In_1525);
nand U8744 (N_8744,In_1841,In_1767);
and U8745 (N_8745,In_253,In_818);
nor U8746 (N_8746,In_982,In_2202);
and U8747 (N_8747,In_1065,In_3120);
nor U8748 (N_8748,In_1094,In_924);
and U8749 (N_8749,In_3020,In_717);
nor U8750 (N_8750,In_3790,In_4848);
nor U8751 (N_8751,In_3258,In_4001);
nand U8752 (N_8752,In_1703,In_1344);
and U8753 (N_8753,In_1162,In_3458);
and U8754 (N_8754,In_783,In_3131);
nand U8755 (N_8755,In_595,In_1704);
or U8756 (N_8756,In_1133,In_3447);
nor U8757 (N_8757,In_1667,In_3962);
nand U8758 (N_8758,In_916,In_4844);
xnor U8759 (N_8759,In_848,In_2472);
nand U8760 (N_8760,In_2599,In_2488);
and U8761 (N_8761,In_2595,In_1727);
and U8762 (N_8762,In_3674,In_4161);
nand U8763 (N_8763,In_202,In_4700);
and U8764 (N_8764,In_3700,In_1346);
and U8765 (N_8765,In_2664,In_4786);
nand U8766 (N_8766,In_2066,In_3392);
xnor U8767 (N_8767,In_1697,In_2623);
nor U8768 (N_8768,In_3599,In_1406);
nor U8769 (N_8769,In_2011,In_1320);
nand U8770 (N_8770,In_3633,In_1818);
xnor U8771 (N_8771,In_4230,In_1571);
nor U8772 (N_8772,In_4319,In_3802);
and U8773 (N_8773,In_3500,In_269);
and U8774 (N_8774,In_3983,In_496);
or U8775 (N_8775,In_2204,In_4154);
and U8776 (N_8776,In_2354,In_4647);
or U8777 (N_8777,In_3576,In_3255);
and U8778 (N_8778,In_1193,In_4312);
nor U8779 (N_8779,In_609,In_3999);
or U8780 (N_8780,In_3450,In_2467);
nand U8781 (N_8781,In_1536,In_1594);
or U8782 (N_8782,In_4088,In_3379);
and U8783 (N_8783,In_2122,In_3656);
and U8784 (N_8784,In_276,In_2694);
or U8785 (N_8785,In_3244,In_4695);
and U8786 (N_8786,In_4772,In_3479);
nor U8787 (N_8787,In_4821,In_2923);
nor U8788 (N_8788,In_4515,In_4474);
nand U8789 (N_8789,In_4708,In_3776);
or U8790 (N_8790,In_1164,In_1775);
nand U8791 (N_8791,In_2709,In_4048);
nor U8792 (N_8792,In_2179,In_2774);
or U8793 (N_8793,In_2597,In_4297);
nand U8794 (N_8794,In_176,In_4523);
nor U8795 (N_8795,In_2614,In_2548);
nor U8796 (N_8796,In_4037,In_1570);
nor U8797 (N_8797,In_4161,In_964);
and U8798 (N_8798,In_3486,In_1690);
nand U8799 (N_8799,In_4465,In_905);
nor U8800 (N_8800,In_1707,In_1699);
and U8801 (N_8801,In_3232,In_340);
nand U8802 (N_8802,In_4964,In_221);
and U8803 (N_8803,In_14,In_1020);
or U8804 (N_8804,In_355,In_274);
nand U8805 (N_8805,In_4468,In_3892);
nor U8806 (N_8806,In_796,In_4702);
or U8807 (N_8807,In_2137,In_1417);
xor U8808 (N_8808,In_1255,In_2848);
and U8809 (N_8809,In_3333,In_3385);
nor U8810 (N_8810,In_2353,In_3013);
nand U8811 (N_8811,In_2267,In_686);
xor U8812 (N_8812,In_3898,In_3107);
or U8813 (N_8813,In_3382,In_1771);
or U8814 (N_8814,In_1677,In_3849);
and U8815 (N_8815,In_4431,In_265);
nor U8816 (N_8816,In_1397,In_1352);
nor U8817 (N_8817,In_803,In_3332);
and U8818 (N_8818,In_1038,In_2681);
nand U8819 (N_8819,In_3416,In_546);
nor U8820 (N_8820,In_3142,In_1555);
nor U8821 (N_8821,In_1006,In_1811);
nand U8822 (N_8822,In_1483,In_1926);
and U8823 (N_8823,In_3673,In_4346);
or U8824 (N_8824,In_9,In_1149);
and U8825 (N_8825,In_4887,In_3919);
or U8826 (N_8826,In_283,In_854);
and U8827 (N_8827,In_235,In_1260);
nand U8828 (N_8828,In_4320,In_2400);
nand U8829 (N_8829,In_3253,In_3337);
nand U8830 (N_8830,In_3662,In_4620);
nand U8831 (N_8831,In_2468,In_4827);
nand U8832 (N_8832,In_3642,In_3177);
nand U8833 (N_8833,In_2336,In_4657);
or U8834 (N_8834,In_3549,In_2969);
and U8835 (N_8835,In_2251,In_1179);
nand U8836 (N_8836,In_3760,In_1019);
nor U8837 (N_8837,In_110,In_4181);
nor U8838 (N_8838,In_2021,In_2761);
nand U8839 (N_8839,In_4845,In_744);
or U8840 (N_8840,In_3838,In_4848);
nor U8841 (N_8841,In_674,In_414);
nand U8842 (N_8842,In_3276,In_4645);
or U8843 (N_8843,In_3066,In_4152);
nor U8844 (N_8844,In_1176,In_127);
nand U8845 (N_8845,In_2134,In_416);
nand U8846 (N_8846,In_1283,In_530);
nor U8847 (N_8847,In_3224,In_4930);
nand U8848 (N_8848,In_4942,In_801);
or U8849 (N_8849,In_1399,In_3067);
xnor U8850 (N_8850,In_4766,In_4616);
nand U8851 (N_8851,In_4207,In_4932);
nand U8852 (N_8852,In_3770,In_3926);
nand U8853 (N_8853,In_579,In_413);
and U8854 (N_8854,In_1470,In_3490);
nand U8855 (N_8855,In_1097,In_1121);
or U8856 (N_8856,In_1055,In_1001);
nor U8857 (N_8857,In_562,In_1549);
or U8858 (N_8858,In_2079,In_3116);
nand U8859 (N_8859,In_1439,In_3933);
nand U8860 (N_8860,In_2716,In_1271);
nor U8861 (N_8861,In_336,In_3522);
nor U8862 (N_8862,In_2121,In_3123);
nand U8863 (N_8863,In_4174,In_511);
or U8864 (N_8864,In_648,In_3119);
nor U8865 (N_8865,In_796,In_1938);
nand U8866 (N_8866,In_1399,In_3577);
nand U8867 (N_8867,In_2605,In_4552);
nor U8868 (N_8868,In_472,In_407);
and U8869 (N_8869,In_644,In_3871);
and U8870 (N_8870,In_1776,In_1981);
nand U8871 (N_8871,In_984,In_556);
or U8872 (N_8872,In_1757,In_3020);
and U8873 (N_8873,In_530,In_3184);
or U8874 (N_8874,In_2527,In_2421);
xnor U8875 (N_8875,In_105,In_3257);
nor U8876 (N_8876,In_2365,In_1070);
nand U8877 (N_8877,In_2863,In_1776);
and U8878 (N_8878,In_2911,In_3775);
or U8879 (N_8879,In_4132,In_4559);
or U8880 (N_8880,In_3485,In_4940);
or U8881 (N_8881,In_4522,In_4704);
and U8882 (N_8882,In_524,In_1578);
and U8883 (N_8883,In_2088,In_4203);
xor U8884 (N_8884,In_140,In_4255);
xor U8885 (N_8885,In_4657,In_3831);
nor U8886 (N_8886,In_3767,In_4077);
nor U8887 (N_8887,In_1217,In_920);
nor U8888 (N_8888,In_254,In_504);
xor U8889 (N_8889,In_4952,In_2544);
nand U8890 (N_8890,In_1140,In_877);
and U8891 (N_8891,In_597,In_2522);
or U8892 (N_8892,In_1390,In_4291);
or U8893 (N_8893,In_381,In_2611);
and U8894 (N_8894,In_1327,In_2635);
nand U8895 (N_8895,In_987,In_1856);
nand U8896 (N_8896,In_2049,In_4873);
nand U8897 (N_8897,In_3471,In_2627);
nand U8898 (N_8898,In_22,In_3371);
and U8899 (N_8899,In_935,In_4897);
or U8900 (N_8900,In_252,In_1572);
nor U8901 (N_8901,In_3032,In_1424);
or U8902 (N_8902,In_3451,In_25);
or U8903 (N_8903,In_3490,In_4216);
nor U8904 (N_8904,In_133,In_4726);
nand U8905 (N_8905,In_680,In_3412);
nand U8906 (N_8906,In_4424,In_3942);
and U8907 (N_8907,In_2803,In_3651);
and U8908 (N_8908,In_350,In_1914);
nor U8909 (N_8909,In_584,In_4271);
and U8910 (N_8910,In_3677,In_4154);
nand U8911 (N_8911,In_4638,In_3655);
or U8912 (N_8912,In_3577,In_529);
and U8913 (N_8913,In_4006,In_1326);
nand U8914 (N_8914,In_1913,In_4818);
or U8915 (N_8915,In_1923,In_4897);
nand U8916 (N_8916,In_4859,In_3024);
nand U8917 (N_8917,In_3064,In_3155);
nand U8918 (N_8918,In_567,In_4042);
and U8919 (N_8919,In_2103,In_2591);
nor U8920 (N_8920,In_3524,In_209);
and U8921 (N_8921,In_2406,In_338);
and U8922 (N_8922,In_2700,In_1699);
or U8923 (N_8923,In_1061,In_223);
xnor U8924 (N_8924,In_1426,In_4831);
or U8925 (N_8925,In_2783,In_4213);
or U8926 (N_8926,In_966,In_3997);
and U8927 (N_8927,In_4671,In_331);
nor U8928 (N_8928,In_303,In_675);
xnor U8929 (N_8929,In_4026,In_3005);
and U8930 (N_8930,In_694,In_957);
xnor U8931 (N_8931,In_776,In_4610);
nor U8932 (N_8932,In_3525,In_3941);
or U8933 (N_8933,In_15,In_2760);
nand U8934 (N_8934,In_2414,In_4744);
nor U8935 (N_8935,In_4390,In_3191);
nand U8936 (N_8936,In_1902,In_934);
and U8937 (N_8937,In_1712,In_2135);
nor U8938 (N_8938,In_354,In_3281);
nor U8939 (N_8939,In_3178,In_1170);
or U8940 (N_8940,In_516,In_3365);
and U8941 (N_8941,In_1091,In_1824);
nand U8942 (N_8942,In_4154,In_4710);
nor U8943 (N_8943,In_4851,In_3497);
nor U8944 (N_8944,In_1707,In_2813);
nor U8945 (N_8945,In_2028,In_870);
or U8946 (N_8946,In_4215,In_354);
or U8947 (N_8947,In_2487,In_1899);
nand U8948 (N_8948,In_4680,In_1130);
nor U8949 (N_8949,In_1544,In_1064);
or U8950 (N_8950,In_728,In_4512);
or U8951 (N_8951,In_157,In_4442);
or U8952 (N_8952,In_4628,In_4062);
nand U8953 (N_8953,In_4757,In_4505);
xor U8954 (N_8954,In_4867,In_203);
and U8955 (N_8955,In_3990,In_3682);
and U8956 (N_8956,In_4558,In_743);
nor U8957 (N_8957,In_1515,In_471);
and U8958 (N_8958,In_532,In_1811);
and U8959 (N_8959,In_3682,In_457);
and U8960 (N_8960,In_2593,In_484);
nor U8961 (N_8961,In_237,In_3846);
nor U8962 (N_8962,In_4506,In_1242);
nand U8963 (N_8963,In_4891,In_1135);
and U8964 (N_8964,In_2496,In_3552);
and U8965 (N_8965,In_2432,In_2807);
or U8966 (N_8966,In_2768,In_4650);
nand U8967 (N_8967,In_3958,In_562);
nand U8968 (N_8968,In_3256,In_2822);
nor U8969 (N_8969,In_4227,In_992);
or U8970 (N_8970,In_4377,In_602);
and U8971 (N_8971,In_4346,In_1476);
and U8972 (N_8972,In_810,In_1434);
nand U8973 (N_8973,In_4093,In_4046);
nand U8974 (N_8974,In_3890,In_3067);
or U8975 (N_8975,In_399,In_1717);
nand U8976 (N_8976,In_675,In_535);
nor U8977 (N_8977,In_1741,In_3153);
nand U8978 (N_8978,In_1854,In_2986);
nor U8979 (N_8979,In_4937,In_1477);
nand U8980 (N_8980,In_4419,In_4777);
xnor U8981 (N_8981,In_825,In_1512);
nor U8982 (N_8982,In_3929,In_2404);
xnor U8983 (N_8983,In_1920,In_1379);
nor U8984 (N_8984,In_1420,In_4492);
nand U8985 (N_8985,In_3950,In_4460);
or U8986 (N_8986,In_2542,In_1847);
or U8987 (N_8987,In_1252,In_1502);
nor U8988 (N_8988,In_3335,In_4918);
or U8989 (N_8989,In_3180,In_4192);
nand U8990 (N_8990,In_1947,In_3230);
nand U8991 (N_8991,In_4040,In_2068);
nor U8992 (N_8992,In_2432,In_1480);
nor U8993 (N_8993,In_2367,In_2861);
nor U8994 (N_8994,In_3406,In_3369);
nand U8995 (N_8995,In_3495,In_3690);
nand U8996 (N_8996,In_4577,In_3570);
and U8997 (N_8997,In_4750,In_3269);
nand U8998 (N_8998,In_4436,In_2168);
and U8999 (N_8999,In_493,In_4522);
and U9000 (N_9000,In_2373,In_3150);
or U9001 (N_9001,In_2971,In_2530);
or U9002 (N_9002,In_4411,In_4754);
xnor U9003 (N_9003,In_1004,In_3433);
nand U9004 (N_9004,In_4688,In_2664);
nor U9005 (N_9005,In_3166,In_4454);
nor U9006 (N_9006,In_4335,In_3097);
nand U9007 (N_9007,In_4145,In_1671);
nand U9008 (N_9008,In_1335,In_1141);
nor U9009 (N_9009,In_2120,In_4088);
or U9010 (N_9010,In_1413,In_3939);
nand U9011 (N_9011,In_3069,In_142);
or U9012 (N_9012,In_1196,In_3406);
and U9013 (N_9013,In_1185,In_939);
nand U9014 (N_9014,In_1906,In_4712);
nand U9015 (N_9015,In_1978,In_1454);
nor U9016 (N_9016,In_2857,In_870);
nor U9017 (N_9017,In_3435,In_4533);
nand U9018 (N_9018,In_1725,In_782);
nor U9019 (N_9019,In_1347,In_4137);
nand U9020 (N_9020,In_1107,In_15);
and U9021 (N_9021,In_169,In_2870);
and U9022 (N_9022,In_4449,In_3820);
nor U9023 (N_9023,In_734,In_2899);
nand U9024 (N_9024,In_963,In_2194);
nor U9025 (N_9025,In_105,In_2024);
nand U9026 (N_9026,In_2577,In_445);
nand U9027 (N_9027,In_4031,In_3222);
nand U9028 (N_9028,In_982,In_4890);
or U9029 (N_9029,In_2262,In_4889);
and U9030 (N_9030,In_3035,In_4474);
nor U9031 (N_9031,In_1748,In_839);
or U9032 (N_9032,In_1813,In_3457);
or U9033 (N_9033,In_4380,In_446);
nand U9034 (N_9034,In_1592,In_2453);
nor U9035 (N_9035,In_4391,In_2184);
nor U9036 (N_9036,In_3675,In_806);
nor U9037 (N_9037,In_949,In_4610);
nor U9038 (N_9038,In_160,In_1668);
nor U9039 (N_9039,In_4534,In_4630);
and U9040 (N_9040,In_4583,In_2637);
nor U9041 (N_9041,In_1510,In_1944);
or U9042 (N_9042,In_3245,In_2249);
and U9043 (N_9043,In_2901,In_3278);
nor U9044 (N_9044,In_684,In_4887);
nand U9045 (N_9045,In_2530,In_4329);
and U9046 (N_9046,In_3030,In_556);
and U9047 (N_9047,In_3940,In_2300);
and U9048 (N_9048,In_2136,In_1511);
and U9049 (N_9049,In_106,In_1665);
or U9050 (N_9050,In_2441,In_2227);
and U9051 (N_9051,In_2105,In_4899);
nor U9052 (N_9052,In_2525,In_553);
nor U9053 (N_9053,In_211,In_1385);
and U9054 (N_9054,In_4927,In_4254);
nor U9055 (N_9055,In_4671,In_1851);
and U9056 (N_9056,In_4727,In_4379);
nor U9057 (N_9057,In_1688,In_349);
or U9058 (N_9058,In_2462,In_554);
nand U9059 (N_9059,In_2978,In_1828);
and U9060 (N_9060,In_1428,In_556);
nor U9061 (N_9061,In_4302,In_3265);
or U9062 (N_9062,In_1532,In_350);
nor U9063 (N_9063,In_3471,In_748);
xor U9064 (N_9064,In_3031,In_476);
or U9065 (N_9065,In_4905,In_273);
xnor U9066 (N_9066,In_2263,In_1856);
nor U9067 (N_9067,In_35,In_1155);
nor U9068 (N_9068,In_1125,In_4412);
or U9069 (N_9069,In_4302,In_934);
nor U9070 (N_9070,In_4043,In_4826);
nor U9071 (N_9071,In_3824,In_3411);
and U9072 (N_9072,In_3047,In_4051);
nand U9073 (N_9073,In_1274,In_3728);
and U9074 (N_9074,In_933,In_466);
nand U9075 (N_9075,In_4319,In_1612);
and U9076 (N_9076,In_107,In_2009);
and U9077 (N_9077,In_2514,In_3825);
and U9078 (N_9078,In_2647,In_953);
nor U9079 (N_9079,In_539,In_4271);
xnor U9080 (N_9080,In_535,In_3797);
nor U9081 (N_9081,In_2684,In_4680);
xnor U9082 (N_9082,In_3237,In_609);
nand U9083 (N_9083,In_196,In_2068);
or U9084 (N_9084,In_224,In_4538);
nor U9085 (N_9085,In_3558,In_1042);
or U9086 (N_9086,In_3789,In_2649);
nand U9087 (N_9087,In_4859,In_3330);
or U9088 (N_9088,In_133,In_2544);
and U9089 (N_9089,In_2648,In_2784);
nand U9090 (N_9090,In_1833,In_2041);
nor U9091 (N_9091,In_1979,In_2003);
nor U9092 (N_9092,In_2406,In_4587);
nor U9093 (N_9093,In_3901,In_1522);
nor U9094 (N_9094,In_967,In_1346);
nand U9095 (N_9095,In_596,In_4438);
or U9096 (N_9096,In_2627,In_2801);
nor U9097 (N_9097,In_1907,In_65);
nand U9098 (N_9098,In_2474,In_1766);
or U9099 (N_9099,In_1494,In_815);
nor U9100 (N_9100,In_2490,In_3420);
nor U9101 (N_9101,In_4147,In_4621);
or U9102 (N_9102,In_2048,In_4398);
nor U9103 (N_9103,In_4741,In_4242);
nand U9104 (N_9104,In_2634,In_4738);
or U9105 (N_9105,In_896,In_3190);
and U9106 (N_9106,In_1874,In_2438);
nand U9107 (N_9107,In_917,In_1763);
and U9108 (N_9108,In_2381,In_4009);
nor U9109 (N_9109,In_4194,In_3114);
xor U9110 (N_9110,In_1861,In_662);
xor U9111 (N_9111,In_2279,In_2253);
nand U9112 (N_9112,In_3537,In_2731);
nor U9113 (N_9113,In_4471,In_3760);
or U9114 (N_9114,In_2243,In_3669);
and U9115 (N_9115,In_3739,In_4903);
or U9116 (N_9116,In_3895,In_4234);
nor U9117 (N_9117,In_3316,In_525);
nor U9118 (N_9118,In_4333,In_2513);
nand U9119 (N_9119,In_2597,In_4119);
or U9120 (N_9120,In_4305,In_3360);
and U9121 (N_9121,In_4754,In_1217);
or U9122 (N_9122,In_2976,In_620);
or U9123 (N_9123,In_175,In_3607);
nand U9124 (N_9124,In_4570,In_3523);
nor U9125 (N_9125,In_1486,In_513);
nand U9126 (N_9126,In_1031,In_2235);
or U9127 (N_9127,In_1888,In_2887);
or U9128 (N_9128,In_3579,In_2457);
nand U9129 (N_9129,In_723,In_2084);
nand U9130 (N_9130,In_952,In_1180);
nand U9131 (N_9131,In_4055,In_732);
and U9132 (N_9132,In_4860,In_3618);
nand U9133 (N_9133,In_3611,In_4950);
nor U9134 (N_9134,In_4508,In_1817);
and U9135 (N_9135,In_2902,In_3773);
or U9136 (N_9136,In_1190,In_2089);
xor U9137 (N_9137,In_2471,In_3805);
and U9138 (N_9138,In_1802,In_3145);
nor U9139 (N_9139,In_1638,In_2533);
nand U9140 (N_9140,In_3007,In_187);
nand U9141 (N_9141,In_4531,In_1768);
or U9142 (N_9142,In_799,In_1611);
nor U9143 (N_9143,In_1779,In_2677);
xor U9144 (N_9144,In_250,In_3939);
or U9145 (N_9145,In_760,In_1784);
and U9146 (N_9146,In_4277,In_65);
nor U9147 (N_9147,In_4334,In_112);
nand U9148 (N_9148,In_1677,In_486);
nand U9149 (N_9149,In_4094,In_4012);
nor U9150 (N_9150,In_327,In_3237);
nor U9151 (N_9151,In_1858,In_1326);
or U9152 (N_9152,In_2702,In_2640);
and U9153 (N_9153,In_78,In_3193);
or U9154 (N_9154,In_3781,In_1931);
nand U9155 (N_9155,In_3445,In_4418);
nor U9156 (N_9156,In_3470,In_3417);
nor U9157 (N_9157,In_581,In_4920);
and U9158 (N_9158,In_330,In_4592);
xnor U9159 (N_9159,In_234,In_4537);
nand U9160 (N_9160,In_2450,In_3801);
nand U9161 (N_9161,In_184,In_4948);
and U9162 (N_9162,In_2586,In_1425);
or U9163 (N_9163,In_2489,In_3880);
and U9164 (N_9164,In_2608,In_3977);
nand U9165 (N_9165,In_4424,In_1193);
xor U9166 (N_9166,In_2562,In_3505);
or U9167 (N_9167,In_3978,In_4655);
nor U9168 (N_9168,In_4581,In_3239);
nor U9169 (N_9169,In_3509,In_2938);
nor U9170 (N_9170,In_4787,In_1826);
nand U9171 (N_9171,In_4776,In_1557);
or U9172 (N_9172,In_2737,In_1572);
nor U9173 (N_9173,In_4386,In_893);
nor U9174 (N_9174,In_3472,In_4838);
and U9175 (N_9175,In_4573,In_314);
nand U9176 (N_9176,In_4080,In_3970);
or U9177 (N_9177,In_3625,In_3853);
nor U9178 (N_9178,In_4691,In_4078);
nand U9179 (N_9179,In_4771,In_3694);
and U9180 (N_9180,In_3514,In_3360);
or U9181 (N_9181,In_488,In_2529);
nand U9182 (N_9182,In_4583,In_248);
xnor U9183 (N_9183,In_3723,In_416);
nor U9184 (N_9184,In_4445,In_1875);
or U9185 (N_9185,In_851,In_4363);
and U9186 (N_9186,In_2677,In_3884);
and U9187 (N_9187,In_2967,In_3858);
nand U9188 (N_9188,In_3654,In_1211);
or U9189 (N_9189,In_4242,In_3635);
and U9190 (N_9190,In_2748,In_1325);
nand U9191 (N_9191,In_4500,In_2746);
nand U9192 (N_9192,In_745,In_3148);
and U9193 (N_9193,In_3601,In_3585);
and U9194 (N_9194,In_727,In_431);
nor U9195 (N_9195,In_1408,In_2721);
xnor U9196 (N_9196,In_3592,In_1669);
nor U9197 (N_9197,In_818,In_1420);
nor U9198 (N_9198,In_1321,In_4005);
nand U9199 (N_9199,In_2098,In_3918);
nor U9200 (N_9200,In_3735,In_4555);
or U9201 (N_9201,In_1475,In_701);
and U9202 (N_9202,In_2606,In_4939);
nor U9203 (N_9203,In_3172,In_2695);
and U9204 (N_9204,In_1979,In_3982);
nand U9205 (N_9205,In_4263,In_1461);
and U9206 (N_9206,In_3571,In_1299);
or U9207 (N_9207,In_1636,In_3163);
nand U9208 (N_9208,In_4631,In_3471);
and U9209 (N_9209,In_4431,In_4870);
nand U9210 (N_9210,In_3516,In_933);
nand U9211 (N_9211,In_2147,In_4223);
or U9212 (N_9212,In_3291,In_961);
or U9213 (N_9213,In_794,In_265);
xnor U9214 (N_9214,In_4998,In_357);
nand U9215 (N_9215,In_2117,In_1104);
nand U9216 (N_9216,In_3298,In_3554);
nor U9217 (N_9217,In_2129,In_72);
and U9218 (N_9218,In_3576,In_4825);
or U9219 (N_9219,In_1159,In_3913);
nand U9220 (N_9220,In_218,In_3845);
nand U9221 (N_9221,In_389,In_1941);
or U9222 (N_9222,In_1526,In_4719);
and U9223 (N_9223,In_3743,In_573);
and U9224 (N_9224,In_349,In_2922);
nor U9225 (N_9225,In_3732,In_721);
nor U9226 (N_9226,In_106,In_4943);
nor U9227 (N_9227,In_3476,In_2799);
nand U9228 (N_9228,In_3299,In_173);
nor U9229 (N_9229,In_1232,In_3903);
nand U9230 (N_9230,In_2140,In_3037);
nand U9231 (N_9231,In_3158,In_2816);
and U9232 (N_9232,In_1046,In_2174);
and U9233 (N_9233,In_4434,In_3041);
or U9234 (N_9234,In_3462,In_1790);
xnor U9235 (N_9235,In_1432,In_1417);
or U9236 (N_9236,In_3266,In_3651);
and U9237 (N_9237,In_3725,In_431);
and U9238 (N_9238,In_3538,In_4602);
or U9239 (N_9239,In_465,In_756);
or U9240 (N_9240,In_2362,In_3717);
nand U9241 (N_9241,In_3588,In_4609);
and U9242 (N_9242,In_4708,In_2802);
and U9243 (N_9243,In_92,In_3072);
nor U9244 (N_9244,In_3710,In_2848);
or U9245 (N_9245,In_1044,In_2247);
and U9246 (N_9246,In_1204,In_732);
and U9247 (N_9247,In_4319,In_4017);
nand U9248 (N_9248,In_2550,In_240);
nand U9249 (N_9249,In_4633,In_1967);
and U9250 (N_9250,In_872,In_1365);
nand U9251 (N_9251,In_1965,In_3291);
nor U9252 (N_9252,In_3280,In_1446);
and U9253 (N_9253,In_4996,In_4461);
and U9254 (N_9254,In_746,In_3503);
or U9255 (N_9255,In_282,In_2040);
nor U9256 (N_9256,In_4783,In_2248);
or U9257 (N_9257,In_319,In_3555);
or U9258 (N_9258,In_4346,In_3402);
or U9259 (N_9259,In_1114,In_2361);
and U9260 (N_9260,In_4091,In_4241);
and U9261 (N_9261,In_3549,In_711);
nor U9262 (N_9262,In_364,In_919);
or U9263 (N_9263,In_1453,In_1151);
or U9264 (N_9264,In_4051,In_2999);
or U9265 (N_9265,In_3239,In_2553);
nand U9266 (N_9266,In_470,In_3338);
nand U9267 (N_9267,In_4301,In_3644);
and U9268 (N_9268,In_891,In_154);
nor U9269 (N_9269,In_4496,In_960);
nor U9270 (N_9270,In_4512,In_2949);
nand U9271 (N_9271,In_3805,In_3147);
and U9272 (N_9272,In_57,In_4023);
or U9273 (N_9273,In_34,In_3195);
nand U9274 (N_9274,In_4026,In_3446);
nand U9275 (N_9275,In_941,In_4476);
nor U9276 (N_9276,In_793,In_4491);
or U9277 (N_9277,In_2851,In_2110);
nor U9278 (N_9278,In_363,In_3607);
nor U9279 (N_9279,In_410,In_2774);
and U9280 (N_9280,In_2659,In_395);
and U9281 (N_9281,In_362,In_1994);
and U9282 (N_9282,In_2107,In_1825);
nand U9283 (N_9283,In_2351,In_400);
nand U9284 (N_9284,In_1323,In_3048);
or U9285 (N_9285,In_3887,In_525);
nor U9286 (N_9286,In_4020,In_2663);
nor U9287 (N_9287,In_1220,In_4704);
nand U9288 (N_9288,In_801,In_1533);
or U9289 (N_9289,In_3422,In_2636);
nor U9290 (N_9290,In_4796,In_2766);
nor U9291 (N_9291,In_1695,In_2395);
and U9292 (N_9292,In_4509,In_3791);
and U9293 (N_9293,In_1444,In_1578);
and U9294 (N_9294,In_220,In_4493);
nand U9295 (N_9295,In_1080,In_4888);
nand U9296 (N_9296,In_2669,In_2558);
xnor U9297 (N_9297,In_4034,In_2415);
or U9298 (N_9298,In_3283,In_3620);
nor U9299 (N_9299,In_1369,In_1715);
nor U9300 (N_9300,In_577,In_2335);
xor U9301 (N_9301,In_3787,In_3503);
nor U9302 (N_9302,In_703,In_4754);
nor U9303 (N_9303,In_1391,In_3573);
or U9304 (N_9304,In_2217,In_3258);
and U9305 (N_9305,In_4870,In_1574);
nand U9306 (N_9306,In_1993,In_2612);
and U9307 (N_9307,In_1395,In_602);
nand U9308 (N_9308,In_352,In_4758);
or U9309 (N_9309,In_3406,In_2852);
nor U9310 (N_9310,In_4913,In_114);
xor U9311 (N_9311,In_1274,In_3007);
nand U9312 (N_9312,In_2576,In_4310);
nor U9313 (N_9313,In_2027,In_171);
or U9314 (N_9314,In_2613,In_4206);
or U9315 (N_9315,In_4720,In_4113);
xnor U9316 (N_9316,In_4207,In_3155);
nand U9317 (N_9317,In_4225,In_1251);
nand U9318 (N_9318,In_1392,In_183);
and U9319 (N_9319,In_1439,In_215);
nor U9320 (N_9320,In_3861,In_2010);
xnor U9321 (N_9321,In_3768,In_1068);
nor U9322 (N_9322,In_2905,In_3481);
nor U9323 (N_9323,In_4042,In_4741);
xor U9324 (N_9324,In_3000,In_2976);
and U9325 (N_9325,In_4726,In_2402);
and U9326 (N_9326,In_4792,In_3718);
and U9327 (N_9327,In_2104,In_3020);
nand U9328 (N_9328,In_3330,In_1339);
or U9329 (N_9329,In_1671,In_4099);
xnor U9330 (N_9330,In_2152,In_3625);
or U9331 (N_9331,In_1543,In_1152);
and U9332 (N_9332,In_2929,In_1363);
nor U9333 (N_9333,In_2247,In_4565);
nor U9334 (N_9334,In_4887,In_485);
nand U9335 (N_9335,In_3809,In_3579);
or U9336 (N_9336,In_2351,In_4963);
and U9337 (N_9337,In_3676,In_2360);
or U9338 (N_9338,In_3643,In_381);
nand U9339 (N_9339,In_4464,In_2810);
and U9340 (N_9340,In_446,In_1183);
nand U9341 (N_9341,In_3171,In_195);
nor U9342 (N_9342,In_1795,In_681);
and U9343 (N_9343,In_3998,In_136);
and U9344 (N_9344,In_428,In_3023);
nor U9345 (N_9345,In_2473,In_98);
nor U9346 (N_9346,In_930,In_4174);
or U9347 (N_9347,In_4713,In_4534);
or U9348 (N_9348,In_4687,In_1734);
or U9349 (N_9349,In_1808,In_2094);
nand U9350 (N_9350,In_793,In_2747);
nor U9351 (N_9351,In_3838,In_397);
nand U9352 (N_9352,In_4423,In_4823);
xnor U9353 (N_9353,In_2497,In_1837);
or U9354 (N_9354,In_2291,In_2213);
and U9355 (N_9355,In_647,In_4994);
or U9356 (N_9356,In_3226,In_3805);
nor U9357 (N_9357,In_3530,In_1643);
xor U9358 (N_9358,In_2201,In_3315);
and U9359 (N_9359,In_1798,In_4292);
xor U9360 (N_9360,In_3321,In_1674);
nor U9361 (N_9361,In_15,In_4974);
xor U9362 (N_9362,In_3253,In_3940);
nand U9363 (N_9363,In_956,In_1581);
nand U9364 (N_9364,In_3814,In_793);
or U9365 (N_9365,In_2281,In_2827);
or U9366 (N_9366,In_3790,In_2363);
and U9367 (N_9367,In_2052,In_167);
nor U9368 (N_9368,In_569,In_371);
and U9369 (N_9369,In_2039,In_1651);
and U9370 (N_9370,In_3568,In_904);
or U9371 (N_9371,In_3331,In_3813);
nor U9372 (N_9372,In_4967,In_4670);
or U9373 (N_9373,In_2553,In_2677);
nor U9374 (N_9374,In_1396,In_3144);
nand U9375 (N_9375,In_3821,In_2091);
or U9376 (N_9376,In_3097,In_2308);
xor U9377 (N_9377,In_3552,In_4360);
nand U9378 (N_9378,In_3644,In_4017);
nor U9379 (N_9379,In_2543,In_2921);
xnor U9380 (N_9380,In_1032,In_3508);
nor U9381 (N_9381,In_3384,In_2422);
nor U9382 (N_9382,In_2870,In_296);
nand U9383 (N_9383,In_3654,In_826);
nand U9384 (N_9384,In_3134,In_1610);
or U9385 (N_9385,In_3519,In_556);
nand U9386 (N_9386,In_2924,In_4911);
or U9387 (N_9387,In_4740,In_760);
and U9388 (N_9388,In_4168,In_3284);
and U9389 (N_9389,In_794,In_226);
nand U9390 (N_9390,In_1808,In_4959);
nor U9391 (N_9391,In_2868,In_2856);
nor U9392 (N_9392,In_2733,In_3620);
xor U9393 (N_9393,In_2146,In_4987);
nand U9394 (N_9394,In_4323,In_1334);
nor U9395 (N_9395,In_3088,In_3890);
nor U9396 (N_9396,In_1431,In_3984);
nand U9397 (N_9397,In_3999,In_4295);
or U9398 (N_9398,In_1697,In_1964);
nand U9399 (N_9399,In_766,In_982);
nor U9400 (N_9400,In_397,In_2684);
or U9401 (N_9401,In_4625,In_1521);
nand U9402 (N_9402,In_425,In_2829);
nor U9403 (N_9403,In_43,In_1227);
nor U9404 (N_9404,In_3050,In_3744);
and U9405 (N_9405,In_584,In_4696);
nor U9406 (N_9406,In_3123,In_2368);
and U9407 (N_9407,In_4441,In_2606);
and U9408 (N_9408,In_4062,In_279);
nor U9409 (N_9409,In_2051,In_938);
and U9410 (N_9410,In_2970,In_354);
or U9411 (N_9411,In_2962,In_808);
and U9412 (N_9412,In_3990,In_1753);
or U9413 (N_9413,In_3450,In_669);
and U9414 (N_9414,In_4645,In_4482);
nand U9415 (N_9415,In_4826,In_696);
and U9416 (N_9416,In_3733,In_3200);
nand U9417 (N_9417,In_1348,In_335);
nand U9418 (N_9418,In_1265,In_2102);
nand U9419 (N_9419,In_3355,In_4455);
nor U9420 (N_9420,In_1429,In_3995);
nor U9421 (N_9421,In_214,In_132);
nand U9422 (N_9422,In_3159,In_937);
nor U9423 (N_9423,In_1203,In_4805);
and U9424 (N_9424,In_3968,In_1695);
nand U9425 (N_9425,In_4470,In_4095);
nand U9426 (N_9426,In_1473,In_3790);
or U9427 (N_9427,In_3855,In_944);
and U9428 (N_9428,In_1774,In_3036);
or U9429 (N_9429,In_4601,In_4103);
xor U9430 (N_9430,In_4777,In_420);
and U9431 (N_9431,In_4689,In_2126);
nor U9432 (N_9432,In_2388,In_4919);
or U9433 (N_9433,In_3462,In_3170);
or U9434 (N_9434,In_1698,In_1482);
nand U9435 (N_9435,In_4780,In_3272);
and U9436 (N_9436,In_3815,In_4884);
nand U9437 (N_9437,In_3164,In_881);
and U9438 (N_9438,In_4817,In_4674);
nor U9439 (N_9439,In_740,In_2313);
nor U9440 (N_9440,In_3810,In_2275);
nor U9441 (N_9441,In_3535,In_2809);
and U9442 (N_9442,In_3179,In_4566);
xnor U9443 (N_9443,In_3881,In_3248);
and U9444 (N_9444,In_3867,In_661);
nand U9445 (N_9445,In_3243,In_3659);
or U9446 (N_9446,In_2811,In_3346);
and U9447 (N_9447,In_2806,In_3583);
nor U9448 (N_9448,In_3286,In_273);
nand U9449 (N_9449,In_4227,In_426);
and U9450 (N_9450,In_880,In_1171);
nand U9451 (N_9451,In_3828,In_4922);
xor U9452 (N_9452,In_1907,In_3799);
or U9453 (N_9453,In_945,In_2534);
xor U9454 (N_9454,In_600,In_3694);
or U9455 (N_9455,In_111,In_1103);
xor U9456 (N_9456,In_587,In_1066);
or U9457 (N_9457,In_929,In_3661);
or U9458 (N_9458,In_4216,In_1043);
xnor U9459 (N_9459,In_4179,In_814);
or U9460 (N_9460,In_229,In_1927);
nor U9461 (N_9461,In_4698,In_1692);
xor U9462 (N_9462,In_1154,In_2253);
nand U9463 (N_9463,In_1643,In_2678);
nor U9464 (N_9464,In_1241,In_4094);
nor U9465 (N_9465,In_1779,In_4851);
and U9466 (N_9466,In_4958,In_2749);
nand U9467 (N_9467,In_880,In_1504);
nand U9468 (N_9468,In_4793,In_3350);
xnor U9469 (N_9469,In_4125,In_818);
or U9470 (N_9470,In_3089,In_1047);
nor U9471 (N_9471,In_532,In_7);
nor U9472 (N_9472,In_1487,In_4468);
and U9473 (N_9473,In_826,In_728);
nor U9474 (N_9474,In_1804,In_230);
nor U9475 (N_9475,In_3208,In_39);
nand U9476 (N_9476,In_210,In_880);
and U9477 (N_9477,In_1638,In_4967);
nor U9478 (N_9478,In_1276,In_4858);
nand U9479 (N_9479,In_1608,In_4839);
nand U9480 (N_9480,In_2779,In_1553);
nand U9481 (N_9481,In_757,In_3915);
nand U9482 (N_9482,In_1790,In_1539);
nand U9483 (N_9483,In_4937,In_4704);
nor U9484 (N_9484,In_3444,In_4345);
xnor U9485 (N_9485,In_2882,In_911);
nand U9486 (N_9486,In_582,In_2361);
and U9487 (N_9487,In_1776,In_788);
nor U9488 (N_9488,In_4923,In_1160);
or U9489 (N_9489,In_4089,In_4348);
or U9490 (N_9490,In_2218,In_4464);
nand U9491 (N_9491,In_4191,In_4258);
nor U9492 (N_9492,In_4950,In_1949);
and U9493 (N_9493,In_63,In_1235);
and U9494 (N_9494,In_1815,In_3848);
nor U9495 (N_9495,In_1992,In_1505);
nor U9496 (N_9496,In_2632,In_1053);
or U9497 (N_9497,In_691,In_4037);
or U9498 (N_9498,In_1630,In_1169);
and U9499 (N_9499,In_764,In_4854);
nor U9500 (N_9500,In_3694,In_532);
or U9501 (N_9501,In_3908,In_548);
nand U9502 (N_9502,In_2104,In_4446);
and U9503 (N_9503,In_2357,In_1703);
or U9504 (N_9504,In_270,In_2655);
and U9505 (N_9505,In_1533,In_908);
nor U9506 (N_9506,In_652,In_1199);
nor U9507 (N_9507,In_1346,In_2181);
or U9508 (N_9508,In_1141,In_4875);
nand U9509 (N_9509,In_2838,In_2495);
and U9510 (N_9510,In_614,In_2632);
nand U9511 (N_9511,In_3887,In_4670);
xor U9512 (N_9512,In_4741,In_1496);
xnor U9513 (N_9513,In_4144,In_1913);
and U9514 (N_9514,In_3635,In_390);
or U9515 (N_9515,In_494,In_4890);
nand U9516 (N_9516,In_3168,In_4413);
xor U9517 (N_9517,In_735,In_3170);
and U9518 (N_9518,In_4007,In_1259);
nand U9519 (N_9519,In_1606,In_2746);
nand U9520 (N_9520,In_1537,In_2988);
nor U9521 (N_9521,In_3048,In_4789);
nor U9522 (N_9522,In_4989,In_640);
nor U9523 (N_9523,In_17,In_3999);
or U9524 (N_9524,In_240,In_4791);
and U9525 (N_9525,In_574,In_3232);
nand U9526 (N_9526,In_1264,In_4813);
nor U9527 (N_9527,In_443,In_675);
or U9528 (N_9528,In_2314,In_3642);
or U9529 (N_9529,In_4592,In_1488);
or U9530 (N_9530,In_269,In_1659);
or U9531 (N_9531,In_3642,In_4653);
nand U9532 (N_9532,In_230,In_582);
nand U9533 (N_9533,In_3712,In_2802);
nand U9534 (N_9534,In_1827,In_3859);
or U9535 (N_9535,In_2207,In_3421);
xnor U9536 (N_9536,In_1486,In_4971);
or U9537 (N_9537,In_4513,In_4799);
and U9538 (N_9538,In_3340,In_292);
and U9539 (N_9539,In_770,In_3976);
or U9540 (N_9540,In_2894,In_3013);
or U9541 (N_9541,In_2722,In_2143);
xnor U9542 (N_9542,In_3090,In_1411);
or U9543 (N_9543,In_2885,In_251);
or U9544 (N_9544,In_855,In_3390);
nand U9545 (N_9545,In_2803,In_1887);
nand U9546 (N_9546,In_4327,In_3548);
nor U9547 (N_9547,In_950,In_4720);
nand U9548 (N_9548,In_808,In_2434);
and U9549 (N_9549,In_3182,In_68);
or U9550 (N_9550,In_3730,In_4461);
and U9551 (N_9551,In_1003,In_383);
nor U9552 (N_9552,In_4074,In_3173);
and U9553 (N_9553,In_4974,In_2542);
xor U9554 (N_9554,In_1326,In_1527);
nand U9555 (N_9555,In_1687,In_3444);
xnor U9556 (N_9556,In_3941,In_4345);
and U9557 (N_9557,In_1830,In_1470);
xor U9558 (N_9558,In_4825,In_3764);
nor U9559 (N_9559,In_4307,In_4739);
and U9560 (N_9560,In_3498,In_2764);
xnor U9561 (N_9561,In_4928,In_902);
nand U9562 (N_9562,In_1866,In_3100);
and U9563 (N_9563,In_1492,In_2914);
or U9564 (N_9564,In_1471,In_1705);
and U9565 (N_9565,In_459,In_1423);
and U9566 (N_9566,In_4443,In_1171);
and U9567 (N_9567,In_3886,In_4207);
or U9568 (N_9568,In_2721,In_832);
nor U9569 (N_9569,In_2634,In_1939);
and U9570 (N_9570,In_4074,In_2785);
or U9571 (N_9571,In_4726,In_1319);
or U9572 (N_9572,In_1518,In_1422);
nand U9573 (N_9573,In_1401,In_2673);
and U9574 (N_9574,In_3615,In_1519);
and U9575 (N_9575,In_3862,In_3278);
and U9576 (N_9576,In_2096,In_1327);
or U9577 (N_9577,In_4957,In_4400);
or U9578 (N_9578,In_3132,In_4690);
or U9579 (N_9579,In_4303,In_4793);
or U9580 (N_9580,In_4046,In_4370);
xnor U9581 (N_9581,In_2708,In_1298);
nand U9582 (N_9582,In_3974,In_1082);
xnor U9583 (N_9583,In_3147,In_64);
nor U9584 (N_9584,In_2577,In_2941);
and U9585 (N_9585,In_3676,In_3318);
and U9586 (N_9586,In_409,In_441);
and U9587 (N_9587,In_845,In_3664);
and U9588 (N_9588,In_2202,In_3759);
or U9589 (N_9589,In_4328,In_680);
or U9590 (N_9590,In_2254,In_2883);
or U9591 (N_9591,In_3835,In_773);
nand U9592 (N_9592,In_3943,In_4060);
nand U9593 (N_9593,In_736,In_1769);
nor U9594 (N_9594,In_2840,In_4224);
nor U9595 (N_9595,In_4153,In_3659);
or U9596 (N_9596,In_3030,In_2223);
nand U9597 (N_9597,In_4984,In_4803);
nand U9598 (N_9598,In_2318,In_3506);
nand U9599 (N_9599,In_3130,In_4677);
and U9600 (N_9600,In_2768,In_1385);
xnor U9601 (N_9601,In_1923,In_3625);
xnor U9602 (N_9602,In_4355,In_4698);
nand U9603 (N_9603,In_2556,In_3459);
nor U9604 (N_9604,In_2228,In_2416);
and U9605 (N_9605,In_4952,In_531);
nor U9606 (N_9606,In_4753,In_3000);
and U9607 (N_9607,In_147,In_4542);
or U9608 (N_9608,In_4542,In_1005);
xnor U9609 (N_9609,In_576,In_2998);
nand U9610 (N_9610,In_2902,In_1237);
or U9611 (N_9611,In_4622,In_4029);
nor U9612 (N_9612,In_1122,In_2731);
xnor U9613 (N_9613,In_3654,In_2110);
and U9614 (N_9614,In_1671,In_3122);
nand U9615 (N_9615,In_1287,In_836);
nand U9616 (N_9616,In_606,In_3928);
or U9617 (N_9617,In_4708,In_1492);
nand U9618 (N_9618,In_773,In_3431);
xor U9619 (N_9619,In_40,In_1391);
nand U9620 (N_9620,In_1992,In_69);
or U9621 (N_9621,In_3110,In_4242);
and U9622 (N_9622,In_4443,In_3570);
nor U9623 (N_9623,In_1111,In_671);
nor U9624 (N_9624,In_919,In_303);
or U9625 (N_9625,In_1734,In_4516);
nand U9626 (N_9626,In_472,In_4977);
xor U9627 (N_9627,In_3423,In_3800);
xnor U9628 (N_9628,In_3498,In_3570);
nor U9629 (N_9629,In_2905,In_3686);
or U9630 (N_9630,In_2681,In_4688);
or U9631 (N_9631,In_1603,In_46);
or U9632 (N_9632,In_3297,In_3545);
and U9633 (N_9633,In_4120,In_905);
nor U9634 (N_9634,In_263,In_837);
nor U9635 (N_9635,In_2508,In_2563);
or U9636 (N_9636,In_4960,In_4765);
or U9637 (N_9637,In_1687,In_2556);
nor U9638 (N_9638,In_154,In_1449);
and U9639 (N_9639,In_3465,In_1757);
nand U9640 (N_9640,In_3701,In_3304);
or U9641 (N_9641,In_2083,In_2973);
or U9642 (N_9642,In_3086,In_47);
nand U9643 (N_9643,In_2209,In_2924);
and U9644 (N_9644,In_3003,In_831);
and U9645 (N_9645,In_4378,In_2162);
nand U9646 (N_9646,In_1096,In_345);
nor U9647 (N_9647,In_2031,In_2512);
nand U9648 (N_9648,In_2091,In_2395);
nor U9649 (N_9649,In_1434,In_4410);
nor U9650 (N_9650,In_2181,In_108);
or U9651 (N_9651,In_473,In_1785);
nand U9652 (N_9652,In_2233,In_764);
nor U9653 (N_9653,In_1356,In_4290);
xnor U9654 (N_9654,In_2455,In_1524);
xnor U9655 (N_9655,In_1593,In_4133);
xnor U9656 (N_9656,In_562,In_1498);
nand U9657 (N_9657,In_1028,In_4700);
or U9658 (N_9658,In_2866,In_3833);
and U9659 (N_9659,In_694,In_955);
nor U9660 (N_9660,In_2433,In_884);
nand U9661 (N_9661,In_3244,In_3590);
nand U9662 (N_9662,In_1546,In_1541);
or U9663 (N_9663,In_371,In_252);
nand U9664 (N_9664,In_3962,In_4129);
xnor U9665 (N_9665,In_3541,In_4065);
nor U9666 (N_9666,In_1515,In_4363);
and U9667 (N_9667,In_1817,In_4603);
nor U9668 (N_9668,In_3734,In_3984);
and U9669 (N_9669,In_4757,In_1171);
or U9670 (N_9670,In_3388,In_3829);
nor U9671 (N_9671,In_454,In_585);
and U9672 (N_9672,In_4370,In_1149);
nand U9673 (N_9673,In_3254,In_4587);
nand U9674 (N_9674,In_3389,In_4392);
nand U9675 (N_9675,In_4238,In_3182);
nor U9676 (N_9676,In_2815,In_1502);
xnor U9677 (N_9677,In_4750,In_1139);
nand U9678 (N_9678,In_4542,In_321);
nor U9679 (N_9679,In_1967,In_4760);
or U9680 (N_9680,In_131,In_2692);
or U9681 (N_9681,In_760,In_4988);
and U9682 (N_9682,In_1864,In_3246);
or U9683 (N_9683,In_2472,In_4804);
and U9684 (N_9684,In_2302,In_4713);
nor U9685 (N_9685,In_4211,In_1698);
nor U9686 (N_9686,In_40,In_1902);
and U9687 (N_9687,In_4655,In_4737);
nand U9688 (N_9688,In_694,In_2667);
or U9689 (N_9689,In_1154,In_4969);
nor U9690 (N_9690,In_1247,In_3696);
nor U9691 (N_9691,In_4654,In_4803);
or U9692 (N_9692,In_951,In_2039);
nor U9693 (N_9693,In_4333,In_3568);
nand U9694 (N_9694,In_2385,In_850);
xnor U9695 (N_9695,In_828,In_2790);
or U9696 (N_9696,In_2579,In_2006);
nand U9697 (N_9697,In_4034,In_126);
and U9698 (N_9698,In_4395,In_1163);
nand U9699 (N_9699,In_2751,In_2528);
or U9700 (N_9700,In_1599,In_1690);
and U9701 (N_9701,In_2382,In_2706);
or U9702 (N_9702,In_369,In_2938);
nor U9703 (N_9703,In_4440,In_1435);
nand U9704 (N_9704,In_2865,In_4865);
xnor U9705 (N_9705,In_1319,In_3101);
and U9706 (N_9706,In_2707,In_983);
nor U9707 (N_9707,In_1014,In_3253);
nand U9708 (N_9708,In_1581,In_3526);
and U9709 (N_9709,In_3438,In_3856);
and U9710 (N_9710,In_1503,In_1448);
nand U9711 (N_9711,In_1160,In_4228);
nand U9712 (N_9712,In_2217,In_4137);
xor U9713 (N_9713,In_2227,In_3830);
or U9714 (N_9714,In_4703,In_4273);
nand U9715 (N_9715,In_207,In_473);
nand U9716 (N_9716,In_4683,In_4150);
nand U9717 (N_9717,In_4570,In_2550);
nand U9718 (N_9718,In_4103,In_2165);
nor U9719 (N_9719,In_4242,In_405);
nand U9720 (N_9720,In_3882,In_3341);
or U9721 (N_9721,In_3628,In_224);
or U9722 (N_9722,In_4626,In_3866);
or U9723 (N_9723,In_123,In_726);
nand U9724 (N_9724,In_4962,In_3883);
or U9725 (N_9725,In_3336,In_3153);
nor U9726 (N_9726,In_4905,In_3372);
nor U9727 (N_9727,In_927,In_4272);
nand U9728 (N_9728,In_1460,In_3096);
and U9729 (N_9729,In_4264,In_1698);
nor U9730 (N_9730,In_3169,In_4734);
or U9731 (N_9731,In_2780,In_617);
nor U9732 (N_9732,In_636,In_4641);
and U9733 (N_9733,In_2308,In_4602);
xor U9734 (N_9734,In_2108,In_3290);
and U9735 (N_9735,In_3841,In_2588);
xnor U9736 (N_9736,In_2877,In_1144);
nor U9737 (N_9737,In_4209,In_2663);
and U9738 (N_9738,In_1349,In_2850);
or U9739 (N_9739,In_3141,In_330);
nor U9740 (N_9740,In_4478,In_4855);
or U9741 (N_9741,In_1044,In_2275);
and U9742 (N_9742,In_4838,In_522);
nor U9743 (N_9743,In_1663,In_776);
nor U9744 (N_9744,In_2933,In_2903);
or U9745 (N_9745,In_4366,In_2448);
and U9746 (N_9746,In_3757,In_4199);
and U9747 (N_9747,In_4913,In_1498);
and U9748 (N_9748,In_28,In_4518);
or U9749 (N_9749,In_2767,In_395);
xor U9750 (N_9750,In_447,In_1436);
and U9751 (N_9751,In_3379,In_817);
and U9752 (N_9752,In_1245,In_4968);
nand U9753 (N_9753,In_3366,In_4780);
and U9754 (N_9754,In_3375,In_4053);
and U9755 (N_9755,In_698,In_3289);
xor U9756 (N_9756,In_3702,In_1591);
or U9757 (N_9757,In_904,In_847);
or U9758 (N_9758,In_3327,In_4484);
or U9759 (N_9759,In_3229,In_805);
nor U9760 (N_9760,In_1158,In_4326);
or U9761 (N_9761,In_3314,In_3698);
or U9762 (N_9762,In_3358,In_1538);
nand U9763 (N_9763,In_2893,In_4438);
nor U9764 (N_9764,In_3065,In_2365);
nand U9765 (N_9765,In_1263,In_1608);
or U9766 (N_9766,In_2032,In_3355);
nor U9767 (N_9767,In_4419,In_3641);
nand U9768 (N_9768,In_489,In_873);
nand U9769 (N_9769,In_4400,In_2936);
xor U9770 (N_9770,In_2844,In_4863);
nand U9771 (N_9771,In_2974,In_2424);
and U9772 (N_9772,In_4713,In_1307);
and U9773 (N_9773,In_64,In_2896);
nor U9774 (N_9774,In_4926,In_3296);
xor U9775 (N_9775,In_1566,In_2702);
nand U9776 (N_9776,In_3396,In_3467);
or U9777 (N_9777,In_169,In_4798);
xor U9778 (N_9778,In_3866,In_2660);
xnor U9779 (N_9779,In_3508,In_2291);
nor U9780 (N_9780,In_1883,In_2036);
and U9781 (N_9781,In_3626,In_2021);
nand U9782 (N_9782,In_517,In_295);
or U9783 (N_9783,In_3879,In_3488);
and U9784 (N_9784,In_3519,In_1018);
or U9785 (N_9785,In_3160,In_1208);
and U9786 (N_9786,In_2450,In_1107);
nand U9787 (N_9787,In_667,In_3774);
nand U9788 (N_9788,In_4972,In_389);
nand U9789 (N_9789,In_1385,In_4375);
or U9790 (N_9790,In_3838,In_601);
nand U9791 (N_9791,In_766,In_754);
nor U9792 (N_9792,In_1696,In_4579);
xor U9793 (N_9793,In_3246,In_1967);
and U9794 (N_9794,In_563,In_3361);
xnor U9795 (N_9795,In_1067,In_4113);
nor U9796 (N_9796,In_4779,In_4337);
or U9797 (N_9797,In_2982,In_4352);
and U9798 (N_9798,In_890,In_3882);
nor U9799 (N_9799,In_2591,In_3427);
nor U9800 (N_9800,In_2545,In_1113);
or U9801 (N_9801,In_4245,In_2892);
nor U9802 (N_9802,In_3219,In_2370);
or U9803 (N_9803,In_4888,In_1055);
nand U9804 (N_9804,In_2440,In_823);
and U9805 (N_9805,In_1521,In_4066);
nand U9806 (N_9806,In_3530,In_1298);
and U9807 (N_9807,In_1189,In_1944);
nor U9808 (N_9808,In_2868,In_57);
and U9809 (N_9809,In_25,In_3101);
or U9810 (N_9810,In_4107,In_1568);
or U9811 (N_9811,In_2980,In_3280);
nor U9812 (N_9812,In_1634,In_1518);
and U9813 (N_9813,In_456,In_1290);
or U9814 (N_9814,In_2587,In_4367);
and U9815 (N_9815,In_3850,In_3594);
or U9816 (N_9816,In_639,In_751);
or U9817 (N_9817,In_223,In_2350);
and U9818 (N_9818,In_1396,In_4724);
or U9819 (N_9819,In_1493,In_834);
or U9820 (N_9820,In_1582,In_1232);
nor U9821 (N_9821,In_3806,In_2424);
xor U9822 (N_9822,In_3041,In_3100);
nor U9823 (N_9823,In_3821,In_155);
nor U9824 (N_9824,In_4336,In_1358);
or U9825 (N_9825,In_3259,In_825);
or U9826 (N_9826,In_301,In_2017);
xnor U9827 (N_9827,In_4165,In_2411);
xor U9828 (N_9828,In_4695,In_1463);
or U9829 (N_9829,In_2571,In_1155);
nor U9830 (N_9830,In_371,In_1371);
nand U9831 (N_9831,In_4464,In_576);
and U9832 (N_9832,In_703,In_4303);
and U9833 (N_9833,In_1489,In_911);
and U9834 (N_9834,In_4174,In_267);
xor U9835 (N_9835,In_4593,In_2373);
and U9836 (N_9836,In_2244,In_2622);
and U9837 (N_9837,In_764,In_1139);
or U9838 (N_9838,In_4305,In_533);
nand U9839 (N_9839,In_3196,In_3432);
nand U9840 (N_9840,In_4249,In_4768);
and U9841 (N_9841,In_225,In_348);
nand U9842 (N_9842,In_2779,In_683);
nor U9843 (N_9843,In_3658,In_4950);
xor U9844 (N_9844,In_2247,In_1610);
xor U9845 (N_9845,In_2238,In_3270);
nand U9846 (N_9846,In_3604,In_3379);
and U9847 (N_9847,In_1864,In_2920);
nand U9848 (N_9848,In_1406,In_1900);
and U9849 (N_9849,In_3785,In_2399);
nand U9850 (N_9850,In_1490,In_4484);
or U9851 (N_9851,In_3254,In_2795);
or U9852 (N_9852,In_520,In_416);
nand U9853 (N_9853,In_736,In_302);
or U9854 (N_9854,In_4017,In_2619);
and U9855 (N_9855,In_602,In_2786);
nor U9856 (N_9856,In_4198,In_3419);
or U9857 (N_9857,In_2678,In_2981);
nand U9858 (N_9858,In_3839,In_4785);
and U9859 (N_9859,In_2993,In_4110);
and U9860 (N_9860,In_3418,In_2452);
nor U9861 (N_9861,In_1946,In_1217);
and U9862 (N_9862,In_4482,In_1260);
or U9863 (N_9863,In_4203,In_4082);
xor U9864 (N_9864,In_2682,In_3605);
nor U9865 (N_9865,In_4914,In_3320);
and U9866 (N_9866,In_2938,In_4335);
nand U9867 (N_9867,In_4489,In_4847);
xor U9868 (N_9868,In_854,In_3285);
nor U9869 (N_9869,In_2958,In_1648);
xnor U9870 (N_9870,In_1845,In_2299);
or U9871 (N_9871,In_4894,In_4917);
and U9872 (N_9872,In_4506,In_2407);
and U9873 (N_9873,In_3515,In_3218);
or U9874 (N_9874,In_3616,In_742);
and U9875 (N_9875,In_3476,In_2996);
nor U9876 (N_9876,In_75,In_4776);
and U9877 (N_9877,In_4170,In_4469);
and U9878 (N_9878,In_3470,In_4099);
and U9879 (N_9879,In_2481,In_1398);
or U9880 (N_9880,In_2422,In_3279);
and U9881 (N_9881,In_2264,In_4853);
and U9882 (N_9882,In_2620,In_2138);
nand U9883 (N_9883,In_3310,In_2198);
and U9884 (N_9884,In_4003,In_283);
xor U9885 (N_9885,In_2566,In_4230);
and U9886 (N_9886,In_574,In_4611);
nand U9887 (N_9887,In_2212,In_4489);
nor U9888 (N_9888,In_2211,In_3975);
nor U9889 (N_9889,In_3898,In_3768);
and U9890 (N_9890,In_973,In_4188);
or U9891 (N_9891,In_4796,In_3308);
and U9892 (N_9892,In_888,In_747);
nand U9893 (N_9893,In_2294,In_4547);
or U9894 (N_9894,In_882,In_2162);
nand U9895 (N_9895,In_708,In_1725);
xor U9896 (N_9896,In_2974,In_4164);
xnor U9897 (N_9897,In_524,In_2028);
nand U9898 (N_9898,In_2674,In_3353);
nand U9899 (N_9899,In_4773,In_1918);
nor U9900 (N_9900,In_2982,In_1700);
or U9901 (N_9901,In_3339,In_387);
nand U9902 (N_9902,In_4478,In_4109);
nor U9903 (N_9903,In_4252,In_4817);
nand U9904 (N_9904,In_3478,In_1747);
nor U9905 (N_9905,In_1883,In_4949);
and U9906 (N_9906,In_2329,In_4937);
xnor U9907 (N_9907,In_508,In_3973);
and U9908 (N_9908,In_2323,In_837);
and U9909 (N_9909,In_1784,In_3145);
nor U9910 (N_9910,In_4869,In_2778);
and U9911 (N_9911,In_584,In_4550);
or U9912 (N_9912,In_664,In_1276);
nor U9913 (N_9913,In_2316,In_687);
nand U9914 (N_9914,In_620,In_839);
nor U9915 (N_9915,In_1084,In_4286);
nor U9916 (N_9916,In_4546,In_1008);
xor U9917 (N_9917,In_3568,In_742);
nand U9918 (N_9918,In_426,In_867);
nor U9919 (N_9919,In_4901,In_931);
xnor U9920 (N_9920,In_1091,In_2623);
nand U9921 (N_9921,In_11,In_2510);
nand U9922 (N_9922,In_2652,In_1444);
nand U9923 (N_9923,In_451,In_701);
nand U9924 (N_9924,In_581,In_4900);
nand U9925 (N_9925,In_2583,In_3584);
xor U9926 (N_9926,In_4967,In_2671);
nand U9927 (N_9927,In_1929,In_4595);
or U9928 (N_9928,In_1098,In_4656);
and U9929 (N_9929,In_784,In_551);
nor U9930 (N_9930,In_1956,In_4047);
nand U9931 (N_9931,In_4980,In_2676);
nor U9932 (N_9932,In_3507,In_1842);
nor U9933 (N_9933,In_1928,In_702);
nand U9934 (N_9934,In_2851,In_4577);
nand U9935 (N_9935,In_3782,In_1969);
xnor U9936 (N_9936,In_2220,In_187);
nand U9937 (N_9937,In_4000,In_1295);
or U9938 (N_9938,In_2934,In_2730);
nor U9939 (N_9939,In_3400,In_3419);
or U9940 (N_9940,In_4898,In_86);
nor U9941 (N_9941,In_3079,In_3043);
or U9942 (N_9942,In_947,In_1631);
nor U9943 (N_9943,In_3891,In_3618);
nor U9944 (N_9944,In_3063,In_3079);
and U9945 (N_9945,In_4237,In_3063);
xnor U9946 (N_9946,In_4627,In_649);
nand U9947 (N_9947,In_426,In_2005);
and U9948 (N_9948,In_1441,In_3792);
xnor U9949 (N_9949,In_2368,In_3067);
nand U9950 (N_9950,In_740,In_734);
xor U9951 (N_9951,In_3858,In_2971);
nor U9952 (N_9952,In_2282,In_4929);
or U9953 (N_9953,In_1074,In_4235);
nand U9954 (N_9954,In_1737,In_4334);
nor U9955 (N_9955,In_2168,In_3123);
nor U9956 (N_9956,In_1430,In_4401);
and U9957 (N_9957,In_3758,In_4462);
or U9958 (N_9958,In_857,In_3041);
nand U9959 (N_9959,In_1794,In_2038);
and U9960 (N_9960,In_3338,In_4136);
xor U9961 (N_9961,In_3556,In_3424);
or U9962 (N_9962,In_3791,In_714);
nor U9963 (N_9963,In_3891,In_1288);
nor U9964 (N_9964,In_1097,In_4158);
nand U9965 (N_9965,In_200,In_2818);
or U9966 (N_9966,In_1002,In_4496);
nand U9967 (N_9967,In_184,In_1805);
nand U9968 (N_9968,In_581,In_899);
nor U9969 (N_9969,In_286,In_399);
and U9970 (N_9970,In_3387,In_4441);
or U9971 (N_9971,In_2481,In_4109);
and U9972 (N_9972,In_207,In_3410);
nand U9973 (N_9973,In_3907,In_2547);
xnor U9974 (N_9974,In_260,In_3355);
nand U9975 (N_9975,In_2704,In_698);
nand U9976 (N_9976,In_1799,In_1917);
nand U9977 (N_9977,In_357,In_1527);
nand U9978 (N_9978,In_1449,In_3552);
nor U9979 (N_9979,In_797,In_3036);
nand U9980 (N_9980,In_3274,In_1640);
or U9981 (N_9981,In_4907,In_1156);
and U9982 (N_9982,In_4129,In_4575);
or U9983 (N_9983,In_847,In_1429);
nor U9984 (N_9984,In_53,In_4004);
and U9985 (N_9985,In_3095,In_3677);
xor U9986 (N_9986,In_1101,In_1090);
nor U9987 (N_9987,In_1785,In_1989);
and U9988 (N_9988,In_2556,In_2227);
and U9989 (N_9989,In_1596,In_475);
nand U9990 (N_9990,In_2944,In_3461);
nand U9991 (N_9991,In_3206,In_2570);
and U9992 (N_9992,In_4922,In_1415);
xor U9993 (N_9993,In_1395,In_4546);
or U9994 (N_9994,In_2027,In_970);
and U9995 (N_9995,In_894,In_3870);
and U9996 (N_9996,In_414,In_3795);
xnor U9997 (N_9997,In_3895,In_4012);
nand U9998 (N_9998,In_531,In_4295);
and U9999 (N_9999,In_3709,In_3516);
nand U10000 (N_10000,N_6254,N_7620);
nor U10001 (N_10001,N_7245,N_2955);
nor U10002 (N_10002,N_7763,N_6791);
or U10003 (N_10003,N_5503,N_5383);
xnor U10004 (N_10004,N_1940,N_2224);
nor U10005 (N_10005,N_4684,N_5778);
nand U10006 (N_10006,N_9567,N_1206);
or U10007 (N_10007,N_228,N_1528);
or U10008 (N_10008,N_8703,N_5686);
nor U10009 (N_10009,N_8083,N_2913);
or U10010 (N_10010,N_3151,N_4421);
xor U10011 (N_10011,N_1453,N_4437);
or U10012 (N_10012,N_3405,N_4668);
nand U10013 (N_10013,N_2502,N_7333);
or U10014 (N_10014,N_1162,N_4530);
nand U10015 (N_10015,N_2265,N_6054);
or U10016 (N_10016,N_6928,N_9723);
nand U10017 (N_10017,N_2139,N_2940);
nor U10018 (N_10018,N_6412,N_9311);
xnor U10019 (N_10019,N_4690,N_2052);
nand U10020 (N_10020,N_4253,N_485);
nand U10021 (N_10021,N_6460,N_1189);
and U10022 (N_10022,N_4044,N_3642);
nor U10023 (N_10023,N_1689,N_773);
nor U10024 (N_10024,N_860,N_8641);
and U10025 (N_10025,N_7986,N_3066);
or U10026 (N_10026,N_1746,N_5488);
nand U10027 (N_10027,N_402,N_8566);
nand U10028 (N_10028,N_7085,N_7789);
nand U10029 (N_10029,N_7140,N_2378);
nor U10030 (N_10030,N_4754,N_6182);
nand U10031 (N_10031,N_2677,N_9324);
nand U10032 (N_10032,N_4389,N_636);
nand U10033 (N_10033,N_9554,N_2309);
xnor U10034 (N_10034,N_9101,N_9408);
xor U10035 (N_10035,N_2275,N_1575);
nor U10036 (N_10036,N_2576,N_4937);
nor U10037 (N_10037,N_9960,N_4468);
xnor U10038 (N_10038,N_5484,N_2365);
or U10039 (N_10039,N_2086,N_6827);
nor U10040 (N_10040,N_4590,N_8306);
or U10041 (N_10041,N_2698,N_2412);
nor U10042 (N_10042,N_5524,N_2811);
nand U10043 (N_10043,N_4896,N_454);
nand U10044 (N_10044,N_1317,N_924);
and U10045 (N_10045,N_2759,N_9159);
or U10046 (N_10046,N_2213,N_6799);
nand U10047 (N_10047,N_6756,N_8624);
or U10048 (N_10048,N_4003,N_415);
or U10049 (N_10049,N_1181,N_9521);
xnor U10050 (N_10050,N_5122,N_4593);
nand U10051 (N_10051,N_6806,N_4326);
xor U10052 (N_10052,N_3490,N_6171);
nor U10053 (N_10053,N_3541,N_4431);
and U10054 (N_10054,N_1769,N_1525);
and U10055 (N_10055,N_6367,N_4779);
nand U10056 (N_10056,N_5663,N_255);
nand U10057 (N_10057,N_4581,N_2226);
nand U10058 (N_10058,N_3413,N_9828);
or U10059 (N_10059,N_6914,N_9420);
nand U10060 (N_10060,N_8226,N_2301);
nand U10061 (N_10061,N_1134,N_2670);
and U10062 (N_10062,N_3650,N_4118);
or U10063 (N_10063,N_1000,N_9556);
nand U10064 (N_10064,N_3379,N_9171);
nand U10065 (N_10065,N_6464,N_4457);
nand U10066 (N_10066,N_9724,N_6225);
xnor U10067 (N_10067,N_4597,N_1192);
and U10068 (N_10068,N_6555,N_9610);
or U10069 (N_10069,N_1813,N_1442);
or U10070 (N_10070,N_721,N_1369);
nand U10071 (N_10071,N_6295,N_5075);
nand U10072 (N_10072,N_4091,N_7677);
nand U10073 (N_10073,N_6110,N_1685);
nor U10074 (N_10074,N_3664,N_4796);
nor U10075 (N_10075,N_263,N_6729);
nand U10076 (N_10076,N_821,N_9224);
nor U10077 (N_10077,N_604,N_6204);
and U10078 (N_10078,N_4699,N_2454);
nor U10079 (N_10079,N_2985,N_4206);
and U10080 (N_10080,N_8396,N_5829);
or U10081 (N_10081,N_8283,N_9249);
xnor U10082 (N_10082,N_199,N_786);
and U10083 (N_10083,N_500,N_5951);
and U10084 (N_10084,N_7290,N_5769);
or U10085 (N_10085,N_9492,N_7775);
nand U10086 (N_10086,N_9764,N_1750);
or U10087 (N_10087,N_2184,N_4346);
nor U10088 (N_10088,N_2656,N_7900);
or U10089 (N_10089,N_245,N_8469);
nor U10090 (N_10090,N_451,N_1721);
nand U10091 (N_10091,N_1016,N_194);
and U10092 (N_10092,N_737,N_3535);
nor U10093 (N_10093,N_9466,N_5556);
or U10094 (N_10094,N_2229,N_6567);
or U10095 (N_10095,N_3231,N_6489);
and U10096 (N_10096,N_8501,N_164);
nor U10097 (N_10097,N_7435,N_8772);
or U10098 (N_10098,N_6701,N_3037);
or U10099 (N_10099,N_287,N_5938);
nor U10100 (N_10100,N_2369,N_1443);
or U10101 (N_10101,N_9499,N_6209);
or U10102 (N_10102,N_9656,N_7631);
nor U10103 (N_10103,N_448,N_8435);
or U10104 (N_10104,N_8602,N_5643);
xnor U10105 (N_10105,N_8471,N_7328);
nor U10106 (N_10106,N_9563,N_2074);
and U10107 (N_10107,N_5196,N_6874);
nor U10108 (N_10108,N_8953,N_2262);
or U10109 (N_10109,N_3636,N_7637);
or U10110 (N_10110,N_7064,N_9445);
nand U10111 (N_10111,N_3499,N_8645);
or U10112 (N_10112,N_1423,N_3601);
nor U10113 (N_10113,N_3171,N_9193);
and U10114 (N_10114,N_6106,N_4405);
and U10115 (N_10115,N_7248,N_7145);
nor U10116 (N_10116,N_672,N_8242);
nor U10117 (N_10117,N_1218,N_2584);
nor U10118 (N_10118,N_6557,N_4612);
and U10119 (N_10119,N_246,N_4004);
nor U10120 (N_10120,N_8672,N_8094);
and U10121 (N_10121,N_2465,N_3433);
or U10122 (N_10122,N_153,N_6396);
nor U10123 (N_10123,N_9534,N_378);
nand U10124 (N_10124,N_2707,N_6379);
xnor U10125 (N_10125,N_7387,N_1451);
nand U10126 (N_10126,N_5294,N_1270);
and U10127 (N_10127,N_7752,N_4343);
nand U10128 (N_10128,N_1679,N_5188);
nand U10129 (N_10129,N_6831,N_2011);
nor U10130 (N_10130,N_2299,N_5976);
nor U10131 (N_10131,N_5699,N_2162);
or U10132 (N_10132,N_7731,N_417);
nand U10133 (N_10133,N_2113,N_4070);
nand U10134 (N_10134,N_6947,N_7303);
nand U10135 (N_10135,N_8150,N_2921);
or U10136 (N_10136,N_1909,N_5943);
nor U10137 (N_10137,N_6271,N_2484);
nor U10138 (N_10138,N_2946,N_4588);
and U10139 (N_10139,N_8520,N_3838);
nand U10140 (N_10140,N_9646,N_1065);
nor U10141 (N_10141,N_4725,N_5641);
and U10142 (N_10142,N_3337,N_3075);
and U10143 (N_10143,N_8541,N_1572);
and U10144 (N_10144,N_1152,N_6824);
nand U10145 (N_10145,N_5844,N_9963);
nor U10146 (N_10146,N_6141,N_1084);
nand U10147 (N_10147,N_7306,N_8764);
xor U10148 (N_10148,N_6351,N_5625);
and U10149 (N_10149,N_1481,N_9872);
and U10150 (N_10150,N_7548,N_2216);
nor U10151 (N_10151,N_1466,N_7479);
nor U10152 (N_10152,N_7963,N_2540);
nand U10153 (N_10153,N_9890,N_41);
nand U10154 (N_10154,N_1511,N_9865);
xnor U10155 (N_10155,N_9292,N_7592);
nor U10156 (N_10156,N_4744,N_8436);
nor U10157 (N_10157,N_2969,N_151);
nand U10158 (N_10158,N_5368,N_8912);
nor U10159 (N_10159,N_8875,N_6278);
nand U10160 (N_10160,N_6046,N_1165);
and U10161 (N_10161,N_4459,N_3966);
xnor U10162 (N_10162,N_9666,N_3939);
or U10163 (N_10163,N_3842,N_6558);
nor U10164 (N_10164,N_9131,N_4930);
xnor U10165 (N_10165,N_6522,N_6703);
nor U10166 (N_10166,N_5030,N_6109);
nor U10167 (N_10167,N_1363,N_862);
and U10168 (N_10168,N_5825,N_7340);
nand U10169 (N_10169,N_5940,N_6499);
xnor U10170 (N_10170,N_6497,N_2911);
nand U10171 (N_10171,N_9071,N_8340);
xnor U10172 (N_10172,N_3869,N_4358);
and U10173 (N_10173,N_7500,N_8379);
or U10174 (N_10174,N_4815,N_2377);
nand U10175 (N_10175,N_4981,N_4578);
nor U10176 (N_10176,N_5884,N_6895);
nand U10177 (N_10177,N_8699,N_9645);
or U10178 (N_10178,N_9954,N_442);
xor U10179 (N_10179,N_9412,N_5013);
or U10180 (N_10180,N_8720,N_3021);
nand U10181 (N_10181,N_1349,N_7608);
nand U10182 (N_10182,N_1148,N_9677);
or U10183 (N_10183,N_9252,N_9941);
xor U10184 (N_10184,N_3539,N_9746);
or U10185 (N_10185,N_9630,N_2725);
nand U10186 (N_10186,N_811,N_4219);
and U10187 (N_10187,N_7337,N_8515);
and U10188 (N_10188,N_5486,N_9273);
xnor U10189 (N_10189,N_6378,N_9075);
and U10190 (N_10190,N_7537,N_7282);
or U10191 (N_10191,N_3773,N_8626);
or U10192 (N_10192,N_9355,N_1615);
nor U10193 (N_10193,N_2679,N_9776);
nand U10194 (N_10194,N_6222,N_8255);
nand U10195 (N_10195,N_6898,N_9018);
nand U10196 (N_10196,N_5813,N_8782);
xor U10197 (N_10197,N_9529,N_3169);
nand U10198 (N_10198,N_5847,N_1147);
and U10199 (N_10199,N_439,N_3924);
nor U10200 (N_10200,N_2882,N_2939);
and U10201 (N_10201,N_5968,N_5793);
nand U10202 (N_10202,N_8884,N_6298);
or U10203 (N_10203,N_2305,N_4341);
nor U10204 (N_10204,N_8911,N_3894);
xor U10205 (N_10205,N_6656,N_1810);
and U10206 (N_10206,N_9548,N_2518);
nor U10207 (N_10207,N_3761,N_5948);
and U10208 (N_10208,N_4085,N_9109);
or U10209 (N_10209,N_6443,N_6749);
nor U10210 (N_10210,N_7645,N_7669);
or U10211 (N_10211,N_4946,N_2346);
xor U10212 (N_10212,N_5722,N_3108);
or U10213 (N_10213,N_7975,N_7120);
nor U10214 (N_10214,N_3166,N_8757);
nor U10215 (N_10215,N_2862,N_602);
nor U10216 (N_10216,N_4702,N_6491);
or U10217 (N_10217,N_6671,N_3242);
nand U10218 (N_10218,N_9036,N_2081);
nand U10219 (N_10219,N_7091,N_2467);
nand U10220 (N_10220,N_3915,N_5192);
nor U10221 (N_10221,N_3055,N_8768);
and U10222 (N_10222,N_5420,N_2401);
or U10223 (N_10223,N_4477,N_7066);
nor U10224 (N_10224,N_4931,N_7440);
nand U10225 (N_10225,N_2239,N_4414);
and U10226 (N_10226,N_5199,N_9932);
nand U10227 (N_10227,N_7054,N_8366);
and U10228 (N_10228,N_4209,N_7933);
or U10229 (N_10229,N_8747,N_5495);
nor U10230 (N_10230,N_8568,N_3307);
xnor U10231 (N_10231,N_1979,N_9837);
nand U10232 (N_10232,N_7401,N_9191);
and U10233 (N_10233,N_5150,N_2522);
and U10234 (N_10234,N_4628,N_1578);
and U10235 (N_10235,N_8742,N_9952);
and U10236 (N_10236,N_2536,N_5953);
and U10237 (N_10237,N_9831,N_1239);
nor U10238 (N_10238,N_3935,N_9429);
xor U10239 (N_10239,N_3571,N_8290);
or U10240 (N_10240,N_385,N_5770);
nand U10241 (N_10241,N_7258,N_870);
xnor U10242 (N_10242,N_2713,N_7902);
and U10243 (N_10243,N_1989,N_8861);
nand U10244 (N_10244,N_8453,N_8837);
and U10245 (N_10245,N_7260,N_3873);
nand U10246 (N_10246,N_8298,N_6542);
or U10247 (N_10247,N_7681,N_9126);
or U10248 (N_10248,N_8456,N_2127);
or U10249 (N_10249,N_7094,N_6334);
nand U10250 (N_10250,N_4146,N_9008);
nand U10251 (N_10251,N_7345,N_9937);
or U10252 (N_10252,N_2871,N_842);
nand U10253 (N_10253,N_8786,N_7257);
xor U10254 (N_10254,N_21,N_3450);
nand U10255 (N_10255,N_7491,N_8955);
nand U10256 (N_10256,N_7795,N_4256);
nor U10257 (N_10257,N_9119,N_2566);
nor U10258 (N_10258,N_7286,N_2787);
or U10259 (N_10259,N_1724,N_4051);
xnor U10260 (N_10260,N_8548,N_1175);
and U10261 (N_10261,N_3787,N_4288);
and U10262 (N_10262,N_123,N_8622);
and U10263 (N_10263,N_5466,N_7720);
or U10264 (N_10264,N_3024,N_8677);
or U10265 (N_10265,N_183,N_6207);
nand U10266 (N_10266,N_6201,N_1786);
nand U10267 (N_10267,N_9857,N_5279);
and U10268 (N_10268,N_9504,N_7873);
and U10269 (N_10269,N_6939,N_3095);
xnor U10270 (N_10270,N_3834,N_6473);
and U10271 (N_10271,N_8274,N_5592);
or U10272 (N_10272,N_1797,N_5520);
nand U10273 (N_10273,N_8897,N_8507);
or U10274 (N_10274,N_3597,N_3440);
nand U10275 (N_10275,N_393,N_4582);
nor U10276 (N_10276,N_5760,N_2119);
nor U10277 (N_10277,N_7612,N_1913);
nand U10278 (N_10278,N_4756,N_6265);
xor U10279 (N_10279,N_5406,N_6150);
or U10280 (N_10280,N_510,N_4800);
xor U10281 (N_10281,N_7061,N_4285);
and U10282 (N_10282,N_192,N_7743);
nor U10283 (N_10283,N_4408,N_3149);
nand U10284 (N_10284,N_2680,N_9508);
nand U10285 (N_10285,N_9417,N_4888);
and U10286 (N_10286,N_5692,N_735);
nor U10287 (N_10287,N_3442,N_8933);
nor U10288 (N_10288,N_7630,N_8365);
or U10289 (N_10289,N_1513,N_148);
nor U10290 (N_10290,N_3871,N_5883);
nor U10291 (N_10291,N_3339,N_9169);
and U10292 (N_10292,N_798,N_9513);
and U10293 (N_10293,N_6640,N_1322);
or U10294 (N_10294,N_6543,N_105);
or U10295 (N_10295,N_8315,N_8798);
nor U10296 (N_10296,N_2782,N_8657);
nor U10297 (N_10297,N_7170,N_9357);
nor U10298 (N_10298,N_4021,N_2355);
or U10299 (N_10299,N_8830,N_3501);
and U10300 (N_10300,N_3395,N_1145);
nand U10301 (N_10301,N_1372,N_3619);
nor U10302 (N_10302,N_6813,N_9869);
nand U10303 (N_10303,N_4489,N_2960);
and U10304 (N_10304,N_9956,N_8107);
nor U10305 (N_10305,N_2555,N_6883);
xnor U10306 (N_10306,N_351,N_994);
nor U10307 (N_10307,N_3796,N_7060);
xor U10308 (N_10308,N_6976,N_976);
or U10309 (N_10309,N_3243,N_1986);
nand U10310 (N_10310,N_3431,N_7105);
or U10311 (N_10311,N_1843,N_6326);
and U10312 (N_10312,N_966,N_138);
xnor U10313 (N_10313,N_1938,N_5066);
or U10314 (N_10314,N_1187,N_2743);
nand U10315 (N_10315,N_8449,N_7126);
nor U10316 (N_10316,N_4507,N_6145);
nor U10317 (N_10317,N_3691,N_8753);
nor U10318 (N_10318,N_4481,N_3759);
nor U10319 (N_10319,N_4830,N_9226);
nand U10320 (N_10320,N_2268,N_2270);
or U10321 (N_10321,N_2036,N_3793);
nor U10322 (N_10322,N_9091,N_5263);
nand U10323 (N_10323,N_4005,N_8674);
or U10324 (N_10324,N_9392,N_9251);
or U10325 (N_10325,N_163,N_1414);
and U10326 (N_10326,N_2741,N_1855);
nand U10327 (N_10327,N_3191,N_1108);
nor U10328 (N_10328,N_1256,N_4592);
nand U10329 (N_10329,N_5243,N_9892);
or U10330 (N_10330,N_6977,N_7143);
nand U10331 (N_10331,N_7147,N_1620);
and U10332 (N_10332,N_7542,N_6935);
and U10333 (N_10333,N_3570,N_3746);
nor U10334 (N_10334,N_7541,N_5664);
nand U10335 (N_10335,N_2009,N_2188);
nand U10336 (N_10336,N_9943,N_95);
nor U10337 (N_10337,N_777,N_5372);
nor U10338 (N_10338,N_6335,N_4040);
nand U10339 (N_10339,N_4281,N_6629);
and U10340 (N_10340,N_8195,N_3953);
and U10341 (N_10341,N_6828,N_4991);
nor U10342 (N_10342,N_2579,N_3212);
xor U10343 (N_10343,N_5756,N_1751);
nor U10344 (N_10344,N_6534,N_2408);
nand U10345 (N_10345,N_7312,N_757);
nor U10346 (N_10346,N_8093,N_2280);
nor U10347 (N_10347,N_1069,N_3366);
xor U10348 (N_10348,N_8258,N_1114);
nor U10349 (N_10349,N_5293,N_4221);
or U10350 (N_10350,N_8136,N_3768);
nor U10351 (N_10351,N_1653,N_4058);
or U10352 (N_10352,N_4910,N_2646);
or U10353 (N_10353,N_3273,N_7729);
nor U10354 (N_10354,N_3950,N_9056);
or U10355 (N_10355,N_6167,N_2187);
or U10356 (N_10356,N_32,N_2855);
nand U10357 (N_10357,N_6600,N_3250);
and U10358 (N_10358,N_7368,N_4988);
and U10359 (N_10359,N_5238,N_7034);
nand U10360 (N_10360,N_883,N_1215);
nand U10361 (N_10361,N_8658,N_6162);
and U10362 (N_10362,N_3685,N_6230);
nand U10363 (N_10363,N_4833,N_2138);
nand U10364 (N_10364,N_2144,N_2409);
or U10365 (N_10365,N_7661,N_2668);
xor U10366 (N_10366,N_2828,N_5442);
and U10367 (N_10367,N_9260,N_3583);
or U10368 (N_10368,N_714,N_8237);
and U10369 (N_10369,N_2423,N_2835);
xnor U10370 (N_10370,N_6197,N_4338);
and U10371 (N_10371,N_2427,N_7380);
nor U10372 (N_10372,N_62,N_7349);
nor U10373 (N_10373,N_8175,N_992);
nor U10374 (N_10374,N_8803,N_9322);
nor U10375 (N_10375,N_5559,N_9544);
and U10376 (N_10376,N_6119,N_7636);
and U10377 (N_10377,N_3623,N_2128);
and U10378 (N_10378,N_9207,N_7448);
or U10379 (N_10379,N_4994,N_4456);
xnor U10380 (N_10380,N_6851,N_5631);
xnor U10381 (N_10381,N_3609,N_8430);
nand U10382 (N_10382,N_9817,N_7182);
xor U10383 (N_10383,N_8654,N_1749);
or U10384 (N_10384,N_5273,N_8969);
xnor U10385 (N_10385,N_6089,N_1139);
nand U10386 (N_10386,N_8606,N_6366);
nand U10387 (N_10387,N_4843,N_57);
nand U10388 (N_10388,N_140,N_1500);
or U10389 (N_10389,N_1088,N_5250);
xnor U10390 (N_10390,N_7334,N_7646);
nand U10391 (N_10391,N_5048,N_1586);
nand U10392 (N_10392,N_7213,N_1561);
nor U10393 (N_10393,N_7800,N_1155);
xnor U10394 (N_10394,N_6773,N_1745);
and U10395 (N_10395,N_3958,N_1567);
nand U10396 (N_10396,N_8527,N_2770);
and U10397 (N_10397,N_4924,N_6730);
or U10398 (N_10398,N_7651,N_468);
and U10399 (N_10399,N_1240,N_2303);
xor U10400 (N_10400,N_9722,N_700);
and U10401 (N_10401,N_8984,N_9367);
xor U10402 (N_10402,N_7294,N_9898);
nor U10403 (N_10403,N_5055,N_1129);
nand U10404 (N_10404,N_3012,N_5833);
and U10405 (N_10405,N_7313,N_655);
nor U10406 (N_10406,N_7002,N_1857);
xor U10407 (N_10407,N_5001,N_1393);
nor U10408 (N_10408,N_1639,N_7960);
nor U10409 (N_10409,N_7081,N_9745);
xor U10410 (N_10410,N_7507,N_9073);
nand U10411 (N_10411,N_2984,N_1600);
and U10412 (N_10412,N_7850,N_6093);
nand U10413 (N_10413,N_4989,N_1335);
nor U10414 (N_10414,N_5343,N_5921);
nor U10415 (N_10415,N_749,N_2282);
nor U10416 (N_10416,N_6525,N_91);
or U10417 (N_10417,N_34,N_5173);
or U10418 (N_10418,N_9195,N_6206);
or U10419 (N_10419,N_3092,N_1761);
nor U10420 (N_10420,N_1957,N_7115);
or U10421 (N_10421,N_8766,N_1936);
and U10422 (N_10422,N_8896,N_9482);
or U10423 (N_10423,N_3743,N_4799);
and U10424 (N_10424,N_6362,N_3270);
or U10425 (N_10425,N_8809,N_4322);
or U10426 (N_10426,N_7240,N_7329);
nor U10427 (N_10427,N_2609,N_5955);
nor U10428 (N_10428,N_8082,N_2846);
nand U10429 (N_10429,N_3819,N_9986);
and U10430 (N_10430,N_9232,N_3982);
or U10431 (N_10431,N_704,N_9069);
or U10432 (N_10432,N_3102,N_4151);
or U10433 (N_10433,N_7087,N_6886);
or U10434 (N_10434,N_5843,N_5816);
nand U10435 (N_10435,N_1559,N_680);
or U10436 (N_10436,N_9961,N_6784);
xor U10437 (N_10437,N_7203,N_7227);
nor U10438 (N_10438,N_2116,N_4311);
nand U10439 (N_10439,N_4733,N_5453);
xnor U10440 (N_10440,N_5511,N_7136);
nor U10441 (N_10441,N_3224,N_6273);
or U10442 (N_10442,N_8944,N_107);
and U10443 (N_10443,N_7019,N_2868);
and U10444 (N_10444,N_1978,N_2788);
and U10445 (N_10445,N_6312,N_428);
and U10446 (N_10446,N_3030,N_5164);
nand U10447 (N_10447,N_7872,N_1827);
nand U10448 (N_10448,N_7351,N_9222);
or U10449 (N_10449,N_5204,N_3641);
xor U10450 (N_10450,N_4783,N_5278);
nor U10451 (N_10451,N_1988,N_2329);
or U10452 (N_10452,N_8752,N_3926);
or U10453 (N_10453,N_3100,N_9518);
nand U10454 (N_10454,N_7642,N_950);
or U10455 (N_10455,N_8026,N_9374);
nor U10456 (N_10456,N_6909,N_4101);
or U10457 (N_10457,N_4920,N_7639);
xnor U10458 (N_10458,N_8659,N_8223);
nor U10459 (N_10459,N_4719,N_4517);
nand U10460 (N_10460,N_2389,N_930);
and U10461 (N_10461,N_816,N_9144);
or U10462 (N_10462,N_8280,N_3375);
nand U10463 (N_10463,N_2874,N_2498);
and U10464 (N_10464,N_4826,N_4381);
nor U10465 (N_10465,N_970,N_8412);
and U10466 (N_10466,N_5029,N_7648);
nand U10467 (N_10467,N_5254,N_1460);
nor U10468 (N_10468,N_2562,N_4672);
and U10469 (N_10469,N_8410,N_3138);
or U10470 (N_10470,N_927,N_1228);
nor U10471 (N_10471,N_6900,N_5277);
nor U10472 (N_10472,N_5257,N_4637);
and U10473 (N_10473,N_5908,N_6921);
nand U10474 (N_10474,N_7177,N_6665);
and U10475 (N_10475,N_7318,N_1966);
nor U10476 (N_10476,N_7922,N_4982);
nand U10477 (N_10477,N_7176,N_4184);
or U10478 (N_10478,N_2819,N_5717);
and U10479 (N_10479,N_5918,N_5915);
nand U10480 (N_10480,N_4724,N_6760);
nor U10481 (N_10481,N_6668,N_7658);
or U10482 (N_10482,N_1632,N_8444);
and U10483 (N_10483,N_1395,N_8231);
xor U10484 (N_10484,N_1116,N_4386);
xnor U10485 (N_10485,N_4138,N_4420);
nand U10486 (N_10486,N_657,N_4079);
nand U10487 (N_10487,N_1174,N_4753);
and U10488 (N_10488,N_6053,N_5726);
nand U10489 (N_10489,N_2934,N_3510);
xnor U10490 (N_10490,N_3398,N_5393);
nand U10491 (N_10491,N_5041,N_8445);
nor U10492 (N_10492,N_5,N_1052);
nor U10493 (N_10493,N_8112,N_7361);
nor U10494 (N_10494,N_1245,N_1506);
and U10495 (N_10495,N_6172,N_1);
nor U10496 (N_10496,N_2927,N_5589);
nor U10497 (N_10497,N_1983,N_2507);
and U10498 (N_10498,N_7896,N_6363);
or U10499 (N_10499,N_5930,N_2165);
xor U10500 (N_10500,N_6342,N_3962);
and U10501 (N_10501,N_3709,N_3071);
and U10502 (N_10502,N_395,N_8029);
nor U10503 (N_10503,N_1484,N_8333);
and U10504 (N_10504,N_2242,N_7906);
or U10505 (N_10505,N_1430,N_1259);
or U10506 (N_10506,N_3513,N_7870);
nand U10507 (N_10507,N_167,N_3059);
nor U10508 (N_10508,N_7848,N_8177);
nor U10509 (N_10509,N_9787,N_6331);
nor U10510 (N_10510,N_5322,N_8995);
or U10511 (N_10511,N_7048,N_2891);
nor U10512 (N_10512,N_7032,N_6468);
or U10513 (N_10513,N_8709,N_692);
and U10514 (N_10514,N_8665,N_8186);
nand U10515 (N_10515,N_4204,N_8097);
nor U10516 (N_10516,N_5605,N_6448);
xnor U10517 (N_10517,N_1151,N_1015);
and U10518 (N_10518,N_5773,N_1930);
nor U10519 (N_10519,N_2368,N_7317);
nor U10520 (N_10520,N_8384,N_5445);
nand U10521 (N_10521,N_6603,N_1555);
or U10522 (N_10522,N_9512,N_159);
nor U10523 (N_10523,N_4728,N_3304);
and U10524 (N_10524,N_1438,N_6708);
and U10525 (N_10525,N_4474,N_707);
and U10526 (N_10526,N_7841,N_1943);
nor U10527 (N_10527,N_7803,N_5473);
and U10528 (N_10528,N_4697,N_9125);
nand U10529 (N_10529,N_1692,N_3081);
nand U10530 (N_10530,N_3692,N_8165);
nand U10531 (N_10531,N_5874,N_3536);
and U10532 (N_10532,N_2418,N_6679);
nor U10533 (N_10533,N_531,N_3705);
nor U10534 (N_10534,N_9919,N_1313);
nor U10535 (N_10535,N_8421,N_2064);
or U10536 (N_10536,N_6919,N_1924);
nor U10537 (N_10537,N_9959,N_4643);
nor U10538 (N_10538,N_738,N_3698);
and U10539 (N_10539,N_6394,N_5378);
and U10540 (N_10540,N_545,N_7942);
nand U10541 (N_10541,N_8392,N_7887);
nor U10542 (N_10542,N_6872,N_6636);
or U10543 (N_10543,N_7528,N_8916);
and U10544 (N_10544,N_9204,N_701);
or U10545 (N_10545,N_4603,N_5914);
nand U10546 (N_10546,N_3369,N_9991);
or U10547 (N_10547,N_3061,N_5078);
and U10548 (N_10548,N_4862,N_3550);
or U10549 (N_10549,N_3420,N_9285);
nor U10550 (N_10550,N_7659,N_1316);
nor U10551 (N_10551,N_6982,N_4987);
or U10552 (N_10552,N_5881,N_9346);
nor U10553 (N_10553,N_5049,N_3031);
nor U10554 (N_10554,N_4497,N_9885);
or U10555 (N_10555,N_4797,N_4669);
or U10556 (N_10556,N_3569,N_2252);
nand U10557 (N_10557,N_9843,N_111);
xor U10558 (N_10558,N_5713,N_3504);
and U10559 (N_10559,N_209,N_6503);
nor U10560 (N_10560,N_3426,N_1385);
nand U10561 (N_10561,N_8569,N_3298);
nor U10562 (N_10562,N_9726,N_9253);
nor U10563 (N_10563,N_6250,N_606);
or U10564 (N_10564,N_9319,N_6893);
or U10565 (N_10565,N_3695,N_7668);
nor U10566 (N_10566,N_1975,N_5081);
and U10567 (N_10567,N_4266,N_1719);
nand U10568 (N_10568,N_8061,N_9203);
or U10569 (N_10569,N_904,N_977);
nor U10570 (N_10570,N_3751,N_9184);
or U10571 (N_10571,N_5802,N_3988);
nor U10572 (N_10572,N_182,N_3844);
and U10573 (N_10573,N_4731,N_1302);
nor U10574 (N_10574,N_3190,N_7157);
xor U10575 (N_10575,N_6074,N_368);
nand U10576 (N_10576,N_5830,N_7384);
and U10577 (N_10577,N_486,N_9989);
nand U10578 (N_10578,N_2457,N_7974);
nor U10579 (N_10579,N_2040,N_3602);
and U10580 (N_10580,N_7302,N_525);
or U10581 (N_10581,N_9942,N_8415);
or U10582 (N_10582,N_5230,N_4899);
and U10583 (N_10583,N_760,N_6233);
or U10584 (N_10584,N_7324,N_8104);
or U10585 (N_10585,N_6487,N_363);
and U10586 (N_10586,N_996,N_6885);
and U10587 (N_10587,N_8835,N_2626);
nor U10588 (N_10588,N_6076,N_4777);
nand U10589 (N_10589,N_1252,N_8836);
and U10590 (N_10590,N_1703,N_3124);
and U10591 (N_10591,N_2712,N_201);
xnor U10592 (N_10592,N_9582,N_6533);
or U10593 (N_10593,N_8004,N_9199);
nor U10594 (N_10594,N_2172,N_109);
and U10595 (N_10595,N_327,N_5868);
or U10596 (N_10596,N_1563,N_2313);
or U10597 (N_10597,N_3207,N_5171);
xnor U10598 (N_10598,N_9465,N_2143);
nand U10599 (N_10599,N_5053,N_8791);
or U10600 (N_10600,N_4249,N_2211);
and U10601 (N_10601,N_418,N_534);
nor U10602 (N_10602,N_9759,N_5835);
nand U10603 (N_10603,N_9781,N_6264);
and U10604 (N_10604,N_7478,N_2784);
nor U10605 (N_10605,N_6240,N_978);
nand U10606 (N_10606,N_6219,N_9325);
nor U10607 (N_10607,N_2145,N_420);
nand U10608 (N_10608,N_3042,N_7080);
or U10609 (N_10609,N_7268,N_9241);
and U10610 (N_10610,N_2995,N_6452);
or U10611 (N_10611,N_9629,N_5353);
nand U10612 (N_10612,N_9416,N_2024);
or U10613 (N_10613,N_2571,N_7649);
and U10614 (N_10614,N_9995,N_1244);
or U10615 (N_10615,N_5581,N_1713);
or U10616 (N_10616,N_9536,N_4010);
nand U10617 (N_10617,N_5619,N_9061);
nand U10618 (N_10618,N_3246,N_7654);
or U10619 (N_10619,N_1850,N_8690);
or U10620 (N_10620,N_7383,N_583);
nor U10621 (N_10621,N_3377,N_1780);
xor U10622 (N_10622,N_6127,N_461);
and U10623 (N_10623,N_8334,N_8592);
or U10624 (N_10624,N_1005,N_2825);
and U10625 (N_10625,N_4679,N_6706);
and U10626 (N_10626,N_5746,N_597);
nor U10627 (N_10627,N_3995,N_1200);
nand U10628 (N_10628,N_1459,N_7216);
and U10629 (N_10629,N_367,N_3117);
and U10630 (N_10630,N_2719,N_9316);
nand U10631 (N_10631,N_7492,N_3856);
nor U10632 (N_10632,N_3652,N_8959);
and U10633 (N_10633,N_7560,N_2154);
and U10634 (N_10634,N_2736,N_7992);
and U10635 (N_10635,N_2883,N_121);
or U10636 (N_10636,N_3595,N_376);
and U10637 (N_10637,N_938,N_13);
or U10638 (N_10638,N_3791,N_6616);
and U10639 (N_10639,N_2971,N_565);
xor U10640 (N_10640,N_3526,N_4917);
or U10641 (N_10641,N_9849,N_8694);
or U10642 (N_10642,N_7705,N_9683);
or U10643 (N_10643,N_2339,N_7434);
and U10644 (N_10644,N_5218,N_5612);
nor U10645 (N_10645,N_6941,N_1712);
nor U10646 (N_10646,N_3621,N_5644);
nor U10647 (N_10647,N_5032,N_8321);
and U10648 (N_10648,N_5822,N_460);
nor U10649 (N_10649,N_3058,N_9501);
nand U10650 (N_10650,N_9969,N_1499);
nand U10651 (N_10651,N_1199,N_3314);
or U10652 (N_10652,N_948,N_3093);
nand U10653 (N_10653,N_3396,N_6761);
nand U10654 (N_10654,N_5172,N_675);
nand U10655 (N_10655,N_1952,N_4027);
and U10656 (N_10656,N_984,N_6344);
nor U10657 (N_10657,N_2010,N_9112);
nand U10658 (N_10658,N_8464,N_9791);
nor U10659 (N_10659,N_5916,N_8673);
nor U10660 (N_10660,N_2122,N_1053);
nand U10661 (N_10661,N_6463,N_2073);
nand U10662 (N_10662,N_7624,N_4246);
xor U10663 (N_10663,N_7450,N_6327);
nor U10664 (N_10664,N_301,N_8182);
or U10665 (N_10665,N_2756,N_5015);
nand U10666 (N_10666,N_6126,N_8152);
nor U10667 (N_10667,N_5611,N_4875);
nor U10668 (N_10668,N_495,N_6694);
or U10669 (N_10669,N_5371,N_1318);
or U10670 (N_10670,N_3945,N_5364);
or U10671 (N_10671,N_8135,N_8976);
and U10672 (N_10672,N_7148,N_5043);
and U10673 (N_10673,N_3449,N_5740);
nand U10674 (N_10674,N_4026,N_8792);
or U10675 (N_10675,N_9296,N_4160);
and U10676 (N_10676,N_2574,N_4192);
or U10677 (N_10677,N_1714,N_1131);
nor U10678 (N_10678,N_3148,N_7829);
nor U10679 (N_10679,N_3423,N_3778);
and U10680 (N_10680,N_1492,N_6612);
or U10681 (N_10681,N_7389,N_9029);
or U10682 (N_10682,N_6689,N_3999);
or U10683 (N_10683,N_6981,N_2472);
and U10684 (N_10684,N_9481,N_3089);
xnor U10685 (N_10685,N_9005,N_7519);
or U10686 (N_10686,N_4105,N_5424);
or U10687 (N_10687,N_5788,N_2254);
nor U10688 (N_10688,N_1802,N_7278);
nand U10689 (N_10689,N_3806,N_4745);
and U10690 (N_10690,N_3113,N_4531);
nand U10691 (N_10691,N_9210,N_1830);
nor U10692 (N_10692,N_2854,N_8589);
and U10693 (N_10693,N_3774,N_1782);
nor U10694 (N_10694,N_6354,N_5695);
nand U10695 (N_10695,N_4524,N_770);
or U10696 (N_10696,N_3755,N_9541);
nor U10697 (N_10697,N_4810,N_756);
and U10698 (N_10698,N_7811,N_4046);
nor U10699 (N_10699,N_2796,N_4908);
or U10700 (N_10700,N_4866,N_9403);
or U10701 (N_10701,N_3931,N_6750);
and U10702 (N_10702,N_1507,N_232);
and U10703 (N_10703,N_3101,N_4509);
or U10704 (N_10704,N_2922,N_7683);
and U10705 (N_10705,N_5019,N_3852);
or U10706 (N_10706,N_218,N_3216);
xnor U10707 (N_10707,N_5467,N_868);
nor U10708 (N_10708,N_1565,N_3973);
and U10709 (N_10709,N_7432,N_5228);
nor U10710 (N_10710,N_1300,N_211);
nand U10711 (N_10711,N_3335,N_3767);
or U10712 (N_10712,N_5669,N_1153);
or U10713 (N_10713,N_158,N_6477);
and U10714 (N_10714,N_4939,N_7741);
or U10715 (N_10715,N_2233,N_7050);
nand U10716 (N_10716,N_5485,N_5934);
xor U10717 (N_10717,N_3088,N_522);
nand U10718 (N_10718,N_3473,N_180);
or U10719 (N_10719,N_3943,N_8363);
or U10720 (N_10720,N_2696,N_2501);
nor U10721 (N_10721,N_2648,N_5342);
and U10722 (N_10722,N_5775,N_2494);
xor U10723 (N_10723,N_9561,N_222);
nor U10724 (N_10724,N_8414,N_1917);
or U10725 (N_10725,N_168,N_2269);
xnor U10726 (N_10726,N_89,N_4383);
xnor U10727 (N_10727,N_6359,N_5472);
xor U10728 (N_10728,N_9140,N_4586);
xor U10729 (N_10729,N_6672,N_9994);
xor U10730 (N_10730,N_3916,N_6287);
and U10731 (N_10731,N_9916,N_7931);
and U10732 (N_10732,N_9017,N_1716);
nand U10733 (N_10733,N_8220,N_8455);
nand U10734 (N_10734,N_4465,N_9568);
or U10735 (N_10735,N_9700,N_9751);
nand U10736 (N_10736,N_6692,N_1535);
or U10737 (N_10737,N_7410,N_8818);
xnor U10738 (N_10738,N_273,N_9879);
nor U10739 (N_10739,N_3593,N_2688);
and U10740 (N_10740,N_1008,N_4020);
and U10741 (N_10741,N_3111,N_9844);
xor U10742 (N_10742,N_5265,N_6792);
nor U10743 (N_10743,N_127,N_6627);
nand U10744 (N_10744,N_4566,N_8863);
and U10745 (N_10745,N_12,N_1059);
and U10746 (N_10746,N_7471,N_4030);
or U10747 (N_10747,N_9609,N_7160);
and U10748 (N_10748,N_6820,N_9797);
nor U10749 (N_10749,N_2519,N_1982);
or U10750 (N_10750,N_394,N_8294);
and U10751 (N_10751,N_8954,N_1480);
xor U10752 (N_10752,N_2704,N_5790);
nand U10753 (N_10753,N_3910,N_6907);
and U10754 (N_10754,N_7633,N_84);
nor U10755 (N_10755,N_2104,N_7454);
or U10756 (N_10756,N_1142,N_5850);
and U10757 (N_10757,N_8966,N_8176);
and U10758 (N_10758,N_7496,N_4995);
nand U10759 (N_10759,N_2331,N_3282);
nor U10760 (N_10760,N_5725,N_8394);
xnor U10761 (N_10761,N_5160,N_6135);
nand U10762 (N_10762,N_8494,N_1832);
nand U10763 (N_10763,N_4819,N_9717);
nor U10764 (N_10764,N_3401,N_4904);
xnor U10765 (N_10765,N_8372,N_8889);
nand U10766 (N_10766,N_8614,N_8200);
nand U10767 (N_10767,N_1276,N_5533);
or U10768 (N_10768,N_3599,N_4033);
nand U10769 (N_10769,N_5255,N_5253);
and U10770 (N_10770,N_3552,N_8914);
and U10771 (N_10771,N_9557,N_6626);
or U10772 (N_10772,N_6724,N_6581);
nand U10773 (N_10773,N_6620,N_53);
nand U10774 (N_10774,N_5547,N_7441);
nor U10775 (N_10775,N_844,N_1104);
nor U10776 (N_10776,N_974,N_6441);
nand U10777 (N_10777,N_8844,N_2135);
nor U10778 (N_10778,N_4778,N_7460);
nand U10779 (N_10779,N_3329,N_4568);
or U10780 (N_10780,N_4916,N_4302);
nand U10781 (N_10781,N_2066,N_9361);
nor U10782 (N_10782,N_6840,N_9712);
nor U10783 (N_10783,N_7884,N_3181);
and U10784 (N_10784,N_305,N_8126);
nor U10785 (N_10785,N_5550,N_373);
and U10786 (N_10786,N_4895,N_1728);
and U10787 (N_10787,N_9435,N_3610);
and U10788 (N_10788,N_855,N_4055);
and U10789 (N_10789,N_8817,N_2544);
nor U10790 (N_10790,N_4348,N_4980);
nor U10791 (N_10791,N_8288,N_5554);
nor U10792 (N_10792,N_3009,N_4495);
or U10793 (N_10793,N_1150,N_9708);
or U10794 (N_10794,N_8230,N_2841);
and U10795 (N_10795,N_780,N_886);
or U10796 (N_10796,N_4767,N_6371);
and U10797 (N_10797,N_6255,N_5623);
and U10798 (N_10798,N_7028,N_5706);
nor U10799 (N_10799,N_3855,N_2530);
and U10800 (N_10800,N_4696,N_205);
nand U10801 (N_10801,N_1094,N_8555);
nand U10802 (N_10802,N_7205,N_7740);
nand U10803 (N_10803,N_6746,N_2203);
nor U10804 (N_10804,N_6666,N_4547);
xor U10805 (N_10805,N_8199,N_845);
and U10806 (N_10806,N_5786,N_1113);
or U10807 (N_10807,N_967,N_8138);
nand U10808 (N_10808,N_6843,N_2959);
nor U10809 (N_10809,N_6556,N_3616);
nor U10810 (N_10810,N_804,N_9675);
and U10811 (N_10811,N_9808,N_3228);
and U10812 (N_10812,N_2381,N_1125);
or U10813 (N_10813,N_2592,N_2754);
or U10814 (N_10814,N_7192,N_8295);
nand U10815 (N_10815,N_705,N_7388);
nand U10816 (N_10816,N_7239,N_3053);
nand U10817 (N_10817,N_1030,N_7909);
or U10818 (N_10818,N_2761,N_3276);
or U10819 (N_10819,N_4485,N_3415);
nand U10820 (N_10820,N_268,N_7212);
nor U10821 (N_10821,N_8197,N_9180);
and U10822 (N_10822,N_3987,N_9010);
nor U10823 (N_10823,N_4828,N_306);
nor U10824 (N_10824,N_491,N_6274);
or U10825 (N_10825,N_177,N_2824);
xnor U10826 (N_10826,N_1512,N_9642);
nor U10827 (N_10827,N_3519,N_6383);
and U10828 (N_10828,N_6816,N_4131);
and U10829 (N_10829,N_908,N_796);
or U10830 (N_10830,N_4580,N_1248);
xnor U10831 (N_10831,N_679,N_456);
and U10832 (N_10832,N_6244,N_9957);
and U10833 (N_10833,N_1914,N_998);
or U10834 (N_10834,N_7934,N_4175);
xnor U10835 (N_10835,N_9001,N_288);
and U10836 (N_10836,N_7877,N_1392);
or U10837 (N_10837,N_8859,N_1223);
and U10838 (N_10838,N_7966,N_4922);
and U10839 (N_10839,N_3370,N_3263);
and U10840 (N_10840,N_9535,N_4997);
xor U10841 (N_10841,N_7842,N_4501);
nand U10842 (N_10842,N_2030,N_3394);
nand U10843 (N_10843,N_2376,N_4073);
nor U10844 (N_10844,N_2945,N_1367);
nand U10845 (N_10845,N_8188,N_5919);
and U10846 (N_10846,N_2003,N_2933);
nand U10847 (N_10847,N_9658,N_3547);
nand U10848 (N_10848,N_3350,N_4259);
or U10849 (N_10849,N_2361,N_2158);
and U10850 (N_10850,N_3617,N_6018);
and U10851 (N_10851,N_8750,N_6280);
xnor U10852 (N_10852,N_4984,N_1357);
nor U10853 (N_10853,N_9744,N_8344);
nor U10854 (N_10854,N_9380,N_3895);
nor U10855 (N_10855,N_5290,N_553);
and U10856 (N_10856,N_9736,N_4847);
nor U10857 (N_10857,N_8679,N_5009);
nor U10858 (N_10858,N_1898,N_9277);
and U10859 (N_10859,N_8656,N_9218);
or U10860 (N_10860,N_3508,N_8637);
and U10861 (N_10861,N_3561,N_4113);
and U10862 (N_10862,N_1741,N_6707);
nand U10863 (N_10863,N_5966,N_2186);
and U10864 (N_10864,N_4992,N_3338);
xnor U10865 (N_10865,N_3107,N_7275);
nor U10866 (N_10866,N_3831,N_9636);
or U10867 (N_10867,N_9031,N_6432);
nor U10868 (N_10868,N_3781,N_3341);
nor U10869 (N_10869,N_9450,N_4563);
or U10870 (N_10870,N_9530,N_9999);
or U10871 (N_10871,N_7042,N_9264);
nand U10872 (N_10872,N_7836,N_3130);
nor U10873 (N_10873,N_7505,N_1698);
or U10874 (N_10874,N_2380,N_4906);
xor U10875 (N_10875,N_6955,N_8684);
and U10876 (N_10876,N_1618,N_8825);
nand U10877 (N_10877,N_6814,N_5969);
nor U10878 (N_10878,N_5694,N_52);
xnor U10879 (N_10879,N_8216,N_1017);
or U10880 (N_10880,N_3786,N_4316);
nand U10881 (N_10881,N_5094,N_9038);
xor U10882 (N_10882,N_4155,N_4953);
xor U10883 (N_10883,N_8607,N_1756);
nor U10884 (N_10884,N_9883,N_1726);
nor U10885 (N_10885,N_6790,N_1537);
nor U10886 (N_10886,N_2615,N_2379);
nand U10887 (N_10887,N_5346,N_1233);
xnor U10888 (N_10888,N_2832,N_1471);
or U10889 (N_10889,N_3447,N_501);
or U10890 (N_10890,N_4857,N_3613);
nor U10891 (N_10891,N_7309,N_7084);
nand U10892 (N_10892,N_4424,N_4496);
or U10893 (N_10893,N_5496,N_9142);
and U10894 (N_10894,N_1046,N_1752);
nor U10895 (N_10895,N_1324,N_2801);
and U10896 (N_10896,N_671,N_1275);
nand U10897 (N_10897,N_8044,N_3769);
nor U10898 (N_10898,N_9938,N_7509);
nand U10899 (N_10899,N_5432,N_8845);
or U10900 (N_10900,N_3223,N_1489);
xor U10901 (N_10901,N_7284,N_8531);
or U10902 (N_10902,N_354,N_1494);
xor U10903 (N_10903,N_5975,N_5917);
or U10904 (N_10904,N_9453,N_326);
or U10905 (N_10905,N_3239,N_9737);
nand U10906 (N_10906,N_8827,N_6674);
nor U10907 (N_10907,N_9711,N_9669);
and U10908 (N_10908,N_6795,N_3789);
nand U10909 (N_10909,N_2120,N_9660);
nand U10910 (N_10910,N_7753,N_2572);
and U10911 (N_10911,N_101,N_7233);
nor U10912 (N_10912,N_8250,N_9804);
nand U10913 (N_10913,N_1831,N_4761);
xnor U10914 (N_10914,N_9050,N_314);
nor U10915 (N_10915,N_5080,N_6316);
nor U10916 (N_10916,N_1210,N_9966);
nor U10917 (N_10917,N_8485,N_2333);
and U10918 (N_10918,N_3997,N_8024);
nand U10919 (N_10919,N_4512,N_2241);
or U10920 (N_10920,N_3858,N_4397);
nand U10921 (N_10921,N_2124,N_7754);
nand U10922 (N_10922,N_1911,N_2398);
and U10923 (N_10923,N_9183,N_2731);
and U10924 (N_10924,N_8418,N_3294);
nand U10925 (N_10925,N_9950,N_4792);
xor U10926 (N_10926,N_1298,N_5099);
nor U10927 (N_10927,N_7394,N_2037);
or U10928 (N_10928,N_5207,N_3047);
nor U10929 (N_10929,N_4212,N_7899);
nor U10930 (N_10930,N_921,N_1120);
nand U10931 (N_10931,N_2253,N_1319);
nand U10932 (N_10932,N_7727,N_8370);
xnor U10933 (N_10933,N_5899,N_6590);
nor U10934 (N_10934,N_1096,N_3327);
nand U10935 (N_10935,N_6067,N_3104);
xnor U10936 (N_10936,N_9045,N_3203);
nand U10937 (N_10937,N_4689,N_5985);
nor U10938 (N_10938,N_6129,N_480);
nor U10939 (N_10939,N_9214,N_1944);
and U10940 (N_10940,N_8615,N_8730);
nand U10941 (N_10941,N_2907,N_6812);
nand U10942 (N_10942,N_1859,N_5169);
or U10943 (N_10943,N_5286,N_1249);
nor U10944 (N_10944,N_9599,N_3913);
and U10945 (N_10945,N_1011,N_6480);
or U10946 (N_10946,N_3800,N_791);
xnor U10947 (N_10947,N_5319,N_479);
nor U10948 (N_10948,N_6402,N_3640);
and U10949 (N_10949,N_3407,N_7005);
and U10950 (N_10950,N_5584,N_3123);
xor U10951 (N_10951,N_9145,N_4979);
and U10952 (N_10952,N_8635,N_5764);
and U10953 (N_10953,N_4809,N_8308);
or U10954 (N_10954,N_449,N_6180);
nand U10955 (N_10955,N_3648,N_8342);
nor U10956 (N_10956,N_7124,N_7576);
nor U10957 (N_10957,N_4140,N_425);
or U10958 (N_10958,N_612,N_239);
xnor U10959 (N_10959,N_876,N_9313);
or U10960 (N_10960,N_7149,N_5670);
xnor U10961 (N_10961,N_4648,N_2450);
nor U10962 (N_10962,N_8739,N_6641);
or U10963 (N_10963,N_550,N_6123);
xor U10964 (N_10964,N_369,N_3684);
and U10965 (N_10965,N_6049,N_2771);
or U10966 (N_10966,N_4337,N_35);
xor U10967 (N_10967,N_5059,N_323);
nor U10968 (N_10968,N_5998,N_1071);
nor U10969 (N_10969,N_7051,N_9594);
and U10970 (N_10970,N_2302,N_8676);
xor U10971 (N_10971,N_3425,N_3468);
and U10972 (N_10972,N_9314,N_2870);
nor U10973 (N_10973,N_6910,N_7074);
or U10974 (N_10974,N_1122,N_413);
nand U10975 (N_10975,N_2222,N_3629);
or U10976 (N_10976,N_5117,N_2155);
or U10977 (N_10977,N_3225,N_706);
nor U10978 (N_10978,N_1526,N_4869);
or U10979 (N_10979,N_9877,N_1285);
and U10980 (N_10980,N_8160,N_6971);
xnor U10981 (N_10981,N_2568,N_4313);
or U10982 (N_10982,N_7700,N_8781);
and U10983 (N_10983,N_8864,N_2671);
nand U10984 (N_10984,N_6094,N_5376);
xor U10985 (N_10985,N_3559,N_8352);
or U10986 (N_10986,N_7876,N_2194);
xnor U10987 (N_10987,N_5879,N_7426);
or U10988 (N_10988,N_685,N_5026);
and U10989 (N_10989,N_5967,N_5033);
nor U10990 (N_10990,N_1916,N_3193);
xor U10991 (N_10991,N_1106,N_1195);
nor U10992 (N_10992,N_1697,N_1060);
and U10993 (N_10993,N_4639,N_8181);
or U10994 (N_10994,N_8629,N_2636);
nand U10995 (N_10995,N_5674,N_8788);
and U10996 (N_10996,N_5023,N_4144);
or U10997 (N_10997,N_7971,N_200);
and U10998 (N_10998,N_3604,N_2111);
and U10999 (N_10999,N_1412,N_7065);
nor U11000 (N_11000,N_9833,N_8754);
nand U11001 (N_11001,N_3227,N_2902);
or U11002 (N_11002,N_971,N_575);
and U11003 (N_11003,N_5104,N_6108);
and U11004 (N_11004,N_2356,N_2002);
nor U11005 (N_11005,N_917,N_4585);
and U11006 (N_11006,N_1320,N_9806);
or U11007 (N_11007,N_9265,N_9352);
or U11008 (N_11008,N_2336,N_8610);
nand U11009 (N_11009,N_1733,N_8267);
nor U11010 (N_11010,N_2695,N_9122);
and U11011 (N_11011,N_4538,N_4680);
xnor U11012 (N_11012,N_8358,N_3940);
and U11013 (N_11013,N_1220,N_2175);
nor U11014 (N_11014,N_4878,N_2228);
and U11015 (N_11015,N_5586,N_6082);
or U11016 (N_11016,N_8206,N_8584);
nor U11017 (N_11017,N_4860,N_8593);
and U11018 (N_11018,N_3980,N_5561);
nor U11019 (N_11019,N_1534,N_5492);
and U11020 (N_11020,N_1556,N_8016);
or U11021 (N_11021,N_7607,N_4966);
nand U11022 (N_11022,N_660,N_4562);
or U11023 (N_11023,N_3162,N_8810);
nand U11024 (N_11024,N_6585,N_7936);
nand U11025 (N_11025,N_9115,N_4416);
or U11026 (N_11026,N_2097,N_1196);
or U11027 (N_11027,N_5971,N_711);
or U11028 (N_11028,N_7845,N_6592);
nand U11029 (N_11029,N_3182,N_8043);
and U11030 (N_11030,N_5246,N_3697);
nand U11031 (N_11031,N_6211,N_8117);
nand U11032 (N_11032,N_4168,N_5128);
or U11033 (N_11033,N_176,N_3810);
or U11034 (N_11034,N_2013,N_3590);
and U11035 (N_11035,N_2115,N_5856);
nand U11036 (N_11036,N_1102,N_8743);
or U11037 (N_11037,N_8285,N_7765);
xnor U11038 (N_11038,N_315,N_1562);
and U11039 (N_11039,N_4954,N_271);
nand U11040 (N_11040,N_2800,N_5601);
and U11041 (N_11041,N_2863,N_2914);
nor U11042 (N_11042,N_4814,N_7422);
nor U11043 (N_11043,N_8122,N_1269);
nand U11044 (N_11044,N_4063,N_3032);
and U11045 (N_11045,N_6459,N_9674);
nor U11046 (N_11046,N_9911,N_1115);
nor U11047 (N_11047,N_2150,N_5545);
nor U11048 (N_11048,N_5562,N_9887);
nor U11049 (N_11049,N_5203,N_518);
or U11050 (N_11050,N_7735,N_6819);
and U11051 (N_11051,N_8292,N_3352);
nand U11052 (N_11052,N_5381,N_2034);
xor U11053 (N_11053,N_3360,N_431);
or U11054 (N_11054,N_1560,N_6193);
nor U11055 (N_11055,N_2126,N_9895);
xor U11056 (N_11056,N_7749,N_9459);
nand U11057 (N_11057,N_8929,N_4726);
or U11058 (N_11058,N_8057,N_2523);
nor U11059 (N_11059,N_8639,N_1533);
nor U11060 (N_11060,N_9200,N_9354);
or U11061 (N_11061,N_7348,N_7371);
nand U11062 (N_11062,N_1584,N_8848);
nor U11063 (N_11063,N_6079,N_1573);
nand U11064 (N_11064,N_8941,N_4029);
nor U11065 (N_11065,N_1361,N_5443);
nand U11066 (N_11066,N_4898,N_7273);
or U11067 (N_11067,N_9583,N_3116);
and U11068 (N_11068,N_6077,N_4519);
nand U11069 (N_11069,N_9298,N_8110);
and U11070 (N_11070,N_2500,N_4240);
nand U11071 (N_11071,N_9605,N_9622);
and U11072 (N_11072,N_9511,N_6347);
nor U11073 (N_11073,N_6901,N_2493);
and U11074 (N_11074,N_3917,N_5534);
nand U11075 (N_11075,N_8535,N_4108);
nand U11076 (N_11076,N_184,N_6490);
nor U11077 (N_11077,N_3060,N_1045);
and U11078 (N_11078,N_9410,N_741);
or U11079 (N_11079,N_1105,N_9526);
nor U11080 (N_11080,N_5046,N_8534);
nor U11081 (N_11081,N_3321,N_8917);
or U11082 (N_11082,N_5810,N_7539);
and U11083 (N_11083,N_7354,N_7593);
or U11084 (N_11084,N_2366,N_3660);
and U11085 (N_11085,N_3159,N_1744);
nor U11086 (N_11086,N_1798,N_175);
or U11087 (N_11087,N_4232,N_3675);
and U11088 (N_11088,N_6368,N_9805);
nor U11089 (N_11089,N_5772,N_6451);
or U11090 (N_11090,N_9187,N_7777);
nand U11091 (N_11091,N_5389,N_7142);
or U11092 (N_11092,N_8202,N_651);
or U11093 (N_11093,N_986,N_76);
nand U11094 (N_11094,N_1959,N_8697);
or U11095 (N_11095,N_7957,N_999);
or U11096 (N_11096,N_5478,N_4837);
or U11097 (N_11097,N_7838,N_8190);
nand U11098 (N_11098,N_6000,N_1570);
or U11099 (N_11099,N_5982,N_8163);
or U11100 (N_11100,N_7953,N_3989);
nor U11101 (N_11101,N_9378,N_805);
or U11102 (N_11102,N_5396,N_3091);
or U11103 (N_11103,N_9379,N_5593);
nand U11104 (N_11104,N_1388,N_2179);
or U11105 (N_11105,N_6978,N_9734);
nand U11106 (N_11106,N_1527,N_3456);
or U11107 (N_11107,N_6745,N_8218);
and U11108 (N_11108,N_7680,N_6818);
and U11109 (N_11109,N_8282,N_6113);
nand U11110 (N_11110,N_4803,N_7167);
nor U11111 (N_11111,N_7398,N_7071);
or U11112 (N_11112,N_991,N_6483);
and U11113 (N_11113,N_1951,N_2686);
or U11114 (N_11114,N_2821,N_8586);
and U11115 (N_11115,N_6377,N_1394);
and U11116 (N_11116,N_30,N_9514);
or U11117 (N_11117,N_9347,N_9284);
nor U11118 (N_11118,N_1614,N_4789);
or U11119 (N_11119,N_139,N_2634);
nor U11120 (N_11120,N_2534,N_5370);
or U11121 (N_11121,N_8387,N_5994);
or U11122 (N_11122,N_8838,N_5206);
and U11123 (N_11123,N_6474,N_1505);
or U11124 (N_11124,N_962,N_4064);
and U11125 (N_11125,N_772,N_4855);
or U11126 (N_11126,N_8530,N_4713);
and U11127 (N_11127,N_4447,N_5347);
and U11128 (N_11128,N_3932,N_4808);
and U11129 (N_11129,N_2630,N_5289);
nand U11130 (N_11130,N_5645,N_1631);
nor U11131 (N_11131,N_1429,N_3070);
nor U11132 (N_11132,N_6718,N_6408);
xnor U11133 (N_11133,N_1579,N_2621);
nand U11134 (N_11134,N_7252,N_5336);
or U11135 (N_11135,N_1040,N_7106);
xor U11136 (N_11136,N_6433,N_8091);
and U11137 (N_11137,N_8876,N_8326);
or U11138 (N_11138,N_6276,N_6216);
nand U11139 (N_11139,N_3711,N_552);
or U11140 (N_11140,N_1166,N_6159);
nor U11141 (N_11141,N_1875,N_2791);
xnor U11142 (N_11142,N_3677,N_9070);
and U11143 (N_11143,N_7742,N_9640);
or U11144 (N_11144,N_5153,N_2802);
or U11145 (N_11145,N_6540,N_2140);
nand U11146 (N_11146,N_3693,N_3065);
and U11147 (N_11147,N_5242,N_7466);
nor U11148 (N_11148,N_7821,N_8756);
nor U11149 (N_11149,N_8120,N_979);
nor U11150 (N_11150,N_2438,N_6275);
xnor U11151 (N_11151,N_815,N_8174);
or U11152 (N_11152,N_7947,N_7769);
nor U11153 (N_11153,N_1937,N_4564);
nand U11154 (N_11154,N_9305,N_3189);
nor U11155 (N_11155,N_8056,N_5227);
or U11156 (N_11156,N_4274,N_7375);
nor U11157 (N_11157,N_611,N_5566);
and U11158 (N_11158,N_3458,N_423);
or U11159 (N_11159,N_7468,N_9004);
nor U11160 (N_11160,N_9490,N_6153);
nor U11161 (N_11161,N_2589,N_5499);
or U11162 (N_11162,N_6242,N_2442);
nor U11163 (N_11163,N_8975,N_2182);
nor U11164 (N_11164,N_9067,N_5528);
and U11165 (N_11165,N_240,N_6878);
nor U11166 (N_11166,N_6853,N_4504);
and U11167 (N_11167,N_1293,N_9129);
nand U11168 (N_11168,N_3937,N_8042);
xor U11169 (N_11169,N_9584,N_6185);
xor U11170 (N_11170,N_2147,N_7472);
nand U11171 (N_11171,N_6740,N_3026);
and U11172 (N_11172,N_2319,N_3158);
nor U11173 (N_11173,N_4291,N_2767);
nor U11174 (N_11174,N_5573,N_1550);
or U11175 (N_11175,N_6484,N_9475);
and U11176 (N_11176,N_4891,N_7869);
nand U11177 (N_11177,N_3452,N_9704);
nand U11178 (N_11178,N_7951,N_7697);
nor U11179 (N_11179,N_6755,N_1098);
nor U11180 (N_11180,N_1772,N_814);
xnor U11181 (N_11181,N_538,N_330);
nand U11182 (N_11182,N_562,N_2745);
or U11183 (N_11183,N_7439,N_9369);
nand U11184 (N_11184,N_8899,N_9834);
or U11185 (N_11185,N_4207,N_9044);
or U11186 (N_11186,N_1895,N_374);
and U11187 (N_11187,N_4790,N_3402);
or U11188 (N_11188,N_5292,N_8219);
nand U11189 (N_11189,N_9391,N_9007);
nand U11190 (N_11190,N_4598,N_7701);
nand U11191 (N_11191,N_3586,N_5845);
nand U11192 (N_11192,N_9886,N_4425);
nor U11193 (N_11193,N_1848,N_889);
and U11194 (N_11194,N_1753,N_8086);
nor U11195 (N_11195,N_8458,N_1305);
xnor U11196 (N_11196,N_7564,N_3986);
xor U11197 (N_11197,N_7269,N_7883);
nand U11198 (N_11198,N_2689,N_5410);
or U11199 (N_11199,N_4476,N_70);
xnor U11200 (N_11200,N_4893,N_3455);
and U11201 (N_11201,N_1410,N_161);
nor U11202 (N_11202,N_5839,N_5536);
nand U11203 (N_11203,N_4164,N_8426);
nand U11204 (N_11204,N_4740,N_3312);
xor U11205 (N_11205,N_3206,N_5272);
or U11206 (N_11206,N_8926,N_1953);
or U11207 (N_11207,N_8011,N_5614);
nor U11208 (N_11208,N_6136,N_9537);
or U11209 (N_11209,N_8302,N_1224);
nor U11210 (N_11210,N_1171,N_2474);
nand U11211 (N_11211,N_6743,N_6306);
and U11212 (N_11212,N_462,N_5045);
xnor U11213 (N_11213,N_7997,N_4560);
nor U11214 (N_11214,N_5502,N_1691);
nor U11215 (N_11215,N_2769,N_4951);
nor U11216 (N_11216,N_4534,N_9143);
xnor U11217 (N_11217,N_7373,N_5477);
and U11218 (N_11218,N_5387,N_3720);
nor U11219 (N_11219,N_1343,N_300);
or U11220 (N_11220,N_6608,N_3068);
or U11221 (N_11221,N_4742,N_3221);
nor U11222 (N_11222,N_1425,N_8971);
or U11223 (N_11223,N_9900,N_1297);
nand U11224 (N_11224,N_5237,N_3798);
xnor U11225 (N_11225,N_7665,N_1980);
and U11226 (N_11226,N_7977,N_920);
or U11227 (N_11227,N_6494,N_3627);
nor U11228 (N_11228,N_3419,N_5064);
nor U11229 (N_11229,N_9971,N_2702);
nor U11230 (N_11230,N_9908,N_4694);
nand U11231 (N_11231,N_9653,N_4851);
nor U11232 (N_11232,N_9235,N_6547);
and U11233 (N_11233,N_2426,N_4426);
and U11234 (N_11234,N_2259,N_2399);
or U11235 (N_11235,N_4487,N_4621);
nand U11236 (N_11236,N_638,N_1479);
and U11237 (N_11237,N_3439,N_9847);
xnor U11238 (N_11238,N_48,N_5553);
xor U11239 (N_11239,N_7994,N_251);
and U11240 (N_11240,N_5803,N_752);
nor U11241 (N_11241,N_2322,N_5365);
nor U11242 (N_11242,N_9234,N_8562);
or U11243 (N_11243,N_5557,N_2941);
xor U11244 (N_11244,N_8522,N_6903);
nor U11245 (N_11245,N_8018,N_7327);
and U11246 (N_11246,N_5005,N_8475);
and U11247 (N_11247,N_9462,N_5926);
nor U11248 (N_11248,N_5797,N_7538);
and U11249 (N_11249,N_1379,N_1727);
nor U11250 (N_11250,N_3864,N_2999);
xor U11251 (N_11251,N_223,N_155);
nor U11252 (N_11252,N_731,N_5730);
nand U11253 (N_11253,N_3646,N_5540);
and U11254 (N_11254,N_4375,N_610);
nor U11255 (N_11255,N_8755,N_9240);
nor U11256 (N_11256,N_625,N_1760);
nand U11257 (N_11257,N_6148,N_9077);
nor U11258 (N_11258,N_5152,N_4097);
or U11259 (N_11259,N_6133,N_9905);
xnor U11260 (N_11260,N_9927,N_2550);
xor U11261 (N_11261,N_2898,N_4398);
and U11262 (N_11262,N_441,N_3013);
or U11263 (N_11263,N_7259,N_3363);
or U11264 (N_11264,N_4060,N_7270);
nand U11265 (N_11265,N_303,N_2463);
xnor U11266 (N_11266,N_8938,N_5397);
nand U11267 (N_11267,N_4543,N_7108);
and U11268 (N_11268,N_2773,N_539);
or U11269 (N_11269,N_6544,N_1431);
xnor U11270 (N_11270,N_8805,N_6258);
nand U11271 (N_11271,N_1932,N_8670);
nand U11272 (N_11272,N_4103,N_1568);
nand U11273 (N_11273,N_6422,N_1472);
xnor U11274 (N_11274,N_5337,N_2292);
and U11275 (N_11275,N_9343,N_1609);
or U11276 (N_11276,N_5313,N_370);
nor U11277 (N_11277,N_6657,N_515);
xnor U11278 (N_11278,N_181,N_7912);
xor U11279 (N_11279,N_7083,N_2942);
nor U11280 (N_11280,N_5241,N_7881);
or U11281 (N_11281,N_4644,N_7622);
and U11282 (N_11282,N_1294,N_8422);
and U11283 (N_11283,N_9280,N_619);
nand U11284 (N_11284,N_9250,N_3577);
xor U11285 (N_11285,N_6144,N_7470);
nand U11286 (N_11286,N_4730,N_455);
or U11287 (N_11287,N_3185,N_9780);
nor U11288 (N_11288,N_3934,N_2974);
or U11289 (N_11289,N_5426,N_1816);
xor U11290 (N_11290,N_4795,N_573);
and U11291 (N_11291,N_4363,N_5456);
or U11292 (N_11292,N_7101,N_5529);
nor U11293 (N_11293,N_2807,N_6526);
xnor U11294 (N_11294,N_3920,N_2090);
nand U11295 (N_11295,N_6072,N_1686);
nor U11296 (N_11296,N_8543,N_2433);
or U11297 (N_11297,N_785,N_4236);
nand U11298 (N_11298,N_9903,N_787);
nor U11299 (N_11299,N_9825,N_4234);
nor U11300 (N_11300,N_8982,N_8820);
and U11301 (N_11301,N_2691,N_494);
nor U11302 (N_11302,N_4571,N_412);
xor U11303 (N_11303,N_8693,N_9638);
or U11304 (N_11304,N_9271,N_9487);
and U11305 (N_11305,N_6691,N_3418);
nor U11306 (N_11306,N_2795,N_3002);
or U11307 (N_11307,N_9968,N_6908);
or U11308 (N_11308,N_1401,N_3622);
and U11309 (N_11309,N_2283,N_8489);
nor U11310 (N_11310,N_9715,N_3718);
and U11311 (N_11311,N_5110,N_7673);
and U11312 (N_11312,N_6115,N_8529);
or U11313 (N_11313,N_4178,N_3594);
and U11314 (N_11314,N_9628,N_5500);
and U11315 (N_11315,N_813,N_7687);
nor U11316 (N_11316,N_1518,N_2888);
nand U11317 (N_11317,N_4110,N_4793);
and U11318 (N_11318,N_7768,N_5997);
or U11319 (N_11319,N_5677,N_3400);
nor U11320 (N_11320,N_4629,N_7261);
xnor U11321 (N_11321,N_6884,N_1915);
or U11322 (N_11322,N_1353,N_7591);
nor U11323 (N_11323,N_476,N_8050);
nor U11324 (N_11324,N_2001,N_7481);
nand U11325 (N_11325,N_3218,N_3556);
nor U11326 (N_11326,N_8600,N_5977);
and U11327 (N_11327,N_6973,N_5777);
and U11328 (N_11328,N_7129,N_8511);
xnor U11329 (N_11329,N_6698,N_9128);
nor U11330 (N_11330,N_3606,N_3961);
or U11331 (N_11331,N_5680,N_2050);
or U11332 (N_11332,N_2991,N_1402);
xor U11333 (N_11333,N_4282,N_4591);
nand U11334 (N_11334,N_2440,N_8313);
nor U11335 (N_11335,N_8429,N_6245);
nand U11336 (N_11336,N_3818,N_9672);
nand U11337 (N_11337,N_4012,N_7503);
or U11338 (N_11338,N_64,N_3167);
and U11339 (N_11339,N_2619,N_259);
nor U11340 (N_11340,N_6044,N_5385);
nand U11341 (N_11341,N_9389,N_5352);
or U11342 (N_11342,N_1768,N_9033);
or U11343 (N_11343,N_520,N_555);
nor U11344 (N_11344,N_6080,N_2561);
nand U11345 (N_11345,N_8336,N_6934);
and U11346 (N_11346,N_2624,N_3126);
xnor U11347 (N_11347,N_616,N_4771);
nand U11348 (N_11348,N_5912,N_414);
and U11349 (N_11349,N_502,N_1033);
xnor U11350 (N_11350,N_3467,N_7287);
nor U11351 (N_11351,N_788,N_5789);
nor U11352 (N_11352,N_1799,N_6783);
nor U11353 (N_11353,N_132,N_7308);
nor U11354 (N_11354,N_3637,N_1095);
or U11355 (N_11355,N_7172,N_9160);
nand U11356 (N_11356,N_932,N_8015);
and U11357 (N_11357,N_6310,N_1963);
xor U11358 (N_11358,N_8506,N_4276);
nand U11359 (N_11359,N_6174,N_7527);
and U11360 (N_11360,N_903,N_5264);
nor U11361 (N_11361,N_8184,N_3025);
or U11362 (N_11362,N_1661,N_6170);
and U11363 (N_11363,N_2176,N_3854);
and U11364 (N_11364,N_3297,N_4072);
and U11365 (N_11365,N_8003,N_4298);
or U11366 (N_11366,N_670,N_3422);
nand U11367 (N_11367,N_6685,N_1611);
nand U11368 (N_11368,N_955,N_6613);
or U11369 (N_11369,N_6325,N_359);
and U11370 (N_11370,N_5701,N_9570);
and U11371 (N_11371,N_1368,N_4973);
and U11372 (N_11372,N_8587,N_3226);
and U11373 (N_11373,N_5113,N_1172);
and U11374 (N_11374,N_9699,N_6027);
or U11375 (N_11375,N_241,N_2740);
and U11376 (N_11376,N_4856,N_9727);
nand U11377 (N_11377,N_9566,N_5379);
and U11378 (N_11378,N_4570,N_7999);
nand U11379 (N_11379,N_4785,N_2808);
nand U11380 (N_11380,N_5341,N_2079);
or U11381 (N_11381,N_9576,N_4154);
nand U11382 (N_11382,N_580,N_5232);
and U11383 (N_11383,N_8521,N_317);
nand U11384 (N_11384,N_4226,N_1377);
nand U11385 (N_11385,N_2818,N_7804);
and U11386 (N_11386,N_5889,N_8075);
nand U11387 (N_11387,N_6196,N_2834);
xnor U11388 (N_11388,N_900,N_6720);
nor U11389 (N_11389,N_5648,N_6669);
nor U11390 (N_11390,N_943,N_3170);
nand U11391 (N_11391,N_6709,N_379);
or U11392 (N_11392,N_2161,N_6846);
and U11393 (N_11393,N_9483,N_4410);
or U11394 (N_11394,N_8185,N_6324);
or U11395 (N_11395,N_8244,N_1706);
nand U11396 (N_11396,N_7353,N_1180);
nand U11397 (N_11397,N_9438,N_5137);
nor U11398 (N_11398,N_8028,N_6979);
nand U11399 (N_11399,N_1164,N_9907);
or U11400 (N_11400,N_8608,N_5134);
nor U11401 (N_11401,N_1415,N_9997);
nand U11402 (N_11402,N_7246,N_18);
or U11403 (N_11403,N_6714,N_5603);
or U11404 (N_11404,N_6502,N_9428);
and U11405 (N_11405,N_8973,N_2035);
and U11406 (N_11406,N_8409,N_4854);
nor U11407 (N_11407,N_3234,N_6286);
nor U11408 (N_11408,N_8996,N_4150);
nand U11409 (N_11409,N_4364,N_46);
nor U11410 (N_11410,N_296,N_7650);
xnor U11411 (N_11411,N_8653,N_4018);
nand U11412 (N_11412,N_7964,N_1288);
nor U11413 (N_11413,N_3217,N_1918);
nor U11414 (N_11414,N_3737,N_1004);
and U11415 (N_11415,N_8312,N_5687);
or U11416 (N_11416,N_6587,N_2088);
or U11417 (N_11417,N_2191,N_9982);
nand U11418 (N_11418,N_2402,N_2058);
and U11419 (N_11419,N_8545,N_1785);
nand U11420 (N_11420,N_887,N_262);
xnor U11421 (N_11421,N_3918,N_3168);
or U11422 (N_11422,N_1054,N_1327);
nand U11423 (N_11423,N_8304,N_6667);
and U11424 (N_11424,N_8952,N_4907);
nor U11425 (N_11425,N_6931,N_5600);
nand U11426 (N_11426,N_8144,N_6595);
xnor U11427 (N_11427,N_104,N_2425);
xor U11428 (N_11428,N_6446,N_5287);
nand U11429 (N_11429,N_154,N_5509);
xnor U11430 (N_11430,N_4305,N_3673);
nand U11431 (N_11431,N_401,N_8194);
or U11432 (N_11432,N_7461,N_906);
xor U11433 (N_11433,N_463,N_405);
or U11434 (N_11434,N_1775,N_9012);
or U11435 (N_11435,N_497,N_8031);
nor U11436 (N_11436,N_5317,N_9479);
nand U11437 (N_11437,N_1109,N_1299);
and U11438 (N_11438,N_2968,N_436);
and U11439 (N_11439,N_1452,N_5011);
nand U11440 (N_11440,N_8137,N_2204);
and U11441 (N_11441,N_5848,N_8908);
or U11442 (N_11442,N_4661,N_2307);
and U11443 (N_11443,N_4258,N_9279);
nand U11444 (N_11444,N_7362,N_5469);
xnor U11445 (N_11445,N_3041,N_6683);
nand U11446 (N_11446,N_9246,N_4645);
xnor U11447 (N_11447,N_1998,N_3710);
and U11448 (N_11448,N_2217,N_8512);
nand U11449 (N_11449,N_9423,N_8514);
and U11450 (N_11450,N_2687,N_6975);
or U11451 (N_11451,N_3388,N_8183);
and U11452 (N_11452,N_5417,N_4392);
or U11453 (N_11453,N_6936,N_725);
nand U11454 (N_11454,N_833,N_2332);
nor U11455 (N_11455,N_7000,N_1574);
nand U11456 (N_11456,N_9559,N_7526);
or U11457 (N_11457,N_3928,N_334);
and U11458 (N_11458,N_7514,N_8891);
nand U11459 (N_11459,N_6320,N_7156);
nand U11460 (N_11460,N_7234,N_2857);
nor U11461 (N_11461,N_4626,N_3967);
nor U11462 (N_11462,N_5042,N_5544);
nor U11463 (N_11463,N_1354,N_4361);
xnor U11464 (N_11464,N_1222,N_6501);
nor U11465 (N_11465,N_3618,N_2107);
nand U11466 (N_11466,N_8779,N_6297);
or U11467 (N_11467,N_1173,N_410);
and U11468 (N_11468,N_5096,N_4215);
or U11469 (N_11469,N_4641,N_4602);
xnor U11470 (N_11470,N_7040,N_4433);
or U11471 (N_11471,N_7062,N_942);
and U11472 (N_11472,N_6246,N_1356);
nand U11473 (N_11473,N_9623,N_9084);
or U11474 (N_11474,N_391,N_8852);
or U11475 (N_11475,N_2471,N_102);
nand U11476 (N_11476,N_7574,N_8726);
and U11477 (N_11477,N_4666,N_4443);
nand U11478 (N_11478,N_1960,N_49);
nand U11479 (N_11479,N_8128,N_286);
and U11480 (N_11480,N_3036,N_7386);
nor U11481 (N_11481,N_25,N_9463);
nand U11482 (N_11482,N_8009,N_7675);
nor U11483 (N_11483,N_5653,N_1309);
nand U11484 (N_11484,N_1708,N_9650);
or U11485 (N_11485,N_8807,N_6821);
and U11486 (N_11486,N_4114,N_2726);
xor U11487 (N_11487,N_3846,N_3390);
xor U11488 (N_11488,N_7130,N_2008);
nand U11489 (N_11489,N_6343,N_7940);
or U11490 (N_11490,N_648,N_4622);
nor U11491 (N_11491,N_9422,N_778);
and U11492 (N_11492,N_9021,N_5395);
nor U11493 (N_11493,N_482,N_1359);
nor U11494 (N_11494,N_2738,N_6375);
nor U11495 (N_11495,N_4166,N_7995);
nand U11496 (N_11496,N_9551,N_2492);
nor U11497 (N_11497,N_9864,N_1462);
nor U11498 (N_11498,N_6257,N_1590);
nor U11499 (N_11499,N_3902,N_3194);
nand U11500 (N_11500,N_4393,N_4655);
nor U11501 (N_11501,N_6844,N_2961);
nor U11502 (N_11502,N_4455,N_8442);
and U11503 (N_11503,N_2169,N_7347);
nand U11504 (N_11504,N_235,N_7766);
nand U11505 (N_11505,N_1358,N_4545);
nand U11506 (N_11506,N_5111,N_8713);
or U11507 (N_11507,N_8909,N_3010);
nor U11508 (N_11508,N_1991,N_8734);
or U11509 (N_11509,N_6247,N_7298);
nand U11510 (N_11510,N_7747,N_6300);
nand U11511 (N_11511,N_6057,N_3145);
or U11512 (N_11512,N_2755,N_7193);
nor U11513 (N_11513,N_2367,N_1179);
nor U11514 (N_11514,N_9621,N_1626);
nor U11515 (N_11515,N_4921,N_1828);
or U11516 (N_11516,N_6938,N_9182);
xnor U11517 (N_11517,N_9089,N_2900);
and U11518 (N_11518,N_5390,N_8212);
and U11519 (N_11519,N_2014,N_1949);
and U11520 (N_11520,N_1456,N_964);
and U11521 (N_11521,N_8054,N_2087);
nand U11522 (N_11522,N_8316,N_9190);
nor U11523 (N_11523,N_4510,N_4438);
nand U11524 (N_11524,N_6374,N_5180);
nand U11525 (N_11525,N_1080,N_1321);
nand U11526 (N_11526,N_9436,N_6887);
and U11527 (N_11527,N_5514,N_6226);
nand U11528 (N_11528,N_1234,N_3374);
nand U11529 (N_11529,N_2552,N_911);
or U11530 (N_11530,N_4864,N_4632);
and U11531 (N_11531,N_6361,N_969);
or U11532 (N_11532,N_4747,N_9274);
and U11533 (N_11533,N_8251,N_4451);
nand U11534 (N_11534,N_965,N_444);
nand U11535 (N_11535,N_3131,N_7490);
or U11536 (N_11536,N_4539,N_3909);
and U11537 (N_11537,N_1390,N_2683);
and U11538 (N_11538,N_9574,N_7073);
and U11539 (N_11539,N_9840,N_7518);
xor U11540 (N_11540,N_1841,N_6205);
nand U11541 (N_11541,N_8192,N_3949);
xnor U11542 (N_11542,N_1729,N_1083);
or U11543 (N_11543,N_3238,N_7184);
nor U11544 (N_11544,N_8055,N_7068);
nand U11545 (N_11545,N_4928,N_7849);
nand U11546 (N_11546,N_3253,N_2963);
and U11547 (N_11547,N_9242,N_128);
and U11548 (N_11548,N_261,N_4422);
xor U11549 (N_11549,N_5312,N_6175);
xor U11550 (N_11550,N_3389,N_3144);
nand U11551 (N_11551,N_73,N_1281);
nor U11552 (N_11552,N_6635,N_5421);
nand U11553 (N_11553,N_1100,N_4870);
nor U11554 (N_11554,N_4940,N_9081);
or U11555 (N_11555,N_396,N_4677);
and U11556 (N_11556,N_3578,N_9446);
or U11557 (N_11557,N_8245,N_8722);
nand U11558 (N_11558,N_4478,N_5000);
nor U11559 (N_11559,N_2559,N_7095);
xor U11560 (N_11560,N_1564,N_2108);
nor U11561 (N_11561,N_2623,N_9528);
nor U11562 (N_11562,N_3861,N_6291);
nand U11563 (N_11563,N_7898,N_9926);
or U11564 (N_11564,N_459,N_8369);
or U11565 (N_11565,N_8552,N_8537);
and U11566 (N_11566,N_5794,N_2285);
and U11567 (N_11567,N_3632,N_9057);
and U11568 (N_11568,N_5494,N_188);
and U11569 (N_11569,N_4711,N_9754);
xnor U11570 (N_11570,N_6551,N_9415);
nor U11571 (N_11571,N_2886,N_5419);
nand U11572 (N_11572,N_8618,N_1197);
and U11573 (N_11573,N_3783,N_7198);
nand U11574 (N_11574,N_5269,N_3289);
nand U11575 (N_11575,N_7546,N_9874);
nor U11576 (N_11576,N_7502,N_6771);
nor U11577 (N_11577,N_6582,N_5455);
and U11578 (N_11578,N_6011,N_5123);
and U11579 (N_11579,N_2200,N_8794);
nand U11580 (N_11580,N_3187,N_1277);
nor U11581 (N_11581,N_2694,N_2360);
nor U11582 (N_11582,N_849,N_3284);
xnor U11583 (N_11583,N_3544,N_1954);
and U11584 (N_11584,N_6776,N_2799);
and U11585 (N_11585,N_9294,N_6987);
or U11586 (N_11586,N_9586,N_3748);
nand U11587 (N_11587,N_7037,N_8987);
nor U11588 (N_11588,N_3688,N_3820);
nor U11589 (N_11589,N_9216,N_9978);
nor U11590 (N_11590,N_2517,N_4147);
nor U11591 (N_11591,N_4948,N_16);
xnor U11592 (N_11592,N_3393,N_6372);
nor U11593 (N_11593,N_9427,N_1110);
nand U11594 (N_11594,N_7853,N_7003);
and U11595 (N_11595,N_3517,N_4373);
or U11596 (N_11596,N_1627,N_5724);
xor U11597 (N_11597,N_790,N_9875);
nand U11598 (N_11598,N_7242,N_7109);
nand U11599 (N_11599,N_8125,N_5970);
or U11600 (N_11600,N_3022,N_6725);
and U11601 (N_11601,N_9041,N_4670);
and U11602 (N_11602,N_7559,N_4737);
and U11603 (N_11603,N_4876,N_4634);
xnor U11604 (N_11604,N_8927,N_3128);
nand U11605 (N_11605,N_489,N_7557);
nand U11606 (N_11606,N_8196,N_7577);
nor U11607 (N_11607,N_5165,N_6549);
and U11608 (N_11608,N_5865,N_9773);
and U11609 (N_11609,N_5834,N_5542);
nand U11610 (N_11610,N_8207,N_3933);
or U11611 (N_11611,N_2345,N_2141);
and U11612 (N_11612,N_8463,N_6970);
and U11613 (N_11613,N_3730,N_6741);
or U11614 (N_11614,N_7244,N_7854);
nand U11615 (N_11615,N_9032,N_116);
xor U11616 (N_11616,N_1587,N_633);
or U11617 (N_11617,N_8325,N_4090);
nand U11618 (N_11618,N_5638,N_9706);
nand U11619 (N_11619,N_6183,N_5329);
and U11620 (N_11620,N_7895,N_9517);
nand U11621 (N_11621,N_6288,N_1237);
nor U11622 (N_11622,N_9569,N_3663);
nor U11623 (N_11623,N_4769,N_2718);
or U11624 (N_11624,N_8095,N_4619);
xnor U11625 (N_11625,N_8525,N_5200);
nand U11626 (N_11626,N_2997,N_8621);
or U11627 (N_11627,N_5457,N_7980);
nand U11628 (N_11628,N_2666,N_9452);
xnor U11629 (N_11629,N_2173,N_2539);
nand U11630 (N_11630,N_956,N_6272);
and U11631 (N_11631,N_2383,N_4290);
nor U11632 (N_11632,N_7987,N_7063);
and U11633 (N_11633,N_5268,N_7782);
nor U11634 (N_11634,N_9467,N_3553);
nor U11635 (N_11635,N_600,N_4061);
or U11636 (N_11636,N_3816,N_8017);
and U11637 (N_11637,N_3657,N_9220);
nand U11638 (N_11638,N_3135,N_4277);
nor U11639 (N_11639,N_7180,N_3801);
or U11640 (N_11640,N_8865,N_2201);
nand U11641 (N_11641,N_6099,N_3277);
nor U11642 (N_11642,N_4163,N_7164);
and U11643 (N_11643,N_45,N_9470);
nand U11644 (N_11644,N_9206,N_7477);
or U11645 (N_11645,N_2390,N_3658);
nor U11646 (N_11646,N_4909,N_2193);
nor U11647 (N_11647,N_4692,N_419);
or U11648 (N_11648,N_2223,N_645);
and U11649 (N_11649,N_6530,N_8564);
or U11650 (N_11650,N_5888,N_5183);
nor U11651 (N_11651,N_2106,N_9105);
nor U11652 (N_11652,N_352,N_9093);
or U11653 (N_11653,N_4962,N_913);
nand U11654 (N_11654,N_7206,N_4839);
xnor U11655 (N_11655,N_1771,N_9692);
or U11656 (N_11656,N_8111,N_7022);
and U11657 (N_11657,N_5597,N_7201);
nor U11658 (N_11658,N_1683,N_1672);
xnor U11659 (N_11659,N_5718,N_8898);
and U11660 (N_11660,N_7311,N_5642);
nand U11661 (N_11661,N_9819,N_6673);
xor U11662 (N_11662,N_1792,N_7615);
and U11663 (N_11663,N_1942,N_546);
or U11664 (N_11664,N_3444,N_4262);
and U11665 (N_11665,N_5588,N_7310);
xnor U11666 (N_11666,N_7879,N_6571);
nor U11667 (N_11667,N_5156,N_934);
or U11668 (N_11668,N_2547,N_2294);
nor U11669 (N_11669,N_1130,N_543);
nand U11670 (N_11670,N_2255,N_618);
and U11671 (N_11671,N_4727,N_6337);
xor U11672 (N_11672,N_9456,N_6078);
xnor U11673 (N_11673,N_1050,N_7606);
and U11674 (N_11674,N_2591,N_7049);
nor U11675 (N_11675,N_8832,N_269);
nor U11676 (N_11676,N_6263,N_1779);
nor U11677 (N_11677,N_5522,N_6882);
or U11678 (N_11678,N_4203,N_767);
xor U11679 (N_11679,N_5109,N_8652);
xor U11680 (N_11680,N_5806,N_6309);
nor U11681 (N_11681,N_8098,N_350);
nand U11682 (N_11682,N_7868,N_1777);
nand U11683 (N_11683,N_6478,N_9014);
nand U11684 (N_11684,N_3886,N_8712);
nand U11685 (N_11685,N_5673,N_8767);
or U11686 (N_11686,N_5826,N_1877);
nor U11687 (N_11687,N_8826,N_7044);
nor U11688 (N_11688,N_4332,N_5074);
or U11689 (N_11689,N_3034,N_7657);
nand U11690 (N_11690,N_9263,N_6815);
nand U11691 (N_11691,N_4448,N_6321);
or U11692 (N_11692,N_9247,N_1464);
and U11693 (N_11693,N_3630,N_2697);
or U11694 (N_11694,N_8256,N_7341);
or U11695 (N_11695,N_4759,N_584);
nor U11696 (N_11696,N_9633,N_676);
or U11697 (N_11697,N_8252,N_9170);
and U11698 (N_11698,N_3963,N_4340);
nand U11699 (N_11699,N_157,N_4270);
nor U11700 (N_11700,N_8069,N_6384);
nand U11701 (N_11701,N_8613,N_9469);
nand U11702 (N_11702,N_4248,N_9310);
xor U11703 (N_11703,N_9028,N_4505);
nor U11704 (N_11704,N_893,N_4370);
or U11705 (N_11705,N_7759,N_854);
nor U11706 (N_11706,N_4239,N_15);
or U11707 (N_11707,N_4273,N_7225);
or U11708 (N_11708,N_7295,N_2076);
or U11709 (N_11709,N_3469,N_789);
and U11710 (N_11710,N_5098,N_4985);
or U11711 (N_11711,N_1308,N_380);
or U11712 (N_11712,N_3725,N_6676);
xnor U11713 (N_11713,N_797,N_6927);
nand U11714 (N_11714,N_2449,N_3722);
and U11715 (N_11715,N_247,N_9850);
or U11716 (N_11716,N_5855,N_2701);
xnor U11717 (N_11717,N_5446,N_5753);
and U11718 (N_11718,N_2007,N_6508);
nor U11719 (N_11719,N_6584,N_7015);
or U11720 (N_11720,N_6329,N_3330);
or U11721 (N_11721,N_3878,N_9611);
and U11722 (N_11722,N_2954,N_4008);
and U11723 (N_11723,N_9860,N_2569);
or U11724 (N_11724,N_9562,N_5807);
and U11725 (N_11725,N_2095,N_7196);
nand U11726 (N_11726,N_847,N_2198);
or U11727 (N_11727,N_3283,N_1531);
nand U11728 (N_11728,N_3133,N_8276);
or U11729 (N_11729,N_3531,N_8423);
or U11730 (N_11730,N_7012,N_7866);
and U11731 (N_11731,N_6002,N_9667);
xor U11732 (N_11732,N_3383,N_923);
nand U11733 (N_11733,N_4915,N_7667);
nand U11734 (N_11734,N_8960,N_4965);
nand U11735 (N_11735,N_6605,N_1022);
or U11736 (N_11736,N_6085,N_7604);
and U11737 (N_11737,N_7939,N_4494);
and U11738 (N_11738,N_740,N_2148);
nand U11739 (N_11739,N_384,N_1693);
and U11740 (N_11740,N_8979,N_6131);
or U11741 (N_11741,N_8888,N_5922);
or U11742 (N_11742,N_1091,N_2230);
nand U11743 (N_11743,N_8777,N_4319);
nand U11744 (N_11744,N_8260,N_3992);
or U11745 (N_11745,N_1304,N_3230);
and U11746 (N_11746,N_7195,N_2545);
xor U11747 (N_11747,N_1640,N_2221);
nand U11748 (N_11748,N_4025,N_5854);
nand U11749 (N_11749,N_6896,N_5925);
and U11750 (N_11750,N_8583,N_5795);
nor U11751 (N_11751,N_4081,N_4134);
and U11752 (N_11752,N_8356,N_7);
and U11753 (N_11753,N_429,N_5220);
nor U11754 (N_11754,N_4611,N_2597);
nand U11755 (N_11755,N_8920,N_1311);
or U11756 (N_11756,N_1006,N_8156);
and U11757 (N_11757,N_528,N_5893);
xor U11758 (N_11758,N_5038,N_321);
and U11759 (N_11759,N_3424,N_9603);
or U11760 (N_11760,N_475,N_193);
nand U11761 (N_11761,N_9928,N_17);
xor U11762 (N_11762,N_9262,N_5990);
and U11763 (N_11763,N_4450,N_4312);
nor U11764 (N_11764,N_6442,N_5436);
nor U11765 (N_11765,N_3978,N_3567);
xnor U11766 (N_11766,N_6045,N_7504);
and U11767 (N_11767,N_8978,N_7706);
nor U11768 (N_11768,N_1598,N_5008);
nor U11769 (N_11769,N_7222,N_4681);
and U11770 (N_11770,N_3753,N_5427);
nand U11771 (N_11771,N_4660,N_331);
nor U11772 (N_11772,N_5537,N_5862);
or U11773 (N_11773,N_9523,N_6059);
and U11774 (N_11774,N_3038,N_31);
and U11775 (N_11775,N_1082,N_4022);
and U11776 (N_11776,N_7415,N_8170);
nand U11777 (N_11777,N_659,N_3115);
and U11778 (N_11778,N_1141,N_5465);
xor U11779 (N_11779,N_5483,N_1759);
or U11780 (N_11780,N_3736,N_9385);
or U11781 (N_11781,N_1667,N_9590);
nand U11782 (N_11782,N_4703,N_1972);
nand U11783 (N_11783,N_8172,N_8849);
nand U11784 (N_11784,N_1596,N_3707);
nor U11785 (N_11785,N_1331,N_5755);
nor U11786 (N_11786,N_5626,N_355);
nor U11787 (N_11787,N_1887,N_9593);
and U11788 (N_11788,N_2549,N_5072);
or U11789 (N_11789,N_8427,N_1364);
nor U11790 (N_11790,N_8078,N_2514);
xnor U11791 (N_11791,N_7739,N_8448);
and U11792 (N_11792,N_9137,N_2117);
nor U11793 (N_11793,N_6435,N_7031);
nand U11794 (N_11794,N_1599,N_9685);
and U11795 (N_11795,N_474,N_6775);
nor U11796 (N_11796,N_6737,N_6829);
and U11797 (N_11797,N_392,N_7447);
or U11798 (N_11798,N_7787,N_4943);
or U11799 (N_11799,N_80,N_7788);
or U11800 (N_11800,N_1400,N_702);
nor U11801 (N_11801,N_6917,N_963);
or U11802 (N_11802,N_3479,N_3644);
nor U11803 (N_11803,N_66,N_8173);
and U11804 (N_11804,N_1348,N_3176);
and U11805 (N_11805,N_827,N_8603);
nand U11806 (N_11806,N_3392,N_4848);
or U11807 (N_11807,N_5799,N_6164);
and U11808 (N_11808,N_1235,N_1866);
nand U11809 (N_11809,N_4675,N_9931);
and U11810 (N_11810,N_4787,N_3763);
nor U11811 (N_11811,N_4032,N_3829);
nor U11812 (N_11812,N_1374,N_3319);
nor U11813 (N_11813,N_8472,N_1844);
nand U11814 (N_11814,N_9873,N_4308);
nand U11815 (N_11815,N_7026,N_7880);
or U11816 (N_11816,N_7264,N_3843);
nand U11817 (N_11817,N_4286,N_4379);
nor U11818 (N_11818,N_3521,N_2727);
nand U11819 (N_11819,N_9821,N_2504);
nor U11820 (N_11820,N_7575,N_1939);
xor U11821 (N_11821,N_5355,N_1232);
or U11822 (N_11822,N_7133,N_4229);
nor U11823 (N_11823,N_4446,N_129);
or U11824 (N_11824,N_8087,N_6929);
xor U11825 (N_11825,N_3639,N_6719);
nor U11826 (N_11826,N_5430,N_9949);
or U11827 (N_11827,N_5792,N_1520);
and U11828 (N_11828,N_9619,N_1968);
xnor U11829 (N_11829,N_2068,N_4272);
and U11830 (N_11830,N_5409,N_5366);
xor U11831 (N_11831,N_9906,N_4049);
nand U11832 (N_11832,N_4542,N_9579);
nor U11833 (N_11833,N_9196,N_5818);
or U11834 (N_11834,N_6062,N_7825);
or U11835 (N_11835,N_7385,N_7010);
nor U11836 (N_11836,N_6933,N_5354);
or U11837 (N_11837,N_7173,N_6071);
or U11838 (N_11838,N_9213,N_3347);
and U11839 (N_11839,N_8800,N_915);
and U11840 (N_11840,N_6188,N_43);
nand U11841 (N_11841,N_9756,N_4706);
xor U11842 (N_11842,N_7813,N_5022);
and U11843 (N_11843,N_5570,N_6731);
nor U11844 (N_11844,N_7493,N_9760);
and U11845 (N_11845,N_6659,N_6863);
or U11846 (N_11846,N_2925,N_1863);
and U11847 (N_11847,N_8362,N_5233);
or U11848 (N_11848,N_2780,N_8706);
nor U11849 (N_11849,N_169,N_1592);
and U11850 (N_11850,N_2480,N_689);
nand U11851 (N_11851,N_7949,N_9970);
or U11852 (N_11852,N_5219,N_3033);
nand U11853 (N_11853,N_7691,N_7534);
and U11854 (N_11854,N_4535,N_4124);
and U11855 (N_11855,N_5411,N_5987);
xnor U11856 (N_11856,N_8870,N_6777);
nand U11857 (N_11857,N_733,N_9769);
and U11858 (N_11858,N_6065,N_8605);
nor U11859 (N_11859,N_560,N_4117);
nand U11860 (N_11860,N_2043,N_7623);
or U11861 (N_11861,N_3680,N_9859);
nand U11862 (N_11862,N_4729,N_1170);
and U11863 (N_11863,N_6642,N_94);
nand U11864 (N_11864,N_5558,N_1515);
or U11865 (N_11865,N_7570,N_1207);
or U11866 (N_11866,N_8885,N_5727);
nor U11867 (N_11867,N_6625,N_4177);
nand U11868 (N_11868,N_5860,N_6350);
nor U11869 (N_11869,N_8919,N_6849);
nor U11870 (N_11870,N_1221,N_8523);
xnor U11871 (N_11871,N_90,N_5262);
nor U11872 (N_11872,N_8279,N_238);
xor U11873 (N_11873,N_28,N_9786);
and U11874 (N_11874,N_6466,N_2779);
nor U11875 (N_11875,N_5988,N_3848);
nor U11876 (N_11876,N_5733,N_7544);
nor U11877 (N_11877,N_7889,N_6318);
or U11878 (N_11878,N_8857,N_6261);
nand U11879 (N_11879,N_1290,N_4802);
nand U11880 (N_11880,N_6168,N_6330);
nor U11881 (N_11881,N_2633,N_1455);
nor U11882 (N_11882,N_5782,N_7113);
and U11883 (N_11883,N_9025,N_7826);
or U11884 (N_11884,N_8517,N_748);
or U11885 (N_11885,N_8263,N_7567);
nand U11886 (N_11886,N_198,N_3481);
or U11887 (N_11887,N_1849,N_9752);
nor U11888 (N_11888,N_6431,N_1934);
nor U11889 (N_11889,N_7799,N_433);
and U11890 (N_11890,N_9955,N_3470);
nand U11891 (N_11891,N_8483,N_1465);
nor U11892 (N_11892,N_2271,N_7828);
nand U11893 (N_11893,N_1503,N_571);
or U11894 (N_11894,N_5191,N_8962);
nor U11895 (N_11895,N_694,N_7609);
nand U11896 (N_11896,N_7923,N_2371);
nor U11897 (N_11897,N_9202,N_3735);
and U11898 (N_11898,N_6860,N_4148);
and U11899 (N_11899,N_224,N_1078);
nand U11900 (N_11900,N_2542,N_1964);
nand U11901 (N_11901,N_9447,N_8923);
nand U11902 (N_11902,N_2511,N_607);
or U11903 (N_11903,N_8271,N_2601);
or U11904 (N_11904,N_6964,N_2809);
nand U11905 (N_11905,N_8301,N_1809);
and U11906 (N_11906,N_3406,N_2413);
and U11907 (N_11907,N_8695,N_2434);
and U11908 (N_11908,N_3713,N_9915);
or U11909 (N_11909,N_4462,N_3367);
nand U11910 (N_11910,N_2214,N_8264);
nor U11911 (N_11911,N_9803,N_4432);
or U11912 (N_11912,N_9902,N_718);
xnor U11913 (N_11913,N_7655,N_1594);
xnor U11914 (N_11914,N_9163,N_372);
or U11915 (N_11915,N_4174,N_7021);
xnor U11916 (N_11916,N_432,N_8683);
xor U11917 (N_11917,N_6661,N_2923);
or U11918 (N_11918,N_4687,N_1839);
nor U11919 (N_11919,N_8678,N_3326);
nor U11920 (N_11920,N_2839,N_2607);
xor U11921 (N_11921,N_6120,N_8052);
or U11922 (N_11922,N_6036,N_2424);
and U11923 (N_11923,N_968,N_260);
or U11924 (N_11924,N_3235,N_9691);
or U11925 (N_11925,N_8080,N_3954);
nor U11926 (N_11926,N_8224,N_7670);
or U11927 (N_11927,N_508,N_1990);
nor U11928 (N_11928,N_8776,N_8936);
nor U11929 (N_11929,N_2721,N_3634);
nand U11930 (N_11930,N_9743,N_1449);
and U11931 (N_11931,N_2676,N_5027);
nor U11932 (N_11932,N_7265,N_4094);
or U11933 (N_11933,N_5866,N_9639);
or U11934 (N_11934,N_9489,N_290);
xnor U11935 (N_11935,N_5986,N_9558);
and U11936 (N_11936,N_7862,N_5245);
or U11937 (N_11937,N_6340,N_720);
and U11938 (N_11938,N_381,N_1351);
or U11939 (N_11939,N_319,N_1251);
nand U11940 (N_11940,N_8994,N_7299);
or U11941 (N_11941,N_3056,N_7601);
nand U11942 (N_11942,N_9580,N_2508);
and U11943 (N_11943,N_793,N_9946);
nand U11944 (N_11944,N_8132,N_697);
or U11945 (N_11945,N_9600,N_58);
and U11946 (N_11946,N_3828,N_7379);
or U11947 (N_11947,N_8784,N_8269);
xor U11948 (N_11948,N_1619,N_8167);
nand U11949 (N_11949,N_1212,N_3969);
nand U11950 (N_11950,N_1018,N_591);
or U11951 (N_11951,N_3662,N_2717);
xnor U11952 (N_11952,N_1981,N_7030);
nor U11953 (N_11953,N_1901,N_5142);
nor U11954 (N_11954,N_9572,N_445);
and U11955 (N_11955,N_3527,N_1422);
or U11956 (N_11956,N_5399,N_2077);
nand U11957 (N_11957,N_51,N_6985);
and U11958 (N_11958,N_4423,N_1403);
nor U11959 (N_11959,N_535,N_452);
nand U11960 (N_11960,N_9054,N_9356);
or U11961 (N_11961,N_6905,N_3797);
or U11962 (N_11962,N_9789,N_4162);
or U11963 (N_11963,N_8076,N_1135);
nor U11964 (N_11964,N_3000,N_2910);
and U11965 (N_11965,N_7920,N_4958);
and U11966 (N_11966,N_7404,N_4801);
nand U11967 (N_11967,N_2528,N_7412);
nand U11968 (N_11968,N_7852,N_7551);
nand U11969 (N_11969,N_759,N_1740);
nand U11970 (N_11970,N_7979,N_2915);
xnor U11971 (N_11971,N_2692,N_3331);
or U11972 (N_11972,N_9538,N_8067);
xor U11973 (N_11973,N_7757,N_2710);
and U11974 (N_11974,N_2286,N_3050);
nor U11975 (N_11975,N_4047,N_1833);
or U11976 (N_11976,N_3592,N_54);
nand U11977 (N_11977,N_7408,N_8675);
and U11978 (N_11978,N_3397,N_7712);
nand U11979 (N_11979,N_7967,N_810);
and U11980 (N_11980,N_1340,N_7767);
nand U11981 (N_11981,N_6675,N_5652);
or U11982 (N_11982,N_8763,N_9164);
and U11983 (N_11983,N_8393,N_4129);
nor U11984 (N_11984,N_9458,N_3074);
nor U11985 (N_11985,N_1715,N_2503);
nand U11986 (N_11986,N_2432,N_9287);
or U11987 (N_11987,N_9003,N_9124);
and U11988 (N_11988,N_9719,N_9377);
and U11989 (N_11989,N_307,N_1705);
or U11990 (N_11990,N_2218,N_9155);
and U11991 (N_11991,N_1803,N_1666);
nor U11992 (N_11992,N_5470,N_8573);
or U11993 (N_11993,N_6747,N_2987);
nand U11994 (N_11994,N_5338,N_2642);
and U11995 (N_11995,N_8317,N_295);
nor U11996 (N_11996,N_2714,N_309);
and U11997 (N_11997,N_390,N_6389);
nand U11998 (N_11998,N_9334,N_8915);
nand U11999 (N_11999,N_1765,N_6456);
or U12000 (N_12000,N_7332,N_1935);
nand U12001 (N_12001,N_4297,N_7690);
and U12002 (N_12002,N_9365,N_1889);
or U12003 (N_12003,N_2278,N_1876);
or U12004 (N_12004,N_8619,N_7714);
or U12005 (N_12005,N_1009,N_5047);
nand U12006 (N_12006,N_6505,N_3154);
xor U12007 (N_12007,N_5904,N_6026);
xnor U12008 (N_12008,N_7016,N_2973);
nand U12009 (N_12009,N_3728,N_9413);
xor U12010 (N_12010,N_8907,N_9668);
or U12011 (N_12011,N_7723,N_5742);
nor U12012 (N_12012,N_2396,N_3057);
nand U12013 (N_12013,N_2937,N_6873);
or U12014 (N_12014,N_9901,N_9110);
nand U12015 (N_12015,N_5720,N_3809);
nor U12016 (N_12016,N_9497,N_2439);
and U12017 (N_12017,N_3826,N_4770);
nor U12018 (N_12018,N_8972,N_905);
nor U12019 (N_12019,N_5632,N_776);
and U12020 (N_12020,N_124,N_83);
nor U12021 (N_12021,N_1260,N_1426);
nand U12022 (N_12022,N_8437,N_5097);
xor U12023 (N_12023,N_2890,N_6798);
or U12024 (N_12024,N_2293,N_884);
or U12025 (N_12025,N_3876,N_5857);
xor U12026 (N_12026,N_9899,N_2563);
nor U12027 (N_12027,N_9689,N_3633);
nor U12028 (N_12028,N_9185,N_6187);
and U12029 (N_12029,N_8918,N_9690);
or U12030 (N_12030,N_1871,N_5688);
nor U12031 (N_12031,N_5523,N_7338);
nand U12032 (N_12032,N_7517,N_297);
nor U12033 (N_12033,N_7930,N_8785);
nor U12034 (N_12034,N_4616,N_179);
or U12035 (N_12035,N_6332,N_2981);
nand U12036 (N_12036,N_6506,N_3795);
and U12037 (N_12037,N_5946,N_9370);
nor U12038 (N_12038,N_3990,N_3208);
nor U12039 (N_12039,N_3232,N_8601);
nand U12040 (N_12040,N_2586,N_3503);
nand U12041 (N_12041,N_5710,N_9948);
nor U12042 (N_12042,N_6161,N_8551);
and U12043 (N_12043,N_8488,N_1743);
and U12044 (N_12044,N_747,N_2153);
and U12045 (N_12045,N_8990,N_3667);
nand U12046 (N_12046,N_2019,N_7790);
nand U12047 (N_12047,N_2325,N_1711);
and U12048 (N_12048,N_9096,N_1823);
nand U12049 (N_12049,N_8354,N_8942);
and U12050 (N_12050,N_3946,N_7671);
nand U12051 (N_12051,N_1617,N_2524);
nor U12052 (N_12052,N_6897,N_6283);
nor U12053 (N_12053,N_5513,N_142);
or U12054 (N_12054,N_2994,N_7784);
nand U12055 (N_12055,N_3944,N_1019);
nand U12056 (N_12056,N_6953,N_9329);
nand U12057 (N_12057,N_3489,N_8666);
and U12058 (N_12058,N_1566,N_6952);
nor U12059 (N_12059,N_4368,N_7554);
and U12060 (N_12060,N_3446,N_2943);
nor U12061 (N_12061,N_6763,N_861);
and U12062 (N_12062,N_7168,N_2889);
or U12063 (N_12063,N_665,N_178);
nand U12064 (N_12064,N_2421,N_5585);
nor U12065 (N_12065,N_5579,N_526);
and U12066 (N_12066,N_9276,N_6778);
nor U12067 (N_12067,N_7356,N_9720);
xor U12068 (N_12068,N_1652,N_1433);
xor U12069 (N_12069,N_324,N_6839);
nand U12070 (N_12070,N_6277,N_4265);
xnor U12071 (N_12071,N_9282,N_9921);
xor U12072 (N_12072,N_5284,N_2541);
and U12073 (N_12073,N_6016,N_7581);
xor U12074 (N_12074,N_7166,N_427);
nor U12075 (N_12075,N_6504,N_3832);
xnor U12076 (N_12076,N_9856,N_8883);
nor U12077 (N_12077,N_8331,N_7663);
and U12078 (N_12078,N_2374,N_6213);
nand U12079 (N_12079,N_1209,N_8796);
xor U12080 (N_12080,N_9800,N_9074);
or U12081 (N_12081,N_2836,N_1739);
or U12082 (N_12082,N_3847,N_1858);
and U12083 (N_12083,N_989,N_4559);
nor U12084 (N_12084,N_11,N_2600);
nand U12085 (N_12085,N_2026,N_5136);
and U12086 (N_12086,N_4235,N_2311);
or U12087 (N_12087,N_6552,N_873);
and U12088 (N_12088,N_6010,N_2475);
and U12089 (N_12089,N_4638,N_6532);
or U12090 (N_12090,N_9060,N_8014);
nand U12091 (N_12091,N_4269,N_9617);
and U12092 (N_12092,N_6682,N_3435);
nor U12093 (N_12093,N_2635,N_1419);
nand U12094 (N_12094,N_206,N_9624);
nand U12095 (N_12095,N_2478,N_4522);
or U12096 (N_12096,N_7346,N_5521);
and U12097 (N_12097,N_7839,N_59);
nand U12098 (N_12098,N_668,N_7189);
or U12099 (N_12099,N_7886,N_4897);
nor U12100 (N_12100,N_6575,N_2996);
nand U12101 (N_12101,N_7728,N_4968);
and U12102 (N_12102,N_6865,N_8187);
or U12103 (N_12103,N_1787,N_703);
nand U12104 (N_12104,N_7013,N_4293);
xnor U12105 (N_12105,N_416,N_8330);
nand U12106 (N_12106,N_5487,N_6234);
nor U12107 (N_12107,N_3496,N_3512);
or U12108 (N_12108,N_5493,N_1931);
nand U12109 (N_12109,N_5252,N_250);
nand U12110 (N_12110,N_6392,N_2628);
or U12111 (N_12111,N_5606,N_8232);
and U12112 (N_12112,N_7802,N_252);
or U12113 (N_12113,N_8089,N_6458);
nand U12114 (N_12114,N_3564,N_1226);
or U12115 (N_12115,N_1681,N_2778);
or U12116 (N_12116,N_7983,N_3174);
and U12117 (N_12117,N_5184,N_885);
and U12118 (N_12118,N_7758,N_2185);
nor U12119 (N_12119,N_6005,N_2560);
xor U12120 (N_12120,N_7874,N_8715);
and U12121 (N_12121,N_6199,N_7756);
and U12122 (N_12122,N_3585,N_8062);
nor U12123 (N_12123,N_7783,N_38);
nand U12124 (N_12124,N_9838,N_8951);
or U12125 (N_12125,N_5282,N_1853);
or U12126 (N_12126,N_3320,N_332);
and U12127 (N_12127,N_6413,N_3463);
nor U12128 (N_12128,N_6231,N_7885);
nand U12129 (N_12129,N_7998,N_6854);
and U12130 (N_12130,N_227,N_5155);
nor U12131 (N_12131,N_4357,N_6832);
or U12132 (N_12132,N_9974,N_2243);
and U12133 (N_12133,N_3959,N_1549);
or U12134 (N_12134,N_7679,N_2244);
nand U12135 (N_12135,N_9290,N_3252);
nand U12136 (N_12136,N_2279,N_7459);
and U12137 (N_12137,N_1804,N_344);
nor U12138 (N_12138,N_5258,N_6842);
and U12139 (N_12139,N_684,N_2098);
or U12140 (N_12140,N_2159,N_1734);
nor U12141 (N_12141,N_1806,N_7656);
and U12142 (N_12142,N_9387,N_8714);
nand U12143 (N_12143,N_2705,N_9882);
or U12144 (N_12144,N_9318,N_6988);
and U12145 (N_12145,N_7501,N_4527);
nor U12146 (N_12146,N_6789,N_2830);
and U12147 (N_12147,N_5784,N_1136);
nand U12148 (N_12148,N_322,N_8425);
and U12149 (N_12149,N_6704,N_7621);
or U12150 (N_12150,N_308,N_9439);
nor U12151 (N_12151,N_6008,N_9913);
and U12152 (N_12152,N_1169,N_2000);
and U12153 (N_12153,N_1329,N_6266);
nor U12154 (N_12154,N_7635,N_2466);
or U12155 (N_12155,N_9765,N_6260);
xnor U12156 (N_12156,N_5980,N_7228);
xnor U12157 (N_12157,N_9211,N_6365);
nor U12158 (N_12158,N_7774,N_5939);
nand U12159 (N_12159,N_3991,N_4532);
or U12160 (N_12160,N_9201,N_1634);
and U12161 (N_12161,N_2452,N_2195);
xor U12162 (N_12162,N_8823,N_4017);
or U12163 (N_12163,N_1688,N_666);
nor U12164 (N_12164,N_9664,N_7014);
nand U12165 (N_12165,N_1612,N_6647);
nor U12166 (N_12166,N_5654,N_729);
and U12167 (N_12167,N_9340,N_5369);
nand U12168 (N_12168,N_3651,N_2678);
or U12169 (N_12169,N_2765,N_1225);
nand U12170 (N_12170,N_9078,N_1532);
nor U12171 (N_12171,N_1101,N_7078);
nand U12172 (N_12172,N_5100,N_1437);
or U12173 (N_12173,N_7703,N_7335);
or U12174 (N_12174,N_6602,N_2156);
xnor U12175 (N_12175,N_7506,N_8155);
or U12176 (N_12176,N_3325,N_1668);
or U12177 (N_12177,N_8038,N_5418);
nor U12178 (N_12178,N_5685,N_4041);
nor U12179 (N_12179,N_3215,N_751);
or U12180 (N_12180,N_3412,N_7990);
or U12181 (N_12181,N_2956,N_5434);
nand U12182 (N_12182,N_8880,N_4693);
and U12183 (N_12183,N_7132,N_9793);
or U12184 (N_12184,N_5851,N_7846);
nand U12185 (N_12185,N_9476,N_3996);
and U12186 (N_12186,N_2082,N_2464);
xor U12187 (N_12187,N_3851,N_5604);
nand U12188 (N_12188,N_3549,N_75);
and U12189 (N_12189,N_430,N_5261);
nor U12190 (N_12190,N_2479,N_6962);
nand U12191 (N_12191,N_5187,N_6406);
nor U12192 (N_12192,N_8289,N_7033);
nand U12193 (N_12193,N_7402,N_4514);
or U12194 (N_12194,N_88,N_678);
xnor U12195 (N_12195,N_5002,N_9098);
nand U12196 (N_12196,N_1328,N_5115);
and U12197 (N_12197,N_8351,N_7981);
and U12198 (N_12198,N_6825,N_337);
nand U12199 (N_12199,N_7781,N_7139);
and U12200 (N_12200,N_1376,N_4268);
and U12201 (N_12201,N_7127,N_4306);
xnor U12202 (N_12202,N_9488,N_2284);
xnor U12203 (N_12203,N_5808,N_8209);
and U12204 (N_12204,N_3461,N_1333);
and U12205 (N_12205,N_5060,N_6357);
or U12206 (N_12206,N_2804,N_6920);
and U12207 (N_12207,N_1476,N_4482);
nor U12208 (N_12208,N_9918,N_4601);
nand U12209 (N_12209,N_898,N_6712);
nand U12210 (N_12210,N_9194,N_1910);
nand U12211 (N_12211,N_4813,N_9058);
or U12212 (N_12212,N_1198,N_6826);
nor U12213 (N_12213,N_6450,N_8686);
nor U12214 (N_12214,N_5897,N_8433);
xnor U12215 (N_12215,N_9552,N_8073);
nand U12216 (N_12216,N_6142,N_8109);
nand U12217 (N_12217,N_6091,N_9753);
nor U12218 (N_12218,N_1474,N_9236);
or U12219 (N_12219,N_9522,N_6415);
nand U12220 (N_12220,N_3659,N_8323);
nor U12221 (N_12221,N_1770,N_3269);
nor U12222 (N_12222,N_2610,N_8833);
nand U12223 (N_12223,N_236,N_7052);
or U12224 (N_12224,N_2664,N_6598);
and U12225 (N_12225,N_2136,N_3598);
nand U12226 (N_12226,N_7292,N_6004);
or U12227 (N_12227,N_1880,N_8327);
or U12228 (N_12228,N_7100,N_3211);
or U12229 (N_12229,N_6944,N_1754);
and U12230 (N_12230,N_1801,N_2023);
or U12231 (N_12231,N_1994,N_2324);
nor U12232 (N_12232,N_850,N_3766);
nor U12233 (N_12233,N_8643,N_3923);
nor U12234 (N_12234,N_9146,N_4158);
nand U12235 (N_12235,N_5548,N_556);
and U12236 (N_12236,N_7686,N_9);
nor U12237 (N_12237,N_6190,N_527);
and U12238 (N_12238,N_2652,N_574);
nand U12239 (N_12239,N_6782,N_8367);
and U12240 (N_12240,N_8513,N_7171);
and U12241 (N_12241,N_5992,N_3256);
xnor U12242 (N_12242,N_1807,N_1593);
nand U12243 (N_12243,N_4210,N_6061);
and U12244 (N_12244,N_8877,N_2509);
nor U12245 (N_12245,N_6654,N_1405);
xor U12246 (N_12246,N_4452,N_7446);
nor U12247 (N_12247,N_213,N_270);
or U12248 (N_12248,N_3620,N_568);
and U12249 (N_12249,N_2606,N_2977);
and U12250 (N_12250,N_7924,N_7211);
or U12251 (N_12251,N_7326,N_7611);
nor U12252 (N_12252,N_134,N_5715);
or U12253 (N_12253,N_6918,N_4428);
and U12254 (N_12254,N_7685,N_7304);
and U12255 (N_12255,N_4473,N_7089);
nor U12256 (N_12256,N_8452,N_9326);
nor U12257 (N_12257,N_5781,N_987);
nand U12258 (N_12258,N_8438,N_937);
nand U12259 (N_12259,N_483,N_5362);
nand U12260 (N_12260,N_3438,N_7453);
nor U12261 (N_12261,N_9426,N_1068);
nand U12262 (N_12262,N_1597,N_3245);
nor U12263 (N_12263,N_687,N_8628);
nor U12264 (N_12264,N_9845,N_9451);
xnor U12265 (N_12265,N_3195,N_6881);
and U12266 (N_12266,N_6655,N_3655);
or U12267 (N_12267,N_5517,N_9894);
nand U12268 (N_12268,N_3143,N_4491);
nor U12269 (N_12269,N_581,N_5575);
nor U12270 (N_12270,N_8070,N_2142);
nand U12271 (N_12271,N_6751,N_7249);
and U12272 (N_12272,N_9601,N_8604);
or U12273 (N_12273,N_839,N_8851);
and U12274 (N_12274,N_2797,N_2613);
or U12275 (N_12275,N_1707,N_4705);
or U12276 (N_12276,N_9500,N_3880);
or U12277 (N_12277,N_8303,N_3268);
or U12278 (N_12278,N_4294,N_8510);
xor U12279 (N_12279,N_2653,N_406);
or U12280 (N_12280,N_9295,N_7730);
or U12281 (N_12281,N_7217,N_6545);
nor U12282 (N_12282,N_726,N_9792);
or U12283 (N_12283,N_8374,N_7123);
or U12284 (N_12284,N_6969,N_7672);
nand U12285 (N_12285,N_7035,N_6586);
and U12286 (N_12286,N_7822,N_4936);
nor U12287 (N_12287,N_6943,N_6805);
or U12288 (N_12288,N_9676,N_5516);
or U12289 (N_12289,N_3699,N_1408);
nor U12290 (N_12290,N_8048,N_3857);
or U12291 (N_12291,N_9474,N_7745);
and U12292 (N_12292,N_9015,N_2772);
nor U12293 (N_12293,N_5984,N_4263);
nor U12294 (N_12294,N_4190,N_642);
nor U12295 (N_12295,N_458,N_677);
and U12296 (N_12296,N_173,N_2783);
and U12297 (N_12297,N_106,N_6097);
nor U12298 (N_12298,N_254,N_7565);
and U12299 (N_12299,N_3732,N_6565);
nor U12300 (N_12300,N_4867,N_3487);
nor U12301 (N_12301,N_8577,N_4483);
and U12302 (N_12302,N_9362,N_8862);
nand U12303 (N_12303,N_3849,N_3210);
or U12304 (N_12304,N_9848,N_7818);
nand U12305 (N_12305,N_2631,N_4772);
nand U12306 (N_12306,N_8503,N_5249);
and U12307 (N_12307,N_9695,N_6165);
and U12308 (N_12308,N_1548,N_4214);
and U12309 (N_12309,N_1542,N_936);
or U12310 (N_12310,N_50,N_7572);
nand U12311 (N_12311,N_2405,N_4513);
nand U12312 (N_12312,N_9777,N_3233);
nand U12313 (N_12313,N_6015,N_9502);
nor U12314 (N_12314,N_120,N_7221);
and U12315 (N_12315,N_4887,N_8724);
and U12316 (N_12316,N_1783,N_2281);
nor U12317 (N_12317,N_1671,N_9547);
and U12318 (N_12318,N_9020,N_8007);
xnor U12319 (N_12319,N_6173,N_5441);
nand U12320 (N_12320,N_7545,N_7086);
nor U12321 (N_12321,N_152,N_4710);
or U12322 (N_12322,N_4444,N_6652);
xor U12323 (N_12323,N_9394,N_3198);
and U12324 (N_12324,N_9424,N_8819);
and U12325 (N_12325,N_4861,N_9304);
and U12326 (N_12326,N_3830,N_2372);
and U12327 (N_12327,N_5161,N_843);
and U12328 (N_12328,N_4320,N_2168);
nor U12329 (N_12329,N_6356,N_6717);
or U12330 (N_12330,N_4180,N_5069);
and U12331 (N_12331,N_807,N_5271);
nor U12332 (N_12332,N_6906,N_8353);
or U12333 (N_12333,N_8630,N_1846);
and U12334 (N_12334,N_264,N_3756);
or U12335 (N_12335,N_3704,N_8740);
and U12336 (N_12336,N_4683,N_5541);
and U12337 (N_12337,N_8222,N_6482);
and U12338 (N_12338,N_2004,N_2151);
or U12339 (N_12339,N_4525,N_1128);
nor U12340 (N_12340,N_7678,N_470);
or U12341 (N_12341,N_9868,N_8332);
or U12342 (N_12342,N_7350,N_8731);
and U12343 (N_12343,N_362,N_196);
nor U12344 (N_12344,N_3173,N_4880);
and U12345 (N_12345,N_8616,N_1791);
and U12346 (N_12346,N_5937,N_1243);
or U12347 (N_12347,N_3668,N_1864);
nand U12348 (N_12348,N_5836,N_7179);
and U12349 (N_12349,N_4344,N_7702);
and U12350 (N_12350,N_7597,N_503);
nand U12351 (N_12351,N_2815,N_9851);
nor U12352 (N_12352,N_7191,N_5656);
nand U12353 (N_12353,N_5891,N_3410);
nor U12354 (N_12354,N_8065,N_2420);
and U12355 (N_12355,N_408,N_4838);
nand U12356 (N_12356,N_7436,N_5963);
nand U12357 (N_12357,N_9088,N_3292);
xnor U12358 (N_12358,N_4013,N_2641);
and U12359 (N_12359,N_5837,N_9382);
and U12360 (N_12360,N_8102,N_5750);
nand U12361 (N_12361,N_2742,N_2393);
or U12362 (N_12362,N_7890,N_3005);
and U12363 (N_12363,N_1079,N_2611);
nand U12364 (N_12364,N_9208,N_7376);
nor U12365 (N_12365,N_590,N_8783);
nor U12366 (N_12366,N_8758,N_7561);
and U12367 (N_12367,N_4011,N_4717);
xor U12368 (N_12368,N_3882,N_4261);
nand U12369 (N_12369,N_3343,N_7652);
nor U12370 (N_12370,N_8872,N_357);
and U12371 (N_12371,N_1517,N_3249);
nand U12372 (N_12372,N_8328,N_4890);
nor U12373 (N_12373,N_2411,N_312);
or U12374 (N_12374,N_8023,N_4901);
nor U12375 (N_12375,N_7253,N_2316);
xor U12376 (N_12376,N_6869,N_4007);
or U12377 (N_12377,N_8749,N_9396);
nand U12378 (N_12378,N_5139,N_9740);
nand U12379 (N_12379,N_766,N_8939);
nand U12380 (N_12380,N_9016,N_1912);
nor U12381 (N_12381,N_6787,N_5297);
nor U12382 (N_12382,N_9775,N_1427);
nor U12383 (N_12383,N_4536,N_9696);
or U12384 (N_12384,N_6485,N_4498);
or U12385 (N_12385,N_6399,N_3079);
nand U12386 (N_12386,N_5576,N_7760);
nand U12387 (N_12387,N_4411,N_8481);
nand U12388 (N_12388,N_2672,N_5655);
or U12389 (N_12389,N_225,N_4933);
nand U12390 (N_12390,N_8578,N_1468);
xor U12391 (N_12391,N_9351,N_5751);
nor U12392 (N_12392,N_3540,N_724);
xor U12393 (N_12393,N_1350,N_9506);
and U12394 (N_12394,N_5202,N_4944);
nand U12395 (N_12395,N_2829,N_7405);
nor U12396 (N_12396,N_5936,N_5311);
nor U12397 (N_12397,N_8329,N_2089);
and U12398 (N_12398,N_2057,N_6619);
and U12399 (N_12399,N_6517,N_9257);
nand U12400 (N_12400,N_3432,N_3029);
or U12401 (N_12401,N_5489,N_3043);
or U12402 (N_12402,N_8101,N_6449);
and U12403 (N_12403,N_5103,N_6237);
or U12404 (N_12404,N_3905,N_1263);
nand U12405 (N_12405,N_8270,N_3348);
xor U12406 (N_12406,N_570,N_8099);
nand U12407 (N_12407,N_6038,N_9965);
nand U12408 (N_12408,N_5061,N_9936);
nand U12409 (N_12409,N_1773,N_7892);
or U12410 (N_12410,N_8021,N_2703);
nor U12411 (N_12411,N_4961,N_282);
or U12412 (N_12412,N_7569,N_2051);
nand U12413 (N_12413,N_8576,N_1543);
or U12414 (N_12414,N_8993,N_1630);
and U12415 (N_12415,N_2681,N_2137);
nand U12416 (N_12416,N_6932,N_4069);
nor U12417 (N_12417,N_8816,N_6877);
or U12418 (N_12418,N_5349,N_5358);
and U12419 (N_12419,N_4245,N_7594);
or U12420 (N_12420,N_6146,N_67);
or U12421 (N_12421,N_8404,N_4990);
and U12422 (N_12422,N_1389,N_4031);
and U12423 (N_12423,N_4986,N_9082);
or U12424 (N_12424,N_8350,N_9985);
or U12425 (N_12425,N_4323,N_4359);
or U12426 (N_12426,N_931,N_9172);
or U12427 (N_12427,N_9515,N_4707);
and U12428 (N_12428,N_4604,N_4844);
nor U12429 (N_12429,N_8829,N_739);
and U12430 (N_12430,N_6403,N_1417);
xor U12431 (N_12431,N_9457,N_5613);
nand U12432 (N_12432,N_7291,N_4941);
and U12433 (N_12433,N_698,N_4384);
nand U12434 (N_12434,N_9345,N_5197);
nor U12435 (N_12435,N_4418,N_113);
xor U12436 (N_12436,N_3045,N_3506);
nand U12437 (N_12437,N_9152,N_4330);
nand U12438 (N_12438,N_5518,N_691);
or U12439 (N_12439,N_4849,N_5201);
and U12440 (N_12440,N_4561,N_4053);
nand U12441 (N_12441,N_4714,N_579);
nand U12442 (N_12442,N_9958,N_2596);
and U12443 (N_12443,N_1190,N_6711);
or U12444 (N_12444,N_2594,N_3862);
or U12445 (N_12445,N_478,N_1735);
xnor U12446 (N_12446,N_9039,N_2516);
xnor U12447 (N_12447,N_2273,N_1158);
nor U12448 (N_12448,N_1085,N_4467);
nor U12449 (N_12449,N_1497,N_2877);
and U12450 (N_12450,N_8834,N_1089);
nand U12451 (N_12451,N_1432,N_7358);
or U12452 (N_12452,N_2708,N_2314);
nor U12453 (N_12453,N_6253,N_7605);
nand U12454 (N_12454,N_3901,N_8719);
and U12455 (N_12455,N_7122,N_6617);
or U12456 (N_12456,N_9893,N_4552);
and U12457 (N_12457,N_7988,N_5163);
and U12458 (N_12458,N_2774,N_1227);
nor U12459 (N_12459,N_869,N_5135);
nor U12460 (N_12460,N_3229,N_1037);
and U12461 (N_12461,N_320,N_5647);
and U12462 (N_12462,N_4515,N_9239);
or U12463 (N_12463,N_6128,N_2337);
and U12464 (N_12464,N_8380,N_7875);
and U12465 (N_12465,N_8508,N_6358);
and U12466 (N_12466,N_2603,N_9048);
nand U12467 (N_12467,N_5051,N_3555);
xnor U12468 (N_12468,N_1675,N_6624);
nor U12469 (N_12469,N_8204,N_133);
or U12470 (N_12470,N_424,N_7589);
nor U12471 (N_12471,N_9320,N_8051);
xor U12472 (N_12472,N_2363,N_9925);
nand U12473 (N_12473,N_281,N_3509);
and U12474 (N_12474,N_7107,N_5649);
nor U12475 (N_12475,N_2370,N_9835);
or U12476 (N_12476,N_9795,N_609);
and U12477 (N_12477,N_7250,N_7186);
or U12478 (N_12478,N_5067,N_6241);
nand U12479 (N_12479,N_7984,N_3716);
nand U12480 (N_12480,N_3960,N_542);
xor U12481 (N_12481,N_1075,N_2049);
or U12482 (N_12482,N_4394,N_2164);
nor U12483 (N_12483,N_819,N_1003);
or U12484 (N_12484,N_9127,N_1255);
nor U12485 (N_12485,N_4971,N_4551);
and U12486 (N_12486,N_529,N_4572);
nor U12487 (N_12487,N_7856,N_1606);
and U12488 (N_12488,N_1043,N_4764);
xnor U12489 (N_12489,N_4034,N_4075);
or U12490 (N_12490,N_5637,N_1478);
or U12491 (N_12491,N_5767,N_2428);
xor U12492 (N_12492,N_498,N_617);
nor U12493 (N_12493,N_5458,N_3476);
and U12494 (N_12494,N_7183,N_7894);
or U12495 (N_12495,N_9151,N_6744);
nand U12496 (N_12496,N_8287,N_2990);
and U12497 (N_12497,N_1519,N_60);
nor U12498 (N_12498,N_8974,N_1341);
and U12499 (N_12499,N_7816,N_3919);
xnor U12500 (N_12500,N_5525,N_951);
nand U12501 (N_12501,N_7617,N_6414);
and U12502 (N_12502,N_985,N_8346);
and U12503 (N_12503,N_6200,N_3214);
and U12504 (N_12504,N_9480,N_6554);
nand U12505 (N_12505,N_3118,N_3775);
or U12506 (N_12506,N_5449,N_1595);
or U12507 (N_12507,N_437,N_1695);
nor U12508 (N_12508,N_7808,N_4331);
or U12509 (N_12509,N_7959,N_8539);
nand U12510 (N_12510,N_1976,N_7224);
nor U12511 (N_12511,N_9283,N_6052);
xor U12512 (N_12512,N_9731,N_7520);
and U12513 (N_12513,N_2246,N_4352);
nand U12514 (N_12514,N_1669,N_2075);
nand U12515 (N_12515,N_3279,N_7625);
and U12516 (N_12516,N_2065,N_7905);
nor U12517 (N_12517,N_3572,N_1873);
or U12518 (N_12518,N_7400,N_6006);
nor U12519 (N_12519,N_7277,N_1176);
or U12520 (N_12520,N_2490,N_2980);
nor U12521 (N_12521,N_1842,N_9023);
nor U12522 (N_12522,N_4299,N_7583);
and U12523 (N_12523,N_639,N_7552);
nand U12524 (N_12524,N_2123,N_9167);
xnor U12525 (N_12525,N_3914,N_7449);
or U12526 (N_12526,N_1344,N_9400);
and U12527 (N_12527,N_7018,N_3241);
nand U12528 (N_12528,N_7956,N_2083);
and U12529 (N_12529,N_3459,N_9631);
and U12530 (N_12530,N_345,N_4969);
or U12531 (N_12531,N_4674,N_5162);
or U12532 (N_12532,N_3180,N_2266);
nor U12533 (N_12533,N_1999,N_3067);
nor U12534 (N_12534,N_8169,N_6963);
nand U12535 (N_12535,N_3205,N_5003);
nand U12536 (N_12536,N_5935,N_5340);
nand U12537 (N_12537,N_5885,N_8447);
or U12538 (N_12538,N_6243,N_2112);
nor U12539 (N_12539,N_682,N_293);
nand U12540 (N_12540,N_1737,N_5088);
xnor U12541 (N_12541,N_2786,N_1454);
or U12542 (N_12542,N_9223,N_5577);
or U12543 (N_12543,N_29,N_4892);
and U12544 (N_12544,N_2538,N_6304);
or U12545 (N_12545,N_6957,N_4794);
or U12546 (N_12546,N_2304,N_5684);
and U12547 (N_12547,N_1058,N_634);
xor U12548 (N_12548,N_3875,N_9197);
nor U12549 (N_12549,N_7535,N_2629);
nor U12550 (N_12550,N_1360,N_7038);
and U12551 (N_12551,N_8428,N_1879);
nand U12552 (N_12552,N_1238,N_2962);
nand U12553 (N_12553,N_6124,N_6681);
and U12554 (N_12554,N_4335,N_1295);
and U12555 (N_12555,N_2873,N_6998);
nand U12556 (N_12556,N_2699,N_9267);
or U12557 (N_12557,N_9493,N_782);
nor U12558 (N_12558,N_6028,N_5210);
and U12559 (N_12559,N_8466,N_1699);
and U12560 (N_12560,N_7489,N_2947);
nor U12561 (N_12561,N_2617,N_2121);
xnor U12562 (N_12562,N_732,N_3865);
and U12563 (N_12563,N_5932,N_7867);
or U12564 (N_12564,N_2750,N_8881);
nand U12565 (N_12565,N_434,N_4750);
and U12566 (N_12566,N_3868,N_147);
and U12567 (N_12567,N_487,N_2251);
nand U12568 (N_12568,N_4002,N_4287);
and U12569 (N_12569,N_5251,N_6768);
or U12570 (N_12570,N_9643,N_3334);
or U12571 (N_12571,N_8134,N_4488);
or U12572 (N_12572,N_6157,N_8146);
nand U12573 (N_12573,N_1477,N_8191);
nand U12574 (N_12574,N_364,N_2032);
or U12575 (N_12575,N_952,N_3964);
nand U12576 (N_12576,N_9461,N_4804);
or U12577 (N_12577,N_6611,N_5583);
nor U12578 (N_12578,N_7494,N_8774);
nand U12579 (N_12579,N_2856,N_7134);
or U12580 (N_12580,N_7549,N_9747);
and U12581 (N_12581,N_5598,N_2441);
nor U12582 (N_12582,N_8638,N_1062);
nor U12583 (N_12583,N_7750,N_1391);
and U12584 (N_12584,N_3437,N_9749);
nor U12585 (N_12585,N_5841,N_3222);
or U12586 (N_12586,N_7390,N_5617);
and U12587 (N_12587,N_9221,N_6034);
or U12588 (N_12588,N_2461,N_4050);
nor U12589 (N_12589,N_8159,N_7146);
or U12590 (N_12590,N_7965,N_6140);
or U12591 (N_12591,N_3251,N_8022);
nand U12592 (N_12592,N_6184,N_7444);
nor U12593 (N_12593,N_628,N_4453);
or U12594 (N_12594,N_8685,N_1701);
and U12595 (N_12595,N_1538,N_8085);
nor U12596 (N_12596,N_7946,N_4781);
nand U12597 (N_12597,N_5440,N_6857);
or U12598 (N_12598,N_1482,N_6447);
nand U12599 (N_12599,N_9245,N_5182);
and U12600 (N_12600,N_8419,N_2206);
nor U12601 (N_12601,N_941,N_4605);
and U12602 (N_12602,N_2497,N_983);
and U12603 (N_12603,N_3324,N_5058);
or U12604 (N_12604,N_3287,N_4157);
or U12605 (N_12605,N_9581,N_5658);
and U12606 (N_12606,N_754,N_2647);
nor U12607 (N_12607,N_1428,N_7272);
and U12608 (N_12608,N_2384,N_3803);
or U12609 (N_12609,N_5933,N_9156);
nand U12610 (N_12610,N_9256,N_2812);
nand U12611 (N_12611,N_2659,N_9665);
and U12612 (N_12612,N_5375,N_2067);
nand U12613 (N_12613,N_1763,N_1838);
nor U12614 (N_12614,N_7296,N_8480);
nand U12615 (N_12615,N_9130,N_8769);
and U12616 (N_12616,N_7973,N_7897);
xor U12617 (N_12617,N_3672,N_7699);
or U12618 (N_12618,N_9527,N_7744);
nor U12619 (N_12619,N_9139,N_464);
or U12620 (N_12620,N_4062,N_8547);
or U12621 (N_12621,N_1168,N_5144);
and U12622 (N_12622,N_2227,N_4111);
nand U12623 (N_12623,N_3750,N_3073);
nor U12624 (N_12624,N_7090,N_1602);
or U12625 (N_12625,N_3734,N_4028);
nand U12626 (N_12626,N_6423,N_3072);
nor U12627 (N_12627,N_4351,N_1271);
and U12628 (N_12628,N_8116,N_8650);
nor U12629 (N_12629,N_6111,N_2469);
and U12630 (N_12630,N_7495,N_1444);
or U12631 (N_12631,N_8229,N_4247);
nor U12632 (N_12632,N_8563,N_187);
nor U12633 (N_12633,N_1684,N_103);
and U12634 (N_12634,N_6913,N_9306);
nand U12635 (N_12635,N_1167,N_6915);
or U12636 (N_12636,N_6453,N_3712);
and U12637 (N_12637,N_6465,N_3770);
or U12638 (N_12638,N_3731,N_2638);
nand U12639 (N_12639,N_1882,N_5303);
and U12640 (N_12640,N_283,N_9608);
nand U12641 (N_12641,N_4464,N_3381);
nor U12642 (N_12642,N_653,N_8147);
nand U12643 (N_12643,N_5675,N_4850);
nand U12644 (N_12644,N_7794,N_8213);
xnor U12645 (N_12645,N_4182,N_3076);
xor U12646 (N_12646,N_5827,N_3147);
and U12647 (N_12647,N_3483,N_7932);
or U12648 (N_12648,N_1467,N_2711);
and U12649 (N_12649,N_2453,N_8375);
xor U12650 (N_12650,N_4932,N_9814);
and U12651 (N_12651,N_916,N_6757);
and U12652 (N_12652,N_3983,N_7274);
nor U12653 (N_12653,N_6593,N_2805);
nor U12654 (N_12654,N_4573,N_8550);
or U12655 (N_12655,N_2094,N_279);
nand U12656 (N_12656,N_2183,N_7972);
nand U12657 (N_12657,N_5660,N_4016);
nor U12658 (N_12658,N_6959,N_3817);
nand U12659 (N_12659,N_6400,N_3120);
nand U12660 (N_12660,N_1254,N_730);
or U12661 (N_12661,N_2585,N_3299);
nand U12662 (N_12662,N_699,N_2022);
nand U12663 (N_12663,N_8457,N_4098);
or U12664 (N_12664,N_9509,N_4419);
and U12665 (N_12665,N_9390,N_8571);
nor U12666 (N_12666,N_1781,N_2790);
xnor U12667 (N_12667,N_1347,N_5535);
and U12668 (N_12668,N_4752,N_9878);
xnor U12669 (N_12669,N_4722,N_4000);
and U12670 (N_12670,N_2860,N_2277);
or U12671 (N_12671,N_6195,N_658);
or U12672 (N_12672,N_6212,N_8324);
nand U12673 (N_12673,N_3264,N_280);
and U12674 (N_12674,N_1885,N_1774);
nand U12675 (N_12675,N_8243,N_37);
nand U12676 (N_12676,N_9807,N_551);
nor U12677 (N_12677,N_7913,N_4035);
or U12678 (N_12678,N_8398,N_959);
or U12679 (N_12679,N_5690,N_2110);
nand U12680 (N_12680,N_559,N_5903);
nand U12681 (N_12681,N_7452,N_6023);
nor U12682 (N_12682,N_8347,N_6723);
nand U12683 (N_12683,N_9842,N_9331);
nor U12684 (N_12684,N_2456,N_2722);
and U12685 (N_12685,N_7289,N_9922);
nand U12686 (N_12686,N_5747,N_6596);
and U12687 (N_12687,N_7736,N_1658);
nand U12688 (N_12688,N_7418,N_8162);
nand U12689 (N_12689,N_3336,N_3956);
nand U12690 (N_12690,N_1362,N_5563);
and U12691 (N_12691,N_9363,N_9701);
nand U12692 (N_12692,N_2416,N_5991);
nor U12693 (N_12693,N_5895,N_6360);
or U12694 (N_12694,N_7300,N_5823);
nor U12695 (N_12695,N_6186,N_9962);
xnor U12696 (N_12696,N_7374,N_3069);
or U12697 (N_12697,N_8339,N_185);
and U12698 (N_12698,N_4395,N_6416);
nor U12699 (N_12699,N_7099,N_2853);
nor U12700 (N_12700,N_217,N_4403);
nor U12701 (N_12701,N_9052,N_1268);
nand U12702 (N_12702,N_243,N_5057);
nand U12703 (N_12703,N_2908,N_7188);
nor U12704 (N_12704,N_4709,N_2764);
nor U12705 (N_12705,N_719,N_5361);
nor U12706 (N_12706,N_6564,N_727);
and U12707 (N_12707,N_2887,N_9647);
and U12708 (N_12708,N_8335,N_2892);
nor U12709 (N_12709,N_2297,N_2485);
xor U12710 (N_12710,N_7780,N_8985);
nor U12711 (N_12711,N_9278,N_1834);
or U12712 (N_12712,N_7525,N_4475);
or U12713 (N_12713,N_2105,N_8581);
nand U12714 (N_12714,N_7055,N_8505);
and U12715 (N_12715,N_4537,N_7200);
nor U12716 (N_12716,N_3701,N_9524);
or U12717 (N_12717,N_8950,N_1629);
nor U12718 (N_12718,N_8716,N_4132);
or U12719 (N_12719,N_3883,N_1027);
or U12720 (N_12720,N_4417,N_736);
nand U12721 (N_12721,N_6017,N_9449);
and U12722 (N_12722,N_5944,N_5308);
or U12723 (N_12723,N_3311,N_6752);
and U12724 (N_12724,N_9649,N_1461);
or U12725 (N_12725,N_3099,N_2928);
nor U12726 (N_12726,N_6875,N_5678);
and U12727 (N_12727,N_7281,N_2535);
xor U12728 (N_12728,N_1020,N_7483);
or U12729 (N_12729,N_3454,N_2992);
and U12730 (N_12730,N_2608,N_36);
nand U12731 (N_12731,N_6967,N_5723);
nand U12732 (N_12732,N_356,N_5398);
and U12733 (N_12733,N_9443,N_1399);
nand U12734 (N_12734,N_9495,N_5291);
or U12735 (N_12735,N_5972,N_3835);
xor U12736 (N_12736,N_6176,N_4820);
nor U12737 (N_12737,N_4865,N_4842);
nor U12738 (N_12738,N_2690,N_6727);
nand U12739 (N_12739,N_9768,N_3132);
nand U12740 (N_12740,N_3346,N_1345);
and U12741 (N_12741,N_9442,N_5744);
nor U12742 (N_12742,N_4087,N_637);
or U12743 (N_12743,N_6922,N_4173);
or U12744 (N_12744,N_2489,N_1554);
xor U12745 (N_12745,N_7562,N_599);
nand U12746 (N_12746,N_9992,N_4903);
or U12747 (N_12747,N_6132,N_7926);
or U12748 (N_12748,N_5085,N_2404);
or U12749 (N_12749,N_4122,N_6651);
nand U12750 (N_12750,N_4613,N_9626);
nor U12751 (N_12751,N_1063,N_2125);
xor U12752 (N_12752,N_6439,N_4093);
xnor U12753 (N_12753,N_343,N_7138);
nand U12754 (N_12754,N_872,N_4374);
nand U12755 (N_12755,N_8233,N_9055);
and U12756 (N_12756,N_212,N_7871);
xor U12757 (N_12757,N_2350,N_8557);
nand U12758 (N_12758,N_5731,N_7036);
nor U12759 (N_12759,N_7185,N_1382);
nor U12760 (N_12760,N_1992,N_3726);
or U12761 (N_12761,N_2924,N_7634);
nor U12762 (N_12762,N_7210,N_3378);
xor U12763 (N_12763,N_5468,N_3027);
nand U12764 (N_12764,N_9693,N_8771);
and U12765 (N_12765,N_5195,N_5198);
nand U12766 (N_12766,N_8599,N_3417);
or U12767 (N_12767,N_9132,N_2918);
nor U12768 (N_12768,N_4952,N_386);
and U12769 (N_12769,N_7641,N_1457);
and U12770 (N_12770,N_7810,N_9168);
and U12771 (N_12771,N_5215,N_5682);
and U12772 (N_12772,N_7497,N_8949);
or U12773 (N_12773,N_6996,N_6236);
or U12774 (N_12774,N_1336,N_5062);
nor U12775 (N_12775,N_3309,N_922);
nand U12776 (N_12776,N_8371,N_4355);
and U12777 (N_12777,N_1273,N_5546);
nand U12778 (N_12778,N_3588,N_4116);
nor U12779 (N_12779,N_3146,N_2794);
nor U12780 (N_12780,N_2612,N_8012);
nand U12781 (N_12781,N_563,N_5363);
and U12782 (N_12782,N_511,N_2735);
or U12783 (N_12783,N_5800,N_7908);
nand U12784 (N_12784,N_1884,N_3837);
nand U12785 (N_12785,N_2616,N_9917);
or U12786 (N_12786,N_1265,N_9177);
nand U12787 (N_12787,N_8893,N_6563);
and U12788 (N_12788,N_4879,N_6876);
and U12789 (N_12789,N_9979,N_888);
and U12790 (N_12790,N_7590,N_834);
and U12791 (N_12791,N_4213,N_7660);
nor U12792 (N_12792,N_6535,N_9684);
and U12793 (N_12793,N_3690,N_4237);
nor U12794 (N_12794,N_7628,N_6628);
or U12795 (N_12795,N_4569,N_3274);
nand U12796 (N_12796,N_7515,N_135);
or U12797 (N_12797,N_7283,N_7725);
nor U12798 (N_12798,N_2414,N_7467);
and U12799 (N_12799,N_2645,N_9106);
and U12800 (N_12800,N_4791,N_646);
or U12801 (N_12801,N_8727,N_7568);
xor U12802 (N_12802,N_7716,N_3643);
nand U12803 (N_12803,N_5928,N_7476);
xnor U12804 (N_12804,N_5832,N_2189);
and U12805 (N_12805,N_2845,N_9657);
nor U12806 (N_12806,N_8556,N_1434);
nor U12807 (N_12807,N_5086,N_7462);
nor U12808 (N_12808,N_7944,N_9620);
or U12809 (N_12809,N_3052,N_3247);
or U12810 (N_12810,N_7643,N_2865);
xnor U12811 (N_12811,N_9788,N_8364);
nand U12812 (N_12812,N_4125,N_2929);
nand U12813 (N_12813,N_1076,N_8871);
and U12814 (N_12814,N_7653,N_3689);
nor U12815 (N_12815,N_9299,N_4307);
nand U12816 (N_12816,N_375,N_3507);
and U12817 (N_12817,N_9553,N_1908);
or U12818 (N_12818,N_8124,N_2499);
nand U12819 (N_12819,N_7331,N_7587);
nand U12820 (N_12820,N_7910,N_3727);
nand U12821 (N_12821,N_3209,N_1545);
nor U12822 (N_12822,N_9393,N_7355);
nor U12823 (N_12823,N_4106,N_5752);
or U12824 (N_12824,N_6809,N_4401);
and U12825 (N_12825,N_1278,N_160);
and U12826 (N_12826,N_7954,N_2739);
nand U12827 (N_12827,N_8632,N_5828);
nand U12828 (N_12828,N_2017,N_960);
nand U12829 (N_12829,N_1896,N_6445);
nor U12830 (N_12830,N_2580,N_9425);
or U12831 (N_12831,N_9053,N_4806);
nor U12832 (N_12832,N_9323,N_1486);
or U12833 (N_12833,N_2909,N_8761);
and U12834 (N_12834,N_4665,N_891);
nand U12835 (N_12835,N_1904,N_7806);
nor U12836 (N_12836,N_9178,N_1450);
xnor U12837 (N_12837,N_2734,N_7301);
and U12838 (N_12838,N_2129,N_291);
and U12839 (N_12839,N_8565,N_5121);
or U12840 (N_12840,N_7831,N_1655);
and U12841 (N_12841,N_6039,N_409);
or U12842 (N_12842,N_6817,N_7442);
nor U12843 (N_12843,N_5106,N_8660);
or U12844 (N_12844,N_8931,N_4244);
or U12845 (N_12845,N_5696,N_9399);
or U12846 (N_12846,N_4947,N_6779);
or U12847 (N_12847,N_9550,N_4170);
nand U12848 (N_12848,N_3017,N_6083);
nor U12849 (N_12849,N_8977,N_9181);
or U12850 (N_12850,N_8246,N_1718);
nor U12851 (N_12851,N_9762,N_220);
or U12852 (N_12852,N_6572,N_3172);
or U12853 (N_12853,N_1817,N_6529);
nor U12854 (N_12854,N_7069,N_1642);
or U12855 (N_12855,N_6601,N_4092);
and U12856 (N_12856,N_6210,N_2673);
nand U12857 (N_12857,N_3608,N_9312);
nand U12858 (N_12858,N_2044,N_4631);
or U12859 (N_12859,N_3286,N_2785);
xor U12860 (N_12860,N_4145,N_1766);
nand U12861 (N_12861,N_2248,N_9244);
or U12862 (N_12862,N_945,N_1504);
nor U12863 (N_12863,N_9430,N_8249);
nor U12864 (N_12864,N_7755,N_9373);
xnor U12865 (N_12865,N_2496,N_6063);
and U12866 (N_12866,N_98,N_4440);
nand U12867 (N_12867,N_6770,N_9889);
or U12868 (N_12868,N_4200,N_8432);
and U12869 (N_12869,N_5804,N_4342);
nor U12870 (N_12870,N_7996,N_19);
nor U12871 (N_12871,N_4378,N_9153);
nor U12872 (N_12872,N_9333,N_7027);
nand U12873 (N_12873,N_9272,N_5666);
or U12874 (N_12874,N_8139,N_397);
and U12875 (N_12875,N_490,N_6064);
nand U12876 (N_12876,N_1825,N_2521);
nand U12877 (N_12877,N_1641,N_5853);
nand U12878 (N_12878,N_2272,N_6911);
nand U12879 (N_12879,N_8189,N_8059);
nand U12880 (N_12880,N_8549,N_1490);
xnor U12881 (N_12881,N_588,N_623);
nor U12882 (N_12882,N_7473,N_1985);
or U12883 (N_12883,N_7263,N_2864);
or U12884 (N_12884,N_3815,N_7417);
nand U12885 (N_12885,N_603,N_8580);
nand U12886 (N_12886,N_5882,N_5738);
xnor U12887 (N_12887,N_1861,N_2152);
and U12888 (N_12888,N_1370,N_3114);
nand U12889 (N_12889,N_231,N_3930);
or U12890 (N_12890,N_6215,N_3202);
nand U12891 (N_12891,N_3484,N_9730);
and U12892 (N_12892,N_5118,N_8071);
nor U12893 (N_12893,N_2235,N_5020);
or U12894 (N_12894,N_4143,N_8476);
or U12895 (N_12895,N_7365,N_4183);
or U12896 (N_12896,N_3782,N_6902);
nand U12897 (N_12897,N_9388,N_361);
xor U12898 (N_12898,N_5973,N_4624);
xor U12899 (N_12899,N_859,N_55);
or U12900 (N_12900,N_867,N_9116);
nor U12901 (N_12901,N_8217,N_8441);
xnor U12902 (N_12902,N_219,N_8728);
nand U12903 (N_12903,N_5307,N_2362);
xnor U12904 (N_12904,N_4318,N_3891);
nand U12905 (N_12905,N_8773,N_3001);
or U12906 (N_12906,N_9533,N_1847);
nor U12907 (N_12907,N_9516,N_848);
and U12908 (N_12908,N_3077,N_4463);
nor U12909 (N_12909,N_2373,N_7798);
nor U12910 (N_12910,N_2715,N_1644);
nor U12911 (N_12911,N_1332,N_2267);
or U12912 (N_12912,N_5754,N_8646);
and U12913 (N_12913,N_7978,N_3984);
or U12914 (N_12914,N_3612,N_3898);
nand U12915 (N_12915,N_6462,N_3019);
or U12916 (N_12916,N_3702,N_8381);
or U12917 (N_12917,N_6797,N_3899);
nor U12918 (N_12918,N_4396,N_8265);
nand U12919 (N_12919,N_6281,N_8524);
and U12920 (N_12920,N_4388,N_7943);
and U12921 (N_12921,N_149,N_8343);
nor U12922 (N_12922,N_8000,N_9855);
xnor U12923 (N_12923,N_909,N_9771);
nor U12924 (N_12924,N_371,N_6548);
xnor U12925 (N_12925,N_5216,N_7571);
and U12926 (N_12926,N_5178,N_4846);
or U12927 (N_12927,N_9841,N_5809);
nor U12928 (N_12928,N_1508,N_2789);
xnor U12929 (N_12929,N_4334,N_99);
or U12930 (N_12930,N_1436,N_5017);
or U12931 (N_12931,N_2256,N_5323);
xnor U12932 (N_12932,N_3199,N_5920);
nand U12933 (N_12933,N_7962,N_7948);
nor U12934 (N_12934,N_6493,N_2685);
nor U12935 (N_12935,N_2537,N_4149);
nand U12936 (N_12936,N_8465,N_3349);
or U12937 (N_12937,N_7425,N_5564);
xor U12938 (N_12938,N_4391,N_830);
and U12939 (N_12939,N_1888,N_933);
or U12940 (N_12940,N_2595,N_7023);
nand U12941 (N_12941,N_9790,N_146);
or U12942 (N_12942,N_4208,N_9189);
nor U12943 (N_12943,N_7666,N_5629);
xnor U12944 (N_12944,N_2578,N_9431);
and U12945 (N_12945,N_9344,N_9035);
nand U12946 (N_12946,N_8558,N_5140);
or U12947 (N_12947,N_4385,N_3105);
nor U12948 (N_12948,N_5506,N_7267);
nor U12949 (N_12949,N_6224,N_8300);
or U12950 (N_12950,N_7053,N_4441);
and U12951 (N_12951,N_7397,N_681);
nand U12952 (N_12952,N_7540,N_8238);
nor U12953 (N_12953,N_5240,N_8905);
and U12954 (N_12954,N_2197,N_818);
or U12955 (N_12955,N_2238,N_5620);
xnor U12956 (N_12956,N_4333,N_6684);
nor U12957 (N_12957,N_2177,N_4863);
and U12958 (N_12958,N_8462,N_6765);
xor U12959 (N_12959,N_2901,N_7243);
nor U12960 (N_12960,N_341,N_4738);
and U12961 (N_12961,N_1851,N_7194);
nor U12962 (N_12962,N_7815,N_4959);
and U12963 (N_12963,N_7059,N_1588);
xor U12964 (N_12964,N_3376,N_2730);
and U12965 (N_12965,N_472,N_2202);
nand U12966 (N_12966,N_4264,N_2709);
nor U12967 (N_12967,N_7830,N_6311);
xor U12968 (N_12968,N_9846,N_4128);
or U12969 (N_12969,N_5332,N_5863);
or U12970 (N_12970,N_897,N_9951);
and U12971 (N_12971,N_972,N_360);
nor U12972 (N_12972,N_3589,N_7485);
nand U12973 (N_12973,N_2986,N_7529);
or U12974 (N_12974,N_1250,N_5295);
or U12975 (N_12975,N_8542,N_8133);
and U12976 (N_12976,N_6726,N_3780);
nand U12977 (N_12977,N_1997,N_3760);
nand U12978 (N_12978,N_7543,N_1967);
nor U12979 (N_12979,N_8582,N_7092);
nor U12980 (N_12980,N_2477,N_6518);
nand U12981 (N_12981,N_5479,N_4284);
and U12982 (N_12982,N_8642,N_8671);
nor U12983 (N_12983,N_8225,N_5913);
nand U12984 (N_12984,N_4821,N_7409);
nand U12985 (N_12985,N_8322,N_5092);
nand U12986 (N_12986,N_9095,N_4599);
nor U12987 (N_12987,N_894,N_9935);
and U12988 (N_12988,N_2029,N_1649);
nand U12989 (N_12989,N_4652,N_3757);
nor U12990 (N_12990,N_4929,N_72);
and U12991 (N_12991,N_6472,N_3516);
nor U12992 (N_12992,N_7314,N_3141);
nor U12993 (N_12993,N_6924,N_4054);
and U12994 (N_12994,N_5451,N_5407);
or U12995 (N_12995,N_3175,N_3872);
xnor U12996 (N_12996,N_289,N_5083);
nor U12997 (N_12997,N_5093,N_4271);
nand U12998 (N_12998,N_42,N_4934);
nor U12999 (N_12999,N_9243,N_4606);
or U13000 (N_13000,N_9820,N_1581);
or U13001 (N_13001,N_3411,N_7901);
nor U13002 (N_13002,N_5736,N_5894);
nor U13003 (N_13003,N_2174,N_4840);
or U13004 (N_13004,N_9503,N_4257);
or U13005 (N_13005,N_4078,N_6833);
or U13006 (N_13006,N_2109,N_6899);
and U13007 (N_13007,N_8348,N_6710);
and U13008 (N_13008,N_8631,N_4671);
or U13009 (N_13009,N_9853,N_8723);
and U13010 (N_13010,N_3345,N_4614);
xnor U13011 (N_13011,N_4080,N_8765);
nand U13012 (N_13012,N_6823,N_6570);
xnor U13013 (N_13013,N_2491,N_1845);
and U13014 (N_13014,N_8736,N_7009);
or U13015 (N_13015,N_4225,N_831);
nor U13016 (N_13016,N_9827,N_1945);
and U13017 (N_13017,N_4596,N_8153);
and U13018 (N_13018,N_9757,N_9571);
or U13019 (N_13019,N_5260,N_6284);
or U13020 (N_13020,N_9046,N_627);
nand U13021 (N_13021,N_1530,N_9964);
nor U13022 (N_13022,N_5405,N_1325);
or U13023 (N_13023,N_593,N_2096);
nor U13024 (N_13024,N_1289,N_5743);
nand U13025 (N_13025,N_4048,N_8579);
and U13026 (N_13026,N_6455,N_435);
nand U13027 (N_13027,N_310,N_3258);
or U13028 (N_13028,N_9575,N_3522);
or U13029 (N_13029,N_1625,N_4086);
nand U13030 (N_13030,N_5539,N_5388);
nand U13031 (N_13031,N_2905,N_7793);
nand U13032 (N_13032,N_3015,N_6968);
nand U13033 (N_13033,N_7153,N_6808);
nor U13034 (N_13034,N_2134,N_6523);
nor U13035 (N_13035,N_7043,N_7664);
and U13036 (N_13036,N_6521,N_3003);
nor U13037 (N_13037,N_649,N_1159);
nor U13038 (N_13038,N_1502,N_9174);
nor U13039 (N_13039,N_9064,N_8574);
nor U13040 (N_13040,N_3248,N_7704);
and U13041 (N_13041,N_6951,N_1112);
nand U13042 (N_13042,N_4490,N_3372);
nand U13043 (N_13043,N_1090,N_5515);
nand U13044 (N_13044,N_5024,N_4292);
nand U13045 (N_13045,N_899,N_3430);
or U13046 (N_13046,N_214,N_9678);
nor U13047 (N_13047,N_2245,N_9733);
and U13048 (N_13048,N_2295,N_576);
nand U13049 (N_13049,N_7352,N_4774);
xnor U13050 (N_13050,N_318,N_2045);
xnor U13051 (N_13051,N_5179,N_2257);
or U13052 (N_13052,N_631,N_5683);
nand U13053 (N_13053,N_9779,N_382);
nand U13054 (N_13054,N_4649,N_7424);
and U13055 (N_13055,N_8965,N_7914);
nor U13056 (N_13056,N_1447,N_4019);
nand U13057 (N_13057,N_3152,N_9444);
nand U13058 (N_13058,N_1758,N_1544);
xor U13059 (N_13059,N_403,N_9641);
nor U13060 (N_13060,N_4607,N_2849);
and U13061 (N_13061,N_7161,N_249);
or U13062 (N_13062,N_875,N_9505);
nand U13063 (N_13063,N_8536,N_9491);
nand U13064 (N_13064,N_566,N_9742);
and U13065 (N_13065,N_4967,N_4627);
and U13066 (N_13066,N_1521,N_5640);
or U13067 (N_13067,N_662,N_1286);
and U13068 (N_13068,N_783,N_7238);
nor U13069 (N_13069,N_8114,N_8208);
nand U13070 (N_13070,N_4663,N_1820);
nor U13071 (N_13071,N_7843,N_829);
nor U13072 (N_13072,N_2757,N_6158);
and U13073 (N_13073,N_4387,N_2658);
and U13074 (N_13074,N_3545,N_9291);
nor U13075 (N_13075,N_4656,N_5401);
and U13076 (N_13076,N_871,N_1380);
nand U13077 (N_13077,N_8477,N_8408);
and U13078 (N_13078,N_248,N_208);
nand U13079 (N_13079,N_3812,N_6427);
or U13080 (N_13080,N_5538,N_750);
nor U13081 (N_13081,N_2446,N_9087);
and U13082 (N_13082,N_7407,N_6267);
nand U13083 (N_13083,N_5267,N_5831);
nor U13084 (N_13084,N_3628,N_5618);
nor U13085 (N_13085,N_3161,N_2548);
or U13086 (N_13086,N_2667,N_2816);
nor U13087 (N_13087,N_5622,N_8341);
and U13088 (N_13088,N_753,N_7202);
xnor U13089 (N_13089,N_2867,N_6945);
and U13090 (N_13090,N_8451,N_8553);
nor U13091 (N_13091,N_3524,N_1107);
xnor U13092 (N_13092,N_8215,N_4695);
nor U13093 (N_13093,N_3262,N_8113);
and U13094 (N_13094,N_9337,N_6994);
and U13095 (N_13095,N_6088,N_6562);
nand U13096 (N_13096,N_2084,N_3805);
nand U13097 (N_13097,N_5702,N_6550);
nand U13098 (N_13098,N_4608,N_6322);
and U13099 (N_13099,N_9209,N_6699);
and U13100 (N_13100,N_3275,N_9100);
nand U13101 (N_13101,N_6621,N_9996);
nor U13102 (N_13102,N_9136,N_2684);
or U13103 (N_13103,N_1723,N_5018);
nor U13104 (N_13104,N_9107,N_3802);
nand U13105 (N_13105,N_6469,N_4130);
or U13106 (N_13106,N_3948,N_4853);
nand U13107 (N_13107,N_2061,N_9836);
xor U13108 (N_13108,N_2192,N_8997);
and U13109 (N_13109,N_1284,N_1878);
or U13110 (N_13110,N_2747,N_8751);
or U13111 (N_13111,N_5437,N_2012);
nand U13112 (N_13112,N_878,N_7423);
nor U13113 (N_13113,N_4084,N_2348);
and U13114 (N_13114,N_5040,N_1473);
nor U13115 (N_13115,N_828,N_9040);
or U13116 (N_13116,N_7693,N_5318);
or U13117 (N_13117,N_5481,N_7644);
and U13118 (N_13118,N_8214,N_3866);
and U13119 (N_13119,N_1722,N_2321);
nor U13120 (N_13120,N_880,N_6166);
or U13121 (N_13121,N_1651,N_1028);
xor U13122 (N_13122,N_9813,N_2486);
or U13123 (N_13123,N_3083,N_8824);
nand U13124 (N_13124,N_6653,N_3511);
xnor U13125 (N_13125,N_601,N_5125);
and U13126 (N_13126,N_3840,N_1496);
or U13127 (N_13127,N_8698,N_5065);
and U13128 (N_13128,N_39,N_8373);
or U13129 (N_13129,N_8027,N_7399);
or U13130 (N_13130,N_3244,N_8046);
or U13131 (N_13131,N_7770,N_2657);
xnor U13132 (N_13132,N_9386,N_6705);
nor U13133 (N_13133,N_1493,N_2533);
xor U13134 (N_13134,N_7600,N_877);
nor U13135 (N_13135,N_806,N_1386);
nand U13136 (N_13136,N_7955,N_9485);
or U13137 (N_13137,N_9158,N_2775);
xor U13138 (N_13138,N_949,N_6417);
xnor U13139 (N_13139,N_1025,N_7175);
nand U13140 (N_13140,N_1893,N_2264);
or U13141 (N_13141,N_1140,N_358);
nand U13142 (N_13142,N_6766,N_621);
nand U13143 (N_13143,N_2936,N_1585);
nor U13144 (N_13144,N_2983,N_5146);
nand U13145 (N_13145,N_3528,N_2495);
nor U13146 (N_13146,N_8575,N_6081);
and U13147 (N_13147,N_8519,N_5983);
nand U13148 (N_13148,N_5689,N_9822);
nor U13149 (N_13149,N_1384,N_8403);
and U13150 (N_13150,N_5923,N_1899);
nand U13151 (N_13151,N_1897,N_2935);
nand U13152 (N_13152,N_8981,N_2858);
nor U13153 (N_13153,N_2431,N_5871);
or U13154 (N_13154,N_5858,N_4230);
and U13155 (N_13155,N_8005,N_5124);
and U13156 (N_13156,N_2527,N_2663);
nor U13157 (N_13157,N_9401,N_5423);
or U13158 (N_13158,N_9225,N_1375);
nor U13159 (N_13159,N_2906,N_3833);
nor U13160 (N_13160,N_9735,N_5050);
or U13161 (N_13161,N_6251,N_6930);
xor U13162 (N_13162,N_8808,N_6177);
xor U13163 (N_13163,N_6030,N_5815);
nand U13164 (N_13164,N_9671,N_93);
or U13165 (N_13165,N_2181,N_8940);
or U13166 (N_13166,N_8762,N_7474);
or U13167 (N_13167,N_5044,N_1547);
nand U13168 (N_13168,N_5305,N_3316);
and U13169 (N_13169,N_8717,N_8148);
nor U13170 (N_13170,N_8986,N_2041);
or U13171 (N_13171,N_2505,N_669);
and U13172 (N_13172,N_3821,N_3318);
nor U13173 (N_13173,N_1977,N_910);
and U13174 (N_13174,N_3611,N_6670);
nand U13175 (N_13175,N_652,N_2583);
nor U13176 (N_13176,N_4121,N_3683);
nor U13177 (N_13177,N_9090,N_9588);
nand U13178 (N_13178,N_7773,N_8733);
and U13179 (N_13179,N_5014,N_9634);
and U13180 (N_13180,N_7945,N_5704);
or U13181 (N_13181,N_5394,N_56);
xor U13182 (N_13182,N_493,N_2118);
and U13183 (N_13183,N_9068,N_4278);
or U13184 (N_13184,N_812,N_2093);
and U13185 (N_13185,N_2385,N_6997);
xor U13186 (N_13186,N_6232,N_6143);
nand U13187 (N_13187,N_3565,N_8538);
nor U13188 (N_13188,N_2781,N_6871);
and U13189 (N_13189,N_6520,N_7223);
or U13190 (N_13190,N_1485,N_9364);
or U13191 (N_13191,N_3495,N_1049);
and U13192 (N_13192,N_10,N_817);
nor U13193 (N_13193,N_6043,N_6217);
nor U13194 (N_13194,N_4135,N_608);
xnor U13195 (N_13195,N_3530,N_7316);
and U13196 (N_13196,N_9440,N_8913);
nor U13197 (N_13197,N_6758,N_7226);
nand U13198 (N_13198,N_8164,N_2171);
nand U13199 (N_13199,N_7366,N_779);
and U13200 (N_13200,N_8006,N_8789);
and U13201 (N_13201,N_7322,N_8559);
nand U13202 (N_13202,N_5628,N_8092);
nor U13203 (N_13203,N_3747,N_2520);
nor U13204 (N_13204,N_6695,N_9637);
and U13205 (N_13205,N_3474,N_9454);
and U13206 (N_13206,N_2944,N_6353);
xor U13207 (N_13207,N_4686,N_117);
or U13208 (N_13208,N_674,N_958);
xor U13209 (N_13209,N_1156,N_6285);
and U13210 (N_13210,N_7463,N_8180);
nor U13211 (N_13211,N_6086,N_9286);
or U13212 (N_13212,N_6437,N_7713);
and U13213 (N_13213,N_8019,N_2793);
nor U13214 (N_13214,N_1264,N_5578);
nand U13215 (N_13215,N_4006,N_8828);
or U13216 (N_13216,N_8039,N_8696);
and U13217 (N_13217,N_8648,N_3086);
xnor U13218 (N_13218,N_6995,N_471);
xor U13219 (N_13219,N_2236,N_8149);
or U13220 (N_13220,N_9802,N_6519);
and U13221 (N_13221,N_2661,N_3064);
and U13222 (N_13222,N_3323,N_9358);
and U13223 (N_13223,N_8405,N_6662);
nand U13224 (N_13224,N_7215,N_6208);
nor U13225 (N_13225,N_5221,N_4227);
nor U13226 (N_13226,N_3941,N_9217);
nor U13227 (N_13227,N_6235,N_3436);
xnor U13228 (N_13228,N_1495,N_6220);
and U13229 (N_13229,N_4529,N_316);
and U13230 (N_13230,N_5582,N_275);
nor U13231 (N_13231,N_2979,N_5236);
and U13232 (N_13232,N_3305,N_6999);
and U13233 (N_13233,N_7039,N_6239);
or U13234 (N_13234,N_7088,N_7370);
nor U13235 (N_13235,N_1314,N_8047);
xnor U13236 (N_13236,N_3889,N_5651);
and U13237 (N_13237,N_1973,N_9065);
or U13238 (N_13238,N_716,N_265);
nand U13239 (N_13239,N_1818,N_4540);
or U13240 (N_13240,N_3342,N_5907);
nand U13241 (N_13241,N_5905,N_4194);
nand U13242 (N_13242,N_1610,N_8700);
nor U13243 (N_13243,N_8947,N_2506);
and U13244 (N_13244,N_8008,N_1824);
and U13245 (N_13245,N_9339,N_130);
nand U13246 (N_13246,N_5247,N_6352);
nand U13247 (N_13247,N_137,N_8319);
xnor U13248 (N_13248,N_3464,N_4356);
nor U13249 (N_13249,N_710,N_2473);
and U13250 (N_13250,N_4911,N_6116);
or U13251 (N_13251,N_9858,N_9175);
xnor U13252 (N_13252,N_8389,N_7585);
nand U13253 (N_13253,N_1355,N_5306);
xnor U13254 (N_13254,N_1279,N_3951);
or U13255 (N_13255,N_3762,N_2948);
nand U13256 (N_13256,N_4885,N_2092);
or U13257 (N_13257,N_5226,N_2310);
or U13258 (N_13258,N_4600,N_5735);
nand U13259 (N_13259,N_5974,N_190);
nor U13260 (N_13260,N_614,N_8526);
nor U13261 (N_13261,N_4548,N_6890);
nand U13262 (N_13262,N_9411,N_2210);
nand U13263 (N_13263,N_3975,N_2063);
and U13264 (N_13264,N_2728,N_5448);
or U13265 (N_13265,N_8053,N_3428);
nor U13266 (N_13266,N_5222,N_1127);
xnor U13267 (N_13267,N_1662,N_5357);
nor U13268 (N_13268,N_4233,N_926);
and U13269 (N_13269,N_4691,N_3877);
or U13270 (N_13270,N_2170,N_7342);
or U13271 (N_13271,N_9944,N_918);
and U13272 (N_13272,N_5709,N_4945);
or U13273 (N_13273,N_6940,N_801);
nor U13274 (N_13274,N_1947,N_9472);
nor U13275 (N_13275,N_2031,N_1829);
nand U13276 (N_13276,N_5739,N_5662);
and U13277 (N_13277,N_6001,N_3717);
xnor U13278 (N_13278,N_2025,N_4360);
or U13279 (N_13279,N_110,N_6407);
nand U13280 (N_13280,N_6801,N_6425);
or U13281 (N_13281,N_9259,N_4682);
and U13282 (N_13282,N_481,N_4623);
and U13283 (N_13283,N_2039,N_8983);
and U13284 (N_13284,N_5785,N_5779);
or U13285 (N_13285,N_7952,N_4400);
or U13286 (N_13286,N_9987,N_9560);
xnor U13287 (N_13287,N_6409,N_7369);
nand U13288 (N_13288,N_6735,N_8868);
or U13289 (N_13289,N_530,N_4935);
or U13290 (N_13290,N_5512,N_1282);
nor U13291 (N_13291,N_266,N_6753);
nand U13292 (N_13292,N_171,N_4127);
and U13293 (N_13293,N_2529,N_3575);
and U13294 (N_13294,N_7851,N_7603);
and U13295 (N_13295,N_3893,N_9519);
and U13296 (N_13296,N_8179,N_8314);
nand U13297 (N_13297,N_9228,N_1073);
nor U13298 (N_13298,N_3266,N_9815);
or U13299 (N_13299,N_5280,N_23);
nand U13300 (N_13300,N_6104,N_1093);
nand U13301 (N_13301,N_6507,N_1558);
or U13302 (N_13302,N_9327,N_9150);
nand U13303 (N_13303,N_9767,N_1012);
xnor U13304 (N_13304,N_6404,N_7993);
nor U13305 (N_13305,N_145,N_8655);
nand U13306 (N_13306,N_5114,N_6578);
or U13307 (N_13307,N_6032,N_9397);
or U13308 (N_13308,N_3518,N_1778);
or U13309 (N_13309,N_2543,N_6025);
nand U13310 (N_13310,N_6573,N_5961);
nor U13311 (N_13311,N_6479,N_1346);
or U13312 (N_13312,N_6764,N_7121);
nand U13313 (N_13313,N_7640,N_9710);
or U13314 (N_13314,N_6475,N_7079);
or U13315 (N_13315,N_1663,N_6888);
or U13316 (N_13316,N_2565,N_7627);
or U13317 (N_13317,N_6009,N_2048);
nand U13318 (N_13318,N_4310,N_4575);
nor U13319 (N_13319,N_2470,N_9799);
nor U13320 (N_13320,N_7364,N_2605);
nand U13321 (N_13321,N_8459,N_5127);
and U13322 (N_13322,N_1541,N_4300);
nor U13323 (N_13323,N_5659,N_6229);
nor U13324 (N_13324,N_6926,N_7135);
and U13325 (N_13325,N_7711,N_5734);
nand U13326 (N_13326,N_85,N_3807);
or U13327 (N_13327,N_9729,N_7692);
nor U13328 (N_13328,N_3542,N_1892);
xnor U13329 (N_13329,N_3929,N_8842);
nand U13330 (N_13330,N_5447,N_8528);
nor U13331 (N_13331,N_6169,N_7047);
or U13332 (N_13332,N_9030,N_6631);
nor U13333 (N_13333,N_353,N_7307);
and U13334 (N_13334,N_1510,N_4460);
or U13335 (N_13335,N_3443,N_8020);
nand U13336 (N_13336,N_4283,N_1242);
nor U13337 (N_13337,N_3892,N_8790);
and U13338 (N_13338,N_1996,N_8804);
nand U13339 (N_13339,N_1424,N_8157);
nand U13340 (N_13340,N_3357,N_7256);
nor U13341 (N_13341,N_9460,N_4427);
xor U13342 (N_13342,N_5798,N_2515);
and U13343 (N_13343,N_6092,N_8168);
and U13344 (N_13344,N_2744,N_4369);
nor U13345 (N_13345,N_8509,N_2644);
xnor U13346 (N_13346,N_7586,N_9227);
or U13347 (N_13347,N_2674,N_1007);
nor U13348 (N_13348,N_8227,N_1928);
nor U13349 (N_13349,N_8257,N_6721);
nand U13350 (N_13350,N_2102,N_6889);
nor U13351 (N_13351,N_4083,N_336);
xor U13352 (N_13352,N_9133,N_8854);
nand U13353 (N_13353,N_995,N_9047);
xor U13354 (N_13354,N_8210,N_6965);
or U13355 (N_13355,N_1835,N_6811);
nand U13356 (N_13356,N_5838,N_7445);
xnor U13357 (N_13357,N_3007,N_8682);
nor U13358 (N_13358,N_8687,N_4409);
xnor U13359 (N_13359,N_4165,N_1144);
or U13360 (N_13360,N_3715,N_6192);
or U13361 (N_13361,N_7279,N_2351);
and U13362 (N_13362,N_1056,N_5374);
or U13363 (N_13363,N_7722,N_4618);
nand U13364 (N_13364,N_594,N_4211);
or U13365 (N_13365,N_3184,N_2966);
or U13366 (N_13366,N_9912,N_1696);
nand U13367 (N_13367,N_8096,N_5415);
xnor U13368 (N_13368,N_532,N_5729);
nand U13369 (N_13369,N_1292,N_4193);
xnor U13370 (N_13370,N_9577,N_9013);
nor U13371 (N_13371,N_2180,N_895);
and U13372 (N_13372,N_7045,N_7547);
or U13373 (N_13373,N_840,N_578);
nor U13374 (N_13374,N_3267,N_6992);
xor U13375 (N_13375,N_881,N_285);
nor U13376 (N_13376,N_3254,N_4218);
nor U13377 (N_13377,N_191,N_2055);
nand U13378 (N_13378,N_9655,N_5728);
and U13379 (N_13379,N_5549,N_8935);
nand U13380 (N_13380,N_4492,N_1326);
nand U13381 (N_13381,N_4912,N_9784);
nand U13382 (N_13382,N_5867,N_743);
nand U13383 (N_13383,N_7357,N_4377);
and U13384 (N_13384,N_136,N_3106);
and U13385 (N_13385,N_4567,N_4137);
and U13386 (N_13386,N_1709,N_5608);
nand U13387 (N_13387,N_234,N_9080);
nand U13388 (N_13388,N_7458,N_4841);
and U13389 (N_13389,N_7336,N_8115);
xor U13390 (N_13390,N_3591,N_4927);
or U13391 (N_13391,N_3825,N_9094);
xnor U13392 (N_13392,N_172,N_4673);
nand U13393 (N_13393,N_3669,N_165);
or U13394 (N_13394,N_1143,N_944);
and U13395 (N_13395,N_3502,N_7724);
xor U13396 (N_13396,N_7174,N_5377);
nand U13397 (N_13397,N_8900,N_544);
or U13398 (N_13398,N_990,N_9539);
or U13399 (N_13399,N_8382,N_2443);
or U13400 (N_13400,N_3280,N_9983);
and U13401 (N_13401,N_9120,N_1886);
nand U13402 (N_13402,N_5572,N_6559);
nand U13403 (N_13403,N_7209,N_7103);
and U13404 (N_13404,N_6112,N_7532);
nor U13405 (N_13405,N_6780,N_7834);
nand U13406 (N_13406,N_5820,N_1048);
nor U13407 (N_13407,N_4152,N_1178);
or U13408 (N_13408,N_505,N_4723);
or U13409 (N_13409,N_1044,N_1536);
or U13410 (N_13410,N_3137,N_4589);
or U13411 (N_13411,N_9148,N_7805);
and U13412 (N_13412,N_1458,N_6891);
nand U13413 (N_13413,N_8504,N_9758);
nor U13414 (N_13414,N_8390,N_8636);
nand U13415 (N_13415,N_1656,N_9027);
or U13416 (N_13416,N_7406,N_7807);
and U13417 (N_13417,N_7151,N_1762);
nor U13418 (N_13418,N_9564,N_4762);
and U13419 (N_13419,N_6013,N_2240);
nor U13420 (N_13420,N_2869,N_446);
nand U13421 (N_13421,N_8718,N_9587);
or U13422 (N_13422,N_744,N_4052);
and U13423 (N_13423,N_9766,N_4996);
nor U13424 (N_13424,N_2429,N_2391);
nand U13425 (N_13425,N_1636,N_6566);
xnor U13426 (N_13426,N_5796,N_8241);
nand U13427 (N_13427,N_5498,N_2872);
and U13428 (N_13428,N_5138,N_914);
and U13429 (N_13429,N_2042,N_3927);
nor U13430 (N_13430,N_7566,N_33);
or U13431 (N_13431,N_4595,N_2879);
nand U13432 (N_13432,N_7330,N_4780);
nor U13433 (N_13433,N_6722,N_8281);
nor U13434 (N_13434,N_5783,N_2593);
or U13435 (N_13435,N_1421,N_1650);
nor U13436 (N_13436,N_2027,N_6302);
xor U13437 (N_13437,N_5979,N_1023);
nand U13438 (N_13438,N_533,N_8273);
and U13439 (N_13439,N_8239,N_6189);
nor U13440 (N_13440,N_5213,N_348);
nor U13441 (N_13441,N_3994,N_9161);
xor U13442 (N_13442,N_7833,N_644);
nand U13443 (N_13443,N_8103,N_9816);
nor U13444 (N_13444,N_8377,N_203);
xnor U13445 (N_13445,N_7860,N_5147);
and U13446 (N_13446,N_5599,N_7937);
or U13447 (N_13447,N_7343,N_2343);
and U13448 (N_13448,N_3313,N_8081);
or U13449 (N_13449,N_4646,N_3087);
or U13450 (N_13450,N_3445,N_5425);
or U13451 (N_13451,N_7598,N_7516);
xor U13452 (N_13452,N_4201,N_1582);
nor U13453 (N_13453,N_5090,N_8554);
nand U13454 (N_13454,N_3163,N_1051);
nand U13455 (N_13455,N_9852,N_6822);
and U13456 (N_13456,N_6179,N_4172);
or U13457 (N_13457,N_7266,N_5565);
and U13458 (N_13458,N_2274,N_9138);
and U13459 (N_13459,N_3679,N_569);
or U13460 (N_13460,N_8035,N_2512);
nor U13461 (N_13461,N_3888,N_8533);
or U13462 (N_13462,N_1645,N_7158);
nor U13463 (N_13463,N_1569,N_5229);
nand U13464 (N_13464,N_5665,N_5101);
nand U13465 (N_13465,N_2103,N_4829);
nand U13466 (N_13466,N_9166,N_8561);
or U13467 (N_13467,N_1132,N_2234);
and U13468 (N_13468,N_1605,N_3301);
nand U13469 (N_13469,N_4493,N_2988);
nand U13470 (N_13470,N_4506,N_5705);
nand U13471 (N_13471,N_3480,N_2926);
or U13472 (N_13472,N_8376,N_5527);
and U13473 (N_13473,N_4768,N_8154);
nand U13474 (N_13474,N_8930,N_519);
nor U13475 (N_13475,N_3534,N_1725);
and U13476 (N_13476,N_6012,N_86);
or U13477 (N_13477,N_3635,N_5327);
nand U13478 (N_13478,N_1266,N_4577);
nand U13479 (N_13479,N_2071,N_9186);
or U13480 (N_13480,N_3237,N_3441);
nand U13481 (N_13481,N_9540,N_1673);
and U13482 (N_13482,N_3014,N_2557);
nor U13483 (N_13483,N_882,N_9867);
and U13484 (N_13484,N_1261,N_763);
nor U13485 (N_13485,N_9705,N_2558);
xnor U13486 (N_13486,N_2899,N_81);
or U13487 (N_13487,N_1664,N_5129);
or U13488 (N_13488,N_4704,N_4223);
nor U13489 (N_13489,N_5091,N_2387);
and U13490 (N_13490,N_5872,N_2100);
xnor U13491 (N_13491,N_2861,N_6904);
nand U13492 (N_13492,N_5174,N_2640);
nand U13493 (N_13493,N_3382,N_1906);
nand U13494 (N_13494,N_2776,N_7844);
or U13495 (N_13495,N_6591,N_9135);
and U13496 (N_13496,N_7580,N_2018);
or U13497 (N_13497,N_792,N_8145);
and U13498 (N_13498,N_6290,N_6650);
or U13499 (N_13499,N_8633,N_9302);
xor U13500 (N_13500,N_6424,N_853);
and U13501 (N_13501,N_6856,N_6090);
nand U13502 (N_13502,N_558,N_4167);
or U13503 (N_13503,N_5012,N_3538);
nand U13504 (N_13504,N_2166,N_2820);
nand U13505 (N_13505,N_9231,N_8746);
nor U13506 (N_13506,N_7305,N_14);
nor U13507 (N_13507,N_8855,N_3165);
nor U13508 (N_13508,N_3082,N_256);
or U13509 (N_13509,N_572,N_5952);
and U13510 (N_13510,N_1608,N_7219);
nor U13511 (N_13511,N_3885,N_27);
nor U13512 (N_13512,N_2551,N_6510);
and U13513 (N_13513,N_4502,N_5676);
and U13514 (N_13514,N_8268,N_615);
nor U13515 (N_13515,N_63,N_7131);
nor U13516 (N_13516,N_8311,N_1516);
nor U13517 (N_13517,N_8349,N_9891);
nand U13518 (N_13518,N_7395,N_5679);
and U13519 (N_13519,N_4399,N_6637);
xor U13520 (N_13520,N_4449,N_9229);
and U13521 (N_13521,N_8123,N_3201);
nand U13522 (N_13522,N_7093,N_1488);
or U13523 (N_13523,N_5805,N_7214);
and U13524 (N_13524,N_6579,N_9254);
nand U13525 (N_13525,N_6428,N_6793);
or U13526 (N_13526,N_3824,N_5259);
nand U13527 (N_13527,N_2263,N_3566);
and U13528 (N_13528,N_349,N_2451);
or U13529 (N_13529,N_2964,N_9478);
nor U13530 (N_13530,N_7709,N_6256);
and U13531 (N_13531,N_5404,N_2976);
nand U13532 (N_13532,N_4202,N_524);
nor U13533 (N_13533,N_1840,N_3974);
or U13534 (N_13534,N_9809,N_6130);
or U13535 (N_13535,N_6732,N_7696);
nor U13536 (N_13536,N_6546,N_5697);
and U13537 (N_13537,N_9418,N_6476);
nor U13538 (N_13538,N_6381,N_6391);
nor U13539 (N_13539,N_4708,N_9123);
nand U13540 (N_13540,N_9486,N_7817);
xnor U13541 (N_13541,N_6373,N_5214);
nand U13542 (N_13542,N_2317,N_2347);
nand U13543 (N_13543,N_2459,N_3296);
or U13544 (N_13544,N_1267,N_329);
or U13545 (N_13545,N_5504,N_3039);
nand U13546 (N_13546,N_2850,N_8822);
xnor U13547 (N_13547,N_7110,N_6019);
or U13548 (N_13548,N_3971,N_1826);
and U13549 (N_13549,N_5887,N_4827);
or U13550 (N_13550,N_399,N_2732);
nor U13551 (N_13551,N_7531,N_8886);
nand U13552 (N_13552,N_6434,N_2167);
or U13553 (N_13553,N_496,N_6693);
or U13554 (N_13554,N_3814,N_3351);
nor U13555 (N_13555,N_7155,N_9663);
nor U13556 (N_13556,N_7710,N_4161);
nor U13557 (N_13557,N_2989,N_9037);
xor U13558 (N_13558,N_9654,N_6810);
nor U13559 (N_13559,N_521,N_7025);
nand U13560 (N_13560,N_8491,N_8780);
nand U13561 (N_13561,N_4220,N_6095);
or U13562 (N_13562,N_7480,N_7941);
and U13563 (N_13563,N_8831,N_8620);
or U13564 (N_13564,N_7733,N_6850);
nand U13565 (N_13565,N_6376,N_874);
and U13566 (N_13566,N_9063,N_1396);
or U13567 (N_13567,N_4224,N_6073);
or U13568 (N_13568,N_4089,N_9134);
or U13569 (N_13569,N_1678,N_3581);
nand U13570 (N_13570,N_5224,N_2260);
and U13571 (N_13571,N_9372,N_5910);
nor U13572 (N_13572,N_7820,N_9980);
or U13573 (N_13573,N_667,N_8591);
nor U13574 (N_13574,N_5239,N_7235);
or U13575 (N_13575,N_9739,N_6481);
or U13576 (N_13576,N_2448,N_8030);
nor U13577 (N_13577,N_3271,N_3938);
and U13578 (N_13578,N_2880,N_9062);
nand U13579 (N_13579,N_4873,N_3870);
and U13580 (N_13580,N_9173,N_3600);
nor U13581 (N_13581,N_2375,N_6639);
and U13582 (N_13582,N_5941,N_3813);
xor U13583 (N_13583,N_8407,N_3236);
nor U13584 (N_13584,N_3344,N_1524);
or U13585 (N_13585,N_1856,N_8906);
nand U13586 (N_13586,N_8496,N_6858);
nor U13587 (N_13587,N_3094,N_9072);
nand U13588 (N_13588,N_6117,N_3373);
and U13589 (N_13589,N_5667,N_6056);
and U13590 (N_13590,N_6401,N_7891);
xor U13591 (N_13591,N_9714,N_6333);
and U13592 (N_13592,N_2752,N_2053);
or U13593 (N_13593,N_3771,N_5510);
nor U13594 (N_13594,N_9414,N_9086);
and U13595 (N_13595,N_8171,N_9300);
and U13596 (N_13596,N_311,N_3177);
nand U13597 (N_13597,N_5947,N_9555);
nand U13598 (N_13598,N_1613,N_4317);
xor U13599 (N_13599,N_5634,N_8259);
and U13600 (N_13600,N_7411,N_1603);
and U13601 (N_13601,N_3708,N_1183);
nor U13602 (N_13602,N_6050,N_4676);
and U13603 (N_13603,N_3358,N_6512);
nand U13604 (N_13604,N_8560,N_2358);
or U13605 (N_13605,N_8360,N_2970);
or U13606 (N_13606,N_2341,N_3605);
nand U13607 (N_13607,N_1795,N_7786);
nor U13608 (N_13608,N_328,N_8594);
nor U13609 (N_13609,N_7797,N_3942);
nand U13610 (N_13610,N_2733,N_769);
or U13611 (N_13611,N_696,N_2553);
nor U13612 (N_13612,N_4350,N_9176);
or U13613 (N_13613,N_1448,N_953);
nand U13614 (N_13614,N_6498,N_9383);
nand U13615 (N_13615,N_8970,N_8738);
and U13616 (N_13616,N_9976,N_3576);
and U13617 (N_13617,N_9149,N_2178);
nor U13618 (N_13618,N_2157,N_5471);
and U13619 (N_13619,N_4077,N_1274);
nand U13620 (N_13620,N_1439,N_6754);
nand U13621 (N_13621,N_4328,N_7487);
nor U13622 (N_13622,N_9102,N_9079);
nor U13623 (N_13623,N_6894,N_4526);
and U13624 (N_13624,N_2662,N_6713);
nor U13625 (N_13625,N_258,N_6528);
and U13626 (N_13626,N_8473,N_4836);
and U13627 (N_13627,N_832,N_1793);
nor U13628 (N_13628,N_3993,N_9289);
and U13629 (N_13629,N_5330,N_7533);
and U13630 (N_13630,N_2912,N_1315);
or U13631 (N_13631,N_6191,N_4658);
or U13632 (N_13632,N_5771,N_3451);
or U13633 (N_13633,N_1971,N_1001);
and U13634 (N_13634,N_5274,N_1665);
or U13635 (N_13635,N_4716,N_4882);
nor U13636 (N_13636,N_9651,N_1283);
and U13637 (N_13637,N_4918,N_929);
nor U13638 (N_13638,N_426,N_1272);
and U13639 (N_13639,N_9525,N_7847);
or U13640 (N_13640,N_8928,N_398);
and U13641 (N_13641,N_2843,N_6051);
or U13642 (N_13642,N_5958,N_8704);
xnor U13643 (N_13643,N_7077,N_826);
nand U13644 (N_13644,N_4039,N_1891);
and U13645 (N_13645,N_7204,N_3136);
or U13646 (N_13646,N_3788,N_3046);
and U13647 (N_13647,N_6467,N_347);
and U13648 (N_13648,N_5422,N_6496);
and U13649 (N_13649,N_7241,N_5151);
or U13650 (N_13650,N_7721,N_3385);
nor U13651 (N_13651,N_4470,N_4942);
nor U13652 (N_13652,N_1633,N_7698);
nand U13653 (N_13653,N_1922,N_7791);
and U13654 (N_13654,N_4831,N_7484);
and U13655 (N_13655,N_3867,N_5812);
and U13656 (N_13656,N_2447,N_7007);
xnor U13657 (N_13657,N_2875,N_6618);
nor U13658 (N_13658,N_2047,N_4782);
or U13659 (N_13659,N_6569,N_5107);
nor U13660 (N_13660,N_189,N_8391);
or U13661 (N_13661,N_8277,N_5301);
or U13662 (N_13662,N_6149,N_3497);
or U13663 (N_13663,N_5007,N_9402);
nand U13664 (N_13664,N_4198,N_2397);
nand U13665 (N_13665,N_112,N_8841);
nand U13666 (N_13666,N_512,N_1883);
nor U13667 (N_13667,N_9266,N_8787);
and U13668 (N_13668,N_8669,N_513);
or U13669 (N_13669,N_4367,N_1659);
or U13670 (N_13670,N_6838,N_9972);
and U13671 (N_13671,N_2072,N_9755);
xor U13672 (N_13672,N_7694,N_6035);
nand U13673 (N_13673,N_1133,N_499);
or U13674 (N_13674,N_8275,N_5159);
nor U13675 (N_13675,N_4289,N_6680);
nor U13676 (N_13676,N_3694,N_587);
or U13677 (N_13677,N_7024,N_8922);
nand U13678 (N_13678,N_4169,N_4250);
or U13679 (N_13679,N_6989,N_3255);
xnor U13680 (N_13680,N_3674,N_3403);
nor U13681 (N_13681,N_5031,N_3596);
and U13682 (N_13682,N_7159,N_2675);
and U13683 (N_13683,N_4254,N_8434);
nor U13684 (N_13684,N_3421,N_8090);
or U13685 (N_13685,N_1607,N_866);
and U13686 (N_13686,N_8681,N_9398);
and U13687 (N_13687,N_8597,N_5068);
and U13688 (N_13688,N_3514,N_2392);
and U13689 (N_13689,N_795,N_9258);
or U13690 (N_13690,N_5296,N_3197);
or U13691 (N_13691,N_4407,N_549);
xnor U13692 (N_13692,N_825,N_8361);
nand U13693 (N_13693,N_365,N_150);
or U13694 (N_13694,N_2070,N_5909);
nand U13695 (N_13695,N_4435,N_9688);
and U13696 (N_13696,N_6984,N_2932);
and U13697 (N_13697,N_9644,N_6576);
nor U13698 (N_13698,N_734,N_1407);
or U13699 (N_13699,N_346,N_6421);
or U13700 (N_13700,N_5552,N_1092);
xor U13701 (N_13701,N_3799,N_2476);
xnor U13702 (N_13702,N_1213,N_6319);
nor U13703 (N_13703,N_9162,N_3140);
or U13704 (N_13704,N_7433,N_6942);
nor U13705 (N_13705,N_1956,N_656);
and U13706 (N_13706,N_3414,N_7734);
nand U13707 (N_13707,N_8060,N_6048);
nor U13708 (N_13708,N_8293,N_4970);
nand U13709 (N_13709,N_6387,N_7512);
or U13710 (N_13710,N_3300,N_7041);
and U13711 (N_13711,N_1700,N_5762);
xor U13712 (N_13712,N_3772,N_1993);
nor U13713 (N_13713,N_8546,N_2748);
and U13714 (N_13714,N_6836,N_4415);
and U13715 (N_13715,N_4913,N_9953);
nand U13716 (N_13716,N_745,N_9330);
nor U13717 (N_13717,N_9308,N_1307);
nand U13718 (N_13718,N_3,N_5476);
or U13719 (N_13719,N_8725,N_7919);
xor U13720 (N_13720,N_2395,N_8815);
nor U13721 (N_13721,N_1865,N_1929);
and U13722 (N_13722,N_7732,N_2763);
or U13723 (N_13723,N_9810,N_8278);
or U13724 (N_13724,N_975,N_9716);
nor U13725 (N_13725,N_2916,N_1805);
and U13726 (N_13726,N_4741,N_4617);
or U13727 (N_13727,N_4825,N_8378);
nor U13728 (N_13728,N_5095,N_5333);
or U13729 (N_13729,N_69,N_1381);
nor U13730 (N_13730,N_9778,N_8988);
or U13731 (N_13731,N_7521,N_8479);
nor U13732 (N_13732,N_77,N_2720);
or U13733 (N_13733,N_6436,N_6364);
nand U13734 (N_13734,N_2091,N_9471);
and U13735 (N_13735,N_9702,N_2570);
nand U13736 (N_13736,N_5077,N_3568);
and U13737 (N_13737,N_9395,N_5741);
nand U13738 (N_13738,N_2364,N_9114);
nor U13739 (N_13739,N_7112,N_6060);
nor U13740 (N_13740,N_507,N_3925);
and U13741 (N_13741,N_8355,N_688);
and U13742 (N_13742,N_215,N_9549);
nor U13743 (N_13743,N_2462,N_4881);
xnor U13744 (N_13744,N_3188,N_5223);
and U13745 (N_13745,N_841,N_3822);
or U13746 (N_13746,N_4429,N_6139);
nand U13747 (N_13747,N_4327,N_6852);
or U13748 (N_13748,N_40,N_8236);
or U13749 (N_13749,N_4765,N_2247);
or U13750 (N_13750,N_114,N_3574);
nor U13751 (N_13751,N_6470,N_1291);
nor U13752 (N_13752,N_2330,N_1378);
and U13753 (N_13753,N_1788,N_663);
or U13754 (N_13754,N_8036,N_6597);
and U13755 (N_13755,N_8839,N_1720);
nor U13756 (N_13756,N_6738,N_4999);
nor U13757 (N_13757,N_564,N_6867);
and U13758 (N_13758,N_4657,N_8058);
xnor U13759 (N_13759,N_1038,N_8041);
and U13760 (N_13760,N_5965,N_9939);
and U13761 (N_13761,N_586,N_3125);
and U13762 (N_13762,N_5633,N_4404);
and U13763 (N_13763,N_1205,N_8882);
nor U13764 (N_13764,N_8867,N_7420);
xnor U13765 (N_13765,N_8383,N_9607);
nor U13766 (N_13766,N_278,N_174);
nand U13767 (N_13767,N_1204,N_5708);
nand U13768 (N_13768,N_9546,N_3257);
xnor U13769 (N_13769,N_635,N_6511);
nand U13770 (N_13770,N_8416,N_9585);
nand U13771 (N_13771,N_6648,N_1974);
nand U13772 (N_13772,N_8627,N_9034);
or U13773 (N_13773,N_2998,N_8129);
and U13774 (N_13774,N_2650,N_3272);
nor U13775 (N_13775,N_7761,N_7882);
or U13776 (N_13776,N_8689,N_8963);
nand U13777 (N_13777,N_774,N_5384);
or U13778 (N_13778,N_4654,N_1236);
xnor U13779 (N_13779,N_9604,N_3485);
and U13780 (N_13780,N_1491,N_3884);
nor U13781 (N_13781,N_9336,N_4812);
nand U13782 (N_13782,N_2276,N_8948);
nor U13783 (N_13783,N_4640,N_4503);
nand U13784 (N_13784,N_338,N_3863);
or U13785 (N_13785,N_5875,N_8943);
nor U13786 (N_13786,N_7451,N_7819);
nand U13787 (N_13787,N_6614,N_8399);
or U13788 (N_13788,N_5193,N_5761);
and U13789 (N_13789,N_9269,N_7056);
nor U13790 (N_13790,N_9335,N_3520);
nor U13791 (N_13791,N_4014,N_3719);
nand U13792 (N_13792,N_4732,N_8400);
nand U13793 (N_13793,N_3745,N_7927);
nor U13794 (N_13794,N_8651,N_1446);
nand U13795 (N_13795,N_1539,N_1194);
nand U13796 (N_13796,N_3907,N_548);
or U13797 (N_13797,N_4059,N_5657);
or U13798 (N_13798,N_6786,N_8001);
nor U13799 (N_13799,N_8497,N_3408);
or U13800 (N_13800,N_557,N_3164);
nor U13801 (N_13801,N_1126,N_541);
or U13802 (N_13802,N_5475,N_3006);
nand U13803 (N_13803,N_1874,N_9404);
nand U13804 (N_13804,N_5672,N_1138);
nor U13805 (N_13805,N_809,N_4587);
or U13806 (N_13806,N_7001,N_9188);
or U13807 (N_13807,N_4301,N_6950);
or U13808 (N_13808,N_554,N_4231);
and U13809 (N_13809,N_216,N_5071);
nand U13810 (N_13810,N_5176,N_5217);
nor U13811 (N_13811,N_5859,N_5877);
nand U13812 (N_13812,N_2532,N_4664);
or U13813 (N_13813,N_4798,N_7888);
nand U13814 (N_13814,N_3649,N_5194);
xor U13815 (N_13815,N_7208,N_1955);
or U13816 (N_13816,N_3921,N_9281);
nor U13817 (N_13817,N_5615,N_4139);
nand U13818 (N_13818,N_761,N_5824);
nor U13819 (N_13819,N_9616,N_5130);
nor U13820 (N_13820,N_5911,N_7610);
xnor U13821 (N_13821,N_4743,N_9434);
nor U13822 (N_13822,N_3472,N_6398);
and U13823 (N_13823,N_8567,N_4303);
nor U13824 (N_13824,N_5880,N_1498);
xor U13825 (N_13825,N_6296,N_7438);
nand U13826 (N_13826,N_8291,N_302);
and U13827 (N_13827,N_469,N_6990);
nand U13828 (N_13828,N_2904,N_6841);
nor U13829 (N_13829,N_6070,N_1862);
nand U13830 (N_13830,N_453,N_3332);
or U13831 (N_13831,N_8992,N_2020);
xor U13832 (N_13832,N_492,N_5567);
nand U13833 (N_13833,N_9824,N_3607);
nor U13834 (N_13834,N_9652,N_7428);
or U13835 (N_13835,N_3543,N_6960);
nor U13836 (N_13836,N_404,N_5635);
nor U13837 (N_13837,N_5707,N_6588);
nor U13838 (N_13838,N_4950,N_5901);
xnor U13839 (N_13839,N_4280,N_4181);
nor U13840 (N_13840,N_6137,N_5391);
and U13841 (N_13841,N_585,N_6380);
nand U13842 (N_13842,N_8142,N_8064);
nand U13843 (N_13843,N_9309,N_2407);
nor U13844 (N_13844,N_2320,N_8946);
nor U13845 (N_13845,N_2777,N_8);
nand U13846 (N_13846,N_1755,N_8118);
nand U13847 (N_13847,N_6426,N_7827);
nor U13848 (N_13848,N_8921,N_2978);
nor U13849 (N_13849,N_8474,N_4442);
and U13850 (N_13850,N_8617,N_6393);
nor U13851 (N_13851,N_9565,N_8968);
and U13852 (N_13852,N_7163,N_3139);
nor U13853 (N_13853,N_8989,N_4845);
nand U13854 (N_13854,N_3631,N_3285);
nand U13855 (N_13855,N_2130,N_1796);
and U13856 (N_13856,N_8680,N_1583);
nand U13857 (N_13857,N_5490,N_1702);
or U13858 (N_13858,N_2665,N_8795);
or U13859 (N_13859,N_3460,N_980);
and U13860 (N_13860,N_8847,N_8625);
nand U13861 (N_13861,N_2099,N_4902);
and U13862 (N_13862,N_4883,N_4187);
or U13863 (N_13863,N_4784,N_4615);
nor U13864 (N_13864,N_6181,N_6194);
nand U13865 (N_13865,N_9494,N_9179);
nor U13866 (N_13866,N_6514,N_2737);
nand U13867 (N_13867,N_2848,N_1919);
or U13868 (N_13868,N_5408,N_3112);
and U13869 (N_13869,N_9862,N_5716);
nand U13870 (N_13870,N_2444,N_9826);
nor U13871 (N_13871,N_122,N_257);
nor U13872 (N_13872,N_2885,N_7125);
xnor U13873 (N_13873,N_8359,N_5898);
nand U13874 (N_13874,N_896,N_6972);
or U13875 (N_13875,N_8856,N_9812);
or U13876 (N_13876,N_9360,N_9421);
or U13877 (N_13877,N_6748,N_1002);
or U13878 (N_13878,N_9484,N_6622);
and U13879 (N_13879,N_7958,N_5531);
and U13880 (N_13880,N_3023,N_6007);
nand U13881 (N_13881,N_9924,N_6788);
and U13882 (N_13882,N_8964,N_1742);
nand U13883 (N_13883,N_3904,N_2196);
or U13884 (N_13884,N_3333,N_2357);
and U13885 (N_13885,N_865,N_7255);
nand U13886 (N_13886,N_1958,N_4480);
nor U13887 (N_13887,N_488,N_9024);
xor U13888 (N_13888,N_3525,N_5334);
and U13889 (N_13889,N_4430,N_3482);
nand U13890 (N_13890,N_4900,N_3874);
xor U13891 (N_13891,N_6862,N_1026);
nand U13892 (N_13892,N_8532,N_7098);
and U13893 (N_13893,N_857,N_7413);
and U13894 (N_13894,N_7772,N_516);
and U13895 (N_13895,N_2349,N_242);
or U13896 (N_13896,N_2975,N_5034);
nor U13897 (N_13897,N_7443,N_7020);
and U13898 (N_13898,N_3362,N_2308);
nor U13899 (N_13899,N_9219,N_9205);
nand U13900 (N_13900,N_3361,N_5560);
and U13901 (N_13901,N_6047,N_4584);
xnor U13902 (N_13902,N_4858,N_5956);
and U13903 (N_13903,N_5978,N_1601);
or U13904 (N_13904,N_7381,N_7114);
and U13905 (N_13905,N_4153,N_6440);
or U13906 (N_13906,N_186,N_1552);
or U13907 (N_13907,N_7746,N_1066);
nand U13908 (N_13908,N_4993,N_4036);
xnor U13909 (N_13909,N_3317,N_3386);
or U13910 (N_13910,N_8903,N_6958);
or U13911 (N_13911,N_7776,N_647);
xnor U13912 (N_13912,N_755,N_6560);
or U13913 (N_13913,N_713,N_366);
nand U13914 (N_13914,N_2021,N_5703);
or U13915 (N_13915,N_939,N_5949);
xor U13916 (N_13916,N_1247,N_9368);
nor U13917 (N_13917,N_5321,N_8732);
and U13918 (N_13918,N_5650,N_4104);
or U13919 (N_13919,N_1514,N_2766);
xor U13920 (N_13920,N_3584,N_8450);
nand U13921 (N_13921,N_6138,N_1409);
nand U13922 (N_13922,N_6021,N_5444);
xor U13923 (N_13923,N_517,N_6762);
or U13924 (N_13924,N_6892,N_4974);
nand U13925 (N_13925,N_536,N_9147);
nor U13926 (N_13926,N_8691,N_1352);
and U13927 (N_13927,N_1398,N_5116);
nand U13928 (N_13928,N_1933,N_1149);
xnor U13929 (N_13929,N_4366,N_864);
nor U13930 (N_13930,N_2085,N_8066);
nand U13931 (N_13931,N_7072,N_8748);
xor U13932 (N_13932,N_3399,N_7152);
nor U13933 (N_13933,N_7008,N_1784);
xor U13934 (N_13934,N_4565,N_3582);
and U13935 (N_13935,N_5360,N_7190);
nand U13936 (N_13936,N_9829,N_1776);
and U13937 (N_13937,N_6395,N_2951);
nand U13938 (N_13938,N_4659,N_1868);
xnor U13939 (N_13939,N_8502,N_1310);
xnor U13940 (N_13940,N_6781,N_126);
or U13941 (N_13941,N_1921,N_5902);
xor U13942 (N_13942,N_4594,N_7046);
nor U13943 (N_13943,N_1041,N_244);
nand U13944 (N_13944,N_7325,N_1365);
nand U13945 (N_13945,N_6101,N_3792);
nor U13946 (N_13946,N_8873,N_4472);
nor U13947 (N_13947,N_7674,N_9103);
nand U13948 (N_13948,N_1965,N_2651);
nand U13949 (N_13949,N_7614,N_6248);
or U13950 (N_13950,N_3110,N_2798);
nand U13951 (N_13951,N_6531,N_6022);
or U13952 (N_13952,N_5821,N_9785);
nor U13953 (N_13953,N_4065,N_68);
and U13954 (N_13954,N_162,N_5344);
and U13955 (N_13955,N_514,N_6020);
or U13956 (N_13956,N_3881,N_620);
nor U13957 (N_13957,N_1869,N_1948);
nor U13958 (N_13958,N_8440,N_5006);
or U13959 (N_13959,N_784,N_3121);
nand U13960 (N_13960,N_537,N_6632);
nand U13961 (N_13961,N_2342,N_5037);
or U13962 (N_13962,N_8490,N_22);
nor U13963 (N_13963,N_3434,N_5348);
xor U13964 (N_13964,N_8544,N_6163);
and U13965 (N_13965,N_6845,N_274);
and U13966 (N_13966,N_9315,N_9026);
and U13967 (N_13967,N_9713,N_1687);
or U13968 (N_13968,N_661,N_1676);
and U13969 (N_13969,N_8661,N_443);
xnor U13970 (N_13970,N_473,N_6227);
nor U13971 (N_13971,N_9043,N_1475);
and U13972 (N_13972,N_5400,N_3062);
nor U13973 (N_13973,N_3134,N_6956);
nor U13974 (N_13974,N_6937,N_1470);
nand U13975 (N_13975,N_8500,N_6983);
and U13976 (N_13976,N_7904,N_1246);
nor U13977 (N_13977,N_7619,N_5555);
nor U13978 (N_13978,N_5981,N_2837);
or U13979 (N_13979,N_9947,N_8401);
nand U13980 (N_13980,N_2972,N_5325);
nand U13981 (N_13981,N_9774,N_272);
or U13982 (N_13982,N_9682,N_8956);
nor U13983 (N_13983,N_4071,N_2753);
or U13984 (N_13984,N_118,N_6794);
or U13985 (N_13985,N_5616,N_7689);
xor U13986 (N_13986,N_5170,N_7070);
nand U13987 (N_13987,N_5302,N_6607);
and U13988 (N_13988,N_5543,N_4500);
or U13989 (N_13989,N_5177,N_4949);
and U13990 (N_13990,N_2403,N_9341);
and U13991 (N_13991,N_477,N_629);
nor U13992 (N_13992,N_6649,N_9896);
nor U13993 (N_13993,N_2768,N_5957);
nand U13994 (N_13994,N_4823,N_6294);
and U13995 (N_13995,N_5950,N_6736);
nand U13996 (N_13996,N_3049,N_4479);
nand U13997 (N_13997,N_4099,N_8623);
or U13998 (N_13998,N_717,N_6084);
and U13999 (N_13999,N_3654,N_6223);
nand U14000 (N_14000,N_7708,N_954);
nor U14001 (N_14001,N_2458,N_4023);
nor U14002 (N_14002,N_8710,N_5532);
and U14003 (N_14003,N_1815,N_4471);
nor U14004 (N_14004,N_5126,N_6270);
nor U14005 (N_14005,N_1483,N_643);
xor U14006 (N_14006,N_6772,N_2080);
and U14007 (N_14007,N_7280,N_6583);
and U14008 (N_14008,N_4009,N_6178);
or U14009 (N_14009,N_7429,N_6385);
nor U14010 (N_14010,N_7430,N_6630);
xor U14011 (N_14011,N_5610,N_5428);
and U14012 (N_14012,N_4228,N_6577);
or U14013 (N_14013,N_673,N_5849);
nand U14014 (N_14014,N_9154,N_2327);
and U14015 (N_14015,N_3020,N_65);
or U14016 (N_14016,N_9861,N_8708);
or U14017 (N_14017,N_7464,N_2838);
xor U14018 (N_14018,N_3981,N_7431);
nand U14019 (N_14019,N_1121,N_2639);
nor U14020 (N_14020,N_4100,N_3700);
and U14021 (N_14021,N_6767,N_2751);
nor U14022 (N_14022,N_630,N_3380);
nand U14023 (N_14023,N_1984,N_5234);
nand U14024 (N_14024,N_5235,N_5878);
and U14025 (N_14025,N_5886,N_7230);
or U14026 (N_14026,N_3724,N_613);
or U14027 (N_14027,N_4372,N_3355);
xor U14028 (N_14028,N_1214,N_8910);
nor U14029 (N_14029,N_9545,N_3478);
or U14030 (N_14030,N_1767,N_5351);
nor U14031 (N_14031,N_9238,N_9543);
nor U14032 (N_14032,N_7082,N_8980);
nor U14033 (N_14033,N_3150,N_2893);
nand U14034 (N_14034,N_6268,N_2445);
nand U14035 (N_14035,N_8127,N_961);
or U14036 (N_14036,N_4096,N_2400);
and U14037 (N_14037,N_8072,N_7285);
and U14038 (N_14038,N_1748,N_2062);
and U14039 (N_14039,N_3179,N_7578);
nand U14040 (N_14040,N_2296,N_7907);
and U14041 (N_14041,N_6102,N_1185);
nor U14042 (N_14042,N_9718,N_9796);
nand U14043 (N_14043,N_7396,N_6301);
nand U14044 (N_14044,N_2054,N_9798);
and U14045 (N_14045,N_7359,N_9049);
or U14046 (N_14046,N_5435,N_1604);
xnor U14047 (N_14047,N_7416,N_2833);
nor U14048 (N_14048,N_9332,N_1103);
and U14049 (N_14049,N_5719,N_3416);
and U14050 (N_14050,N_6068,N_9111);
nand U14051 (N_14051,N_457,N_1418);
xnor U14052 (N_14052,N_5433,N_4554);
xor U14053 (N_14053,N_3387,N_197);
and U14054 (N_14054,N_9338,N_2258);
nor U14055 (N_14055,N_9085,N_4324);
nor U14056 (N_14056,N_3220,N_8119);
nor U14057 (N_14057,N_6993,N_9632);
or U14058 (N_14058,N_3465,N_4436);
nand U14059 (N_14059,N_9375,N_8887);
or U14060 (N_14060,N_8211,N_3533);
nand U14061 (N_14061,N_1067,N_7573);
nor U14062 (N_14062,N_9998,N_7254);
and U14063 (N_14063,N_2382,N_9839);
and U14064 (N_14064,N_4365,N_6524);
and U14065 (N_14065,N_4260,N_589);
and U14066 (N_14066,N_6066,N_7779);
xor U14067 (N_14067,N_4528,N_8424);
or U14068 (N_14068,N_973,N_5158);
or U14069 (N_14069,N_5328,N_5551);
nand U14070 (N_14070,N_6855,N_2693);
or U14071 (N_14071,N_7457,N_6369);
nand U14072 (N_14072,N_1680,N_3486);
nor U14073 (N_14073,N_6759,N_4775);
xnor U14074 (N_14074,N_3122,N_96);
or U14075 (N_14075,N_1032,N_1061);
or U14076 (N_14076,N_2056,N_7523);
or U14077 (N_14077,N_8032,N_5460);
nand U14078 (N_14078,N_4868,N_6610);
nand U14079 (N_14079,N_6107,N_5590);
or U14080 (N_14080,N_2844,N_9083);
nor U14081 (N_14081,N_2895,N_2531);
nand U14082 (N_14082,N_7935,N_1731);
and U14083 (N_14083,N_7748,N_276);
or U14084 (N_14084,N_5141,N_5993);
nor U14085 (N_14085,N_125,N_9830);
or U14086 (N_14086,N_3671,N_3303);
and U14087 (N_14087,N_4066,N_9929);
or U14088 (N_14088,N_1404,N_8705);
nor U14089 (N_14089,N_9000,N_1509);
nor U14090 (N_14090,N_6262,N_1657);
and U14091 (N_14091,N_4042,N_2344);
nor U14092 (N_14092,N_4082,N_5693);
or U14093 (N_14093,N_3498,N_7181);
and U14094 (N_14094,N_5530,N_9782);
nor U14095 (N_14095,N_3084,N_9407);
or U14096 (N_14096,N_9328,N_1589);
and U14097 (N_14097,N_1690,N_1624);
or U14098 (N_14098,N_8895,N_3681);
and U14099 (N_14099,N_2289,N_6299);
or U14100 (N_14100,N_8077,N_5211);
nand U14101 (N_14101,N_3051,N_8878);
nand U14102 (N_14102,N_2655,N_1717);
or U14103 (N_14103,N_9597,N_2207);
and U14104 (N_14104,N_1445,N_9248);
and U14105 (N_14105,N_1070,N_2406);
nor U14106 (N_14106,N_7632,N_3011);
and U14107 (N_14107,N_6303,N_7915);
nor U14108 (N_14108,N_2599,N_5594);
and U14109 (N_14109,N_1961,N_6382);
or U14110 (N_14110,N_2205,N_2005);
nand U14111 (N_14111,N_9738,N_9993);
nand U14112 (N_14112,N_9973,N_8205);
nand U14113 (N_14113,N_5931,N_9818);
xor U14114 (N_14114,N_8198,N_2930);
nand U14115 (N_14115,N_9578,N_5876);
nor U14116 (N_14116,N_4574,N_4191);
xnor U14117 (N_14117,N_3922,N_3404);
and U14118 (N_14118,N_7499,N_7119);
nor U14119 (N_14119,N_3785,N_6486);
nor U14120 (N_14120,N_4171,N_5054);
and U14121 (N_14121,N_2133,N_5416);
xnor U14122 (N_14122,N_946,N_9419);
or U14123 (N_14123,N_226,N_2814);
nand U14124 (N_14124,N_2952,N_8540);
and U14125 (N_14125,N_9384,N_3900);
nand U14126 (N_14126,N_3308,N_1941);
xor U14127 (N_14127,N_1926,N_1469);
or U14128 (N_14128,N_9881,N_6880);
xor U14129 (N_14129,N_3529,N_1342);
or U14130 (N_14130,N_5464,N_1622);
nand U14131 (N_14131,N_5491,N_1064);
or U14132 (N_14132,N_2455,N_981);
and U14133 (N_14133,N_6623,N_8460);
and U14134 (N_14134,N_2232,N_4133);
nor U14135 (N_14135,N_24,N_7522);
or U14136 (N_14136,N_8025,N_7638);
or U14137 (N_14137,N_3661,N_4817);
or U14138 (N_14138,N_3626,N_8248);
nor U14139 (N_14139,N_1812,N_5501);
xor U14140 (N_14140,N_1035,N_5505);
nor U14141 (N_14141,N_8812,N_4109);
nand U14142 (N_14142,N_7969,N_9350);
xor U14143 (N_14143,N_2291,N_8013);
and U14144 (N_14144,N_5133,N_7863);
nor U14145 (N_14145,N_4620,N_3744);
nor U14146 (N_14146,N_4015,N_6033);
and U14147 (N_14147,N_2967,N_5569);
nor U14148 (N_14148,N_8253,N_8702);
and U14149 (N_14149,N_2625,N_7878);
or U14150 (N_14150,N_2590,N_6228);
xor U14151 (N_14151,N_9923,N_3466);
nor U14152 (N_14152,N_9520,N_2876);
nor U14153 (N_14153,N_3004,N_982);
nor U14154 (N_14154,N_7372,N_1704);
nor U14155 (N_14155,N_7595,N_6336);
nor U14156 (N_14156,N_6804,N_4486);
and U14157 (N_14157,N_9406,N_3368);
xnor U14158 (N_14158,N_8925,N_5711);
or U14159 (N_14159,N_1822,N_5960);
or U14160 (N_14160,N_6087,N_6830);
or U14161 (N_14161,N_7288,N_6733);
and U14162 (N_14162,N_6160,N_8467);
or U14163 (N_14163,N_1557,N_7486);
nor U14164 (N_14164,N_9990,N_8151);
nand U14165 (N_14165,N_230,N_4748);
and U14166 (N_14166,N_1387,N_2567);
nor U14167 (N_14167,N_7097,N_8958);
and U14168 (N_14168,N_8667,N_4279);
nor U14169 (N_14169,N_9772,N_7737);
nor U14170 (N_14170,N_6633,N_3471);
or U14171 (N_14171,N_8084,N_6500);
nor U14172 (N_14172,N_2810,N_1257);
nor U14173 (N_14173,N_4095,N_325);
and U14174 (N_14174,N_5225,N_9595);
and U14175 (N_14175,N_7832,N_8612);
and U14176 (N_14176,N_7588,N_3119);
nor U14177 (N_14177,N_6420,N_1014);
and U14178 (N_14178,N_4960,N_3409);
and U14179 (N_14179,N_3340,N_592);
and U14180 (N_14180,N_4074,N_4362);
nand U14181 (N_14181,N_207,N_6282);
or U14182 (N_14182,N_3008,N_8904);
and U14183 (N_14183,N_824,N_781);
and U14184 (N_14184,N_5326,N_5079);
or U14185 (N_14185,N_4955,N_6156);
nand U14186 (N_14186,N_7482,N_3676);
or U14187 (N_14187,N_5906,N_7403);
or U14188 (N_14188,N_7150,N_3647);
or U14189 (N_14189,N_7840,N_8121);
nor U14190 (N_14190,N_8307,N_708);
and U14191 (N_14191,N_7771,N_2847);
or U14192 (N_14192,N_4662,N_1523);
and U14193 (N_14193,N_4579,N_8499);
xnor U14194 (N_14194,N_4736,N_9662);
and U14195 (N_14195,N_7393,N_92);
nand U14196 (N_14196,N_5759,N_6388);
nor U14197 (N_14197,N_1637,N_7118);
xor U14198 (N_14198,N_8492,N_3764);
or U14199 (N_14199,N_1137,N_2353);
nand U14200 (N_14200,N_5231,N_8310);
or U14201 (N_14201,N_1208,N_3811);
nand U14202 (N_14202,N_7929,N_1821);
or U14203 (N_14203,N_4434,N_6785);
and U14204 (N_14204,N_5373,N_1230);
nor U14205 (N_14205,N_3281,N_3860);
and U14206 (N_14206,N_3976,N_2422);
xor U14207 (N_14207,N_8284,N_5749);
and U14208 (N_14208,N_1571,N_3200);
nor U14209 (N_14209,N_447,N_3085);
or U14210 (N_14210,N_9981,N_6098);
or U14211 (N_14211,N_1860,N_2660);
nand U14212 (N_14212,N_143,N_9707);
or U14213 (N_14213,N_2149,N_8647);
nand U14214 (N_14214,N_4329,N_9371);
nor U14215 (N_14215,N_3696,N_6259);
and U14216 (N_14216,N_1647,N_7982);
xor U14217 (N_14217,N_5817,N_4766);
xor U14218 (N_14218,N_6041,N_4926);
and U14219 (N_14219,N_4688,N_9076);
or U14220 (N_14220,N_204,N_4550);
xor U14221 (N_14221,N_3384,N_5300);
nor U14222 (N_14222,N_4199,N_9042);
and U14223 (N_14223,N_5959,N_7004);
nor U14224 (N_14224,N_852,N_907);
nand U14225 (N_14225,N_8901,N_1411);
and U14226 (N_14226,N_1757,N_6643);
nand U14227 (N_14227,N_8570,N_768);
nand U14228 (N_14228,N_9904,N_3028);
or U14229 (N_14229,N_7662,N_9118);
nor U14230 (N_14230,N_9823,N_7738);
or U14231 (N_14231,N_4553,N_484);
nand U14232 (N_14232,N_7814,N_3776);
or U14233 (N_14233,N_5774,N_1330);
xnor U14234 (N_14234,N_5929,N_5439);
nor U14235 (N_14235,N_4556,N_4205);
nor U14236 (N_14236,N_4088,N_2919);
nand U14237 (N_14237,N_7796,N_7647);
and U14238 (N_14238,N_5636,N_1635);
nor U14239 (N_14239,N_7232,N_4353);
nor U14240 (N_14240,N_771,N_4650);
nand U14241 (N_14241,N_8945,N_1124);
and U14242 (N_14242,N_8010,N_1119);
nor U14243 (N_14243,N_2287,N_6100);
and U14244 (N_14244,N_7067,N_6609);
nor U14245 (N_14245,N_2620,N_6870);
nand U14246 (N_14246,N_1962,N_8701);
nor U14247 (N_14247,N_9215,N_7751);
or U14248 (N_14248,N_7950,N_3153);
or U14249 (N_14249,N_6252,N_9967);
or U14250 (N_14250,N_4859,N_5288);
nand U14251 (N_14251,N_8309,N_342);
or U14252 (N_14252,N_3656,N_5331);
or U14253 (N_14253,N_1182,N_2706);
nor U14254 (N_14254,N_504,N_6125);
nor U14255 (N_14255,N_6606,N_6042);
nand U14256 (N_14256,N_1193,N_5840);
nor U14257 (N_14257,N_6868,N_9602);
or U14258 (N_14258,N_3912,N_1303);
nand U14259 (N_14259,N_3035,N_1970);
xor U14260 (N_14260,N_44,N_1836);
or U14261 (N_14261,N_6075,N_5698);
nand U14262 (N_14262,N_6339,N_7602);
and U14263 (N_14263,N_6986,N_6948);
nand U14264 (N_14264,N_9606,N_8221);
or U14265 (N_14265,N_2468,N_6658);
nand U14266 (N_14266,N_3563,N_9307);
or U14267 (N_14267,N_3666,N_3488);
nand U14268 (N_14268,N_695,N_5607);
nor U14269 (N_14269,N_5392,N_1881);
nor U14270 (N_14270,N_3947,N_6800);
and U14271 (N_14271,N_6837,N_654);
and U14272 (N_14272,N_803,N_1029);
nor U14273 (N_14273,N_3790,N_3741);
nor U14274 (N_14274,N_8357,N_835);
or U14275 (N_14275,N_641,N_3779);
or U14276 (N_14276,N_1580,N_595);
and U14277 (N_14277,N_2323,N_6663);
nor U14278 (N_14278,N_1576,N_7918);
and U14279 (N_14279,N_7144,N_3952);
and U14280 (N_14280,N_299,N_890);
and U14281 (N_14281,N_9681,N_5414);
xor U14282 (N_14282,N_8572,N_8869);
nand U14283 (N_14283,N_9317,N_6515);
nand U14284 (N_14284,N_4919,N_304);
or U14285 (N_14285,N_2300,N_892);
nand U14286 (N_14286,N_709,N_3739);
xor U14287 (N_14287,N_78,N_20);
and U14288 (N_14288,N_6279,N_1097);
and U14289 (N_14289,N_4115,N_9661);
and U14290 (N_14290,N_1338,N_411);
nand U14291 (N_14291,N_7717,N_1674);
and U14292 (N_14292,N_5995,N_4884);
nor U14293 (N_14293,N_2700,N_7293);
nand U14294 (N_14294,N_2487,N_8890);
and U14295 (N_14295,N_9880,N_1814);
nand U14296 (N_14296,N_6405,N_2419);
and U14297 (N_14297,N_229,N_9468);
nand U14298 (N_14298,N_7688,N_7726);
xor U14299 (N_14299,N_9353,N_6495);
nor U14300 (N_14300,N_5519,N_4001);
nand U14301 (N_14301,N_1646,N_4499);
xor U14302 (N_14302,N_4176,N_6152);
nor U14303 (N_14303,N_8688,N_5861);
and U14304 (N_14304,N_2060,N_8874);
nor U14305 (N_14305,N_4558,N_9977);
and U14306 (N_14306,N_2298,N_3109);
or U14307 (N_14307,N_8235,N_5700);
nand U14308 (N_14308,N_407,N_1546);
nor U14309 (N_14309,N_6687,N_1323);
nand U14310 (N_14310,N_4805,N_4746);
nand U14311 (N_14311,N_6848,N_3573);
xor U14312 (N_14312,N_4120,N_2237);
nand U14313 (N_14313,N_7865,N_8649);
nand U14314 (N_14314,N_4871,N_4);
or U14315 (N_14315,N_6410,N_7801);
or U14316 (N_14316,N_7360,N_4376);
nand U14317 (N_14317,N_7320,N_762);
nor U14318 (N_14318,N_5748,N_1811);
xor U14319 (N_14319,N_856,N_4976);
nand U14320 (N_14320,N_6345,N_6058);
or U14321 (N_14321,N_2582,N_5737);
nor U14322 (N_14322,N_3558,N_8590);
nor U14323 (N_14323,N_1969,N_3157);
xor U14324 (N_14324,N_5714,N_3896);
xor U14325 (N_14325,N_7550,N_7029);
and U14326 (N_14326,N_1371,N_6346);
and U14327 (N_14327,N_8516,N_4045);
nand U14328 (N_14328,N_4712,N_9909);
nor U14329 (N_14329,N_5367,N_928);
or U14330 (N_14330,N_9884,N_6923);
nand U14331 (N_14331,N_2160,N_8585);
or U14332 (N_14332,N_1201,N_7363);
and U14333 (N_14333,N_3240,N_4142);
or U14334 (N_14334,N_5063,N_3044);
xnor U14335 (N_14335,N_3353,N_7116);
nand U14336 (N_14336,N_9648,N_1487);
or U14337 (N_14337,N_8932,N_119);
nand U14338 (N_14338,N_6594,N_3784);
and U14339 (N_14339,N_8439,N_2729);
and U14340 (N_14340,N_6803,N_837);
or U14341 (N_14341,N_4576,N_3841);
nor U14342 (N_14342,N_5431,N_8668);
xnor U14343 (N_14343,N_2581,N_7616);
nand U14344 (N_14344,N_5768,N_313);
or U14345 (N_14345,N_5087,N_5157);
and U14346 (N_14346,N_1790,N_2823);
nand U14347 (N_14347,N_957,N_3127);
or U14348 (N_14348,N_7378,N_8088);
or U14349 (N_14349,N_8843,N_1435);
and U14350 (N_14350,N_3427,N_4380);
nor U14351 (N_14351,N_4186,N_800);
nor U14352 (N_14352,N_6348,N_2513);
nor U14353 (N_14353,N_1055,N_5244);
and U14354 (N_14354,N_1732,N_6688);
or U14355 (N_14355,N_9297,N_6615);
xor U14356 (N_14356,N_640,N_6105);
and U14357 (N_14357,N_9694,N_6096);
and U14358 (N_14358,N_7824,N_4304);
or U14359 (N_14359,N_8707,N_400);
xnor U14360 (N_14360,N_5335,N_7169);
or U14361 (N_14361,N_5463,N_6411);
xnor U14362 (N_14362,N_8320,N_8588);
nor U14363 (N_14363,N_9573,N_7925);
nor U14364 (N_14364,N_294,N_6966);
or U14365 (N_14365,N_3897,N_5285);
xor U14366 (N_14366,N_1177,N_3429);
nand U14367 (N_14367,N_7247,N_4818);
and U14368 (N_14368,N_1694,N_3078);
nor U14369 (N_14369,N_4413,N_9288);
nor U14370 (N_14370,N_2415,N_7513);
and U14371 (N_14371,N_2306,N_9897);
nand U14372 (N_14372,N_2219,N_8879);
xor U14373 (N_14373,N_7718,N_7921);
and U14374 (N_14374,N_4678,N_9728);
nor U14375 (N_14375,N_8484,N_3587);
and U14376 (N_14376,N_8486,N_6328);
nand U14377 (N_14377,N_9498,N_5438);
and U14378 (N_14378,N_9432,N_5497);
and U14379 (N_14379,N_1628,N_3859);
or U14380 (N_14380,N_1670,N_1800);
and U14381 (N_14381,N_3979,N_8074);
or U14382 (N_14382,N_6305,N_5119);
nand U14383 (N_14383,N_3315,N_7141);
nor U14384 (N_14384,N_4189,N_2078);
nor U14385 (N_14385,N_2749,N_1894);
and U14386 (N_14386,N_3359,N_5462);
or U14387 (N_14387,N_6574,N_8338);
nand U14388 (N_14388,N_9009,N_8892);
and U14389 (N_14389,N_7344,N_2598);
and U14390 (N_14390,N_8737,N_8240);
and U14391 (N_14391,N_3850,N_5474);
nor U14392 (N_14392,N_3448,N_3142);
nor U14393 (N_14393,N_7117,N_6961);
nor U14394 (N_14394,N_3491,N_9230);
and U14395 (N_14395,N_9376,N_3749);
or U14396 (N_14396,N_2649,N_1253);
nor U14397 (N_14397,N_3523,N_3365);
nand U14398 (N_14398,N_422,N_2435);
or U14399 (N_14399,N_3977,N_5089);
nor U14400 (N_14400,N_6029,N_2826);
nor U14401 (N_14401,N_6341,N_3354);
or U14402 (N_14402,N_3204,N_9783);
nand U14403 (N_14403,N_879,N_8443);
or U14404 (N_14404,N_7469,N_2215);
and U14405 (N_14405,N_7682,N_2813);
or U14406 (N_14406,N_9099,N_4625);
nor U14407 (N_14407,N_9945,N_3178);
nor U14408 (N_14408,N_1117,N_3291);
nor U14409 (N_14409,N_690,N_8850);
or U14410 (N_14410,N_5275,N_421);
or U14411 (N_14411,N_3500,N_4402);
and U14412 (N_14412,N_4874,N_6457);
nor U14413 (N_14413,N_9542,N_993);
nand U14414 (N_14414,N_5964,N_7178);
nand U14415 (N_14415,N_9598,N_7058);
or U14416 (N_14416,N_5757,N_5765);
or U14417 (N_14417,N_9303,N_2746);
nand U14418 (N_14418,N_9698,N_6734);
or U14419 (N_14419,N_7715,N_1638);
or U14420 (N_14420,N_8793,N_6134);
nor U14421 (N_14421,N_4067,N_2762);
and U14422 (N_14422,N_7465,N_7991);
and U14423 (N_14423,N_8385,N_3048);
nor U14424 (N_14424,N_7556,N_3562);
nand U14425 (N_14425,N_1118,N_2033);
nand U14426 (N_14426,N_7251,N_9104);
nor U14427 (N_14427,N_1161,N_1081);
nor U14428 (N_14428,N_5310,N_440);
nor U14429 (N_14429,N_6561,N_2894);
or U14430 (N_14430,N_2437,N_6834);
or U14431 (N_14431,N_6527,N_7197);
or U14432 (N_14432,N_7392,N_3965);
nand U14433 (N_14433,N_746,N_4255);
and U14434 (N_14434,N_9589,N_3665);
and U14435 (N_14435,N_2851,N_2577);
and U14436 (N_14436,N_2953,N_202);
nor U14437 (N_14437,N_7011,N_9381);
nor U14438 (N_14438,N_1923,N_2842);
and U14439 (N_14439,N_1334,N_7321);
and U14440 (N_14440,N_823,N_5450);
and U14441 (N_14441,N_8846,N_5386);
and U14442 (N_14442,N_6954,N_6513);
and U14443 (N_14443,N_6742,N_1927);
xnor U14444 (N_14444,N_4889,N_4123);
or U14445 (N_14445,N_3985,N_8079);
or U14446 (N_14446,N_7858,N_6802);
nand U14447 (N_14447,N_9686,N_1111);
nand U14448 (N_14448,N_3729,N_333);
and U14449 (N_14449,N_6055,N_5924);
nor U14450 (N_14450,N_4544,N_6014);
nor U14451 (N_14451,N_4188,N_820);
and U14452 (N_14452,N_166,N_3097);
nand U14453 (N_14453,N_2602,N_4685);
xnor U14454 (N_14454,N_4242,N_1522);
nand U14455 (N_14455,N_5989,N_2340);
or U14456 (N_14456,N_9268,N_8203);
nand U14457 (N_14457,N_1203,N_3457);
xnor U14458 (N_14458,N_9933,N_4516);
nand U14459 (N_14459,N_2896,N_6912);
and U14460 (N_14460,N_723,N_4923);
nor U14461 (N_14461,N_2949,N_388);
or U14462 (N_14462,N_450,N_2318);
nand U14463 (N_14463,N_6307,N_2131);
xor U14464 (N_14464,N_1794,N_0);
nand U14465 (N_14465,N_4609,N_5036);
and U14466 (N_14466,N_8495,N_233);
nand U14467 (N_14467,N_6696,N_4630);
nand U14468 (N_14468,N_5819,N_339);
and U14469 (N_14469,N_4651,N_6539);
or U14470 (N_14470,N_8821,N_5304);
or U14471 (N_14471,N_6599,N_9473);
or U14472 (N_14472,N_4852,N_7323);
nor U14473 (N_14473,N_4998,N_6471);
or U14474 (N_14474,N_8858,N_4978);
and U14475 (N_14475,N_4549,N_9920);
and U14476 (N_14476,N_2637,N_8595);
nor U14477 (N_14477,N_3742,N_5143);
xor U14478 (N_14478,N_7762,N_7676);
nor U14479 (N_14479,N_8131,N_9888);
nor U14480 (N_14480,N_4647,N_9876);
nand U14481 (N_14481,N_9157,N_3462);
nor U14482 (N_14482,N_8178,N_8934);
nor U14483 (N_14483,N_2046,N_284);
or U14484 (N_14484,N_467,N_858);
nor U14485 (N_14485,N_7558,N_2315);
nor U14486 (N_14486,N_7498,N_156);
nand U14487 (N_14487,N_5266,N_1160);
nor U14488 (N_14488,N_4068,N_9770);
nand U14489 (N_14489,N_1074,N_1366);
nor U14490 (N_14490,N_5574,N_7017);
nand U14491 (N_14491,N_1157,N_5270);
and U14492 (N_14492,N_5526,N_4720);
nor U14493 (N_14493,N_2209,N_3998);
and U14494 (N_14494,N_3129,N_4251);
nor U14495 (N_14495,N_8853,N_4336);
nor U14496 (N_14496,N_1987,N_1660);
and U14497 (N_14497,N_6916,N_8247);
and U14498 (N_14498,N_9477,N_4642);
xor U14499 (N_14499,N_4382,N_7911);
nand U14500 (N_14500,N_3356,N_4541);
and U14501 (N_14501,N_9255,N_2866);
nor U14502 (N_14502,N_210,N_5359);
nor U14503 (N_14503,N_3957,N_7857);
and U14504 (N_14504,N_3908,N_2920);
or U14505 (N_14505,N_6114,N_8745);
nor U14506 (N_14506,N_4749,N_1057);
nand U14507 (N_14507,N_5076,N_97);
nor U14508 (N_14508,N_2950,N_8161);
or U14509 (N_14509,N_1087,N_5212);
nor U14510 (N_14510,N_6370,N_5070);
and U14511 (N_14511,N_2290,N_8140);
xor U14512 (N_14512,N_5004,N_5758);
nor U14513 (N_14513,N_1441,N_4315);
nor U14514 (N_14514,N_4755,N_3970);
or U14515 (N_14515,N_5380,N_9212);
nor U14516 (N_14516,N_5681,N_5345);
or U14517 (N_14517,N_4056,N_9914);
nand U14518 (N_14518,N_9293,N_8840);
and U14519 (N_14519,N_1339,N_4872);
or U14520 (N_14520,N_2806,N_3625);
nand U14521 (N_14521,N_4484,N_4957);
nand U14522 (N_14522,N_8397,N_5403);
nand U14523 (N_14523,N_9615,N_1710);
or U14524 (N_14524,N_3603,N_9342);
nand U14525 (N_14525,N_8664,N_4886);
nor U14526 (N_14526,N_3758,N_2483);
and U14527 (N_14527,N_5413,N_4956);
nand U14528 (N_14528,N_6355,N_7855);
and U14529 (N_14529,N_1146,N_1501);
nor U14530 (N_14530,N_2354,N_836);
or U14531 (N_14531,N_6677,N_2881);
and U14532 (N_14532,N_1047,N_1072);
nor U14533 (N_14533,N_4057,N_6040);
nand U14534 (N_14534,N_5587,N_1738);
nand U14535 (N_14535,N_6308,N_4390);
xnor U14536 (N_14536,N_2831,N_7511);
or U14537 (N_14537,N_9618,N_567);
or U14538 (N_14538,N_6835,N_8498);
nor U14539 (N_14539,N_9721,N_3453);
nor U14540 (N_14540,N_8406,N_5763);
nand U14541 (N_14541,N_1021,N_9763);
or U14542 (N_14542,N_1216,N_1280);
nor U14543 (N_14543,N_5256,N_3738);
or U14544 (N_14544,N_2015,N_2006);
nor U14545 (N_14545,N_6949,N_7419);
nand U14546 (N_14546,N_8999,N_6715);
and U14547 (N_14547,N_8799,N_9165);
or U14548 (N_14548,N_9496,N_4179);
and U14549 (N_14549,N_5314,N_9709);
xor U14550 (N_14550,N_2917,N_2199);
nor U14551 (N_14551,N_3645,N_6796);
nor U14552 (N_14552,N_5021,N_2038);
or U14553 (N_14553,N_383,N_1682);
and U14554 (N_14554,N_596,N_1925);
nand U14555 (N_14555,N_6664,N_5661);
xor U14556 (N_14556,N_851,N_7530);
and U14557 (N_14557,N_764,N_1296);
nor U14558 (N_14558,N_715,N_6118);
or U14559 (N_14559,N_3546,N_7864);
xnor U14560 (N_14560,N_7104,N_2958);
and U14561 (N_14561,N_5016,N_8034);
nand U14562 (N_14562,N_775,N_8454);
nand U14563 (N_14563,N_799,N_9697);
nand U14564 (N_14564,N_141,N_6861);
nand U14565 (N_14565,N_9301,N_3686);
or U14566 (N_14566,N_925,N_8860);
nand U14567 (N_14567,N_1036,N_4807);
nand U14568 (N_14568,N_9934,N_5787);
nor U14569 (N_14569,N_3278,N_9359);
or U14570 (N_14570,N_5890,N_5842);
or U14571 (N_14571,N_8318,N_5927);
or U14572 (N_14572,N_5811,N_1643);
and U14573 (N_14573,N_8286,N_3391);
or U14574 (N_14574,N_6313,N_9613);
or U14575 (N_14575,N_5324,N_4776);
and U14576 (N_14576,N_2760,N_5962);
xor U14577 (N_14577,N_5507,N_5208);
xor U14578 (N_14578,N_7809,N_5276);
and U14579 (N_14579,N_3721,N_8482);
nand U14580 (N_14580,N_7297,N_4760);
nor U14581 (N_14581,N_5084,N_8262);
and U14582 (N_14582,N_2249,N_3063);
and U14583 (N_14583,N_5776,N_7455);
and U14584 (N_14584,N_5382,N_6638);
or U14585 (N_14585,N_2526,N_7778);
and U14586 (N_14586,N_3752,N_3777);
nor U14587 (N_14587,N_5073,N_5039);
nor U14588 (N_14588,N_7199,N_8234);
nor U14589 (N_14589,N_9794,N_3972);
and U14590 (N_14590,N_8296,N_1553);
nand U14591 (N_14591,N_1337,N_4721);
and U14592 (N_14592,N_438,N_3290);
and U14593 (N_14593,N_4267,N_4546);
nand U14594 (N_14594,N_9673,N_79);
and U14595 (N_14595,N_2359,N_6859);
nand U14596 (N_14596,N_6,N_7968);
or U14597 (N_14597,N_8596,N_3322);
xnor U14598 (N_14598,N_8487,N_1413);
nand U14599 (N_14599,N_6147,N_3477);
or U14600 (N_14600,N_8040,N_540);
and U14601 (N_14601,N_4734,N_4533);
or U14602 (N_14602,N_4309,N_4636);
nor U14603 (N_14603,N_8998,N_7938);
and U14604 (N_14604,N_5459,N_6702);
nor U14605 (N_14605,N_4275,N_2028);
or U14606 (N_14606,N_808,N_5102);
and U14607 (N_14607,N_6430,N_4102);
nor U14608 (N_14608,N_4043,N_5814);
or U14609 (N_14609,N_7916,N_683);
nand U14610 (N_14610,N_9022,N_5745);
nand U14611 (N_14611,N_1077,N_340);
nand U14612 (N_14612,N_7989,N_6847);
or U14613 (N_14613,N_7057,N_912);
nor U14614 (N_14614,N_6069,N_3968);
nand U14615 (N_14615,N_4325,N_8106);
and U14616 (N_14616,N_902,N_8100);
nand U14617 (N_14617,N_1747,N_6646);
nor U14618 (N_14618,N_2588,N_8037);
nand U14619 (N_14619,N_9680,N_4735);
and U14620 (N_14620,N_3903,N_9863);
nor U14621 (N_14621,N_3706,N_5712);
nor U14622 (N_14622,N_5112,N_9059);
or U14623 (N_14623,N_8368,N_7917);
or U14624 (N_14624,N_5954,N_919);
or U14625 (N_14625,N_5209,N_4832);
nor U14626 (N_14626,N_8468,N_9532);
and U14627 (N_14627,N_335,N_1099);
nand U14628 (N_14628,N_1217,N_9930);
nand U14629 (N_14629,N_7584,N_3018);
nand U14630 (N_14630,N_5108,N_7579);
and U14631 (N_14631,N_7812,N_1154);
nand U14632 (N_14632,N_4835,N_8395);
and U14633 (N_14633,N_8143,N_2114);
nand U14634 (N_14634,N_9832,N_7555);
or U14635 (N_14635,N_7508,N_9627);
and U14636 (N_14636,N_8813,N_4252);
or U14637 (N_14637,N_9871,N_5167);
xnor U14638 (N_14638,N_5248,N_5482);
or U14639 (N_14639,N_5864,N_9198);
or U14640 (N_14640,N_5412,N_5105);
or U14641 (N_14641,N_3192,N_4633);
nor U14642 (N_14642,N_5609,N_5766);
nor U14643 (N_14643,N_6536,N_5052);
and U14644 (N_14644,N_6864,N_9531);
and U14645 (N_14645,N_3156,N_2897);
nor U14646 (N_14646,N_3740,N_1551);
nor U14647 (N_14647,N_4751,N_9687);
and U14648 (N_14648,N_5154,N_4963);
or U14649 (N_14649,N_1540,N_2546);
nor U14650 (N_14650,N_8634,N_4758);
and U14651 (N_14651,N_4126,N_9097);
xnor U14652 (N_14652,N_6338,N_2190);
or U14653 (N_14653,N_5791,N_2225);
and U14654 (N_14654,N_9596,N_4222);
nand U14655 (N_14655,N_170,N_1730);
nor U14656 (N_14656,N_2840,N_9801);
nor U14657 (N_14657,N_3213,N_6390);
nand U14658 (N_14658,N_4243,N_74);
and U14659 (N_14659,N_4296,N_2482);
xor U14660 (N_14660,N_3906,N_131);
and U14661 (N_14661,N_2817,N_2460);
or U14662 (N_14662,N_6644,N_1219);
and U14663 (N_14663,N_6454,N_3183);
xnor U14664 (N_14664,N_9975,N_4824);
or U14665 (N_14665,N_6774,N_2884);
or U14666 (N_14666,N_2288,N_1406);
nor U14667 (N_14667,N_7823,N_4718);
or U14668 (N_14668,N_6991,N_6739);
and U14669 (N_14669,N_9366,N_1186);
and U14670 (N_14670,N_822,N_4345);
or U14671 (N_14671,N_5132,N_2803);
nor U14672 (N_14672,N_1262,N_9448);
or U14673 (N_14673,N_8692,N_4983);
xor U14674 (N_14674,N_3475,N_2554);
and U14675 (N_14675,N_4197,N_267);
xnor U14676 (N_14676,N_4700,N_5596);
xor U14677 (N_14677,N_3560,N_5801);
nand U14678 (N_14678,N_9121,N_8741);
xor U14679 (N_14679,N_6154,N_686);
nor U14680 (N_14680,N_5869,N_9741);
or U14681 (N_14681,N_8866,N_3936);
nand U14682 (N_14682,N_1191,N_7475);
and U14683 (N_14683,N_1854,N_3098);
and U14684 (N_14684,N_7764,N_3537);
or U14685 (N_14685,N_8446,N_2564);
and U14686 (N_14686,N_4141,N_5508);
nand U14687 (N_14687,N_7006,N_5452);
nand U14688 (N_14688,N_9117,N_765);
nor U14689 (N_14689,N_1905,N_6568);
or U14690 (N_14690,N_7154,N_3096);
nor U14691 (N_14691,N_3836,N_4523);
nand U14692 (N_14692,N_3733,N_1420);
nor U14693 (N_14693,N_4406,N_1736);
nand U14694 (N_14694,N_1024,N_7599);
nor U14695 (N_14695,N_2556,N_6516);
nand U14696 (N_14696,N_4557,N_2965);
or U14697 (N_14697,N_87,N_4196);
nand U14698 (N_14698,N_5945,N_5131);
nor U14699 (N_14699,N_8937,N_4972);
xor U14700 (N_14700,N_6678,N_997);
nor U14701 (N_14701,N_5846,N_465);
or U14702 (N_14702,N_1440,N_2859);
nand U14703 (N_14703,N_1677,N_7488);
or U14704 (N_14704,N_605,N_3853);
nand U14705 (N_14705,N_7695,N_3624);
or U14706 (N_14706,N_8130,N_9866);
or U14707 (N_14707,N_3955,N_8272);
nor U14708 (N_14708,N_5028,N_1903);
nand U14709 (N_14709,N_7928,N_5595);
or U14710 (N_14710,N_1010,N_1907);
nand U14711 (N_14711,N_4914,N_8345);
and U14712 (N_14712,N_7861,N_4321);
and U14713 (N_14713,N_509,N_3090);
or U14714 (N_14714,N_4461,N_6397);
and U14715 (N_14715,N_8266,N_5149);
and U14716 (N_14716,N_9464,N_6293);
nor U14717 (N_14717,N_9703,N_2016);
nand U14718 (N_14718,N_6589,N_9002);
or U14719 (N_14719,N_7315,N_6203);
or U14720 (N_14720,N_5145,N_1870);
or U14721 (N_14721,N_3492,N_8902);
and U14722 (N_14722,N_6037,N_8105);
and U14723 (N_14723,N_8108,N_6289);
and U14724 (N_14724,N_7111,N_7427);
or U14725 (N_14725,N_3261,N_9659);
or U14726 (N_14726,N_7596,N_9748);
nand U14727 (N_14727,N_7236,N_4136);
or U14728 (N_14728,N_9984,N_626);
nor U14729 (N_14729,N_1920,N_4757);
or U14730 (N_14730,N_935,N_2261);
and U14731 (N_14731,N_7985,N_108);
or U14732 (N_14732,N_9433,N_1577);
and U14733 (N_14733,N_2338,N_5624);
and U14734 (N_14734,N_7792,N_9441);
nor U14735 (N_14735,N_2957,N_1301);
and U14736 (N_14736,N_6214,N_253);
xor U14737 (N_14737,N_6429,N_6488);
and U14738 (N_14738,N_5205,N_6269);
and U14739 (N_14739,N_4521,N_5350);
and U14740 (N_14740,N_6509,N_4925);
nand U14741 (N_14741,N_4024,N_794);
nand U14742 (N_14742,N_9811,N_2903);
nand U14743 (N_14743,N_3196,N_3080);
or U14744 (N_14744,N_3827,N_9108);
or U14745 (N_14745,N_3054,N_4834);
or U14746 (N_14746,N_1184,N_1529);
nor U14747 (N_14747,N_6249,N_4786);
or U14748 (N_14748,N_7220,N_2792);
nand U14749 (N_14749,N_2146,N_2669);
xnor U14750 (N_14750,N_6980,N_3879);
nand U14751 (N_14751,N_8991,N_9011);
nand U14752 (N_14752,N_7707,N_8744);
and U14753 (N_14753,N_4469,N_8598);
nor U14754 (N_14754,N_4037,N_5999);
nand U14755 (N_14755,N_7271,N_5900);
nand U14756 (N_14756,N_6538,N_9679);
nand U14757 (N_14757,N_7207,N_5309);
and U14758 (N_14758,N_4788,N_4555);
nand U14759 (N_14759,N_6660,N_2069);
nor U14760 (N_14760,N_4822,N_1995);
nor U14761 (N_14761,N_9051,N_4763);
nand U14762 (N_14762,N_2938,N_2326);
nand U14763 (N_14763,N_728,N_8431);
nand U14764 (N_14764,N_8760,N_5996);
nor U14765 (N_14765,N_5454,N_4508);
or U14766 (N_14766,N_9612,N_6386);
or U14767 (N_14767,N_4339,N_6697);
or U14768 (N_14768,N_8778,N_3670);
xor U14769 (N_14769,N_4347,N_863);
and U14770 (N_14770,N_8797,N_8228);
nand U14771 (N_14771,N_3653,N_9349);
and U14772 (N_14772,N_144,N_8337);
nor U14773 (N_14773,N_5568,N_3016);
and U14774 (N_14774,N_5189,N_6151);
nand U14775 (N_14775,N_8711,N_3295);
nor U14776 (N_14776,N_2328,N_2388);
xor U14777 (N_14777,N_8814,N_4412);
or U14778 (N_14778,N_2618,N_3765);
or U14779 (N_14779,N_7563,N_5571);
nor U14780 (N_14780,N_3638,N_9591);
xor U14781 (N_14781,N_1039,N_8924);
nor U14782 (N_14782,N_7719,N_8663);
or U14783 (N_14783,N_1852,N_2163);
and U14784 (N_14784,N_1231,N_9988);
or U14785 (N_14785,N_624,N_3754);
and U14786 (N_14786,N_3804,N_901);
and U14787 (N_14787,N_2208,N_1306);
nor U14788 (N_14788,N_5339,N_7524);
nand U14789 (N_14789,N_4610,N_3687);
and U14790 (N_14790,N_9141,N_5873);
or U14791 (N_14791,N_6238,N_4653);
nand U14792 (N_14792,N_1463,N_1086);
or U14793 (N_14793,N_632,N_2654);
nand U14794 (N_14794,N_5630,N_2410);
and U14795 (N_14795,N_2101,N_6314);
nor U14796 (N_14796,N_3494,N_5621);
and U14797 (N_14797,N_2993,N_7162);
nand U14798 (N_14798,N_7553,N_9510);
nor U14799 (N_14799,N_3260,N_7421);
or U14800 (N_14800,N_2723,N_6537);
nor U14801 (N_14801,N_5732,N_7229);
nand U14802 (N_14802,N_3845,N_4156);
and U14803 (N_14803,N_3155,N_561);
nor U14804 (N_14804,N_5639,N_7231);
and U14805 (N_14805,N_3580,N_5691);
nor U14806 (N_14806,N_2573,N_7276);
and U14807 (N_14807,N_2386,N_8729);
nor U14808 (N_14808,N_2627,N_5166);
nand U14809 (N_14809,N_1211,N_6317);
nor U14810 (N_14810,N_6879,N_9750);
or U14811 (N_14811,N_742,N_598);
xor U14812 (N_14812,N_6728,N_650);
or U14813 (N_14813,N_387,N_6866);
xnor U14814 (N_14814,N_466,N_4185);
nand U14815 (N_14815,N_4811,N_988);
nand U14816 (N_14816,N_1188,N_7391);
or U14817 (N_14817,N_2220,N_4216);
nand U14818 (N_14818,N_6292,N_2575);
nand U14819 (N_14819,N_2430,N_6634);
or U14820 (N_14820,N_5870,N_2352);
nand U14821 (N_14821,N_6700,N_622);
xor U14822 (N_14822,N_8033,N_9405);
or U14823 (N_14823,N_6418,N_4877);
or U14824 (N_14824,N_5668,N_1202);
and U14825 (N_14825,N_693,N_8201);
and U14826 (N_14826,N_9066,N_1946);
and U14827 (N_14827,N_1373,N_1872);
nor U14828 (N_14828,N_7613,N_4701);
or U14829 (N_14829,N_3328,N_2724);
and U14830 (N_14830,N_6003,N_7961);
xnor U14831 (N_14831,N_3890,N_1163);
and U14832 (N_14832,N_277,N_5181);
and U14833 (N_14833,N_4112,N_8193);
and U14834 (N_14834,N_4894,N_8961);
and U14835 (N_14835,N_2587,N_5120);
and U14836 (N_14836,N_4583,N_5186);
and U14837 (N_14837,N_3371,N_6645);
nand U14838 (N_14838,N_1621,N_5283);
or U14839 (N_14839,N_7582,N_8894);
nand U14840 (N_14840,N_1890,N_9732);
or U14841 (N_14841,N_2250,N_4977);
nor U14842 (N_14842,N_1042,N_3293);
nor U14843 (N_14843,N_6541,N_6122);
nand U14844 (N_14844,N_100,N_4119);
or U14845 (N_14845,N_3310,N_6604);
xor U14846 (N_14846,N_2822,N_9854);
nand U14847 (N_14847,N_9614,N_5281);
xnor U14848 (N_14848,N_9670,N_8611);
or U14849 (N_14849,N_8254,N_5480);
or U14850 (N_14850,N_5591,N_4454);
and U14851 (N_14851,N_8305,N_5780);
or U14852 (N_14852,N_4715,N_1591);
or U14853 (N_14853,N_2488,N_5461);
nor U14854 (N_14854,N_3505,N_7218);
nor U14855 (N_14855,N_61,N_5315);
and U14856 (N_14856,N_6444,N_4667);
and U14857 (N_14857,N_8478,N_3557);
xor U14858 (N_14858,N_9261,N_2);
and U14859 (N_14859,N_8402,N_5320);
and U14860 (N_14860,N_7237,N_5190);
nor U14861 (N_14861,N_3714,N_5175);
and U14862 (N_14862,N_2525,N_9348);
or U14863 (N_14863,N_8802,N_4241);
and U14864 (N_14864,N_2682,N_7075);
nor U14865 (N_14865,N_8806,N_7626);
nand U14866 (N_14866,N_47,N_802);
nor U14867 (N_14867,N_3548,N_5721);
nand U14868 (N_14868,N_6769,N_6553);
or U14869 (N_14869,N_6438,N_3703);
and U14870 (N_14870,N_2417,N_8417);
and U14871 (N_14871,N_1383,N_2827);
and U14872 (N_14872,N_7382,N_7339);
and U14873 (N_14873,N_1950,N_3887);
xnor U14874 (N_14874,N_8518,N_5082);
or U14875 (N_14875,N_4195,N_3682);
nand U14876 (N_14876,N_5185,N_6690);
or U14877 (N_14877,N_3532,N_5402);
xor U14878 (N_14878,N_7377,N_722);
and U14879 (N_14879,N_4520,N_9019);
and U14880 (N_14880,N_4314,N_7437);
and U14881 (N_14881,N_2982,N_9192);
nand U14882 (N_14882,N_6103,N_8420);
and U14883 (N_14883,N_712,N_4739);
or U14884 (N_14884,N_6121,N_4458);
or U14885 (N_14885,N_5602,N_5896);
or U14886 (N_14886,N_4905,N_838);
or U14887 (N_14887,N_26,N_4238);
nand U14888 (N_14888,N_8609,N_4371);
nor U14889 (N_14889,N_6925,N_115);
or U14890 (N_14890,N_5580,N_9409);
nor U14891 (N_14891,N_1031,N_9092);
and U14892 (N_14892,N_3103,N_71);
or U14893 (N_14893,N_5035,N_1867);
nand U14894 (N_14894,N_4038,N_7837);
or U14895 (N_14895,N_2614,N_1900);
or U14896 (N_14896,N_3911,N_5316);
nor U14897 (N_14897,N_5010,N_4107);
or U14898 (N_14898,N_7165,N_582);
nand U14899 (N_14899,N_7367,N_1312);
nand U14900 (N_14900,N_3723,N_2643);
and U14901 (N_14901,N_2878,N_2312);
nand U14902 (N_14902,N_8386,N_4773);
and U14903 (N_14903,N_4635,N_1654);
or U14904 (N_14904,N_9006,N_8413);
or U14905 (N_14905,N_8002,N_5148);
nor U14906 (N_14906,N_2481,N_1258);
or U14907 (N_14907,N_3794,N_1623);
nor U14908 (N_14908,N_6716,N_7510);
or U14909 (N_14909,N_8770,N_8721);
or U14910 (N_14910,N_5168,N_5429);
or U14911 (N_14911,N_6492,N_758);
and U14912 (N_14912,N_2632,N_506);
or U14913 (N_14913,N_7618,N_3493);
nor U14914 (N_14914,N_2335,N_1616);
or U14915 (N_14915,N_8158,N_8299);
and U14916 (N_14916,N_3515,N_577);
nand U14917 (N_14917,N_4349,N_8297);
nand U14918 (N_14918,N_7629,N_4354);
and U14919 (N_14919,N_2231,N_2132);
or U14920 (N_14920,N_5892,N_4076);
and U14921 (N_14921,N_9233,N_9507);
nor U14922 (N_14922,N_7076,N_1034);
nor U14923 (N_14923,N_7319,N_3302);
xor U14924 (N_14924,N_8141,N_237);
and U14925 (N_14925,N_8493,N_3040);
nor U14926 (N_14926,N_5852,N_4511);
and U14927 (N_14927,N_1397,N_523);
xnor U14928 (N_14928,N_5646,N_7096);
or U14929 (N_14929,N_4445,N_389);
nand U14930 (N_14930,N_1416,N_8967);
nand U14931 (N_14931,N_8068,N_7893);
nand U14932 (N_14932,N_6580,N_7262);
nor U14933 (N_14933,N_7785,N_6419);
xnor U14934 (N_14934,N_3288,N_9761);
nor U14935 (N_14935,N_9237,N_2212);
nand U14936 (N_14936,N_1241,N_3678);
nor U14937 (N_14937,N_8759,N_5627);
nand U14938 (N_14938,N_3186,N_1819);
xnor U14939 (N_14939,N_298,N_846);
nand U14940 (N_14940,N_8801,N_6155);
and U14941 (N_14941,N_9635,N_4698);
nor U14942 (N_14942,N_292,N_3839);
and U14943 (N_14943,N_2622,N_7684);
xnor U14944 (N_14944,N_82,N_3808);
nor U14945 (N_14945,N_6202,N_8166);
and U14946 (N_14946,N_3823,N_8735);
or U14947 (N_14947,N_7187,N_2394);
and U14948 (N_14948,N_5942,N_2436);
and U14949 (N_14949,N_8461,N_221);
or U14950 (N_14950,N_6218,N_8811);
xnor U14951 (N_14951,N_8063,N_8957);
nand U14952 (N_14952,N_1229,N_1764);
or U14953 (N_14953,N_7456,N_8049);
or U14954 (N_14954,N_1648,N_2758);
and U14955 (N_14955,N_6974,N_2604);
nor U14956 (N_14956,N_6031,N_9870);
nand U14957 (N_14957,N_8640,N_3259);
and U14958 (N_14958,N_664,N_6221);
xor U14959 (N_14959,N_8662,N_9625);
xor U14960 (N_14960,N_4518,N_5671);
nand U14961 (N_14961,N_5356,N_6198);
or U14962 (N_14962,N_8045,N_7835);
and U14963 (N_14963,N_7859,N_5025);
or U14964 (N_14964,N_5056,N_8644);
nor U14965 (N_14965,N_6686,N_2334);
nor U14966 (N_14966,N_6807,N_3306);
and U14967 (N_14967,N_6461,N_4938);
and U14968 (N_14968,N_9275,N_7102);
nor U14969 (N_14969,N_4159,N_1013);
nor U14970 (N_14970,N_9592,N_9437);
or U14971 (N_14971,N_8388,N_7536);
nand U14972 (N_14972,N_4816,N_7128);
nand U14973 (N_14973,N_195,N_2510);
nand U14974 (N_14974,N_4295,N_1123);
nand U14975 (N_14975,N_9455,N_3364);
or U14976 (N_14976,N_940,N_3615);
xor U14977 (N_14977,N_3265,N_5298);
and U14978 (N_14978,N_4217,N_6349);
nand U14979 (N_14979,N_2059,N_4439);
nor U14980 (N_14980,N_1287,N_3579);
and U14981 (N_14981,N_3219,N_947);
nand U14982 (N_14982,N_3551,N_6323);
and U14983 (N_14983,N_9321,N_8775);
xnor U14984 (N_14984,N_6024,N_6946);
and U14985 (N_14985,N_7976,N_1808);
or U14986 (N_14986,N_3554,N_8411);
nor U14987 (N_14987,N_9113,N_3160);
nand U14988 (N_14988,N_4964,N_4975);
or U14989 (N_14989,N_7137,N_547);
xnor U14990 (N_14990,N_3614,N_2931);
and U14991 (N_14991,N_9940,N_9270);
nor U14992 (N_14992,N_1837,N_377);
nand U14993 (N_14993,N_7970,N_7903);
or U14994 (N_14994,N_6315,N_8470);
and U14995 (N_14995,N_2716,N_5299);
or U14996 (N_14996,N_1902,N_9910);
nor U14997 (N_14997,N_8261,N_1789);
and U14998 (N_14998,N_4466,N_7414);
xnor U14999 (N_14999,N_9725,N_2852);
and U15000 (N_15000,N_2230,N_8962);
xnor U15001 (N_15001,N_9236,N_3052);
nor U15002 (N_15002,N_3882,N_4703);
or U15003 (N_15003,N_9124,N_294);
or U15004 (N_15004,N_2722,N_341);
and U15005 (N_15005,N_6167,N_7190);
or U15006 (N_15006,N_2401,N_9950);
nand U15007 (N_15007,N_6734,N_7003);
or U15008 (N_15008,N_1767,N_1139);
nand U15009 (N_15009,N_2158,N_8468);
nand U15010 (N_15010,N_4679,N_7338);
or U15011 (N_15011,N_4315,N_555);
xnor U15012 (N_15012,N_5698,N_2726);
nor U15013 (N_15013,N_6878,N_7886);
xnor U15014 (N_15014,N_2612,N_6426);
nor U15015 (N_15015,N_7373,N_8989);
and U15016 (N_15016,N_2773,N_6819);
xnor U15017 (N_15017,N_6352,N_7818);
nor U15018 (N_15018,N_4636,N_3387);
nor U15019 (N_15019,N_6290,N_6127);
nand U15020 (N_15020,N_2524,N_6159);
nor U15021 (N_15021,N_2282,N_8254);
nor U15022 (N_15022,N_5291,N_1109);
xnor U15023 (N_15023,N_8313,N_3720);
xor U15024 (N_15024,N_4773,N_2711);
nand U15025 (N_15025,N_1383,N_8031);
nand U15026 (N_15026,N_6217,N_8022);
and U15027 (N_15027,N_5992,N_1362);
nor U15028 (N_15028,N_6101,N_3668);
nor U15029 (N_15029,N_4092,N_6439);
nor U15030 (N_15030,N_2628,N_2081);
nand U15031 (N_15031,N_1447,N_8194);
xor U15032 (N_15032,N_1194,N_3414);
and U15033 (N_15033,N_6790,N_3671);
nor U15034 (N_15034,N_7694,N_2089);
nand U15035 (N_15035,N_6511,N_6662);
or U15036 (N_15036,N_1808,N_410);
or U15037 (N_15037,N_3852,N_7290);
or U15038 (N_15038,N_4772,N_2779);
or U15039 (N_15039,N_8862,N_3877);
and U15040 (N_15040,N_2707,N_7092);
nor U15041 (N_15041,N_7895,N_7447);
and U15042 (N_15042,N_4641,N_3709);
xor U15043 (N_15043,N_3754,N_6556);
nor U15044 (N_15044,N_3568,N_7484);
or U15045 (N_15045,N_5283,N_7987);
or U15046 (N_15046,N_9249,N_7453);
and U15047 (N_15047,N_4487,N_8779);
or U15048 (N_15048,N_8433,N_2597);
nand U15049 (N_15049,N_4691,N_7728);
nand U15050 (N_15050,N_3525,N_7854);
nor U15051 (N_15051,N_2160,N_6591);
nor U15052 (N_15052,N_1552,N_6295);
nand U15053 (N_15053,N_6498,N_9723);
or U15054 (N_15054,N_9366,N_8526);
and U15055 (N_15055,N_1927,N_9297);
and U15056 (N_15056,N_8351,N_872);
and U15057 (N_15057,N_3469,N_9802);
and U15058 (N_15058,N_1864,N_1300);
xor U15059 (N_15059,N_1981,N_5087);
nor U15060 (N_15060,N_5627,N_3230);
nand U15061 (N_15061,N_8672,N_8951);
and U15062 (N_15062,N_2022,N_6147);
and U15063 (N_15063,N_7624,N_4259);
nand U15064 (N_15064,N_969,N_2631);
and U15065 (N_15065,N_9525,N_8801);
and U15066 (N_15066,N_9765,N_7237);
nor U15067 (N_15067,N_8157,N_7534);
and U15068 (N_15068,N_4333,N_8555);
and U15069 (N_15069,N_6314,N_9797);
nor U15070 (N_15070,N_8497,N_174);
and U15071 (N_15071,N_3945,N_4804);
nor U15072 (N_15072,N_2075,N_5644);
nand U15073 (N_15073,N_9520,N_4849);
nand U15074 (N_15074,N_1070,N_3017);
nand U15075 (N_15075,N_8528,N_1097);
nand U15076 (N_15076,N_3022,N_6114);
nor U15077 (N_15077,N_2772,N_7944);
and U15078 (N_15078,N_559,N_6996);
or U15079 (N_15079,N_5616,N_582);
nor U15080 (N_15080,N_4463,N_3131);
or U15081 (N_15081,N_9717,N_519);
nand U15082 (N_15082,N_6663,N_8959);
and U15083 (N_15083,N_5238,N_6149);
nor U15084 (N_15084,N_8431,N_5747);
nand U15085 (N_15085,N_6125,N_5295);
nor U15086 (N_15086,N_8087,N_3556);
nor U15087 (N_15087,N_1285,N_1877);
nor U15088 (N_15088,N_9565,N_7254);
nor U15089 (N_15089,N_2010,N_7743);
or U15090 (N_15090,N_3608,N_8168);
nor U15091 (N_15091,N_4655,N_508);
nand U15092 (N_15092,N_4335,N_6694);
xor U15093 (N_15093,N_3206,N_3958);
and U15094 (N_15094,N_8215,N_3056);
nor U15095 (N_15095,N_3701,N_1771);
xor U15096 (N_15096,N_349,N_9935);
and U15097 (N_15097,N_1854,N_1127);
nand U15098 (N_15098,N_9499,N_8695);
nand U15099 (N_15099,N_2021,N_7705);
and U15100 (N_15100,N_1707,N_1924);
nand U15101 (N_15101,N_4885,N_9976);
or U15102 (N_15102,N_3464,N_8001);
and U15103 (N_15103,N_6619,N_5252);
and U15104 (N_15104,N_8980,N_9198);
or U15105 (N_15105,N_6489,N_7067);
and U15106 (N_15106,N_5370,N_1927);
nand U15107 (N_15107,N_1116,N_1780);
or U15108 (N_15108,N_6704,N_895);
or U15109 (N_15109,N_3996,N_2132);
nor U15110 (N_15110,N_9102,N_3684);
and U15111 (N_15111,N_5663,N_5091);
xnor U15112 (N_15112,N_2871,N_6618);
or U15113 (N_15113,N_2266,N_9930);
nor U15114 (N_15114,N_2008,N_1223);
or U15115 (N_15115,N_9496,N_894);
nor U15116 (N_15116,N_6609,N_6205);
nor U15117 (N_15117,N_8579,N_1212);
or U15118 (N_15118,N_8974,N_6374);
nand U15119 (N_15119,N_2281,N_3643);
nor U15120 (N_15120,N_6307,N_4835);
nand U15121 (N_15121,N_1623,N_6249);
nand U15122 (N_15122,N_2579,N_3907);
nand U15123 (N_15123,N_212,N_2256);
nand U15124 (N_15124,N_5645,N_7562);
nor U15125 (N_15125,N_4985,N_7919);
xnor U15126 (N_15126,N_9782,N_579);
nand U15127 (N_15127,N_6278,N_352);
and U15128 (N_15128,N_6591,N_8405);
nand U15129 (N_15129,N_7961,N_3718);
or U15130 (N_15130,N_2423,N_5814);
nor U15131 (N_15131,N_2881,N_2922);
xor U15132 (N_15132,N_2243,N_6511);
nor U15133 (N_15133,N_1364,N_5656);
or U15134 (N_15134,N_9670,N_2169);
xnor U15135 (N_15135,N_9320,N_6838);
nor U15136 (N_15136,N_3171,N_9755);
nor U15137 (N_15137,N_7869,N_2927);
or U15138 (N_15138,N_459,N_7735);
or U15139 (N_15139,N_715,N_8215);
and U15140 (N_15140,N_8290,N_6022);
or U15141 (N_15141,N_8542,N_7856);
nor U15142 (N_15142,N_6089,N_7812);
nand U15143 (N_15143,N_5643,N_4729);
nand U15144 (N_15144,N_2510,N_8310);
or U15145 (N_15145,N_1792,N_3911);
and U15146 (N_15146,N_5310,N_4396);
and U15147 (N_15147,N_8862,N_6639);
nand U15148 (N_15148,N_9547,N_1715);
nand U15149 (N_15149,N_2829,N_9648);
or U15150 (N_15150,N_1242,N_9672);
nand U15151 (N_15151,N_1008,N_8045);
nor U15152 (N_15152,N_8082,N_717);
nor U15153 (N_15153,N_2922,N_5794);
nor U15154 (N_15154,N_9844,N_4421);
nor U15155 (N_15155,N_6008,N_970);
nand U15156 (N_15156,N_1921,N_9849);
xor U15157 (N_15157,N_4031,N_9905);
or U15158 (N_15158,N_1297,N_8363);
or U15159 (N_15159,N_5052,N_6163);
nand U15160 (N_15160,N_6381,N_8626);
or U15161 (N_15161,N_2218,N_5385);
and U15162 (N_15162,N_33,N_3986);
nand U15163 (N_15163,N_7005,N_822);
and U15164 (N_15164,N_850,N_695);
and U15165 (N_15165,N_679,N_1140);
nor U15166 (N_15166,N_759,N_7237);
xor U15167 (N_15167,N_6388,N_8987);
and U15168 (N_15168,N_4252,N_4496);
nand U15169 (N_15169,N_9399,N_4280);
and U15170 (N_15170,N_5140,N_9322);
and U15171 (N_15171,N_4724,N_9585);
nor U15172 (N_15172,N_2245,N_374);
nor U15173 (N_15173,N_3686,N_2754);
xor U15174 (N_15174,N_3568,N_3610);
nor U15175 (N_15175,N_988,N_4301);
or U15176 (N_15176,N_5225,N_8643);
or U15177 (N_15177,N_4991,N_4838);
nor U15178 (N_15178,N_1594,N_3079);
nand U15179 (N_15179,N_5837,N_5660);
or U15180 (N_15180,N_7071,N_157);
nor U15181 (N_15181,N_9036,N_1784);
nand U15182 (N_15182,N_4527,N_4416);
nand U15183 (N_15183,N_6752,N_7258);
nor U15184 (N_15184,N_1492,N_7398);
or U15185 (N_15185,N_4165,N_8460);
nand U15186 (N_15186,N_7438,N_582);
nand U15187 (N_15187,N_3996,N_2150);
and U15188 (N_15188,N_7852,N_3145);
nand U15189 (N_15189,N_9847,N_7659);
nand U15190 (N_15190,N_6220,N_3432);
nand U15191 (N_15191,N_9021,N_6004);
nand U15192 (N_15192,N_2875,N_7350);
xor U15193 (N_15193,N_7822,N_3168);
or U15194 (N_15194,N_6791,N_9856);
and U15195 (N_15195,N_2059,N_1129);
or U15196 (N_15196,N_9007,N_4704);
nand U15197 (N_15197,N_4563,N_2035);
or U15198 (N_15198,N_7471,N_2383);
nand U15199 (N_15199,N_7030,N_6083);
or U15200 (N_15200,N_2587,N_5751);
xor U15201 (N_15201,N_7230,N_8966);
xnor U15202 (N_15202,N_1540,N_3322);
nand U15203 (N_15203,N_9016,N_3847);
nand U15204 (N_15204,N_9945,N_2775);
nand U15205 (N_15205,N_8263,N_5656);
nand U15206 (N_15206,N_5829,N_8620);
nor U15207 (N_15207,N_3387,N_3968);
nor U15208 (N_15208,N_121,N_8442);
nor U15209 (N_15209,N_1438,N_1190);
nand U15210 (N_15210,N_2745,N_3681);
xor U15211 (N_15211,N_5250,N_1593);
nand U15212 (N_15212,N_7349,N_7956);
or U15213 (N_15213,N_2209,N_7438);
or U15214 (N_15214,N_5678,N_716);
or U15215 (N_15215,N_4152,N_3953);
and U15216 (N_15216,N_6947,N_8241);
and U15217 (N_15217,N_4625,N_1310);
nand U15218 (N_15218,N_2742,N_596);
nor U15219 (N_15219,N_6161,N_7632);
nor U15220 (N_15220,N_9129,N_7024);
or U15221 (N_15221,N_6421,N_5859);
xnor U15222 (N_15222,N_6337,N_1117);
xor U15223 (N_15223,N_9834,N_512);
and U15224 (N_15224,N_2353,N_9701);
nand U15225 (N_15225,N_3545,N_1840);
nor U15226 (N_15226,N_215,N_9720);
nand U15227 (N_15227,N_8861,N_307);
or U15228 (N_15228,N_9522,N_9935);
or U15229 (N_15229,N_5079,N_6849);
nor U15230 (N_15230,N_8396,N_8911);
nand U15231 (N_15231,N_1328,N_4871);
xor U15232 (N_15232,N_2530,N_4000);
or U15233 (N_15233,N_3722,N_2005);
and U15234 (N_15234,N_441,N_9788);
nor U15235 (N_15235,N_1498,N_8928);
nand U15236 (N_15236,N_6351,N_5439);
or U15237 (N_15237,N_2589,N_1071);
and U15238 (N_15238,N_8907,N_8756);
nand U15239 (N_15239,N_4354,N_8570);
and U15240 (N_15240,N_107,N_9040);
nor U15241 (N_15241,N_31,N_3519);
or U15242 (N_15242,N_9632,N_9771);
or U15243 (N_15243,N_3410,N_4239);
nand U15244 (N_15244,N_6383,N_7154);
or U15245 (N_15245,N_4766,N_252);
nand U15246 (N_15246,N_2080,N_6714);
nor U15247 (N_15247,N_5513,N_5250);
and U15248 (N_15248,N_6479,N_9775);
and U15249 (N_15249,N_4520,N_9500);
nand U15250 (N_15250,N_8173,N_2865);
nor U15251 (N_15251,N_8640,N_1521);
and U15252 (N_15252,N_459,N_9242);
nand U15253 (N_15253,N_1074,N_1800);
nand U15254 (N_15254,N_3159,N_6163);
nand U15255 (N_15255,N_233,N_1881);
or U15256 (N_15256,N_3218,N_4123);
nor U15257 (N_15257,N_5826,N_5526);
xnor U15258 (N_15258,N_5405,N_6102);
and U15259 (N_15259,N_6917,N_7786);
xnor U15260 (N_15260,N_363,N_5837);
and U15261 (N_15261,N_9015,N_856);
xnor U15262 (N_15262,N_3736,N_6974);
or U15263 (N_15263,N_6630,N_3517);
xnor U15264 (N_15264,N_9788,N_9909);
nand U15265 (N_15265,N_9048,N_832);
and U15266 (N_15266,N_8170,N_8634);
nor U15267 (N_15267,N_3573,N_6440);
and U15268 (N_15268,N_7521,N_9172);
and U15269 (N_15269,N_9736,N_654);
or U15270 (N_15270,N_1563,N_3084);
nor U15271 (N_15271,N_907,N_5514);
and U15272 (N_15272,N_1768,N_3970);
and U15273 (N_15273,N_7302,N_6569);
or U15274 (N_15274,N_6691,N_2008);
xor U15275 (N_15275,N_8253,N_6155);
and U15276 (N_15276,N_3011,N_6900);
or U15277 (N_15277,N_1159,N_8283);
and U15278 (N_15278,N_1356,N_7421);
nand U15279 (N_15279,N_3732,N_2193);
nand U15280 (N_15280,N_3937,N_981);
nor U15281 (N_15281,N_3294,N_8715);
and U15282 (N_15282,N_5240,N_2774);
and U15283 (N_15283,N_1234,N_9124);
nor U15284 (N_15284,N_2695,N_1390);
and U15285 (N_15285,N_3738,N_6268);
xor U15286 (N_15286,N_8114,N_9364);
nor U15287 (N_15287,N_5620,N_6523);
nor U15288 (N_15288,N_8201,N_5350);
or U15289 (N_15289,N_3776,N_1795);
nand U15290 (N_15290,N_6306,N_9412);
nor U15291 (N_15291,N_3979,N_4674);
xor U15292 (N_15292,N_9103,N_6325);
nor U15293 (N_15293,N_9398,N_1422);
nand U15294 (N_15294,N_993,N_7509);
nor U15295 (N_15295,N_2086,N_7258);
xnor U15296 (N_15296,N_7537,N_3653);
or U15297 (N_15297,N_7307,N_2662);
and U15298 (N_15298,N_4286,N_9484);
nor U15299 (N_15299,N_6386,N_4651);
or U15300 (N_15300,N_9785,N_7641);
nor U15301 (N_15301,N_9371,N_7973);
nor U15302 (N_15302,N_2256,N_8437);
nand U15303 (N_15303,N_6882,N_9903);
xnor U15304 (N_15304,N_2689,N_6509);
xnor U15305 (N_15305,N_6751,N_2680);
or U15306 (N_15306,N_2324,N_9494);
nor U15307 (N_15307,N_9380,N_4678);
and U15308 (N_15308,N_552,N_3441);
nor U15309 (N_15309,N_6525,N_4371);
xor U15310 (N_15310,N_6267,N_4132);
or U15311 (N_15311,N_9559,N_883);
or U15312 (N_15312,N_8961,N_5571);
or U15313 (N_15313,N_8253,N_9797);
nor U15314 (N_15314,N_5433,N_2985);
nand U15315 (N_15315,N_1432,N_2976);
xor U15316 (N_15316,N_5899,N_5931);
nand U15317 (N_15317,N_5231,N_2198);
and U15318 (N_15318,N_302,N_3584);
nand U15319 (N_15319,N_1010,N_3750);
and U15320 (N_15320,N_2582,N_3986);
or U15321 (N_15321,N_1283,N_678);
nand U15322 (N_15322,N_3966,N_8258);
xor U15323 (N_15323,N_9039,N_2465);
nor U15324 (N_15324,N_271,N_5396);
and U15325 (N_15325,N_4831,N_8638);
and U15326 (N_15326,N_2861,N_6615);
nor U15327 (N_15327,N_3637,N_5806);
nand U15328 (N_15328,N_5297,N_6068);
or U15329 (N_15329,N_3664,N_4978);
nor U15330 (N_15330,N_6272,N_4855);
nand U15331 (N_15331,N_1333,N_3143);
nand U15332 (N_15332,N_9893,N_5813);
and U15333 (N_15333,N_7415,N_4478);
nand U15334 (N_15334,N_5416,N_8995);
or U15335 (N_15335,N_3881,N_7775);
xor U15336 (N_15336,N_3253,N_7057);
and U15337 (N_15337,N_1214,N_556);
or U15338 (N_15338,N_6645,N_1709);
and U15339 (N_15339,N_6576,N_3769);
xor U15340 (N_15340,N_4818,N_8075);
xor U15341 (N_15341,N_7021,N_5379);
nand U15342 (N_15342,N_7138,N_3821);
or U15343 (N_15343,N_6853,N_3477);
nand U15344 (N_15344,N_3030,N_5930);
nand U15345 (N_15345,N_3200,N_9227);
and U15346 (N_15346,N_8417,N_4415);
or U15347 (N_15347,N_6249,N_8867);
nor U15348 (N_15348,N_1964,N_5655);
nor U15349 (N_15349,N_1303,N_1384);
and U15350 (N_15350,N_233,N_5112);
nand U15351 (N_15351,N_1305,N_1044);
or U15352 (N_15352,N_9666,N_1363);
xnor U15353 (N_15353,N_1668,N_6584);
nor U15354 (N_15354,N_9475,N_2694);
nand U15355 (N_15355,N_5111,N_4947);
nand U15356 (N_15356,N_1295,N_9387);
nand U15357 (N_15357,N_6616,N_9980);
nand U15358 (N_15358,N_6878,N_375);
and U15359 (N_15359,N_817,N_3794);
nor U15360 (N_15360,N_2064,N_8179);
nand U15361 (N_15361,N_1344,N_7590);
and U15362 (N_15362,N_7157,N_2963);
nand U15363 (N_15363,N_5881,N_5626);
nand U15364 (N_15364,N_5547,N_6894);
xnor U15365 (N_15365,N_4679,N_1308);
xor U15366 (N_15366,N_6224,N_9762);
and U15367 (N_15367,N_170,N_8103);
nor U15368 (N_15368,N_4603,N_4239);
and U15369 (N_15369,N_5818,N_7170);
xor U15370 (N_15370,N_2001,N_4426);
nor U15371 (N_15371,N_1234,N_3947);
and U15372 (N_15372,N_8868,N_8972);
or U15373 (N_15373,N_5375,N_9582);
nand U15374 (N_15374,N_3210,N_250);
and U15375 (N_15375,N_6541,N_7403);
nand U15376 (N_15376,N_4517,N_688);
or U15377 (N_15377,N_4265,N_6099);
nor U15378 (N_15378,N_3514,N_4930);
and U15379 (N_15379,N_2257,N_1312);
and U15380 (N_15380,N_8614,N_6990);
nand U15381 (N_15381,N_6006,N_535);
nor U15382 (N_15382,N_9173,N_4620);
nor U15383 (N_15383,N_7548,N_4267);
nor U15384 (N_15384,N_1318,N_9783);
xor U15385 (N_15385,N_4334,N_628);
and U15386 (N_15386,N_4340,N_6833);
nand U15387 (N_15387,N_8837,N_8498);
and U15388 (N_15388,N_4739,N_4281);
and U15389 (N_15389,N_3272,N_4386);
or U15390 (N_15390,N_6817,N_6672);
nor U15391 (N_15391,N_9362,N_5564);
and U15392 (N_15392,N_1131,N_4080);
or U15393 (N_15393,N_7970,N_972);
and U15394 (N_15394,N_2187,N_8718);
or U15395 (N_15395,N_5483,N_8456);
nor U15396 (N_15396,N_3853,N_4669);
and U15397 (N_15397,N_5001,N_5671);
or U15398 (N_15398,N_5301,N_657);
nand U15399 (N_15399,N_5069,N_6555);
nor U15400 (N_15400,N_391,N_8640);
nand U15401 (N_15401,N_4314,N_4249);
or U15402 (N_15402,N_535,N_3692);
nor U15403 (N_15403,N_7946,N_458);
nor U15404 (N_15404,N_777,N_2078);
nand U15405 (N_15405,N_3884,N_715);
and U15406 (N_15406,N_6512,N_3091);
nand U15407 (N_15407,N_8048,N_7381);
and U15408 (N_15408,N_307,N_7497);
and U15409 (N_15409,N_1258,N_3499);
or U15410 (N_15410,N_522,N_4179);
and U15411 (N_15411,N_2549,N_3560);
nor U15412 (N_15412,N_6473,N_9017);
or U15413 (N_15413,N_6249,N_5188);
nor U15414 (N_15414,N_7253,N_8204);
or U15415 (N_15415,N_3165,N_1935);
xor U15416 (N_15416,N_206,N_880);
nand U15417 (N_15417,N_3843,N_7068);
xnor U15418 (N_15418,N_9641,N_4969);
nand U15419 (N_15419,N_748,N_2653);
nand U15420 (N_15420,N_8085,N_3318);
nor U15421 (N_15421,N_658,N_2134);
and U15422 (N_15422,N_4621,N_2056);
or U15423 (N_15423,N_3452,N_2974);
nand U15424 (N_15424,N_1160,N_7196);
nand U15425 (N_15425,N_2451,N_533);
nand U15426 (N_15426,N_4221,N_943);
nand U15427 (N_15427,N_2116,N_8004);
or U15428 (N_15428,N_4880,N_7294);
or U15429 (N_15429,N_6614,N_3241);
xnor U15430 (N_15430,N_7893,N_3958);
or U15431 (N_15431,N_1020,N_1018);
and U15432 (N_15432,N_4601,N_6398);
or U15433 (N_15433,N_4064,N_7147);
nand U15434 (N_15434,N_8933,N_3512);
or U15435 (N_15435,N_1350,N_1623);
nand U15436 (N_15436,N_1200,N_8701);
xor U15437 (N_15437,N_6649,N_7840);
nor U15438 (N_15438,N_6541,N_7802);
nand U15439 (N_15439,N_1556,N_7429);
nor U15440 (N_15440,N_3709,N_5508);
and U15441 (N_15441,N_5206,N_5229);
xor U15442 (N_15442,N_617,N_3788);
nor U15443 (N_15443,N_8233,N_1983);
nand U15444 (N_15444,N_8945,N_8992);
nand U15445 (N_15445,N_2034,N_510);
xnor U15446 (N_15446,N_7410,N_617);
and U15447 (N_15447,N_5837,N_1086);
nand U15448 (N_15448,N_6483,N_4284);
and U15449 (N_15449,N_1718,N_4885);
and U15450 (N_15450,N_7287,N_639);
nand U15451 (N_15451,N_9672,N_1358);
and U15452 (N_15452,N_6385,N_3080);
or U15453 (N_15453,N_5176,N_6364);
xor U15454 (N_15454,N_5001,N_9517);
nand U15455 (N_15455,N_3202,N_2517);
nor U15456 (N_15456,N_2084,N_8845);
nand U15457 (N_15457,N_8839,N_9262);
nand U15458 (N_15458,N_93,N_7475);
nor U15459 (N_15459,N_8206,N_7110);
xor U15460 (N_15460,N_9708,N_9173);
and U15461 (N_15461,N_9036,N_1814);
or U15462 (N_15462,N_8677,N_2195);
xnor U15463 (N_15463,N_1731,N_1941);
nor U15464 (N_15464,N_4156,N_2231);
nand U15465 (N_15465,N_2299,N_2260);
or U15466 (N_15466,N_9421,N_6515);
nand U15467 (N_15467,N_1103,N_9469);
nor U15468 (N_15468,N_2460,N_2474);
nor U15469 (N_15469,N_8016,N_3240);
or U15470 (N_15470,N_7818,N_1235);
nor U15471 (N_15471,N_5774,N_9033);
or U15472 (N_15472,N_4925,N_5958);
and U15473 (N_15473,N_2691,N_6994);
and U15474 (N_15474,N_1517,N_8416);
nor U15475 (N_15475,N_8576,N_7534);
and U15476 (N_15476,N_7775,N_1805);
and U15477 (N_15477,N_6804,N_9948);
nor U15478 (N_15478,N_3446,N_9389);
and U15479 (N_15479,N_8876,N_572);
and U15480 (N_15480,N_3532,N_3780);
nand U15481 (N_15481,N_6001,N_9082);
or U15482 (N_15482,N_2091,N_4620);
or U15483 (N_15483,N_5225,N_4896);
xnor U15484 (N_15484,N_2277,N_1486);
or U15485 (N_15485,N_558,N_4009);
nand U15486 (N_15486,N_568,N_600);
and U15487 (N_15487,N_4767,N_8702);
or U15488 (N_15488,N_3854,N_7337);
nand U15489 (N_15489,N_6935,N_227);
nand U15490 (N_15490,N_1386,N_6694);
nor U15491 (N_15491,N_9613,N_721);
and U15492 (N_15492,N_6199,N_6737);
nand U15493 (N_15493,N_6296,N_5176);
nor U15494 (N_15494,N_4901,N_49);
nor U15495 (N_15495,N_7060,N_9757);
or U15496 (N_15496,N_1803,N_8523);
nor U15497 (N_15497,N_738,N_1812);
and U15498 (N_15498,N_6251,N_5508);
nand U15499 (N_15499,N_6219,N_3164);
or U15500 (N_15500,N_7844,N_5040);
nor U15501 (N_15501,N_3092,N_8291);
or U15502 (N_15502,N_4458,N_6003);
nor U15503 (N_15503,N_4468,N_3950);
and U15504 (N_15504,N_468,N_6933);
or U15505 (N_15505,N_5161,N_6478);
nor U15506 (N_15506,N_9815,N_1491);
nor U15507 (N_15507,N_361,N_6875);
and U15508 (N_15508,N_7366,N_8227);
nand U15509 (N_15509,N_7487,N_7157);
and U15510 (N_15510,N_9431,N_3634);
nor U15511 (N_15511,N_7784,N_1216);
or U15512 (N_15512,N_5376,N_5037);
nand U15513 (N_15513,N_2038,N_8991);
nand U15514 (N_15514,N_9465,N_7141);
or U15515 (N_15515,N_6895,N_1060);
nand U15516 (N_15516,N_1147,N_5837);
xor U15517 (N_15517,N_1181,N_7501);
xnor U15518 (N_15518,N_1041,N_6903);
nor U15519 (N_15519,N_9684,N_356);
nor U15520 (N_15520,N_9403,N_4823);
or U15521 (N_15521,N_9328,N_3395);
and U15522 (N_15522,N_1612,N_4);
or U15523 (N_15523,N_6777,N_3514);
or U15524 (N_15524,N_8580,N_3876);
or U15525 (N_15525,N_7780,N_634);
and U15526 (N_15526,N_2336,N_5765);
or U15527 (N_15527,N_6019,N_8021);
and U15528 (N_15528,N_2766,N_4421);
nand U15529 (N_15529,N_6025,N_5345);
and U15530 (N_15530,N_1213,N_8990);
nor U15531 (N_15531,N_6887,N_3050);
and U15532 (N_15532,N_672,N_9131);
or U15533 (N_15533,N_8326,N_3142);
and U15534 (N_15534,N_2127,N_8989);
xor U15535 (N_15535,N_5000,N_3649);
and U15536 (N_15536,N_8555,N_4432);
or U15537 (N_15537,N_3523,N_8136);
and U15538 (N_15538,N_5047,N_6943);
nor U15539 (N_15539,N_6573,N_343);
xnor U15540 (N_15540,N_8505,N_6289);
nand U15541 (N_15541,N_2593,N_4806);
nand U15542 (N_15542,N_5717,N_8556);
or U15543 (N_15543,N_2647,N_7036);
xnor U15544 (N_15544,N_9822,N_8845);
nor U15545 (N_15545,N_8808,N_1515);
or U15546 (N_15546,N_1380,N_739);
or U15547 (N_15547,N_9198,N_6712);
nand U15548 (N_15548,N_621,N_8584);
and U15549 (N_15549,N_7273,N_6237);
nor U15550 (N_15550,N_5200,N_6603);
or U15551 (N_15551,N_6058,N_6952);
nor U15552 (N_15552,N_4544,N_1341);
nand U15553 (N_15553,N_3103,N_3687);
or U15554 (N_15554,N_4294,N_6692);
xnor U15555 (N_15555,N_8601,N_4026);
nand U15556 (N_15556,N_7807,N_8137);
nand U15557 (N_15557,N_9765,N_1803);
nor U15558 (N_15558,N_6137,N_1235);
nand U15559 (N_15559,N_9076,N_8628);
and U15560 (N_15560,N_244,N_836);
nand U15561 (N_15561,N_933,N_8158);
nor U15562 (N_15562,N_7956,N_6682);
or U15563 (N_15563,N_4312,N_6245);
and U15564 (N_15564,N_5160,N_3920);
or U15565 (N_15565,N_7146,N_8295);
or U15566 (N_15566,N_3423,N_6057);
or U15567 (N_15567,N_4317,N_273);
and U15568 (N_15568,N_4902,N_5629);
and U15569 (N_15569,N_2548,N_463);
and U15570 (N_15570,N_6527,N_2524);
nand U15571 (N_15571,N_9804,N_2158);
or U15572 (N_15572,N_917,N_2453);
nand U15573 (N_15573,N_980,N_6182);
and U15574 (N_15574,N_1287,N_9498);
xor U15575 (N_15575,N_6165,N_6979);
xnor U15576 (N_15576,N_6813,N_8442);
and U15577 (N_15577,N_305,N_7053);
xnor U15578 (N_15578,N_2332,N_5516);
nor U15579 (N_15579,N_7649,N_6163);
nand U15580 (N_15580,N_4882,N_560);
or U15581 (N_15581,N_7215,N_5159);
nand U15582 (N_15582,N_448,N_3525);
nand U15583 (N_15583,N_3691,N_7564);
or U15584 (N_15584,N_1323,N_8739);
xnor U15585 (N_15585,N_3792,N_6526);
nor U15586 (N_15586,N_210,N_2895);
or U15587 (N_15587,N_5455,N_9021);
and U15588 (N_15588,N_9187,N_4931);
and U15589 (N_15589,N_1414,N_5696);
nand U15590 (N_15590,N_8256,N_8720);
nand U15591 (N_15591,N_4611,N_2471);
nand U15592 (N_15592,N_2970,N_8029);
xor U15593 (N_15593,N_2306,N_9343);
nand U15594 (N_15594,N_2362,N_4534);
and U15595 (N_15595,N_1726,N_2421);
or U15596 (N_15596,N_868,N_8700);
or U15597 (N_15597,N_9858,N_6657);
or U15598 (N_15598,N_4495,N_2834);
nand U15599 (N_15599,N_6537,N_7763);
and U15600 (N_15600,N_1402,N_3069);
nand U15601 (N_15601,N_8026,N_2276);
and U15602 (N_15602,N_891,N_3859);
xor U15603 (N_15603,N_5251,N_6916);
nand U15604 (N_15604,N_1345,N_5000);
xnor U15605 (N_15605,N_4335,N_2711);
nand U15606 (N_15606,N_3219,N_7503);
nor U15607 (N_15607,N_5953,N_4721);
and U15608 (N_15608,N_3704,N_2278);
and U15609 (N_15609,N_3063,N_7967);
nor U15610 (N_15610,N_7403,N_9962);
and U15611 (N_15611,N_4909,N_3727);
nand U15612 (N_15612,N_7801,N_8958);
or U15613 (N_15613,N_9405,N_8915);
and U15614 (N_15614,N_8691,N_5698);
and U15615 (N_15615,N_6818,N_827);
xnor U15616 (N_15616,N_4684,N_8841);
and U15617 (N_15617,N_9919,N_8529);
and U15618 (N_15618,N_5380,N_5534);
nor U15619 (N_15619,N_1038,N_9942);
or U15620 (N_15620,N_4517,N_3055);
nand U15621 (N_15621,N_6841,N_178);
and U15622 (N_15622,N_4540,N_1644);
nor U15623 (N_15623,N_8624,N_2973);
nand U15624 (N_15624,N_2547,N_9886);
nand U15625 (N_15625,N_3232,N_6627);
xnor U15626 (N_15626,N_2778,N_8642);
and U15627 (N_15627,N_5507,N_2720);
or U15628 (N_15628,N_8417,N_9848);
and U15629 (N_15629,N_6781,N_9651);
nand U15630 (N_15630,N_4227,N_6117);
nor U15631 (N_15631,N_5977,N_2350);
nand U15632 (N_15632,N_9678,N_4127);
nand U15633 (N_15633,N_7380,N_7859);
nand U15634 (N_15634,N_4334,N_6802);
nand U15635 (N_15635,N_6816,N_3121);
nor U15636 (N_15636,N_4771,N_4788);
xor U15637 (N_15637,N_9935,N_9878);
and U15638 (N_15638,N_1790,N_1411);
or U15639 (N_15639,N_2227,N_5622);
nor U15640 (N_15640,N_5611,N_4832);
xor U15641 (N_15641,N_9834,N_7123);
nand U15642 (N_15642,N_6494,N_6799);
and U15643 (N_15643,N_1998,N_8737);
xor U15644 (N_15644,N_748,N_1558);
xnor U15645 (N_15645,N_1866,N_6492);
or U15646 (N_15646,N_1096,N_150);
nor U15647 (N_15647,N_4307,N_6006);
or U15648 (N_15648,N_7446,N_1523);
nand U15649 (N_15649,N_2833,N_6338);
xor U15650 (N_15650,N_5618,N_5957);
xor U15651 (N_15651,N_6597,N_9453);
or U15652 (N_15652,N_5570,N_8093);
nand U15653 (N_15653,N_2232,N_9623);
and U15654 (N_15654,N_4037,N_2175);
nand U15655 (N_15655,N_4397,N_9632);
nand U15656 (N_15656,N_7587,N_3301);
and U15657 (N_15657,N_366,N_5031);
nand U15658 (N_15658,N_8724,N_6917);
and U15659 (N_15659,N_8261,N_8276);
nor U15660 (N_15660,N_8168,N_3357);
nand U15661 (N_15661,N_6593,N_2218);
nand U15662 (N_15662,N_6105,N_9786);
xor U15663 (N_15663,N_2452,N_9041);
and U15664 (N_15664,N_5288,N_606);
or U15665 (N_15665,N_6667,N_1378);
and U15666 (N_15666,N_5323,N_6200);
or U15667 (N_15667,N_5246,N_5735);
nand U15668 (N_15668,N_9913,N_8117);
and U15669 (N_15669,N_2633,N_3431);
or U15670 (N_15670,N_7790,N_3694);
xnor U15671 (N_15671,N_4998,N_7611);
nor U15672 (N_15672,N_7797,N_5329);
xnor U15673 (N_15673,N_1059,N_3191);
or U15674 (N_15674,N_5909,N_4105);
nor U15675 (N_15675,N_6120,N_8217);
or U15676 (N_15676,N_5441,N_7642);
and U15677 (N_15677,N_1497,N_6845);
or U15678 (N_15678,N_9424,N_4249);
and U15679 (N_15679,N_5742,N_4491);
nor U15680 (N_15680,N_9260,N_337);
nor U15681 (N_15681,N_2309,N_7685);
or U15682 (N_15682,N_383,N_5081);
nor U15683 (N_15683,N_6530,N_5679);
and U15684 (N_15684,N_1790,N_859);
or U15685 (N_15685,N_5475,N_1671);
nand U15686 (N_15686,N_585,N_8062);
and U15687 (N_15687,N_792,N_4070);
nand U15688 (N_15688,N_846,N_261);
nand U15689 (N_15689,N_99,N_3231);
and U15690 (N_15690,N_3020,N_5570);
or U15691 (N_15691,N_11,N_1860);
and U15692 (N_15692,N_8431,N_5052);
and U15693 (N_15693,N_9800,N_9445);
xnor U15694 (N_15694,N_7733,N_7928);
nand U15695 (N_15695,N_7997,N_6110);
nand U15696 (N_15696,N_7243,N_2464);
or U15697 (N_15697,N_3989,N_5229);
nand U15698 (N_15698,N_8842,N_6667);
nor U15699 (N_15699,N_7817,N_9898);
nor U15700 (N_15700,N_6133,N_3549);
nor U15701 (N_15701,N_7415,N_3697);
nor U15702 (N_15702,N_9590,N_3306);
nand U15703 (N_15703,N_66,N_9839);
nor U15704 (N_15704,N_3299,N_8429);
and U15705 (N_15705,N_7902,N_758);
nor U15706 (N_15706,N_165,N_6769);
nand U15707 (N_15707,N_7052,N_7492);
nor U15708 (N_15708,N_4071,N_3359);
and U15709 (N_15709,N_4213,N_794);
xnor U15710 (N_15710,N_5056,N_3101);
and U15711 (N_15711,N_3945,N_9931);
xor U15712 (N_15712,N_2058,N_6519);
or U15713 (N_15713,N_5970,N_9376);
and U15714 (N_15714,N_1786,N_5349);
nand U15715 (N_15715,N_7995,N_5372);
and U15716 (N_15716,N_9376,N_2456);
nand U15717 (N_15717,N_8898,N_7671);
nand U15718 (N_15718,N_4863,N_3567);
nor U15719 (N_15719,N_5848,N_7888);
xor U15720 (N_15720,N_8219,N_365);
nand U15721 (N_15721,N_6499,N_1864);
nand U15722 (N_15722,N_306,N_9868);
and U15723 (N_15723,N_5409,N_6260);
xor U15724 (N_15724,N_8017,N_6984);
and U15725 (N_15725,N_3979,N_1787);
or U15726 (N_15726,N_8817,N_885);
nor U15727 (N_15727,N_8224,N_9280);
or U15728 (N_15728,N_9415,N_4650);
nor U15729 (N_15729,N_5656,N_8594);
nor U15730 (N_15730,N_418,N_1423);
nand U15731 (N_15731,N_669,N_5560);
or U15732 (N_15732,N_4088,N_924);
nor U15733 (N_15733,N_5890,N_1662);
and U15734 (N_15734,N_7703,N_1123);
or U15735 (N_15735,N_5027,N_4515);
or U15736 (N_15736,N_7453,N_594);
nor U15737 (N_15737,N_6543,N_3706);
nor U15738 (N_15738,N_7973,N_4146);
or U15739 (N_15739,N_9008,N_5923);
and U15740 (N_15740,N_5714,N_3216);
or U15741 (N_15741,N_4841,N_174);
or U15742 (N_15742,N_9387,N_3287);
or U15743 (N_15743,N_5577,N_5642);
xor U15744 (N_15744,N_7054,N_821);
xor U15745 (N_15745,N_8543,N_6797);
nand U15746 (N_15746,N_3817,N_2680);
nand U15747 (N_15747,N_4418,N_1111);
nand U15748 (N_15748,N_8270,N_4105);
and U15749 (N_15749,N_6259,N_3971);
or U15750 (N_15750,N_389,N_1178);
nand U15751 (N_15751,N_2488,N_1643);
nor U15752 (N_15752,N_8486,N_386);
nand U15753 (N_15753,N_3449,N_7232);
nand U15754 (N_15754,N_9259,N_71);
and U15755 (N_15755,N_4375,N_9102);
and U15756 (N_15756,N_9224,N_1040);
nor U15757 (N_15757,N_5239,N_5190);
or U15758 (N_15758,N_4300,N_3496);
nand U15759 (N_15759,N_9078,N_3997);
and U15760 (N_15760,N_614,N_9011);
nor U15761 (N_15761,N_7260,N_8775);
nand U15762 (N_15762,N_5294,N_8179);
xnor U15763 (N_15763,N_3037,N_891);
and U15764 (N_15764,N_8014,N_3112);
or U15765 (N_15765,N_169,N_3442);
nor U15766 (N_15766,N_7528,N_4516);
or U15767 (N_15767,N_4540,N_3690);
and U15768 (N_15768,N_5640,N_7593);
nand U15769 (N_15769,N_7220,N_9953);
nor U15770 (N_15770,N_4480,N_13);
and U15771 (N_15771,N_9698,N_8250);
xnor U15772 (N_15772,N_2884,N_2554);
nand U15773 (N_15773,N_7058,N_5957);
or U15774 (N_15774,N_4212,N_4773);
xnor U15775 (N_15775,N_2558,N_6859);
and U15776 (N_15776,N_9106,N_5235);
or U15777 (N_15777,N_6239,N_1685);
or U15778 (N_15778,N_3743,N_8884);
xnor U15779 (N_15779,N_1846,N_9725);
xnor U15780 (N_15780,N_4558,N_1885);
nand U15781 (N_15781,N_5110,N_7107);
nor U15782 (N_15782,N_322,N_6805);
or U15783 (N_15783,N_3981,N_9295);
nor U15784 (N_15784,N_9866,N_8440);
or U15785 (N_15785,N_9086,N_5994);
xor U15786 (N_15786,N_6002,N_1841);
nor U15787 (N_15787,N_512,N_1393);
xnor U15788 (N_15788,N_6159,N_1113);
or U15789 (N_15789,N_9222,N_3974);
and U15790 (N_15790,N_5538,N_7293);
and U15791 (N_15791,N_4733,N_9364);
and U15792 (N_15792,N_1165,N_4051);
or U15793 (N_15793,N_3775,N_6142);
or U15794 (N_15794,N_2341,N_1316);
nand U15795 (N_15795,N_6733,N_3905);
nor U15796 (N_15796,N_1249,N_9682);
and U15797 (N_15797,N_257,N_5244);
or U15798 (N_15798,N_3757,N_6175);
or U15799 (N_15799,N_8812,N_8614);
or U15800 (N_15800,N_5659,N_7791);
and U15801 (N_15801,N_2348,N_5859);
nor U15802 (N_15802,N_8085,N_7848);
nand U15803 (N_15803,N_4712,N_2191);
nor U15804 (N_15804,N_9657,N_1642);
nor U15805 (N_15805,N_4940,N_2599);
nand U15806 (N_15806,N_87,N_463);
or U15807 (N_15807,N_4428,N_9969);
xnor U15808 (N_15808,N_3996,N_9359);
nor U15809 (N_15809,N_3979,N_9247);
nand U15810 (N_15810,N_3970,N_8921);
xnor U15811 (N_15811,N_3163,N_4698);
xor U15812 (N_15812,N_9827,N_3148);
nor U15813 (N_15813,N_2655,N_7347);
or U15814 (N_15814,N_5973,N_707);
nand U15815 (N_15815,N_5221,N_9028);
or U15816 (N_15816,N_6729,N_4466);
nand U15817 (N_15817,N_1727,N_7283);
xor U15818 (N_15818,N_8270,N_5480);
nand U15819 (N_15819,N_9534,N_704);
nor U15820 (N_15820,N_4394,N_6181);
xnor U15821 (N_15821,N_8760,N_2329);
nand U15822 (N_15822,N_2075,N_8141);
and U15823 (N_15823,N_66,N_1953);
nor U15824 (N_15824,N_1760,N_4411);
nand U15825 (N_15825,N_3523,N_2492);
nand U15826 (N_15826,N_1032,N_101);
nor U15827 (N_15827,N_640,N_5511);
or U15828 (N_15828,N_7850,N_6699);
nor U15829 (N_15829,N_1508,N_8844);
or U15830 (N_15830,N_3955,N_7016);
xor U15831 (N_15831,N_4866,N_3220);
and U15832 (N_15832,N_3053,N_6868);
nand U15833 (N_15833,N_9237,N_5246);
nand U15834 (N_15834,N_4025,N_5735);
and U15835 (N_15835,N_408,N_7378);
xnor U15836 (N_15836,N_821,N_448);
nor U15837 (N_15837,N_8888,N_9018);
and U15838 (N_15838,N_4450,N_844);
and U15839 (N_15839,N_5433,N_262);
and U15840 (N_15840,N_2615,N_9764);
nor U15841 (N_15841,N_7623,N_6525);
or U15842 (N_15842,N_1700,N_2401);
nand U15843 (N_15843,N_8403,N_8423);
nand U15844 (N_15844,N_7761,N_5308);
or U15845 (N_15845,N_274,N_9909);
and U15846 (N_15846,N_6572,N_3734);
nand U15847 (N_15847,N_7497,N_7453);
and U15848 (N_15848,N_8049,N_7025);
nand U15849 (N_15849,N_8357,N_223);
xnor U15850 (N_15850,N_7805,N_9248);
or U15851 (N_15851,N_21,N_675);
nand U15852 (N_15852,N_8002,N_9853);
xor U15853 (N_15853,N_5111,N_805);
nor U15854 (N_15854,N_2040,N_2637);
nand U15855 (N_15855,N_360,N_3859);
or U15856 (N_15856,N_7213,N_4365);
nor U15857 (N_15857,N_1890,N_9110);
nand U15858 (N_15858,N_9547,N_342);
xnor U15859 (N_15859,N_9179,N_1537);
nor U15860 (N_15860,N_4683,N_5289);
nand U15861 (N_15861,N_2155,N_439);
or U15862 (N_15862,N_5246,N_1650);
and U15863 (N_15863,N_4235,N_637);
or U15864 (N_15864,N_2205,N_330);
and U15865 (N_15865,N_9301,N_33);
xor U15866 (N_15866,N_385,N_7557);
nor U15867 (N_15867,N_1845,N_803);
xnor U15868 (N_15868,N_6913,N_1139);
nor U15869 (N_15869,N_6924,N_5412);
nor U15870 (N_15870,N_5992,N_104);
or U15871 (N_15871,N_7078,N_3606);
nor U15872 (N_15872,N_2801,N_7107);
and U15873 (N_15873,N_9909,N_6943);
nand U15874 (N_15874,N_2699,N_3723);
and U15875 (N_15875,N_4464,N_8451);
nor U15876 (N_15876,N_7752,N_4075);
nor U15877 (N_15877,N_2222,N_9854);
xnor U15878 (N_15878,N_8798,N_7909);
nand U15879 (N_15879,N_9870,N_84);
nor U15880 (N_15880,N_6782,N_3712);
nand U15881 (N_15881,N_25,N_6923);
or U15882 (N_15882,N_340,N_3531);
xor U15883 (N_15883,N_7017,N_8388);
or U15884 (N_15884,N_8335,N_7621);
or U15885 (N_15885,N_2311,N_3474);
nor U15886 (N_15886,N_7960,N_1104);
xnor U15887 (N_15887,N_6169,N_3678);
nor U15888 (N_15888,N_2308,N_9153);
nor U15889 (N_15889,N_6191,N_9384);
and U15890 (N_15890,N_3695,N_458);
xor U15891 (N_15891,N_7973,N_761);
nor U15892 (N_15892,N_1078,N_8293);
and U15893 (N_15893,N_1781,N_2609);
or U15894 (N_15894,N_604,N_174);
nor U15895 (N_15895,N_4462,N_1452);
and U15896 (N_15896,N_786,N_8632);
nor U15897 (N_15897,N_4619,N_239);
nor U15898 (N_15898,N_221,N_9890);
or U15899 (N_15899,N_7242,N_690);
nand U15900 (N_15900,N_8291,N_4369);
nor U15901 (N_15901,N_8088,N_7397);
and U15902 (N_15902,N_689,N_7846);
and U15903 (N_15903,N_4983,N_4694);
and U15904 (N_15904,N_375,N_995);
nand U15905 (N_15905,N_4166,N_572);
or U15906 (N_15906,N_8690,N_720);
or U15907 (N_15907,N_4780,N_3534);
nor U15908 (N_15908,N_8178,N_2700);
nor U15909 (N_15909,N_4538,N_5185);
nor U15910 (N_15910,N_8562,N_1189);
and U15911 (N_15911,N_3665,N_3754);
and U15912 (N_15912,N_7849,N_2177);
and U15913 (N_15913,N_8723,N_7583);
and U15914 (N_15914,N_6914,N_2701);
and U15915 (N_15915,N_5704,N_3782);
or U15916 (N_15916,N_2079,N_2215);
and U15917 (N_15917,N_6874,N_1990);
or U15918 (N_15918,N_3462,N_9739);
or U15919 (N_15919,N_5024,N_8889);
nand U15920 (N_15920,N_5662,N_5939);
or U15921 (N_15921,N_8548,N_8807);
nor U15922 (N_15922,N_8076,N_8467);
nand U15923 (N_15923,N_5497,N_5713);
nand U15924 (N_15924,N_2971,N_1180);
xnor U15925 (N_15925,N_3582,N_9551);
and U15926 (N_15926,N_9627,N_4333);
nand U15927 (N_15927,N_8689,N_6820);
nand U15928 (N_15928,N_5114,N_8299);
and U15929 (N_15929,N_8725,N_5658);
and U15930 (N_15930,N_576,N_3090);
or U15931 (N_15931,N_4277,N_7941);
nor U15932 (N_15932,N_6980,N_5700);
or U15933 (N_15933,N_283,N_714);
nor U15934 (N_15934,N_5176,N_788);
nand U15935 (N_15935,N_5068,N_5451);
or U15936 (N_15936,N_251,N_2833);
nor U15937 (N_15937,N_7471,N_8629);
nand U15938 (N_15938,N_9456,N_7099);
and U15939 (N_15939,N_3799,N_2133);
nor U15940 (N_15940,N_7578,N_3162);
and U15941 (N_15941,N_277,N_3521);
nor U15942 (N_15942,N_306,N_154);
nand U15943 (N_15943,N_149,N_3422);
nand U15944 (N_15944,N_9745,N_1961);
nor U15945 (N_15945,N_2310,N_100);
nor U15946 (N_15946,N_2152,N_5982);
xor U15947 (N_15947,N_4293,N_2156);
nand U15948 (N_15948,N_8493,N_6089);
nand U15949 (N_15949,N_6407,N_7882);
nor U15950 (N_15950,N_7736,N_597);
nand U15951 (N_15951,N_4200,N_3469);
and U15952 (N_15952,N_7712,N_6246);
or U15953 (N_15953,N_8660,N_4729);
or U15954 (N_15954,N_7741,N_8279);
xor U15955 (N_15955,N_5289,N_2339);
nor U15956 (N_15956,N_8516,N_8970);
xor U15957 (N_15957,N_9012,N_5481);
nand U15958 (N_15958,N_7493,N_5386);
xor U15959 (N_15959,N_7273,N_1093);
nor U15960 (N_15960,N_5561,N_7387);
nand U15961 (N_15961,N_8781,N_7854);
nand U15962 (N_15962,N_8337,N_6147);
nand U15963 (N_15963,N_9576,N_6561);
and U15964 (N_15964,N_5110,N_7204);
or U15965 (N_15965,N_9416,N_912);
and U15966 (N_15966,N_8281,N_7889);
or U15967 (N_15967,N_4504,N_2228);
nor U15968 (N_15968,N_9369,N_4193);
xor U15969 (N_15969,N_4415,N_6341);
nor U15970 (N_15970,N_4086,N_9363);
xnor U15971 (N_15971,N_8530,N_461);
nand U15972 (N_15972,N_8382,N_7453);
or U15973 (N_15973,N_5255,N_4975);
and U15974 (N_15974,N_4797,N_5672);
nor U15975 (N_15975,N_9701,N_3003);
and U15976 (N_15976,N_6783,N_8253);
and U15977 (N_15977,N_8760,N_8330);
and U15978 (N_15978,N_644,N_7065);
or U15979 (N_15979,N_6321,N_1763);
xor U15980 (N_15980,N_3265,N_1020);
nand U15981 (N_15981,N_7529,N_2156);
nor U15982 (N_15982,N_7649,N_2601);
and U15983 (N_15983,N_9913,N_2518);
nand U15984 (N_15984,N_7138,N_6203);
nand U15985 (N_15985,N_2307,N_6637);
nand U15986 (N_15986,N_7498,N_6685);
and U15987 (N_15987,N_9223,N_425);
and U15988 (N_15988,N_1933,N_2461);
nor U15989 (N_15989,N_9976,N_7816);
nor U15990 (N_15990,N_1410,N_366);
nand U15991 (N_15991,N_5680,N_1939);
nor U15992 (N_15992,N_5530,N_5930);
nor U15993 (N_15993,N_3518,N_9249);
xor U15994 (N_15994,N_3992,N_8594);
nand U15995 (N_15995,N_2590,N_6797);
and U15996 (N_15996,N_3289,N_7483);
and U15997 (N_15997,N_5956,N_6230);
nand U15998 (N_15998,N_2777,N_4559);
and U15999 (N_15999,N_6335,N_5682);
or U16000 (N_16000,N_8712,N_8495);
and U16001 (N_16001,N_8323,N_5604);
and U16002 (N_16002,N_1751,N_5227);
or U16003 (N_16003,N_9463,N_3937);
and U16004 (N_16004,N_7002,N_8888);
nor U16005 (N_16005,N_7125,N_394);
or U16006 (N_16006,N_3675,N_9596);
xor U16007 (N_16007,N_1188,N_3791);
nand U16008 (N_16008,N_9075,N_4250);
and U16009 (N_16009,N_2475,N_1016);
nor U16010 (N_16010,N_6442,N_742);
nor U16011 (N_16011,N_6351,N_3567);
nor U16012 (N_16012,N_4562,N_3408);
or U16013 (N_16013,N_9034,N_1293);
nand U16014 (N_16014,N_6707,N_6944);
nor U16015 (N_16015,N_7214,N_4546);
and U16016 (N_16016,N_276,N_122);
or U16017 (N_16017,N_4084,N_9631);
and U16018 (N_16018,N_4140,N_5133);
nor U16019 (N_16019,N_2628,N_2204);
and U16020 (N_16020,N_5474,N_6934);
or U16021 (N_16021,N_94,N_8973);
and U16022 (N_16022,N_6708,N_2457);
and U16023 (N_16023,N_757,N_6794);
nand U16024 (N_16024,N_373,N_3189);
or U16025 (N_16025,N_2633,N_4651);
nor U16026 (N_16026,N_3057,N_2643);
nand U16027 (N_16027,N_9099,N_6793);
or U16028 (N_16028,N_8943,N_5508);
nor U16029 (N_16029,N_9937,N_9202);
and U16030 (N_16030,N_9301,N_940);
and U16031 (N_16031,N_7792,N_3466);
nand U16032 (N_16032,N_604,N_1692);
and U16033 (N_16033,N_6087,N_6507);
or U16034 (N_16034,N_7168,N_8466);
nor U16035 (N_16035,N_2175,N_3057);
and U16036 (N_16036,N_4188,N_6856);
or U16037 (N_16037,N_1093,N_3385);
and U16038 (N_16038,N_4935,N_2997);
and U16039 (N_16039,N_7118,N_217);
or U16040 (N_16040,N_2669,N_3379);
and U16041 (N_16041,N_2947,N_3219);
nand U16042 (N_16042,N_2032,N_8903);
or U16043 (N_16043,N_2181,N_1772);
or U16044 (N_16044,N_1515,N_7503);
and U16045 (N_16045,N_677,N_7015);
nor U16046 (N_16046,N_4865,N_3330);
xnor U16047 (N_16047,N_6725,N_9195);
and U16048 (N_16048,N_1909,N_8912);
or U16049 (N_16049,N_9532,N_4352);
or U16050 (N_16050,N_4764,N_2391);
nor U16051 (N_16051,N_9604,N_9467);
and U16052 (N_16052,N_2290,N_3541);
and U16053 (N_16053,N_827,N_4707);
nand U16054 (N_16054,N_7985,N_4060);
xnor U16055 (N_16055,N_5615,N_3650);
and U16056 (N_16056,N_8133,N_6096);
or U16057 (N_16057,N_6549,N_1232);
or U16058 (N_16058,N_937,N_7701);
or U16059 (N_16059,N_6145,N_7828);
nor U16060 (N_16060,N_9460,N_7700);
xor U16061 (N_16061,N_8030,N_1087);
nand U16062 (N_16062,N_2922,N_1449);
nand U16063 (N_16063,N_413,N_6647);
nor U16064 (N_16064,N_4279,N_417);
nor U16065 (N_16065,N_6640,N_6797);
and U16066 (N_16066,N_7833,N_9161);
nand U16067 (N_16067,N_5781,N_8803);
xnor U16068 (N_16068,N_9902,N_4856);
nor U16069 (N_16069,N_590,N_1132);
nand U16070 (N_16070,N_1193,N_9492);
or U16071 (N_16071,N_8555,N_9138);
nand U16072 (N_16072,N_2875,N_9926);
or U16073 (N_16073,N_2185,N_9470);
nand U16074 (N_16074,N_9563,N_3103);
nand U16075 (N_16075,N_3814,N_2964);
nor U16076 (N_16076,N_5166,N_5185);
nand U16077 (N_16077,N_4378,N_6070);
and U16078 (N_16078,N_2018,N_5423);
and U16079 (N_16079,N_8285,N_9048);
nor U16080 (N_16080,N_8070,N_7139);
nand U16081 (N_16081,N_5625,N_107);
nand U16082 (N_16082,N_30,N_6361);
nor U16083 (N_16083,N_117,N_7907);
or U16084 (N_16084,N_5840,N_3077);
nor U16085 (N_16085,N_1484,N_5006);
nor U16086 (N_16086,N_6581,N_9798);
nand U16087 (N_16087,N_1246,N_8813);
and U16088 (N_16088,N_6429,N_9993);
nand U16089 (N_16089,N_4507,N_5688);
nand U16090 (N_16090,N_2320,N_4336);
or U16091 (N_16091,N_1499,N_2631);
or U16092 (N_16092,N_6748,N_7291);
nor U16093 (N_16093,N_9706,N_125);
and U16094 (N_16094,N_9767,N_4424);
nand U16095 (N_16095,N_5304,N_8130);
and U16096 (N_16096,N_5207,N_9550);
nand U16097 (N_16097,N_9341,N_6762);
or U16098 (N_16098,N_5644,N_5070);
nand U16099 (N_16099,N_5534,N_4394);
and U16100 (N_16100,N_6031,N_8736);
nor U16101 (N_16101,N_1940,N_6749);
or U16102 (N_16102,N_2765,N_8480);
or U16103 (N_16103,N_6706,N_5751);
nor U16104 (N_16104,N_2617,N_6235);
xor U16105 (N_16105,N_5334,N_8425);
nor U16106 (N_16106,N_8272,N_2727);
or U16107 (N_16107,N_2226,N_3716);
nor U16108 (N_16108,N_1,N_803);
and U16109 (N_16109,N_9027,N_2293);
nor U16110 (N_16110,N_4405,N_2674);
and U16111 (N_16111,N_845,N_800);
nor U16112 (N_16112,N_6482,N_4716);
or U16113 (N_16113,N_926,N_652);
xnor U16114 (N_16114,N_8896,N_2894);
nand U16115 (N_16115,N_3625,N_916);
and U16116 (N_16116,N_2948,N_6788);
or U16117 (N_16117,N_2337,N_8480);
and U16118 (N_16118,N_590,N_3349);
nand U16119 (N_16119,N_6346,N_962);
nor U16120 (N_16120,N_7659,N_5684);
nand U16121 (N_16121,N_7845,N_5621);
nand U16122 (N_16122,N_5242,N_9334);
and U16123 (N_16123,N_59,N_7320);
nor U16124 (N_16124,N_4534,N_8822);
and U16125 (N_16125,N_7441,N_5152);
nor U16126 (N_16126,N_9242,N_7726);
and U16127 (N_16127,N_5254,N_4952);
xor U16128 (N_16128,N_2866,N_2102);
nand U16129 (N_16129,N_6764,N_318);
nor U16130 (N_16130,N_6726,N_8990);
or U16131 (N_16131,N_9400,N_9621);
nor U16132 (N_16132,N_8749,N_337);
or U16133 (N_16133,N_4997,N_9130);
nand U16134 (N_16134,N_1786,N_1524);
or U16135 (N_16135,N_4993,N_6714);
nand U16136 (N_16136,N_2865,N_1244);
or U16137 (N_16137,N_5128,N_3673);
or U16138 (N_16138,N_6958,N_7154);
and U16139 (N_16139,N_9786,N_5672);
or U16140 (N_16140,N_372,N_6635);
nor U16141 (N_16141,N_5468,N_2121);
nand U16142 (N_16142,N_3975,N_1643);
and U16143 (N_16143,N_1261,N_9348);
or U16144 (N_16144,N_7131,N_7057);
and U16145 (N_16145,N_1400,N_2877);
and U16146 (N_16146,N_5903,N_4177);
nor U16147 (N_16147,N_1794,N_2944);
or U16148 (N_16148,N_7560,N_1298);
and U16149 (N_16149,N_3123,N_3217);
nand U16150 (N_16150,N_8531,N_7364);
xor U16151 (N_16151,N_5413,N_5575);
nand U16152 (N_16152,N_6734,N_9682);
or U16153 (N_16153,N_3367,N_4458);
and U16154 (N_16154,N_6757,N_5580);
nor U16155 (N_16155,N_6849,N_2411);
nand U16156 (N_16156,N_4861,N_4416);
or U16157 (N_16157,N_337,N_707);
and U16158 (N_16158,N_4022,N_3175);
or U16159 (N_16159,N_3424,N_6233);
nand U16160 (N_16160,N_854,N_5784);
nand U16161 (N_16161,N_7941,N_7140);
or U16162 (N_16162,N_3435,N_4866);
nand U16163 (N_16163,N_3132,N_1486);
nor U16164 (N_16164,N_1532,N_5328);
xnor U16165 (N_16165,N_6011,N_5938);
nor U16166 (N_16166,N_9326,N_4352);
and U16167 (N_16167,N_7395,N_903);
nand U16168 (N_16168,N_8785,N_4494);
nor U16169 (N_16169,N_2768,N_9773);
nand U16170 (N_16170,N_7866,N_2296);
or U16171 (N_16171,N_1644,N_3074);
nor U16172 (N_16172,N_1298,N_7684);
nor U16173 (N_16173,N_2392,N_7629);
and U16174 (N_16174,N_3836,N_2112);
or U16175 (N_16175,N_2501,N_6145);
nand U16176 (N_16176,N_7557,N_3501);
xnor U16177 (N_16177,N_8207,N_1361);
xor U16178 (N_16178,N_3512,N_8214);
nor U16179 (N_16179,N_1497,N_1514);
or U16180 (N_16180,N_3478,N_308);
xor U16181 (N_16181,N_4394,N_1371);
nor U16182 (N_16182,N_8723,N_5299);
and U16183 (N_16183,N_7234,N_9148);
and U16184 (N_16184,N_9371,N_4135);
nand U16185 (N_16185,N_8477,N_4673);
and U16186 (N_16186,N_5902,N_7789);
nand U16187 (N_16187,N_1307,N_7819);
or U16188 (N_16188,N_8043,N_9898);
nor U16189 (N_16189,N_6215,N_1527);
nand U16190 (N_16190,N_5461,N_6294);
or U16191 (N_16191,N_9738,N_5818);
nand U16192 (N_16192,N_670,N_3454);
and U16193 (N_16193,N_3841,N_1170);
or U16194 (N_16194,N_1088,N_4083);
xor U16195 (N_16195,N_4777,N_4582);
nor U16196 (N_16196,N_7567,N_4095);
nor U16197 (N_16197,N_2258,N_2636);
nand U16198 (N_16198,N_2277,N_3169);
and U16199 (N_16199,N_335,N_3837);
nor U16200 (N_16200,N_5173,N_5697);
and U16201 (N_16201,N_4598,N_5446);
nand U16202 (N_16202,N_1451,N_4233);
and U16203 (N_16203,N_4455,N_8396);
nor U16204 (N_16204,N_5382,N_4004);
or U16205 (N_16205,N_7167,N_653);
or U16206 (N_16206,N_2495,N_8501);
nand U16207 (N_16207,N_7312,N_9563);
nand U16208 (N_16208,N_3996,N_6317);
or U16209 (N_16209,N_2502,N_6622);
and U16210 (N_16210,N_2392,N_4828);
nor U16211 (N_16211,N_9360,N_138);
nand U16212 (N_16212,N_8815,N_1348);
nor U16213 (N_16213,N_7045,N_917);
nor U16214 (N_16214,N_425,N_8324);
nor U16215 (N_16215,N_1223,N_6097);
and U16216 (N_16216,N_7386,N_4935);
xor U16217 (N_16217,N_937,N_2613);
nor U16218 (N_16218,N_3993,N_779);
nand U16219 (N_16219,N_4002,N_2749);
nor U16220 (N_16220,N_8826,N_6143);
xor U16221 (N_16221,N_9292,N_8612);
and U16222 (N_16222,N_3712,N_3201);
nor U16223 (N_16223,N_6512,N_35);
and U16224 (N_16224,N_171,N_3374);
and U16225 (N_16225,N_1207,N_9715);
and U16226 (N_16226,N_6341,N_9147);
or U16227 (N_16227,N_9140,N_3034);
or U16228 (N_16228,N_7586,N_5830);
or U16229 (N_16229,N_4231,N_8749);
nor U16230 (N_16230,N_8631,N_5107);
or U16231 (N_16231,N_2263,N_9974);
or U16232 (N_16232,N_7566,N_3857);
and U16233 (N_16233,N_2643,N_5697);
or U16234 (N_16234,N_8548,N_8015);
nor U16235 (N_16235,N_6277,N_6527);
or U16236 (N_16236,N_1266,N_8278);
and U16237 (N_16237,N_6559,N_6086);
nand U16238 (N_16238,N_3626,N_4145);
nor U16239 (N_16239,N_7447,N_6038);
and U16240 (N_16240,N_9595,N_320);
or U16241 (N_16241,N_7398,N_2722);
nor U16242 (N_16242,N_234,N_9320);
or U16243 (N_16243,N_8088,N_3997);
nand U16244 (N_16244,N_6679,N_1305);
nor U16245 (N_16245,N_9359,N_5589);
nand U16246 (N_16246,N_1807,N_2702);
nor U16247 (N_16247,N_2839,N_6088);
nor U16248 (N_16248,N_7676,N_9515);
nand U16249 (N_16249,N_4447,N_3122);
and U16250 (N_16250,N_440,N_5612);
or U16251 (N_16251,N_4691,N_2086);
nand U16252 (N_16252,N_5961,N_9370);
or U16253 (N_16253,N_7684,N_7744);
and U16254 (N_16254,N_3601,N_4109);
nand U16255 (N_16255,N_1835,N_66);
nand U16256 (N_16256,N_4887,N_785);
and U16257 (N_16257,N_9551,N_4548);
nand U16258 (N_16258,N_684,N_9266);
or U16259 (N_16259,N_7499,N_4542);
and U16260 (N_16260,N_8198,N_470);
and U16261 (N_16261,N_8036,N_2077);
and U16262 (N_16262,N_725,N_9471);
nand U16263 (N_16263,N_5557,N_6503);
and U16264 (N_16264,N_6831,N_3156);
nor U16265 (N_16265,N_4366,N_9681);
nor U16266 (N_16266,N_983,N_7319);
nor U16267 (N_16267,N_6020,N_2147);
nor U16268 (N_16268,N_963,N_3982);
nand U16269 (N_16269,N_4135,N_1335);
or U16270 (N_16270,N_4623,N_6358);
or U16271 (N_16271,N_5577,N_8688);
and U16272 (N_16272,N_2814,N_6518);
nand U16273 (N_16273,N_7317,N_7476);
nor U16274 (N_16274,N_9481,N_5817);
and U16275 (N_16275,N_4981,N_9662);
nor U16276 (N_16276,N_2102,N_3040);
or U16277 (N_16277,N_6038,N_6030);
xor U16278 (N_16278,N_9728,N_1786);
nand U16279 (N_16279,N_6362,N_2868);
or U16280 (N_16280,N_2879,N_1705);
and U16281 (N_16281,N_2049,N_28);
nor U16282 (N_16282,N_8338,N_1391);
and U16283 (N_16283,N_915,N_5978);
or U16284 (N_16284,N_4335,N_3228);
or U16285 (N_16285,N_4362,N_2523);
nor U16286 (N_16286,N_9636,N_9707);
xor U16287 (N_16287,N_7944,N_773);
nand U16288 (N_16288,N_1807,N_1066);
or U16289 (N_16289,N_2458,N_90);
nand U16290 (N_16290,N_1963,N_3515);
or U16291 (N_16291,N_1115,N_5818);
and U16292 (N_16292,N_604,N_8491);
or U16293 (N_16293,N_4465,N_9297);
or U16294 (N_16294,N_234,N_4781);
nor U16295 (N_16295,N_5267,N_2805);
xor U16296 (N_16296,N_5049,N_3435);
nand U16297 (N_16297,N_9201,N_7494);
xor U16298 (N_16298,N_1818,N_1372);
and U16299 (N_16299,N_3179,N_4734);
nand U16300 (N_16300,N_3058,N_7957);
nand U16301 (N_16301,N_2172,N_2445);
or U16302 (N_16302,N_8702,N_2018);
or U16303 (N_16303,N_5000,N_4817);
xnor U16304 (N_16304,N_2120,N_4724);
or U16305 (N_16305,N_354,N_8752);
or U16306 (N_16306,N_6799,N_1129);
and U16307 (N_16307,N_7350,N_4232);
nor U16308 (N_16308,N_1614,N_6395);
and U16309 (N_16309,N_9030,N_5742);
and U16310 (N_16310,N_2975,N_2148);
or U16311 (N_16311,N_2740,N_4258);
nor U16312 (N_16312,N_3393,N_1233);
nor U16313 (N_16313,N_2523,N_5196);
and U16314 (N_16314,N_5868,N_9674);
and U16315 (N_16315,N_1819,N_1574);
nand U16316 (N_16316,N_1626,N_4910);
nand U16317 (N_16317,N_537,N_9308);
or U16318 (N_16318,N_323,N_7610);
nand U16319 (N_16319,N_290,N_3960);
nor U16320 (N_16320,N_1973,N_5126);
xor U16321 (N_16321,N_3802,N_4688);
or U16322 (N_16322,N_8717,N_3947);
nor U16323 (N_16323,N_209,N_5172);
nor U16324 (N_16324,N_2309,N_7639);
nor U16325 (N_16325,N_2881,N_7250);
or U16326 (N_16326,N_7842,N_9221);
or U16327 (N_16327,N_2240,N_931);
or U16328 (N_16328,N_2665,N_2162);
nor U16329 (N_16329,N_475,N_5730);
or U16330 (N_16330,N_4994,N_2733);
and U16331 (N_16331,N_5906,N_7099);
and U16332 (N_16332,N_6264,N_6916);
nand U16333 (N_16333,N_7016,N_3519);
nor U16334 (N_16334,N_136,N_6594);
or U16335 (N_16335,N_3230,N_4337);
nand U16336 (N_16336,N_8910,N_1007);
and U16337 (N_16337,N_5282,N_4673);
nor U16338 (N_16338,N_4566,N_9193);
nand U16339 (N_16339,N_7040,N_7595);
or U16340 (N_16340,N_9772,N_8081);
and U16341 (N_16341,N_9635,N_2434);
or U16342 (N_16342,N_5947,N_3781);
nor U16343 (N_16343,N_9946,N_7236);
xnor U16344 (N_16344,N_7102,N_1389);
and U16345 (N_16345,N_1704,N_7888);
xor U16346 (N_16346,N_4455,N_6641);
nand U16347 (N_16347,N_9814,N_8023);
nand U16348 (N_16348,N_2925,N_7403);
or U16349 (N_16349,N_3648,N_5425);
nor U16350 (N_16350,N_9606,N_8430);
or U16351 (N_16351,N_7410,N_8930);
nor U16352 (N_16352,N_576,N_8914);
or U16353 (N_16353,N_5157,N_1177);
nor U16354 (N_16354,N_5229,N_9606);
nor U16355 (N_16355,N_8859,N_1195);
nor U16356 (N_16356,N_8342,N_1636);
or U16357 (N_16357,N_4812,N_6710);
xnor U16358 (N_16358,N_1515,N_2004);
or U16359 (N_16359,N_1748,N_7381);
and U16360 (N_16360,N_8663,N_5232);
nor U16361 (N_16361,N_2463,N_8693);
or U16362 (N_16362,N_7623,N_5786);
nor U16363 (N_16363,N_5521,N_3253);
and U16364 (N_16364,N_3304,N_7071);
nand U16365 (N_16365,N_2877,N_1260);
nand U16366 (N_16366,N_7860,N_4211);
and U16367 (N_16367,N_3463,N_8974);
or U16368 (N_16368,N_7391,N_6511);
or U16369 (N_16369,N_577,N_789);
and U16370 (N_16370,N_4534,N_6313);
nor U16371 (N_16371,N_540,N_9883);
nand U16372 (N_16372,N_7209,N_1879);
xor U16373 (N_16373,N_880,N_2395);
nand U16374 (N_16374,N_1150,N_5428);
or U16375 (N_16375,N_2270,N_8503);
nor U16376 (N_16376,N_3683,N_3607);
nand U16377 (N_16377,N_7371,N_8283);
or U16378 (N_16378,N_1076,N_5431);
nor U16379 (N_16379,N_7849,N_2104);
or U16380 (N_16380,N_2690,N_3101);
nand U16381 (N_16381,N_8647,N_5426);
nor U16382 (N_16382,N_9434,N_1559);
and U16383 (N_16383,N_5980,N_8403);
or U16384 (N_16384,N_8871,N_4237);
or U16385 (N_16385,N_6418,N_1348);
nor U16386 (N_16386,N_4377,N_7693);
nor U16387 (N_16387,N_6556,N_4622);
nor U16388 (N_16388,N_2201,N_9521);
or U16389 (N_16389,N_4656,N_6819);
xnor U16390 (N_16390,N_7361,N_5304);
nand U16391 (N_16391,N_5625,N_6098);
nor U16392 (N_16392,N_6887,N_5763);
or U16393 (N_16393,N_8989,N_2745);
nor U16394 (N_16394,N_6141,N_7078);
and U16395 (N_16395,N_8580,N_5765);
nor U16396 (N_16396,N_2752,N_1060);
xnor U16397 (N_16397,N_4525,N_7852);
xnor U16398 (N_16398,N_948,N_1838);
nand U16399 (N_16399,N_269,N_4129);
nand U16400 (N_16400,N_7567,N_3111);
xnor U16401 (N_16401,N_9513,N_613);
and U16402 (N_16402,N_6117,N_6946);
nand U16403 (N_16403,N_4878,N_4432);
and U16404 (N_16404,N_5681,N_2369);
or U16405 (N_16405,N_4252,N_4108);
nor U16406 (N_16406,N_5600,N_3366);
or U16407 (N_16407,N_3295,N_6029);
nor U16408 (N_16408,N_3761,N_3301);
and U16409 (N_16409,N_8262,N_9537);
nor U16410 (N_16410,N_3196,N_4806);
or U16411 (N_16411,N_4001,N_4130);
nor U16412 (N_16412,N_5965,N_7185);
nor U16413 (N_16413,N_4771,N_356);
nand U16414 (N_16414,N_520,N_2480);
or U16415 (N_16415,N_7667,N_7185);
nor U16416 (N_16416,N_8079,N_5195);
nand U16417 (N_16417,N_5390,N_6794);
nand U16418 (N_16418,N_4147,N_7014);
and U16419 (N_16419,N_735,N_7748);
or U16420 (N_16420,N_6691,N_981);
nor U16421 (N_16421,N_9486,N_4021);
nand U16422 (N_16422,N_6103,N_5580);
xor U16423 (N_16423,N_7025,N_3301);
or U16424 (N_16424,N_6749,N_2416);
and U16425 (N_16425,N_3618,N_7198);
nand U16426 (N_16426,N_8641,N_2853);
or U16427 (N_16427,N_4580,N_2891);
or U16428 (N_16428,N_2457,N_9302);
and U16429 (N_16429,N_9016,N_2931);
and U16430 (N_16430,N_8771,N_6761);
or U16431 (N_16431,N_4259,N_4501);
nor U16432 (N_16432,N_2955,N_4706);
and U16433 (N_16433,N_9998,N_235);
and U16434 (N_16434,N_9783,N_8836);
nand U16435 (N_16435,N_112,N_1558);
nand U16436 (N_16436,N_6077,N_5205);
nand U16437 (N_16437,N_5006,N_3353);
or U16438 (N_16438,N_9738,N_2218);
and U16439 (N_16439,N_159,N_7892);
or U16440 (N_16440,N_2980,N_9465);
and U16441 (N_16441,N_6996,N_369);
nand U16442 (N_16442,N_9316,N_5832);
or U16443 (N_16443,N_6781,N_8194);
nor U16444 (N_16444,N_311,N_1225);
nor U16445 (N_16445,N_1823,N_9074);
or U16446 (N_16446,N_3340,N_3583);
or U16447 (N_16447,N_7714,N_4852);
and U16448 (N_16448,N_8211,N_2370);
and U16449 (N_16449,N_4341,N_7807);
and U16450 (N_16450,N_4914,N_5994);
or U16451 (N_16451,N_9100,N_9729);
or U16452 (N_16452,N_7901,N_8864);
nor U16453 (N_16453,N_2528,N_2265);
or U16454 (N_16454,N_9798,N_958);
nand U16455 (N_16455,N_7247,N_7640);
and U16456 (N_16456,N_3727,N_4497);
and U16457 (N_16457,N_8665,N_3712);
or U16458 (N_16458,N_8955,N_6548);
nor U16459 (N_16459,N_4149,N_8697);
nor U16460 (N_16460,N_893,N_287);
and U16461 (N_16461,N_67,N_1557);
or U16462 (N_16462,N_6362,N_7863);
nor U16463 (N_16463,N_406,N_9883);
and U16464 (N_16464,N_7613,N_7961);
or U16465 (N_16465,N_9554,N_1240);
nor U16466 (N_16466,N_4462,N_2019);
or U16467 (N_16467,N_1613,N_9877);
and U16468 (N_16468,N_3120,N_9697);
or U16469 (N_16469,N_2008,N_1532);
or U16470 (N_16470,N_1198,N_2416);
nand U16471 (N_16471,N_6536,N_6489);
and U16472 (N_16472,N_7552,N_6573);
nand U16473 (N_16473,N_6789,N_6144);
nor U16474 (N_16474,N_4208,N_4407);
nand U16475 (N_16475,N_9081,N_9450);
nor U16476 (N_16476,N_3258,N_9310);
and U16477 (N_16477,N_8456,N_7585);
and U16478 (N_16478,N_7930,N_7057);
and U16479 (N_16479,N_4866,N_2389);
or U16480 (N_16480,N_3098,N_6647);
nor U16481 (N_16481,N_9518,N_8233);
nor U16482 (N_16482,N_1519,N_1906);
nor U16483 (N_16483,N_5193,N_2725);
nand U16484 (N_16484,N_5108,N_2379);
and U16485 (N_16485,N_8910,N_2581);
or U16486 (N_16486,N_31,N_9119);
nor U16487 (N_16487,N_7226,N_241);
nand U16488 (N_16488,N_7584,N_8077);
or U16489 (N_16489,N_8353,N_7054);
and U16490 (N_16490,N_4386,N_5441);
nor U16491 (N_16491,N_3305,N_9752);
and U16492 (N_16492,N_4766,N_4051);
and U16493 (N_16493,N_9967,N_9664);
nor U16494 (N_16494,N_2812,N_1115);
or U16495 (N_16495,N_6955,N_4885);
or U16496 (N_16496,N_488,N_2391);
nor U16497 (N_16497,N_3064,N_2566);
or U16498 (N_16498,N_443,N_8049);
or U16499 (N_16499,N_8188,N_8753);
and U16500 (N_16500,N_8715,N_5228);
nor U16501 (N_16501,N_6815,N_4095);
nor U16502 (N_16502,N_4879,N_7347);
nor U16503 (N_16503,N_1713,N_424);
nand U16504 (N_16504,N_9700,N_4524);
nor U16505 (N_16505,N_4160,N_3787);
and U16506 (N_16506,N_2746,N_3964);
or U16507 (N_16507,N_7867,N_7007);
or U16508 (N_16508,N_1949,N_895);
and U16509 (N_16509,N_1148,N_7968);
and U16510 (N_16510,N_2916,N_6598);
nand U16511 (N_16511,N_4882,N_3716);
or U16512 (N_16512,N_372,N_4903);
or U16513 (N_16513,N_8645,N_3872);
or U16514 (N_16514,N_3630,N_8134);
nor U16515 (N_16515,N_2041,N_2953);
nand U16516 (N_16516,N_1575,N_8572);
nor U16517 (N_16517,N_2852,N_1092);
or U16518 (N_16518,N_5809,N_2836);
nor U16519 (N_16519,N_841,N_150);
and U16520 (N_16520,N_1614,N_1172);
and U16521 (N_16521,N_2384,N_2621);
and U16522 (N_16522,N_7732,N_6080);
or U16523 (N_16523,N_8562,N_3543);
nand U16524 (N_16524,N_7779,N_3952);
or U16525 (N_16525,N_48,N_2493);
or U16526 (N_16526,N_2688,N_8101);
nand U16527 (N_16527,N_1607,N_9293);
or U16528 (N_16528,N_3493,N_5564);
xnor U16529 (N_16529,N_2522,N_3584);
or U16530 (N_16530,N_5344,N_8906);
nand U16531 (N_16531,N_6320,N_820);
xnor U16532 (N_16532,N_8556,N_6009);
and U16533 (N_16533,N_9093,N_3107);
and U16534 (N_16534,N_9202,N_3219);
nand U16535 (N_16535,N_1617,N_4689);
or U16536 (N_16536,N_772,N_3948);
nor U16537 (N_16537,N_8643,N_8405);
xnor U16538 (N_16538,N_5557,N_2196);
xor U16539 (N_16539,N_4235,N_6679);
and U16540 (N_16540,N_4641,N_5588);
nand U16541 (N_16541,N_8712,N_4864);
and U16542 (N_16542,N_6889,N_2642);
nor U16543 (N_16543,N_211,N_1854);
or U16544 (N_16544,N_2417,N_8392);
or U16545 (N_16545,N_8996,N_6419);
and U16546 (N_16546,N_8200,N_7829);
nor U16547 (N_16547,N_1918,N_4698);
and U16548 (N_16548,N_397,N_883);
and U16549 (N_16549,N_9527,N_3356);
or U16550 (N_16550,N_465,N_6386);
and U16551 (N_16551,N_7137,N_3027);
nor U16552 (N_16552,N_809,N_580);
or U16553 (N_16553,N_8866,N_5337);
or U16554 (N_16554,N_3873,N_9500);
xor U16555 (N_16555,N_4670,N_7270);
nor U16556 (N_16556,N_2122,N_7753);
or U16557 (N_16557,N_7760,N_5359);
and U16558 (N_16558,N_1606,N_9416);
nand U16559 (N_16559,N_3768,N_898);
nor U16560 (N_16560,N_9982,N_4783);
nand U16561 (N_16561,N_7794,N_1523);
nor U16562 (N_16562,N_4805,N_1549);
nor U16563 (N_16563,N_5972,N_9572);
or U16564 (N_16564,N_1307,N_961);
nand U16565 (N_16565,N_2505,N_6330);
and U16566 (N_16566,N_6073,N_3709);
nor U16567 (N_16567,N_4415,N_8969);
nand U16568 (N_16568,N_5233,N_1131);
or U16569 (N_16569,N_7692,N_8852);
or U16570 (N_16570,N_5443,N_7161);
nor U16571 (N_16571,N_4705,N_9048);
nor U16572 (N_16572,N_630,N_2834);
or U16573 (N_16573,N_2293,N_9877);
nor U16574 (N_16574,N_777,N_8881);
nor U16575 (N_16575,N_1786,N_2127);
nor U16576 (N_16576,N_3235,N_9252);
nor U16577 (N_16577,N_4664,N_5559);
or U16578 (N_16578,N_6356,N_9782);
and U16579 (N_16579,N_2873,N_3024);
nor U16580 (N_16580,N_2883,N_42);
and U16581 (N_16581,N_4743,N_9095);
nand U16582 (N_16582,N_4770,N_3529);
xor U16583 (N_16583,N_7232,N_1474);
nand U16584 (N_16584,N_5992,N_4789);
nor U16585 (N_16585,N_3009,N_7899);
nor U16586 (N_16586,N_7941,N_2150);
nand U16587 (N_16587,N_30,N_4466);
xnor U16588 (N_16588,N_4244,N_8700);
xnor U16589 (N_16589,N_6370,N_7644);
or U16590 (N_16590,N_789,N_8982);
or U16591 (N_16591,N_5640,N_1311);
or U16592 (N_16592,N_2267,N_4457);
and U16593 (N_16593,N_3740,N_7313);
nand U16594 (N_16594,N_6510,N_9606);
nor U16595 (N_16595,N_1175,N_7621);
or U16596 (N_16596,N_2160,N_9134);
nand U16597 (N_16597,N_1810,N_5484);
nand U16598 (N_16598,N_2351,N_6390);
xor U16599 (N_16599,N_6867,N_3744);
or U16600 (N_16600,N_5350,N_5037);
and U16601 (N_16601,N_5525,N_6860);
nor U16602 (N_16602,N_922,N_8668);
or U16603 (N_16603,N_32,N_6359);
or U16604 (N_16604,N_6916,N_1453);
and U16605 (N_16605,N_5298,N_6527);
nor U16606 (N_16606,N_8108,N_7330);
nor U16607 (N_16607,N_5659,N_4209);
nor U16608 (N_16608,N_6161,N_8382);
and U16609 (N_16609,N_4260,N_1528);
xnor U16610 (N_16610,N_4102,N_3813);
nor U16611 (N_16611,N_2474,N_6457);
and U16612 (N_16612,N_4757,N_7610);
and U16613 (N_16613,N_1605,N_9034);
nand U16614 (N_16614,N_481,N_796);
nor U16615 (N_16615,N_357,N_4683);
nand U16616 (N_16616,N_327,N_1672);
or U16617 (N_16617,N_9423,N_6582);
nor U16618 (N_16618,N_9303,N_2018);
and U16619 (N_16619,N_2769,N_1746);
xor U16620 (N_16620,N_8645,N_1289);
nand U16621 (N_16621,N_5173,N_9106);
nand U16622 (N_16622,N_1527,N_2896);
and U16623 (N_16623,N_4607,N_1755);
and U16624 (N_16624,N_2296,N_8375);
and U16625 (N_16625,N_4732,N_7902);
and U16626 (N_16626,N_1727,N_6846);
nand U16627 (N_16627,N_6235,N_1903);
and U16628 (N_16628,N_6495,N_9081);
nor U16629 (N_16629,N_3526,N_8108);
and U16630 (N_16630,N_1059,N_5301);
xnor U16631 (N_16631,N_5868,N_8446);
and U16632 (N_16632,N_6058,N_2186);
and U16633 (N_16633,N_4999,N_138);
xnor U16634 (N_16634,N_437,N_9147);
nand U16635 (N_16635,N_6182,N_3238);
xnor U16636 (N_16636,N_5849,N_2569);
nor U16637 (N_16637,N_814,N_6239);
and U16638 (N_16638,N_8894,N_3784);
nand U16639 (N_16639,N_9768,N_7866);
nor U16640 (N_16640,N_7211,N_7482);
nand U16641 (N_16641,N_8688,N_6639);
nor U16642 (N_16642,N_9265,N_7021);
and U16643 (N_16643,N_4072,N_4623);
xnor U16644 (N_16644,N_1534,N_5382);
or U16645 (N_16645,N_2598,N_456);
nor U16646 (N_16646,N_996,N_7247);
nor U16647 (N_16647,N_221,N_9795);
or U16648 (N_16648,N_1422,N_7796);
and U16649 (N_16649,N_7439,N_3989);
nand U16650 (N_16650,N_9633,N_8326);
nand U16651 (N_16651,N_8513,N_6406);
nand U16652 (N_16652,N_8739,N_4154);
nand U16653 (N_16653,N_3745,N_6399);
nand U16654 (N_16654,N_2972,N_2730);
nor U16655 (N_16655,N_8060,N_9803);
nand U16656 (N_16656,N_7867,N_2171);
nand U16657 (N_16657,N_8321,N_8554);
nor U16658 (N_16658,N_4164,N_4701);
nand U16659 (N_16659,N_6355,N_9829);
or U16660 (N_16660,N_9405,N_1292);
or U16661 (N_16661,N_2097,N_8266);
and U16662 (N_16662,N_639,N_8788);
and U16663 (N_16663,N_4966,N_194);
xor U16664 (N_16664,N_7657,N_4210);
and U16665 (N_16665,N_9076,N_1293);
or U16666 (N_16666,N_6972,N_9595);
and U16667 (N_16667,N_6882,N_2507);
and U16668 (N_16668,N_5505,N_1716);
and U16669 (N_16669,N_723,N_7529);
or U16670 (N_16670,N_4640,N_4835);
xor U16671 (N_16671,N_3613,N_3991);
and U16672 (N_16672,N_3533,N_2992);
nand U16673 (N_16673,N_9856,N_4603);
nand U16674 (N_16674,N_4369,N_6784);
and U16675 (N_16675,N_7349,N_7123);
and U16676 (N_16676,N_287,N_4491);
xor U16677 (N_16677,N_4092,N_8708);
or U16678 (N_16678,N_9751,N_2691);
xor U16679 (N_16679,N_9935,N_4307);
xnor U16680 (N_16680,N_5357,N_7382);
nor U16681 (N_16681,N_9728,N_2700);
nor U16682 (N_16682,N_5601,N_705);
and U16683 (N_16683,N_3813,N_5897);
nor U16684 (N_16684,N_2148,N_6318);
xnor U16685 (N_16685,N_912,N_7430);
nor U16686 (N_16686,N_4310,N_2228);
nand U16687 (N_16687,N_4590,N_5541);
and U16688 (N_16688,N_8332,N_5363);
nor U16689 (N_16689,N_1767,N_9132);
xor U16690 (N_16690,N_1145,N_9516);
or U16691 (N_16691,N_4981,N_4613);
nor U16692 (N_16692,N_9762,N_776);
nand U16693 (N_16693,N_8983,N_4627);
nand U16694 (N_16694,N_4823,N_6846);
and U16695 (N_16695,N_2206,N_482);
nor U16696 (N_16696,N_7856,N_143);
nand U16697 (N_16697,N_5773,N_3617);
and U16698 (N_16698,N_7934,N_4188);
nor U16699 (N_16699,N_4797,N_2602);
and U16700 (N_16700,N_7782,N_6046);
or U16701 (N_16701,N_9925,N_6203);
or U16702 (N_16702,N_1450,N_2597);
and U16703 (N_16703,N_8134,N_9348);
or U16704 (N_16704,N_3172,N_6730);
or U16705 (N_16705,N_72,N_7674);
nor U16706 (N_16706,N_9075,N_911);
or U16707 (N_16707,N_6261,N_5275);
nand U16708 (N_16708,N_8868,N_2350);
nor U16709 (N_16709,N_9365,N_705);
nand U16710 (N_16710,N_2708,N_8485);
nand U16711 (N_16711,N_84,N_4340);
and U16712 (N_16712,N_949,N_9247);
or U16713 (N_16713,N_6378,N_6431);
and U16714 (N_16714,N_1378,N_8427);
nor U16715 (N_16715,N_758,N_8768);
nor U16716 (N_16716,N_7804,N_9526);
or U16717 (N_16717,N_416,N_7296);
nand U16718 (N_16718,N_2432,N_640);
or U16719 (N_16719,N_7571,N_628);
nand U16720 (N_16720,N_8332,N_8748);
or U16721 (N_16721,N_6132,N_4499);
nand U16722 (N_16722,N_5825,N_5169);
and U16723 (N_16723,N_567,N_4316);
and U16724 (N_16724,N_9130,N_2236);
nor U16725 (N_16725,N_9124,N_5312);
nor U16726 (N_16726,N_6136,N_7986);
nand U16727 (N_16727,N_5705,N_4487);
xor U16728 (N_16728,N_2554,N_2669);
nand U16729 (N_16729,N_4073,N_807);
xnor U16730 (N_16730,N_8954,N_4614);
nor U16731 (N_16731,N_5124,N_9551);
nor U16732 (N_16732,N_8301,N_3087);
nor U16733 (N_16733,N_6680,N_3400);
nand U16734 (N_16734,N_2944,N_4379);
nor U16735 (N_16735,N_8872,N_8533);
nand U16736 (N_16736,N_6501,N_9442);
and U16737 (N_16737,N_3762,N_3564);
nor U16738 (N_16738,N_976,N_6780);
nand U16739 (N_16739,N_867,N_2817);
or U16740 (N_16740,N_5932,N_7095);
or U16741 (N_16741,N_5204,N_8097);
and U16742 (N_16742,N_1327,N_3940);
and U16743 (N_16743,N_7892,N_8041);
nand U16744 (N_16744,N_4316,N_4542);
nand U16745 (N_16745,N_5656,N_691);
or U16746 (N_16746,N_1238,N_2312);
nand U16747 (N_16747,N_9011,N_3642);
or U16748 (N_16748,N_1440,N_3778);
or U16749 (N_16749,N_7947,N_7244);
nor U16750 (N_16750,N_237,N_2678);
or U16751 (N_16751,N_477,N_9343);
and U16752 (N_16752,N_6167,N_194);
or U16753 (N_16753,N_4631,N_5627);
xnor U16754 (N_16754,N_4417,N_7987);
nor U16755 (N_16755,N_109,N_3833);
nand U16756 (N_16756,N_8138,N_9666);
xor U16757 (N_16757,N_6087,N_7105);
nand U16758 (N_16758,N_229,N_1663);
nand U16759 (N_16759,N_3011,N_4540);
nand U16760 (N_16760,N_7072,N_5847);
and U16761 (N_16761,N_4008,N_4365);
nand U16762 (N_16762,N_9121,N_8891);
nor U16763 (N_16763,N_1028,N_8503);
or U16764 (N_16764,N_4103,N_8529);
nor U16765 (N_16765,N_5121,N_342);
nand U16766 (N_16766,N_4876,N_2435);
and U16767 (N_16767,N_7781,N_1559);
nor U16768 (N_16768,N_4215,N_5114);
nor U16769 (N_16769,N_8848,N_5608);
or U16770 (N_16770,N_3109,N_7166);
and U16771 (N_16771,N_4565,N_545);
and U16772 (N_16772,N_1668,N_1758);
and U16773 (N_16773,N_3328,N_5290);
or U16774 (N_16774,N_8571,N_7950);
nor U16775 (N_16775,N_7180,N_3613);
nor U16776 (N_16776,N_7338,N_7603);
nand U16777 (N_16777,N_9140,N_5514);
nor U16778 (N_16778,N_8897,N_3362);
or U16779 (N_16779,N_4296,N_2212);
nand U16780 (N_16780,N_3816,N_1250);
nor U16781 (N_16781,N_3178,N_9934);
nor U16782 (N_16782,N_6405,N_5849);
nand U16783 (N_16783,N_1027,N_6945);
nand U16784 (N_16784,N_3027,N_5645);
and U16785 (N_16785,N_9340,N_3575);
nand U16786 (N_16786,N_8402,N_9171);
and U16787 (N_16787,N_2195,N_4787);
and U16788 (N_16788,N_1379,N_4795);
nor U16789 (N_16789,N_9042,N_7107);
nor U16790 (N_16790,N_5708,N_4668);
and U16791 (N_16791,N_6992,N_2423);
nor U16792 (N_16792,N_2785,N_4805);
and U16793 (N_16793,N_9209,N_5781);
nand U16794 (N_16794,N_8691,N_2334);
nand U16795 (N_16795,N_1480,N_9727);
or U16796 (N_16796,N_4560,N_2383);
nor U16797 (N_16797,N_5134,N_3656);
and U16798 (N_16798,N_2649,N_6968);
and U16799 (N_16799,N_1363,N_4619);
nor U16800 (N_16800,N_1655,N_7057);
nand U16801 (N_16801,N_3396,N_7275);
nor U16802 (N_16802,N_8077,N_9249);
or U16803 (N_16803,N_7229,N_3102);
xnor U16804 (N_16804,N_3773,N_2544);
nor U16805 (N_16805,N_1068,N_6221);
or U16806 (N_16806,N_9408,N_9601);
or U16807 (N_16807,N_5148,N_1276);
or U16808 (N_16808,N_1491,N_910);
nor U16809 (N_16809,N_7958,N_8078);
nand U16810 (N_16810,N_7488,N_5010);
nor U16811 (N_16811,N_7513,N_6914);
or U16812 (N_16812,N_7750,N_3306);
nand U16813 (N_16813,N_1187,N_5627);
nor U16814 (N_16814,N_7869,N_2355);
and U16815 (N_16815,N_8519,N_6395);
or U16816 (N_16816,N_4159,N_7865);
nand U16817 (N_16817,N_9666,N_5553);
and U16818 (N_16818,N_9482,N_8625);
nor U16819 (N_16819,N_8434,N_1763);
and U16820 (N_16820,N_3721,N_133);
or U16821 (N_16821,N_151,N_2445);
nand U16822 (N_16822,N_30,N_5211);
nor U16823 (N_16823,N_5443,N_5077);
nor U16824 (N_16824,N_2949,N_6296);
nor U16825 (N_16825,N_4218,N_6405);
and U16826 (N_16826,N_7322,N_1345);
or U16827 (N_16827,N_3499,N_648);
and U16828 (N_16828,N_9907,N_5403);
nor U16829 (N_16829,N_4263,N_4827);
nor U16830 (N_16830,N_728,N_2433);
xor U16831 (N_16831,N_1443,N_432);
xnor U16832 (N_16832,N_5500,N_123);
and U16833 (N_16833,N_4870,N_2103);
nor U16834 (N_16834,N_3386,N_3119);
or U16835 (N_16835,N_6247,N_6925);
or U16836 (N_16836,N_1170,N_2568);
nor U16837 (N_16837,N_7168,N_5407);
or U16838 (N_16838,N_7423,N_266);
or U16839 (N_16839,N_2173,N_2189);
or U16840 (N_16840,N_4876,N_7407);
and U16841 (N_16841,N_4014,N_5260);
or U16842 (N_16842,N_1318,N_1664);
nor U16843 (N_16843,N_3921,N_6232);
nor U16844 (N_16844,N_2811,N_7657);
nand U16845 (N_16845,N_3224,N_4869);
or U16846 (N_16846,N_6743,N_8635);
nor U16847 (N_16847,N_9297,N_855);
nor U16848 (N_16848,N_4645,N_9827);
nand U16849 (N_16849,N_6727,N_2031);
nor U16850 (N_16850,N_1877,N_8159);
xnor U16851 (N_16851,N_7249,N_4126);
or U16852 (N_16852,N_7215,N_4436);
nand U16853 (N_16853,N_9527,N_9022);
xnor U16854 (N_16854,N_6219,N_7087);
xor U16855 (N_16855,N_9553,N_7205);
nor U16856 (N_16856,N_5704,N_8159);
xor U16857 (N_16857,N_4176,N_1115);
nor U16858 (N_16858,N_5438,N_7368);
and U16859 (N_16859,N_1230,N_8381);
and U16860 (N_16860,N_9409,N_2396);
xnor U16861 (N_16861,N_6833,N_9047);
or U16862 (N_16862,N_8074,N_2040);
nand U16863 (N_16863,N_8451,N_8283);
nand U16864 (N_16864,N_4331,N_188);
or U16865 (N_16865,N_2068,N_9650);
nand U16866 (N_16866,N_7711,N_8179);
xor U16867 (N_16867,N_4212,N_7641);
and U16868 (N_16868,N_3145,N_2770);
or U16869 (N_16869,N_4454,N_7067);
and U16870 (N_16870,N_9255,N_1665);
xor U16871 (N_16871,N_8698,N_8228);
or U16872 (N_16872,N_7089,N_9875);
nor U16873 (N_16873,N_664,N_7374);
xnor U16874 (N_16874,N_2963,N_6589);
nand U16875 (N_16875,N_3262,N_7431);
nand U16876 (N_16876,N_4013,N_7376);
nand U16877 (N_16877,N_9108,N_9689);
xnor U16878 (N_16878,N_1528,N_9870);
nand U16879 (N_16879,N_8587,N_3848);
xor U16880 (N_16880,N_138,N_3669);
nand U16881 (N_16881,N_8483,N_9293);
xnor U16882 (N_16882,N_6424,N_1808);
nand U16883 (N_16883,N_5986,N_683);
nand U16884 (N_16884,N_9810,N_5602);
nor U16885 (N_16885,N_3290,N_8626);
and U16886 (N_16886,N_7451,N_220);
and U16887 (N_16887,N_8355,N_7959);
nor U16888 (N_16888,N_2018,N_5201);
nor U16889 (N_16889,N_6773,N_1510);
nand U16890 (N_16890,N_9422,N_5027);
nor U16891 (N_16891,N_4355,N_768);
and U16892 (N_16892,N_7776,N_2650);
or U16893 (N_16893,N_1214,N_3660);
nor U16894 (N_16894,N_8657,N_5637);
nand U16895 (N_16895,N_1099,N_7237);
nand U16896 (N_16896,N_4863,N_9345);
nor U16897 (N_16897,N_7407,N_3660);
nand U16898 (N_16898,N_3506,N_4863);
or U16899 (N_16899,N_8588,N_7815);
or U16900 (N_16900,N_2960,N_7246);
or U16901 (N_16901,N_40,N_33);
and U16902 (N_16902,N_3069,N_9263);
nor U16903 (N_16903,N_3981,N_8973);
nand U16904 (N_16904,N_8599,N_3917);
and U16905 (N_16905,N_5704,N_8127);
or U16906 (N_16906,N_2860,N_8891);
nand U16907 (N_16907,N_9739,N_6432);
nand U16908 (N_16908,N_6265,N_4977);
or U16909 (N_16909,N_5547,N_2224);
and U16910 (N_16910,N_9458,N_1780);
and U16911 (N_16911,N_8805,N_4316);
or U16912 (N_16912,N_9420,N_2184);
nor U16913 (N_16913,N_1444,N_6041);
nor U16914 (N_16914,N_625,N_9287);
and U16915 (N_16915,N_5556,N_5965);
nand U16916 (N_16916,N_369,N_1558);
or U16917 (N_16917,N_8733,N_2306);
xor U16918 (N_16918,N_8333,N_4228);
or U16919 (N_16919,N_4395,N_2916);
nor U16920 (N_16920,N_5414,N_1681);
or U16921 (N_16921,N_2374,N_9185);
and U16922 (N_16922,N_9060,N_4445);
and U16923 (N_16923,N_970,N_160);
nor U16924 (N_16924,N_9404,N_4648);
nor U16925 (N_16925,N_5372,N_6476);
or U16926 (N_16926,N_6234,N_9433);
and U16927 (N_16927,N_7542,N_1023);
xnor U16928 (N_16928,N_5269,N_3831);
nor U16929 (N_16929,N_9334,N_3193);
nand U16930 (N_16930,N_4162,N_2089);
or U16931 (N_16931,N_1489,N_1703);
and U16932 (N_16932,N_7510,N_2380);
nor U16933 (N_16933,N_9729,N_4828);
and U16934 (N_16934,N_3366,N_7641);
xnor U16935 (N_16935,N_9264,N_8812);
and U16936 (N_16936,N_5545,N_9996);
nor U16937 (N_16937,N_4589,N_974);
nand U16938 (N_16938,N_8358,N_5267);
xnor U16939 (N_16939,N_5895,N_4388);
nor U16940 (N_16940,N_693,N_2328);
or U16941 (N_16941,N_1996,N_5170);
nor U16942 (N_16942,N_9410,N_6454);
xor U16943 (N_16943,N_3015,N_9133);
nor U16944 (N_16944,N_7985,N_3858);
nor U16945 (N_16945,N_9498,N_6761);
and U16946 (N_16946,N_3142,N_8227);
xor U16947 (N_16947,N_4697,N_3390);
xor U16948 (N_16948,N_9682,N_4616);
nor U16949 (N_16949,N_1825,N_6846);
or U16950 (N_16950,N_7604,N_7698);
nand U16951 (N_16951,N_7020,N_9294);
xor U16952 (N_16952,N_6664,N_1969);
or U16953 (N_16953,N_4647,N_6511);
or U16954 (N_16954,N_742,N_8958);
nor U16955 (N_16955,N_6907,N_1241);
or U16956 (N_16956,N_7963,N_8326);
or U16957 (N_16957,N_4982,N_3425);
nand U16958 (N_16958,N_5581,N_7638);
nor U16959 (N_16959,N_3728,N_5185);
nand U16960 (N_16960,N_7715,N_5747);
nand U16961 (N_16961,N_6240,N_7079);
and U16962 (N_16962,N_172,N_950);
nor U16963 (N_16963,N_2776,N_472);
and U16964 (N_16964,N_3064,N_7104);
nor U16965 (N_16965,N_4177,N_1131);
or U16966 (N_16966,N_2340,N_2450);
xor U16967 (N_16967,N_2863,N_1049);
nand U16968 (N_16968,N_5831,N_8742);
nand U16969 (N_16969,N_9764,N_6492);
xor U16970 (N_16970,N_8653,N_2889);
or U16971 (N_16971,N_139,N_3552);
xnor U16972 (N_16972,N_5143,N_4980);
nor U16973 (N_16973,N_8051,N_6948);
nand U16974 (N_16974,N_6425,N_2087);
xnor U16975 (N_16975,N_717,N_7506);
and U16976 (N_16976,N_5182,N_8832);
nor U16977 (N_16977,N_1407,N_8877);
and U16978 (N_16978,N_113,N_8785);
and U16979 (N_16979,N_9148,N_4983);
nor U16980 (N_16980,N_658,N_7711);
nor U16981 (N_16981,N_6261,N_9496);
and U16982 (N_16982,N_2833,N_3229);
nand U16983 (N_16983,N_9254,N_555);
nor U16984 (N_16984,N_3797,N_7344);
and U16985 (N_16985,N_5263,N_791);
nand U16986 (N_16986,N_1799,N_7781);
nand U16987 (N_16987,N_8995,N_9218);
nand U16988 (N_16988,N_4487,N_5794);
or U16989 (N_16989,N_3001,N_11);
and U16990 (N_16990,N_4639,N_7716);
nor U16991 (N_16991,N_6136,N_8179);
nand U16992 (N_16992,N_4355,N_6725);
xnor U16993 (N_16993,N_5900,N_5826);
and U16994 (N_16994,N_4036,N_5540);
nor U16995 (N_16995,N_6522,N_1722);
nand U16996 (N_16996,N_2642,N_3899);
or U16997 (N_16997,N_8968,N_6047);
nand U16998 (N_16998,N_5451,N_6359);
nand U16999 (N_16999,N_3469,N_7690);
nor U17000 (N_17000,N_8583,N_6528);
nor U17001 (N_17001,N_5674,N_7323);
or U17002 (N_17002,N_5102,N_1992);
nor U17003 (N_17003,N_8338,N_2086);
and U17004 (N_17004,N_5291,N_1174);
nor U17005 (N_17005,N_2586,N_4743);
or U17006 (N_17006,N_3208,N_8808);
and U17007 (N_17007,N_8010,N_3365);
xnor U17008 (N_17008,N_1350,N_2321);
nor U17009 (N_17009,N_6030,N_5763);
nand U17010 (N_17010,N_7563,N_305);
and U17011 (N_17011,N_9086,N_3678);
and U17012 (N_17012,N_408,N_2089);
or U17013 (N_17013,N_5841,N_980);
nor U17014 (N_17014,N_9467,N_9709);
and U17015 (N_17015,N_8293,N_7789);
and U17016 (N_17016,N_8198,N_2726);
or U17017 (N_17017,N_5788,N_2672);
or U17018 (N_17018,N_1687,N_6516);
nor U17019 (N_17019,N_5890,N_3852);
nor U17020 (N_17020,N_7250,N_6769);
and U17021 (N_17021,N_4678,N_584);
and U17022 (N_17022,N_2319,N_795);
nor U17023 (N_17023,N_5038,N_8680);
or U17024 (N_17024,N_8772,N_297);
nor U17025 (N_17025,N_3325,N_3526);
nor U17026 (N_17026,N_8040,N_5141);
and U17027 (N_17027,N_6132,N_7120);
xnor U17028 (N_17028,N_9812,N_9770);
and U17029 (N_17029,N_8259,N_3086);
nand U17030 (N_17030,N_4105,N_6776);
and U17031 (N_17031,N_9162,N_8071);
and U17032 (N_17032,N_7898,N_5985);
nor U17033 (N_17033,N_4296,N_1649);
or U17034 (N_17034,N_6375,N_198);
and U17035 (N_17035,N_6984,N_9683);
nor U17036 (N_17036,N_3598,N_2693);
nor U17037 (N_17037,N_5134,N_279);
nor U17038 (N_17038,N_6540,N_2382);
nor U17039 (N_17039,N_3206,N_5080);
nor U17040 (N_17040,N_6240,N_5869);
and U17041 (N_17041,N_6028,N_1027);
or U17042 (N_17042,N_951,N_4256);
nand U17043 (N_17043,N_940,N_2025);
or U17044 (N_17044,N_2742,N_1090);
nand U17045 (N_17045,N_5122,N_4444);
nor U17046 (N_17046,N_7552,N_4063);
or U17047 (N_17047,N_4034,N_4539);
xnor U17048 (N_17048,N_6032,N_1387);
nand U17049 (N_17049,N_9006,N_8660);
nor U17050 (N_17050,N_6849,N_7848);
nor U17051 (N_17051,N_7395,N_9928);
nand U17052 (N_17052,N_7075,N_8864);
xnor U17053 (N_17053,N_8333,N_8116);
nand U17054 (N_17054,N_598,N_314);
nor U17055 (N_17055,N_9200,N_7537);
nand U17056 (N_17056,N_5273,N_3059);
nand U17057 (N_17057,N_6712,N_8568);
and U17058 (N_17058,N_8284,N_5305);
nand U17059 (N_17059,N_6706,N_4691);
and U17060 (N_17060,N_4556,N_9205);
nor U17061 (N_17061,N_4514,N_39);
nand U17062 (N_17062,N_1716,N_4449);
nor U17063 (N_17063,N_349,N_6072);
or U17064 (N_17064,N_9589,N_6717);
nor U17065 (N_17065,N_903,N_3958);
xnor U17066 (N_17066,N_6126,N_4841);
and U17067 (N_17067,N_8810,N_8737);
nor U17068 (N_17068,N_6795,N_2137);
and U17069 (N_17069,N_2382,N_8504);
nor U17070 (N_17070,N_2756,N_5209);
or U17071 (N_17071,N_8296,N_3533);
xnor U17072 (N_17072,N_7473,N_5169);
or U17073 (N_17073,N_2994,N_611);
and U17074 (N_17074,N_9432,N_1370);
or U17075 (N_17075,N_3492,N_8181);
or U17076 (N_17076,N_7154,N_7934);
or U17077 (N_17077,N_127,N_2709);
nand U17078 (N_17078,N_7868,N_2554);
and U17079 (N_17079,N_416,N_6848);
and U17080 (N_17080,N_4011,N_8193);
or U17081 (N_17081,N_93,N_2943);
or U17082 (N_17082,N_8614,N_5048);
nand U17083 (N_17083,N_5586,N_1662);
and U17084 (N_17084,N_7592,N_1360);
nand U17085 (N_17085,N_2857,N_8720);
and U17086 (N_17086,N_652,N_7422);
and U17087 (N_17087,N_7484,N_6693);
nor U17088 (N_17088,N_4560,N_6780);
nand U17089 (N_17089,N_2519,N_9392);
or U17090 (N_17090,N_179,N_9052);
or U17091 (N_17091,N_8851,N_2946);
nand U17092 (N_17092,N_8788,N_2377);
xnor U17093 (N_17093,N_469,N_806);
and U17094 (N_17094,N_9857,N_9178);
or U17095 (N_17095,N_4561,N_1788);
nand U17096 (N_17096,N_5807,N_8710);
nand U17097 (N_17097,N_7004,N_6631);
nor U17098 (N_17098,N_5549,N_4069);
xor U17099 (N_17099,N_5514,N_496);
or U17100 (N_17100,N_2239,N_2156);
nand U17101 (N_17101,N_805,N_6086);
and U17102 (N_17102,N_5172,N_3032);
nor U17103 (N_17103,N_7527,N_132);
or U17104 (N_17104,N_4480,N_616);
nor U17105 (N_17105,N_7578,N_8144);
xor U17106 (N_17106,N_9196,N_3083);
nand U17107 (N_17107,N_6120,N_9600);
xor U17108 (N_17108,N_751,N_1467);
xor U17109 (N_17109,N_265,N_8617);
and U17110 (N_17110,N_51,N_1091);
nand U17111 (N_17111,N_518,N_8599);
xor U17112 (N_17112,N_7319,N_6974);
or U17113 (N_17113,N_2198,N_3258);
or U17114 (N_17114,N_1049,N_2542);
or U17115 (N_17115,N_5763,N_4070);
or U17116 (N_17116,N_1804,N_3444);
nor U17117 (N_17117,N_6978,N_7544);
nand U17118 (N_17118,N_8974,N_2030);
nand U17119 (N_17119,N_5391,N_5173);
nand U17120 (N_17120,N_1656,N_9280);
and U17121 (N_17121,N_825,N_6453);
or U17122 (N_17122,N_3453,N_5327);
and U17123 (N_17123,N_3924,N_3966);
nor U17124 (N_17124,N_5276,N_3267);
and U17125 (N_17125,N_2912,N_124);
nand U17126 (N_17126,N_4882,N_9997);
and U17127 (N_17127,N_5411,N_6775);
or U17128 (N_17128,N_9819,N_6404);
nor U17129 (N_17129,N_1896,N_4176);
or U17130 (N_17130,N_1796,N_3787);
or U17131 (N_17131,N_3639,N_2700);
and U17132 (N_17132,N_7950,N_8141);
nand U17133 (N_17133,N_6174,N_3524);
or U17134 (N_17134,N_297,N_4261);
nand U17135 (N_17135,N_7583,N_8117);
and U17136 (N_17136,N_4930,N_9663);
xor U17137 (N_17137,N_9961,N_322);
xnor U17138 (N_17138,N_1476,N_1673);
and U17139 (N_17139,N_8483,N_1226);
and U17140 (N_17140,N_3401,N_1321);
nand U17141 (N_17141,N_9602,N_1554);
nand U17142 (N_17142,N_234,N_3751);
or U17143 (N_17143,N_6792,N_1850);
and U17144 (N_17144,N_9381,N_8700);
nor U17145 (N_17145,N_1609,N_3869);
nor U17146 (N_17146,N_9187,N_5723);
and U17147 (N_17147,N_750,N_1696);
or U17148 (N_17148,N_4243,N_8608);
xnor U17149 (N_17149,N_4984,N_9553);
nor U17150 (N_17150,N_7187,N_8036);
nor U17151 (N_17151,N_1518,N_4677);
and U17152 (N_17152,N_6630,N_2004);
nor U17153 (N_17153,N_9314,N_2715);
nand U17154 (N_17154,N_5568,N_42);
and U17155 (N_17155,N_2074,N_6678);
and U17156 (N_17156,N_5718,N_4994);
or U17157 (N_17157,N_4885,N_379);
and U17158 (N_17158,N_8349,N_4958);
nor U17159 (N_17159,N_5304,N_177);
xnor U17160 (N_17160,N_2170,N_7871);
nand U17161 (N_17161,N_5211,N_5401);
or U17162 (N_17162,N_3925,N_5457);
nand U17163 (N_17163,N_6191,N_508);
and U17164 (N_17164,N_3263,N_6956);
and U17165 (N_17165,N_3252,N_5502);
nand U17166 (N_17166,N_1512,N_5107);
or U17167 (N_17167,N_796,N_2019);
and U17168 (N_17168,N_8098,N_654);
or U17169 (N_17169,N_9671,N_4406);
nand U17170 (N_17170,N_9786,N_2736);
and U17171 (N_17171,N_4754,N_9936);
nand U17172 (N_17172,N_3022,N_9655);
xor U17173 (N_17173,N_4357,N_8690);
or U17174 (N_17174,N_2642,N_9360);
nor U17175 (N_17175,N_9334,N_8866);
nor U17176 (N_17176,N_6840,N_3053);
or U17177 (N_17177,N_5047,N_7290);
xnor U17178 (N_17178,N_8601,N_815);
and U17179 (N_17179,N_5061,N_1135);
nor U17180 (N_17180,N_8816,N_1902);
or U17181 (N_17181,N_5200,N_9234);
or U17182 (N_17182,N_1712,N_7105);
or U17183 (N_17183,N_9208,N_6130);
nor U17184 (N_17184,N_7479,N_1157);
xor U17185 (N_17185,N_4966,N_6916);
or U17186 (N_17186,N_3574,N_2966);
or U17187 (N_17187,N_6320,N_7895);
nand U17188 (N_17188,N_7529,N_4154);
or U17189 (N_17189,N_3962,N_2049);
nand U17190 (N_17190,N_9720,N_1146);
nand U17191 (N_17191,N_4570,N_2355);
nand U17192 (N_17192,N_9630,N_7290);
nor U17193 (N_17193,N_2969,N_992);
nand U17194 (N_17194,N_6233,N_3650);
and U17195 (N_17195,N_2046,N_349);
nor U17196 (N_17196,N_3595,N_9162);
or U17197 (N_17197,N_7096,N_3931);
nor U17198 (N_17198,N_8986,N_8227);
nor U17199 (N_17199,N_4507,N_3650);
xnor U17200 (N_17200,N_5628,N_6852);
and U17201 (N_17201,N_4026,N_4184);
or U17202 (N_17202,N_4247,N_3988);
and U17203 (N_17203,N_6178,N_6399);
or U17204 (N_17204,N_7413,N_1069);
and U17205 (N_17205,N_8658,N_4526);
nand U17206 (N_17206,N_9178,N_72);
or U17207 (N_17207,N_9298,N_799);
and U17208 (N_17208,N_9597,N_1197);
nor U17209 (N_17209,N_2792,N_723);
xnor U17210 (N_17210,N_1715,N_615);
nand U17211 (N_17211,N_7658,N_7627);
nor U17212 (N_17212,N_4539,N_3421);
or U17213 (N_17213,N_5821,N_1328);
nand U17214 (N_17214,N_5346,N_3607);
and U17215 (N_17215,N_3993,N_6422);
or U17216 (N_17216,N_3931,N_6660);
and U17217 (N_17217,N_180,N_2349);
nand U17218 (N_17218,N_7631,N_6143);
nand U17219 (N_17219,N_2459,N_4992);
nor U17220 (N_17220,N_4216,N_9403);
and U17221 (N_17221,N_8974,N_3189);
or U17222 (N_17222,N_6210,N_8289);
nand U17223 (N_17223,N_5628,N_9431);
xor U17224 (N_17224,N_3741,N_5889);
and U17225 (N_17225,N_7112,N_8628);
or U17226 (N_17226,N_9893,N_7224);
nor U17227 (N_17227,N_3715,N_25);
and U17228 (N_17228,N_7997,N_5555);
or U17229 (N_17229,N_7936,N_4886);
nand U17230 (N_17230,N_8794,N_9273);
or U17231 (N_17231,N_6344,N_3736);
nor U17232 (N_17232,N_2579,N_6740);
nor U17233 (N_17233,N_1247,N_1363);
nand U17234 (N_17234,N_3024,N_7221);
and U17235 (N_17235,N_5233,N_5492);
nand U17236 (N_17236,N_7634,N_6503);
xor U17237 (N_17237,N_4254,N_5271);
nor U17238 (N_17238,N_3860,N_3388);
xor U17239 (N_17239,N_1125,N_2150);
or U17240 (N_17240,N_1303,N_3499);
nor U17241 (N_17241,N_1609,N_5701);
and U17242 (N_17242,N_6319,N_9651);
or U17243 (N_17243,N_6964,N_4091);
and U17244 (N_17244,N_6186,N_8465);
or U17245 (N_17245,N_1709,N_1569);
or U17246 (N_17246,N_2287,N_5072);
or U17247 (N_17247,N_4559,N_5095);
and U17248 (N_17248,N_9063,N_2552);
or U17249 (N_17249,N_381,N_6810);
and U17250 (N_17250,N_4566,N_9079);
and U17251 (N_17251,N_5285,N_9841);
xor U17252 (N_17252,N_2422,N_7327);
nand U17253 (N_17253,N_400,N_6122);
or U17254 (N_17254,N_1732,N_4748);
and U17255 (N_17255,N_1056,N_7609);
nand U17256 (N_17256,N_7694,N_4905);
nor U17257 (N_17257,N_149,N_4649);
and U17258 (N_17258,N_4174,N_2905);
nand U17259 (N_17259,N_946,N_5115);
and U17260 (N_17260,N_2142,N_844);
nor U17261 (N_17261,N_7135,N_1173);
nor U17262 (N_17262,N_1138,N_9909);
nor U17263 (N_17263,N_1579,N_1742);
nand U17264 (N_17264,N_5514,N_4124);
or U17265 (N_17265,N_3572,N_6601);
or U17266 (N_17266,N_5944,N_8851);
nor U17267 (N_17267,N_9905,N_9500);
xor U17268 (N_17268,N_8777,N_6440);
or U17269 (N_17269,N_6829,N_8359);
xor U17270 (N_17270,N_8999,N_6805);
xor U17271 (N_17271,N_6223,N_9887);
xor U17272 (N_17272,N_7161,N_8616);
xor U17273 (N_17273,N_5596,N_5650);
and U17274 (N_17274,N_9249,N_2314);
nand U17275 (N_17275,N_7580,N_8203);
and U17276 (N_17276,N_6611,N_2328);
or U17277 (N_17277,N_1530,N_2619);
or U17278 (N_17278,N_7578,N_2278);
nor U17279 (N_17279,N_5564,N_2800);
and U17280 (N_17280,N_4650,N_8752);
xnor U17281 (N_17281,N_1629,N_1730);
nand U17282 (N_17282,N_3156,N_666);
or U17283 (N_17283,N_9575,N_2492);
or U17284 (N_17284,N_6836,N_2490);
or U17285 (N_17285,N_1694,N_3163);
xor U17286 (N_17286,N_6219,N_9012);
nor U17287 (N_17287,N_2815,N_9095);
and U17288 (N_17288,N_7022,N_9189);
xnor U17289 (N_17289,N_7077,N_5850);
nor U17290 (N_17290,N_6003,N_6393);
nor U17291 (N_17291,N_5050,N_1716);
nor U17292 (N_17292,N_4240,N_4968);
nand U17293 (N_17293,N_1642,N_7161);
or U17294 (N_17294,N_6027,N_4953);
and U17295 (N_17295,N_4027,N_1361);
nand U17296 (N_17296,N_2921,N_585);
or U17297 (N_17297,N_3209,N_7422);
or U17298 (N_17298,N_157,N_8341);
nand U17299 (N_17299,N_5499,N_6415);
or U17300 (N_17300,N_3837,N_4382);
nand U17301 (N_17301,N_9595,N_9574);
nand U17302 (N_17302,N_2468,N_6490);
and U17303 (N_17303,N_7189,N_9035);
or U17304 (N_17304,N_4186,N_713);
or U17305 (N_17305,N_6763,N_2852);
and U17306 (N_17306,N_2895,N_8681);
or U17307 (N_17307,N_8331,N_7878);
or U17308 (N_17308,N_1617,N_4800);
and U17309 (N_17309,N_7285,N_1503);
nor U17310 (N_17310,N_4029,N_4425);
and U17311 (N_17311,N_4338,N_8138);
or U17312 (N_17312,N_1559,N_7149);
nand U17313 (N_17313,N_6902,N_4006);
or U17314 (N_17314,N_402,N_4307);
xor U17315 (N_17315,N_8993,N_3184);
xnor U17316 (N_17316,N_8726,N_7058);
xnor U17317 (N_17317,N_6805,N_4514);
nor U17318 (N_17318,N_5270,N_1695);
nor U17319 (N_17319,N_6715,N_5337);
nor U17320 (N_17320,N_589,N_4432);
xor U17321 (N_17321,N_6715,N_5430);
nand U17322 (N_17322,N_692,N_4576);
nand U17323 (N_17323,N_7839,N_3298);
xor U17324 (N_17324,N_5857,N_9220);
nand U17325 (N_17325,N_1833,N_108);
or U17326 (N_17326,N_9773,N_1993);
nor U17327 (N_17327,N_5182,N_4596);
nand U17328 (N_17328,N_2178,N_3652);
nor U17329 (N_17329,N_2460,N_5067);
nand U17330 (N_17330,N_1028,N_5414);
and U17331 (N_17331,N_6702,N_4253);
nor U17332 (N_17332,N_8547,N_5071);
or U17333 (N_17333,N_5227,N_7753);
or U17334 (N_17334,N_4685,N_1937);
and U17335 (N_17335,N_5142,N_8436);
xnor U17336 (N_17336,N_2645,N_4365);
nor U17337 (N_17337,N_6884,N_931);
and U17338 (N_17338,N_6132,N_9722);
nand U17339 (N_17339,N_4645,N_8699);
nand U17340 (N_17340,N_9389,N_4867);
xor U17341 (N_17341,N_6310,N_2843);
or U17342 (N_17342,N_5415,N_6465);
or U17343 (N_17343,N_8301,N_427);
nand U17344 (N_17344,N_7907,N_3319);
or U17345 (N_17345,N_2011,N_4438);
or U17346 (N_17346,N_2293,N_2097);
or U17347 (N_17347,N_7466,N_3624);
nor U17348 (N_17348,N_8466,N_5524);
nor U17349 (N_17349,N_6755,N_1734);
nor U17350 (N_17350,N_270,N_5338);
nor U17351 (N_17351,N_6758,N_2261);
nor U17352 (N_17352,N_3890,N_3130);
nand U17353 (N_17353,N_3252,N_8938);
xor U17354 (N_17354,N_4928,N_2944);
or U17355 (N_17355,N_7096,N_803);
nor U17356 (N_17356,N_8609,N_2608);
and U17357 (N_17357,N_6765,N_7464);
or U17358 (N_17358,N_8048,N_8655);
nand U17359 (N_17359,N_8524,N_9218);
nor U17360 (N_17360,N_6835,N_4891);
nand U17361 (N_17361,N_4884,N_8729);
xnor U17362 (N_17362,N_1477,N_1595);
nand U17363 (N_17363,N_9397,N_8962);
or U17364 (N_17364,N_3650,N_72);
nand U17365 (N_17365,N_5773,N_6728);
nor U17366 (N_17366,N_6210,N_786);
or U17367 (N_17367,N_8985,N_5796);
or U17368 (N_17368,N_5888,N_7632);
nor U17369 (N_17369,N_8248,N_3452);
nand U17370 (N_17370,N_8408,N_107);
and U17371 (N_17371,N_2180,N_3392);
nor U17372 (N_17372,N_6485,N_2472);
or U17373 (N_17373,N_3741,N_2479);
or U17374 (N_17374,N_1138,N_885);
or U17375 (N_17375,N_800,N_3129);
or U17376 (N_17376,N_8371,N_3786);
nor U17377 (N_17377,N_8314,N_677);
or U17378 (N_17378,N_1379,N_6914);
and U17379 (N_17379,N_2745,N_9271);
nand U17380 (N_17380,N_965,N_4225);
or U17381 (N_17381,N_9584,N_3511);
nand U17382 (N_17382,N_8533,N_129);
or U17383 (N_17383,N_3089,N_8082);
or U17384 (N_17384,N_4994,N_3074);
and U17385 (N_17385,N_7306,N_4725);
nand U17386 (N_17386,N_2389,N_3679);
or U17387 (N_17387,N_220,N_5759);
nor U17388 (N_17388,N_9783,N_3353);
xor U17389 (N_17389,N_6411,N_2597);
or U17390 (N_17390,N_3858,N_8392);
or U17391 (N_17391,N_2011,N_1040);
xnor U17392 (N_17392,N_6387,N_5767);
nand U17393 (N_17393,N_4751,N_4887);
and U17394 (N_17394,N_3677,N_1701);
or U17395 (N_17395,N_1025,N_2002);
nand U17396 (N_17396,N_4556,N_5521);
or U17397 (N_17397,N_2384,N_5844);
xor U17398 (N_17398,N_4899,N_9532);
nand U17399 (N_17399,N_1609,N_3057);
xnor U17400 (N_17400,N_4444,N_2259);
or U17401 (N_17401,N_2883,N_9134);
nor U17402 (N_17402,N_9557,N_6297);
or U17403 (N_17403,N_1309,N_2693);
nor U17404 (N_17404,N_7620,N_6943);
or U17405 (N_17405,N_3615,N_8253);
or U17406 (N_17406,N_8186,N_1166);
and U17407 (N_17407,N_7473,N_6502);
xor U17408 (N_17408,N_315,N_3132);
or U17409 (N_17409,N_7455,N_7880);
nand U17410 (N_17410,N_485,N_9818);
nand U17411 (N_17411,N_4210,N_4378);
and U17412 (N_17412,N_1100,N_1970);
and U17413 (N_17413,N_6626,N_5217);
and U17414 (N_17414,N_8217,N_7168);
nand U17415 (N_17415,N_8974,N_9102);
and U17416 (N_17416,N_320,N_2228);
nor U17417 (N_17417,N_169,N_7632);
nor U17418 (N_17418,N_2178,N_6026);
or U17419 (N_17419,N_6406,N_2654);
nor U17420 (N_17420,N_4565,N_6480);
nor U17421 (N_17421,N_3863,N_7920);
and U17422 (N_17422,N_5661,N_4567);
and U17423 (N_17423,N_4646,N_6694);
nand U17424 (N_17424,N_1366,N_1828);
nor U17425 (N_17425,N_4953,N_5329);
and U17426 (N_17426,N_7721,N_1530);
nor U17427 (N_17427,N_29,N_6278);
nor U17428 (N_17428,N_9289,N_6525);
and U17429 (N_17429,N_7800,N_8971);
nand U17430 (N_17430,N_1794,N_7449);
and U17431 (N_17431,N_7306,N_5236);
or U17432 (N_17432,N_1979,N_9258);
nand U17433 (N_17433,N_8464,N_9547);
nor U17434 (N_17434,N_7151,N_3026);
nand U17435 (N_17435,N_9679,N_7222);
and U17436 (N_17436,N_9262,N_7396);
nor U17437 (N_17437,N_2685,N_4649);
and U17438 (N_17438,N_9988,N_7023);
or U17439 (N_17439,N_2562,N_2836);
nand U17440 (N_17440,N_7437,N_6512);
xor U17441 (N_17441,N_6845,N_337);
nor U17442 (N_17442,N_929,N_2346);
nor U17443 (N_17443,N_6676,N_2445);
nor U17444 (N_17444,N_6310,N_6279);
nand U17445 (N_17445,N_1430,N_8083);
nand U17446 (N_17446,N_5200,N_8797);
nor U17447 (N_17447,N_4487,N_1974);
nand U17448 (N_17448,N_3568,N_5843);
or U17449 (N_17449,N_4676,N_7636);
nor U17450 (N_17450,N_4575,N_297);
nor U17451 (N_17451,N_7146,N_5684);
and U17452 (N_17452,N_9711,N_9259);
nand U17453 (N_17453,N_3073,N_960);
or U17454 (N_17454,N_6735,N_4089);
xor U17455 (N_17455,N_288,N_9552);
nand U17456 (N_17456,N_4720,N_4742);
or U17457 (N_17457,N_9293,N_825);
nand U17458 (N_17458,N_3702,N_623);
xor U17459 (N_17459,N_8320,N_6408);
xor U17460 (N_17460,N_8595,N_999);
nand U17461 (N_17461,N_1692,N_4318);
and U17462 (N_17462,N_9064,N_8110);
and U17463 (N_17463,N_8432,N_5276);
or U17464 (N_17464,N_4245,N_1249);
nor U17465 (N_17465,N_1064,N_8137);
nor U17466 (N_17466,N_4084,N_2542);
nand U17467 (N_17467,N_787,N_6041);
and U17468 (N_17468,N_9646,N_8742);
and U17469 (N_17469,N_6136,N_7885);
or U17470 (N_17470,N_3284,N_4607);
or U17471 (N_17471,N_6480,N_6073);
or U17472 (N_17472,N_8130,N_555);
nor U17473 (N_17473,N_2353,N_4243);
nand U17474 (N_17474,N_6925,N_2186);
or U17475 (N_17475,N_496,N_7650);
nor U17476 (N_17476,N_4357,N_6647);
and U17477 (N_17477,N_7039,N_9947);
and U17478 (N_17478,N_4372,N_8194);
xor U17479 (N_17479,N_6712,N_4474);
nor U17480 (N_17480,N_9231,N_9860);
or U17481 (N_17481,N_9724,N_2574);
and U17482 (N_17482,N_703,N_8541);
nor U17483 (N_17483,N_118,N_7206);
xor U17484 (N_17484,N_4452,N_8311);
and U17485 (N_17485,N_6376,N_2493);
and U17486 (N_17486,N_2534,N_7032);
nand U17487 (N_17487,N_2954,N_6529);
xnor U17488 (N_17488,N_9382,N_9307);
nor U17489 (N_17489,N_8797,N_9590);
nand U17490 (N_17490,N_5308,N_2955);
nor U17491 (N_17491,N_5034,N_360);
and U17492 (N_17492,N_4453,N_7609);
nor U17493 (N_17493,N_1946,N_5435);
nand U17494 (N_17494,N_4915,N_5404);
xor U17495 (N_17495,N_9843,N_8707);
or U17496 (N_17496,N_920,N_1962);
nor U17497 (N_17497,N_9329,N_6628);
xor U17498 (N_17498,N_9434,N_443);
nor U17499 (N_17499,N_9993,N_5878);
nand U17500 (N_17500,N_761,N_2181);
or U17501 (N_17501,N_3803,N_3673);
xor U17502 (N_17502,N_6496,N_2744);
nor U17503 (N_17503,N_5903,N_7476);
nor U17504 (N_17504,N_9650,N_3714);
nor U17505 (N_17505,N_6452,N_3611);
nor U17506 (N_17506,N_2144,N_7697);
or U17507 (N_17507,N_3141,N_5092);
and U17508 (N_17508,N_3443,N_8014);
and U17509 (N_17509,N_3822,N_2762);
and U17510 (N_17510,N_7627,N_9468);
nor U17511 (N_17511,N_1313,N_6743);
and U17512 (N_17512,N_5141,N_9598);
nor U17513 (N_17513,N_3705,N_5746);
and U17514 (N_17514,N_5977,N_8426);
xor U17515 (N_17515,N_7354,N_1076);
nor U17516 (N_17516,N_3172,N_6611);
xnor U17517 (N_17517,N_4586,N_8888);
nor U17518 (N_17518,N_536,N_5329);
and U17519 (N_17519,N_2642,N_1136);
xor U17520 (N_17520,N_9473,N_5035);
or U17521 (N_17521,N_1912,N_509);
or U17522 (N_17522,N_4644,N_1338);
xor U17523 (N_17523,N_6960,N_603);
nor U17524 (N_17524,N_7667,N_3624);
or U17525 (N_17525,N_1447,N_9584);
nor U17526 (N_17526,N_9185,N_9944);
and U17527 (N_17527,N_2169,N_4782);
and U17528 (N_17528,N_3889,N_566);
nand U17529 (N_17529,N_4324,N_6078);
nor U17530 (N_17530,N_2646,N_6397);
or U17531 (N_17531,N_1066,N_9771);
and U17532 (N_17532,N_8872,N_8625);
nand U17533 (N_17533,N_5056,N_3241);
or U17534 (N_17534,N_3244,N_6445);
nor U17535 (N_17535,N_9963,N_5281);
nor U17536 (N_17536,N_5500,N_2869);
xnor U17537 (N_17537,N_2369,N_2816);
nand U17538 (N_17538,N_7593,N_2098);
xor U17539 (N_17539,N_2135,N_1);
nor U17540 (N_17540,N_5573,N_4385);
nor U17541 (N_17541,N_5058,N_5640);
and U17542 (N_17542,N_5032,N_8818);
xnor U17543 (N_17543,N_532,N_5619);
nor U17544 (N_17544,N_5987,N_3782);
nand U17545 (N_17545,N_4390,N_4590);
nor U17546 (N_17546,N_8684,N_6983);
nor U17547 (N_17547,N_8257,N_7354);
or U17548 (N_17548,N_6401,N_3919);
nand U17549 (N_17549,N_7959,N_2398);
nor U17550 (N_17550,N_9843,N_9176);
or U17551 (N_17551,N_7762,N_2873);
or U17552 (N_17552,N_6121,N_6091);
nand U17553 (N_17553,N_1642,N_1373);
nor U17554 (N_17554,N_5409,N_3489);
nor U17555 (N_17555,N_969,N_3118);
or U17556 (N_17556,N_5738,N_7268);
xnor U17557 (N_17557,N_376,N_9844);
nand U17558 (N_17558,N_1049,N_6924);
nor U17559 (N_17559,N_4649,N_435);
and U17560 (N_17560,N_7437,N_7399);
nor U17561 (N_17561,N_3052,N_3851);
or U17562 (N_17562,N_5059,N_9806);
xor U17563 (N_17563,N_7355,N_5800);
nand U17564 (N_17564,N_2947,N_9672);
or U17565 (N_17565,N_4169,N_6807);
nand U17566 (N_17566,N_9484,N_3421);
or U17567 (N_17567,N_5088,N_9467);
and U17568 (N_17568,N_3224,N_24);
and U17569 (N_17569,N_6671,N_3564);
or U17570 (N_17570,N_6704,N_5842);
nand U17571 (N_17571,N_6159,N_9040);
nor U17572 (N_17572,N_461,N_4602);
nand U17573 (N_17573,N_9786,N_5070);
nor U17574 (N_17574,N_2321,N_2181);
and U17575 (N_17575,N_2711,N_7222);
and U17576 (N_17576,N_2235,N_883);
or U17577 (N_17577,N_8073,N_6249);
xnor U17578 (N_17578,N_3421,N_229);
or U17579 (N_17579,N_6747,N_2477);
nor U17580 (N_17580,N_1431,N_7446);
nand U17581 (N_17581,N_7776,N_4206);
or U17582 (N_17582,N_1835,N_6689);
xor U17583 (N_17583,N_2854,N_895);
nand U17584 (N_17584,N_4594,N_4291);
or U17585 (N_17585,N_9818,N_716);
or U17586 (N_17586,N_5450,N_2426);
or U17587 (N_17587,N_5253,N_6173);
nand U17588 (N_17588,N_2240,N_2595);
nand U17589 (N_17589,N_3086,N_5696);
nand U17590 (N_17590,N_4179,N_3178);
and U17591 (N_17591,N_4637,N_6009);
nor U17592 (N_17592,N_3255,N_81);
nor U17593 (N_17593,N_3401,N_1677);
nand U17594 (N_17594,N_227,N_4847);
nand U17595 (N_17595,N_4685,N_9496);
and U17596 (N_17596,N_5049,N_1537);
nand U17597 (N_17597,N_5781,N_7969);
or U17598 (N_17598,N_5003,N_4229);
nor U17599 (N_17599,N_6080,N_2963);
or U17600 (N_17600,N_5110,N_5695);
nor U17601 (N_17601,N_4954,N_9724);
nand U17602 (N_17602,N_7239,N_5290);
xnor U17603 (N_17603,N_2532,N_4079);
and U17604 (N_17604,N_4635,N_7352);
nor U17605 (N_17605,N_2940,N_7802);
or U17606 (N_17606,N_3627,N_251);
and U17607 (N_17607,N_2666,N_5699);
or U17608 (N_17608,N_6740,N_8337);
and U17609 (N_17609,N_7013,N_6529);
nand U17610 (N_17610,N_3043,N_5256);
nand U17611 (N_17611,N_784,N_3107);
and U17612 (N_17612,N_3601,N_6550);
nor U17613 (N_17613,N_9993,N_5705);
nor U17614 (N_17614,N_4216,N_5609);
and U17615 (N_17615,N_8627,N_3030);
nand U17616 (N_17616,N_5465,N_1618);
nand U17617 (N_17617,N_2097,N_2555);
nor U17618 (N_17618,N_5655,N_1608);
nand U17619 (N_17619,N_4369,N_543);
nand U17620 (N_17620,N_2688,N_804);
nor U17621 (N_17621,N_6830,N_1873);
or U17622 (N_17622,N_1924,N_5025);
and U17623 (N_17623,N_1961,N_1317);
nand U17624 (N_17624,N_8,N_3592);
or U17625 (N_17625,N_7121,N_5587);
or U17626 (N_17626,N_2851,N_8022);
or U17627 (N_17627,N_6051,N_9903);
or U17628 (N_17628,N_7424,N_7480);
nand U17629 (N_17629,N_1250,N_9612);
xor U17630 (N_17630,N_7310,N_2887);
or U17631 (N_17631,N_137,N_6576);
and U17632 (N_17632,N_1630,N_7887);
nor U17633 (N_17633,N_3322,N_4566);
nand U17634 (N_17634,N_2379,N_160);
and U17635 (N_17635,N_4947,N_4334);
xor U17636 (N_17636,N_6676,N_9497);
or U17637 (N_17637,N_6780,N_475);
nor U17638 (N_17638,N_990,N_9577);
or U17639 (N_17639,N_3385,N_8607);
nand U17640 (N_17640,N_4576,N_1070);
nand U17641 (N_17641,N_4893,N_2650);
nor U17642 (N_17642,N_4181,N_6149);
nand U17643 (N_17643,N_8600,N_5139);
or U17644 (N_17644,N_8074,N_1546);
nor U17645 (N_17645,N_3702,N_4815);
nand U17646 (N_17646,N_5290,N_917);
nor U17647 (N_17647,N_4132,N_6242);
nand U17648 (N_17648,N_7524,N_5411);
xnor U17649 (N_17649,N_8557,N_5570);
xor U17650 (N_17650,N_6749,N_7420);
and U17651 (N_17651,N_9369,N_8506);
and U17652 (N_17652,N_3532,N_1550);
or U17653 (N_17653,N_4819,N_4407);
xnor U17654 (N_17654,N_2112,N_8423);
or U17655 (N_17655,N_928,N_5529);
xor U17656 (N_17656,N_8503,N_2941);
nand U17657 (N_17657,N_1375,N_626);
xnor U17658 (N_17658,N_2299,N_5322);
nand U17659 (N_17659,N_9596,N_4227);
nand U17660 (N_17660,N_492,N_5712);
xor U17661 (N_17661,N_3640,N_2699);
and U17662 (N_17662,N_5091,N_5585);
or U17663 (N_17663,N_1418,N_8478);
and U17664 (N_17664,N_3653,N_9404);
or U17665 (N_17665,N_6707,N_5871);
nor U17666 (N_17666,N_6383,N_3447);
and U17667 (N_17667,N_8015,N_1310);
and U17668 (N_17668,N_5442,N_5007);
or U17669 (N_17669,N_6129,N_6785);
nor U17670 (N_17670,N_3119,N_5775);
or U17671 (N_17671,N_7134,N_6144);
nor U17672 (N_17672,N_9583,N_2747);
nand U17673 (N_17673,N_5312,N_6761);
nor U17674 (N_17674,N_3848,N_5835);
xor U17675 (N_17675,N_2856,N_971);
nor U17676 (N_17676,N_5300,N_2802);
or U17677 (N_17677,N_4450,N_8985);
nor U17678 (N_17678,N_9317,N_3816);
nor U17679 (N_17679,N_1866,N_7759);
nor U17680 (N_17680,N_4956,N_7245);
xnor U17681 (N_17681,N_4050,N_4696);
and U17682 (N_17682,N_1092,N_8272);
and U17683 (N_17683,N_1823,N_6291);
and U17684 (N_17684,N_4024,N_3341);
nand U17685 (N_17685,N_5391,N_6097);
nand U17686 (N_17686,N_6487,N_1208);
and U17687 (N_17687,N_4947,N_8300);
nor U17688 (N_17688,N_5874,N_951);
or U17689 (N_17689,N_2989,N_9688);
or U17690 (N_17690,N_3904,N_2617);
nor U17691 (N_17691,N_3122,N_8575);
or U17692 (N_17692,N_3758,N_8531);
or U17693 (N_17693,N_4656,N_8877);
nor U17694 (N_17694,N_9997,N_3522);
and U17695 (N_17695,N_5092,N_3735);
nand U17696 (N_17696,N_4741,N_8232);
nand U17697 (N_17697,N_8527,N_2400);
xnor U17698 (N_17698,N_6299,N_4484);
and U17699 (N_17699,N_3352,N_1495);
and U17700 (N_17700,N_951,N_1525);
or U17701 (N_17701,N_6472,N_513);
nor U17702 (N_17702,N_7407,N_9925);
or U17703 (N_17703,N_9986,N_6301);
nand U17704 (N_17704,N_8462,N_7076);
nand U17705 (N_17705,N_4141,N_7432);
and U17706 (N_17706,N_3583,N_4539);
nand U17707 (N_17707,N_5475,N_5694);
or U17708 (N_17708,N_3134,N_9065);
xnor U17709 (N_17709,N_1336,N_7585);
nor U17710 (N_17710,N_1379,N_5751);
and U17711 (N_17711,N_8595,N_4164);
and U17712 (N_17712,N_879,N_2319);
and U17713 (N_17713,N_9609,N_9280);
nor U17714 (N_17714,N_7217,N_9056);
nand U17715 (N_17715,N_483,N_2719);
xnor U17716 (N_17716,N_6037,N_2186);
nor U17717 (N_17717,N_5343,N_2939);
and U17718 (N_17718,N_3674,N_1974);
nand U17719 (N_17719,N_6986,N_7727);
nor U17720 (N_17720,N_5768,N_4717);
nand U17721 (N_17721,N_5859,N_3331);
nor U17722 (N_17722,N_6579,N_2053);
and U17723 (N_17723,N_4712,N_9201);
nand U17724 (N_17724,N_5652,N_5383);
nand U17725 (N_17725,N_6188,N_6346);
nor U17726 (N_17726,N_3509,N_5302);
and U17727 (N_17727,N_309,N_8971);
and U17728 (N_17728,N_5927,N_255);
or U17729 (N_17729,N_7612,N_2328);
nor U17730 (N_17730,N_688,N_7739);
and U17731 (N_17731,N_9129,N_7292);
nand U17732 (N_17732,N_6049,N_7011);
nand U17733 (N_17733,N_6032,N_9981);
and U17734 (N_17734,N_2488,N_5605);
nand U17735 (N_17735,N_9195,N_597);
nor U17736 (N_17736,N_4766,N_7745);
nand U17737 (N_17737,N_7508,N_6459);
and U17738 (N_17738,N_3225,N_8317);
and U17739 (N_17739,N_5840,N_818);
or U17740 (N_17740,N_2424,N_2297);
nor U17741 (N_17741,N_4650,N_2426);
and U17742 (N_17742,N_6870,N_4491);
and U17743 (N_17743,N_9234,N_7550);
and U17744 (N_17744,N_2859,N_5535);
or U17745 (N_17745,N_4928,N_4147);
xnor U17746 (N_17746,N_9704,N_5311);
or U17747 (N_17747,N_8857,N_7666);
or U17748 (N_17748,N_656,N_6227);
xnor U17749 (N_17749,N_9873,N_2885);
xor U17750 (N_17750,N_5422,N_9118);
nor U17751 (N_17751,N_2752,N_726);
nor U17752 (N_17752,N_18,N_3598);
nand U17753 (N_17753,N_6863,N_5122);
or U17754 (N_17754,N_2031,N_9139);
nor U17755 (N_17755,N_8743,N_1987);
nor U17756 (N_17756,N_434,N_5585);
nand U17757 (N_17757,N_5209,N_4552);
nor U17758 (N_17758,N_187,N_6790);
or U17759 (N_17759,N_2953,N_4090);
or U17760 (N_17760,N_361,N_7095);
nor U17761 (N_17761,N_6869,N_4080);
nand U17762 (N_17762,N_9279,N_5030);
nor U17763 (N_17763,N_2544,N_8664);
and U17764 (N_17764,N_410,N_9948);
nor U17765 (N_17765,N_1153,N_8127);
nand U17766 (N_17766,N_3276,N_8518);
nand U17767 (N_17767,N_8756,N_7406);
nor U17768 (N_17768,N_8477,N_6292);
or U17769 (N_17769,N_8879,N_2233);
and U17770 (N_17770,N_6762,N_9412);
xor U17771 (N_17771,N_3584,N_7677);
nor U17772 (N_17772,N_7742,N_8171);
or U17773 (N_17773,N_8284,N_9204);
nor U17774 (N_17774,N_7384,N_3608);
xor U17775 (N_17775,N_9184,N_8858);
or U17776 (N_17776,N_4841,N_4289);
nor U17777 (N_17777,N_8972,N_6319);
nand U17778 (N_17778,N_5686,N_3932);
nand U17779 (N_17779,N_4387,N_2621);
and U17780 (N_17780,N_5346,N_7501);
and U17781 (N_17781,N_768,N_2244);
nor U17782 (N_17782,N_6194,N_1422);
and U17783 (N_17783,N_5749,N_5355);
nand U17784 (N_17784,N_6453,N_2339);
nand U17785 (N_17785,N_2155,N_4807);
nand U17786 (N_17786,N_5995,N_4583);
xnor U17787 (N_17787,N_5625,N_6937);
nor U17788 (N_17788,N_1369,N_1483);
nor U17789 (N_17789,N_2451,N_4517);
nor U17790 (N_17790,N_5628,N_3478);
or U17791 (N_17791,N_7537,N_3409);
nor U17792 (N_17792,N_9260,N_6427);
and U17793 (N_17793,N_3434,N_814);
and U17794 (N_17794,N_8625,N_4589);
or U17795 (N_17795,N_9538,N_2920);
and U17796 (N_17796,N_8427,N_7971);
nand U17797 (N_17797,N_8458,N_517);
nor U17798 (N_17798,N_2556,N_4680);
nand U17799 (N_17799,N_6808,N_7770);
and U17800 (N_17800,N_8952,N_2284);
and U17801 (N_17801,N_1048,N_8429);
xnor U17802 (N_17802,N_9169,N_2650);
and U17803 (N_17803,N_1696,N_7169);
nand U17804 (N_17804,N_7986,N_1590);
xnor U17805 (N_17805,N_7211,N_4343);
nand U17806 (N_17806,N_1898,N_8137);
and U17807 (N_17807,N_5026,N_7006);
nand U17808 (N_17808,N_2520,N_6245);
and U17809 (N_17809,N_9488,N_121);
nand U17810 (N_17810,N_548,N_589);
and U17811 (N_17811,N_1633,N_1295);
nor U17812 (N_17812,N_7504,N_6820);
or U17813 (N_17813,N_64,N_6282);
and U17814 (N_17814,N_8080,N_2097);
nor U17815 (N_17815,N_4778,N_6054);
nor U17816 (N_17816,N_6450,N_738);
or U17817 (N_17817,N_5527,N_3278);
nor U17818 (N_17818,N_6260,N_4181);
nor U17819 (N_17819,N_7616,N_2449);
nand U17820 (N_17820,N_1651,N_1427);
nand U17821 (N_17821,N_749,N_1509);
nand U17822 (N_17822,N_712,N_8263);
nand U17823 (N_17823,N_3975,N_9463);
nand U17824 (N_17824,N_2696,N_6567);
and U17825 (N_17825,N_4695,N_7284);
or U17826 (N_17826,N_1705,N_9106);
nand U17827 (N_17827,N_1049,N_1909);
or U17828 (N_17828,N_3685,N_2004);
nand U17829 (N_17829,N_8003,N_7564);
xor U17830 (N_17830,N_8585,N_3261);
nor U17831 (N_17831,N_8765,N_4171);
nand U17832 (N_17832,N_4265,N_3820);
nor U17833 (N_17833,N_7083,N_7112);
xor U17834 (N_17834,N_7793,N_2335);
or U17835 (N_17835,N_5644,N_2424);
and U17836 (N_17836,N_7074,N_2328);
and U17837 (N_17837,N_9153,N_2730);
or U17838 (N_17838,N_5858,N_5394);
or U17839 (N_17839,N_4802,N_8448);
and U17840 (N_17840,N_5410,N_8067);
nand U17841 (N_17841,N_7755,N_381);
xor U17842 (N_17842,N_9666,N_3408);
nand U17843 (N_17843,N_8831,N_2028);
and U17844 (N_17844,N_520,N_2953);
xor U17845 (N_17845,N_9432,N_9683);
nand U17846 (N_17846,N_598,N_7110);
nand U17847 (N_17847,N_5268,N_2539);
and U17848 (N_17848,N_9351,N_5251);
xor U17849 (N_17849,N_1783,N_4747);
and U17850 (N_17850,N_4791,N_3451);
or U17851 (N_17851,N_489,N_3063);
and U17852 (N_17852,N_7577,N_269);
xor U17853 (N_17853,N_3153,N_366);
nand U17854 (N_17854,N_9653,N_8016);
or U17855 (N_17855,N_2910,N_8619);
nor U17856 (N_17856,N_7429,N_9660);
and U17857 (N_17857,N_9264,N_201);
or U17858 (N_17858,N_1007,N_1980);
and U17859 (N_17859,N_656,N_6367);
xor U17860 (N_17860,N_7779,N_1660);
and U17861 (N_17861,N_5136,N_4647);
xnor U17862 (N_17862,N_4406,N_9878);
nor U17863 (N_17863,N_3440,N_9050);
nand U17864 (N_17864,N_1456,N_6899);
or U17865 (N_17865,N_7754,N_587);
nor U17866 (N_17866,N_3767,N_8775);
nand U17867 (N_17867,N_8089,N_20);
or U17868 (N_17868,N_3899,N_9814);
nand U17869 (N_17869,N_4282,N_2530);
xnor U17870 (N_17870,N_7688,N_9285);
and U17871 (N_17871,N_7487,N_21);
nand U17872 (N_17872,N_1064,N_1136);
nand U17873 (N_17873,N_8347,N_1812);
and U17874 (N_17874,N_6961,N_1552);
or U17875 (N_17875,N_6733,N_7218);
and U17876 (N_17876,N_1542,N_5615);
and U17877 (N_17877,N_6700,N_443);
and U17878 (N_17878,N_9935,N_1547);
or U17879 (N_17879,N_8119,N_1643);
nand U17880 (N_17880,N_4482,N_9303);
or U17881 (N_17881,N_3369,N_5502);
nand U17882 (N_17882,N_2653,N_5563);
nor U17883 (N_17883,N_7603,N_4987);
nand U17884 (N_17884,N_4680,N_2309);
nand U17885 (N_17885,N_3955,N_2657);
xor U17886 (N_17886,N_830,N_1759);
nand U17887 (N_17887,N_2880,N_3877);
nor U17888 (N_17888,N_928,N_8713);
or U17889 (N_17889,N_4847,N_2564);
nor U17890 (N_17890,N_8932,N_6406);
xor U17891 (N_17891,N_1031,N_6000);
and U17892 (N_17892,N_4050,N_129);
and U17893 (N_17893,N_4985,N_2514);
nor U17894 (N_17894,N_8153,N_5766);
nor U17895 (N_17895,N_928,N_9622);
and U17896 (N_17896,N_7758,N_6414);
or U17897 (N_17897,N_8505,N_5581);
or U17898 (N_17898,N_7342,N_2032);
and U17899 (N_17899,N_5074,N_2590);
xnor U17900 (N_17900,N_7861,N_1530);
xnor U17901 (N_17901,N_7407,N_4222);
nand U17902 (N_17902,N_5957,N_7957);
nor U17903 (N_17903,N_1164,N_1425);
nor U17904 (N_17904,N_5824,N_1425);
and U17905 (N_17905,N_5737,N_4265);
or U17906 (N_17906,N_3372,N_3240);
nor U17907 (N_17907,N_2250,N_679);
and U17908 (N_17908,N_4301,N_1942);
nand U17909 (N_17909,N_9997,N_9998);
nor U17910 (N_17910,N_3716,N_2079);
xnor U17911 (N_17911,N_8466,N_1836);
and U17912 (N_17912,N_5348,N_1413);
nor U17913 (N_17913,N_3068,N_1051);
nor U17914 (N_17914,N_2075,N_1484);
nand U17915 (N_17915,N_7984,N_3285);
nor U17916 (N_17916,N_1447,N_8772);
xor U17917 (N_17917,N_5724,N_2144);
or U17918 (N_17918,N_1830,N_8802);
or U17919 (N_17919,N_9039,N_5294);
or U17920 (N_17920,N_7144,N_3654);
nand U17921 (N_17921,N_7028,N_8119);
xnor U17922 (N_17922,N_9220,N_8267);
nand U17923 (N_17923,N_7563,N_6346);
or U17924 (N_17924,N_4617,N_5795);
and U17925 (N_17925,N_2946,N_8530);
nand U17926 (N_17926,N_3136,N_5679);
xnor U17927 (N_17927,N_2983,N_8325);
nand U17928 (N_17928,N_8572,N_9824);
xnor U17929 (N_17929,N_6284,N_2309);
xor U17930 (N_17930,N_9175,N_1111);
and U17931 (N_17931,N_7231,N_8504);
or U17932 (N_17932,N_3193,N_6189);
and U17933 (N_17933,N_3899,N_4414);
nor U17934 (N_17934,N_2493,N_451);
nand U17935 (N_17935,N_5891,N_8841);
and U17936 (N_17936,N_6702,N_3692);
nand U17937 (N_17937,N_3660,N_9330);
xnor U17938 (N_17938,N_3512,N_4065);
and U17939 (N_17939,N_5449,N_2284);
nand U17940 (N_17940,N_8321,N_4501);
xnor U17941 (N_17941,N_6843,N_4515);
or U17942 (N_17942,N_673,N_7189);
nand U17943 (N_17943,N_75,N_7953);
nor U17944 (N_17944,N_629,N_3582);
or U17945 (N_17945,N_5673,N_7766);
nand U17946 (N_17946,N_2158,N_4304);
or U17947 (N_17947,N_4572,N_7586);
and U17948 (N_17948,N_9770,N_3885);
xor U17949 (N_17949,N_8293,N_2907);
xnor U17950 (N_17950,N_3977,N_1558);
nor U17951 (N_17951,N_361,N_2731);
and U17952 (N_17952,N_4522,N_5901);
and U17953 (N_17953,N_4526,N_4439);
nor U17954 (N_17954,N_5721,N_3729);
nand U17955 (N_17955,N_8300,N_474);
or U17956 (N_17956,N_119,N_867);
and U17957 (N_17957,N_2519,N_5714);
nor U17958 (N_17958,N_9319,N_1334);
and U17959 (N_17959,N_4305,N_739);
and U17960 (N_17960,N_4740,N_8746);
nor U17961 (N_17961,N_1219,N_5325);
nor U17962 (N_17962,N_5411,N_4324);
or U17963 (N_17963,N_363,N_508);
nor U17964 (N_17964,N_1312,N_225);
and U17965 (N_17965,N_2784,N_8277);
nor U17966 (N_17966,N_7726,N_5818);
or U17967 (N_17967,N_5162,N_3229);
nor U17968 (N_17968,N_9609,N_6789);
nand U17969 (N_17969,N_387,N_62);
or U17970 (N_17970,N_7588,N_8744);
xor U17971 (N_17971,N_135,N_968);
and U17972 (N_17972,N_2005,N_3239);
nor U17973 (N_17973,N_2375,N_5270);
xor U17974 (N_17974,N_2787,N_8180);
xnor U17975 (N_17975,N_1007,N_7934);
nor U17976 (N_17976,N_8694,N_441);
nand U17977 (N_17977,N_2477,N_3923);
nand U17978 (N_17978,N_5452,N_6028);
nor U17979 (N_17979,N_1716,N_8043);
nand U17980 (N_17980,N_9300,N_354);
nor U17981 (N_17981,N_4283,N_9687);
nor U17982 (N_17982,N_4639,N_390);
nor U17983 (N_17983,N_6171,N_7377);
and U17984 (N_17984,N_7956,N_1867);
nor U17985 (N_17985,N_1877,N_1269);
xor U17986 (N_17986,N_4177,N_6857);
nand U17987 (N_17987,N_7476,N_8832);
or U17988 (N_17988,N_3726,N_2073);
and U17989 (N_17989,N_2440,N_595);
and U17990 (N_17990,N_7987,N_4241);
nand U17991 (N_17991,N_3429,N_6650);
nand U17992 (N_17992,N_9039,N_5629);
nor U17993 (N_17993,N_4097,N_1885);
nor U17994 (N_17994,N_5573,N_6872);
nand U17995 (N_17995,N_6906,N_7850);
nand U17996 (N_17996,N_7556,N_2992);
or U17997 (N_17997,N_818,N_7812);
and U17998 (N_17998,N_8346,N_9355);
nor U17999 (N_17999,N_7033,N_3694);
nor U18000 (N_18000,N_2350,N_4024);
or U18001 (N_18001,N_1913,N_5688);
or U18002 (N_18002,N_9748,N_6417);
nand U18003 (N_18003,N_8413,N_532);
nor U18004 (N_18004,N_1300,N_9570);
nor U18005 (N_18005,N_5436,N_6102);
and U18006 (N_18006,N_3269,N_2554);
and U18007 (N_18007,N_6870,N_1276);
nand U18008 (N_18008,N_49,N_7224);
nand U18009 (N_18009,N_6978,N_2565);
and U18010 (N_18010,N_1575,N_2283);
nor U18011 (N_18011,N_6657,N_7042);
nor U18012 (N_18012,N_4257,N_7504);
and U18013 (N_18013,N_8168,N_5719);
or U18014 (N_18014,N_4766,N_1804);
or U18015 (N_18015,N_4112,N_8033);
or U18016 (N_18016,N_611,N_7707);
nor U18017 (N_18017,N_1018,N_5931);
or U18018 (N_18018,N_8554,N_958);
nor U18019 (N_18019,N_9639,N_2817);
nor U18020 (N_18020,N_2023,N_2228);
nand U18021 (N_18021,N_2258,N_6221);
nor U18022 (N_18022,N_8420,N_5032);
or U18023 (N_18023,N_9702,N_7597);
nor U18024 (N_18024,N_3523,N_5908);
nor U18025 (N_18025,N_904,N_2057);
or U18026 (N_18026,N_6744,N_5781);
and U18027 (N_18027,N_5706,N_7686);
or U18028 (N_18028,N_8707,N_3725);
or U18029 (N_18029,N_3894,N_5142);
or U18030 (N_18030,N_4902,N_9186);
and U18031 (N_18031,N_9373,N_1304);
or U18032 (N_18032,N_1489,N_4199);
and U18033 (N_18033,N_9964,N_9132);
and U18034 (N_18034,N_6969,N_9569);
nor U18035 (N_18035,N_2243,N_1351);
nand U18036 (N_18036,N_521,N_4371);
nor U18037 (N_18037,N_439,N_1951);
and U18038 (N_18038,N_9337,N_8714);
xnor U18039 (N_18039,N_7364,N_5131);
and U18040 (N_18040,N_8180,N_7010);
nand U18041 (N_18041,N_329,N_3608);
and U18042 (N_18042,N_5657,N_5096);
nor U18043 (N_18043,N_3672,N_8206);
nand U18044 (N_18044,N_7383,N_5974);
and U18045 (N_18045,N_6976,N_3005);
nand U18046 (N_18046,N_5526,N_9516);
or U18047 (N_18047,N_216,N_4052);
and U18048 (N_18048,N_3018,N_5740);
and U18049 (N_18049,N_5598,N_5070);
or U18050 (N_18050,N_5322,N_6872);
xnor U18051 (N_18051,N_3989,N_9610);
nand U18052 (N_18052,N_5853,N_4324);
and U18053 (N_18053,N_7649,N_5087);
nand U18054 (N_18054,N_7651,N_8358);
or U18055 (N_18055,N_5571,N_7171);
or U18056 (N_18056,N_6672,N_9070);
nand U18057 (N_18057,N_8613,N_6781);
nor U18058 (N_18058,N_1087,N_4041);
nor U18059 (N_18059,N_1787,N_6320);
and U18060 (N_18060,N_2652,N_4588);
and U18061 (N_18061,N_3197,N_771);
nand U18062 (N_18062,N_8970,N_8065);
nor U18063 (N_18063,N_3501,N_4356);
nand U18064 (N_18064,N_8311,N_616);
or U18065 (N_18065,N_9789,N_2892);
or U18066 (N_18066,N_6838,N_3841);
nor U18067 (N_18067,N_8362,N_7650);
nand U18068 (N_18068,N_6623,N_1026);
and U18069 (N_18069,N_2981,N_7214);
xnor U18070 (N_18070,N_3898,N_3954);
or U18071 (N_18071,N_6173,N_5011);
nor U18072 (N_18072,N_2881,N_4941);
nor U18073 (N_18073,N_52,N_9073);
and U18074 (N_18074,N_4592,N_1403);
nand U18075 (N_18075,N_3976,N_4932);
or U18076 (N_18076,N_9021,N_5576);
or U18077 (N_18077,N_7813,N_9467);
nor U18078 (N_18078,N_1874,N_2375);
or U18079 (N_18079,N_8856,N_5216);
nor U18080 (N_18080,N_7324,N_6738);
nand U18081 (N_18081,N_8,N_470);
and U18082 (N_18082,N_5028,N_553);
nor U18083 (N_18083,N_9633,N_6471);
nor U18084 (N_18084,N_5298,N_1312);
nor U18085 (N_18085,N_9833,N_4842);
nor U18086 (N_18086,N_5011,N_6516);
and U18087 (N_18087,N_8147,N_157);
or U18088 (N_18088,N_1803,N_1799);
xnor U18089 (N_18089,N_7311,N_7647);
and U18090 (N_18090,N_5670,N_9086);
and U18091 (N_18091,N_2838,N_304);
nand U18092 (N_18092,N_5772,N_1658);
nor U18093 (N_18093,N_5632,N_6081);
nand U18094 (N_18094,N_6010,N_3698);
nor U18095 (N_18095,N_8062,N_4321);
and U18096 (N_18096,N_9982,N_9272);
nor U18097 (N_18097,N_2079,N_4842);
xnor U18098 (N_18098,N_1827,N_6630);
xor U18099 (N_18099,N_5291,N_7336);
and U18100 (N_18100,N_4173,N_7756);
nand U18101 (N_18101,N_5235,N_1025);
nand U18102 (N_18102,N_9667,N_5919);
nand U18103 (N_18103,N_3748,N_7748);
nand U18104 (N_18104,N_4289,N_7696);
nor U18105 (N_18105,N_3112,N_4236);
nand U18106 (N_18106,N_2526,N_9404);
and U18107 (N_18107,N_2346,N_1474);
xor U18108 (N_18108,N_8925,N_2665);
or U18109 (N_18109,N_2081,N_5386);
nand U18110 (N_18110,N_838,N_1829);
nor U18111 (N_18111,N_2431,N_424);
nor U18112 (N_18112,N_4411,N_2627);
or U18113 (N_18113,N_569,N_195);
or U18114 (N_18114,N_2129,N_148);
nor U18115 (N_18115,N_9920,N_5672);
or U18116 (N_18116,N_9550,N_5881);
nand U18117 (N_18117,N_9532,N_1907);
xnor U18118 (N_18118,N_3320,N_3191);
nand U18119 (N_18119,N_3032,N_8575);
nor U18120 (N_18120,N_2342,N_3520);
and U18121 (N_18121,N_7764,N_5669);
nor U18122 (N_18122,N_4163,N_7038);
nand U18123 (N_18123,N_5222,N_2366);
and U18124 (N_18124,N_5611,N_146);
nor U18125 (N_18125,N_3644,N_4277);
and U18126 (N_18126,N_9847,N_1741);
or U18127 (N_18127,N_5733,N_2879);
nand U18128 (N_18128,N_2701,N_5431);
nand U18129 (N_18129,N_5332,N_9373);
nand U18130 (N_18130,N_933,N_9325);
nand U18131 (N_18131,N_1678,N_4194);
or U18132 (N_18132,N_9349,N_6558);
nor U18133 (N_18133,N_1914,N_9851);
nand U18134 (N_18134,N_3313,N_4333);
and U18135 (N_18135,N_9983,N_7778);
nand U18136 (N_18136,N_9071,N_4334);
nor U18137 (N_18137,N_9901,N_5131);
or U18138 (N_18138,N_574,N_3254);
and U18139 (N_18139,N_1272,N_8589);
and U18140 (N_18140,N_6193,N_8944);
nand U18141 (N_18141,N_9119,N_4708);
or U18142 (N_18142,N_7979,N_7299);
or U18143 (N_18143,N_8464,N_2514);
nor U18144 (N_18144,N_6825,N_4602);
and U18145 (N_18145,N_6723,N_1362);
xnor U18146 (N_18146,N_4631,N_2328);
nor U18147 (N_18147,N_8761,N_1410);
and U18148 (N_18148,N_9963,N_5737);
nand U18149 (N_18149,N_2724,N_9846);
and U18150 (N_18150,N_9617,N_2088);
xor U18151 (N_18151,N_9607,N_765);
nor U18152 (N_18152,N_6280,N_5739);
nor U18153 (N_18153,N_1673,N_3097);
and U18154 (N_18154,N_4196,N_2264);
nor U18155 (N_18155,N_1855,N_2862);
nor U18156 (N_18156,N_4398,N_6014);
and U18157 (N_18157,N_4010,N_1282);
nand U18158 (N_18158,N_2648,N_9051);
nor U18159 (N_18159,N_7347,N_4087);
or U18160 (N_18160,N_6854,N_7165);
and U18161 (N_18161,N_6916,N_5226);
nand U18162 (N_18162,N_6789,N_2885);
and U18163 (N_18163,N_4533,N_1601);
nor U18164 (N_18164,N_5171,N_3223);
nor U18165 (N_18165,N_5399,N_8568);
nand U18166 (N_18166,N_5172,N_2713);
and U18167 (N_18167,N_2946,N_5727);
and U18168 (N_18168,N_9483,N_11);
or U18169 (N_18169,N_917,N_3431);
and U18170 (N_18170,N_5696,N_8618);
xnor U18171 (N_18171,N_9892,N_7351);
or U18172 (N_18172,N_8291,N_9607);
or U18173 (N_18173,N_6956,N_3197);
xnor U18174 (N_18174,N_599,N_1592);
nand U18175 (N_18175,N_3396,N_5198);
nor U18176 (N_18176,N_847,N_6523);
xnor U18177 (N_18177,N_8746,N_6947);
or U18178 (N_18178,N_7095,N_2051);
nand U18179 (N_18179,N_8745,N_4534);
and U18180 (N_18180,N_2023,N_3544);
or U18181 (N_18181,N_4676,N_1209);
and U18182 (N_18182,N_807,N_4897);
nor U18183 (N_18183,N_6769,N_3602);
or U18184 (N_18184,N_5676,N_8584);
nand U18185 (N_18185,N_5882,N_1335);
nand U18186 (N_18186,N_2692,N_3568);
and U18187 (N_18187,N_2358,N_6274);
nand U18188 (N_18188,N_4997,N_1104);
nand U18189 (N_18189,N_8899,N_9506);
xnor U18190 (N_18190,N_1140,N_1912);
xor U18191 (N_18191,N_1325,N_4433);
xnor U18192 (N_18192,N_8913,N_2253);
nor U18193 (N_18193,N_574,N_9779);
nor U18194 (N_18194,N_2092,N_7043);
nor U18195 (N_18195,N_5113,N_7111);
nor U18196 (N_18196,N_4809,N_9508);
nor U18197 (N_18197,N_3761,N_6127);
nand U18198 (N_18198,N_1074,N_3064);
or U18199 (N_18199,N_5368,N_6058);
nand U18200 (N_18200,N_5848,N_1722);
xnor U18201 (N_18201,N_4512,N_305);
nand U18202 (N_18202,N_667,N_8337);
xor U18203 (N_18203,N_810,N_3462);
or U18204 (N_18204,N_4435,N_304);
nor U18205 (N_18205,N_9111,N_6895);
nor U18206 (N_18206,N_1032,N_9872);
nand U18207 (N_18207,N_9602,N_5026);
and U18208 (N_18208,N_2579,N_8909);
nor U18209 (N_18209,N_1008,N_8567);
and U18210 (N_18210,N_4929,N_8212);
nor U18211 (N_18211,N_1548,N_96);
and U18212 (N_18212,N_2527,N_2672);
and U18213 (N_18213,N_428,N_5874);
nand U18214 (N_18214,N_5304,N_1305);
or U18215 (N_18215,N_7289,N_8841);
or U18216 (N_18216,N_2891,N_6063);
nor U18217 (N_18217,N_1934,N_3097);
nor U18218 (N_18218,N_9779,N_8770);
and U18219 (N_18219,N_4963,N_8821);
nand U18220 (N_18220,N_8644,N_1627);
or U18221 (N_18221,N_3739,N_2267);
and U18222 (N_18222,N_9940,N_539);
and U18223 (N_18223,N_6271,N_7571);
nor U18224 (N_18224,N_5567,N_3283);
or U18225 (N_18225,N_8153,N_6474);
and U18226 (N_18226,N_8526,N_6606);
and U18227 (N_18227,N_1368,N_9084);
xor U18228 (N_18228,N_6908,N_1490);
or U18229 (N_18229,N_7019,N_1614);
xor U18230 (N_18230,N_7839,N_4418);
nor U18231 (N_18231,N_3502,N_9022);
nand U18232 (N_18232,N_8473,N_7840);
or U18233 (N_18233,N_878,N_445);
and U18234 (N_18234,N_9615,N_4065);
nand U18235 (N_18235,N_8047,N_4722);
and U18236 (N_18236,N_4932,N_902);
and U18237 (N_18237,N_3650,N_2171);
nand U18238 (N_18238,N_7613,N_56);
nor U18239 (N_18239,N_849,N_4474);
nand U18240 (N_18240,N_5716,N_4952);
and U18241 (N_18241,N_5454,N_9583);
nor U18242 (N_18242,N_9819,N_4674);
or U18243 (N_18243,N_5260,N_4817);
and U18244 (N_18244,N_280,N_5121);
and U18245 (N_18245,N_4769,N_1337);
or U18246 (N_18246,N_261,N_826);
and U18247 (N_18247,N_9904,N_6141);
or U18248 (N_18248,N_7059,N_7135);
nand U18249 (N_18249,N_9226,N_8903);
nand U18250 (N_18250,N_7182,N_8460);
and U18251 (N_18251,N_1086,N_5472);
nor U18252 (N_18252,N_9074,N_8331);
xor U18253 (N_18253,N_3320,N_7333);
nor U18254 (N_18254,N_4187,N_4847);
or U18255 (N_18255,N_6154,N_1832);
or U18256 (N_18256,N_4058,N_2335);
nor U18257 (N_18257,N_9451,N_3138);
xor U18258 (N_18258,N_1299,N_336);
nand U18259 (N_18259,N_6879,N_5016);
or U18260 (N_18260,N_4504,N_8533);
nor U18261 (N_18261,N_1298,N_6871);
and U18262 (N_18262,N_2355,N_1912);
and U18263 (N_18263,N_5225,N_4212);
xor U18264 (N_18264,N_2920,N_3646);
or U18265 (N_18265,N_9512,N_8253);
nor U18266 (N_18266,N_6695,N_3026);
and U18267 (N_18267,N_4874,N_6700);
nand U18268 (N_18268,N_6614,N_9957);
xnor U18269 (N_18269,N_5061,N_2042);
nor U18270 (N_18270,N_2787,N_2092);
nand U18271 (N_18271,N_2707,N_9896);
nand U18272 (N_18272,N_489,N_9090);
xor U18273 (N_18273,N_1342,N_3710);
and U18274 (N_18274,N_8249,N_3007);
nor U18275 (N_18275,N_7909,N_1092);
nor U18276 (N_18276,N_904,N_1876);
nand U18277 (N_18277,N_159,N_3093);
nor U18278 (N_18278,N_7225,N_5788);
and U18279 (N_18279,N_4431,N_4491);
or U18280 (N_18280,N_3814,N_2786);
or U18281 (N_18281,N_1201,N_4423);
nor U18282 (N_18282,N_7784,N_5663);
or U18283 (N_18283,N_4981,N_9586);
nand U18284 (N_18284,N_8566,N_1480);
nand U18285 (N_18285,N_6271,N_4281);
or U18286 (N_18286,N_9316,N_1459);
nand U18287 (N_18287,N_5218,N_8006);
and U18288 (N_18288,N_2214,N_4113);
or U18289 (N_18289,N_2540,N_6772);
and U18290 (N_18290,N_3530,N_743);
nand U18291 (N_18291,N_6759,N_3497);
or U18292 (N_18292,N_2284,N_7002);
xor U18293 (N_18293,N_4124,N_6608);
xor U18294 (N_18294,N_2608,N_8503);
xor U18295 (N_18295,N_2010,N_3325);
and U18296 (N_18296,N_9498,N_9236);
and U18297 (N_18297,N_6642,N_1983);
and U18298 (N_18298,N_304,N_4348);
xor U18299 (N_18299,N_3673,N_2430);
nor U18300 (N_18300,N_2388,N_5696);
nand U18301 (N_18301,N_4886,N_7149);
xor U18302 (N_18302,N_3620,N_130);
and U18303 (N_18303,N_3901,N_7834);
xor U18304 (N_18304,N_5441,N_2806);
and U18305 (N_18305,N_5481,N_3505);
and U18306 (N_18306,N_5458,N_9495);
or U18307 (N_18307,N_8563,N_7078);
nand U18308 (N_18308,N_4083,N_8780);
and U18309 (N_18309,N_8213,N_9128);
nand U18310 (N_18310,N_2605,N_8096);
and U18311 (N_18311,N_6096,N_2621);
nor U18312 (N_18312,N_3954,N_1860);
or U18313 (N_18313,N_1372,N_1954);
and U18314 (N_18314,N_7384,N_7298);
or U18315 (N_18315,N_2804,N_7740);
or U18316 (N_18316,N_8160,N_3394);
nor U18317 (N_18317,N_2258,N_5929);
nand U18318 (N_18318,N_9822,N_2654);
or U18319 (N_18319,N_6355,N_3460);
or U18320 (N_18320,N_2994,N_5966);
nand U18321 (N_18321,N_7708,N_6975);
nand U18322 (N_18322,N_5945,N_2327);
nor U18323 (N_18323,N_730,N_8924);
and U18324 (N_18324,N_4921,N_8445);
or U18325 (N_18325,N_1822,N_1275);
nand U18326 (N_18326,N_3842,N_8408);
and U18327 (N_18327,N_3671,N_6760);
nand U18328 (N_18328,N_6525,N_7282);
or U18329 (N_18329,N_1070,N_8569);
nor U18330 (N_18330,N_871,N_456);
nand U18331 (N_18331,N_9927,N_8044);
nand U18332 (N_18332,N_7097,N_7606);
xnor U18333 (N_18333,N_8535,N_4577);
nand U18334 (N_18334,N_5348,N_8039);
xor U18335 (N_18335,N_5982,N_5408);
or U18336 (N_18336,N_491,N_8366);
xor U18337 (N_18337,N_54,N_7141);
and U18338 (N_18338,N_2146,N_5849);
nor U18339 (N_18339,N_5937,N_1748);
or U18340 (N_18340,N_6107,N_3889);
or U18341 (N_18341,N_2885,N_340);
or U18342 (N_18342,N_7533,N_3905);
or U18343 (N_18343,N_1423,N_9966);
or U18344 (N_18344,N_4424,N_3345);
nor U18345 (N_18345,N_8234,N_1407);
and U18346 (N_18346,N_5696,N_6175);
nor U18347 (N_18347,N_6668,N_7904);
and U18348 (N_18348,N_5033,N_2902);
or U18349 (N_18349,N_9006,N_7982);
nor U18350 (N_18350,N_1710,N_1477);
and U18351 (N_18351,N_8201,N_9358);
and U18352 (N_18352,N_6692,N_5474);
xnor U18353 (N_18353,N_1988,N_4465);
nand U18354 (N_18354,N_5237,N_4824);
nor U18355 (N_18355,N_8649,N_4789);
nor U18356 (N_18356,N_1280,N_7112);
nor U18357 (N_18357,N_5200,N_3418);
and U18358 (N_18358,N_7459,N_5225);
and U18359 (N_18359,N_103,N_7026);
nand U18360 (N_18360,N_608,N_367);
and U18361 (N_18361,N_5167,N_6822);
or U18362 (N_18362,N_459,N_9829);
and U18363 (N_18363,N_7636,N_547);
or U18364 (N_18364,N_8792,N_5940);
xor U18365 (N_18365,N_9429,N_8295);
nor U18366 (N_18366,N_9905,N_4425);
nor U18367 (N_18367,N_5278,N_992);
nor U18368 (N_18368,N_2069,N_5038);
and U18369 (N_18369,N_9739,N_9362);
xnor U18370 (N_18370,N_3321,N_8326);
nor U18371 (N_18371,N_5000,N_1835);
or U18372 (N_18372,N_7950,N_7225);
and U18373 (N_18373,N_9714,N_3544);
nand U18374 (N_18374,N_7850,N_8314);
nand U18375 (N_18375,N_4448,N_9511);
or U18376 (N_18376,N_3847,N_8997);
nor U18377 (N_18377,N_4512,N_7874);
xor U18378 (N_18378,N_7654,N_600);
nand U18379 (N_18379,N_2178,N_2033);
or U18380 (N_18380,N_4084,N_6642);
nor U18381 (N_18381,N_4963,N_5562);
and U18382 (N_18382,N_9919,N_9982);
and U18383 (N_18383,N_6270,N_667);
nor U18384 (N_18384,N_3601,N_8117);
and U18385 (N_18385,N_8909,N_3380);
or U18386 (N_18386,N_2832,N_8864);
nand U18387 (N_18387,N_8147,N_5701);
xor U18388 (N_18388,N_723,N_5772);
and U18389 (N_18389,N_6918,N_499);
nand U18390 (N_18390,N_7447,N_6538);
and U18391 (N_18391,N_6687,N_183);
or U18392 (N_18392,N_8230,N_2091);
xnor U18393 (N_18393,N_6680,N_8723);
nand U18394 (N_18394,N_1262,N_6073);
nor U18395 (N_18395,N_6428,N_2104);
xor U18396 (N_18396,N_3523,N_6251);
nand U18397 (N_18397,N_5886,N_3554);
or U18398 (N_18398,N_3545,N_2758);
or U18399 (N_18399,N_8222,N_2849);
and U18400 (N_18400,N_8606,N_8123);
nor U18401 (N_18401,N_9004,N_1005);
nor U18402 (N_18402,N_6179,N_7095);
and U18403 (N_18403,N_4582,N_4909);
nand U18404 (N_18404,N_2897,N_8362);
and U18405 (N_18405,N_9694,N_6925);
xor U18406 (N_18406,N_9178,N_4034);
nand U18407 (N_18407,N_6548,N_4771);
nand U18408 (N_18408,N_9620,N_6829);
xor U18409 (N_18409,N_6995,N_5436);
or U18410 (N_18410,N_9445,N_7290);
nor U18411 (N_18411,N_6714,N_6236);
nor U18412 (N_18412,N_4664,N_131);
nand U18413 (N_18413,N_3761,N_708);
and U18414 (N_18414,N_1396,N_8513);
nand U18415 (N_18415,N_9499,N_6317);
or U18416 (N_18416,N_6394,N_484);
or U18417 (N_18417,N_708,N_1970);
nor U18418 (N_18418,N_6465,N_8138);
nand U18419 (N_18419,N_873,N_7462);
nor U18420 (N_18420,N_1440,N_5101);
nor U18421 (N_18421,N_5532,N_2881);
nor U18422 (N_18422,N_2639,N_4934);
and U18423 (N_18423,N_6314,N_5205);
or U18424 (N_18424,N_1670,N_6761);
nand U18425 (N_18425,N_8935,N_7206);
and U18426 (N_18426,N_9089,N_9814);
and U18427 (N_18427,N_6638,N_9276);
nand U18428 (N_18428,N_6751,N_8358);
and U18429 (N_18429,N_8048,N_214);
or U18430 (N_18430,N_9866,N_31);
nor U18431 (N_18431,N_49,N_1159);
nand U18432 (N_18432,N_8032,N_8669);
and U18433 (N_18433,N_4216,N_8471);
nor U18434 (N_18434,N_7698,N_8792);
xor U18435 (N_18435,N_8701,N_3587);
xnor U18436 (N_18436,N_157,N_810);
nand U18437 (N_18437,N_762,N_9183);
xor U18438 (N_18438,N_4775,N_2896);
nor U18439 (N_18439,N_6300,N_7728);
nand U18440 (N_18440,N_5938,N_6553);
nand U18441 (N_18441,N_4403,N_4091);
or U18442 (N_18442,N_3816,N_758);
or U18443 (N_18443,N_8577,N_8707);
or U18444 (N_18444,N_9385,N_9595);
and U18445 (N_18445,N_3679,N_7729);
and U18446 (N_18446,N_7167,N_9669);
and U18447 (N_18447,N_3372,N_4444);
nand U18448 (N_18448,N_8828,N_64);
nor U18449 (N_18449,N_541,N_8635);
or U18450 (N_18450,N_7454,N_6178);
or U18451 (N_18451,N_8597,N_4107);
nand U18452 (N_18452,N_4797,N_1150);
or U18453 (N_18453,N_8074,N_4207);
or U18454 (N_18454,N_3756,N_4693);
and U18455 (N_18455,N_1122,N_447);
and U18456 (N_18456,N_5675,N_3070);
and U18457 (N_18457,N_3607,N_9990);
nor U18458 (N_18458,N_3918,N_3620);
nor U18459 (N_18459,N_8997,N_7013);
or U18460 (N_18460,N_7168,N_3214);
nand U18461 (N_18461,N_1601,N_2075);
nand U18462 (N_18462,N_8750,N_9135);
xor U18463 (N_18463,N_7022,N_3813);
nand U18464 (N_18464,N_7679,N_3751);
nand U18465 (N_18465,N_6437,N_9632);
and U18466 (N_18466,N_4690,N_5338);
and U18467 (N_18467,N_5449,N_1052);
or U18468 (N_18468,N_469,N_6027);
and U18469 (N_18469,N_9748,N_6228);
xor U18470 (N_18470,N_3434,N_5607);
or U18471 (N_18471,N_7359,N_1750);
and U18472 (N_18472,N_3982,N_8900);
or U18473 (N_18473,N_6408,N_6135);
nand U18474 (N_18474,N_9481,N_5247);
nor U18475 (N_18475,N_1968,N_9666);
and U18476 (N_18476,N_3188,N_9032);
nor U18477 (N_18477,N_1743,N_4342);
nor U18478 (N_18478,N_753,N_5923);
or U18479 (N_18479,N_9966,N_8032);
and U18480 (N_18480,N_8571,N_8594);
xnor U18481 (N_18481,N_2566,N_5266);
or U18482 (N_18482,N_6245,N_9097);
nor U18483 (N_18483,N_3077,N_6450);
nor U18484 (N_18484,N_4332,N_1787);
and U18485 (N_18485,N_6870,N_9243);
and U18486 (N_18486,N_9806,N_4857);
nor U18487 (N_18487,N_8820,N_5599);
nand U18488 (N_18488,N_1047,N_2153);
nor U18489 (N_18489,N_8283,N_7240);
or U18490 (N_18490,N_4984,N_273);
and U18491 (N_18491,N_490,N_7898);
or U18492 (N_18492,N_3537,N_5769);
nor U18493 (N_18493,N_8088,N_8996);
xor U18494 (N_18494,N_5094,N_3034);
or U18495 (N_18495,N_2256,N_3410);
xnor U18496 (N_18496,N_4189,N_3213);
nand U18497 (N_18497,N_8503,N_8104);
nor U18498 (N_18498,N_3997,N_60);
and U18499 (N_18499,N_5978,N_8414);
and U18500 (N_18500,N_4116,N_1687);
and U18501 (N_18501,N_4586,N_5132);
nand U18502 (N_18502,N_4638,N_6251);
and U18503 (N_18503,N_8607,N_3075);
and U18504 (N_18504,N_17,N_6256);
or U18505 (N_18505,N_7603,N_9492);
nand U18506 (N_18506,N_3312,N_842);
or U18507 (N_18507,N_8569,N_3626);
or U18508 (N_18508,N_4166,N_7416);
or U18509 (N_18509,N_7420,N_8258);
nor U18510 (N_18510,N_251,N_7568);
and U18511 (N_18511,N_2010,N_1168);
nand U18512 (N_18512,N_4356,N_9727);
or U18513 (N_18513,N_7942,N_1677);
and U18514 (N_18514,N_5831,N_370);
or U18515 (N_18515,N_5897,N_5182);
nand U18516 (N_18516,N_4973,N_9009);
nor U18517 (N_18517,N_2489,N_4199);
xor U18518 (N_18518,N_4104,N_7798);
and U18519 (N_18519,N_6825,N_2560);
nand U18520 (N_18520,N_4879,N_7933);
and U18521 (N_18521,N_183,N_5368);
nand U18522 (N_18522,N_3378,N_9498);
xor U18523 (N_18523,N_3275,N_2222);
and U18524 (N_18524,N_3290,N_4342);
or U18525 (N_18525,N_2970,N_4648);
and U18526 (N_18526,N_5532,N_3473);
and U18527 (N_18527,N_27,N_6733);
nor U18528 (N_18528,N_1320,N_6012);
nor U18529 (N_18529,N_2621,N_8271);
or U18530 (N_18530,N_2368,N_672);
nand U18531 (N_18531,N_4086,N_3791);
or U18532 (N_18532,N_5131,N_208);
and U18533 (N_18533,N_4734,N_9410);
nand U18534 (N_18534,N_7477,N_1801);
nor U18535 (N_18535,N_5252,N_7364);
or U18536 (N_18536,N_7738,N_8114);
nor U18537 (N_18537,N_2262,N_5287);
xor U18538 (N_18538,N_6483,N_9394);
nor U18539 (N_18539,N_7810,N_2620);
or U18540 (N_18540,N_6305,N_2558);
nand U18541 (N_18541,N_6831,N_8395);
and U18542 (N_18542,N_3119,N_4985);
and U18543 (N_18543,N_1385,N_4635);
and U18544 (N_18544,N_7728,N_7618);
nand U18545 (N_18545,N_8722,N_9106);
nor U18546 (N_18546,N_3986,N_9207);
and U18547 (N_18547,N_81,N_7178);
or U18548 (N_18548,N_911,N_4153);
or U18549 (N_18549,N_63,N_1504);
and U18550 (N_18550,N_9007,N_1590);
nand U18551 (N_18551,N_8895,N_6981);
nand U18552 (N_18552,N_9401,N_7840);
and U18553 (N_18553,N_7190,N_5192);
or U18554 (N_18554,N_1811,N_5528);
and U18555 (N_18555,N_4743,N_2123);
and U18556 (N_18556,N_9562,N_1837);
or U18557 (N_18557,N_1329,N_6811);
nand U18558 (N_18558,N_2479,N_2038);
and U18559 (N_18559,N_4278,N_6415);
nor U18560 (N_18560,N_4864,N_3199);
and U18561 (N_18561,N_7408,N_4196);
xnor U18562 (N_18562,N_1083,N_1567);
and U18563 (N_18563,N_1460,N_7155);
and U18564 (N_18564,N_3363,N_3881);
xnor U18565 (N_18565,N_2913,N_4150);
nand U18566 (N_18566,N_4584,N_4290);
xor U18567 (N_18567,N_7277,N_2839);
nor U18568 (N_18568,N_2514,N_1341);
xor U18569 (N_18569,N_6997,N_2068);
and U18570 (N_18570,N_8394,N_3638);
or U18571 (N_18571,N_3458,N_5732);
nand U18572 (N_18572,N_7538,N_7785);
nand U18573 (N_18573,N_7261,N_163);
or U18574 (N_18574,N_6573,N_6907);
nor U18575 (N_18575,N_8860,N_8606);
nor U18576 (N_18576,N_8944,N_3412);
nor U18577 (N_18577,N_8031,N_7602);
and U18578 (N_18578,N_7454,N_8687);
nor U18579 (N_18579,N_9802,N_2600);
nor U18580 (N_18580,N_6233,N_4937);
xor U18581 (N_18581,N_1037,N_5596);
xnor U18582 (N_18582,N_7781,N_6902);
or U18583 (N_18583,N_5490,N_3050);
or U18584 (N_18584,N_7153,N_9630);
xor U18585 (N_18585,N_6888,N_2482);
nand U18586 (N_18586,N_1498,N_781);
or U18587 (N_18587,N_9294,N_7281);
nor U18588 (N_18588,N_374,N_1088);
nand U18589 (N_18589,N_2427,N_8564);
or U18590 (N_18590,N_7930,N_3174);
nor U18591 (N_18591,N_7715,N_4573);
nand U18592 (N_18592,N_8547,N_5653);
nor U18593 (N_18593,N_1538,N_7333);
nor U18594 (N_18594,N_4189,N_7749);
and U18595 (N_18595,N_2101,N_922);
or U18596 (N_18596,N_5869,N_6480);
and U18597 (N_18597,N_921,N_3409);
nand U18598 (N_18598,N_254,N_1087);
nor U18599 (N_18599,N_1850,N_9306);
or U18600 (N_18600,N_9655,N_5226);
and U18601 (N_18601,N_6981,N_8833);
nor U18602 (N_18602,N_2909,N_6119);
xnor U18603 (N_18603,N_3980,N_9022);
nor U18604 (N_18604,N_6193,N_713);
and U18605 (N_18605,N_6622,N_6934);
nand U18606 (N_18606,N_6744,N_7502);
nand U18607 (N_18607,N_9596,N_5242);
xnor U18608 (N_18608,N_3380,N_7860);
nor U18609 (N_18609,N_2724,N_5313);
nor U18610 (N_18610,N_2029,N_8050);
nand U18611 (N_18611,N_7409,N_6900);
xor U18612 (N_18612,N_5767,N_8751);
and U18613 (N_18613,N_7054,N_334);
nor U18614 (N_18614,N_5289,N_3096);
and U18615 (N_18615,N_6392,N_1813);
nand U18616 (N_18616,N_4459,N_1929);
or U18617 (N_18617,N_511,N_4298);
or U18618 (N_18618,N_1497,N_955);
nor U18619 (N_18619,N_7345,N_3366);
nor U18620 (N_18620,N_6549,N_6041);
xor U18621 (N_18621,N_392,N_4485);
or U18622 (N_18622,N_6436,N_8923);
nand U18623 (N_18623,N_315,N_4481);
or U18624 (N_18624,N_9245,N_7559);
and U18625 (N_18625,N_7809,N_9720);
xor U18626 (N_18626,N_9013,N_4194);
nand U18627 (N_18627,N_9345,N_4149);
and U18628 (N_18628,N_7184,N_2184);
nor U18629 (N_18629,N_359,N_7025);
and U18630 (N_18630,N_4531,N_4782);
and U18631 (N_18631,N_7570,N_7544);
xnor U18632 (N_18632,N_7092,N_3718);
and U18633 (N_18633,N_9457,N_8934);
xnor U18634 (N_18634,N_9965,N_5794);
or U18635 (N_18635,N_1086,N_741);
and U18636 (N_18636,N_5335,N_9118);
and U18637 (N_18637,N_9677,N_2942);
nand U18638 (N_18638,N_5488,N_5766);
or U18639 (N_18639,N_7127,N_2761);
nand U18640 (N_18640,N_2100,N_319);
nand U18641 (N_18641,N_9810,N_4914);
and U18642 (N_18642,N_9791,N_3750);
nor U18643 (N_18643,N_5700,N_6593);
xnor U18644 (N_18644,N_5543,N_7755);
and U18645 (N_18645,N_8776,N_6436);
nor U18646 (N_18646,N_4322,N_215);
nand U18647 (N_18647,N_4281,N_7213);
xor U18648 (N_18648,N_876,N_9506);
nand U18649 (N_18649,N_5588,N_1707);
or U18650 (N_18650,N_7071,N_6312);
nor U18651 (N_18651,N_4390,N_1211);
nand U18652 (N_18652,N_7477,N_4199);
and U18653 (N_18653,N_7791,N_8035);
nand U18654 (N_18654,N_4282,N_2032);
nand U18655 (N_18655,N_7392,N_2925);
or U18656 (N_18656,N_4820,N_1144);
and U18657 (N_18657,N_8343,N_4210);
nor U18658 (N_18658,N_2216,N_3257);
and U18659 (N_18659,N_8664,N_9596);
nand U18660 (N_18660,N_7179,N_7033);
or U18661 (N_18661,N_3190,N_9778);
nor U18662 (N_18662,N_4545,N_8324);
nand U18663 (N_18663,N_3801,N_7077);
nand U18664 (N_18664,N_3739,N_114);
or U18665 (N_18665,N_8734,N_486);
nand U18666 (N_18666,N_1640,N_4291);
xnor U18667 (N_18667,N_2949,N_5718);
nand U18668 (N_18668,N_1538,N_2005);
and U18669 (N_18669,N_3313,N_3924);
nor U18670 (N_18670,N_100,N_5026);
nor U18671 (N_18671,N_2582,N_5433);
nor U18672 (N_18672,N_5120,N_2433);
and U18673 (N_18673,N_1659,N_6913);
nand U18674 (N_18674,N_2452,N_5110);
nand U18675 (N_18675,N_4981,N_9525);
nor U18676 (N_18676,N_5728,N_6937);
and U18677 (N_18677,N_6225,N_7095);
xnor U18678 (N_18678,N_9107,N_6369);
nor U18679 (N_18679,N_9097,N_1580);
and U18680 (N_18680,N_4154,N_880);
nor U18681 (N_18681,N_2830,N_8287);
nand U18682 (N_18682,N_3662,N_544);
and U18683 (N_18683,N_6553,N_3734);
and U18684 (N_18684,N_3064,N_9851);
nor U18685 (N_18685,N_5191,N_7650);
and U18686 (N_18686,N_6471,N_5404);
xnor U18687 (N_18687,N_8970,N_1160);
nand U18688 (N_18688,N_6672,N_5603);
nor U18689 (N_18689,N_4536,N_8778);
and U18690 (N_18690,N_5242,N_475);
or U18691 (N_18691,N_5759,N_1878);
nor U18692 (N_18692,N_7816,N_3122);
nand U18693 (N_18693,N_4643,N_9147);
and U18694 (N_18694,N_511,N_4640);
and U18695 (N_18695,N_848,N_2063);
xor U18696 (N_18696,N_3585,N_5661);
nor U18697 (N_18697,N_1731,N_8475);
xnor U18698 (N_18698,N_3478,N_988);
nor U18699 (N_18699,N_7335,N_4413);
nand U18700 (N_18700,N_6944,N_1595);
or U18701 (N_18701,N_2242,N_6952);
and U18702 (N_18702,N_8851,N_3854);
xor U18703 (N_18703,N_2558,N_4636);
nand U18704 (N_18704,N_736,N_3610);
or U18705 (N_18705,N_1336,N_4702);
nor U18706 (N_18706,N_96,N_2648);
and U18707 (N_18707,N_1593,N_5445);
or U18708 (N_18708,N_281,N_5680);
and U18709 (N_18709,N_2685,N_5021);
or U18710 (N_18710,N_5749,N_3120);
and U18711 (N_18711,N_9644,N_3064);
nor U18712 (N_18712,N_8775,N_3310);
or U18713 (N_18713,N_7511,N_643);
or U18714 (N_18714,N_3938,N_1363);
nor U18715 (N_18715,N_7936,N_7992);
nand U18716 (N_18716,N_7658,N_6637);
and U18717 (N_18717,N_3385,N_2429);
or U18718 (N_18718,N_7068,N_1237);
nor U18719 (N_18719,N_445,N_8209);
and U18720 (N_18720,N_5734,N_4022);
nand U18721 (N_18721,N_3957,N_9860);
nor U18722 (N_18722,N_6332,N_7071);
and U18723 (N_18723,N_8212,N_5245);
nand U18724 (N_18724,N_345,N_2706);
and U18725 (N_18725,N_9084,N_6296);
nor U18726 (N_18726,N_2264,N_7855);
or U18727 (N_18727,N_5849,N_9535);
or U18728 (N_18728,N_2031,N_9875);
nor U18729 (N_18729,N_9164,N_8672);
nand U18730 (N_18730,N_4016,N_5180);
or U18731 (N_18731,N_4905,N_398);
nand U18732 (N_18732,N_2464,N_5272);
nand U18733 (N_18733,N_10,N_9999);
nor U18734 (N_18734,N_8577,N_9571);
nand U18735 (N_18735,N_6488,N_4457);
and U18736 (N_18736,N_2828,N_464);
xor U18737 (N_18737,N_9615,N_8677);
nand U18738 (N_18738,N_1592,N_7961);
or U18739 (N_18739,N_1744,N_1235);
and U18740 (N_18740,N_4390,N_8887);
nor U18741 (N_18741,N_5738,N_983);
or U18742 (N_18742,N_4464,N_9749);
xnor U18743 (N_18743,N_4069,N_6624);
or U18744 (N_18744,N_4868,N_8859);
and U18745 (N_18745,N_5409,N_517);
or U18746 (N_18746,N_6202,N_5158);
nand U18747 (N_18747,N_7602,N_6013);
or U18748 (N_18748,N_4225,N_7046);
or U18749 (N_18749,N_7036,N_8997);
or U18750 (N_18750,N_560,N_3338);
nand U18751 (N_18751,N_3496,N_1710);
and U18752 (N_18752,N_9670,N_7236);
or U18753 (N_18753,N_8601,N_9088);
and U18754 (N_18754,N_3859,N_1227);
nand U18755 (N_18755,N_6266,N_2558);
or U18756 (N_18756,N_2175,N_5961);
and U18757 (N_18757,N_7009,N_9669);
nor U18758 (N_18758,N_5671,N_7768);
nand U18759 (N_18759,N_2492,N_1699);
xor U18760 (N_18760,N_8680,N_9915);
and U18761 (N_18761,N_5869,N_9800);
nor U18762 (N_18762,N_3958,N_7288);
nand U18763 (N_18763,N_6060,N_4599);
nand U18764 (N_18764,N_8644,N_4706);
xor U18765 (N_18765,N_6013,N_1445);
nand U18766 (N_18766,N_6894,N_5746);
nor U18767 (N_18767,N_239,N_6372);
xnor U18768 (N_18768,N_7021,N_1564);
nor U18769 (N_18769,N_3445,N_811);
or U18770 (N_18770,N_9732,N_5093);
or U18771 (N_18771,N_536,N_2576);
xor U18772 (N_18772,N_6475,N_4438);
nor U18773 (N_18773,N_562,N_3984);
nand U18774 (N_18774,N_8052,N_4350);
nand U18775 (N_18775,N_4101,N_7674);
or U18776 (N_18776,N_5084,N_4665);
nand U18777 (N_18777,N_8122,N_8865);
or U18778 (N_18778,N_8976,N_5054);
and U18779 (N_18779,N_9901,N_1045);
and U18780 (N_18780,N_6291,N_590);
nand U18781 (N_18781,N_231,N_4440);
and U18782 (N_18782,N_7811,N_6944);
or U18783 (N_18783,N_7539,N_84);
xor U18784 (N_18784,N_5296,N_5437);
nand U18785 (N_18785,N_3061,N_4076);
nor U18786 (N_18786,N_459,N_4112);
or U18787 (N_18787,N_5955,N_3673);
xor U18788 (N_18788,N_2987,N_6174);
nor U18789 (N_18789,N_10,N_4304);
xor U18790 (N_18790,N_5081,N_6972);
nor U18791 (N_18791,N_4368,N_2315);
xnor U18792 (N_18792,N_6805,N_2266);
nor U18793 (N_18793,N_5408,N_3709);
and U18794 (N_18794,N_9810,N_7588);
nand U18795 (N_18795,N_1792,N_1844);
nor U18796 (N_18796,N_8769,N_542);
nand U18797 (N_18797,N_4436,N_8265);
nor U18798 (N_18798,N_7480,N_977);
and U18799 (N_18799,N_1035,N_7840);
and U18800 (N_18800,N_4012,N_182);
or U18801 (N_18801,N_6096,N_381);
nor U18802 (N_18802,N_8781,N_4683);
and U18803 (N_18803,N_6326,N_5770);
nor U18804 (N_18804,N_7858,N_9860);
and U18805 (N_18805,N_220,N_7826);
nor U18806 (N_18806,N_6430,N_5419);
nor U18807 (N_18807,N_6302,N_2442);
nand U18808 (N_18808,N_7785,N_672);
or U18809 (N_18809,N_6640,N_8351);
xor U18810 (N_18810,N_5689,N_9454);
nor U18811 (N_18811,N_3272,N_8361);
xor U18812 (N_18812,N_5370,N_6233);
nor U18813 (N_18813,N_381,N_1443);
and U18814 (N_18814,N_338,N_9565);
xnor U18815 (N_18815,N_1330,N_5917);
nor U18816 (N_18816,N_9667,N_998);
nor U18817 (N_18817,N_5428,N_5936);
nand U18818 (N_18818,N_9962,N_212);
xnor U18819 (N_18819,N_7757,N_118);
or U18820 (N_18820,N_9711,N_1176);
or U18821 (N_18821,N_5800,N_3187);
nor U18822 (N_18822,N_5246,N_5336);
nor U18823 (N_18823,N_9478,N_7104);
nand U18824 (N_18824,N_6668,N_9994);
and U18825 (N_18825,N_5751,N_8036);
and U18826 (N_18826,N_6499,N_4754);
or U18827 (N_18827,N_8024,N_1723);
nor U18828 (N_18828,N_9621,N_9958);
or U18829 (N_18829,N_2238,N_3469);
or U18830 (N_18830,N_1709,N_2532);
xor U18831 (N_18831,N_5093,N_2149);
and U18832 (N_18832,N_1235,N_1182);
nand U18833 (N_18833,N_7224,N_3747);
nor U18834 (N_18834,N_1208,N_6718);
nand U18835 (N_18835,N_1489,N_42);
nand U18836 (N_18836,N_8162,N_4681);
or U18837 (N_18837,N_7778,N_7673);
or U18838 (N_18838,N_8559,N_8587);
nor U18839 (N_18839,N_3833,N_8963);
nor U18840 (N_18840,N_8301,N_8081);
nor U18841 (N_18841,N_6477,N_7983);
or U18842 (N_18842,N_8224,N_7151);
nor U18843 (N_18843,N_7707,N_6899);
or U18844 (N_18844,N_3435,N_6482);
nand U18845 (N_18845,N_3352,N_720);
or U18846 (N_18846,N_4827,N_7110);
nand U18847 (N_18847,N_3300,N_6427);
or U18848 (N_18848,N_3637,N_433);
nor U18849 (N_18849,N_8581,N_3479);
xnor U18850 (N_18850,N_1339,N_3395);
and U18851 (N_18851,N_9825,N_2802);
xnor U18852 (N_18852,N_5193,N_8611);
nand U18853 (N_18853,N_7699,N_7817);
xnor U18854 (N_18854,N_1167,N_8657);
nand U18855 (N_18855,N_5960,N_3509);
and U18856 (N_18856,N_9275,N_4671);
or U18857 (N_18857,N_4288,N_7878);
and U18858 (N_18858,N_5697,N_3932);
and U18859 (N_18859,N_896,N_9191);
nor U18860 (N_18860,N_5609,N_4657);
xnor U18861 (N_18861,N_4335,N_7584);
nor U18862 (N_18862,N_1045,N_4263);
nand U18863 (N_18863,N_7308,N_6720);
and U18864 (N_18864,N_5116,N_9476);
nor U18865 (N_18865,N_587,N_6375);
nand U18866 (N_18866,N_3495,N_711);
or U18867 (N_18867,N_403,N_7996);
and U18868 (N_18868,N_1558,N_2161);
xnor U18869 (N_18869,N_8772,N_9065);
xor U18870 (N_18870,N_6812,N_3573);
and U18871 (N_18871,N_3876,N_5265);
and U18872 (N_18872,N_5911,N_6805);
or U18873 (N_18873,N_702,N_8039);
or U18874 (N_18874,N_6231,N_8160);
and U18875 (N_18875,N_6401,N_3610);
or U18876 (N_18876,N_3235,N_2712);
nor U18877 (N_18877,N_5849,N_2003);
nand U18878 (N_18878,N_6245,N_519);
nor U18879 (N_18879,N_8469,N_7613);
xor U18880 (N_18880,N_6762,N_7891);
nor U18881 (N_18881,N_7193,N_1440);
xor U18882 (N_18882,N_1351,N_2597);
or U18883 (N_18883,N_2831,N_5392);
or U18884 (N_18884,N_1679,N_3168);
nor U18885 (N_18885,N_2146,N_7276);
nor U18886 (N_18886,N_9121,N_3325);
or U18887 (N_18887,N_9838,N_4295);
nor U18888 (N_18888,N_8333,N_5405);
and U18889 (N_18889,N_9638,N_8298);
or U18890 (N_18890,N_9668,N_714);
nand U18891 (N_18891,N_383,N_9338);
nor U18892 (N_18892,N_8589,N_6566);
nand U18893 (N_18893,N_9506,N_4511);
nor U18894 (N_18894,N_1646,N_7284);
nand U18895 (N_18895,N_2210,N_8533);
nor U18896 (N_18896,N_6453,N_6601);
or U18897 (N_18897,N_4384,N_9286);
nand U18898 (N_18898,N_4058,N_1847);
nand U18899 (N_18899,N_9257,N_9685);
and U18900 (N_18900,N_8038,N_9501);
xnor U18901 (N_18901,N_111,N_5830);
or U18902 (N_18902,N_8139,N_5334);
or U18903 (N_18903,N_3998,N_8644);
nand U18904 (N_18904,N_9797,N_7324);
and U18905 (N_18905,N_1112,N_8706);
and U18906 (N_18906,N_2655,N_1583);
nand U18907 (N_18907,N_1520,N_1621);
nand U18908 (N_18908,N_7131,N_96);
nand U18909 (N_18909,N_7851,N_8507);
nand U18910 (N_18910,N_1253,N_6576);
or U18911 (N_18911,N_6295,N_507);
or U18912 (N_18912,N_4447,N_807);
or U18913 (N_18913,N_4986,N_2192);
nand U18914 (N_18914,N_5225,N_5933);
nand U18915 (N_18915,N_1460,N_5442);
and U18916 (N_18916,N_3661,N_8999);
nand U18917 (N_18917,N_6826,N_6457);
nand U18918 (N_18918,N_7491,N_2842);
or U18919 (N_18919,N_1949,N_2350);
nand U18920 (N_18920,N_2534,N_1546);
xor U18921 (N_18921,N_7625,N_5112);
xnor U18922 (N_18922,N_2718,N_5175);
and U18923 (N_18923,N_4199,N_437);
nand U18924 (N_18924,N_2950,N_3187);
or U18925 (N_18925,N_1958,N_3088);
nor U18926 (N_18926,N_8503,N_166);
nand U18927 (N_18927,N_985,N_7404);
and U18928 (N_18928,N_7744,N_8846);
nand U18929 (N_18929,N_5399,N_1175);
or U18930 (N_18930,N_5708,N_5747);
nand U18931 (N_18931,N_1381,N_6659);
xnor U18932 (N_18932,N_7025,N_47);
nor U18933 (N_18933,N_7624,N_2292);
or U18934 (N_18934,N_1592,N_5194);
nand U18935 (N_18935,N_6963,N_3963);
nand U18936 (N_18936,N_4193,N_1270);
and U18937 (N_18937,N_7816,N_6971);
and U18938 (N_18938,N_794,N_1353);
nand U18939 (N_18939,N_8323,N_2399);
and U18940 (N_18940,N_893,N_1603);
nand U18941 (N_18941,N_8668,N_128);
and U18942 (N_18942,N_3979,N_2133);
or U18943 (N_18943,N_757,N_8854);
nand U18944 (N_18944,N_553,N_1016);
or U18945 (N_18945,N_2523,N_4515);
nor U18946 (N_18946,N_6923,N_4179);
and U18947 (N_18947,N_5734,N_7067);
xnor U18948 (N_18948,N_999,N_3083);
and U18949 (N_18949,N_1336,N_2094);
nor U18950 (N_18950,N_8628,N_8232);
nor U18951 (N_18951,N_8942,N_1257);
nand U18952 (N_18952,N_7908,N_905);
and U18953 (N_18953,N_7321,N_1904);
and U18954 (N_18954,N_8292,N_9976);
and U18955 (N_18955,N_9682,N_3208);
nand U18956 (N_18956,N_3963,N_8303);
nor U18957 (N_18957,N_9519,N_257);
and U18958 (N_18958,N_1843,N_3696);
and U18959 (N_18959,N_5880,N_6688);
or U18960 (N_18960,N_8945,N_2073);
or U18961 (N_18961,N_3967,N_3198);
and U18962 (N_18962,N_1095,N_5866);
or U18963 (N_18963,N_7099,N_7265);
nor U18964 (N_18964,N_2842,N_5813);
nor U18965 (N_18965,N_7475,N_3208);
and U18966 (N_18966,N_9747,N_5036);
and U18967 (N_18967,N_9581,N_1538);
nand U18968 (N_18968,N_4002,N_9523);
nand U18969 (N_18969,N_5090,N_7340);
or U18970 (N_18970,N_4471,N_2374);
or U18971 (N_18971,N_1956,N_1554);
xor U18972 (N_18972,N_3591,N_5170);
and U18973 (N_18973,N_2589,N_8073);
and U18974 (N_18974,N_3697,N_2791);
nor U18975 (N_18975,N_6154,N_6007);
or U18976 (N_18976,N_2795,N_9861);
nand U18977 (N_18977,N_2276,N_1490);
or U18978 (N_18978,N_3327,N_6478);
nand U18979 (N_18979,N_2065,N_6512);
or U18980 (N_18980,N_3554,N_9232);
nand U18981 (N_18981,N_5498,N_7459);
xnor U18982 (N_18982,N_9894,N_6970);
nor U18983 (N_18983,N_2478,N_5466);
and U18984 (N_18984,N_2290,N_4148);
nor U18985 (N_18985,N_3721,N_3830);
and U18986 (N_18986,N_6799,N_7691);
nand U18987 (N_18987,N_5362,N_5519);
nor U18988 (N_18988,N_9371,N_1614);
nand U18989 (N_18989,N_8946,N_1785);
nor U18990 (N_18990,N_698,N_2198);
nand U18991 (N_18991,N_90,N_4763);
nor U18992 (N_18992,N_8181,N_5089);
nand U18993 (N_18993,N_5510,N_4778);
nand U18994 (N_18994,N_29,N_467);
or U18995 (N_18995,N_7366,N_9888);
nand U18996 (N_18996,N_5475,N_5748);
xor U18997 (N_18997,N_2161,N_9613);
and U18998 (N_18998,N_2447,N_7509);
xnor U18999 (N_18999,N_1512,N_3967);
and U19000 (N_19000,N_4542,N_1319);
or U19001 (N_19001,N_6893,N_8212);
nand U19002 (N_19002,N_7383,N_5222);
xnor U19003 (N_19003,N_646,N_1780);
and U19004 (N_19004,N_8326,N_5739);
nor U19005 (N_19005,N_2467,N_8540);
and U19006 (N_19006,N_4052,N_261);
or U19007 (N_19007,N_219,N_3851);
nor U19008 (N_19008,N_9376,N_8546);
or U19009 (N_19009,N_2007,N_7257);
nand U19010 (N_19010,N_8894,N_3828);
and U19011 (N_19011,N_8930,N_4499);
and U19012 (N_19012,N_8901,N_7328);
nor U19013 (N_19013,N_9891,N_4557);
nand U19014 (N_19014,N_8593,N_1080);
or U19015 (N_19015,N_2553,N_6018);
and U19016 (N_19016,N_5299,N_6349);
nand U19017 (N_19017,N_9444,N_4053);
nand U19018 (N_19018,N_7596,N_5338);
nand U19019 (N_19019,N_5814,N_1502);
nor U19020 (N_19020,N_5130,N_1977);
nand U19021 (N_19021,N_9152,N_8741);
nand U19022 (N_19022,N_3826,N_2049);
xor U19023 (N_19023,N_4248,N_8427);
or U19024 (N_19024,N_3050,N_9319);
and U19025 (N_19025,N_6445,N_1848);
nor U19026 (N_19026,N_8642,N_17);
xnor U19027 (N_19027,N_8226,N_3960);
nand U19028 (N_19028,N_2432,N_1127);
xor U19029 (N_19029,N_23,N_9897);
or U19030 (N_19030,N_3808,N_9479);
and U19031 (N_19031,N_4108,N_5392);
and U19032 (N_19032,N_8917,N_2266);
xnor U19033 (N_19033,N_811,N_6710);
or U19034 (N_19034,N_2075,N_6686);
nor U19035 (N_19035,N_1355,N_2166);
nand U19036 (N_19036,N_5942,N_467);
or U19037 (N_19037,N_392,N_9197);
or U19038 (N_19038,N_8982,N_8011);
or U19039 (N_19039,N_23,N_6080);
and U19040 (N_19040,N_7305,N_8177);
and U19041 (N_19041,N_9169,N_2960);
and U19042 (N_19042,N_262,N_9923);
or U19043 (N_19043,N_3307,N_8639);
or U19044 (N_19044,N_9830,N_5582);
xnor U19045 (N_19045,N_5710,N_6001);
nor U19046 (N_19046,N_7774,N_2990);
or U19047 (N_19047,N_9809,N_6506);
nand U19048 (N_19048,N_9757,N_9584);
and U19049 (N_19049,N_8052,N_3068);
xnor U19050 (N_19050,N_9159,N_576);
or U19051 (N_19051,N_1316,N_4826);
nand U19052 (N_19052,N_112,N_3329);
nor U19053 (N_19053,N_653,N_1674);
or U19054 (N_19054,N_6963,N_8287);
and U19055 (N_19055,N_2212,N_2230);
nand U19056 (N_19056,N_9576,N_35);
and U19057 (N_19057,N_2381,N_1031);
or U19058 (N_19058,N_7548,N_8431);
nor U19059 (N_19059,N_9051,N_2145);
or U19060 (N_19060,N_5794,N_5508);
and U19061 (N_19061,N_6778,N_4193);
nor U19062 (N_19062,N_4742,N_1114);
nor U19063 (N_19063,N_4620,N_3632);
nand U19064 (N_19064,N_8295,N_7875);
nor U19065 (N_19065,N_6015,N_9442);
or U19066 (N_19066,N_2605,N_1385);
nand U19067 (N_19067,N_90,N_6878);
or U19068 (N_19068,N_1734,N_9245);
nor U19069 (N_19069,N_813,N_4486);
or U19070 (N_19070,N_9355,N_9149);
nor U19071 (N_19071,N_6891,N_7156);
nor U19072 (N_19072,N_5217,N_3174);
nand U19073 (N_19073,N_9471,N_2353);
nand U19074 (N_19074,N_7240,N_4889);
nand U19075 (N_19075,N_8656,N_4453);
nor U19076 (N_19076,N_6207,N_330);
and U19077 (N_19077,N_9420,N_4369);
nand U19078 (N_19078,N_386,N_1374);
nand U19079 (N_19079,N_5858,N_5137);
nand U19080 (N_19080,N_7791,N_4487);
or U19081 (N_19081,N_2677,N_5806);
and U19082 (N_19082,N_2380,N_7946);
nand U19083 (N_19083,N_6031,N_7692);
and U19084 (N_19084,N_2124,N_5407);
or U19085 (N_19085,N_6026,N_3919);
or U19086 (N_19086,N_4164,N_8482);
or U19087 (N_19087,N_1748,N_2172);
nand U19088 (N_19088,N_1906,N_2881);
and U19089 (N_19089,N_6891,N_8607);
or U19090 (N_19090,N_844,N_9895);
nand U19091 (N_19091,N_6368,N_9613);
or U19092 (N_19092,N_662,N_1788);
or U19093 (N_19093,N_6863,N_117);
or U19094 (N_19094,N_9583,N_285);
nand U19095 (N_19095,N_6824,N_4331);
and U19096 (N_19096,N_2093,N_1048);
nor U19097 (N_19097,N_3021,N_373);
nor U19098 (N_19098,N_1582,N_4587);
and U19099 (N_19099,N_1189,N_2710);
and U19100 (N_19100,N_6950,N_3129);
and U19101 (N_19101,N_9630,N_2714);
and U19102 (N_19102,N_6903,N_1754);
nor U19103 (N_19103,N_7487,N_5038);
nand U19104 (N_19104,N_8465,N_1036);
nor U19105 (N_19105,N_7356,N_3340);
nor U19106 (N_19106,N_6156,N_1918);
nor U19107 (N_19107,N_4151,N_341);
or U19108 (N_19108,N_4296,N_9403);
or U19109 (N_19109,N_9234,N_4483);
nor U19110 (N_19110,N_7770,N_8997);
nor U19111 (N_19111,N_6947,N_8100);
or U19112 (N_19112,N_5986,N_5495);
xor U19113 (N_19113,N_2828,N_9609);
nor U19114 (N_19114,N_7,N_7343);
nor U19115 (N_19115,N_5892,N_1787);
or U19116 (N_19116,N_9504,N_8631);
nand U19117 (N_19117,N_2658,N_4868);
nor U19118 (N_19118,N_4497,N_5650);
nor U19119 (N_19119,N_8209,N_4050);
nand U19120 (N_19120,N_6157,N_8581);
nand U19121 (N_19121,N_3928,N_7144);
nor U19122 (N_19122,N_9415,N_4920);
nand U19123 (N_19123,N_1414,N_14);
and U19124 (N_19124,N_2244,N_4077);
and U19125 (N_19125,N_6033,N_350);
or U19126 (N_19126,N_6273,N_5717);
nor U19127 (N_19127,N_3095,N_3221);
nor U19128 (N_19128,N_9214,N_1225);
or U19129 (N_19129,N_6988,N_8048);
nor U19130 (N_19130,N_4444,N_8465);
and U19131 (N_19131,N_4664,N_3199);
nand U19132 (N_19132,N_1390,N_5877);
nor U19133 (N_19133,N_9393,N_755);
or U19134 (N_19134,N_1427,N_1559);
nor U19135 (N_19135,N_3356,N_329);
nor U19136 (N_19136,N_8393,N_8967);
nand U19137 (N_19137,N_5054,N_3147);
or U19138 (N_19138,N_1012,N_6471);
nor U19139 (N_19139,N_9869,N_3976);
or U19140 (N_19140,N_2701,N_1524);
nor U19141 (N_19141,N_7521,N_5104);
or U19142 (N_19142,N_7085,N_8696);
or U19143 (N_19143,N_9380,N_851);
or U19144 (N_19144,N_7937,N_6253);
nor U19145 (N_19145,N_9037,N_1973);
nand U19146 (N_19146,N_1906,N_3181);
or U19147 (N_19147,N_2659,N_5139);
xor U19148 (N_19148,N_1581,N_3745);
or U19149 (N_19149,N_6267,N_3505);
and U19150 (N_19150,N_6591,N_4460);
nand U19151 (N_19151,N_4760,N_5612);
or U19152 (N_19152,N_7409,N_7760);
or U19153 (N_19153,N_1252,N_2508);
and U19154 (N_19154,N_4654,N_7163);
or U19155 (N_19155,N_5630,N_6246);
and U19156 (N_19156,N_8500,N_6533);
xor U19157 (N_19157,N_7536,N_5481);
and U19158 (N_19158,N_5941,N_9274);
and U19159 (N_19159,N_6481,N_9158);
and U19160 (N_19160,N_3607,N_8119);
and U19161 (N_19161,N_9747,N_4414);
nor U19162 (N_19162,N_4682,N_757);
nand U19163 (N_19163,N_7319,N_4626);
nand U19164 (N_19164,N_1449,N_1783);
or U19165 (N_19165,N_5487,N_6560);
and U19166 (N_19166,N_6468,N_8556);
nor U19167 (N_19167,N_9925,N_4417);
xor U19168 (N_19168,N_3388,N_8327);
and U19169 (N_19169,N_4765,N_4091);
or U19170 (N_19170,N_317,N_5565);
or U19171 (N_19171,N_3169,N_435);
nand U19172 (N_19172,N_5015,N_1718);
nor U19173 (N_19173,N_6853,N_7504);
nand U19174 (N_19174,N_2149,N_2336);
or U19175 (N_19175,N_8968,N_9181);
or U19176 (N_19176,N_2613,N_8281);
nor U19177 (N_19177,N_387,N_963);
and U19178 (N_19178,N_5546,N_5733);
or U19179 (N_19179,N_2614,N_768);
nand U19180 (N_19180,N_4169,N_8995);
and U19181 (N_19181,N_5820,N_4158);
and U19182 (N_19182,N_4120,N_373);
xor U19183 (N_19183,N_2054,N_7414);
or U19184 (N_19184,N_1040,N_2569);
nand U19185 (N_19185,N_8778,N_7878);
nand U19186 (N_19186,N_7205,N_3413);
and U19187 (N_19187,N_3248,N_9610);
nor U19188 (N_19188,N_2217,N_5589);
nand U19189 (N_19189,N_5487,N_1932);
or U19190 (N_19190,N_4775,N_2594);
nand U19191 (N_19191,N_6106,N_6756);
and U19192 (N_19192,N_875,N_6604);
nor U19193 (N_19193,N_7451,N_9621);
nand U19194 (N_19194,N_2715,N_2115);
and U19195 (N_19195,N_5846,N_3672);
xor U19196 (N_19196,N_1226,N_3045);
nor U19197 (N_19197,N_8013,N_4412);
nand U19198 (N_19198,N_5421,N_7947);
nor U19199 (N_19199,N_894,N_3946);
nand U19200 (N_19200,N_2223,N_3567);
and U19201 (N_19201,N_1488,N_1685);
nor U19202 (N_19202,N_9152,N_3927);
nor U19203 (N_19203,N_2597,N_8292);
or U19204 (N_19204,N_7724,N_1128);
nand U19205 (N_19205,N_9750,N_5772);
and U19206 (N_19206,N_7028,N_8328);
and U19207 (N_19207,N_9188,N_1000);
or U19208 (N_19208,N_6159,N_4746);
or U19209 (N_19209,N_2938,N_9448);
nor U19210 (N_19210,N_4191,N_5983);
or U19211 (N_19211,N_1576,N_106);
and U19212 (N_19212,N_6103,N_2004);
nor U19213 (N_19213,N_3465,N_3161);
or U19214 (N_19214,N_3668,N_3667);
xnor U19215 (N_19215,N_9441,N_1929);
and U19216 (N_19216,N_8036,N_2373);
nand U19217 (N_19217,N_5896,N_8292);
nor U19218 (N_19218,N_0,N_8793);
nor U19219 (N_19219,N_8280,N_627);
or U19220 (N_19220,N_2577,N_2517);
nand U19221 (N_19221,N_8136,N_2833);
and U19222 (N_19222,N_4118,N_3060);
or U19223 (N_19223,N_3258,N_3236);
xnor U19224 (N_19224,N_6258,N_7619);
xor U19225 (N_19225,N_2251,N_434);
or U19226 (N_19226,N_1861,N_9226);
and U19227 (N_19227,N_4628,N_1933);
or U19228 (N_19228,N_5962,N_5113);
or U19229 (N_19229,N_1494,N_3716);
or U19230 (N_19230,N_7904,N_1714);
nand U19231 (N_19231,N_4096,N_7144);
nand U19232 (N_19232,N_22,N_5093);
or U19233 (N_19233,N_6748,N_5348);
nor U19234 (N_19234,N_5059,N_3878);
nand U19235 (N_19235,N_676,N_6800);
and U19236 (N_19236,N_8567,N_9973);
and U19237 (N_19237,N_959,N_3494);
and U19238 (N_19238,N_2562,N_5664);
nand U19239 (N_19239,N_6686,N_4962);
or U19240 (N_19240,N_7395,N_8878);
nor U19241 (N_19241,N_3183,N_8969);
nand U19242 (N_19242,N_9072,N_6794);
nor U19243 (N_19243,N_5734,N_5212);
nor U19244 (N_19244,N_9513,N_2726);
or U19245 (N_19245,N_449,N_3932);
and U19246 (N_19246,N_351,N_8750);
or U19247 (N_19247,N_2568,N_6777);
nand U19248 (N_19248,N_4913,N_5720);
nand U19249 (N_19249,N_5964,N_8399);
xnor U19250 (N_19250,N_1776,N_8509);
nand U19251 (N_19251,N_4843,N_4758);
xor U19252 (N_19252,N_9366,N_8172);
nor U19253 (N_19253,N_7485,N_3875);
and U19254 (N_19254,N_111,N_2450);
xor U19255 (N_19255,N_3525,N_994);
nor U19256 (N_19256,N_4378,N_7086);
nand U19257 (N_19257,N_8722,N_7993);
nand U19258 (N_19258,N_3591,N_921);
or U19259 (N_19259,N_1818,N_4882);
nand U19260 (N_19260,N_9042,N_413);
or U19261 (N_19261,N_4996,N_2992);
and U19262 (N_19262,N_9811,N_6320);
and U19263 (N_19263,N_8192,N_8198);
nor U19264 (N_19264,N_9484,N_2425);
and U19265 (N_19265,N_442,N_2381);
nand U19266 (N_19266,N_209,N_5664);
or U19267 (N_19267,N_8850,N_8604);
xnor U19268 (N_19268,N_9049,N_3245);
xnor U19269 (N_19269,N_8977,N_3202);
nand U19270 (N_19270,N_6760,N_8313);
nand U19271 (N_19271,N_8443,N_9244);
nand U19272 (N_19272,N_3888,N_7280);
nand U19273 (N_19273,N_6528,N_4406);
nand U19274 (N_19274,N_7061,N_6344);
nand U19275 (N_19275,N_5842,N_2221);
and U19276 (N_19276,N_2505,N_2988);
nor U19277 (N_19277,N_2211,N_7387);
nand U19278 (N_19278,N_8043,N_8320);
and U19279 (N_19279,N_614,N_3747);
nand U19280 (N_19280,N_3016,N_5822);
and U19281 (N_19281,N_3922,N_4984);
nor U19282 (N_19282,N_2659,N_1050);
xnor U19283 (N_19283,N_8997,N_2832);
xnor U19284 (N_19284,N_2178,N_6810);
or U19285 (N_19285,N_1665,N_6920);
nand U19286 (N_19286,N_4261,N_3508);
or U19287 (N_19287,N_5800,N_7794);
nand U19288 (N_19288,N_6041,N_3166);
and U19289 (N_19289,N_152,N_7614);
nor U19290 (N_19290,N_5964,N_1348);
nand U19291 (N_19291,N_8635,N_8090);
nand U19292 (N_19292,N_6061,N_6913);
nand U19293 (N_19293,N_4258,N_3525);
nand U19294 (N_19294,N_4762,N_1774);
xnor U19295 (N_19295,N_7996,N_1259);
and U19296 (N_19296,N_7329,N_7315);
nor U19297 (N_19297,N_5713,N_560);
or U19298 (N_19298,N_4561,N_7121);
nor U19299 (N_19299,N_5712,N_1168);
or U19300 (N_19300,N_9313,N_6547);
nor U19301 (N_19301,N_2171,N_5342);
or U19302 (N_19302,N_8077,N_5505);
and U19303 (N_19303,N_6464,N_7735);
or U19304 (N_19304,N_7453,N_2155);
and U19305 (N_19305,N_2001,N_4965);
or U19306 (N_19306,N_560,N_9334);
nor U19307 (N_19307,N_3740,N_3863);
nand U19308 (N_19308,N_8750,N_5100);
nor U19309 (N_19309,N_8141,N_5680);
xor U19310 (N_19310,N_4282,N_9242);
or U19311 (N_19311,N_260,N_486);
and U19312 (N_19312,N_7152,N_7242);
nor U19313 (N_19313,N_8703,N_6456);
and U19314 (N_19314,N_9779,N_922);
nor U19315 (N_19315,N_6250,N_9042);
and U19316 (N_19316,N_254,N_6284);
or U19317 (N_19317,N_9065,N_2362);
nand U19318 (N_19318,N_3088,N_9861);
nor U19319 (N_19319,N_6532,N_494);
or U19320 (N_19320,N_2448,N_9681);
or U19321 (N_19321,N_991,N_9117);
xnor U19322 (N_19322,N_7524,N_2349);
nand U19323 (N_19323,N_6487,N_6147);
nand U19324 (N_19324,N_6289,N_2186);
nand U19325 (N_19325,N_128,N_4104);
nand U19326 (N_19326,N_1820,N_7643);
and U19327 (N_19327,N_9280,N_9973);
nand U19328 (N_19328,N_2603,N_905);
nor U19329 (N_19329,N_4912,N_7195);
and U19330 (N_19330,N_3270,N_6926);
and U19331 (N_19331,N_4345,N_8434);
nor U19332 (N_19332,N_9822,N_8504);
or U19333 (N_19333,N_337,N_7924);
or U19334 (N_19334,N_6388,N_8648);
nor U19335 (N_19335,N_7670,N_5351);
and U19336 (N_19336,N_100,N_2486);
or U19337 (N_19337,N_492,N_7119);
or U19338 (N_19338,N_1392,N_852);
or U19339 (N_19339,N_2630,N_9668);
and U19340 (N_19340,N_4760,N_3457);
nand U19341 (N_19341,N_3950,N_7140);
or U19342 (N_19342,N_3492,N_7108);
and U19343 (N_19343,N_2518,N_2456);
and U19344 (N_19344,N_5497,N_3922);
nor U19345 (N_19345,N_9402,N_3844);
and U19346 (N_19346,N_5267,N_1436);
or U19347 (N_19347,N_4038,N_4892);
or U19348 (N_19348,N_1572,N_8775);
nor U19349 (N_19349,N_982,N_3285);
xor U19350 (N_19350,N_3371,N_1513);
nand U19351 (N_19351,N_6839,N_4872);
nor U19352 (N_19352,N_8718,N_1230);
nor U19353 (N_19353,N_5852,N_6736);
xor U19354 (N_19354,N_2513,N_643);
or U19355 (N_19355,N_9707,N_4701);
nor U19356 (N_19356,N_3924,N_4359);
nand U19357 (N_19357,N_5450,N_6692);
and U19358 (N_19358,N_4783,N_249);
and U19359 (N_19359,N_5711,N_1189);
xor U19360 (N_19360,N_3522,N_1673);
nor U19361 (N_19361,N_7805,N_5403);
or U19362 (N_19362,N_3349,N_9975);
nor U19363 (N_19363,N_5086,N_452);
or U19364 (N_19364,N_2007,N_7210);
and U19365 (N_19365,N_9173,N_2991);
and U19366 (N_19366,N_4412,N_6409);
nand U19367 (N_19367,N_9124,N_4729);
and U19368 (N_19368,N_1610,N_4799);
and U19369 (N_19369,N_1098,N_6433);
and U19370 (N_19370,N_9552,N_5221);
xnor U19371 (N_19371,N_7967,N_5976);
nor U19372 (N_19372,N_233,N_4400);
nand U19373 (N_19373,N_2237,N_3524);
nor U19374 (N_19374,N_6644,N_7602);
xor U19375 (N_19375,N_5698,N_7118);
or U19376 (N_19376,N_9364,N_4647);
nand U19377 (N_19377,N_3048,N_718);
or U19378 (N_19378,N_4597,N_802);
nand U19379 (N_19379,N_8197,N_7087);
or U19380 (N_19380,N_3978,N_7025);
xnor U19381 (N_19381,N_5708,N_7453);
or U19382 (N_19382,N_5303,N_1855);
nor U19383 (N_19383,N_1290,N_4969);
nand U19384 (N_19384,N_4815,N_5994);
and U19385 (N_19385,N_7716,N_7383);
nor U19386 (N_19386,N_5826,N_7075);
nor U19387 (N_19387,N_3309,N_2027);
and U19388 (N_19388,N_603,N_9449);
or U19389 (N_19389,N_4565,N_2210);
nand U19390 (N_19390,N_6002,N_4015);
nand U19391 (N_19391,N_6519,N_5444);
nor U19392 (N_19392,N_7667,N_1553);
and U19393 (N_19393,N_4143,N_6871);
and U19394 (N_19394,N_7270,N_8976);
or U19395 (N_19395,N_1450,N_6761);
or U19396 (N_19396,N_9108,N_5310);
or U19397 (N_19397,N_845,N_1587);
and U19398 (N_19398,N_6649,N_4857);
or U19399 (N_19399,N_9186,N_8244);
nor U19400 (N_19400,N_8160,N_4115);
or U19401 (N_19401,N_3567,N_7359);
or U19402 (N_19402,N_7321,N_1011);
and U19403 (N_19403,N_4027,N_9589);
or U19404 (N_19404,N_563,N_572);
nor U19405 (N_19405,N_8724,N_5995);
nor U19406 (N_19406,N_3378,N_8346);
or U19407 (N_19407,N_278,N_5270);
and U19408 (N_19408,N_7462,N_4575);
or U19409 (N_19409,N_5248,N_1664);
nand U19410 (N_19410,N_6775,N_3729);
or U19411 (N_19411,N_950,N_4476);
and U19412 (N_19412,N_6907,N_6063);
and U19413 (N_19413,N_3353,N_5614);
nor U19414 (N_19414,N_8303,N_4872);
or U19415 (N_19415,N_4775,N_5184);
and U19416 (N_19416,N_261,N_2058);
and U19417 (N_19417,N_8912,N_2976);
and U19418 (N_19418,N_9579,N_9754);
nand U19419 (N_19419,N_1204,N_4316);
and U19420 (N_19420,N_4722,N_5651);
nor U19421 (N_19421,N_745,N_7681);
and U19422 (N_19422,N_908,N_3177);
or U19423 (N_19423,N_915,N_8873);
nand U19424 (N_19424,N_5422,N_9705);
and U19425 (N_19425,N_3881,N_4423);
or U19426 (N_19426,N_4744,N_9955);
and U19427 (N_19427,N_6045,N_3920);
nor U19428 (N_19428,N_2054,N_8737);
nand U19429 (N_19429,N_112,N_6832);
nor U19430 (N_19430,N_3350,N_6033);
and U19431 (N_19431,N_5519,N_4371);
or U19432 (N_19432,N_2240,N_6238);
and U19433 (N_19433,N_1772,N_918);
and U19434 (N_19434,N_8921,N_7258);
xnor U19435 (N_19435,N_4308,N_2266);
and U19436 (N_19436,N_4270,N_3998);
or U19437 (N_19437,N_7802,N_6418);
and U19438 (N_19438,N_9558,N_3007);
nand U19439 (N_19439,N_2808,N_9830);
nor U19440 (N_19440,N_9206,N_8052);
and U19441 (N_19441,N_722,N_4987);
or U19442 (N_19442,N_5456,N_4736);
and U19443 (N_19443,N_3751,N_1359);
nor U19444 (N_19444,N_7843,N_433);
nor U19445 (N_19445,N_6814,N_7261);
nand U19446 (N_19446,N_5332,N_8091);
or U19447 (N_19447,N_5569,N_9822);
or U19448 (N_19448,N_7430,N_4752);
nor U19449 (N_19449,N_2352,N_1651);
nor U19450 (N_19450,N_8680,N_701);
nand U19451 (N_19451,N_5171,N_8224);
and U19452 (N_19452,N_316,N_4003);
nor U19453 (N_19453,N_9226,N_7818);
or U19454 (N_19454,N_8561,N_2872);
and U19455 (N_19455,N_9198,N_7915);
nand U19456 (N_19456,N_7244,N_8961);
or U19457 (N_19457,N_8291,N_1749);
and U19458 (N_19458,N_7240,N_8157);
nand U19459 (N_19459,N_6102,N_3607);
or U19460 (N_19460,N_245,N_8411);
xnor U19461 (N_19461,N_1024,N_9651);
or U19462 (N_19462,N_306,N_1972);
and U19463 (N_19463,N_8899,N_800);
or U19464 (N_19464,N_4685,N_9249);
and U19465 (N_19465,N_845,N_9123);
xnor U19466 (N_19466,N_5208,N_8486);
and U19467 (N_19467,N_3847,N_2121);
or U19468 (N_19468,N_2342,N_6492);
or U19469 (N_19469,N_2639,N_343);
nor U19470 (N_19470,N_3447,N_2957);
nand U19471 (N_19471,N_7527,N_6869);
xnor U19472 (N_19472,N_4965,N_9237);
nand U19473 (N_19473,N_2457,N_6687);
nor U19474 (N_19474,N_3461,N_729);
and U19475 (N_19475,N_818,N_1253);
xor U19476 (N_19476,N_9687,N_9870);
nor U19477 (N_19477,N_922,N_7152);
or U19478 (N_19478,N_6412,N_1871);
xor U19479 (N_19479,N_7035,N_9366);
or U19480 (N_19480,N_3487,N_6267);
and U19481 (N_19481,N_6168,N_1339);
or U19482 (N_19482,N_6889,N_1310);
nor U19483 (N_19483,N_6912,N_3775);
and U19484 (N_19484,N_1188,N_9656);
nand U19485 (N_19485,N_1169,N_9033);
and U19486 (N_19486,N_1525,N_7888);
nor U19487 (N_19487,N_3254,N_5457);
nand U19488 (N_19488,N_1814,N_2390);
nand U19489 (N_19489,N_2268,N_8655);
xor U19490 (N_19490,N_5073,N_9597);
nor U19491 (N_19491,N_7474,N_4009);
and U19492 (N_19492,N_9214,N_2418);
and U19493 (N_19493,N_8997,N_1290);
nor U19494 (N_19494,N_1056,N_746);
nand U19495 (N_19495,N_7885,N_6300);
or U19496 (N_19496,N_9960,N_7585);
nand U19497 (N_19497,N_904,N_6151);
nor U19498 (N_19498,N_4053,N_5757);
nor U19499 (N_19499,N_8548,N_9467);
nand U19500 (N_19500,N_6909,N_677);
and U19501 (N_19501,N_7204,N_2087);
nor U19502 (N_19502,N_4857,N_8878);
xor U19503 (N_19503,N_7152,N_5412);
nand U19504 (N_19504,N_8220,N_6561);
nand U19505 (N_19505,N_8395,N_6398);
or U19506 (N_19506,N_5362,N_4899);
nand U19507 (N_19507,N_5922,N_6839);
or U19508 (N_19508,N_5122,N_7319);
nor U19509 (N_19509,N_4859,N_9214);
xnor U19510 (N_19510,N_9587,N_4764);
and U19511 (N_19511,N_7550,N_567);
and U19512 (N_19512,N_9232,N_6864);
nor U19513 (N_19513,N_5006,N_7679);
and U19514 (N_19514,N_2818,N_3689);
nor U19515 (N_19515,N_3851,N_2881);
xor U19516 (N_19516,N_522,N_9034);
and U19517 (N_19517,N_863,N_8654);
nor U19518 (N_19518,N_9858,N_9559);
nand U19519 (N_19519,N_9958,N_5639);
nor U19520 (N_19520,N_1257,N_2239);
xnor U19521 (N_19521,N_2408,N_1102);
nand U19522 (N_19522,N_4774,N_4950);
nor U19523 (N_19523,N_7540,N_1151);
and U19524 (N_19524,N_7065,N_4179);
nand U19525 (N_19525,N_8328,N_4568);
nor U19526 (N_19526,N_6408,N_7686);
nand U19527 (N_19527,N_3329,N_2554);
or U19528 (N_19528,N_4991,N_7147);
or U19529 (N_19529,N_3584,N_5316);
or U19530 (N_19530,N_6829,N_5744);
and U19531 (N_19531,N_1601,N_8840);
or U19532 (N_19532,N_1175,N_675);
xnor U19533 (N_19533,N_4584,N_5320);
nand U19534 (N_19534,N_3563,N_6040);
xor U19535 (N_19535,N_8689,N_9418);
or U19536 (N_19536,N_5527,N_1133);
nand U19537 (N_19537,N_5569,N_5489);
nor U19538 (N_19538,N_32,N_1510);
nor U19539 (N_19539,N_5109,N_4338);
or U19540 (N_19540,N_1567,N_5960);
nor U19541 (N_19541,N_5538,N_9299);
nand U19542 (N_19542,N_295,N_9392);
or U19543 (N_19543,N_7497,N_2312);
nor U19544 (N_19544,N_1013,N_6427);
nand U19545 (N_19545,N_1069,N_506);
nand U19546 (N_19546,N_6272,N_4748);
nand U19547 (N_19547,N_9441,N_7011);
or U19548 (N_19548,N_576,N_9570);
xnor U19549 (N_19549,N_7626,N_9458);
and U19550 (N_19550,N_6942,N_9747);
or U19551 (N_19551,N_3213,N_1411);
nand U19552 (N_19552,N_2089,N_9054);
nor U19553 (N_19553,N_3750,N_4722);
nor U19554 (N_19554,N_1165,N_1051);
nor U19555 (N_19555,N_847,N_4215);
or U19556 (N_19556,N_3200,N_6653);
and U19557 (N_19557,N_6730,N_6907);
or U19558 (N_19558,N_1115,N_2908);
and U19559 (N_19559,N_1363,N_6096);
nand U19560 (N_19560,N_5483,N_8071);
xor U19561 (N_19561,N_1047,N_5957);
or U19562 (N_19562,N_77,N_542);
xor U19563 (N_19563,N_7317,N_1172);
or U19564 (N_19564,N_538,N_3478);
xor U19565 (N_19565,N_9588,N_6285);
or U19566 (N_19566,N_4997,N_8146);
nand U19567 (N_19567,N_8644,N_8617);
nor U19568 (N_19568,N_3617,N_280);
nor U19569 (N_19569,N_2122,N_5561);
xor U19570 (N_19570,N_5205,N_4524);
nor U19571 (N_19571,N_3815,N_4559);
and U19572 (N_19572,N_8570,N_8264);
nand U19573 (N_19573,N_2358,N_9963);
nor U19574 (N_19574,N_4110,N_2834);
and U19575 (N_19575,N_5935,N_3099);
nor U19576 (N_19576,N_2060,N_3097);
nand U19577 (N_19577,N_6885,N_3856);
nor U19578 (N_19578,N_8349,N_6317);
and U19579 (N_19579,N_6608,N_2258);
nor U19580 (N_19580,N_5800,N_42);
xnor U19581 (N_19581,N_5833,N_2243);
and U19582 (N_19582,N_808,N_1935);
nor U19583 (N_19583,N_99,N_7564);
nor U19584 (N_19584,N_6933,N_2623);
nor U19585 (N_19585,N_3721,N_180);
xor U19586 (N_19586,N_5935,N_9082);
nand U19587 (N_19587,N_2266,N_5398);
and U19588 (N_19588,N_5054,N_265);
and U19589 (N_19589,N_4814,N_8172);
nand U19590 (N_19590,N_90,N_2024);
nor U19591 (N_19591,N_9736,N_3995);
nand U19592 (N_19592,N_5774,N_4653);
xnor U19593 (N_19593,N_3393,N_5648);
and U19594 (N_19594,N_4357,N_4926);
or U19595 (N_19595,N_1954,N_2000);
and U19596 (N_19596,N_8005,N_1199);
and U19597 (N_19597,N_1430,N_1442);
nor U19598 (N_19598,N_9712,N_7057);
or U19599 (N_19599,N_2337,N_4155);
and U19600 (N_19600,N_8149,N_6366);
nand U19601 (N_19601,N_3771,N_4094);
and U19602 (N_19602,N_7448,N_1641);
or U19603 (N_19603,N_4508,N_1032);
nor U19604 (N_19604,N_3460,N_9996);
and U19605 (N_19605,N_1940,N_3941);
nand U19606 (N_19606,N_4678,N_202);
and U19607 (N_19607,N_2389,N_7410);
or U19608 (N_19608,N_4368,N_3030);
nor U19609 (N_19609,N_5466,N_6080);
xor U19610 (N_19610,N_3029,N_1440);
and U19611 (N_19611,N_2100,N_8120);
nand U19612 (N_19612,N_5077,N_3348);
or U19613 (N_19613,N_6631,N_5836);
or U19614 (N_19614,N_5639,N_7854);
nand U19615 (N_19615,N_6400,N_5124);
nand U19616 (N_19616,N_2523,N_2855);
and U19617 (N_19617,N_3276,N_1015);
xor U19618 (N_19618,N_2106,N_4355);
xor U19619 (N_19619,N_1385,N_9745);
xnor U19620 (N_19620,N_9434,N_2282);
nand U19621 (N_19621,N_4965,N_431);
nand U19622 (N_19622,N_6563,N_4238);
and U19623 (N_19623,N_2881,N_4969);
nand U19624 (N_19624,N_8982,N_3055);
or U19625 (N_19625,N_3209,N_7213);
xor U19626 (N_19626,N_2163,N_8576);
and U19627 (N_19627,N_7734,N_2067);
or U19628 (N_19628,N_8778,N_8627);
xnor U19629 (N_19629,N_4406,N_3857);
xor U19630 (N_19630,N_9732,N_6496);
or U19631 (N_19631,N_864,N_7963);
or U19632 (N_19632,N_3602,N_614);
and U19633 (N_19633,N_1106,N_1192);
or U19634 (N_19634,N_5730,N_8724);
and U19635 (N_19635,N_2392,N_4361);
nor U19636 (N_19636,N_3741,N_7870);
nand U19637 (N_19637,N_6385,N_1469);
and U19638 (N_19638,N_5979,N_1872);
or U19639 (N_19639,N_5074,N_4784);
or U19640 (N_19640,N_2421,N_1393);
xor U19641 (N_19641,N_5362,N_4821);
nand U19642 (N_19642,N_2380,N_4595);
nand U19643 (N_19643,N_3390,N_8758);
or U19644 (N_19644,N_8135,N_4691);
nand U19645 (N_19645,N_4470,N_7369);
nor U19646 (N_19646,N_4309,N_6666);
nor U19647 (N_19647,N_6881,N_8354);
nor U19648 (N_19648,N_641,N_9076);
and U19649 (N_19649,N_2032,N_20);
or U19650 (N_19650,N_9981,N_6585);
nand U19651 (N_19651,N_5546,N_3234);
or U19652 (N_19652,N_8094,N_4781);
and U19653 (N_19653,N_3982,N_4940);
or U19654 (N_19654,N_5489,N_4451);
xor U19655 (N_19655,N_7638,N_2528);
nor U19656 (N_19656,N_7003,N_6996);
nor U19657 (N_19657,N_5297,N_4749);
nand U19658 (N_19658,N_3816,N_5718);
nand U19659 (N_19659,N_2561,N_9775);
and U19660 (N_19660,N_3759,N_1452);
xor U19661 (N_19661,N_4415,N_2232);
nand U19662 (N_19662,N_225,N_1708);
or U19663 (N_19663,N_5307,N_2993);
or U19664 (N_19664,N_9776,N_8945);
nor U19665 (N_19665,N_5461,N_1923);
and U19666 (N_19666,N_4532,N_2295);
or U19667 (N_19667,N_3286,N_533);
and U19668 (N_19668,N_3220,N_5306);
and U19669 (N_19669,N_9085,N_949);
or U19670 (N_19670,N_7464,N_8813);
nand U19671 (N_19671,N_6206,N_6434);
and U19672 (N_19672,N_6458,N_7585);
nand U19673 (N_19673,N_8433,N_3648);
xnor U19674 (N_19674,N_5848,N_7510);
nand U19675 (N_19675,N_9699,N_5207);
nor U19676 (N_19676,N_7258,N_9781);
or U19677 (N_19677,N_8841,N_1810);
or U19678 (N_19678,N_8405,N_3419);
and U19679 (N_19679,N_7275,N_268);
nand U19680 (N_19680,N_3318,N_8416);
nand U19681 (N_19681,N_4770,N_3886);
nor U19682 (N_19682,N_7459,N_9427);
nor U19683 (N_19683,N_3815,N_8847);
nor U19684 (N_19684,N_2729,N_3923);
nor U19685 (N_19685,N_6735,N_6382);
nor U19686 (N_19686,N_9956,N_3322);
nor U19687 (N_19687,N_4164,N_6527);
nand U19688 (N_19688,N_558,N_2714);
nand U19689 (N_19689,N_5521,N_326);
nand U19690 (N_19690,N_7232,N_7919);
and U19691 (N_19691,N_7612,N_8481);
nor U19692 (N_19692,N_4463,N_5459);
nand U19693 (N_19693,N_1602,N_311);
or U19694 (N_19694,N_3686,N_3189);
nand U19695 (N_19695,N_6247,N_5998);
nand U19696 (N_19696,N_1633,N_9714);
and U19697 (N_19697,N_4205,N_4089);
or U19698 (N_19698,N_8914,N_8526);
or U19699 (N_19699,N_1924,N_4332);
nand U19700 (N_19700,N_8040,N_2076);
nor U19701 (N_19701,N_3812,N_4792);
and U19702 (N_19702,N_6950,N_2204);
and U19703 (N_19703,N_611,N_1501);
and U19704 (N_19704,N_7846,N_6805);
nor U19705 (N_19705,N_4848,N_507);
nand U19706 (N_19706,N_6883,N_3692);
xor U19707 (N_19707,N_2502,N_3430);
nand U19708 (N_19708,N_2594,N_6362);
and U19709 (N_19709,N_1215,N_4075);
nand U19710 (N_19710,N_6847,N_1014);
nand U19711 (N_19711,N_1250,N_1941);
xnor U19712 (N_19712,N_3590,N_8627);
and U19713 (N_19713,N_4207,N_9003);
nor U19714 (N_19714,N_3072,N_1371);
and U19715 (N_19715,N_4312,N_9549);
xor U19716 (N_19716,N_3392,N_8195);
nor U19717 (N_19717,N_4583,N_5850);
nand U19718 (N_19718,N_6817,N_1663);
xor U19719 (N_19719,N_2764,N_4166);
and U19720 (N_19720,N_6358,N_9675);
or U19721 (N_19721,N_2797,N_1826);
and U19722 (N_19722,N_6702,N_4227);
nand U19723 (N_19723,N_6747,N_363);
nand U19724 (N_19724,N_5835,N_6490);
xnor U19725 (N_19725,N_2152,N_1656);
nand U19726 (N_19726,N_6731,N_3952);
nand U19727 (N_19727,N_661,N_4855);
nand U19728 (N_19728,N_1685,N_1911);
and U19729 (N_19729,N_1025,N_4034);
or U19730 (N_19730,N_488,N_4419);
xor U19731 (N_19731,N_8686,N_6240);
and U19732 (N_19732,N_4969,N_7084);
or U19733 (N_19733,N_5152,N_8675);
nor U19734 (N_19734,N_6405,N_7028);
or U19735 (N_19735,N_8193,N_9496);
nor U19736 (N_19736,N_8611,N_5521);
nand U19737 (N_19737,N_1335,N_6737);
and U19738 (N_19738,N_1745,N_6712);
nor U19739 (N_19739,N_6261,N_2582);
nand U19740 (N_19740,N_6710,N_4208);
nor U19741 (N_19741,N_8616,N_7341);
or U19742 (N_19742,N_5771,N_9655);
or U19743 (N_19743,N_899,N_7013);
or U19744 (N_19744,N_6347,N_9351);
and U19745 (N_19745,N_7700,N_2572);
nor U19746 (N_19746,N_518,N_3707);
or U19747 (N_19747,N_9974,N_9832);
and U19748 (N_19748,N_6847,N_3296);
nor U19749 (N_19749,N_5407,N_700);
or U19750 (N_19750,N_8568,N_3772);
or U19751 (N_19751,N_9987,N_858);
nand U19752 (N_19752,N_8296,N_8514);
nor U19753 (N_19753,N_8740,N_8203);
and U19754 (N_19754,N_5175,N_2913);
and U19755 (N_19755,N_9231,N_1239);
or U19756 (N_19756,N_1203,N_7920);
nand U19757 (N_19757,N_5026,N_4391);
nor U19758 (N_19758,N_2727,N_9397);
and U19759 (N_19759,N_5786,N_5400);
nor U19760 (N_19760,N_7731,N_9878);
xor U19761 (N_19761,N_5262,N_501);
nand U19762 (N_19762,N_9887,N_1595);
xor U19763 (N_19763,N_3179,N_902);
nor U19764 (N_19764,N_912,N_2162);
and U19765 (N_19765,N_7313,N_5403);
or U19766 (N_19766,N_1691,N_2337);
or U19767 (N_19767,N_4231,N_8180);
nor U19768 (N_19768,N_2454,N_1142);
and U19769 (N_19769,N_9760,N_9511);
nor U19770 (N_19770,N_8904,N_3334);
or U19771 (N_19771,N_315,N_9331);
and U19772 (N_19772,N_1456,N_3436);
and U19773 (N_19773,N_2969,N_3623);
nand U19774 (N_19774,N_1261,N_5217);
and U19775 (N_19775,N_922,N_2306);
nor U19776 (N_19776,N_3674,N_4219);
nand U19777 (N_19777,N_3785,N_5538);
nor U19778 (N_19778,N_5224,N_7632);
or U19779 (N_19779,N_7869,N_8275);
nand U19780 (N_19780,N_4871,N_3500);
and U19781 (N_19781,N_9283,N_2391);
and U19782 (N_19782,N_1606,N_3607);
or U19783 (N_19783,N_7356,N_888);
xnor U19784 (N_19784,N_5709,N_2382);
nor U19785 (N_19785,N_7831,N_5606);
nor U19786 (N_19786,N_2245,N_4527);
or U19787 (N_19787,N_1005,N_3897);
nor U19788 (N_19788,N_2906,N_6298);
and U19789 (N_19789,N_8466,N_302);
xor U19790 (N_19790,N_5827,N_6313);
nor U19791 (N_19791,N_6843,N_8209);
nand U19792 (N_19792,N_8575,N_2417);
and U19793 (N_19793,N_2327,N_6062);
nand U19794 (N_19794,N_1645,N_5039);
or U19795 (N_19795,N_2249,N_7484);
nor U19796 (N_19796,N_9232,N_5079);
or U19797 (N_19797,N_917,N_1395);
xor U19798 (N_19798,N_9312,N_8754);
nor U19799 (N_19799,N_1240,N_1261);
or U19800 (N_19800,N_3938,N_9981);
nor U19801 (N_19801,N_9394,N_7447);
xor U19802 (N_19802,N_2686,N_3754);
and U19803 (N_19803,N_3909,N_6756);
or U19804 (N_19804,N_3604,N_721);
nor U19805 (N_19805,N_952,N_9430);
and U19806 (N_19806,N_3149,N_1972);
or U19807 (N_19807,N_6716,N_7558);
and U19808 (N_19808,N_781,N_1968);
or U19809 (N_19809,N_1382,N_7462);
or U19810 (N_19810,N_166,N_6652);
or U19811 (N_19811,N_4081,N_99);
and U19812 (N_19812,N_3314,N_460);
nor U19813 (N_19813,N_4595,N_6320);
xnor U19814 (N_19814,N_7458,N_6413);
or U19815 (N_19815,N_986,N_9588);
xnor U19816 (N_19816,N_7656,N_2044);
or U19817 (N_19817,N_9149,N_7076);
nand U19818 (N_19818,N_8018,N_9807);
nand U19819 (N_19819,N_3347,N_7167);
and U19820 (N_19820,N_315,N_896);
nor U19821 (N_19821,N_7626,N_911);
and U19822 (N_19822,N_6337,N_9192);
and U19823 (N_19823,N_2744,N_9487);
or U19824 (N_19824,N_7772,N_7086);
and U19825 (N_19825,N_253,N_5323);
nor U19826 (N_19826,N_6653,N_4302);
and U19827 (N_19827,N_557,N_7837);
or U19828 (N_19828,N_4635,N_4204);
nor U19829 (N_19829,N_9298,N_4419);
nor U19830 (N_19830,N_7959,N_9039);
or U19831 (N_19831,N_5331,N_350);
or U19832 (N_19832,N_1633,N_732);
nand U19833 (N_19833,N_4302,N_300);
and U19834 (N_19834,N_2919,N_4733);
and U19835 (N_19835,N_9617,N_2314);
nor U19836 (N_19836,N_1003,N_1096);
and U19837 (N_19837,N_7894,N_4806);
or U19838 (N_19838,N_9325,N_8600);
or U19839 (N_19839,N_8381,N_9573);
or U19840 (N_19840,N_214,N_8795);
or U19841 (N_19841,N_4693,N_5432);
nand U19842 (N_19842,N_4720,N_5225);
nor U19843 (N_19843,N_5732,N_5587);
nor U19844 (N_19844,N_1165,N_9771);
nor U19845 (N_19845,N_4142,N_2498);
and U19846 (N_19846,N_8149,N_9896);
and U19847 (N_19847,N_5141,N_9185);
nor U19848 (N_19848,N_404,N_7622);
nand U19849 (N_19849,N_2187,N_9468);
or U19850 (N_19850,N_9263,N_9370);
and U19851 (N_19851,N_8493,N_7184);
and U19852 (N_19852,N_4730,N_6983);
and U19853 (N_19853,N_4872,N_5498);
or U19854 (N_19854,N_9402,N_7324);
nor U19855 (N_19855,N_4518,N_231);
nor U19856 (N_19856,N_8822,N_2165);
nand U19857 (N_19857,N_3301,N_6582);
nor U19858 (N_19858,N_703,N_7562);
or U19859 (N_19859,N_2470,N_5485);
or U19860 (N_19860,N_8238,N_6190);
or U19861 (N_19861,N_1091,N_4275);
nor U19862 (N_19862,N_4574,N_4289);
and U19863 (N_19863,N_7213,N_8852);
or U19864 (N_19864,N_1963,N_8999);
xor U19865 (N_19865,N_3000,N_7982);
nand U19866 (N_19866,N_9591,N_5820);
or U19867 (N_19867,N_8202,N_7408);
or U19868 (N_19868,N_2088,N_4433);
nor U19869 (N_19869,N_7025,N_1523);
nand U19870 (N_19870,N_8467,N_1390);
nand U19871 (N_19871,N_624,N_5981);
and U19872 (N_19872,N_637,N_1930);
or U19873 (N_19873,N_1611,N_1305);
or U19874 (N_19874,N_4762,N_1873);
nor U19875 (N_19875,N_2435,N_9987);
and U19876 (N_19876,N_2957,N_1784);
and U19877 (N_19877,N_1205,N_3110);
and U19878 (N_19878,N_8438,N_3454);
and U19879 (N_19879,N_3273,N_2248);
nor U19880 (N_19880,N_1135,N_878);
nor U19881 (N_19881,N_3369,N_26);
nand U19882 (N_19882,N_7932,N_7703);
or U19883 (N_19883,N_5603,N_6408);
xnor U19884 (N_19884,N_8871,N_7688);
nor U19885 (N_19885,N_6731,N_2287);
and U19886 (N_19886,N_5716,N_4176);
or U19887 (N_19887,N_6449,N_2344);
xor U19888 (N_19888,N_2147,N_7210);
and U19889 (N_19889,N_1785,N_977);
nand U19890 (N_19890,N_3912,N_3149);
xnor U19891 (N_19891,N_8479,N_8361);
nand U19892 (N_19892,N_4208,N_7981);
nor U19893 (N_19893,N_2327,N_7190);
or U19894 (N_19894,N_765,N_7946);
and U19895 (N_19895,N_6534,N_9163);
nand U19896 (N_19896,N_8612,N_536);
and U19897 (N_19897,N_3599,N_6102);
or U19898 (N_19898,N_9370,N_4471);
nor U19899 (N_19899,N_6976,N_2298);
nand U19900 (N_19900,N_9823,N_9826);
and U19901 (N_19901,N_1795,N_9593);
xor U19902 (N_19902,N_3499,N_9596);
or U19903 (N_19903,N_5975,N_796);
and U19904 (N_19904,N_1187,N_2664);
xor U19905 (N_19905,N_767,N_5580);
nand U19906 (N_19906,N_4386,N_9327);
nand U19907 (N_19907,N_6560,N_5656);
or U19908 (N_19908,N_3209,N_3187);
nand U19909 (N_19909,N_6573,N_2330);
and U19910 (N_19910,N_4214,N_546);
nor U19911 (N_19911,N_6595,N_261);
nand U19912 (N_19912,N_530,N_2807);
or U19913 (N_19913,N_7172,N_9832);
or U19914 (N_19914,N_3184,N_7424);
nand U19915 (N_19915,N_1139,N_2765);
or U19916 (N_19916,N_45,N_8583);
nand U19917 (N_19917,N_2326,N_7731);
and U19918 (N_19918,N_3061,N_840);
and U19919 (N_19919,N_9680,N_2100);
nor U19920 (N_19920,N_612,N_9262);
and U19921 (N_19921,N_4631,N_7632);
nor U19922 (N_19922,N_6551,N_4465);
nand U19923 (N_19923,N_1879,N_9724);
nor U19924 (N_19924,N_8487,N_1679);
nand U19925 (N_19925,N_8000,N_1579);
nor U19926 (N_19926,N_3511,N_5591);
nand U19927 (N_19927,N_6240,N_6452);
and U19928 (N_19928,N_4576,N_9851);
and U19929 (N_19929,N_982,N_9719);
and U19930 (N_19930,N_579,N_9216);
nand U19931 (N_19931,N_8377,N_443);
and U19932 (N_19932,N_5128,N_3012);
xor U19933 (N_19933,N_8457,N_1326);
and U19934 (N_19934,N_6460,N_1720);
nand U19935 (N_19935,N_9814,N_632);
or U19936 (N_19936,N_8093,N_9435);
nor U19937 (N_19937,N_8876,N_1791);
or U19938 (N_19938,N_4891,N_4102);
and U19939 (N_19939,N_7111,N_3177);
nor U19940 (N_19940,N_9122,N_2081);
xor U19941 (N_19941,N_1073,N_7528);
and U19942 (N_19942,N_3864,N_949);
nor U19943 (N_19943,N_7545,N_7363);
nor U19944 (N_19944,N_8349,N_2303);
and U19945 (N_19945,N_2831,N_164);
nor U19946 (N_19946,N_5517,N_1533);
nor U19947 (N_19947,N_7690,N_6993);
nor U19948 (N_19948,N_8595,N_8965);
and U19949 (N_19949,N_6983,N_4417);
nor U19950 (N_19950,N_296,N_8661);
nor U19951 (N_19951,N_9343,N_9501);
nor U19952 (N_19952,N_2221,N_639);
nand U19953 (N_19953,N_1003,N_6174);
nor U19954 (N_19954,N_2360,N_9489);
or U19955 (N_19955,N_3303,N_4482);
nand U19956 (N_19956,N_5577,N_625);
and U19957 (N_19957,N_7836,N_7673);
or U19958 (N_19958,N_5414,N_220);
xnor U19959 (N_19959,N_574,N_1095);
and U19960 (N_19960,N_7566,N_8518);
nor U19961 (N_19961,N_9466,N_5105);
xor U19962 (N_19962,N_1291,N_7320);
and U19963 (N_19963,N_5895,N_1652);
or U19964 (N_19964,N_1786,N_5655);
nor U19965 (N_19965,N_2665,N_3970);
and U19966 (N_19966,N_4952,N_1471);
or U19967 (N_19967,N_6651,N_5960);
and U19968 (N_19968,N_9227,N_7958);
and U19969 (N_19969,N_2675,N_1692);
or U19970 (N_19970,N_4807,N_4630);
nand U19971 (N_19971,N_3897,N_1139);
or U19972 (N_19972,N_9701,N_6526);
or U19973 (N_19973,N_6081,N_7235);
and U19974 (N_19974,N_8493,N_2305);
nand U19975 (N_19975,N_4473,N_1905);
and U19976 (N_19976,N_6114,N_1636);
or U19977 (N_19977,N_6490,N_4878);
or U19978 (N_19978,N_401,N_3689);
nor U19979 (N_19979,N_3494,N_6384);
nor U19980 (N_19980,N_4612,N_1874);
nand U19981 (N_19981,N_4976,N_6083);
nand U19982 (N_19982,N_9245,N_2936);
or U19983 (N_19983,N_2832,N_1975);
nor U19984 (N_19984,N_6390,N_5234);
and U19985 (N_19985,N_8960,N_1337);
nand U19986 (N_19986,N_4319,N_2214);
and U19987 (N_19987,N_4984,N_3126);
or U19988 (N_19988,N_8047,N_2182);
or U19989 (N_19989,N_8579,N_7153);
nand U19990 (N_19990,N_1587,N_3938);
nand U19991 (N_19991,N_9959,N_9737);
nand U19992 (N_19992,N_2380,N_504);
nand U19993 (N_19993,N_9739,N_461);
nand U19994 (N_19994,N_4340,N_2422);
nand U19995 (N_19995,N_8624,N_3802);
nand U19996 (N_19996,N_1849,N_3071);
and U19997 (N_19997,N_4944,N_2436);
nor U19998 (N_19998,N_3093,N_1287);
nand U19999 (N_19999,N_5614,N_3391);
nand U20000 (N_20000,N_18248,N_18640);
or U20001 (N_20001,N_11740,N_12886);
or U20002 (N_20002,N_16920,N_15140);
and U20003 (N_20003,N_17342,N_10950);
nor U20004 (N_20004,N_16302,N_16877);
nor U20005 (N_20005,N_14256,N_18861);
nand U20006 (N_20006,N_16164,N_16671);
nand U20007 (N_20007,N_18084,N_10702);
xnor U20008 (N_20008,N_14724,N_16637);
xnor U20009 (N_20009,N_13670,N_17271);
or U20010 (N_20010,N_18060,N_15805);
nand U20011 (N_20011,N_17936,N_18443);
or U20012 (N_20012,N_17671,N_11530);
and U20013 (N_20013,N_13816,N_13290);
or U20014 (N_20014,N_12214,N_12089);
or U20015 (N_20015,N_12487,N_15504);
and U20016 (N_20016,N_19635,N_17590);
xor U20017 (N_20017,N_14632,N_13633);
nand U20018 (N_20018,N_11482,N_16474);
or U20019 (N_20019,N_17270,N_17012);
and U20020 (N_20020,N_13729,N_18730);
nor U20021 (N_20021,N_11967,N_17319);
and U20022 (N_20022,N_11010,N_10169);
and U20023 (N_20023,N_11420,N_18438);
xnor U20024 (N_20024,N_11802,N_10616);
and U20025 (N_20025,N_18340,N_16396);
nand U20026 (N_20026,N_17388,N_19953);
nand U20027 (N_20027,N_10333,N_16694);
or U20028 (N_20028,N_18641,N_12553);
or U20029 (N_20029,N_16228,N_14783);
or U20030 (N_20030,N_11697,N_16995);
or U20031 (N_20031,N_13712,N_16518);
xnor U20032 (N_20032,N_11952,N_15439);
nor U20033 (N_20033,N_14085,N_13409);
nand U20034 (N_20034,N_11619,N_18965);
nand U20035 (N_20035,N_13149,N_18552);
or U20036 (N_20036,N_15577,N_10152);
and U20037 (N_20037,N_14268,N_11483);
or U20038 (N_20038,N_18910,N_11507);
and U20039 (N_20039,N_10649,N_19462);
nor U20040 (N_20040,N_13175,N_16197);
xnor U20041 (N_20041,N_11661,N_11291);
nor U20042 (N_20042,N_10407,N_16574);
nor U20043 (N_20043,N_14584,N_10971);
or U20044 (N_20044,N_14689,N_10339);
nand U20045 (N_20045,N_19310,N_18367);
and U20046 (N_20046,N_12787,N_12692);
nor U20047 (N_20047,N_18960,N_13225);
or U20048 (N_20048,N_14966,N_18122);
nor U20049 (N_20049,N_17364,N_10260);
or U20050 (N_20050,N_17332,N_12765);
nor U20051 (N_20051,N_17172,N_12119);
and U20052 (N_20052,N_13580,N_19941);
and U20053 (N_20053,N_13692,N_10193);
xor U20054 (N_20054,N_14940,N_15114);
nand U20055 (N_20055,N_19902,N_18170);
nor U20056 (N_20056,N_16374,N_14761);
xnor U20057 (N_20057,N_12714,N_19457);
nor U20058 (N_20058,N_12223,N_15860);
or U20059 (N_20059,N_15564,N_13595);
or U20060 (N_20060,N_15502,N_14368);
nand U20061 (N_20061,N_16315,N_19086);
and U20062 (N_20062,N_13344,N_12754);
or U20063 (N_20063,N_13251,N_14103);
nor U20064 (N_20064,N_18288,N_16918);
or U20065 (N_20065,N_11873,N_12306);
nand U20066 (N_20066,N_18653,N_13393);
nor U20067 (N_20067,N_18554,N_16800);
nor U20068 (N_20068,N_10944,N_11641);
or U20069 (N_20069,N_11701,N_14246);
or U20070 (N_20070,N_17031,N_11643);
nand U20071 (N_20071,N_12622,N_12684);
nand U20072 (N_20072,N_19245,N_15138);
nand U20073 (N_20073,N_11819,N_13226);
and U20074 (N_20074,N_14800,N_14281);
or U20075 (N_20075,N_14189,N_14307);
and U20076 (N_20076,N_17761,N_15496);
nand U20077 (N_20077,N_19639,N_16073);
nand U20078 (N_20078,N_14359,N_17223);
nor U20079 (N_20079,N_12870,N_18390);
and U20080 (N_20080,N_11073,N_10610);
nor U20081 (N_20081,N_11469,N_19063);
or U20082 (N_20082,N_14471,N_19216);
or U20083 (N_20083,N_17589,N_16466);
or U20084 (N_20084,N_14944,N_13492);
nand U20085 (N_20085,N_13497,N_17431);
nand U20086 (N_20086,N_13521,N_11850);
or U20087 (N_20087,N_18987,N_14916);
nor U20088 (N_20088,N_16099,N_18949);
nand U20089 (N_20089,N_17913,N_15836);
xnor U20090 (N_20090,N_12663,N_19071);
nor U20091 (N_20091,N_13807,N_15802);
xnor U20092 (N_20092,N_16236,N_17969);
or U20093 (N_20093,N_13914,N_16125);
and U20094 (N_20094,N_16705,N_11976);
nor U20095 (N_20095,N_15563,N_14133);
nor U20096 (N_20096,N_12300,N_14329);
and U20097 (N_20097,N_11058,N_11508);
nand U20098 (N_20098,N_19599,N_15680);
or U20099 (N_20099,N_18755,N_10886);
and U20100 (N_20100,N_12128,N_13183);
and U20101 (N_20101,N_12875,N_16757);
nor U20102 (N_20102,N_19495,N_18792);
nor U20103 (N_20103,N_12361,N_17766);
and U20104 (N_20104,N_19302,N_11197);
or U20105 (N_20105,N_12731,N_19858);
nand U20106 (N_20106,N_17281,N_17410);
or U20107 (N_20107,N_13618,N_12073);
or U20108 (N_20108,N_12149,N_17113);
or U20109 (N_20109,N_13493,N_11353);
nor U20110 (N_20110,N_15253,N_11553);
nor U20111 (N_20111,N_12415,N_15832);
and U20112 (N_20112,N_14493,N_15491);
and U20113 (N_20113,N_10862,N_10483);
or U20114 (N_20114,N_11229,N_12613);
xor U20115 (N_20115,N_17494,N_10527);
nand U20116 (N_20116,N_16308,N_18754);
nor U20117 (N_20117,N_10929,N_17227);
nor U20118 (N_20118,N_11209,N_14848);
or U20119 (N_20119,N_17507,N_17219);
or U20120 (N_20120,N_15735,N_16301);
xnor U20121 (N_20121,N_15488,N_19783);
nor U20122 (N_20122,N_11360,N_19368);
or U20123 (N_20123,N_13390,N_16990);
and U20124 (N_20124,N_15905,N_18068);
or U20125 (N_20125,N_13323,N_11236);
xnor U20126 (N_20126,N_15745,N_17579);
nand U20127 (N_20127,N_18293,N_10437);
or U20128 (N_20128,N_18079,N_18400);
nor U20129 (N_20129,N_13498,N_19905);
and U20130 (N_20130,N_17194,N_16536);
and U20131 (N_20131,N_15196,N_13810);
or U20132 (N_20132,N_17192,N_12810);
and U20133 (N_20133,N_19002,N_11940);
nor U20134 (N_20134,N_17749,N_10191);
or U20135 (N_20135,N_10392,N_13177);
and U20136 (N_20136,N_15125,N_15009);
or U20137 (N_20137,N_16468,N_18875);
and U20138 (N_20138,N_13252,N_19722);
or U20139 (N_20139,N_18059,N_11866);
nand U20140 (N_20140,N_17620,N_14156);
nor U20141 (N_20141,N_15049,N_11301);
or U20142 (N_20142,N_17122,N_14529);
or U20143 (N_20143,N_15139,N_12228);
or U20144 (N_20144,N_10073,N_18114);
nor U20145 (N_20145,N_12541,N_11936);
nand U20146 (N_20146,N_17720,N_13241);
nand U20147 (N_20147,N_16475,N_18954);
or U20148 (N_20148,N_13714,N_17242);
or U20149 (N_20149,N_13327,N_10672);
nor U20150 (N_20150,N_15963,N_10298);
nor U20151 (N_20151,N_15409,N_18610);
and U20152 (N_20152,N_18865,N_10291);
or U20153 (N_20153,N_15547,N_19480);
xor U20154 (N_20154,N_12166,N_13439);
nor U20155 (N_20155,N_16741,N_17696);
nor U20156 (N_20156,N_16887,N_12769);
nor U20157 (N_20157,N_14324,N_17167);
and U20158 (N_20158,N_16435,N_13775);
nor U20159 (N_20159,N_16392,N_18631);
and U20160 (N_20160,N_19373,N_18428);
nor U20161 (N_20161,N_16847,N_16379);
or U20162 (N_20162,N_19637,N_13533);
nor U20163 (N_20163,N_11259,N_10074);
or U20164 (N_20164,N_15320,N_16003);
nand U20165 (N_20165,N_18729,N_13785);
and U20166 (N_20166,N_12456,N_10151);
nand U20167 (N_20167,N_17970,N_10962);
nor U20168 (N_20168,N_17309,N_15069);
nor U20169 (N_20169,N_10079,N_12463);
or U20170 (N_20170,N_14150,N_14045);
or U20171 (N_20171,N_11849,N_16166);
nor U20172 (N_20172,N_14962,N_14975);
nand U20173 (N_20173,N_15782,N_15800);
nor U20174 (N_20174,N_14861,N_12389);
xnor U20175 (N_20175,N_14625,N_11309);
and U20176 (N_20176,N_10268,N_12177);
nor U20177 (N_20177,N_18587,N_13683);
nand U20178 (N_20178,N_15904,N_14597);
and U20179 (N_20179,N_19167,N_16141);
xnor U20180 (N_20180,N_17591,N_10102);
nor U20181 (N_20181,N_11723,N_11835);
nor U20182 (N_20182,N_11329,N_13347);
nor U20183 (N_20183,N_19991,N_16018);
nand U20184 (N_20184,N_14267,N_12885);
or U20185 (N_20185,N_18284,N_17041);
or U20186 (N_20186,N_15042,N_17793);
and U20187 (N_20187,N_16034,N_17274);
nor U20188 (N_20188,N_18734,N_11698);
and U20189 (N_20189,N_11522,N_19734);
nand U20190 (N_20190,N_19698,N_16794);
nor U20191 (N_20191,N_11974,N_11574);
or U20192 (N_20192,N_18147,N_13564);
xor U20193 (N_20193,N_11511,N_12724);
nor U20194 (N_20194,N_15672,N_13250);
or U20195 (N_20195,N_14193,N_18991);
and U20196 (N_20196,N_17797,N_13228);
and U20197 (N_20197,N_14185,N_19388);
nor U20198 (N_20198,N_18869,N_19037);
or U20199 (N_20199,N_17030,N_14575);
nor U20200 (N_20200,N_19260,N_15464);
and U20201 (N_20201,N_19828,N_10590);
or U20202 (N_20202,N_13106,N_14637);
nor U20203 (N_20203,N_15168,N_18789);
and U20204 (N_20204,N_18990,N_12318);
xnor U20205 (N_20205,N_15667,N_16978);
and U20206 (N_20206,N_19837,N_13287);
xnor U20207 (N_20207,N_10372,N_11141);
nor U20208 (N_20208,N_13898,N_13457);
or U20209 (N_20209,N_13018,N_10632);
and U20210 (N_20210,N_15354,N_17770);
or U20211 (N_20211,N_19419,N_14518);
or U20212 (N_20212,N_19735,N_13757);
nor U20213 (N_20213,N_16597,N_11671);
or U20214 (N_20214,N_15821,N_14726);
nand U20215 (N_20215,N_11855,N_11818);
or U20216 (N_20216,N_14473,N_15005);
nand U20217 (N_20217,N_11251,N_18778);
xnor U20218 (N_20218,N_13306,N_18576);
or U20219 (N_20219,N_10229,N_18224);
or U20220 (N_20220,N_10824,N_19272);
or U20221 (N_20221,N_13219,N_17385);
nand U20222 (N_20222,N_11039,N_18444);
or U20223 (N_20223,N_10168,N_16243);
and U20224 (N_20224,N_10438,N_15734);
nor U20225 (N_20225,N_19608,N_11061);
and U20226 (N_20226,N_17175,N_11402);
and U20227 (N_20227,N_18983,N_15273);
and U20228 (N_20228,N_10237,N_16838);
and U20229 (N_20229,N_14224,N_15131);
and U20230 (N_20230,N_19056,N_13236);
or U20231 (N_20231,N_16378,N_18590);
nand U20232 (N_20232,N_15119,N_15789);
nor U20233 (N_20233,N_18155,N_12010);
and U20234 (N_20234,N_13234,N_19728);
or U20235 (N_20235,N_13075,N_18593);
xor U20236 (N_20236,N_12403,N_12657);
xor U20237 (N_20237,N_14757,N_14439);
nand U20238 (N_20238,N_13561,N_16304);
nor U20239 (N_20239,N_16805,N_10978);
or U20240 (N_20240,N_15780,N_17341);
nand U20241 (N_20241,N_18484,N_19155);
or U20242 (N_20242,N_16085,N_17047);
nand U20243 (N_20243,N_17107,N_11627);
and U20244 (N_20244,N_11930,N_11665);
and U20245 (N_20245,N_16987,N_16780);
xor U20246 (N_20246,N_17977,N_17790);
nand U20247 (N_20247,N_19811,N_17644);
or U20248 (N_20248,N_13639,N_16495);
nand U20249 (N_20249,N_15787,N_19697);
nand U20250 (N_20250,N_14852,N_17256);
nor U20251 (N_20251,N_14688,N_11862);
xor U20252 (N_20252,N_17756,N_12619);
or U20253 (N_20253,N_10968,N_15791);
nor U20254 (N_20254,N_17209,N_13191);
nor U20255 (N_20255,N_10119,N_15418);
and U20256 (N_20256,N_14499,N_10382);
or U20257 (N_20257,N_10373,N_11231);
and U20258 (N_20258,N_18320,N_12240);
nand U20259 (N_20259,N_15869,N_13966);
and U20260 (N_20260,N_18324,N_19823);
nand U20261 (N_20261,N_13356,N_10424);
nand U20262 (N_20262,N_12921,N_18900);
xnor U20263 (N_20263,N_15096,N_14040);
nand U20264 (N_20264,N_11812,N_12156);
nand U20265 (N_20265,N_11751,N_11765);
and U20266 (N_20266,N_15285,N_13360);
xnor U20267 (N_20267,N_11100,N_13253);
or U20268 (N_20268,N_15443,N_19113);
nor U20269 (N_20269,N_10953,N_14260);
nor U20270 (N_20270,N_11026,N_12586);
and U20271 (N_20271,N_19426,N_16989);
or U20272 (N_20272,N_14673,N_11768);
nor U20273 (N_20273,N_17779,N_13845);
and U20274 (N_20274,N_17964,N_11924);
xor U20275 (N_20275,N_18223,N_19282);
and U20276 (N_20276,N_12347,N_19038);
or U20277 (N_20277,N_15662,N_15848);
xor U20278 (N_20278,N_18595,N_10288);
or U20279 (N_20279,N_18636,N_15030);
xor U20280 (N_20280,N_14259,N_17940);
or U20281 (N_20281,N_16101,N_11846);
or U20282 (N_20282,N_16562,N_14098);
and U20283 (N_20283,N_18879,N_19505);
or U20284 (N_20284,N_12579,N_17066);
or U20285 (N_20285,N_12862,N_10835);
or U20286 (N_20286,N_12175,N_15959);
and U20287 (N_20287,N_16948,N_10469);
nor U20288 (N_20288,N_18659,N_18495);
nor U20289 (N_20289,N_12367,N_18748);
nor U20290 (N_20290,N_15639,N_11869);
and U20291 (N_20291,N_17515,N_12880);
nand U20292 (N_20292,N_12062,N_18855);
nand U20293 (N_20293,N_15580,N_16114);
or U20294 (N_20294,N_12797,N_17445);
nor U20295 (N_20295,N_11839,N_12064);
nand U20296 (N_20296,N_12445,N_14312);
xor U20297 (N_20297,N_15484,N_15307);
and U20298 (N_20298,N_17234,N_15663);
nand U20299 (N_20299,N_10426,N_12668);
nand U20300 (N_20300,N_10751,N_15445);
and U20301 (N_20301,N_14500,N_16909);
nand U20302 (N_20302,N_13419,N_10493);
xor U20303 (N_20303,N_15703,N_12493);
and U20304 (N_20304,N_15562,N_15083);
xor U20305 (N_20305,N_15644,N_18821);
nor U20306 (N_20306,N_15766,N_18185);
nand U20307 (N_20307,N_15152,N_13593);
nor U20308 (N_20308,N_12491,N_16727);
or U20309 (N_20309,N_17626,N_13658);
and U20310 (N_20310,N_19927,N_17017);
and U20311 (N_20311,N_11993,N_16258);
or U20312 (N_20312,N_19416,N_17942);
xnor U20313 (N_20313,N_17144,N_18193);
and U20314 (N_20314,N_15775,N_11386);
and U20315 (N_20315,N_14340,N_12337);
nor U20316 (N_20316,N_19672,N_14441);
and U20317 (N_20317,N_12653,N_12798);
or U20318 (N_20318,N_12977,N_10986);
nand U20319 (N_20319,N_19725,N_16430);
xor U20320 (N_20320,N_19704,N_18795);
or U20321 (N_20321,N_18623,N_10252);
xnor U20322 (N_20322,N_19447,N_13477);
and U20323 (N_20323,N_17432,N_13044);
and U20324 (N_20324,N_15723,N_18429);
nor U20325 (N_20325,N_15180,N_16211);
nor U20326 (N_20326,N_18322,N_12947);
or U20327 (N_20327,N_11461,N_19138);
xor U20328 (N_20328,N_10982,N_12395);
or U20329 (N_20329,N_12178,N_13152);
and U20330 (N_20330,N_17948,N_18230);
nor U20331 (N_20331,N_17472,N_16496);
and U20332 (N_20332,N_15726,N_11599);
or U20333 (N_20333,N_15010,N_10351);
nor U20334 (N_20334,N_16016,N_18117);
or U20335 (N_20335,N_12323,N_10271);
nand U20336 (N_20336,N_17759,N_19846);
and U20337 (N_20337,N_16604,N_19985);
and U20338 (N_20338,N_17391,N_17393);
xor U20339 (N_20339,N_15317,N_14347);
nand U20340 (N_20340,N_15919,N_17551);
xor U20341 (N_20341,N_16583,N_11826);
nand U20342 (N_20342,N_17982,N_18758);
xor U20343 (N_20343,N_12509,N_14044);
nand U20344 (N_20344,N_10366,N_10566);
and U20345 (N_20345,N_13850,N_18621);
or U20346 (N_20346,N_13599,N_10661);
and U20347 (N_20347,N_11535,N_15906);
or U20348 (N_20348,N_10870,N_10421);
and U20349 (N_20349,N_18442,N_14389);
or U20350 (N_20350,N_15157,N_17555);
xnor U20351 (N_20351,N_18401,N_11738);
xnor U20352 (N_20352,N_15795,N_12015);
and U20353 (N_20353,N_17794,N_13259);
nand U20354 (N_20354,N_11234,N_17814);
nand U20355 (N_20355,N_15252,N_16412);
nor U20356 (N_20356,N_10265,N_10432);
nand U20357 (N_20357,N_12567,N_16157);
nand U20358 (N_20358,N_19893,N_13624);
nor U20359 (N_20359,N_18108,N_11016);
or U20360 (N_20360,N_17003,N_12258);
or U20361 (N_20361,N_18677,N_12560);
or U20362 (N_20362,N_19098,N_14484);
nor U20363 (N_20363,N_15438,N_17803);
or U20364 (N_20364,N_12049,N_16541);
nand U20365 (N_20365,N_17263,N_15308);
or U20366 (N_20366,N_13743,N_17745);
or U20367 (N_20367,N_19726,N_17034);
nand U20368 (N_20368,N_19350,N_13166);
and U20369 (N_20369,N_18012,N_13040);
or U20370 (N_20370,N_12908,N_17447);
and U20371 (N_20371,N_10524,N_17450);
nor U20372 (N_20372,N_10510,N_15687);
nand U20373 (N_20373,N_14911,N_12628);
and U20374 (N_20374,N_16487,N_11052);
nand U20375 (N_20375,N_10980,N_17389);
or U20376 (N_20376,N_16365,N_17430);
nor U20377 (N_20377,N_19771,N_13938);
or U20378 (N_20378,N_14328,N_15094);
nor U20379 (N_20379,N_14686,N_11921);
or U20380 (N_20380,N_14405,N_19409);
xor U20381 (N_20381,N_19361,N_16963);
nand U20382 (N_20382,N_11700,N_14165);
nand U20383 (N_20383,N_12410,N_12350);
xor U20384 (N_20384,N_15322,N_19981);
nand U20385 (N_20385,N_17593,N_11875);
xnor U20386 (N_20386,N_11926,N_10940);
nand U20387 (N_20387,N_19948,N_19178);
xnor U20388 (N_20388,N_19879,N_11813);
and U20389 (N_20389,N_16815,N_18159);
and U20390 (N_20390,N_18948,N_17486);
and U20391 (N_20391,N_16590,N_11983);
nand U20392 (N_20392,N_10383,N_13589);
or U20393 (N_20393,N_13935,N_16086);
or U20394 (N_20394,N_10367,N_19317);
and U20395 (N_20395,N_14535,N_17191);
nor U20396 (N_20396,N_17306,N_13482);
or U20397 (N_20397,N_13636,N_19355);
nand U20398 (N_20398,N_19449,N_17369);
or U20399 (N_20399,N_15421,N_14947);
xor U20400 (N_20400,N_16158,N_11218);
xnor U20401 (N_20401,N_17024,N_13846);
and U20402 (N_20402,N_15804,N_11097);
or U20403 (N_20403,N_14901,N_13544);
nand U20404 (N_20404,N_17606,N_17748);
and U20405 (N_20405,N_16443,N_14558);
nand U20406 (N_20406,N_14554,N_10001);
nand U20407 (N_20407,N_19857,N_15211);
nand U20408 (N_20408,N_14228,N_19912);
or U20409 (N_20409,N_18163,N_10642);
and U20410 (N_20410,N_19108,N_12369);
or U20411 (N_20411,N_11636,N_18505);
or U20412 (N_20412,N_19966,N_17864);
or U20413 (N_20413,N_11409,N_17880);
nand U20414 (N_20414,N_16651,N_11210);
xor U20415 (N_20415,N_19533,N_16032);
nand U20416 (N_20416,N_13456,N_11648);
nand U20417 (N_20417,N_12784,N_11650);
xnor U20418 (N_20418,N_18373,N_12506);
and U20419 (N_20419,N_11472,N_19024);
and U20420 (N_20420,N_11799,N_14690);
xnor U20421 (N_20421,N_13427,N_13706);
nor U20422 (N_20422,N_17233,N_15377);
nand U20423 (N_20423,N_15936,N_15428);
and U20424 (N_20424,N_19179,N_18784);
nor U20425 (N_20425,N_11961,N_15319);
nand U20426 (N_20426,N_15235,N_17534);
and U20427 (N_20427,N_12416,N_10647);
nor U20428 (N_20428,N_16662,N_17096);
and U20429 (N_20429,N_10473,N_17147);
or U20430 (N_20430,N_11895,N_14397);
and U20431 (N_20431,N_11326,N_18984);
nand U20432 (N_20432,N_19943,N_16448);
and U20433 (N_20433,N_10547,N_13527);
nor U20434 (N_20434,N_18346,N_16103);
and U20435 (N_20435,N_18329,N_18289);
or U20436 (N_20436,N_19538,N_14177);
nor U20437 (N_20437,N_18029,N_10007);
or U20438 (N_20438,N_15255,N_12927);
and U20439 (N_20439,N_14196,N_18162);
nand U20440 (N_20440,N_13540,N_17188);
or U20441 (N_20441,N_18024,N_16936);
or U20442 (N_20442,N_14360,N_12325);
nor U20443 (N_20443,N_11677,N_17289);
or U20444 (N_20444,N_19052,N_19122);
or U20445 (N_20445,N_17726,N_15524);
or U20446 (N_20446,N_16769,N_16875);
nand U20447 (N_20447,N_14434,N_17953);
and U20448 (N_20448,N_15654,N_12785);
or U20449 (N_20449,N_13543,N_12530);
nor U20450 (N_20450,N_19968,N_19314);
nand U20451 (N_20451,N_12336,N_15259);
or U20452 (N_20452,N_19978,N_17298);
or U20453 (N_20453,N_15286,N_14404);
nor U20454 (N_20454,N_17828,N_17776);
and U20455 (N_20455,N_10687,N_16001);
xnor U20456 (N_20456,N_12171,N_19579);
nand U20457 (N_20457,N_15493,N_18536);
xor U20458 (N_20458,N_13483,N_19170);
xor U20459 (N_20459,N_10925,N_16093);
or U20460 (N_20460,N_10630,N_17042);
nor U20461 (N_20461,N_18057,N_10577);
or U20462 (N_20462,N_12618,N_19861);
nor U20463 (N_20463,N_19048,N_12414);
nand U20464 (N_20464,N_11998,N_11364);
and U20465 (N_20465,N_12006,N_16009);
and U20466 (N_20466,N_17873,N_15121);
nor U20467 (N_20467,N_12025,N_13433);
and U20468 (N_20468,N_14334,N_14282);
nand U20469 (N_20469,N_10928,N_12262);
or U20470 (N_20470,N_18871,N_16578);
nor U20471 (N_20471,N_13053,N_11805);
nor U20472 (N_20472,N_14609,N_10124);
and U20473 (N_20473,N_16097,N_14876);
xor U20474 (N_20474,N_10126,N_17867);
nand U20475 (N_20475,N_18175,N_15934);
or U20476 (N_20476,N_12867,N_11515);
and U20477 (N_20477,N_19564,N_18834);
nand U20478 (N_20478,N_11506,N_11022);
and U20479 (N_20479,N_18249,N_17625);
nand U20480 (N_20480,N_10419,N_15036);
nor U20481 (N_20481,N_16762,N_19625);
xnor U20482 (N_20482,N_17339,N_17724);
or U20483 (N_20483,N_11897,N_12747);
or U20484 (N_20484,N_15424,N_11132);
and U20485 (N_20485,N_16038,N_17655);
nor U20486 (N_20486,N_12946,N_11966);
nand U20487 (N_20487,N_16550,N_19194);
nand U20488 (N_20488,N_10606,N_12855);
and U20489 (N_20489,N_10192,N_18014);
or U20490 (N_20490,N_11017,N_16270);
nor U20491 (N_20491,N_16993,N_19573);
or U20492 (N_20492,N_12597,N_13311);
or U20493 (N_20493,N_15113,N_13854);
nand U20494 (N_20494,N_12770,N_10045);
nand U20495 (N_20495,N_12656,N_13317);
nand U20496 (N_20496,N_13731,N_10858);
nand U20497 (N_20497,N_11504,N_19191);
nand U20498 (N_20498,N_17313,N_19645);
and U20499 (N_20499,N_19745,N_14204);
nor U20500 (N_20500,N_15684,N_10253);
nor U20501 (N_20501,N_17524,N_17753);
and U20502 (N_20502,N_10792,N_11934);
or U20503 (N_20503,N_14564,N_19971);
nor U20504 (N_20504,N_15655,N_13224);
or U20505 (N_20505,N_14013,N_13213);
nor U20506 (N_20506,N_16137,N_13141);
or U20507 (N_20507,N_10917,N_10141);
nor U20508 (N_20508,N_18389,N_18840);
xnor U20509 (N_20509,N_17347,N_17433);
nor U20510 (N_20510,N_16789,N_15506);
nand U20511 (N_20511,N_18509,N_11725);
nand U20512 (N_20512,N_13552,N_19969);
xor U20513 (N_20513,N_14873,N_19988);
or U20514 (N_20514,N_19010,N_13376);
and U20515 (N_20515,N_19566,N_11638);
or U20516 (N_20516,N_19676,N_10827);
nand U20517 (N_20517,N_17865,N_14006);
and U20518 (N_20518,N_16007,N_14481);
nor U20519 (N_20519,N_10771,N_16556);
nand U20520 (N_20520,N_14247,N_17334);
and U20521 (N_20521,N_16015,N_17376);
nand U20522 (N_20522,N_18810,N_14664);
or U20523 (N_20523,N_16732,N_13724);
nand U20524 (N_20524,N_18276,N_14828);
or U20525 (N_20525,N_19934,N_10589);
xor U20526 (N_20526,N_11247,N_14351);
nand U20527 (N_20527,N_14756,N_10429);
and U20528 (N_20528,N_10280,N_13489);
and U20529 (N_20529,N_16765,N_11576);
xor U20530 (N_20530,N_10914,N_14407);
or U20531 (N_20531,N_15623,N_10177);
or U20532 (N_20532,N_18571,N_16706);
or U20533 (N_20533,N_12302,N_15587);
nor U20534 (N_20534,N_15198,N_17403);
nand U20535 (N_20535,N_18534,N_10361);
and U20536 (N_20536,N_15607,N_19099);
or U20537 (N_20537,N_16748,N_17597);
or U20538 (N_20538,N_17657,N_17894);
or U20539 (N_20539,N_16328,N_19940);
nand U20540 (N_20540,N_13004,N_16292);
nand U20541 (N_20541,N_11228,N_19693);
nand U20542 (N_20542,N_12802,N_12189);
nor U20543 (N_20543,N_13116,N_12232);
and U20544 (N_20544,N_12353,N_14137);
nand U20545 (N_20545,N_12080,N_14083);
nand U20546 (N_20546,N_18258,N_16791);
nor U20547 (N_20547,N_11348,N_16839);
and U20548 (N_20548,N_10997,N_17139);
or U20549 (N_20549,N_16061,N_10664);
nor U20550 (N_20550,N_11912,N_13331);
or U20551 (N_20551,N_15194,N_12683);
xnor U20552 (N_20552,N_15454,N_16021);
nor U20553 (N_20553,N_12470,N_17646);
and U20554 (N_20554,N_10657,N_17660);
or U20555 (N_20555,N_13608,N_12922);
nand U20556 (N_20556,N_15529,N_18519);
and U20557 (N_20557,N_15422,N_10217);
nor U20558 (N_20558,N_11944,N_13610);
nor U20559 (N_20559,N_17285,N_14790);
nand U20560 (N_20560,N_14074,N_10240);
nand U20561 (N_20561,N_16454,N_10084);
nand U20562 (N_20562,N_12960,N_10695);
and U20563 (N_20563,N_12161,N_17496);
or U20564 (N_20564,N_15343,N_15227);
and U20565 (N_20565,N_13737,N_17891);
or U20566 (N_20566,N_18507,N_13425);
nand U20567 (N_20567,N_13643,N_15345);
xor U20568 (N_20568,N_13911,N_16686);
or U20569 (N_20569,N_15191,N_10528);
nor U20570 (N_20570,N_15626,N_17386);
nand U20571 (N_20571,N_11831,N_14482);
and U20572 (N_20572,N_15873,N_14301);
or U20573 (N_20573,N_15758,N_18398);
nand U20574 (N_20574,N_18626,N_10520);
or U20575 (N_20575,N_11374,N_10201);
and U20576 (N_20576,N_15231,N_16783);
nand U20577 (N_20577,N_15633,N_14701);
and U20578 (N_20578,N_11324,N_12041);
nand U20579 (N_20579,N_15862,N_11937);
and U20580 (N_20580,N_19558,N_15759);
nand U20581 (N_20581,N_16124,N_19660);
or U20582 (N_20582,N_17027,N_16170);
or U20583 (N_20583,N_13755,N_13782);
and U20584 (N_20584,N_19757,N_10207);
nor U20585 (N_20585,N_12623,N_17036);
and U20586 (N_20586,N_15704,N_16644);
and U20587 (N_20587,N_12996,N_13038);
nand U20588 (N_20588,N_17249,N_11724);
nor U20589 (N_20589,N_18654,N_12974);
nand U20590 (N_20590,N_13201,N_11134);
nor U20591 (N_20591,N_11756,N_10703);
or U20592 (N_20592,N_17333,N_13022);
and U20593 (N_20593,N_10562,N_12422);
nand U20594 (N_20594,N_10415,N_11688);
or U20595 (N_20595,N_15412,N_16053);
or U20596 (N_20596,N_11115,N_11321);
nor U20597 (N_20597,N_15291,N_10778);
nand U20598 (N_20598,N_14502,N_19849);
nor U20599 (N_20599,N_18857,N_13353);
and U20600 (N_20600,N_12468,N_18424);
and U20601 (N_20601,N_14955,N_13517);
nor U20602 (N_20602,N_10420,N_13908);
and U20603 (N_20603,N_17015,N_11587);
and U20604 (N_20604,N_14959,N_19019);
and U20605 (N_20605,N_10042,N_15147);
nor U20606 (N_20606,N_18544,N_13959);
nor U20607 (N_20607,N_18449,N_18776);
xor U20608 (N_20608,N_13171,N_14257);
nor U20609 (N_20609,N_10855,N_15846);
xnor U20610 (N_20610,N_19824,N_19659);
nand U20611 (N_20611,N_17752,N_14336);
nand U20612 (N_20612,N_12693,N_18023);
nand U20613 (N_20613,N_18408,N_10831);
or U20614 (N_20614,N_11298,N_11302);
nor U20615 (N_20615,N_14781,N_10156);
xnor U20616 (N_20616,N_18589,N_12896);
or U20617 (N_20617,N_14871,N_14795);
or U20618 (N_20618,N_15844,N_18678);
or U20619 (N_20619,N_18150,N_13851);
or U20620 (N_20620,N_15811,N_16675);
nand U20621 (N_20621,N_16362,N_13461);
nand U20622 (N_20622,N_18956,N_19816);
nand U20623 (N_20623,N_11891,N_16372);
and U20624 (N_20624,N_14727,N_12349);
or U20625 (N_20625,N_11354,N_15794);
and U20626 (N_20626,N_12687,N_15625);
nand U20627 (N_20627,N_13453,N_15369);
or U20628 (N_20628,N_15542,N_10212);
and U20629 (N_20629,N_10865,N_11293);
xor U20630 (N_20630,N_12039,N_14740);
and U20631 (N_20631,N_18411,N_10508);
nand U20632 (N_20632,N_19939,N_14341);
and U20633 (N_20633,N_10388,N_13368);
or U20634 (N_20634,N_16870,N_14212);
nor U20635 (N_20635,N_15948,N_16689);
nor U20636 (N_20636,N_11565,N_19999);
or U20637 (N_20637,N_14109,N_15012);
or U20638 (N_20638,N_13058,N_14429);
or U20639 (N_20639,N_11696,N_10770);
nand U20640 (N_20640,N_13604,N_14318);
nor U20641 (N_20641,N_16979,N_14854);
xnor U20642 (N_20642,N_10815,N_11851);
nor U20643 (N_20643,N_12447,N_16189);
or U20644 (N_20644,N_11297,N_15411);
xor U20645 (N_20645,N_16497,N_15997);
nand U20646 (N_20646,N_15385,N_18118);
nor U20647 (N_20647,N_15358,N_19621);
and U20648 (N_20648,N_10451,N_15634);
nand U20649 (N_20649,N_15059,N_12352);
or U20650 (N_20650,N_14326,N_13229);
nor U20651 (N_20651,N_18696,N_10840);
and U20652 (N_20652,N_14060,N_15419);
and U20653 (N_20653,N_17573,N_16133);
and U20654 (N_20654,N_10721,N_16628);
and U20655 (N_20655,N_10360,N_12750);
nand U20656 (N_20656,N_18427,N_14017);
or U20657 (N_20657,N_17000,N_13870);
and U20658 (N_20658,N_14807,N_17451);
and U20659 (N_20659,N_18283,N_11313);
xnor U20660 (N_20660,N_18096,N_18637);
or U20661 (N_20661,N_16059,N_17697);
nor U20662 (N_20662,N_14754,N_15330);
and U20663 (N_20663,N_17109,N_17782);
nor U20664 (N_20664,N_18694,N_12666);
xnor U20665 (N_20665,N_12796,N_12297);
and U20666 (N_20666,N_15999,N_10089);
and U20667 (N_20667,N_15670,N_18420);
or U20668 (N_20668,N_17295,N_16077);
nor U20669 (N_20669,N_11468,N_15556);
and U20670 (N_20670,N_13820,N_18781);
nor U20671 (N_20671,N_12170,N_16983);
and U20672 (N_20672,N_11797,N_14810);
nand U20673 (N_20673,N_15870,N_14320);
xnor U20674 (N_20674,N_17939,N_19784);
nand U20675 (N_20675,N_10542,N_19381);
nand U20676 (N_20676,N_16303,N_11013);
nor U20677 (N_20677,N_14900,N_13741);
xnor U20678 (N_20678,N_14782,N_17988);
xor U20679 (N_20679,N_15392,N_13089);
or U20680 (N_20680,N_15470,N_19644);
xnor U20681 (N_20681,N_15062,N_19569);
nor U20682 (N_20682,N_18351,N_11180);
xnor U20683 (N_20683,N_19132,N_13684);
and U20684 (N_20684,N_12734,N_18194);
xor U20685 (N_20685,N_16773,N_15554);
and U20686 (N_20686,N_19496,N_18709);
nor U20687 (N_20687,N_17359,N_11994);
and U20688 (N_20688,N_13506,N_17094);
or U20689 (N_20689,N_18977,N_15019);
and U20690 (N_20690,N_16247,N_11282);
nor U20691 (N_20691,N_17801,N_19765);
or U20692 (N_20692,N_12289,N_13210);
and U20693 (N_20693,N_15217,N_18978);
nand U20694 (N_20694,N_14758,N_13982);
or U20695 (N_20695,N_15151,N_18905);
nor U20696 (N_20696,N_16614,N_19414);
nand U20697 (N_20697,N_12878,N_18808);
and U20698 (N_20698,N_14415,N_10348);
and U20699 (N_20699,N_19226,N_19684);
nand U20700 (N_20700,N_17143,N_13486);
nand U20701 (N_20701,N_18457,N_12385);
or U20702 (N_20702,N_12743,N_11493);
nor U20703 (N_20703,N_11634,N_16609);
and U20704 (N_20704,N_13537,N_15082);
nand U20705 (N_20705,N_19339,N_11342);
or U20706 (N_20706,N_13420,N_16923);
nand U20707 (N_20707,N_15292,N_13857);
or U20708 (N_20708,N_11042,N_13951);
nand U20709 (N_20709,N_17110,N_16535);
or U20710 (N_20710,N_19227,N_13342);
or U20711 (N_20711,N_15315,N_14672);
or U20712 (N_20712,N_12595,N_12632);
nand U20713 (N_20713,N_13157,N_10880);
and U20714 (N_20714,N_16058,N_12142);
and U20715 (N_20715,N_14366,N_19095);
or U20716 (N_20716,N_18881,N_17519);
nor U20717 (N_20717,N_13965,N_18388);
and U20718 (N_20718,N_19295,N_14080);
nand U20719 (N_20719,N_17126,N_14601);
nand U20720 (N_20720,N_10241,N_16795);
or U20721 (N_20721,N_11267,N_11911);
and U20722 (N_20722,N_10924,N_15309);
or U20723 (N_20723,N_13375,N_13827);
xor U20724 (N_20724,N_10902,N_14460);
and U20725 (N_20725,N_17743,N_18158);
nor U20726 (N_20726,N_14128,N_16876);
nor U20727 (N_20727,N_11673,N_16709);
nor U20728 (N_20728,N_14780,N_11902);
nor U20729 (N_20729,N_12901,N_12805);
xnor U20730 (N_20730,N_15047,N_10307);
or U20731 (N_20731,N_12846,N_10668);
and U20732 (N_20732,N_17629,N_13667);
nor U20733 (N_20733,N_11336,N_11382);
or U20734 (N_20734,N_14089,N_17628);
nand U20735 (N_20735,N_12838,N_16615);
xnor U20736 (N_20736,N_19133,N_11760);
nor U20737 (N_20737,N_12407,N_15892);
nand U20738 (N_20738,N_15175,N_16878);
and U20739 (N_20739,N_17783,N_15288);
or U20740 (N_20740,N_18204,N_16575);
xnor U20741 (N_20741,N_19120,N_15574);
and U20742 (N_20742,N_10503,N_12114);
nor U20743 (N_20743,N_11263,N_11459);
or U20744 (N_20744,N_12941,N_12633);
nor U20745 (N_20745,N_16460,N_11957);
and U20746 (N_20746,N_18315,N_13937);
nand U20747 (N_20747,N_19481,N_19458);
and U20748 (N_20748,N_13838,N_17876);
nand U20749 (N_20749,N_13017,N_15316);
and U20750 (N_20750,N_15666,N_12198);
nand U20751 (N_20751,N_14496,N_17908);
or U20752 (N_20752,N_16519,N_15393);
nand U20753 (N_20753,N_15947,N_12740);
and U20754 (N_20754,N_16284,N_14933);
nand U20755 (N_20755,N_18972,N_15399);
nand U20756 (N_20756,N_19200,N_12125);
xor U20757 (N_20757,N_17520,N_14579);
or U20758 (N_20758,N_18588,N_13932);
or U20759 (N_20759,N_16648,N_15110);
nand U20760 (N_20760,N_11678,N_16215);
xnor U20761 (N_20761,N_14935,N_12503);
and U20762 (N_20762,N_19012,N_10995);
and U20763 (N_20763,N_17043,N_11979);
xor U20764 (N_20764,N_14262,N_16343);
nor U20765 (N_20765,N_18785,N_17158);
and U20766 (N_20766,N_16070,N_17881);
and U20767 (N_20767,N_12449,N_15342);
and U20768 (N_20768,N_16723,N_12431);
or U20769 (N_20769,N_17899,N_10443);
nor U20770 (N_20770,N_12115,N_12488);
nand U20771 (N_20771,N_10741,N_17740);
nand U20772 (N_20772,N_10898,N_11165);
nor U20773 (N_20773,N_12699,N_10724);
nand U20774 (N_20774,N_19478,N_17764);
nor U20775 (N_20775,N_18993,N_17130);
and U20776 (N_20776,N_17448,N_16739);
and U20777 (N_20777,N_10248,N_16245);
or U20778 (N_20778,N_18581,N_10393);
nand U20779 (N_20779,N_16095,N_13232);
xor U20780 (N_20780,N_11034,N_11113);
or U20781 (N_20781,N_10478,N_19657);
nand U20782 (N_20782,N_18852,N_15079);
nor U20783 (N_20783,N_17038,N_14938);
nand U20784 (N_20784,N_18473,N_12308);
xor U20785 (N_20785,N_15265,N_19246);
nor U20786 (N_20786,N_11306,N_18197);
and U20787 (N_20787,N_14731,N_14160);
nand U20788 (N_20788,N_13995,N_19499);
nor U20789 (N_20789,N_18402,N_19348);
or U20790 (N_20790,N_10012,N_17259);
or U20791 (N_20791,N_18027,N_17019);
nor U20792 (N_20792,N_11163,N_11280);
xor U20793 (N_20793,N_17884,N_11580);
or U20794 (N_20794,N_10629,N_15533);
or U20795 (N_20795,N_12230,N_10321);
or U20796 (N_20796,N_19582,N_12137);
nand U20797 (N_20797,N_17173,N_18343);
nand U20798 (N_20798,N_18898,N_14587);
nand U20799 (N_20799,N_13451,N_15521);
nor U20800 (N_20800,N_12013,N_19548);
or U20801 (N_20801,N_16751,N_18548);
and U20802 (N_20802,N_17654,N_14483);
and U20803 (N_20803,N_14142,N_16966);
or U20804 (N_20804,N_19607,N_10023);
xor U20805 (N_20805,N_19908,N_12123);
or U20806 (N_20806,N_18935,N_17405);
or U20807 (N_20807,N_18146,N_16325);
xor U20808 (N_20808,N_19557,N_13128);
nor U20809 (N_20809,N_10378,N_17762);
nor U20810 (N_20810,N_18009,N_11235);
and U20811 (N_20811,N_16833,N_17833);
nor U20812 (N_20812,N_16013,N_10639);
or U20813 (N_20813,N_13003,N_19870);
nand U20814 (N_20814,N_15238,N_13818);
nand U20815 (N_20815,N_17968,N_18471);
or U20816 (N_20816,N_16429,N_12997);
nand U20817 (N_20817,N_12176,N_14591);
nand U20818 (N_20818,N_14730,N_13787);
or U20819 (N_20819,N_14117,N_12281);
or U20820 (N_20820,N_13950,N_15866);
xor U20821 (N_20821,N_11816,N_16224);
nand U20822 (N_20822,N_14578,N_19169);
xnor U20823 (N_20823,N_16673,N_17033);
nor U20824 (N_20824,N_13925,N_14008);
nand U20825 (N_20825,N_12439,N_11728);
nand U20826 (N_20826,N_14408,N_14158);
nand U20827 (N_20827,N_16947,N_19383);
nor U20828 (N_20828,N_11253,N_15164);
nand U20829 (N_20829,N_14923,N_10409);
nor U20830 (N_20830,N_16559,N_12540);
nor U20831 (N_20831,N_17205,N_12280);
nor U20832 (N_20832,N_13736,N_14530);
nand U20833 (N_20833,N_11307,N_19797);
and U20834 (N_20834,N_13068,N_17254);
or U20835 (N_20835,N_10517,N_13397);
nor U20836 (N_20836,N_11719,N_19915);
nor U20837 (N_20837,N_17817,N_19891);
or U20838 (N_20838,N_19758,N_11104);
nand U20839 (N_20839,N_15415,N_13266);
xor U20840 (N_20840,N_12576,N_13654);
or U20841 (N_20841,N_17612,N_11220);
nand U20842 (N_20842,N_18516,N_12843);
nand U20843 (N_20843,N_10176,N_10092);
and U20844 (N_20844,N_12249,N_12498);
nand U20845 (N_20845,N_11153,N_17852);
or U20846 (N_20846,N_16768,N_10910);
nor U20847 (N_20847,N_16814,N_17732);
and U20848 (N_20848,N_11963,N_16052);
xor U20849 (N_20849,N_14014,N_18051);
xnor U20850 (N_20850,N_13127,N_18615);
and U20851 (N_20851,N_13717,N_10070);
nand U20852 (N_20852,N_11775,N_19959);
and U20853 (N_20853,N_13647,N_19109);
and U20854 (N_20854,N_14925,N_17201);
and U20855 (N_20855,N_13515,N_11537);
or U20856 (N_20856,N_19671,N_13585);
and U20857 (N_20857,N_12158,N_15881);
or U20858 (N_20858,N_15241,N_14501);
and U20859 (N_20859,N_15995,N_17198);
nand U20860 (N_20860,N_18254,N_19759);
or U20861 (N_20861,N_18648,N_12165);
nor U20862 (N_20862,N_15485,N_17845);
and U20863 (N_20863,N_17056,N_14651);
nor U20864 (N_20864,N_11540,N_16745);
and U20865 (N_20865,N_11863,N_19418);
nand U20866 (N_20866,N_10149,N_11618);
or U20867 (N_20867,N_14707,N_11299);
or U20868 (N_20868,N_18488,N_12715);
nor U20869 (N_20869,N_15526,N_14718);
xor U20870 (N_20870,N_17292,N_13790);
xor U20871 (N_20871,N_15613,N_10662);
nor U20872 (N_20872,N_18218,N_11666);
nor U20873 (N_20873,N_15266,N_19228);
and U20874 (N_20874,N_16913,N_12751);
and U20875 (N_20875,N_13606,N_19474);
and U20876 (N_20876,N_11046,N_19790);
or U20877 (N_20877,N_18368,N_12342);
nand U20878 (N_20878,N_15102,N_18700);
or U20879 (N_20879,N_11006,N_11712);
and U20880 (N_20880,N_10067,N_14905);
and U20881 (N_20881,N_17068,N_15335);
and U20882 (N_20882,N_17429,N_15760);
or U20883 (N_20883,N_14170,N_16585);
nor U20884 (N_20884,N_13546,N_13863);
nand U20885 (N_20885,N_13733,N_15956);
xor U20886 (N_20886,N_19139,N_18535);
nand U20887 (N_20887,N_12146,N_10285);
nand U20888 (N_20888,N_18704,N_13660);
nand U20889 (N_20889,N_18690,N_18547);
nor U20890 (N_20890,N_10756,N_16679);
or U20891 (N_20891,N_10624,N_11249);
xor U20892 (N_20892,N_10873,N_13432);
or U20893 (N_20893,N_16109,N_13920);
xnor U20894 (N_20894,N_10399,N_14239);
nand U20895 (N_20895,N_12523,N_11822);
and U20896 (N_20896,N_15681,N_16929);
and U20897 (N_20897,N_14043,N_13247);
nand U20898 (N_20898,N_10390,N_17371);
or U20899 (N_20899,N_16714,N_10033);
nand U20900 (N_20900,N_12890,N_15746);
and U20901 (N_20901,N_15301,N_12070);
xnor U20902 (N_20902,N_18236,N_18459);
nor U20903 (N_20903,N_14639,N_19057);
nand U20904 (N_20904,N_19128,N_16921);
or U20905 (N_20905,N_15410,N_12283);
xnor U20906 (N_20906,N_13024,N_15636);
and U20907 (N_20907,N_16796,N_10258);
and U20908 (N_20908,N_10836,N_12259);
nor U20909 (N_20909,N_15025,N_16617);
xor U20910 (N_20910,N_13312,N_10157);
xor U20911 (N_20911,N_17739,N_18803);
and U20912 (N_20912,N_13150,N_12900);
nand U20913 (N_20913,N_19320,N_19327);
nand U20914 (N_20914,N_13962,N_12381);
or U20915 (N_20915,N_10466,N_14992);
nand U20916 (N_20916,N_15381,N_16121);
or U20917 (N_20917,N_14184,N_13394);
and U20918 (N_20918,N_17806,N_19025);
nor U20919 (N_20919,N_13143,N_11244);
and U20920 (N_20920,N_15080,N_16869);
or U20921 (N_20921,N_11232,N_15511);
xor U20922 (N_20922,N_19020,N_17011);
or U20923 (N_20923,N_19627,N_11442);
and U20924 (N_20924,N_19325,N_16230);
or U20925 (N_20925,N_12630,N_12427);
or U20926 (N_20926,N_15022,N_16314);
nand U20927 (N_20927,N_16173,N_14048);
or U20928 (N_20928,N_12879,N_10637);
nand U20929 (N_20929,N_15968,N_18933);
nand U20930 (N_20930,N_16040,N_19266);
or U20931 (N_20931,N_15508,N_16216);
nand U20932 (N_20932,N_14596,N_15616);
or U20933 (N_20933,N_11095,N_10352);
nor U20934 (N_20934,N_19332,N_13961);
xor U20935 (N_20935,N_16653,N_12237);
nand U20936 (N_20936,N_19937,N_15272);
or U20937 (N_20937,N_12826,N_19465);
nand U20938 (N_20938,N_15294,N_14614);
xor U20939 (N_20939,N_17228,N_16389);
and U20940 (N_20940,N_12046,N_14175);
or U20941 (N_20941,N_17945,N_18752);
nand U20942 (N_20942,N_16564,N_19618);
or U20943 (N_20943,N_16187,N_16199);
nor U20944 (N_20944,N_14229,N_19376);
nor U20945 (N_20945,N_10228,N_15961);
or U20946 (N_20946,N_10916,N_15064);
nand U20947 (N_20947,N_19198,N_10573);
nor U20948 (N_20948,N_15589,N_10678);
and U20949 (N_20949,N_16643,N_15002);
nand U20950 (N_20950,N_11790,N_15658);
nand U20951 (N_20951,N_18490,N_16729);
and U20952 (N_20952,N_15689,N_13817);
nor U20953 (N_20953,N_15365,N_10896);
nor U20954 (N_20954,N_11838,N_14568);
or U20955 (N_20955,N_15207,N_16788);
nand U20956 (N_20956,N_18968,N_12912);
nand U20957 (N_20957,N_14381,N_16511);
xor U20958 (N_20958,N_14713,N_17427);
nand U20959 (N_20959,N_10894,N_16504);
nand U20960 (N_20960,N_14641,N_17400);
nand U20961 (N_20961,N_18822,N_18103);
xnor U20962 (N_20962,N_15974,N_11667);
and U20963 (N_20963,N_14988,N_14338);
and U20964 (N_20964,N_16296,N_12188);
and U20965 (N_20965,N_10435,N_11589);
and U20966 (N_20966,N_13085,N_17564);
nand U20967 (N_20967,N_13108,N_10656);
and U20968 (N_20968,N_11077,N_18359);
and U20969 (N_20969,N_18966,N_17648);
nor U20970 (N_20970,N_13964,N_12859);
or U20971 (N_20971,N_15925,N_16411);
and U20972 (N_20972,N_12256,N_14321);
and U20973 (N_20973,N_18085,N_14019);
xor U20974 (N_20974,N_13246,N_14820);
nor U20975 (N_20975,N_11541,N_13491);
or U20976 (N_20976,N_18133,N_16400);
or U20977 (N_20977,N_14929,N_19655);
xnor U20978 (N_20978,N_19203,N_18681);
or U20979 (N_20979,N_18365,N_13207);
nand U20980 (N_20980,N_16664,N_13968);
nor U20981 (N_20981,N_11843,N_11154);
nor U20982 (N_20982,N_10890,N_18335);
and U20983 (N_20983,N_17595,N_16737);
nor U20984 (N_20984,N_17956,N_19572);
nand U20985 (N_20985,N_19341,N_11642);
and U20986 (N_20986,N_18295,N_16000);
and U20987 (N_20987,N_13015,N_13973);
and U20988 (N_20988,N_10638,N_17471);
or U20989 (N_20989,N_13632,N_12524);
and U20990 (N_20990,N_13277,N_10530);
nor U20991 (N_20991,N_10118,N_10887);
or U20992 (N_20992,N_18833,N_13194);
nand U20993 (N_20993,N_15173,N_14344);
or U20994 (N_20994,N_14414,N_18275);
xnor U20995 (N_20995,N_14837,N_11311);
nand U20996 (N_20996,N_11071,N_11355);
and U20997 (N_20997,N_16080,N_14714);
and U20998 (N_20998,N_14372,N_11000);
or U20999 (N_20999,N_13678,N_12756);
or U21000 (N_21000,N_16974,N_10099);
nor U21001 (N_21001,N_14546,N_10861);
or U21002 (N_21002,N_12032,N_18813);
xor U21003 (N_21003,N_12134,N_11594);
nor U21004 (N_21004,N_15652,N_13447);
and U21005 (N_21005,N_17398,N_19860);
nor U21006 (N_21006,N_13488,N_16453);
and U21007 (N_21007,N_10143,N_14571);
or U21008 (N_21008,N_18182,N_16801);
or U21009 (N_21009,N_19154,N_18376);
nor U21010 (N_21010,N_19732,N_17772);
nand U21011 (N_21011,N_12948,N_15895);
xor U21012 (N_21012,N_11467,N_12647);
nand U21013 (N_21013,N_15851,N_13844);
xnor U21014 (N_21014,N_19782,N_15597);
or U21015 (N_21015,N_13197,N_11213);
nand U21016 (N_21016,N_11543,N_15189);
nor U21017 (N_21017,N_16806,N_17875);
and U21018 (N_21018,N_19527,N_13577);
and U21019 (N_21019,N_17675,N_12665);
nor U21020 (N_21020,N_10923,N_15465);
and U21021 (N_21021,N_13700,N_18164);
nor U21022 (N_21022,N_11458,N_15624);
and U21023 (N_21023,N_16573,N_16469);
nor U21024 (N_21024,N_19795,N_18090);
or U21025 (N_21025,N_16627,N_17926);
and U21026 (N_21026,N_15063,N_11200);
or U21027 (N_21027,N_10484,N_18605);
and U21028 (N_21028,N_11075,N_17460);
and U21029 (N_21029,N_10462,N_11152);
nand U21030 (N_21030,N_17991,N_17975);
and U21031 (N_21031,N_12703,N_14113);
nor U21032 (N_21032,N_12874,N_17266);
and U21033 (N_21033,N_15039,N_10790);
nor U21034 (N_21034,N_13217,N_14486);
xor U21035 (N_21035,N_12242,N_10786);
and U21036 (N_21036,N_11439,N_11941);
and U21037 (N_21037,N_13570,N_10326);
and U21038 (N_21038,N_15790,N_11123);
nand U21039 (N_21039,N_17679,N_15098);
nor U21040 (N_21040,N_14273,N_16281);
or U21041 (N_21041,N_11384,N_17632);
and U21042 (N_21042,N_10044,N_18502);
or U21043 (N_21043,N_14950,N_16265);
and U21044 (N_21044,N_16782,N_11363);
or U21045 (N_21045,N_17615,N_17335);
nor U21046 (N_21046,N_10801,N_12676);
or U21047 (N_21047,N_16540,N_11987);
or U21048 (N_21048,N_13773,N_10883);
or U21049 (N_21049,N_13975,N_16033);
and U21050 (N_21050,N_16633,N_17730);
xnor U21051 (N_21051,N_14264,N_12139);
or U21052 (N_21052,N_15858,N_11452);
xor U21053 (N_21053,N_11652,N_12477);
nor U21054 (N_21054,N_15572,N_12555);
and U21055 (N_21055,N_19877,N_17065);
nand U21056 (N_21056,N_13438,N_13711);
or U21057 (N_21057,N_13934,N_16539);
xnor U21058 (N_21058,N_18923,N_19296);
xor U21059 (N_21059,N_11914,N_12075);
xor U21060 (N_21060,N_16692,N_18081);
nand U21061 (N_21061,N_17255,N_18676);
or U21062 (N_21062,N_16742,N_11992);
nor U21063 (N_21063,N_14495,N_17990);
nor U21064 (N_21064,N_16649,N_10791);
nand U21065 (N_21065,N_13274,N_19367);
or U21066 (N_21066,N_19856,N_11396);
or U21067 (N_21067,N_11207,N_12388);
nand U21068 (N_21068,N_11683,N_16702);
nand U21069 (N_21069,N_19401,N_18596);
and U21070 (N_21070,N_19403,N_12962);
nand U21071 (N_21071,N_14555,N_19177);
xnor U21072 (N_21072,N_11065,N_15220);
or U21073 (N_21073,N_12636,N_12270);
xor U21074 (N_21074,N_18695,N_14447);
nand U21075 (N_21075,N_16902,N_18310);
nand U21076 (N_21076,N_16441,N_12721);
or U21077 (N_21077,N_15475,N_11625);
nor U21078 (N_21078,N_18213,N_18374);
nand U21079 (N_21079,N_14190,N_18743);
or U21080 (N_21080,N_12961,N_17650);
or U21081 (N_21081,N_16366,N_11516);
and U21082 (N_21082,N_14660,N_17581);
or U21083 (N_21083,N_12939,N_15825);
and U21084 (N_21084,N_13359,N_14903);
nor U21085 (N_21085,N_10262,N_18269);
nand U21086 (N_21086,N_18985,N_15258);
nor U21087 (N_21087,N_15246,N_15447);
nand U21088 (N_21088,N_15352,N_12469);
or U21089 (N_21089,N_16755,N_18070);
nand U21090 (N_21090,N_15431,N_10003);
or U21091 (N_21091,N_14613,N_16772);
or U21092 (N_21092,N_13370,N_11377);
nand U21093 (N_21093,N_18167,N_16200);
or U21094 (N_21094,N_17446,N_12517);
or U21095 (N_21095,N_12127,N_15774);
or U21096 (N_21096,N_11945,N_11370);
or U21097 (N_21097,N_14515,N_17588);
and U21098 (N_21098,N_17979,N_16447);
or U21099 (N_21099,N_14053,N_12023);
and U21100 (N_21100,N_10282,N_12608);
and U21101 (N_21101,N_18298,N_13212);
nor U21102 (N_21102,N_15053,N_10145);
xor U21103 (N_21103,N_17316,N_17356);
or U21104 (N_21104,N_11771,N_17553);
nor U21105 (N_21105,N_14497,N_12076);
nand U21106 (N_21106,N_10203,N_11868);
or U21107 (N_21107,N_11959,N_12164);
and U21108 (N_21108,N_19103,N_14606);
or U21109 (N_21109,N_16347,N_17006);
or U21110 (N_21110,N_14474,N_19581);
nand U21111 (N_21111,N_17118,N_15478);
nor U21112 (N_21112,N_10502,N_10457);
nor U21113 (N_21113,N_19264,N_12771);
nor U21114 (N_21114,N_16512,N_11438);
or U21115 (N_21115,N_10180,N_15706);
and U21116 (N_21116,N_10355,N_13444);
or U21117 (N_21117,N_19006,N_16370);
nor U21118 (N_21118,N_13993,N_15017);
nand U21119 (N_21119,N_12122,N_16641);
xnor U21120 (N_21120,N_18902,N_18297);
and U21121 (N_21121,N_11050,N_12117);
and U21122 (N_21122,N_13841,N_11371);
or U21123 (N_21123,N_18256,N_11753);
xor U21124 (N_21124,N_14995,N_15909);
xor U21125 (N_21125,N_16257,N_13470);
and U21126 (N_21126,N_11048,N_18698);
or U21127 (N_21127,N_10641,N_14866);
nor U21128 (N_21128,N_18466,N_16925);
and U21129 (N_21129,N_19238,N_12133);
or U21130 (N_21130,N_19623,N_12084);
nor U21131 (N_21131,N_14395,N_10736);
and U21132 (N_21132,N_10652,N_13132);
nor U21133 (N_21133,N_12008,N_13550);
nor U21134 (N_21134,N_13786,N_12931);
nor U21135 (N_21135,N_10423,N_10057);
xor U21136 (N_21136,N_15531,N_13231);
nor U21137 (N_21137,N_11429,N_17857);
nor U21138 (N_21138,N_14695,N_19283);
and U21139 (N_21139,N_19719,N_16168);
nand U21140 (N_21140,N_12428,N_13742);
nor U21141 (N_21141,N_19290,N_18064);
nand U21142 (N_21142,N_14186,N_14202);
or U21143 (N_21143,N_15133,N_14149);
nor U21144 (N_21144,N_14024,N_10901);
nor U21145 (N_21145,N_19326,N_14155);
nor U21146 (N_21146,N_18083,N_19652);
xnor U21147 (N_21147,N_19954,N_18927);
nand U21148 (N_21148,N_10113,N_11586);
and U21149 (N_21149,N_14478,N_13635);
nor U21150 (N_21150,N_18851,N_13977);
nor U21151 (N_21151,N_15818,N_16828);
nand U21152 (N_21152,N_15219,N_18619);
xnor U21153 (N_21153,N_18559,N_12099);
nand U21154 (N_21154,N_10766,N_19404);
and U21155 (N_21155,N_11573,N_11659);
and U21156 (N_21156,N_11135,N_16688);
and U21157 (N_21157,N_17208,N_14561);
xor U21158 (N_21158,N_11008,N_18540);
nor U21159 (N_21159,N_19172,N_10060);
nor U21160 (N_21160,N_16901,N_14005);
and U21161 (N_21161,N_19729,N_18912);
xnor U21162 (N_21162,N_17971,N_10094);
and U21163 (N_21163,N_16083,N_18279);
nor U21164 (N_21164,N_19351,N_17300);
nor U21165 (N_21165,N_11876,N_14337);
nor U21166 (N_21166,N_16740,N_14373);
nor U21167 (N_21167,N_16489,N_12118);
nand U21168 (N_21168,N_14676,N_17485);
xor U21169 (N_21169,N_13799,N_19904);
and U21170 (N_21170,N_15209,N_10261);
and U21171 (N_21171,N_12460,N_10735);
nand U21172 (N_21172,N_14671,N_15856);
and U21173 (N_21173,N_18762,N_10585);
xor U21174 (N_21174,N_17692,N_14583);
xnor U21175 (N_21175,N_10609,N_11588);
and U21176 (N_21176,N_14288,N_19933);
nand U21177 (N_21177,N_16254,N_15770);
nor U21178 (N_21178,N_19895,N_19307);
nand U21179 (N_21179,N_10716,N_11549);
or U21180 (N_21180,N_14056,N_11203);
nand U21181 (N_21181,N_16226,N_10553);
or U21182 (N_21182,N_13500,N_12500);
and U21183 (N_21183,N_13695,N_18701);
and U21184 (N_21184,N_19707,N_19793);
nand U21185 (N_21185,N_18950,N_10852);
or U21186 (N_21186,N_10495,N_14922);
or U21187 (N_21187,N_10471,N_19013);
nand U21188 (N_21188,N_17757,N_18649);
and U21189 (N_21189,N_14766,N_10014);
nand U21190 (N_21190,N_14086,N_13458);
and U21191 (N_21191,N_18290,N_16312);
nand U21192 (N_21192,N_14677,N_13190);
xnor U21193 (N_21193,N_11668,N_12679);
nor U21194 (N_21194,N_18474,N_10368);
nor U21195 (N_21195,N_19651,N_19251);
or U21196 (N_21196,N_13882,N_11221);
xnor U21197 (N_21197,N_14654,N_16834);
and U21198 (N_21198,N_16180,N_11946);
and U21199 (N_21199,N_13739,N_18013);
nor U21200 (N_21200,N_10224,N_12443);
or U21201 (N_21201,N_13200,N_18839);
xor U21202 (N_21202,N_15736,N_11932);
nor U21203 (N_21203,N_12869,N_15159);
or U21204 (N_21204,N_17102,N_16248);
and U21205 (N_21205,N_13578,N_13020);
nand U21206 (N_21206,N_19990,N_15719);
nand U21207 (N_21207,N_17196,N_12818);
and U21208 (N_21208,N_14102,N_11989);
nor U21209 (N_21209,N_16659,N_15697);
nand U21210 (N_21210,N_10316,N_14842);
nand U21211 (N_21211,N_14131,N_16613);
xor U21212 (N_21212,N_13441,N_10586);
xor U21213 (N_21213,N_17703,N_16998);
nand U21214 (N_21214,N_14436,N_19931);
and U21215 (N_21215,N_11111,N_15222);
nand U21216 (N_21216,N_15091,N_16588);
nand U21217 (N_21217,N_13605,N_14744);
and U21218 (N_21218,N_10714,N_10499);
and U21219 (N_21219,N_18208,N_18569);
and U21220 (N_21220,N_16088,N_14619);
nor U21221 (N_21221,N_18591,N_11155);
nor U21222 (N_21222,N_17847,N_10186);
nor U21223 (N_21223,N_15112,N_16928);
nor U21224 (N_21224,N_17075,N_13826);
nor U21225 (N_21225,N_19788,N_16566);
and U21226 (N_21226,N_15084,N_14691);
and U21227 (N_21227,N_15202,N_19899);
nand U21228 (N_21228,N_18529,N_14463);
nand U21229 (N_21229,N_14572,N_10061);
or U21230 (N_21230,N_16359,N_19256);
or U21231 (N_21231,N_11053,N_12390);
xnor U21232 (N_21232,N_18212,N_14041);
and U21233 (N_21233,N_11059,N_12907);
or U21234 (N_21234,N_14121,N_17001);
nor U21235 (N_21235,N_18757,N_18198);
nand U21236 (N_21236,N_15467,N_17721);
and U21237 (N_21237,N_15690,N_16821);
or U21238 (N_21238,N_10030,N_11288);
nor U21239 (N_21239,N_18280,N_11066);
nand U21240 (N_21240,N_11713,N_12620);
nand U21241 (N_21241,N_15376,N_10539);
xnor U21242 (N_21242,N_15237,N_14937);
nand U21243 (N_21243,N_18574,N_10446);
or U21244 (N_21244,N_12744,N_17769);
and U21245 (N_21245,N_15967,N_15973);
nand U21246 (N_21246,N_14433,N_18016);
or U21247 (N_21247,N_12942,N_10309);
nor U21248 (N_21248,N_15370,N_12224);
nand U21249 (N_21249,N_17744,N_14335);
and U21250 (N_21250,N_17200,N_18613);
or U21251 (N_21251,N_12924,N_17954);
or U21252 (N_21252,N_12452,N_14918);
or U21253 (N_21253,N_19156,N_16997);
xnor U21254 (N_21254,N_12789,N_17406);
nor U21255 (N_21255,N_10740,N_10787);
or U21256 (N_21256,N_10076,N_18277);
or U21257 (N_21257,N_10385,N_15027);
xnor U21258 (N_21258,N_19839,N_13062);
or U21259 (N_21259,N_12940,N_19918);
nand U21260 (N_21260,N_14948,N_14799);
and U21261 (N_21261,N_18921,N_15329);
or U21262 (N_21262,N_14220,N_11927);
nand U21263 (N_21263,N_18362,N_10682);
nor U21264 (N_21264,N_13549,N_17965);
nor U21265 (N_21265,N_12698,N_12973);
or U21266 (N_21266,N_19111,N_16708);
nor U21267 (N_21267,N_17861,N_11037);
and U21268 (N_21268,N_16822,N_12368);
nor U21269 (N_21269,N_16577,N_11607);
nor U21270 (N_21270,N_17128,N_16724);
nor U21271 (N_21271,N_13707,N_19011);
nor U21272 (N_21272,N_14375,N_17513);
or U21273 (N_21273,N_14961,N_19127);
and U21274 (N_21274,N_14505,N_10660);
nor U21275 (N_21275,N_16098,N_13332);
nor U21276 (N_21276,N_13158,N_18382);
nand U21277 (N_21277,N_10117,N_11174);
nand U21278 (N_21278,N_15660,N_14755);
and U21279 (N_21279,N_18462,N_11804);
and U21280 (N_21280,N_18773,N_13689);
xnor U21281 (N_21281,N_13631,N_16611);
nor U21282 (N_21282,N_17176,N_19786);
nor U21283 (N_21283,N_11999,N_17584);
nor U21284 (N_21284,N_11176,N_16377);
xnor U21285 (N_21285,N_17442,N_11752);
xor U21286 (N_21286,N_19512,N_19157);
and U21287 (N_21287,N_18338,N_18093);
xor U21288 (N_21288,N_18618,N_17449);
and U21289 (N_21289,N_15363,N_16274);
xnor U21290 (N_21290,N_12781,N_14844);
xor U21291 (N_21291,N_14386,N_10171);
and U21292 (N_21292,N_13861,N_19225);
xor U21293 (N_21293,N_17537,N_12102);
or U21294 (N_21294,N_15582,N_10627);
nand U21295 (N_21295,N_12244,N_10431);
nor U21296 (N_21296,N_18041,N_19596);
and U21297 (N_21297,N_19045,N_13094);
or U21298 (N_21298,N_10760,N_11476);
or U21299 (N_21299,N_18363,N_14919);
or U21300 (N_21300,N_15933,N_10041);
xnor U21301 (N_21301,N_12210,N_18988);
nand U21302 (N_21302,N_15879,N_18877);
nor U21303 (N_21303,N_18226,N_12411);
or U21304 (N_21304,N_17587,N_17687);
nand U21305 (N_21305,N_11252,N_10842);
nand U21306 (N_21306,N_11939,N_12587);
xnor U21307 (N_21307,N_11456,N_15855);
or U21308 (N_21308,N_16132,N_10296);
and U21309 (N_21309,N_16203,N_17268);
or U21310 (N_21310,N_15792,N_16100);
xor U21311 (N_21311,N_15664,N_13686);
or U21312 (N_21312,N_10623,N_11566);
nor U21313 (N_21313,N_11105,N_16227);
or U21314 (N_21314,N_17312,N_19977);
nor U21315 (N_21315,N_18918,N_14181);
nor U21316 (N_21316,N_10558,N_16984);
or U21317 (N_21317,N_16960,N_17663);
and U21318 (N_21318,N_14029,N_11036);
nand U21319 (N_21319,N_11281,N_13969);
or U21320 (N_21320,N_18005,N_16894);
and U21321 (N_21321,N_15360,N_11693);
and U21322 (N_21322,N_13263,N_11497);
or U21323 (N_21323,N_17479,N_19778);
or U21324 (N_21324,N_16895,N_15274);
and U21325 (N_21325,N_18989,N_16712);
nor U21326 (N_21326,N_13400,N_14604);
nor U21327 (N_21327,N_13812,N_15737);
nand U21328 (N_21328,N_18531,N_19492);
nor U21329 (N_21329,N_11918,N_19700);
nand U21330 (N_21330,N_19232,N_15199);
nand U21331 (N_21331,N_15620,N_14409);
nand U21332 (N_21332,N_12462,N_19094);
xnor U21333 (N_21333,N_19540,N_14791);
nor U21334 (N_21334,N_12949,N_17469);
or U21335 (N_21335,N_14769,N_18489);
and U21336 (N_21336,N_18321,N_17736);
and U21337 (N_21337,N_17601,N_19922);
nand U21338 (N_21338,N_11590,N_13082);
and U21339 (N_21339,N_13468,N_15321);
and U21340 (N_21340,N_17461,N_17838);
nor U21341 (N_21341,N_13760,N_15095);
and U21342 (N_21342,N_16326,N_13727);
and U21343 (N_21343,N_15071,N_15013);
nand U21344 (N_21344,N_18570,N_10794);
and U21345 (N_21345,N_12640,N_15143);
nand U21346 (N_21346,N_15109,N_12298);
or U21347 (N_21347,N_15738,N_13336);
nor U21348 (N_21348,N_16835,N_11644);
or U21349 (N_21349,N_15169,N_11069);
or U21350 (N_21350,N_18015,N_16354);
nand U21351 (N_21351,N_11766,N_10701);
or U21352 (N_21352,N_11748,N_19087);
nor U21353 (N_21353,N_10533,N_15713);
or U21354 (N_21354,N_16560,N_13321);
nand U21355 (N_21355,N_15819,N_12050);
or U21356 (N_21356,N_10798,N_13487);
nor U21357 (N_21357,N_14453,N_17470);
nor U21358 (N_21358,N_18141,N_10738);
and U21359 (N_21359,N_11901,N_18019);
and U21360 (N_21360,N_17293,N_18862);
or U21361 (N_21361,N_18819,N_16022);
nand U21362 (N_21362,N_10251,N_14287);
and U21363 (N_21363,N_11984,N_17087);
xnor U21364 (N_21364,N_12998,N_17775);
xor U21365 (N_21365,N_14065,N_15724);
nor U21366 (N_21366,N_15721,N_13954);
and U21367 (N_21367,N_12695,N_18625);
nand U21368 (N_21368,N_14139,N_10375);
xor U21369 (N_21369,N_10022,N_14274);
and U21370 (N_21370,N_19342,N_12093);
nor U21371 (N_21371,N_10857,N_14112);
nand U21372 (N_21372,N_13221,N_10278);
nand U21373 (N_21373,N_11749,N_10202);
nand U21374 (N_21374,N_16020,N_16786);
and U21375 (N_21375,N_12821,N_18717);
nor U21376 (N_21376,N_17310,N_15334);
nand U21377 (N_21377,N_10211,N_19888);
xnor U21378 (N_21378,N_11047,N_17004);
and U21379 (N_21379,N_18616,N_18684);
or U21380 (N_21380,N_11136,N_19036);
or U21381 (N_21381,N_13381,N_19522);
nand U21382 (N_21382,N_15918,N_14817);
and U21383 (N_21383,N_15861,N_11879);
xor U21384 (N_21384,N_13244,N_11502);
nand U21385 (N_21385,N_19259,N_19926);
xor U21386 (N_21386,N_14488,N_11091);
or U21387 (N_21387,N_17600,N_16850);
nand U21388 (N_21388,N_11900,N_17499);
nor U21389 (N_21389,N_12993,N_10397);
xnor U21390 (N_21390,N_16606,N_14882);
or U21391 (N_21391,N_16357,N_18033);
or U21392 (N_21392,N_18183,N_19254);
or U21393 (N_21393,N_16293,N_14537);
nor U21394 (N_21394,N_17637,N_18682);
and U21395 (N_21395,N_17711,N_13758);
and U21396 (N_21396,N_19402,N_11308);
or U21397 (N_21397,N_11692,N_11907);
nor U21398 (N_21398,N_16176,N_11350);
nand U21399 (N_21399,N_10922,N_18890);
or U21400 (N_21400,N_16531,N_14130);
xor U21401 (N_21401,N_13984,N_12441);
nor U21402 (N_21402,N_13395,N_17754);
and U21403 (N_21403,N_11817,N_11496);
and U21404 (N_21404,N_17108,N_19164);
nand U21405 (N_21405,N_14291,N_17904);
and U21406 (N_21406,N_13291,N_13602);
and U21407 (N_21407,N_16699,N_15886);
nand U21408 (N_21408,N_13798,N_18061);
nand U21409 (N_21409,N_14026,N_16143);
nand U21410 (N_21410,N_18740,N_18077);
or U21411 (N_21411,N_12362,N_17791);
or U21412 (N_21412,N_19027,N_16722);
or U21413 (N_21413,N_11206,N_19281);
xor U21414 (N_21414,N_14728,N_13117);
or U21415 (N_21415,N_16803,N_17841);
and U21416 (N_21416,N_10949,N_19626);
and U21417 (N_21417,N_11148,N_15104);
and U21418 (N_21418,N_16696,N_15423);
nor U21419 (N_21419,N_18669,N_16975);
or U21420 (N_21420,N_10318,N_15117);
nor U21421 (N_21421,N_11569,N_17458);
nand U21422 (N_21422,N_12326,N_11028);
nor U21423 (N_21423,N_16678,N_12521);
and U21424 (N_21424,N_12895,N_18381);
nand U21425 (N_21425,N_10727,N_11733);
nand U21426 (N_21426,N_15461,N_15691);
or U21427 (N_21427,N_18568,N_16135);
xor U21428 (N_21428,N_14406,N_18883);
xor U21429 (N_21429,N_14203,N_13084);
nand U21430 (N_21430,N_16761,N_14191);
nand U21431 (N_21431,N_19470,N_10449);
or U21432 (N_21432,N_17774,N_17559);
nor U21433 (N_21433,N_10723,N_18092);
or U21434 (N_21434,N_13778,N_15420);
or U21435 (N_21435,N_19354,N_10371);
nor U21436 (N_21436,N_18632,N_10274);
nand U21437 (N_21437,N_15441,N_17647);
nand U21438 (N_21438,N_11758,N_19434);
nor U21439 (N_21439,N_17856,N_14388);
nor U21440 (N_21440,N_11557,N_13080);
xnor U21441 (N_21441,N_16542,N_12187);
xnor U21442 (N_21442,N_18008,N_19654);
and U21443 (N_21443,N_18647,N_12732);
and U21444 (N_21444,N_18523,N_12168);
xnor U21445 (N_21445,N_14804,N_15122);
or U21446 (N_21446,N_14063,N_17418);
nor U21447 (N_21447,N_10040,N_12320);
or U21448 (N_21448,N_10250,N_14119);
nand U21449 (N_21449,N_11194,N_10370);
nand U21450 (N_21450,N_18511,N_10775);
and U21451 (N_21451,N_15657,N_15406);
xnor U21452 (N_21452,N_11560,N_14687);
and U21453 (N_21453,N_16369,N_16733);
and U21454 (N_21454,N_15817,N_17476);
nand U21455 (N_21455,N_13673,N_14678);
and U21456 (N_21456,N_16128,N_11903);
or U21457 (N_21457,N_17677,N_17918);
nor U21458 (N_21458,N_11800,N_19468);
nor U21459 (N_21459,N_19901,N_14551);
nor U21460 (N_21460,N_12989,N_19436);
nand U21461 (N_21461,N_14234,N_13260);
nor U21462 (N_21462,N_19752,N_11548);
and U21463 (N_21463,N_17302,N_16829);
or U21464 (N_21464,N_18099,N_10455);
or U21465 (N_21465,N_19067,N_15642);
nor U21466 (N_21466,N_18130,N_10391);
nor U21467 (N_21467,N_11794,N_19524);
or U21468 (N_21468,N_13528,N_17883);
nor U21469 (N_21469,N_11020,N_17835);
and U21470 (N_21470,N_16300,N_12274);
or U21471 (N_21471,N_10788,N_16484);
or U21472 (N_21472,N_17084,N_10167);
and U21473 (N_21473,N_18671,N_13680);
or U21474 (N_21474,N_12195,N_15507);
nand U21475 (N_21475,N_12218,N_13866);
or U21476 (N_21476,N_18751,N_19484);
or U21477 (N_21477,N_14093,N_15224);
or U21478 (N_21478,N_10053,N_13848);
xor U21479 (N_21479,N_13262,N_18825);
and U21480 (N_21480,N_15499,N_13367);
or U21481 (N_21481,N_16120,N_15092);
and U21482 (N_21482,N_10932,N_19334);
or U21483 (N_21483,N_14811,N_10416);
or U21484 (N_21484,N_18688,N_17284);
or U21485 (N_21485,N_17018,N_16464);
or U21486 (N_21486,N_16784,N_16940);
and U21487 (N_21487,N_15108,N_13822);
nand U21488 (N_21488,N_13936,N_19984);
nand U21489 (N_21489,N_16867,N_18385);
xor U21490 (N_21490,N_18168,N_14897);
nand U21491 (N_21491,N_17462,N_17630);
nand U21492 (N_21492,N_16218,N_11358);
nand U21493 (N_21493,N_17611,N_16042);
or U21494 (N_21494,N_13092,N_18724);
and U21495 (N_21495,N_18959,N_18318);
nor U21496 (N_21496,N_11680,N_15816);
or U21497 (N_21497,N_17493,N_18721);
and U21498 (N_21498,N_13110,N_19785);
or U21499 (N_21499,N_17683,N_10066);
and U21500 (N_21500,N_19662,N_12357);
and U21501 (N_21501,N_19420,N_19219);
nand U21502 (N_21502,N_11585,N_11315);
and U21503 (N_21503,N_11558,N_19776);
or U21504 (N_21504,N_19118,N_13385);
nand U21505 (N_21505,N_13187,N_15781);
and U21506 (N_21506,N_12100,N_11312);
or U21507 (N_21507,N_16235,N_18657);
nor U21508 (N_21508,N_10096,N_18658);
or U21509 (N_21509,N_16652,N_19911);
and U21510 (N_21510,N_11485,N_17558);
xnor U21511 (N_21511,N_13565,N_12094);
nand U21512 (N_21512,N_19145,N_12184);
and U21513 (N_21513,N_16886,N_13837);
and U21514 (N_21514,N_13884,N_16953);
nand U21515 (N_21515,N_16581,N_12816);
or U21516 (N_21516,N_12629,N_12652);
xnor U21517 (N_21517,N_16717,N_12906);
nand U21518 (N_21518,N_15715,N_13271);
nor U21519 (N_21519,N_17607,N_13365);
or U21520 (N_21520,N_11995,N_13382);
nand U21521 (N_21521,N_19741,N_15161);
and U21522 (N_21522,N_11432,N_15516);
nand U21523 (N_21523,N_15353,N_12807);
or U21524 (N_21524,N_17478,N_11164);
or U21525 (N_21525,N_17129,N_14970);
nor U21526 (N_21526,N_15801,N_11922);
nor U21527 (N_21527,N_11001,N_12758);
nand U21528 (N_21528,N_15809,N_16672);
or U21529 (N_21529,N_13445,N_11331);
or U21530 (N_21530,N_14832,N_16506);
xnor U21531 (N_21531,N_19815,N_19680);
nor U21532 (N_21532,N_18354,N_17182);
nor U21533 (N_21533,N_11596,N_12253);
xor U21534 (N_21534,N_14490,N_17532);
nor U21535 (N_21535,N_10136,N_18135);
and U21536 (N_21536,N_17688,N_12162);
or U21537 (N_21537,N_10709,N_11969);
nor U21538 (N_21538,N_18782,N_12109);
and U21539 (N_21539,N_18187,N_18946);
nand U21540 (N_21540,N_16855,N_16758);
or U21541 (N_21541,N_19324,N_13391);
or U21542 (N_21542,N_19641,N_14843);
nand U21543 (N_21543,N_18291,N_17645);
nand U21544 (N_21544,N_18222,N_12645);
or U21545 (N_21545,N_15512,N_14507);
nand U21546 (N_21546,N_19005,N_14680);
nand U21547 (N_21547,N_17708,N_16885);
nor U21548 (N_21548,N_11349,N_14840);
or U21549 (N_21549,N_16138,N_19665);
or U21550 (N_21550,N_13285,N_17331);
nor U21551 (N_21551,N_17021,N_18190);
nor U21552 (N_21552,N_10468,N_11620);
or U21553 (N_21553,N_18307,N_17100);
xor U21554 (N_21554,N_11019,N_17252);
nand U21555 (N_21555,N_19475,N_17664);
and U21556 (N_21556,N_14084,N_17375);
nor U21557 (N_21557,N_13295,N_13467);
and U21558 (N_21558,N_15014,N_14333);
and U21559 (N_21559,N_17291,N_15260);
or U21560 (N_21560,N_14777,N_17877);
or U21561 (N_21561,N_16107,N_17702);
or U21562 (N_21562,N_19265,N_14379);
or U21563 (N_21563,N_14365,N_12017);
and U21564 (N_21564,N_14803,N_13479);
nand U21565 (N_21565,N_17272,N_19105);
or U21566 (N_21566,N_19916,N_14164);
and U21567 (N_21567,N_10531,N_13186);
nor U21568 (N_21568,N_10340,N_12191);
nor U21569 (N_21569,N_12110,N_10091);
nor U21570 (N_21570,N_19315,N_13539);
xor U21571 (N_21571,N_15299,N_16691);
and U21572 (N_21572,N_15812,N_16544);
or U21573 (N_21573,N_17951,N_14503);
nand U21574 (N_21574,N_19488,N_12234);
nand U21575 (N_21575,N_16610,N_14417);
or U21576 (N_21576,N_14465,N_16467);
and U21577 (N_21577,N_10535,N_17718);
and U21578 (N_21578,N_17712,N_15640);
nor U21579 (N_21579,N_16526,N_12079);
and U21580 (N_21580,N_14363,N_17557);
and U21581 (N_21581,N_15603,N_19250);
and U21582 (N_21582,N_18344,N_17325);
xor U21583 (N_21583,N_19622,N_15137);
nor U21584 (N_21584,N_18460,N_12733);
nor U21585 (N_21585,N_18771,N_10511);
xor U21586 (N_21586,N_13079,N_12034);
nand U21587 (N_21587,N_17401,N_16968);
nor U21588 (N_21588,N_12593,N_16452);
nand U21589 (N_21589,N_10259,N_19142);
nor U21590 (N_21590,N_19875,N_12612);
nor U21591 (N_21591,N_19486,N_10847);
xnor U21592 (N_21592,N_14681,N_12020);
xor U21593 (N_21593,N_16569,N_18358);
nor U21594 (N_21594,N_15395,N_16450);
xor U21595 (N_21595,N_12892,N_14261);
or U21596 (N_21596,N_13413,N_18148);
nor U21597 (N_21597,N_13240,N_14648);
and U21598 (N_21598,N_13218,N_12858);
and U21599 (N_21599,N_11414,N_12464);
nand U21600 (N_21600,N_18518,N_15337);
or U21601 (N_21601,N_16295,N_16646);
nand U21602 (N_21602,N_15889,N_14603);
nand U21603 (N_21603,N_16185,N_15328);
xor U21604 (N_21604,N_12685,N_14034);
and U21605 (N_21605,N_11935,N_18216);
and U21606 (N_21606,N_18838,N_17871);
or U21607 (N_21607,N_18287,N_16900);
nand U21608 (N_21608,N_14353,N_15050);
nand U21609 (N_21609,N_12584,N_13416);
xor U21610 (N_21610,N_18714,N_10867);
nand U21611 (N_21611,N_10762,N_12105);
nor U21612 (N_21612,N_15021,N_14271);
nor U21613 (N_21613,N_18286,N_19945);
or U21614 (N_21614,N_10215,N_18970);
or U21615 (N_21615,N_12658,N_16612);
xor U21616 (N_21616,N_13185,N_13028);
and U21617 (N_21617,N_13307,N_18010);
nand U21618 (N_21618,N_19210,N_14574);
nand U21619 (N_21619,N_13745,N_12535);
nand U21620 (N_21620,N_13442,N_11054);
and U21621 (N_21621,N_12126,N_12066);
nand U21622 (N_21622,N_15078,N_13708);
nand U21623 (N_21623,N_15449,N_10651);
or U21624 (N_21624,N_17354,N_13107);
or U21625 (N_21625,N_12520,N_15532);
nor U21626 (N_21626,N_15324,N_13662);
nor U21627 (N_21627,N_13173,N_16593);
nand U21628 (N_21628,N_13480,N_18436);
nor U21629 (N_21629,N_16401,N_17232);
nand U21630 (N_21630,N_16942,N_19632);
or U21631 (N_21631,N_18201,N_11167);
nor U21632 (N_21632,N_13188,N_12920);
or U21633 (N_21633,N_18205,N_17685);
or U21634 (N_21634,N_15218,N_10846);
and U21635 (N_21635,N_19181,N_15857);
nand U21636 (N_21636,N_13193,N_16337);
and U21637 (N_21637,N_10072,N_17456);
or U21638 (N_21638,N_18634,N_10364);
nand U21639 (N_21639,N_11694,N_17722);
and U21640 (N_21640,N_10743,N_15628);
xor U21641 (N_21641,N_14833,N_16957);
and U21642 (N_21642,N_11403,N_14725);
and U21643 (N_21643,N_12205,N_10275);
nand U21644 (N_21644,N_11874,N_19199);
and U21645 (N_21645,N_12284,N_14050);
and U21646 (N_21646,N_12651,N_15327);
and U21647 (N_21647,N_13855,N_16603);
and U21648 (N_21648,N_16291,N_12299);
or U21649 (N_21649,N_10670,N_16624);
and U21650 (N_21650,N_13762,N_13808);
nor U21651 (N_21651,N_15240,N_19755);
or U21652 (N_21652,N_15705,N_10557);
nor U21653 (N_21653,N_15675,N_19078);
and U21654 (N_21654,N_16237,N_13716);
or U21655 (N_21655,N_18818,N_12557);
nand U21656 (N_21656,N_15135,N_15480);
and U21657 (N_21657,N_12272,N_17443);
nor U21658 (N_21658,N_14920,N_18467);
xnor U21659 (N_21659,N_11798,N_19305);
nor U21660 (N_21660,N_18448,N_17503);
and U21661 (N_21661,N_17276,N_16816);
and U21662 (N_21662,N_13626,N_10396);
or U21663 (N_21663,N_18044,N_10489);
nand U21664 (N_21664,N_12472,N_15938);
nand U21665 (N_21665,N_14346,N_12930);
and U21666 (N_21666,N_18255,N_16269);
and U21667 (N_21667,N_17190,N_17244);
and U21668 (N_21668,N_16289,N_17531);
or U21669 (N_21669,N_19992,N_14424);
and U21670 (N_21670,N_13825,N_17928);
and U21671 (N_21671,N_15256,N_14835);
and U21672 (N_21672,N_13434,N_15733);
nand U21673 (N_21673,N_16525,N_18493);
or U21674 (N_21674,N_14403,N_13286);
nor U21675 (N_21675,N_14549,N_11243);
and U21676 (N_21676,N_16777,N_12502);
nor U21677 (N_21677,N_16964,N_17053);
or U21678 (N_21678,N_10807,N_15247);
nand U21679 (N_21679,N_14508,N_16971);
or U21680 (N_21680,N_15578,N_16756);
nor U21681 (N_21681,N_12933,N_17993);
and U21682 (N_21682,N_13145,N_10884);
xnor U21683 (N_21683,N_17178,N_15585);
or U21684 (N_21684,N_12157,N_13591);
and U21685 (N_21685,N_12704,N_18513);
nand U21686 (N_21686,N_13349,N_10776);
nor U21687 (N_21687,N_16790,N_13874);
nand U21688 (N_21688,N_19380,N_19472);
nor U21689 (N_21689,N_10433,N_13027);
or U21690 (N_21690,N_16767,N_15295);
nor U21691 (N_21691,N_12916,N_15551);
or U21692 (N_21692,N_18125,N_14094);
or U21693 (N_21693,N_17682,N_14605);
and U21694 (N_21694,N_19197,N_11398);
or U21695 (N_21695,N_15998,N_14221);
or U21696 (N_21696,N_12348,N_11906);
or U21697 (N_21697,N_18567,N_17516);
and U21698 (N_21698,N_18271,N_16567);
or U21699 (N_21699,N_14180,N_13115);
nor U21700 (N_21700,N_15651,N_16212);
xor U21701 (N_21701,N_14608,N_11275);
nor U21702 (N_21702,N_17567,N_12957);
nand U21703 (N_21703,N_18885,N_13761);
nand U21704 (N_21704,N_13414,N_12690);
nor U21705 (N_21705,N_18246,N_14894);
nand U21706 (N_21706,N_12694,N_13902);
or U21707 (N_21707,N_14135,N_15455);
nand U21708 (N_21708,N_12689,N_10472);
nor U21709 (N_21709,N_13867,N_17235);
nand U21710 (N_21710,N_18553,N_19550);
or U21711 (N_21711,N_19196,N_17986);
xnor U21712 (N_21712,N_14610,N_11139);
nand U21713 (N_21713,N_12398,N_11960);
nand U21714 (N_21714,N_11003,N_17269);
or U21715 (N_21715,N_10346,N_18111);
or U21716 (N_21716,N_10565,N_15638);
or U21717 (N_21717,N_13806,N_11368);
nand U21718 (N_21718,N_19743,N_12600);
xnor U21719 (N_21719,N_17536,N_11915);
or U21720 (N_21720,N_18738,N_12043);
nand U21721 (N_21721,N_18174,N_13675);
or U21722 (N_21722,N_18036,N_13502);
nand U21723 (N_21723,N_10475,N_19186);
nor U21724 (N_21724,N_10206,N_18292);
or U21725 (N_21725,N_16119,N_19775);
or U21726 (N_21726,N_15426,N_16959);
or U21727 (N_21727,N_10238,N_13978);
nand U21728 (N_21728,N_10197,N_18098);
or U21729 (N_21729,N_11536,N_11375);
or U21730 (N_21730,N_12174,N_19744);
or U21731 (N_21731,N_14127,N_10458);
nand U21732 (N_21732,N_14892,N_18425);
nor U21733 (N_21733,N_15676,N_15615);
or U21734 (N_21734,N_16914,N_14055);
and U21735 (N_21735,N_17961,N_10603);
and U21736 (N_21736,N_19188,N_14670);
nor U21737 (N_21737,N_16367,N_16485);
and U21738 (N_21738,N_15969,N_12678);
nor U21739 (N_21739,N_12705,N_15300);
nand U21740 (N_21740,N_19370,N_13620);
and U21741 (N_21741,N_18800,N_19537);
and U21742 (N_21742,N_19826,N_19042);
nand U21743 (N_21743,N_19192,N_14039);
nor U21744 (N_21744,N_10442,N_15957);
and U21745 (N_21745,N_15648,N_14534);
nor U21746 (N_21746,N_19808,N_18323);
or U21747 (N_21747,N_13652,N_15134);
nand U21748 (N_21748,N_18261,N_18831);
or U21749 (N_21749,N_11933,N_15167);
or U21750 (N_21750,N_18038,N_14748);
nor U21751 (N_21751,N_13474,N_13301);
nor U21752 (N_21752,N_10196,N_17505);
and U21753 (N_21753,N_11791,N_15318);
and U21754 (N_21754,N_19444,N_17322);
nand U21755 (N_21755,N_10717,N_12682);
nand U21756 (N_21756,N_18017,N_13016);
nor U21757 (N_21757,N_19791,N_17150);
or U21758 (N_21758,N_18089,N_11269);
or U21759 (N_21759,N_10998,N_19411);
and U21760 (N_21760,N_17154,N_12204);
nor U21761 (N_21761,N_18922,N_15557);
nor U21762 (N_21762,N_17552,N_12016);
nand U21763 (N_21763,N_19658,N_18860);
and U21764 (N_21764,N_19168,N_12723);
nand U21765 (N_21765,N_10138,N_19134);
nand U21766 (N_21766,N_17092,N_11675);
or U21767 (N_21767,N_15375,N_15404);
nor U21768 (N_21768,N_14773,N_16019);
and U21769 (N_21769,N_12047,N_18004);
nor U21770 (N_21770,N_12497,N_13860);
nand U21771 (N_21771,N_13410,N_18759);
nand U21772 (N_21772,N_19207,N_16505);
nor U21773 (N_21773,N_10029,N_12113);
and U21774 (N_21774,N_15123,N_12366);
or U21775 (N_21775,N_15868,N_10744);
nand U21776 (N_21776,N_14567,N_11886);
and U21777 (N_21777,N_19072,N_16944);
nand U21778 (N_21778,N_13674,N_17577);
or U21779 (N_21779,N_15555,N_15863);
nor U21780 (N_21780,N_15332,N_15520);
nor U21781 (N_21781,N_13522,N_16444);
xor U21782 (N_21782,N_16584,N_10719);
nand U21783 (N_21783,N_12442,N_12292);
or U21784 (N_21784,N_10814,N_12229);
xor U21785 (N_21785,N_13373,N_17967);
nor U21786 (N_21786,N_15798,N_16861);
and U21787 (N_21787,N_18478,N_13923);
or U21788 (N_21788,N_18305,N_17734);
nand U21789 (N_21789,N_17311,N_12211);
or U21790 (N_21790,N_15203,N_12271);
nor U21791 (N_21791,N_10123,N_11489);
or U21792 (N_21792,N_15743,N_12024);
nand U21793 (N_21793,N_16129,N_10567);
or U21794 (N_21794,N_10999,N_17185);
nor U21795 (N_21795,N_16220,N_14300);
nand U21796 (N_21796,N_10255,N_15940);
nand U21797 (N_21797,N_19014,N_14847);
xnor U21798 (N_21798,N_10948,N_14623);
nor U21799 (N_21799,N_18439,N_13873);
nor U21800 (N_21800,N_15590,N_11572);
and U21801 (N_21801,N_11457,N_17915);
nand U21802 (N_21802,N_12036,N_14787);
nor U21803 (N_21803,N_16549,N_16841);
nor U21804 (N_21804,N_15631,N_16208);
nor U21805 (N_21805,N_16091,N_17521);
nand U21806 (N_21806,N_14126,N_10599);
nor U21807 (N_21807,N_12735,N_13705);
nand U21808 (N_21808,N_18002,N_12026);
and U21809 (N_21809,N_13520,N_13358);
and U21810 (N_21810,N_14985,N_13856);
nand U21811 (N_21811,N_18349,N_16747);
nor U21812 (N_21812,N_13114,N_12021);
nand U21813 (N_21813,N_14577,N_18319);
nand U21814 (N_21814,N_19043,N_18604);
or U21815 (N_21815,N_14659,N_13074);
and U21816 (N_21816,N_18560,N_15000);
nand U21817 (N_21817,N_16514,N_10501);
xor U21818 (N_21818,N_13169,N_19713);
nor U21819 (N_21819,N_10276,N_15060);
nand U21820 (N_21820,N_13310,N_15463);
xor U21821 (N_21821,N_11949,N_17349);
nand U21822 (N_21822,N_13770,N_11137);
nand U21823 (N_21823,N_16932,N_13945);
nor U21824 (N_21824,N_19500,N_15913);
nor U21825 (N_21825,N_12077,N_15248);
nor U21826 (N_21826,N_11195,N_11718);
nor U21827 (N_21827,N_13587,N_18360);
nor U21828 (N_21828,N_14699,N_18244);
nor U21829 (N_21829,N_17527,N_10860);
nand U21830 (N_21830,N_15236,N_19670);
and U21831 (N_21831,N_14602,N_11090);
and U21832 (N_21832,N_14930,N_11397);
or U21833 (N_21833,N_18131,N_16537);
or U21834 (N_21834,N_15614,N_14857);
nand U21835 (N_21835,N_16547,N_17938);
nand U21836 (N_21836,N_11246,N_15984);
and U21837 (N_21837,N_15700,N_14325);
nor U21838 (N_21838,N_15271,N_13628);
nand U21839 (N_21839,N_15384,N_15935);
nor U21840 (N_21840,N_10242,N_14110);
nor U21841 (N_21841,N_15081,N_19487);
and U21842 (N_21842,N_18074,N_13842);
or U21843 (N_21843,N_19736,N_16310);
nand U21844 (N_21844,N_17893,N_10479);
and U21845 (N_21845,N_17010,N_16177);
xnor U21846 (N_21846,N_11615,N_15326);
nor U21847 (N_21847,N_19352,N_19935);
nand U21848 (N_21848,N_12343,N_14051);
or U21849 (N_21849,N_15586,N_19331);
nand U21850 (N_21850,N_11204,N_15922);
nand U21851 (N_21851,N_18069,N_19498);
or U21852 (N_21852,N_10526,N_19077);
or U21853 (N_21853,N_16799,N_15727);
or U21854 (N_21854,N_17976,N_14633);
nand U21855 (N_21855,N_19549,N_14941);
nor U21856 (N_21856,N_18844,N_19616);
nand U21857 (N_21857,N_13567,N_14667);
or U21858 (N_21858,N_14104,N_11248);
nand U21859 (N_21859,N_16781,N_11441);
nand U21860 (N_21860,N_17624,N_14831);
nand U21861 (N_21861,N_11787,N_15950);
and U21862 (N_21862,N_16728,N_19963);
or U21863 (N_21863,N_14562,N_15917);
or U21864 (N_21864,N_17222,N_14542);
and U21865 (N_21865,N_19298,N_13354);
nor U21866 (N_21866,N_17355,N_17985);
xnor U21867 (N_21867,N_15088,N_16503);
xor U21868 (N_21868,N_12981,N_11304);
and U21869 (N_21869,N_15987,N_11747);
xnor U21870 (N_21870,N_10560,N_15155);
nand U21871 (N_21871,N_18662,N_13042);
nor U21872 (N_21872,N_14816,N_19592);
or U21873 (N_21873,N_19859,N_11545);
and U21874 (N_21874,N_13459,N_18975);
nand U21875 (N_21875,N_12923,N_14979);
nand U21876 (N_21876,N_14958,N_11844);
nand U21877 (N_21877,N_12091,N_14161);
nor U21878 (N_21878,N_13100,N_10374);
and U21879 (N_21879,N_19760,N_10080);
and U21880 (N_21880,N_13655,N_13696);
or U21881 (N_21881,N_15618,N_16820);
nor U21882 (N_21882,N_13713,N_18608);
nand U21883 (N_21883,N_11405,N_17575);
and U21884 (N_21884,N_19827,N_11662);
xor U21885 (N_21885,N_16941,N_15368);
nand U21886 (N_21886,N_11792,N_16903);
or U21887 (N_21887,N_18071,N_17378);
nor U21888 (N_21888,N_15311,N_19328);
nor U21889 (N_21889,N_14276,N_16219);
or U21890 (N_21890,N_10048,N_14411);
and U21891 (N_21891,N_14999,N_14367);
nor U21892 (N_21892,N_13881,N_11717);
or U21893 (N_21893,N_10698,N_10247);
nor U21894 (N_21894,N_10349,N_14994);
or U21895 (N_21895,N_19009,N_15254);
xor U21896 (N_21896,N_19853,N_18943);
xnor U21897 (N_21897,N_15699,N_18925);
or U21898 (N_21898,N_13421,N_16360);
nor U21899 (N_21899,N_11762,N_16524);
and U21900 (N_21900,N_16418,N_13088);
nor U21901 (N_21901,N_12909,N_16349);
nand U21902 (N_21902,N_18799,N_13824);
nand U21903 (N_21903,N_19742,N_18210);
xnor U21904 (N_21904,N_18973,N_17510);
nand U21905 (N_21905,N_14253,N_14470);
or U21906 (N_21906,N_17638,N_10777);
nand U21907 (N_21907,N_15807,N_15239);
or U21908 (N_21908,N_13568,N_11121);
or U21909 (N_21909,N_17317,N_13101);
and U21910 (N_21910,N_12792,N_16579);
or U21911 (N_21911,N_10604,N_15622);
nor U21912 (N_21912,N_14830,N_18775);
xor U21913 (N_21913,N_16179,N_10622);
xnor U21914 (N_21914,N_10737,N_12937);
or U21915 (N_21915,N_18482,N_17944);
nor U21916 (N_21916,N_14972,N_17086);
or U21917 (N_21917,N_13249,N_10946);
and U21918 (N_21918,N_17413,N_10803);
and U21919 (N_21919,N_14179,N_11769);
nor U21920 (N_21920,N_17467,N_11824);
nor U21921 (N_21921,N_15170,N_11779);
or U21922 (N_21922,N_19638,N_12448);
nand U21923 (N_21923,N_19897,N_14926);
nor U21924 (N_21924,N_18882,N_17080);
and U21925 (N_21925,N_14354,N_16044);
and U21926 (N_21926,N_10987,N_10575);
or U21927 (N_21927,N_10797,N_12707);
nand U21928 (N_21928,N_13180,N_12887);
nor U21929 (N_21929,N_15612,N_11774);
or U21930 (N_21930,N_16382,N_12994);
or U21931 (N_21931,N_18909,N_15710);
and U21932 (N_21932,N_19184,N_11425);
nand U21933 (N_21933,N_19928,N_18635);
nor U21934 (N_21934,N_18030,N_14143);
xnor U21935 (N_21935,N_10401,N_12709);
or U21936 (N_21936,N_19114,N_13429);
nand U21937 (N_21937,N_11784,N_15763);
nor U21938 (N_21938,N_12290,N_10300);
or U21939 (N_21939,N_16882,N_19392);
or U21940 (N_21940,N_17580,N_14969);
nand U21941 (N_21941,N_15223,N_18073);
or U21942 (N_21942,N_11064,N_10952);
nor U21943 (N_21943,N_19171,N_13545);
nand U21944 (N_21944,N_19445,N_19125);
nor U21945 (N_21945,N_12314,N_13204);
nor U21946 (N_21946,N_13847,N_14931);
or U21947 (N_21947,N_19073,N_17955);
and U21948 (N_21948,N_18876,N_19531);
xnor U21949 (N_21949,N_17689,N_19150);
nor U21950 (N_21950,N_17422,N_19391);
or U21951 (N_21951,N_17681,N_17197);
xnor U21952 (N_21952,N_12988,N_10726);
nor U21953 (N_21953,N_19026,N_10574);
or U21954 (N_21954,N_19806,N_14240);
nor U21955 (N_21955,N_17844,N_12401);
or U21956 (N_21956,N_17037,N_12492);
nand U21957 (N_21957,N_14636,N_16368);
nor U21958 (N_21958,N_12729,N_16521);
nor U21959 (N_21959,N_11142,N_18600);
nor U21960 (N_21960,N_10782,N_13999);
nand U21961 (N_21961,N_10945,N_15434);
nand U21962 (N_21962,N_12954,N_16341);
xnor U21963 (N_21963,N_19408,N_18282);
and U21964 (N_21964,N_10514,N_14401);
nor U21965 (N_21965,N_17771,N_12801);
and U21966 (N_21966,N_10534,N_11514);
or U21967 (N_21967,N_15593,N_13093);
xnor U21968 (N_21968,N_14255,N_16470);
nand U21969 (N_21969,N_18859,N_11750);
and U21970 (N_21970,N_17411,N_19421);
nor U21971 (N_21971,N_10135,N_14455);
and U21972 (N_21972,N_14909,N_11392);
and U21973 (N_21973,N_14921,N_16010);
nand U21974 (N_21974,N_13843,N_17862);
or U21975 (N_21975,N_15208,N_15190);
and U21976 (N_21976,N_16713,N_11498);
or U21977 (N_21977,N_18403,N_12042);
nor U21978 (N_21978,N_17963,N_10906);
or U21979 (N_21979,N_11635,N_14786);
xor U21980 (N_21980,N_19364,N_10715);
and U21981 (N_21981,N_10731,N_12007);
xor U21982 (N_21982,N_19964,N_16743);
nor U21983 (N_21983,N_18312,N_10595);
and U21984 (N_21984,N_12512,N_13644);
nand U21985 (N_21985,N_16922,N_11554);
nor U21986 (N_21986,N_13871,N_17658);
or U21987 (N_21987,N_16149,N_18455);
nand U21988 (N_21988,N_16421,N_11260);
and U21989 (N_21989,N_19724,N_11859);
nand U21990 (N_21990,N_14957,N_11239);
nor U21991 (N_21991,N_11757,N_11528);
nor U21992 (N_21992,N_13272,N_10284);
and U21993 (N_21993,N_17863,N_15785);
xnor U21994 (N_21994,N_10506,N_17737);
xnor U21995 (N_21995,N_17023,N_16438);
nand U21996 (N_21996,N_13455,N_17698);
and U21997 (N_21997,N_13341,N_10733);
nand U21998 (N_21998,N_14369,N_12625);
xnor U21999 (N_21999,N_12561,N_10216);
nor U22000 (N_22000,N_18522,N_15955);
or U22001 (N_22001,N_16307,N_19182);
and U22002 (N_22002,N_16502,N_19050);
xnor U22003 (N_22003,N_14976,N_10461);
and U22004 (N_22004,N_14088,N_10209);
nor U22005 (N_22005,N_18646,N_17888);
nand U22006 (N_22006,N_15698,N_13801);
xor U22007 (N_22007,N_11928,N_15717);
and U22008 (N_22008,N_18171,N_15055);
nand U22009 (N_22009,N_13694,N_11009);
and U22010 (N_22010,N_11138,N_16592);
nor U22011 (N_22011,N_14850,N_14669);
nand U22012 (N_22012,N_11463,N_19051);
nor U22013 (N_22013,N_19960,N_15519);
or U22014 (N_22014,N_14232,N_13910);
or U22015 (N_22015,N_17299,N_18599);
xnor U22016 (N_22016,N_16988,N_12005);
nand U22017 (N_22017,N_13630,N_13803);
nand U22018 (N_22018,N_13641,N_15494);
or U22019 (N_22019,N_14951,N_11257);
or U22020 (N_22020,N_13176,N_12635);
and U22021 (N_22021,N_10311,N_17819);
and U22022 (N_22022,N_19262,N_17874);
xor U22023 (N_22023,N_18153,N_12273);
or U22024 (N_22024,N_10353,N_13627);
and U22025 (N_22025,N_10521,N_12822);
nand U22026 (N_22026,N_13579,N_11190);
and U22027 (N_22027,N_10970,N_13065);
nor U22028 (N_22028,N_14893,N_15490);
or U22029 (N_22029,N_15136,N_11372);
or U22030 (N_22030,N_18999,N_12841);
xor U22031 (N_22031,N_19812,N_10498);
or U22032 (N_22032,N_17742,N_18498);
or U22033 (N_22033,N_13768,N_11404);
or U22034 (N_22034,N_14550,N_18886);
or U22035 (N_22035,N_18578,N_13122);
and U22036 (N_22036,N_16283,N_18916);
nand U22037 (N_22037,N_15629,N_19507);
or U22038 (N_22038,N_11109,N_13594);
and U22039 (N_22039,N_14784,N_10120);
nand U22040 (N_22040,N_12434,N_19881);
xor U22041 (N_22041,N_19649,N_12519);
or U22042 (N_22042,N_17104,N_10347);
and U22043 (N_22043,N_13205,N_16522);
and U22044 (N_22044,N_15893,N_19764);
nor U22045 (N_22045,N_13181,N_10189);
and U22046 (N_22046,N_13505,N_19612);
or U22047 (N_22047,N_16854,N_14430);
nand U22048 (N_22048,N_15471,N_14531);
nor U22049 (N_22049,N_10257,N_12399);
and U22050 (N_22050,N_10765,N_13077);
nand U22051 (N_22051,N_11380,N_18733);
nor U22052 (N_22052,N_13557,N_11413);
or U22053 (N_22053,N_12626,N_11214);
and U22054 (N_22054,N_11857,N_12966);
nand U22055 (N_22055,N_19718,N_18142);
nor U22056 (N_22056,N_15606,N_17224);
and U22057 (N_22057,N_13006,N_10793);
xor U22058 (N_22058,N_16071,N_17345);
nand U22059 (N_22059,N_11534,N_16005);
nand U22060 (N_22060,N_19998,N_18697);
nor U22061 (N_22061,N_13814,N_14292);
or U22062 (N_22062,N_11803,N_14400);
and U22063 (N_22063,N_19754,N_12387);
and U22064 (N_22064,N_10463,N_10504);
nand U22065 (N_22065,N_10178,N_13997);
nor U22066 (N_22066,N_14553,N_17239);
xor U22067 (N_22067,N_19535,N_15405);
or U22068 (N_22068,N_16108,N_12539);
nor U22069 (N_22069,N_16831,N_13536);
or U22070 (N_22070,N_19686,N_11970);
nor U22071 (N_22071,N_14140,N_11250);
and U22072 (N_22072,N_18609,N_16186);
or U22073 (N_22073,N_13859,N_11561);
nand U22074 (N_22074,N_13072,N_19479);
and U22075 (N_22075,N_14052,N_18143);
or U22076 (N_22076,N_16632,N_17351);
xnor U22077 (N_22077,N_19069,N_14964);
and U22078 (N_22078,N_10663,N_15732);
xnor U22079 (N_22079,N_15386,N_10757);
xnor U22080 (N_22080,N_10287,N_10204);
nor U22081 (N_22081,N_18583,N_12267);
nor U22082 (N_22082,N_19929,N_11947);
and U22083 (N_22083,N_10689,N_16725);
and U22084 (N_22084,N_16402,N_15298);
or U22085 (N_22085,N_19923,N_15748);
nand U22086 (N_22086,N_18189,N_19574);
xnor U22087 (N_22087,N_13646,N_18491);
nand U22088 (N_22088,N_17554,N_13913);
nand U22089 (N_22089,N_14082,N_14658);
or U22090 (N_22090,N_16272,N_12934);
or U22091 (N_22091,N_15914,N_13125);
nand U22092 (N_22092,N_11149,N_16339);
and U22093 (N_22093,N_19871,N_18311);
xnor U22094 (N_22094,N_12534,N_16045);
nor U22095 (N_22095,N_17911,N_13155);
nor U22096 (N_22096,N_16700,N_11942);
nand U22097 (N_22097,N_10055,N_13835);
nand U22098 (N_22098,N_19688,N_12276);
or U22099 (N_22099,N_10704,N_16719);
or U22100 (N_22100,N_11977,N_17996);
and U22101 (N_22101,N_18233,N_10607);
or U22102 (N_22102,N_14851,N_10165);
nor U22103 (N_22103,N_10728,N_18760);
nor U22104 (N_22104,N_16600,N_12601);
or U22105 (N_22105,N_12700,N_13091);
nor U22106 (N_22106,N_19279,N_14998);
nor U22107 (N_22107,N_13868,N_15827);
and U22108 (N_22108,N_16242,N_17512);
and U22109 (N_22109,N_18630,N_10540);
nand U22110 (N_22110,N_10386,N_15599);
xnor U22111 (N_22111,N_10692,N_12394);
nor U22112 (N_22112,N_12551,N_12929);
nor U22113 (N_22113,N_11773,N_11024);
or U22114 (N_22114,N_10761,N_13140);
and U22115 (N_22115,N_10556,N_11807);
and U22116 (N_22116,N_18791,N_14827);
xnor U22117 (N_22117,N_14869,N_17686);
nor U22118 (N_22118,N_15543,N_19878);
or U22119 (N_22119,N_11836,N_18327);
nand U22120 (N_22120,N_11510,N_13424);
nand U22121 (N_22121,N_11014,N_11385);
or U22122 (N_22122,N_14789,N_19938);
and U22123 (N_22123,N_11810,N_12696);
or U22124 (N_22124,N_11330,N_15591);
or U22125 (N_22125,N_10941,N_17402);
nand U22126 (N_22126,N_17788,N_16445);
or U22127 (N_22127,N_11333,N_10507);
nor U22128 (N_22128,N_18934,N_11651);
or U22129 (N_22129,N_12800,N_10665);
or U22130 (N_22130,N_15323,N_17408);
nor U22131 (N_22131,N_12011,N_17013);
or U22132 (N_22132,N_12494,N_19982);
or U22133 (N_22133,N_11193,N_17614);
or U22134 (N_22134,N_10129,N_12544);
nand U22135 (N_22135,N_11023,N_18353);
xor U22136 (N_22136,N_15481,N_12386);
nor U22137 (N_22137,N_18078,N_15127);
nor U22138 (N_22138,N_17966,N_11689);
or U22139 (N_22139,N_10243,N_11997);
and U22140 (N_22140,N_13355,N_18617);
and U22141 (N_22141,N_11198,N_18903);
nand U22142 (N_22142,N_16261,N_14194);
nor U22143 (N_22143,N_13047,N_11437);
and U22144 (N_22144,N_17250,N_16616);
nor U22145 (N_22145,N_12817,N_14855);
and U22146 (N_22146,N_13656,N_17631);
and U22147 (N_22147,N_14152,N_14536);
and U22148 (N_22148,N_19242,N_18463);
nor U22149 (N_22149,N_16439,N_10576);
nor U22150 (N_22150,N_17914,N_13029);
or U22151 (N_22151,N_16568,N_11991);
nor U22152 (N_22152,N_15085,N_16589);
and U22153 (N_22153,N_18673,N_15487);
nand U22154 (N_22154,N_12691,N_13926);
nor U22155 (N_22155,N_12287,N_15592);
and U22156 (N_22156,N_11551,N_12022);
xnor U22157 (N_22157,N_11162,N_16864);
nand U22158 (N_22158,N_18066,N_13531);
nor U22159 (N_22159,N_14100,N_11931);
or U22160 (N_22160,N_11737,N_16062);
or U22161 (N_22161,N_13612,N_11335);
or U22162 (N_22162,N_10973,N_11448);
and U22163 (N_22163,N_12872,N_19035);
and U22164 (N_22164,N_16640,N_14010);
nor U22165 (N_22165,N_12830,N_19748);
xor U22166 (N_22166,N_13275,N_12201);
nor U22167 (N_22167,N_11145,N_15571);
nor U22168 (N_22168,N_14734,N_16426);
or U22169 (N_22169,N_15402,N_15090);
nor U22170 (N_22170,N_13529,N_17678);
or U22171 (N_22171,N_18348,N_14456);
nor U22172 (N_22172,N_14884,N_14472);
and U22173 (N_22173,N_12529,N_18301);
nand U22174 (N_22174,N_11343,N_11707);
and U22175 (N_22175,N_12315,N_10829);
nor U22176 (N_22176,N_10363,N_12069);
nor U22177 (N_22177,N_17618,N_14580);
nor U22178 (N_22178,N_10802,N_14656);
nor U22179 (N_22179,N_17093,N_19146);
xor U22180 (N_22180,N_18299,N_10713);
nor U22181 (N_22181,N_15281,N_10895);
nor U22182 (N_22182,N_15838,N_19349);
nor U22183 (N_22183,N_19689,N_16682);
or U22184 (N_22184,N_19715,N_17522);
and U22185 (N_22185,N_12373,N_11272);
nor U22186 (N_22186,N_19357,N_12150);
nand U22187 (N_22187,N_10680,N_12863);
or U22188 (N_22188,N_13305,N_12322);
nor U22189 (N_22189,N_16239,N_17241);
or U22190 (N_22190,N_16027,N_12078);
or U22191 (N_22191,N_12038,N_16866);
nor U22192 (N_22192,N_12112,N_10905);
nand U22193 (N_22193,N_16171,N_16538);
and U22194 (N_22194,N_10341,N_12902);
xor U22195 (N_22195,N_15718,N_17514);
nand U22196 (N_22196,N_16160,N_15901);
or U22197 (N_22197,N_11378,N_12891);
nor U22198 (N_22198,N_12655,N_13011);
or U22199 (N_22199,N_13245,N_12662);
nand U22200 (N_22200,N_14270,N_18456);
or U22201 (N_22201,N_12432,N_12943);
xnor U22202 (N_22202,N_10004,N_14802);
nand U22203 (N_22203,N_15417,N_13095);
or U22204 (N_22204,N_18703,N_17039);
nand U22205 (N_22205,N_17649,N_16404);
xor U22206 (N_22206,N_16907,N_15407);
or U22207 (N_22207,N_15966,N_10035);
xnor U22208 (N_22208,N_18938,N_19532);
nand U22209 (N_22209,N_14492,N_10594);
nor U22210 (N_22210,N_19323,N_17755);
and U22211 (N_22211,N_17746,N_19294);
nand U22212 (N_22212,N_15215,N_13494);
xnor U22213 (N_22213,N_10938,N_19946);
nor U22214 (N_22214,N_13924,N_19131);
nand U22215 (N_22215,N_14867,N_11067);
nand U22216 (N_22216,N_17399,N_14607);
nand U22217 (N_22217,N_14009,N_11893);
nand U22218 (N_22218,N_10549,N_11764);
or U22219 (N_22219,N_13496,N_15432);
nand U22220 (N_22220,N_14047,N_10222);
and U22221 (N_22221,N_12583,N_18546);
or U22222 (N_22222,N_11925,N_12037);
or U22223 (N_22223,N_18761,N_17161);
nor U22224 (N_22224,N_14459,N_15842);
or U22225 (N_22225,N_10358,N_13791);
and U22226 (N_22226,N_10047,N_17455);
or U22227 (N_22227,N_11346,N_13555);
nor U22228 (N_22228,N_13659,N_13137);
nand U22229 (N_22229,N_18897,N_13828);
nor U22230 (N_22230,N_11546,N_10685);
nor U22231 (N_22231,N_13976,N_17989);
and U22232 (N_22232,N_15875,N_14168);
nand U22233 (N_22233,N_15765,N_14076);
nand U22234 (N_22234,N_13836,N_17949);
nand U22235 (N_22235,N_16798,N_11562);
nor U22236 (N_22236,N_16771,N_19278);
and U22237 (N_22237,N_13308,N_11240);
xor U22238 (N_22238,N_16718,N_11649);
and U22239 (N_22239,N_16704,N_18378);
or U22240 (N_22240,N_11415,N_13067);
nand U22241 (N_22241,N_18464,N_10674);
or U22242 (N_22242,N_19415,N_16424);
nand U22243 (N_22243,N_19456,N_18056);
and U22244 (N_22244,N_14945,N_17049);
nor U22245 (N_22245,N_10447,N_14167);
and U22246 (N_22246,N_19303,N_16398);
nor U22247 (N_22247,N_19454,N_11532);
nand U22248 (N_22248,N_13931,N_13629);
nor U22249 (N_22249,N_15145,N_14653);
nand U22250 (N_22250,N_10850,N_19556);
nor U22251 (N_22251,N_14025,N_18739);
xor U22252 (N_22252,N_17616,N_16457);
and U22253 (N_22253,N_18517,N_11854);
nor U22254 (N_22254,N_19333,N_19611);
or U22255 (N_22255,N_15476,N_16937);
or U22256 (N_22256,N_11005,N_14733);
nor U22257 (N_22257,N_13050,N_16687);
or U22258 (N_22258,N_14290,N_11303);
nor U22259 (N_22259,N_14145,N_18964);
and U22260 (N_22260,N_14533,N_14067);
and U22261 (N_22261,N_14586,N_15346);
nor U22262 (N_22262,N_19841,N_14209);
or U22263 (N_22263,N_14949,N_16507);
nor U22264 (N_22264,N_12803,N_13763);
or U22265 (N_22265,N_11359,N_13063);
nand U22266 (N_22266,N_10799,N_17674);
xor U22267 (N_22267,N_17098,N_14462);
and U22268 (N_22268,N_17016,N_13463);
and U22269 (N_22269,N_19185,N_15820);
and U22270 (N_22270,N_16110,N_17353);
nand U22271 (N_22271,N_10889,N_16065);
nor U22272 (N_22272,N_11287,N_19586);
and U22273 (N_22273,N_14298,N_12346);
nand U22274 (N_22274,N_18145,N_13510);
nor U22275 (N_22275,N_19321,N_18665);
xor U22276 (N_22276,N_16840,N_17885);
or U22277 (N_22277,N_12252,N_10185);
and U22278 (N_22278,N_14068,N_13563);
or U22279 (N_22279,N_14036,N_16409);
or U22280 (N_22280,N_13886,N_12481);
or U22281 (N_22281,N_12111,N_19075);
nor U22282 (N_22282,N_18181,N_13485);
nand U22283 (N_22283,N_12767,N_13235);
and U22284 (N_22284,N_17125,N_11245);
or U22285 (N_22285,N_11739,N_19443);
and U22286 (N_22286,N_19594,N_14446);
nor U22287 (N_22287,N_15779,N_19453);
nand U22288 (N_22288,N_12532,N_12985);
nand U22289 (N_22289,N_19506,N_12451);
or U22290 (N_22290,N_18453,N_10954);
nor U22291 (N_22291,N_16551,N_13892);
xnor U22292 (N_22292,N_10445,N_13440);
or U22293 (N_22293,N_18562,N_12845);
and U22294 (N_22294,N_18043,N_19777);
nand U22295 (N_22295,N_10959,N_13035);
and U22296 (N_22296,N_13609,N_19107);
nor U22297 (N_22297,N_10772,N_11783);
or U22298 (N_22298,N_18206,N_12338);
or U22299 (N_22299,N_13070,N_18986);
or U22300 (N_22300,N_14657,N_12791);
or U22301 (N_22301,N_19976,N_12233);
and U22302 (N_22302,N_19842,N_17374);
nor U22303 (N_22303,N_19539,N_18563);
nor U22304 (N_22304,N_17680,N_10913);
nand U22305 (N_22305,N_12670,N_16746);
or U22306 (N_22306,N_10773,N_11447);
or U22307 (N_22307,N_11433,N_19643);
or U22308 (N_22308,N_14138,N_12986);
or U22309 (N_22309,N_12227,N_19979);
nand U22310 (N_22310,N_18496,N_12179);
or U22311 (N_22311,N_16055,N_18242);
nor U22312 (N_22312,N_11044,N_10256);
nand U22313 (N_22313,N_17404,N_10369);
nand U22314 (N_22314,N_11418,N_16647);
nand U22315 (N_22315,N_14477,N_19455);
nand U22316 (N_22316,N_15205,N_11531);
nor U22317 (N_22317,N_11746,N_16703);
or U22318 (N_22318,N_10452,N_16552);
or U22319 (N_22319,N_18564,N_11062);
and U22320 (N_22320,N_10991,N_19664);
xor U22321 (N_22321,N_14627,N_13318);
nand U22322 (N_22322,N_16500,N_15026);
and U22323 (N_22323,N_19153,N_18577);
and U22324 (N_22324,N_18380,N_10961);
nand U22325 (N_22325,N_10584,N_12911);
and U22326 (N_22326,N_19514,N_13907);
and U22327 (N_22327,N_14319,N_13372);
or U22328 (N_22328,N_11722,N_17778);
and U22329 (N_22329,N_15097,N_10254);
nor U22330 (N_22330,N_19353,N_18787);
nor U22331 (N_22331,N_13590,N_18899);
nand U22332 (N_22332,N_18251,N_12871);
nor U22333 (N_22333,N_11732,N_19822);
xnor U22334 (N_22334,N_11080,N_17962);
xor U22335 (N_22335,N_13303,N_10314);
or U22336 (N_22336,N_18967,N_18132);
nand U22337 (N_22337,N_13105,N_19668);
nand U22338 (N_22338,N_14977,N_16072);
nor U22339 (N_22339,N_13000,N_16872);
and U22340 (N_22340,N_19876,N_14087);
nor U22341 (N_22341,N_16690,N_16863);
or U22342 (N_22342,N_12358,N_14860);
nand U22343 (N_22343,N_18417,N_13685);
nand U22344 (N_22344,N_16231,N_11027);
nand U22345 (N_22345,N_13033,N_15728);
nand U22346 (N_22346,N_16792,N_17151);
or U22347 (N_22347,N_12591,N_15182);
nand U22348 (N_22348,N_13518,N_11919);
xor U22349 (N_22349,N_13329,N_13120);
and U22350 (N_22350,N_12282,N_10172);
or U22351 (N_22351,N_18337,N_15492);
or U22352 (N_22352,N_16419,N_11070);
xnor U22353 (N_22353,N_12938,N_18214);
and U22354 (N_22354,N_16428,N_16992);
xor U22355 (N_22355,N_16667,N_15249);
or U22356 (N_22356,N_15383,N_11710);
nor U22357 (N_22357,N_18745,N_13709);
nor U22358 (N_22358,N_17855,N_16565);
and U22359 (N_22359,N_15915,N_15845);
and U22360 (N_22360,N_14115,N_13399);
nor U22361 (N_22361,N_13690,N_19803);
or U22362 (N_22362,N_15195,N_10097);
nor U22363 (N_22363,N_10354,N_14764);
xnor U22364 (N_22364,N_13772,N_19386);
and U22365 (N_22365,N_14111,N_13014);
or U22366 (N_22366,N_15550,N_16793);
and U22367 (N_22367,N_10394,N_19768);
nand U22368 (N_22368,N_11098,N_10969);
nor U22369 (N_22369,N_14350,N_13998);
xnor U22370 (N_22370,N_12248,N_17805);
xnor U22371 (N_22371,N_19588,N_15806);
and U22372 (N_22372,N_18735,N_12293);
nor U22373 (N_22373,N_19865,N_16155);
nand U22374 (N_22374,N_19685,N_17152);
or U22375 (N_22375,N_13121,N_10183);
and U22376 (N_22376,N_10068,N_11178);
nand U22377 (N_22377,N_15541,N_18829);
and U22378 (N_22378,N_11292,N_10582);
nand U22379 (N_22379,N_13715,N_15518);
xnor U22380 (N_22380,N_17438,N_16408);
nor U22381 (N_22381,N_19060,N_18687);
or U22382 (N_22382,N_18628,N_13064);
or U22383 (N_22383,N_19394,N_11045);
or U22384 (N_22384,N_12438,N_14188);
or U22385 (N_22385,N_18597,N_10979);
or U22386 (N_22386,N_11778,N_13203);
or U22387 (N_22387,N_14886,N_13071);
nor U22388 (N_22388,N_13523,N_15707);
nor U22389 (N_22389,N_19159,N_13499);
and U22390 (N_22390,N_18347,N_17729);
nand U22391 (N_22391,N_16327,N_17381);
nor U22392 (N_22392,N_17164,N_13767);
or U22393 (N_22393,N_13273,N_12574);
nor U22394 (N_22394,N_10190,N_10377);
nor U22395 (N_22395,N_13507,N_16563);
nand U22396 (N_22396,N_19509,N_18426);
or U22397 (N_22397,N_15165,N_19874);
nor U22398 (N_22398,N_11305,N_15537);
or U22399 (N_22399,N_12365,N_16393);
nand U22400 (N_22400,N_18939,N_18549);
xnor U22401 (N_22401,N_19629,N_18313);
xnor U22402 (N_22402,N_18470,N_13534);
nand U22403 (N_22403,N_12190,N_15174);
nor U22404 (N_22404,N_16206,N_13426);
and U22405 (N_22405,N_12238,N_10939);
xnor U22406 (N_22406,N_19371,N_13146);
and U22407 (N_22407,N_17097,N_13380);
and U22408 (N_22408,N_15671,N_10548);
nor U22409 (N_22409,N_10086,N_11481);
or U22410 (N_22410,N_17459,N_15269);
nand U22411 (N_22411,N_19270,N_15144);
nand U22412 (N_22412,N_14069,N_16290);
or U22413 (N_22413,N_17465,N_13215);
or U22414 (N_22414,N_10696,N_17804);
nor U22415 (N_22415,N_19218,N_17892);
nor U22416 (N_22416,N_16263,N_19463);
or U22417 (N_22417,N_13649,N_10813);
nor U22418 (N_22418,N_16977,N_12646);
nor U22419 (N_22419,N_17384,N_17273);
nand U22420 (N_22420,N_11227,N_11527);
nand U22421 (N_22421,N_11279,N_15632);
and U22422 (N_22422,N_19947,N_16471);
or U22423 (N_22423,N_11188,N_12364);
nor U22424 (N_22424,N_18196,N_15983);
or U22425 (N_22425,N_11256,N_11422);
and U22426 (N_22426,N_11978,N_18273);
nand U22427 (N_22427,N_15245,N_13687);
and U22428 (N_22428,N_19907,N_10919);
nor U22429 (N_22429,N_13289,N_13699);
and U22430 (N_22430,N_14304,N_13464);
xor U22431 (N_22431,N_19545,N_18842);
or U22432 (N_22432,N_12286,N_17700);
nand U22433 (N_22433,N_15996,N_18521);
nand U22434 (N_22434,N_17253,N_11150);
or U22435 (N_22435,N_17020,N_17796);
nand U22436 (N_22436,N_19630,N_11814);
or U22437 (N_22437,N_17821,N_17189);
xor U22438 (N_22438,N_16249,N_15958);
or U22439 (N_22439,N_19840,N_16331);
xor U22440 (N_22440,N_14049,N_10064);
nor U22441 (N_22441,N_17379,N_14569);
nor U22442 (N_22442,N_15552,N_13906);
and U22443 (N_22443,N_12058,N_14868);
and U22444 (N_22444,N_18655,N_13415);
and U22445 (N_22445,N_18864,N_17523);
nor U22446 (N_22446,N_11114,N_15442);
xnor U22447 (N_22447,N_19501,N_15539);
xor U22448 (N_22448,N_14696,N_18774);
and U22449 (N_22449,N_17878,N_15503);
or U22450 (N_22450,N_18601,N_18926);
nor U22451 (N_22451,N_13900,N_10564);
or U22452 (N_22452,N_14487,N_16856);
or U22453 (N_22453,N_18997,N_10410);
and U22454 (N_22454,N_19678,N_11780);
nand U22455 (N_22455,N_13242,N_19587);
nand U22456 (N_22456,N_10881,N_19585);
xnor U22457 (N_22457,N_16049,N_15716);
nor U22458 (N_22458,N_15823,N_17346);
nor U22459 (N_22459,N_13160,N_10844);
nand U22460 (N_22460,N_12200,N_16316);
nand U22461 (N_22461,N_16345,N_19101);
nor U22462 (N_22462,N_16150,N_15282);
or U22463 (N_22463,N_17709,N_15688);
and U22464 (N_22464,N_11129,N_13023);
nor U22465 (N_22465,N_19022,N_14971);
nand U22466 (N_22466,N_12795,N_18514);
xnor U22467 (N_22467,N_12572,N_13435);
and U22468 (N_22468,N_14323,N_14981);
or U22469 (N_22469,N_14997,N_14308);
nor U22470 (N_22470,N_15505,N_17849);
nor U22471 (N_22471,N_16163,N_18753);
nor U22472 (N_22472,N_12746,N_19683);
and U22473 (N_22473,N_18884,N_15594);
or U22474 (N_22474,N_10608,N_10304);
nand U22475 (N_22475,N_12090,N_19311);
or U22476 (N_22476,N_17081,N_13672);
nor U22477 (N_22477,N_18835,N_18732);
or U22478 (N_22478,N_15452,N_10146);
nor U22479 (N_22479,N_17787,N_15627);
nor U22480 (N_22480,N_11905,N_16680);
or U22481 (N_22481,N_13364,N_10329);
nor U22482 (N_22482,N_10459,N_16188);
nand U22483 (N_22483,N_11362,N_13864);
or U22484 (N_22484,N_12374,N_13268);
nand U22485 (N_22485,N_14775,N_10052);
or U22486 (N_22486,N_17480,N_11185);
and U22487 (N_22487,N_10505,N_12919);
nand U22488 (N_22488,N_14904,N_19792);
nand U22489 (N_22489,N_10181,N_19261);
nor U22490 (N_22490,N_10002,N_17326);
or U22491 (N_22491,N_16394,N_18718);
xor U22492 (N_22492,N_13811,N_18931);
or U22493 (N_22493,N_19624,N_14092);
nand U22494 (N_22494,N_19682,N_17090);
or U22495 (N_22495,N_15878,N_15730);
or U22496 (N_22496,N_10646,N_14915);
nand U22497 (N_22497,N_10653,N_13732);
or U22498 (N_22498,N_19809,N_17840);
nand U22499 (N_22499,N_19614,N_14980);
and U22500 (N_22500,N_11834,N_19485);
or U22501 (N_22501,N_19590,N_19074);
nor U22502 (N_22502,N_14279,N_12138);
and U22503 (N_22503,N_15382,N_17202);
nand U22504 (N_22504,N_16655,N_13019);
nor U22505 (N_22505,N_12950,N_16843);
xor U22506 (N_22506,N_17820,N_16446);
nor U22507 (N_22507,N_18874,N_12722);
and U22508 (N_22508,N_14506,N_11226);
and U22509 (N_22509,N_17777,N_12061);
or U22510 (N_22510,N_18958,N_16499);
nand U22511 (N_22511,N_18154,N_15056);
nand U22512 (N_22512,N_11691,N_15960);
nor U22513 (N_22513,N_19385,N_16832);
nand U22514 (N_22514,N_13671,N_15341);
xor U22515 (N_22515,N_13815,N_16685);
nor U22516 (N_22516,N_12959,N_17248);
nor U22517 (N_22517,N_16634,N_15602);
nor U22518 (N_22518,N_16229,N_15686);
and U22519 (N_22519,N_15183,N_15921);
nand U22520 (N_22520,N_16760,N_11056);
nand U22521 (N_22521,N_19363,N_11443);
and U22522 (N_22522,N_13512,N_17598);
nand U22523 (N_22523,N_10310,N_10227);
nor U22524 (N_22524,N_10105,N_10046);
nor U22525 (N_22525,N_16221,N_12182);
nand U22526 (N_22526,N_19617,N_15416);
and U22527 (N_22527,N_15538,N_15535);
nor U22528 (N_22528,N_15290,N_11427);
nor U22529 (N_22529,N_12384,N_15338);
and U22530 (N_22530,N_14560,N_13983);
nand U22531 (N_22531,N_11099,N_16750);
nand U22532 (N_22532,N_16147,N_17827);
and U22533 (N_22533,N_14197,N_13448);
nor U22534 (N_22534,N_12319,N_18545);
nand U22535 (N_22535,N_13346,N_16461);
or U22536 (N_22536,N_14124,N_19378);
and U22537 (N_22537,N_15702,N_14762);
or U22538 (N_22538,N_12429,N_17525);
nand U22539 (N_22539,N_16162,N_10006);
nor U22540 (N_22540,N_11274,N_18932);
nor U22541 (N_22541,N_17509,N_10194);
xnor U22542 (N_22542,N_12433,N_18031);
and U22543 (N_22543,N_16351,N_17246);
nand U22544 (N_22544,N_17112,N_11913);
or U22545 (N_22545,N_11140,N_11593);
or U22546 (N_22546,N_18565,N_11087);
nand U22547 (N_22547,N_16280,N_17426);
nor U22548 (N_22548,N_17117,N_17014);
nand U22549 (N_22549,N_15756,N_15181);
nor U22550 (N_22550,N_10125,N_15630);
nand U22551 (N_22551,N_16770,N_13443);
nand U22552 (N_22552,N_12475,N_13865);
nand U22553 (N_22553,N_16842,N_16191);
and U22554 (N_22554,N_13650,N_12903);
or U22555 (N_22555,N_18794,N_16639);
or U22556 (N_22556,N_11156,N_12779);
and U22557 (N_22557,N_12766,N_11614);
and U22558 (N_22558,N_12155,N_19523);
nor U22559 (N_22559,N_10926,N_15972);
nand U22560 (N_22560,N_13809,N_16051);
or U22561 (N_22561,N_16473,N_16698);
nor U22562 (N_22562,N_18849,N_17846);
or U22563 (N_22563,N_18930,N_10620);
nor U22564 (N_22564,N_11294,N_19213);
and U22565 (N_22565,N_10518,N_10299);
xnor U22566 (N_22566,N_16488,N_10018);
nand U22567 (N_22567,N_11088,N_15068);
nand U22568 (N_22568,N_19100,N_14863);
or U22569 (N_22569,N_18479,N_15942);
nand U22570 (N_22570,N_15885,N_14412);
nand U22571 (N_22571,N_15797,N_17572);
and U22572 (N_22572,N_12527,N_15924);
nor U22573 (N_22573,N_19551,N_15350);
or U22574 (N_22574,N_11632,N_16969);
and U22575 (N_22575,N_10305,N_17350);
nand U22576 (N_22576,N_16482,N_12649);
nor U22577 (N_22577,N_13944,N_17946);
and U22578 (N_22578,N_19910,N_19263);
nor U22579 (N_22579,N_10750,N_10957);
nor U22580 (N_22580,N_15101,N_10659);
xnor U22581 (N_22581,N_15073,N_18202);
or U22582 (N_22582,N_16849,N_10219);
nor U22583 (N_22583,N_17187,N_12339);
nor U22584 (N_22584,N_12044,N_14547);
or U22585 (N_22585,N_11394,N_19000);
nor U22586 (N_22586,N_15263,N_15803);
xnor U22587 (N_22587,N_12418,N_12726);
nand U22588 (N_22588,N_18891,N_12664);
xor U22589 (N_22589,N_15394,N_14265);
or U22590 (N_22590,N_15466,N_18614);
nor U22591 (N_22591,N_19015,N_14557);
nand U22592 (N_22592,N_15980,N_15046);
xor U22593 (N_22593,N_18234,N_15912);
nor U22594 (N_22594,N_15367,N_17262);
or U22595 (N_22595,N_19515,N_13131);
nand U22596 (N_22596,N_12991,N_17483);
nor U22597 (N_22597,N_11955,N_17800);
nand U22598 (N_22598,N_19215,N_15793);
nand U22599 (N_22599,N_12852,N_17127);
or U22600 (N_22600,N_12773,N_19008);
nor U22601 (N_22601,N_10088,N_13378);
nor U22602 (N_22602,N_15581,N_14934);
and U22603 (N_22603,N_12096,N_13940);
nand U22604 (N_22604,N_16151,N_18268);
nand U22605 (N_22605,N_18539,N_15057);
nand U22606 (N_22606,N_12686,N_11408);
xor U22607 (N_22607,N_13165,N_11830);
xor U22608 (N_22608,N_11265,N_17972);
nand U22609 (N_22609,N_18850,N_10008);
or U22610 (N_22610,N_19309,N_16420);
xor U22611 (N_22611,N_15854,N_12971);
nand U22612 (N_22612,N_10024,N_11133);
nor U22613 (N_22613,N_13562,N_16967);
and U22614 (N_22614,N_19366,N_13269);
nand U22615 (N_22615,N_14046,N_18639);
and U22616 (N_22616,N_11177,N_19727);
and U22617 (N_22617,N_15979,N_13710);
nand U22618 (N_22618,N_11183,N_12718);
or U22619 (N_22619,N_17174,N_11320);
and U22620 (N_22620,N_13718,N_16802);
or U22621 (N_22621,N_13142,N_14442);
and U22622 (N_22622,N_10931,N_17691);
nand U22623 (N_22623,N_17981,N_14743);
and U22624 (N_22624,N_11670,N_18476);
xnor U22625 (N_22625,N_13103,N_13947);
nor U22626 (N_22626,N_12925,N_13988);
or U22627 (N_22627,N_14513,N_18828);
or U22628 (N_22628,N_15596,N_15124);
and U22629 (N_22629,N_10188,N_19211);
nor U22630 (N_22630,N_13386,N_13462);
nor U22631 (N_22631,N_18707,N_19268);
nor U22632 (N_22632,N_10208,N_14064);
nor U22633 (N_22633,N_19957,N_14213);
nand U22634 (N_22634,N_11212,N_17602);
nand U22635 (N_22635,N_18303,N_17627);
nand U22636 (N_22636,N_19656,N_13726);
nand U22637 (N_22637,N_11318,N_14509);
nor U22638 (N_22638,N_19648,N_19287);
nand U22639 (N_22639,N_15243,N_14967);
or U22640 (N_22640,N_12839,N_12136);
nand U22641 (N_22641,N_18006,N_19819);
and U22642 (N_22642,N_11356,N_10218);
xor U22643 (N_22643,N_16275,N_16102);
nor U22644 (N_22644,N_11041,N_18180);
nand U22645 (N_22645,N_11411,N_17105);
and U22646 (N_22646,N_10163,N_14277);
xnor U22647 (N_22647,N_18768,N_14963);
nand U22648 (N_22648,N_19190,N_16118);
nand U22649 (N_22649,N_13124,N_19116);
and U22650 (N_22650,N_13056,N_19845);
and U22651 (N_22651,N_14096,N_11682);
nor U22652 (N_22652,N_14612,N_19913);
nand U22653 (N_22653,N_13930,N_18764);
and U22654 (N_22654,N_15347,N_13051);
or U22655 (N_22655,N_18830,N_16576);
xor U22656 (N_22656,N_14858,N_11631);
xor U22657 (N_22657,N_15344,N_19802);
or U22658 (N_22658,N_14839,N_14898);
nor U22659 (N_22659,N_12952,N_18062);
nand U22660 (N_22660,N_17811,N_17009);
and U22661 (N_22661,N_14428,N_17140);
and U22662 (N_22662,N_19699,N_19520);
nor U22663 (N_22663,N_14792,N_15226);
or U22664 (N_22664,N_18375,N_14198);
and U22665 (N_22665,N_10037,N_14200);
nor U22666 (N_22666,N_12002,N_14295);
or U22667 (N_22667,N_14735,N_13634);
nand U22668 (N_22668,N_12221,N_18127);
xnor U22669 (N_22669,N_15489,N_11564);
nand U22670 (N_22670,N_19433,N_15831);
and U22671 (N_22671,N_13597,N_11622);
and U22672 (N_22672,N_18123,N_16493);
and U22673 (N_22673,N_19798,N_18737);
or U22674 (N_22674,N_11715,N_12857);
nand U22675 (N_22675,N_16605,N_19914);
xor U22676 (N_22676,N_16530,N_13538);
nand U22677 (N_22677,N_15077,N_11453);
nor U22678 (N_22678,N_13387,N_14173);
and U22679 (N_22679,N_19119,N_12435);
or U22680 (N_22680,N_11254,N_14846);
and U22681 (N_22681,N_19359,N_13912);
or U22682 (N_22682,N_11811,N_11389);
xor U22683 (N_22683,N_18561,N_15843);
nor U22684 (N_22684,N_17992,N_13909);
nor U22685 (N_22685,N_19023,N_13877);
and U22686 (N_22686,N_13264,N_14559);
and U22687 (N_22687,N_14004,N_16571);
or U22688 (N_22688,N_17064,N_19661);
xor U22689 (N_22689,N_19906,N_16030);
nor U22690 (N_22690,N_19956,N_17502);
and U22691 (N_22691,N_12823,N_13300);
nor U22692 (N_22692,N_14845,N_13299);
nor U22693 (N_22693,N_17434,N_12473);
nor U22694 (N_22694,N_13254,N_15425);
nand U22695 (N_22695,N_10903,N_14978);
nor U22696 (N_22696,N_13361,N_11055);
or U22697 (N_22697,N_14616,N_10187);
and U22698 (N_22698,N_16734,N_10877);
xor U22699 (N_22699,N_12893,N_15397);
nor U22700 (N_22700,N_12071,N_15850);
nand U22701 (N_22701,N_17054,N_18477);
and U22702 (N_22702,N_12505,N_17297);
and U22703 (N_22703,N_18624,N_17676);
nor U22704 (N_22704,N_15696,N_15829);
nor U22705 (N_22705,N_16970,N_10235);
and U22706 (N_22706,N_17490,N_14226);
and U22707 (N_22707,N_16848,N_12951);
and U22708 (N_22708,N_15853,N_10350);
nor U22709 (N_22709,N_15206,N_16962);
nor U22710 (N_22710,N_19429,N_17717);
nor U22711 (N_22711,N_12160,N_12811);
and U22712 (N_22712,N_12404,N_12926);
nand U22713 (N_22713,N_10414,N_14523);
and U22714 (N_22714,N_16397,N_14956);
or U22715 (N_22715,N_10600,N_11624);
and U22716 (N_22716,N_16399,N_16543);
xnor U22717 (N_22717,N_17725,N_14953);
and U22718 (N_22718,N_12291,N_16416);
nor U22719 (N_22719,N_15665,N_19080);
and U22720 (N_22720,N_18504,N_11840);
nor U22721 (N_22721,N_15230,N_17085);
and U22722 (N_22722,N_13895,N_12701);
or U22723 (N_22723,N_16217,N_19223);
nor U22724 (N_22724,N_19691,N_18195);
and U22725 (N_22725,N_10545,N_18025);
or U22726 (N_22726,N_16385,N_13611);
nor U22727 (N_22727,N_19843,N_16094);
nor U22728 (N_22728,N_15588,N_18598);
and U22729 (N_22729,N_14423,N_19983);
or U22730 (N_22730,N_12860,N_17099);
xnor U22731 (N_22731,N_11578,N_11057);
nor U22732 (N_22732,N_13833,N_13049);
or U22733 (N_22733,N_19542,N_16749);
xnor U22734 (N_22734,N_18345,N_16520);
nand U22735 (N_22735,N_10640,N_14451);
xnor U22736 (N_22736,N_10273,N_11676);
nand U22737 (N_22737,N_10301,N_12086);
nand U22738 (N_22738,N_12621,N_17106);
or U22739 (N_22739,N_18440,N_19423);
nor U22740 (N_22740,N_19749,N_19469);
nand U22741 (N_22741,N_14141,N_17215);
and U22742 (N_22742,N_12450,N_18178);
nor U22743 (N_22743,N_19180,N_15100);
xor U22744 (N_22744,N_13294,N_14435);
or U22745 (N_22745,N_14396,N_13725);
nand U22746 (N_22746,N_17155,N_18812);
or U22747 (N_22747,N_11861,N_10722);
nand U22748 (N_22748,N_15609,N_10434);
nand U22749 (N_22749,N_17392,N_13511);
nor U22750 (N_22750,N_13096,N_17453);
nand U22751 (N_22751,N_10417,N_19716);
xnor U22752 (N_22752,N_13888,N_15761);
or U22753 (N_22753,N_19606,N_19952);
nor U22754 (N_22754,N_14655,N_13697);
nor U22755 (N_22755,N_17617,N_11954);
nor U22756 (N_22756,N_14532,N_17570);
and U22757 (N_22757,N_13292,N_12035);
and U22758 (N_22758,N_12116,N_18809);
or U22759 (N_22759,N_15018,N_11431);
or U22760 (N_22760,N_10888,N_19003);
nand U22761 (N_22761,N_17439,N_16477);
or U22762 (N_22762,N_13698,N_16620);
and U22763 (N_22763,N_11582,N_12749);
and U22764 (N_22764,N_14420,N_15052);
and U22765 (N_22765,N_11151,N_11943);
nor U22766 (N_22766,N_12048,N_12120);
or U22767 (N_22767,N_14382,N_17069);
nor U22768 (N_22768,N_16681,N_11166);
or U22769 (N_22769,N_18397,N_16145);
or U22770 (N_22770,N_11663,N_18116);
nand U22771 (N_22771,N_18129,N_14592);
nand U22772 (N_22772,N_10571,N_15067);
or U22773 (N_22773,N_13086,N_13832);
and U22774 (N_22774,N_16695,N_14924);
nand U22775 (N_22775,N_11735,N_12321);
or U22776 (N_22776,N_14392,N_17218);
and U22777 (N_22777,N_10236,N_14993);
and U22778 (N_22778,N_16115,N_13334);
nor U22779 (N_22779,N_15435,N_19600);
nor U22780 (N_22780,N_19555,N_15762);
nor U22781 (N_22781,N_11465,N_10666);
nand U22782 (N_22782,N_10712,N_11373);
or U22783 (N_22783,N_16011,N_17870);
nor U22784 (N_22784,N_16763,N_14316);
or U22785 (N_22785,N_14075,N_15474);
or U22786 (N_22786,N_17357,N_14468);
nand U22787 (N_22787,N_11904,N_10032);
or U22788 (N_22788,N_18045,N_11317);
nor U22789 (N_22789,N_14836,N_12638);
or U22790 (N_22790,N_18638,N_11709);
nand U22791 (N_22791,N_10313,N_19695);
or U22792 (N_22792,N_11314,N_10592);
or U22793 (N_22793,N_16436,N_18683);
nor U22794 (N_22794,N_19424,N_12775);
nor U22795 (N_22795,N_10992,N_16256);
xnor U22796 (N_22796,N_16766,N_10214);
nor U22797 (N_22797,N_11786,N_18128);
nand U22798 (N_22798,N_17290,N_11172);
nand U22799 (N_22799,N_14358,N_15949);
nand U22800 (N_22800,N_17170,N_11332);
or U22801 (N_22801,N_10838,N_17810);
and U22802 (N_22802,N_16759,N_10308);
nand U22803 (N_22803,N_18055,N_11089);
or U22804 (N_22804,N_10500,N_16323);
or U22805 (N_22805,N_11690,N_19733);
nor U22806 (N_22806,N_12474,N_18532);
nor U22807 (N_22807,N_18350,N_10626);
nor U22808 (N_22808,N_13057,N_15312);
and U22809 (N_22809,N_11082,N_17275);
nor U22810 (N_22810,N_16184,N_17636);
and U22811 (N_22811,N_18747,N_19711);
nor U22812 (N_22812,N_10697,N_14322);
and U22813 (N_22813,N_16553,N_11720);
or U22814 (N_22814,N_13135,N_19372);
nand U22815 (N_22815,N_13601,N_12672);
nand U22816 (N_22816,N_10440,N_17372);
and U22817 (N_22817,N_14099,N_17826);
or U22818 (N_22818,N_14902,N_19619);
and U22819 (N_22819,N_17854,N_10667);
nor U22820 (N_22820,N_18843,N_19140);
and U22821 (N_22821,N_16084,N_15561);
nor U22822 (N_22822,N_13054,N_19053);
or U22823 (N_22823,N_11890,N_18917);
and U22824 (N_22824,N_19202,N_16591);
nand U22825 (N_22825,N_19240,N_11479);
and U22826 (N_22826,N_17693,N_12558);
or U22827 (N_22827,N_14022,N_13288);
and U22828 (N_22828,N_10753,N_13138);
nand U22829 (N_22829,N_18072,N_17206);
nand U22830 (N_22830,N_18404,N_11334);
nand U22831 (N_22831,N_15859,N_10199);
nand U22832 (N_22832,N_11423,N_15045);
or U22833 (N_22833,N_10764,N_11962);
xnor U22834 (N_22834,N_11381,N_14516);
and U22835 (N_22835,N_10673,N_10107);
or U22836 (N_22836,N_14717,N_17415);
nor U22837 (N_22837,N_12471,N_12598);
nand U22838 (N_22838,N_16298,N_12332);
and U22839 (N_22839,N_12828,N_19692);
or U22840 (N_22840,N_18807,N_15006);
nor U22841 (N_22841,N_15796,N_14101);
nand U22842 (N_22842,N_15939,N_10334);
and U22843 (N_22843,N_11679,N_19030);
nor U22844 (N_22844,N_11122,N_18001);
or U22845 (N_22845,N_13941,N_16670);
or U22846 (N_22846,N_11262,N_12085);
nand U22847 (N_22847,N_18893,N_11219);
nand U22848 (N_22848,N_18497,N_11376);
xnor U22849 (N_22849,N_12904,N_16425);
and U22850 (N_22850,N_13663,N_10536);
nand U22851 (N_22851,N_15764,N_11923);
nand U22852 (N_22852,N_16113,N_14003);
or U22853 (N_22853,N_12819,N_10476);
nand U22854 (N_22854,N_19746,N_19866);
or U22855 (N_22855,N_10160,N_11120);
nand U22856 (N_22856,N_10487,N_11475);
and U22857 (N_22857,N_19088,N_14205);
nor U22858 (N_22858,N_17652,N_18465);
or U22859 (N_22859,N_10809,N_12413);
and U22860 (N_22860,N_11130,N_18481);
and U22861 (N_22861,N_18454,N_12659);
nor U22862 (N_22862,N_18854,N_10098);
and U22863 (N_22863,N_13126,N_19091);
xor U22864 (N_22864,N_18650,N_13688);
and U22865 (N_22865,N_10264,N_15186);
xor U22866 (N_22866,N_17518,N_18237);
nor U22867 (N_22867,N_15371,N_10550);
and U22868 (N_22868,N_12033,N_15569);
and U22869 (N_22869,N_19761,N_10200);
or U22870 (N_22870,N_13894,N_12604);
nand U22871 (N_22871,N_17952,N_10747);
nor U22872 (N_22872,N_15364,N_13614);
xnor U22873 (N_22873,N_15993,N_16130);
and U22874 (N_22874,N_10781,N_15472);
nand U22875 (N_22875,N_12577,N_18431);
nand U22876 (N_22876,N_14899,N_18797);
nand U22877 (N_22877,N_16202,N_18107);
nor U22878 (N_22878,N_14765,N_15204);
or U22879 (N_22879,N_16684,N_19578);
nand U22880 (N_22880,N_17604,N_17277);
nand U22881 (N_22881,N_18302,N_13679);
or U22882 (N_22882,N_14475,N_15087);
and U22883 (N_22883,N_12455,N_13248);
xor U22884 (N_22884,N_10628,N_14356);
nor U22885 (N_22885,N_19955,N_10789);
nor U22886 (N_22886,N_10387,N_16527);
and U22887 (N_22887,N_16533,N_11538);
or U22888 (N_22888,N_19518,N_10963);
nand U22889 (N_22889,N_19863,N_11081);
and U22890 (N_22890,N_18533,N_13366);
and U22891 (N_22891,N_10739,N_18633);
nand U22892 (N_22892,N_15477,N_13398);
or U22893 (N_22893,N_18330,N_16933);
nand U22894 (N_22894,N_16660,N_18028);
nor U22895 (N_22895,N_16927,N_13267);
nand U22896 (N_22896,N_12152,N_17124);
or U22897 (N_22897,N_16824,N_18620);
nand U22898 (N_22898,N_18606,N_16985);
nor U22899 (N_22899,N_19892,N_11171);
and U22900 (N_22900,N_12206,N_14421);
nand U22901 (N_22901,N_19112,N_18708);
and U22902 (N_22902,N_16333,N_16494);
nand U22903 (N_22903,N_15673,N_17171);
nand U22904 (N_22904,N_17091,N_12222);
xor U22905 (N_22905,N_13946,N_19405);
xnor U22906 (N_22906,N_12132,N_15146);
nor U22907 (N_22907,N_13405,N_10338);
nand U22908 (N_22908,N_17468,N_15994);
or U22909 (N_22909,N_11845,N_14514);
xor U22910 (N_22910,N_10272,N_11630);
xnor U22911 (N_22911,N_13216,N_18607);
nand U22912 (N_22912,N_11877,N_13535);
nand U22913 (N_22913,N_13905,N_16046);
or U22914 (N_22914,N_15920,N_18265);
nor U22915 (N_22915,N_17808,N_16481);
nand U22916 (N_22916,N_12027,N_15359);
nor U22917 (N_22917,N_15669,N_18086);
nand U22918 (N_22918,N_19530,N_16106);
nand U22919 (N_22919,N_16873,N_12193);
and U22920 (N_22920,N_13719,N_10267);
or U22921 (N_22921,N_15567,N_11487);
and U22922 (N_22922,N_12794,N_19237);
xnor U22923 (N_22923,N_15978,N_13744);
nor U22924 (N_22924,N_16014,N_16797);
nand U22925 (N_22925,N_17561,N_19064);
nand U22926 (N_22926,N_12018,N_19820);
and U22927 (N_22927,N_11509,N_17243);
nand U22928 (N_22928,N_17932,N_11669);
xnor U22929 (N_22929,N_19285,N_11519);
nand U22930 (N_22930,N_14986,N_19148);
xnor U22931 (N_22931,N_14907,N_15400);
and U22932 (N_22932,N_10036,N_15391);
and U22933 (N_22933,N_16677,N_19390);
or U22934 (N_22934,N_16413,N_17162);
nor U22935 (N_22935,N_12982,N_18942);
nor U22936 (N_22936,N_14116,N_17872);
and U22937 (N_22937,N_12514,N_11916);
nor U22938 (N_22938,N_13151,N_10005);
nand U22939 (N_22939,N_17882,N_10295);
xnor U22940 (N_22940,N_11079,N_14311);
nand U22941 (N_22941,N_12333,N_16024);
xor U22942 (N_22942,N_12831,N_15040);
or U22943 (N_22943,N_15560,N_13524);
nor U22944 (N_22944,N_12063,N_19345);
and U22945 (N_22945,N_14932,N_12203);
and U22946 (N_22946,N_17338,N_10444);
and U22947 (N_22947,N_12310,N_14286);
or U22948 (N_22948,N_13885,N_12563);
or U22949 (N_22949,N_11300,N_16654);
nand U22950 (N_22950,N_13796,N_13099);
or U22951 (N_22951,N_12483,N_17165);
or U22952 (N_22952,N_15573,N_17466);
nor U22953 (N_22953,N_18722,N_18391);
or U22954 (N_22954,N_16196,N_12978);
xor U22955 (N_22955,N_17716,N_10864);
and U22956 (N_22956,N_11040,N_15828);
nand U22957 (N_22957,N_16152,N_15008);
nor U22958 (N_22958,N_16089,N_10019);
xor U22959 (N_22959,N_18992,N_16067);
xor U22960 (N_22960,N_17529,N_12159);
and U22961 (N_22961,N_10601,N_10496);
nand U22962 (N_22962,N_16142,N_17639);
xor U22963 (N_22963,N_11393,N_18974);
xor U22964 (N_22964,N_12607,N_19615);
or U22965 (N_22965,N_10428,N_18370);
or U22966 (N_22966,N_12081,N_17818);
nand U22967 (N_22967,N_17216,N_12172);
nor U22968 (N_22968,N_10784,N_17661);
nand U22969 (N_22969,N_18837,N_14230);
nand U22970 (N_22970,N_12208,N_10021);
nor U22971 (N_22971,N_10754,N_11708);
and U22972 (N_22972,N_17917,N_12257);
and U22973 (N_22973,N_19903,N_17238);
nor U22974 (N_22974,N_18982,N_11880);
xnor U22975 (N_22975,N_12329,N_17504);
xnor U22976 (N_22976,N_19106,N_18120);
or U22977 (N_22977,N_13953,N_12045);
and U22978 (N_22978,N_16111,N_16255);
or U22979 (N_22979,N_13407,N_10474);
nand U22980 (N_22980,N_11096,N_17159);
and U22981 (N_22981,N_10984,N_14494);
nor U22982 (N_22982,N_11128,N_10742);
xor U22983 (N_22983,N_19316,N_15283);
or U22984 (N_22984,N_19779,N_19560);
nand U22985 (N_22985,N_11608,N_10832);
and U22986 (N_22986,N_10645,N_19855);
nand U22987 (N_22987,N_17983,N_14697);
nand U22988 (N_22988,N_16483,N_19773);
nor U22989 (N_22989,N_13747,N_18963);
nor U22990 (N_22990,N_11609,N_16810);
and U22991 (N_22991,N_14706,N_11858);
nor U22992 (N_22992,N_15468,N_11606);
nand U22993 (N_22993,N_10081,N_10381);
or U22994 (N_22994,N_13436,N_16279);
xnor U22995 (N_22995,N_15177,N_15148);
or U22996 (N_22996,N_19312,N_18065);
nand U22997 (N_22997,N_14617,N_10115);
and U22998 (N_22998,N_18176,N_19032);
nor U22999 (N_22999,N_13777,N_17166);
nand U23000 (N_23000,N_18727,N_15600);
nor U23001 (N_23001,N_16701,N_18788);
nand U23002 (N_23002,N_13209,N_12260);
and U23003 (N_23003,N_15118,N_15015);
or U23004 (N_23004,N_12515,N_12196);
nor U23005 (N_23005,N_11035,N_18767);
or U23006 (N_23006,N_14398,N_13383);
xnor U23007 (N_23007,N_18240,N_17690);
or U23008 (N_23008,N_13677,N_14887);
nand U23009 (N_23009,N_10911,N_17710);
and U23010 (N_23010,N_19335,N_14705);
or U23011 (N_23011,N_18736,N_10043);
nand U23012 (N_23012,N_11289,N_15988);
nand U23013 (N_23013,N_13668,N_13298);
nand U23014 (N_23014,N_12969,N_10570);
nor U23015 (N_23015,N_17937,N_19306);
xnor U23016 (N_23016,N_18058,N_11445);
or U23017 (N_23017,N_12835,N_12760);
nand U23018 (N_23018,N_12444,N_17296);
or U23019 (N_23019,N_13746,N_17035);
and U23020 (N_23020,N_16253,N_10059);
nand U23021 (N_23021,N_13343,N_18892);
nor U23022 (N_23022,N_10700,N_16123);
nand U23023 (N_23023,N_15293,N_10675);
xor U23024 (N_23024,N_16383,N_14238);
and U23025 (N_23025,N_14647,N_14675);
nand U23026 (N_23026,N_17943,N_15540);
and U23027 (N_23027,N_15086,N_16434);
or U23028 (N_23028,N_16626,N_10513);
nand U23029 (N_23029,N_13469,N_15621);
or U23030 (N_23030,N_15261,N_19580);
nand U23031 (N_23031,N_13279,N_15280);
or U23032 (N_23032,N_10077,N_17454);
nor U23033 (N_23033,N_15130,N_11182);
or U23034 (N_23034,N_14712,N_11772);
xnor U23035 (N_23035,N_12570,N_19442);
nor U23036 (N_23036,N_10058,N_16738);
nor U23037 (N_23037,N_18895,N_12606);
and U23038 (N_23038,N_15495,N_15171);
or U23039 (N_23039,N_14199,N_14207);
xor U23040 (N_23040,N_10405,N_16492);
nand U23041 (N_23041,N_19065,N_17592);
nand U23042 (N_23042,N_17635,N_19921);
and U23043 (N_23043,N_12980,N_17135);
and U23044 (N_23044,N_14485,N_11416);
nor U23045 (N_23045,N_12279,N_12236);
nor U23046 (N_23046,N_14809,N_12932);
and U23047 (N_23047,N_15926,N_14105);
nor U23048 (N_23048,N_13730,N_14015);
or U23049 (N_23049,N_14856,N_10866);
and U23050 (N_23050,N_14527,N_18231);
xnor U23051 (N_23051,N_19669,N_19365);
xor U23052 (N_23052,N_10000,N_14163);
nand U23053 (N_23053,N_19395,N_13625);
and U23054 (N_23054,N_14122,N_10767);
nand U23055 (N_23055,N_17541,N_18087);
nand U23056 (N_23056,N_10994,N_10244);
nand U23057 (N_23057,N_12741,N_12547);
and U23058 (N_23058,N_14679,N_16004);
nor U23059 (N_23059,N_18040,N_10150);
nor U23060 (N_23060,N_15390,N_11179);
nor U23061 (N_23061,N_10210,N_13195);
or U23062 (N_23062,N_13794,N_10854);
xor U23063 (N_23063,N_16650,N_16532);
nor U23064 (N_23064,N_18199,N_15374);
nand U23065 (N_23065,N_10231,N_17142);
nand U23066 (N_23066,N_10148,N_14598);
nand U23067 (N_23067,N_14187,N_19193);
nor U23068 (N_23068,N_13738,N_12617);
or U23069 (N_23069,N_15469,N_16182);
or U23070 (N_23070,N_15184,N_18446);
nand U23071 (N_23071,N_10362,N_12181);
nand U23072 (N_23072,N_13238,N_10706);
or U23073 (N_23073,N_13202,N_11552);
nand U23074 (N_23074,N_18105,N_17148);
or U23075 (N_23075,N_16209,N_14588);
nand U23076 (N_23076,N_13514,N_17028);
and U23077 (N_23077,N_16222,N_15768);
or U23078 (N_23078,N_18364,N_19869);
nor U23079 (N_23079,N_18661,N_12251);
or U23080 (N_23080,N_15549,N_12209);
nor U23081 (N_23081,N_14785,N_12135);
nor U23082 (N_23082,N_19489,N_16056);
xor U23083 (N_23083,N_12476,N_12095);
and U23084 (N_23084,N_19438,N_14821);
nand U23085 (N_23085,N_15989,N_16883);
nor U23086 (N_23086,N_17060,N_18119);
and U23087 (N_23087,N_17839,N_16352);
nor U23088 (N_23088,N_12753,N_13917);
nor U23089 (N_23089,N_13043,N_10785);
nor U23090 (N_23090,N_19041,N_11223);
and U23091 (N_23091,N_16234,N_13637);
nor U23092 (N_23092,N_14834,N_10874);
or U23093 (N_23093,N_12882,N_17395);
and U23094 (N_23094,N_17741,N_16092);
nand U23095 (N_23095,N_15210,N_18104);
and U23096 (N_23096,N_16297,N_18149);
nand U23097 (N_23097,N_11345,N_16064);
xor U23098 (N_23098,N_10804,N_14280);
and U23099 (N_23099,N_14385,N_15264);
or U23100 (N_23100,N_16427,N_13098);
nand U23101 (N_23101,N_15619,N_12737);
or U23102 (N_23102,N_19432,N_16267);
or U23103 (N_23103,N_15437,N_16587);
nand U23104 (N_23104,N_10140,N_14823);
and U23105 (N_23105,N_10090,N_13130);
and U23106 (N_23106,N_19890,N_14021);
xnor U23107 (N_23107,N_12217,N_16982);
or U23108 (N_23108,N_17078,N_18126);
or U23109 (N_23109,N_16726,N_19867);
xor U23110 (N_23110,N_18603,N_10245);
and U23111 (N_23111,N_17307,N_15212);
nand U23112 (N_23112,N_16375,N_17727);
or U23113 (N_23113,N_14888,N_16939);
nand U23114 (N_23114,N_15890,N_17083);
nor U23115 (N_23115,N_11015,N_11258);
or U23116 (N_23116,N_19589,N_19344);
or U23117 (N_23117,N_19299,N_10614);
nand U23118 (N_23118,N_11637,N_10062);
nor U23119 (N_23119,N_17957,N_19362);
nor U23120 (N_23120,N_18806,N_19970);
and U23121 (N_23121,N_11116,N_10519);
nand U23122 (N_23122,N_10871,N_11500);
and U23123 (N_23123,N_10147,N_13097);
nand U23124 (N_23124,N_10818,N_10578);
nand U23125 (N_23125,N_10808,N_14144);
xor U23126 (N_23126,N_19288,N_15103);
xor U23127 (N_23127,N_17699,N_10292);
or U23128 (N_23128,N_17344,N_11705);
or U23129 (N_23129,N_10650,N_18325);
and U23130 (N_23130,N_17160,N_18642);
nor U23131 (N_23131,N_19217,N_17040);
nor U23132 (N_23132,N_16431,N_17315);
and U23133 (N_23133,N_17481,N_12392);
xor U23134 (N_23134,N_13960,N_14698);
or U23135 (N_23135,N_12331,N_14383);
xnor U23136 (N_23136,N_10552,N_17046);
or U23137 (N_23137,N_17195,N_12728);
nand U23138 (N_23138,N_17052,N_14454);
nor U23139 (N_23139,N_13012,N_14284);
nand U23140 (N_23140,N_14825,N_15043);
and U23141 (N_23141,N_17747,N_13330);
and U23142 (N_23142,N_18414,N_12935);
or U23143 (N_23143,N_16104,N_19375);
or U23144 (N_23144,N_13839,N_18034);
nor U23145 (N_23145,N_10816,N_14182);
nor U23146 (N_23146,N_19329,N_13584);
and U23147 (N_23147,N_16980,N_12738);
nor U23148 (N_23148,N_11781,N_14517);
or U23149 (N_23149,N_10974,N_14283);
or U23150 (N_23150,N_13265,N_11124);
or U23151 (N_23151,N_12465,N_13918);
nand U23152 (N_23152,N_11860,N_11478);
nor U23153 (N_23153,N_16934,N_17896);
or U23154 (N_23154,N_16338,N_16999);
nand U23155 (N_23155,N_12412,N_18021);
and U23156 (N_23156,N_13316,N_18192);
and U23157 (N_23157,N_18300,N_17114);
xor U23158 (N_23158,N_11878,N_18566);
xor U23159 (N_23159,N_12419,N_14426);
nor U23160 (N_23160,N_11754,N_17889);
and U23161 (N_23161,N_16952,N_16074);
nand U23162 (N_23162,N_11714,N_13473);
and U23163 (N_23163,N_11695,N_12054);
or U23164 (N_23164,N_13890,N_15970);
nor U23165 (N_23165,N_14875,N_11990);
nand U23166 (N_23166,N_12602,N_17706);
or U23167 (N_23167,N_11971,N_17823);
and U23168 (N_23168,N_18422,N_13504);
xnor U23169 (N_23169,N_13371,N_12736);
nor U23170 (N_23170,N_17179,N_19062);
nor U23171 (N_23171,N_14362,N_15479);
xnor U23172 (N_23172,N_17980,N_13990);
and U23173 (N_23173,N_13740,N_13430);
or U23174 (N_23174,N_19993,N_15436);
or U23175 (N_23175,N_10195,N_16169);
nor U23176 (N_23176,N_13963,N_18121);
nor U23177 (N_23177,N_13362,N_18629);
xor U23178 (N_23178,N_15923,N_12106);
xor U23179 (N_23179,N_17230,N_11820);
or U23180 (N_23180,N_14391,N_13721);
xnor U23181 (N_23181,N_12461,N_18026);
nor U23182 (N_23182,N_13283,N_12554);
nand U23183 (N_23183,N_18063,N_12268);
or U23184 (N_23184,N_12417,N_10233);
and U23185 (N_23185,N_12490,N_18395);
or U23186 (N_23186,N_10828,N_11865);
nand U23187 (N_23187,N_19204,N_15267);
and U23188 (N_23188,N_17348,N_18689);
or U23189 (N_23189,N_15776,N_17987);
nand U23190 (N_23190,N_16463,N_16140);
xor U23191 (N_23191,N_19061,N_17088);
or U23192 (N_23192,N_18705,N_16954);
or U23193 (N_23193,N_16508,N_11600);
nor U23194 (N_23194,N_11296,N_15566);
nand U23195 (N_23195,N_14540,N_10538);
nor U23196 (N_23196,N_19459,N_17765);
and U23197 (N_23197,N_18712,N_19396);
and U23198 (N_23198,N_13418,N_10711);
or U23199 (N_23199,N_18217,N_19410);
xnor U23200 (N_23200,N_17768,N_10078);
and U23201 (N_23201,N_18341,N_10465);
nand U23202 (N_23202,N_19417,N_18680);
nor U23203 (N_23203,N_19399,N_19271);
or U23204 (N_23204,N_10234,N_10900);
xnor U23205 (N_23205,N_13829,N_17665);
xnor U23206 (N_23206,N_19631,N_14342);
or U23207 (N_23207,N_17859,N_13073);
or U23208 (N_23208,N_15427,N_10494);
nand U23209 (N_23209,N_16994,N_14694);
and U23210 (N_23210,N_13319,N_10615);
or U23211 (N_23211,N_11255,N_16407);
nand U23212 (N_23212,N_19561,N_16154);
xor U23213 (N_23213,N_19174,N_19358);
and U23214 (N_23214,N_10485,N_19747);
and U23215 (N_23215,N_17199,N_10306);
nor U23216 (N_23216,N_15221,N_14751);
and U23217 (N_23217,N_17643,N_15971);
nand U23218 (N_23218,N_11175,N_11604);
nand U23219 (N_23219,N_11455,N_12154);
nor U23220 (N_23220,N_16194,N_15943);
and U23221 (N_23221,N_13980,N_18947);
xor U23222 (N_23222,N_15747,N_16608);
or U23223 (N_23223,N_18000,N_15750);
nor U23224 (N_23224,N_12397,N_12285);
and U23225 (N_23225,N_19886,N_19687);
nand U23226 (N_23226,N_17387,N_15179);
xor U23227 (N_23227,N_18396,N_11454);
and U23228 (N_23228,N_10412,N_18749);
and U23229 (N_23229,N_19805,N_13351);
nor U23230 (N_23230,N_16905,N_12983);
nor U23231 (N_23231,N_10159,N_15302);
xor U23232 (N_23232,N_11038,N_19141);
nor U23233 (N_23233,N_14983,N_17237);
or U23234 (N_23234,N_16105,N_13396);
nor U23235 (N_23235,N_17825,N_11742);
and U23236 (N_23236,N_14023,N_12250);
nand U23237 (N_23237,N_13669,N_11777);
nor U23238 (N_23238,N_15509,N_17816);
or U23239 (N_23239,N_12317,N_10671);
or U23240 (N_23240,N_11711,N_17180);
or U23241 (N_23241,N_16924,N_15946);
and U23242 (N_23242,N_15708,N_19516);
or U23243 (N_23243,N_10708,N_16451);
nor U23244 (N_23244,N_17623,N_18342);
nand U23245 (N_23245,N_17705,N_17280);
and U23246 (N_23246,N_18207,N_16181);
or U23247 (N_23247,N_10826,N_13402);
and U23248 (N_23248,N_12762,N_13338);
nand U23249 (N_23249,N_18228,N_11571);
nor U23250 (N_23250,N_12928,N_13255);
and U23251 (N_23251,N_15044,N_16159);
nand U23252 (N_23252,N_16938,N_16405);
nor U23253 (N_23253,N_19249,N_12673);
and U23254 (N_23254,N_10718,N_14250);
nand U23255 (N_23255,N_16060,N_13958);
nand U23256 (N_23256,N_12067,N_14476);
nand U23257 (N_23257,N_13987,N_15668);
and U23258 (N_23258,N_11501,N_14425);
nand U23259 (N_23259,N_10942,N_12813);
nor U23260 (N_23260,N_18314,N_19413);
nand U23261 (N_23261,N_19377,N_12180);
nor U23262 (N_23262,N_16334,N_16561);
xnor U23263 (N_23263,N_10882,N_11399);
and U23264 (N_23264,N_10039,N_10691);
nor U23265 (N_23265,N_15440,N_11929);
or U23266 (N_23266,N_16961,N_16008);
and U23267 (N_23267,N_16406,N_16082);
nor U23268 (N_23268,N_17301,N_19930);
nand U23269 (N_23269,N_16910,N_11102);
or U23270 (N_23270,N_19511,N_10400);
nor U23271 (N_23271,N_19598,N_11117);
or U23272 (N_23272,N_16631,N_15679);
nand U23273 (N_23273,N_14552,N_18969);
nand U23274 (N_23274,N_18221,N_11449);
nand U23275 (N_23275,N_11290,N_17278);
nand U23276 (N_23276,N_13750,N_17543);
or U23277 (N_23277,N_17177,N_17251);
nand U23278 (N_23278,N_10996,N_19723);
or U23279 (N_23279,N_14638,N_11525);
nand U23280 (N_23280,N_12642,N_10427);
or U23281 (N_23281,N_13471,N_16403);
nor U23282 (N_23282,N_12881,N_16825);
or U23283 (N_23283,N_11266,N_18995);
nor U23284 (N_23284,N_19102,N_19085);
nand U23285 (N_23285,N_12029,N_18415);
xor U23286 (N_23286,N_17670,N_12324);
or U23287 (N_23287,N_19338,N_13211);
nor U23288 (N_23288,N_12725,N_12192);
xor U23289 (N_23289,N_15871,N_19534);
nand U23290 (N_23290,N_10028,N_14772);
xnor U23291 (N_23291,N_14942,N_15313);
or U23292 (N_23292,N_18580,N_14123);
or U23293 (N_23293,N_12103,N_18441);
xor U23294 (N_23294,N_15813,N_14332);
nor U23295 (N_23295,N_10891,N_17436);
and U23296 (N_23296,N_10636,N_10796);
nand U23297 (N_23297,N_12976,N_18499);
or U23298 (N_23298,N_13196,N_17076);
xor U23299 (N_23299,N_17071,N_11785);
or U23300 (N_23300,N_16193,N_19650);
and U23301 (N_23301,N_11870,N_18675);
xnor U23302 (N_23302,N_17156,N_11721);
or U23303 (N_23303,N_15653,N_14624);
nand U23304 (N_23304,N_13134,N_16958);
xnor U23305 (N_23305,N_14779,N_15751);
or U23306 (N_23306,N_16572,N_18951);
nor U23307 (N_23307,N_14841,N_10725);
or U23308 (N_23308,N_16674,N_15769);
and U23309 (N_23309,N_14174,N_10270);
nand U23310 (N_23310,N_18668,N_12782);
nand U23311 (N_23311,N_10330,N_15366);
nand U23312 (N_23312,N_18692,N_14136);
nor U23313 (N_23313,N_11492,N_12955);
nand U23314 (N_23314,N_16844,N_13408);
nand U23315 (N_23315,N_11086,N_11084);
or U23316 (N_23316,N_12564,N_10293);
and U23317 (N_23317,N_17207,N_15310);
nand U23318 (N_23318,N_12235,N_11201);
nand U23319 (N_23319,N_11273,N_10933);
or U23320 (N_23320,N_13083,N_19832);
nand U23321 (N_23321,N_18409,N_17417);
nand U23322 (N_23322,N_17920,N_16683);
and U23323 (N_23323,N_12708,N_10101);
nand U23324 (N_23324,N_19789,N_14629);
and U23325 (N_23325,N_13167,N_18304);
nor U23326 (N_23326,N_12030,N_19068);
and U23327 (N_23327,N_15033,N_10989);
nand U23328 (N_23328,N_16880,N_12582);
nor U23329 (N_23329,N_11517,N_18361);
and U23330 (N_23330,N_18769,N_19460);
and U23331 (N_23331,N_10155,N_19852);
and U23332 (N_23332,N_11369,N_17959);
nand U23333 (N_23333,N_14285,N_12894);
or U23334 (N_23334,N_14987,N_11592);
nand U23335 (N_23335,N_17082,N_11327);
and U23336 (N_23336,N_19129,N_17079);
nor U23337 (N_23337,N_15154,N_16006);
or U23338 (N_23338,N_15041,N_14166);
or U23339 (N_23339,N_19640,N_11196);
or U23340 (N_23340,N_19135,N_12581);
nor U23341 (N_23341,N_17994,N_16048);
nor U23342 (N_23342,N_18908,N_19494);
nand U23343 (N_23343,N_16491,N_16223);
nand U23344 (N_23344,N_10011,N_17565);
and U23345 (N_23345,N_19435,N_15694);
and U23346 (N_23346,N_18082,N_14146);
or U23347 (N_23347,N_12542,N_13179);
nand U23348 (N_23348,N_12421,N_16116);
or U23349 (N_23349,N_19543,N_13214);
or U23350 (N_23350,N_17858,N_18551);
or U23351 (N_23351,N_16286,N_17380);
and U23352 (N_23352,N_19642,N_10561);
nand U23353 (N_23353,N_11068,N_17327);
nor U23354 (N_23354,N_11616,N_11520);
nand U23355 (N_23355,N_13041,N_15007);
nor U23356 (N_23356,N_14693,N_19510);
or U23357 (N_23357,N_12083,N_16955);
nor U23358 (N_23358,N_19830,N_14237);
nor U23359 (N_23359,N_18113,N_12014);
xor U23360 (N_23360,N_18572,N_15020);
nand U23361 (N_23361,N_18805,N_10612);
nor U23362 (N_23362,N_16774,N_12340);
nor U23363 (N_23363,N_18670,N_18032);
xor U23364 (N_23364,N_15900,N_16002);
and U23365 (N_23365,N_10010,N_13133);
and U23366 (N_23366,N_17184,N_15244);
or U23367 (N_23367,N_10269,N_14151);
and U23368 (N_23368,N_11579,N_18853);
nor U23369 (N_23369,N_16195,N_12814);
nand U23370 (N_23370,N_11965,N_16916);
nor U23371 (N_23371,N_10579,N_18907);
or U23372 (N_23372,N_19920,N_13651);
nand U23373 (N_23373,N_15546,N_15501);
and U23374 (N_23374,N_12565,N_17373);
nor U23375 (N_23375,N_17425,N_17366);
nor U23376 (N_23376,N_16381,N_13849);
or U23377 (N_23377,N_11146,N_19583);
nor U23378 (N_23378,N_16156,N_13573);
nand U23379 (N_23379,N_11379,N_10106);
or U23380 (N_23380,N_19104,N_12876);
xor U23381 (N_23381,N_13753,N_16663);
nand U23382 (N_23382,N_17562,N_14011);
nor U23383 (N_23383,N_15874,N_15833);
or U23384 (N_23384,N_19308,N_19369);
nor U23385 (N_23385,N_11745,N_14666);
nor U23386 (N_23386,N_11106,N_14770);
and U23387 (N_23387,N_17974,N_12832);
nand U23388 (N_23388,N_14374,N_19007);
xor U23389 (N_23389,N_13230,N_19525);
xnor U23390 (N_23390,N_16893,N_16174);
or U23391 (N_23391,N_19900,N_12436);
nor U23392 (N_23392,N_10100,N_18136);
or U23393 (N_23393,N_18952,N_12575);
and U23394 (N_23394,N_16744,N_19880);
or U23395 (N_23395,N_15460,N_12508);
and U23396 (N_23396,N_19995,N_16260);
and U23397 (N_23397,N_19528,N_12504);
or U23398 (N_23398,N_18901,N_15162);
and U23399 (N_23399,N_14685,N_11390);
nor U23400 (N_23400,N_14774,N_16241);
and U23401 (N_23401,N_16320,N_12305);
or U23402 (N_23402,N_10063,N_10026);
and U23403 (N_23403,N_18239,N_15339);
nor U23404 (N_23404,N_15911,N_13243);
nand U23405 (N_23405,N_19517,N_11853);
nand U23406 (N_23406,N_12675,N_17267);
or U23407 (N_23407,N_19221,N_10912);
and U23408 (N_23408,N_18485,N_11391);
or U23409 (N_23409,N_19121,N_19563);
nand U23410 (N_23410,N_13985,N_10174);
nor U23411 (N_23411,N_14413,N_13278);
nand U23412 (N_23412,N_14788,N_10034);
nor U23413 (N_23413,N_14643,N_17733);
and U23414 (N_23414,N_13766,N_12220);
nor U23415 (N_23415,N_18790,N_12151);
or U23416 (N_23416,N_11383,N_16449);
or U23417 (N_23417,N_18847,N_12379);
nor U23418 (N_23418,N_17585,N_15650);
nand U23419 (N_23419,N_16545,N_17666);
xor U23420 (N_23420,N_13503,N_17487);
or U23421 (N_23421,N_12866,N_14719);
and U23422 (N_23422,N_10634,N_12376);
or U23423 (N_23423,N_13681,N_16501);
nor U23424 (N_23424,N_13921,N_10885);
nor U23425 (N_23425,N_18527,N_15579);
nor U23426 (N_23426,N_15115,N_17226);
or U23427 (N_23427,N_16340,N_17247);
nand U23428 (N_23428,N_10976,N_13374);
and U23429 (N_23429,N_10109,N_14838);
or U23430 (N_23430,N_12031,N_10559);
or U23431 (N_23431,N_19123,N_16214);
or U23432 (N_23432,N_19554,N_13172);
xor U23433 (N_23433,N_11917,N_15035);
and U23434 (N_23434,N_16879,N_13357);
xor U23435 (N_23435,N_16204,N_13554);
and U23436 (N_23436,N_16287,N_19825);
or U23437 (N_23437,N_19610,N_12899);
and U23438 (N_23438,N_10618,N_18896);
nor U23439 (N_23439,N_11310,N_16364);
or U23440 (N_23440,N_19070,N_10380);
and U23441 (N_23441,N_17528,N_12806);
nor U23442 (N_23442,N_12537,N_17832);
xnor U23443 (N_23443,N_18530,N_19222);
and U23444 (N_23444,N_18169,N_14233);
nor U23445 (N_23445,N_16642,N_17538);
and U23446 (N_23446,N_14661,N_16721);
and U23447 (N_23447,N_12173,N_10869);
nand U23448 (N_23448,N_14079,N_11160);
xnor U23449 (N_23449,N_18468,N_17978);
and U23450 (N_23450,N_10966,N_19962);
or U23451 (N_23451,N_17397,N_16509);
nand U23452 (N_23452,N_15156,N_13541);
and U23453 (N_23453,N_13258,N_12055);
nand U23454 (N_23454,N_19253,N_15810);
or U23455 (N_23455,N_17785,N_14528);
nand U23456 (N_23456,N_17070,N_16513);
nand U23457 (N_23457,N_14960,N_17897);
or U23458 (N_23458,N_19258,N_12780);
and U23459 (N_23459,N_10142,N_10324);
nand U23460 (N_23460,N_12615,N_18278);
and U23461 (N_23461,N_18245,N_18691);
xnor U23462 (N_23462,N_14249,N_16516);
nor U23463 (N_23463,N_16294,N_11110);
and U23464 (N_23464,N_19577,N_12799);
nor U23465 (N_23465,N_16529,N_19212);
and U23466 (N_23466,N_14511,N_14721);
xor U23467 (N_23467,N_10337,N_13581);
nand U23468 (N_23468,N_14437,N_15954);
nor U23469 (N_23469,N_13929,N_12068);
nand U23470 (N_23470,N_12833,N_14973);
and U23471 (N_23471,N_16621,N_14464);
and U23472 (N_23472,N_14824,N_12856);
nand U23473 (N_23473,N_12667,N_15429);
nand U23474 (N_23474,N_18211,N_14479);
or U23475 (N_23475,N_16198,N_11277);
and U23476 (N_23476,N_18110,N_13136);
nand U23477 (N_23477,N_10795,N_18685);
or U23478 (N_23478,N_15601,N_12964);
xnor U23479 (N_23479,N_12108,N_15483);
nor U23480 (N_23480,N_11613,N_10993);
nand U23481 (N_23481,N_15176,N_16716);
or U23482 (N_23482,N_16285,N_16601);
nor U23483 (N_23483,N_11848,N_12360);
and U23484 (N_23484,N_14258,N_12074);
and U23485 (N_23485,N_14716,N_18720);
and U23486 (N_23486,N_10783,N_19924);
nand U23487 (N_23487,N_12536,N_18225);
or U23488 (N_23488,N_11410,N_10182);
and U23489 (N_23489,N_18483,N_18765);
and U23490 (N_23490,N_17560,N_17599);
or U23491 (N_23491,N_16819,N_18172);
and U23492 (N_23492,N_11191,N_18719);
xor U23493 (N_23493,N_12717,N_19989);
and U23494 (N_23494,N_12391,N_15962);
nor U23495 (N_23495,N_10082,N_19521);
nand U23496 (N_23496,N_16172,N_11216);
and U23497 (N_23497,N_16386,N_12992);
or U23498 (N_23498,N_19476,N_15907);
or U23499 (N_23499,N_13490,N_19787);
nand U23500 (N_23500,N_19289,N_18542);
or U23501 (N_23501,N_19679,N_17435);
xor U23502 (N_23502,N_14309,N_16472);
nand U23503 (N_23503,N_13967,N_18243);
nand U23504 (N_23504,N_15837,N_10221);
and U23505 (N_23505,N_11605,N_13161);
nand U23506 (N_23506,N_19340,N_10893);
and U23507 (N_23507,N_15166,N_11996);
and U23508 (N_23508,N_11894,N_15387);
nand U23509 (N_23509,N_17119,N_15742);
and U23510 (N_23510,N_10833,N_13576);
and U23511 (N_23511,N_12053,N_18134);
nor U23512 (N_23512,N_19079,N_16811);
xor U23513 (N_23513,N_17089,N_15945);
and U23514 (N_23514,N_10406,N_18020);
and U23515 (N_23515,N_19425,N_17474);
nand U23516 (N_23516,N_14345,N_10454);
nand U23517 (N_23517,N_16023,N_19766);
xor U23518 (N_23518,N_18856,N_14626);
nor U23519 (N_23519,N_16517,N_11645);
nand U23520 (N_23520,N_18823,N_15692);
or U23521 (N_23521,N_13592,N_15430);
and U23522 (N_23522,N_11956,N_15739);
and U23523 (N_23523,N_15880,N_12578);
nand U23524 (N_23524,N_18306,N_15576);
and U23525 (N_23525,N_15985,N_19058);
nand U23526 (N_23526,N_16891,N_18779);
or U23527 (N_23527,N_17115,N_19706);
or U23528 (N_23528,N_10811,N_12307);
nand U23529 (N_23529,N_11887,N_18525);
and U23530 (N_23530,N_16665,N_17935);
nand U23531 (N_23531,N_19526,N_13756);
and U23532 (N_23532,N_13170,N_17922);
nor U23533 (N_23533,N_17414,N_17902);
nor U23534 (N_23534,N_11049,N_14313);
nor U23535 (N_23535,N_17428,N_12511);
nor U23536 (N_23536,N_11464,N_16391);
nand U23537 (N_23537,N_17407,N_15214);
nand U23538 (N_23538,N_17850,N_17294);
and U23539 (N_23539,N_17145,N_18815);
nand U23540 (N_23540,N_17760,N_12864);
or U23541 (N_23541,N_19817,N_18863);
or U23542 (N_23542,N_17506,N_19054);
nor U23543 (N_23543,N_10213,N_15388);
and U23544 (N_23544,N_13328,N_19224);
nand U23545 (N_23545,N_13401,N_10759);
and U23546 (N_23546,N_15608,N_16035);
and U23547 (N_23547,N_10625,N_18054);
nand U23548 (N_23548,N_14563,N_13090);
or U23549 (N_23549,N_15150,N_16087);
nor U23550 (N_23550,N_13345,N_12351);
or U23551 (N_23551,N_14216,N_18866);
and U23552 (N_23552,N_13069,N_15929);
or U23553 (N_23553,N_18579,N_10491);
or U23554 (N_23554,N_16669,N_12219);
and U23555 (N_23555,N_12549,N_14331);
and U23556 (N_23556,N_12088,N_12316);
or U23557 (N_23557,N_16313,N_15372);
nand U23558 (N_23558,N_13472,N_18541);
xor U23559 (N_23559,N_12328,N_14315);
nand U23560 (N_23560,N_13112,N_12641);
nor U23561 (N_23561,N_18816,N_15898);
nor U23562 (N_23562,N_11988,N_19838);
nand U23563 (N_23563,N_10920,N_15910);
nand U23564 (N_23564,N_15839,N_10232);
and U23565 (N_23565,N_16852,N_13615);
nand U23566 (N_23566,N_12533,N_14512);
and U23567 (N_23567,N_17792,N_17212);
nor U23568 (N_23568,N_16890,N_15444);
nand U23569 (N_23569,N_14815,N_15534);
nand U23570 (N_23570,N_13569,N_14649);
nor U23571 (N_23571,N_13600,N_19975);
or U23572 (N_23572,N_15752,N_16976);
and U23573 (N_23573,N_14576,N_18914);
or U23574 (N_23574,N_19862,N_13957);
and U23575 (N_23575,N_16845,N_18622);
and U23576 (N_23576,N_12185,N_13182);
nand U23577 (N_23577,N_11421,N_11230);
xnor U23578 (N_23578,N_14538,N_12124);
and U23579 (N_23579,N_12275,N_18003);
nand U23580 (N_23580,N_13779,N_19949);
nand U23581 (N_23581,N_11222,N_13774);
nand U23582 (N_23582,N_14543,N_19163);
nor U23583 (N_23583,N_17260,N_10512);
xor U23584 (N_23584,N_10075,N_10294);
or U23585 (N_23585,N_11833,N_12953);
nand U23586 (N_23586,N_15172,N_19575);
nand U23587 (N_23587,N_18726,N_18594);
and U23588 (N_23588,N_10848,N_15396);
and U23589 (N_23589,N_12241,N_11093);
nand U23590 (N_23590,N_18186,N_12914);
nor U23591 (N_23591,N_18331,N_15899);
nor U23592 (N_23592,N_15799,N_18500);
and U23593 (N_23593,N_10729,N_17488);
and U23594 (N_23594,N_12278,N_10655);
nand U23595 (N_23595,N_13876,N_14159);
or U23596 (N_23596,N_13974,N_17610);
and U23597 (N_23597,N_19829,N_15711);
or U23598 (N_23598,N_16271,N_18980);
nor U23599 (N_23599,N_11435,N_19152);
or U23600 (N_23600,N_11211,N_13889);
nor U23601 (N_23601,N_16422,N_13113);
or U23602 (N_23602,N_13048,N_10509);
or U23603 (N_23603,N_12644,N_13164);
nand U23604 (N_23604,N_19471,N_18955);
xor U23605 (N_23605,N_16778,N_13392);
and U23606 (N_23606,N_16178,N_16047);
nor U23607 (N_23607,N_17358,N_12141);
nand U23608 (N_23608,N_11112,N_18528);
and U23609 (N_23609,N_13666,N_17352);
or U23610 (N_23610,N_18888,N_17477);
or U23611 (N_23611,N_12516,N_14042);
or U23612 (N_23612,N_14222,N_10281);
or U23613 (N_23613,N_12979,N_11159);
or U23614 (N_23614,N_10935,N_14683);
nor U23615 (N_23615,N_18053,N_11029);
and U23616 (N_23616,N_10069,N_14548);
or U23617 (N_23617,N_14703,N_13891);
and U23618 (N_23618,N_19161,N_15604);
nor U23619 (N_23619,N_10763,N_14078);
nand U23620 (N_23620,N_13996,N_18944);
or U23621 (N_23621,N_18804,N_16930);
nor U23622 (N_23622,N_15570,N_16904);
nor U23623 (N_23623,N_16139,N_14611);
or U23624 (N_23624,N_19144,N_15277);
nor U23625 (N_23625,N_14753,N_13572);
xor U23626 (N_23626,N_12243,N_19374);
nor U23627 (N_23627,N_15500,N_11827);
nor U23628 (N_23628,N_14936,N_12772);
or U23629 (N_23629,N_19972,N_16205);
or U23630 (N_23630,N_17695,N_15773);
or U23631 (N_23631,N_18317,N_17997);
and U23632 (N_23632,N_14566,N_13682);
and U23633 (N_23633,N_15251,N_19628);
nor U23634 (N_23634,N_16830,N_11406);
xor U23635 (N_23635,N_14201,N_16787);
or U23636 (N_23636,N_14996,N_15229);
and U23637 (N_23637,N_16707,N_13320);
or U23638 (N_23638,N_15610,N_18328);
and U23639 (N_23639,N_18407,N_16809);
nand U23640 (N_23640,N_13823,N_19814);
and U23641 (N_23641,N_10065,N_16697);
nor U23642 (N_23642,N_14544,N_11352);
or U23643 (N_23643,N_16355,N_16167);
nand U23644 (N_23644,N_11344,N_14711);
nor U23645 (N_23645,N_13148,N_16865);
and U23646 (N_23646,N_15778,N_19997);
nor U23647 (N_23647,N_15883,N_11796);
nand U23648 (N_23648,N_13037,N_17758);
or U23649 (N_23649,N_15070,N_13036);
nor U23650 (N_23650,N_19081,N_12865);
xnor U23651 (N_23651,N_15023,N_16859);
or U23652 (N_23652,N_12861,N_18393);
and U23653 (N_23653,N_19677,N_15037);
or U23654 (N_23654,N_13284,N_12247);
and U23655 (N_23655,N_16078,N_14302);
or U23656 (N_23656,N_19293,N_19483);
xor U23657 (N_23657,N_11601,N_11577);
nor U23658 (N_23658,N_10020,N_13154);
nor U23659 (N_23659,N_11107,N_17829);
nor U23660 (N_23660,N_15720,N_18510);
and U23661 (N_23661,N_18780,N_12129);
nor U23662 (N_23662,N_16246,N_19284);
or U23663 (N_23663,N_18868,N_15822);
nand U23664 (N_23664,N_17556,N_16912);
xnor U23665 (N_23665,N_12727,N_19774);
nand U23666 (N_23666,N_10112,N_16414);
nor U23667 (N_23667,N_18602,N_19620);
nand U23668 (N_23668,N_18880,N_13896);
nand U23669 (N_23669,N_11825,N_11684);
nor U23670 (N_23670,N_17383,N_17489);
nand U23671 (N_23671,N_12482,N_12383);
or U23672 (N_23672,N_19066,N_10872);
and U23673 (N_23673,N_11018,N_10956);
and U23674 (N_23674,N_17287,N_11597);
nor U23675 (N_23675,N_16812,N_18957);
or U23676 (N_23676,N_10239,N_11674);
nor U23677 (N_23677,N_13704,N_17984);
xor U23678 (N_23678,N_17851,N_15637);
and U23679 (N_23679,N_14114,N_18109);
nor U23680 (N_23680,N_12868,N_11702);
and U23681 (N_23681,N_19126,N_10752);
nor U23682 (N_23682,N_18919,N_17578);
and U23683 (N_23683,N_13702,N_19570);
nand U23684 (N_23684,N_15731,N_15284);
nor U23685 (N_23685,N_13007,N_11672);
or U23686 (N_23686,N_10225,N_12143);
nor U23687 (N_23687,N_12377,N_17853);
and U23688 (N_23688,N_17929,N_14172);
nand U23689 (N_23689,N_19412,N_12674);
nor U23690 (N_23690,N_10780,N_17583);
nor U23691 (N_23691,N_11763,N_17062);
nand U23692 (N_23692,N_10568,N_15722);
and U23693 (N_23693,N_18022,N_17225);
nand U23694 (N_23694,N_14870,N_15712);
nand U23695 (N_23695,N_14236,N_19384);
and U23696 (N_23696,N_13046,N_14914);
or U23697 (N_23697,N_18937,N_15771);
or U23698 (N_23698,N_17539,N_13571);
and U23699 (N_23699,N_13793,N_19343);
nand U23700 (N_23700,N_10658,N_10908);
nand U23701 (N_23701,N_11964,N_13623);
and U23702 (N_23702,N_19304,N_18410);
nor U23703 (N_23703,N_14590,N_16122);
nand U23704 (N_23704,N_19529,N_16676);
or U23705 (N_23705,N_16807,N_18693);
nor U23706 (N_23706,N_16775,N_17586);
nor U23707 (N_23707,N_15276,N_11215);
xor U23708 (N_23708,N_11581,N_17535);
nand U23709 (N_23709,N_15977,N_11948);
nor U23710 (N_23710,N_11101,N_16596);
or U23711 (N_23711,N_14371,N_10821);
and U23712 (N_23712,N_14349,N_12712);
or U23713 (N_23713,N_12169,N_13548);
nand U23714 (N_23714,N_13325,N_16911);
nor U23715 (N_23715,N_12101,N_13192);
or U23716 (N_23716,N_15054,N_18101);
nand U23717 (N_23717,N_14219,N_18867);
nand U23718 (N_23718,N_18557,N_10031);
nand U23719 (N_23719,N_15714,N_17906);
nand U23720 (N_23720,N_10128,N_17763);
or U23721 (N_23721,N_17613,N_15031);
nand U23722 (N_23722,N_13087,N_19546);
or U23723 (N_23723,N_13403,N_15099);
and U23724 (N_23724,N_16330,N_12716);
nand U23725 (N_23725,N_11419,N_18915);
nor U23726 (N_23726,N_15279,N_10297);
or U23727 (N_23727,N_18555,N_13076);
nor U23728 (N_23728,N_16582,N_12910);
nand U23729 (N_23729,N_11899,N_11741);
or U23730 (N_23730,N_14422,N_18741);
nand U23731 (N_23731,N_12501,N_13198);
xnor U23732 (N_23732,N_18355,N_12972);
nand U23733 (N_23733,N_16823,N_16433);
nor U23734 (N_23734,N_15142,N_14038);
nor U23735 (N_23735,N_15458,N_17475);
xnor U23736 (N_23736,N_14812,N_14134);
nor U23737 (N_23737,N_14263,N_18339);
xnor U23738 (N_23738,N_18827,N_17055);
and U23739 (N_23739,N_10137,N_15725);
nor U23740 (N_23740,N_10450,N_14299);
or U23741 (N_23741,N_12764,N_19382);
and U23742 (N_23742,N_18011,N_14522);
xor U23743 (N_23743,N_19731,N_14750);
or U23744 (N_23744,N_13045,N_14524);
nand U23745 (N_23745,N_12423,N_16846);
and U23746 (N_23746,N_19393,N_16432);
nand U23747 (N_23747,N_17072,N_19039);
or U23748 (N_23748,N_11051,N_16456);
or U23749 (N_23749,N_12594,N_13915);
and U23750 (N_23750,N_19322,N_15457);
nor U23751 (N_23751,N_15847,N_11563);
and U23752 (N_23752,N_15814,N_12130);
nor U23753 (N_23753,N_11434,N_13943);
nand U23754 (N_23754,N_11704,N_11867);
nor U23755 (N_23755,N_17781,N_14352);
nor U23756 (N_23756,N_11428,N_19093);
nor U23757 (N_23757,N_13722,N_18188);
or U23758 (N_23758,N_13784,N_10823);
nor U23759 (N_23759,N_10095,N_11617);
or U23760 (N_23760,N_12596,N_16335);
xnor U23761 (N_23761,N_16329,N_19441);
and U23762 (N_23762,N_18102,N_16201);
nor U23763 (N_23763,N_17834,N_14243);
nor U23764 (N_23764,N_12370,N_11021);
nand U23765 (N_23765,N_13454,N_13111);
or U23766 (N_23766,N_16390,N_19714);
xnor U23767 (N_23767,N_12380,N_17029);
or U23768 (N_23768,N_16555,N_10402);
and U23769 (N_23769,N_19137,N_13728);
xnor U23770 (N_23770,N_19883,N_14364);
or U23771 (N_23771,N_15362,N_18399);
nand U23772 (N_23772,N_12677,N_10154);
and U23773 (N_23773,N_14526,N_18039);
or U23774 (N_23774,N_16264,N_19769);
nor U23775 (N_23775,N_18435,N_12098);
or U23776 (N_23776,N_19467,N_10633);
nand U23777 (N_23777,N_17738,N_10332);
nor U23778 (N_23778,N_14984,N_16079);
nand U23779 (N_23779,N_15163,N_10943);
nand U23780 (N_23780,N_10312,N_19553);
and U23781 (N_23781,N_11973,N_10779);
nand U23782 (N_23782,N_17905,N_17320);
xnor U23783 (N_23783,N_11430,N_12354);
nand U23784 (N_23784,N_11829,N_18352);
nand U23785 (N_23785,N_13516,N_12763);
nor U23786 (N_23786,N_15565,N_14872);
nor U23787 (N_23787,N_10810,N_19571);
xor U23788 (N_23788,N_10477,N_15340);
or U23789 (N_23789,N_13559,N_18820);
nor U23790 (N_23790,N_13437,N_19028);
or U23791 (N_23791,N_17831,N_19431);
nand U23792 (N_23792,N_15336,N_11491);
and U23793 (N_23793,N_19844,N_11189);
xnor U23794 (N_23794,N_17116,N_16889);
or U23795 (N_23795,N_10336,N_19885);
nand U23796 (N_23796,N_10425,N_13333);
or U23797 (N_23797,N_12730,N_19898);
xor U23798 (N_23798,N_11186,N_11612);
or U23799 (N_23799,N_11063,N_10654);
nor U23800 (N_23800,N_15275,N_17329);
and U23801 (N_23801,N_14314,N_12526);
nand U23802 (N_23802,N_16192,N_11094);
nand U23803 (N_23803,N_11761,N_16043);
or U23804 (N_23804,N_14466,N_11365);
and U23805 (N_23805,N_19076,N_19209);
xnor U23806 (N_23806,N_13030,N_18270);
xnor U23807 (N_23807,N_19300,N_17497);
or U23808 (N_23808,N_14218,N_17324);
nand U23809 (N_23809,N_11242,N_14646);
or U23810 (N_23810,N_18332,N_17282);
and U23811 (N_23811,N_11103,N_12335);
or U23812 (N_23812,N_18508,N_19884);
or U23813 (N_23813,N_19248,N_17836);
or U23814 (N_23814,N_18238,N_17576);
nand U23815 (N_23815,N_15701,N_11806);
xnor U23816 (N_23816,N_13922,N_15355);
nand U23817 (N_23817,N_17032,N_10705);
or U23818 (N_23818,N_19189,N_14539);
nor U23819 (N_23819,N_11471,N_13972);
or U23820 (N_23820,N_11556,N_11490);
nand U23821 (N_23821,N_16908,N_10619);
nand U23822 (N_23822,N_11192,N_16127);
nand U23823 (N_23823,N_19818,N_15129);
nor U23824 (N_23824,N_19925,N_18173);
xor U23825 (N_23825,N_10972,N_10482);
xor U23826 (N_23826,N_19292,N_12719);
xor U23827 (N_23827,N_17394,N_17007);
xnor U23828 (N_23828,N_19239,N_17547);
or U23829 (N_23829,N_15141,N_13352);
or U23830 (N_23830,N_16785,N_11734);
and U23831 (N_23831,N_19717,N_11286);
and U23832 (N_23832,N_17662,N_13066);
xnor U23833 (N_23833,N_11920,N_15128);
nor U23834 (N_23834,N_16570,N_15527);
xnor U23835 (N_23835,N_17203,N_13530);
and U23836 (N_23836,N_10572,N_14545);
nor U23837 (N_23837,N_17240,N_16144);
or U23838 (N_23838,N_12965,N_18067);
or U23839 (N_23839,N_10071,N_10325);
nor U23840 (N_23840,N_11158,N_10676);
and U23841 (N_23841,N_16858,N_15024);
xor U23842 (N_23842,N_18075,N_15132);
nor U23843 (N_23843,N_12226,N_10839);
or U23844 (N_23844,N_16851,N_18257);
and U23845 (N_23845,N_15262,N_16054);
and U23846 (N_23846,N_14266,N_12486);
nor U23847 (N_23847,N_13475,N_15641);
nor U23848 (N_23848,N_11366,N_10551);
nor U23849 (N_23849,N_17798,N_17134);
or U23850 (N_23850,N_14806,N_11144);
or U23851 (N_23851,N_19124,N_19854);
or U23852 (N_23852,N_13431,N_13887);
and U23853 (N_23853,N_19737,N_10868);
or U23854 (N_23854,N_14297,N_11881);
and U23855 (N_23855,N_15187,N_15193);
or U23856 (N_23856,N_16131,N_14210);
nor U23857 (N_23857,N_10819,N_11499);
and U23858 (N_23858,N_19482,N_15617);
or U23859 (N_23859,N_11815,N_19117);
xnor U23860 (N_23860,N_19347,N_19247);
and U23861 (N_23861,N_10161,N_13752);
or U23862 (N_23862,N_13813,N_10490);
nand U23863 (N_23863,N_12518,N_14520);
nand U23864 (N_23864,N_10749,N_17133);
nor U23865 (N_23865,N_15379,N_19330);
nor U23866 (N_23866,N_19781,N_13147);
and U23867 (N_23867,N_19318,N_15659);
nor U23868 (N_23868,N_14037,N_17186);
nand U23869 (N_23869,N_11328,N_12147);
and U23870 (N_23870,N_17633,N_12264);
and U23871 (N_23871,N_18166,N_14822);
nand U23872 (N_23872,N_17714,N_10379);
nor U23873 (N_23873,N_18215,N_14622);
or U23874 (N_23874,N_17314,N_12400);
nand U23875 (N_23875,N_12984,N_13621);
and U23876 (N_23876,N_13754,N_14864);
and U23877 (N_23877,N_18371,N_12710);
nand U23878 (N_23878,N_14908,N_12479);
and U23879 (N_23879,N_19872,N_12255);
or U23880 (N_23880,N_18998,N_12783);
or U23881 (N_23881,N_17750,N_17168);
and U23882 (N_23882,N_10116,N_12834);
nand U23883 (N_23883,N_18710,N_18124);
or U23884 (N_23884,N_15992,N_15351);
xnor U23885 (N_23885,N_18911,N_15011);
nor U23886 (N_23886,N_10320,N_16250);
nand U23887 (N_23887,N_12513,N_10899);
and U23888 (N_23888,N_13734,N_18384);
xnor U23889 (N_23889,N_15451,N_16277);
nor U23890 (N_23890,N_17370,N_11085);
or U23891 (N_23891,N_12446,N_16557);
and U23892 (N_23892,N_16350,N_13021);
nor U23893 (N_23893,N_10768,N_16817);
nand U23894 (N_23894,N_12294,N_14001);
or U23895 (N_23895,N_15729,N_16853);
nor U23896 (N_23896,N_12599,N_18585);
nor U23897 (N_23897,N_17214,N_10130);
and U23898 (N_23898,N_11477,N_17659);
nand U23899 (N_23899,N_17571,N_12545);
or U23900 (N_23900,N_18475,N_18050);
and U23901 (N_23901,N_15646,N_16657);
xnor U23902 (N_23902,N_18766,N_14741);
nor U23903 (N_23903,N_10748,N_17131);
nand U23904 (N_23904,N_19493,N_12254);
and U23905 (N_23905,N_10583,N_11647);
nor U23906 (N_23906,N_15558,N_16595);
or U23907 (N_23907,N_13348,N_12263);
and U23908 (N_23908,N_11776,N_19504);
nor U23909 (N_23909,N_13586,N_13971);
and U23910 (N_23910,N_18386,N_16711);
or U23911 (N_23911,N_19001,N_12052);
nor U23912 (N_23912,N_19236,N_16776);
or U23913 (N_23913,N_17802,N_12060);
nand U23914 (N_23914,N_10015,N_19397);
nand U23915 (N_23915,N_12610,N_13751);
nor U23916 (N_23916,N_14178,N_11387);
and U23917 (N_23917,N_10683,N_15257);
or U23918 (N_23918,N_14504,N_11199);
and U23919 (N_23919,N_10166,N_18191);
or U23920 (N_23920,N_10581,N_11202);
and U23921 (N_23921,N_17437,N_13783);
nor U23922 (N_23922,N_11583,N_16906);
or U23923 (N_23923,N_14991,N_13322);
nand U23924 (N_23924,N_12661,N_19703);
nor U23925 (N_23925,N_14303,N_14431);
or U23926 (N_23926,N_18802,N_14767);
and U23927 (N_23927,N_14147,N_18253);
nor U23928 (N_23928,N_15304,N_15105);
or U23929 (N_23929,N_14702,N_10769);
nor U23930 (N_23930,N_13293,N_10017);
nor U23931 (N_23931,N_12345,N_13897);
and U23932 (N_23932,N_17707,N_18725);
and U23933 (N_23933,N_16666,N_13789);
nand U23934 (N_23934,N_12999,N_16554);
nor U23935 (N_23935,N_11621,N_18461);
and U23936 (N_23936,N_19110,N_17059);
and U23937 (N_23937,N_19255,N_17511);
or U23938 (N_23938,N_18786,N_15695);
nor U23939 (N_23939,N_12776,N_12531);
and U23940 (N_23940,N_11322,N_18437);
xnor U23941 (N_23941,N_11270,N_13765);
nor U23942 (N_23942,N_15605,N_11495);
xor U23943 (N_23943,N_16479,N_13237);
or U23944 (N_23944,N_19234,N_18035);
nand U23945 (N_23945,N_16233,N_13582);
nor U23946 (N_23946,N_12087,N_10173);
xor U23947 (N_23947,N_10016,N_15897);
and U23948 (N_23948,N_10470,N_12478);
or U23949 (N_23949,N_13109,N_19633);
nand U23950 (N_23950,N_10343,N_11285);
and U23951 (N_23951,N_17960,N_10104);
and U23952 (N_23952,N_10834,N_13795);
nor U23953 (N_23953,N_19800,N_13804);
or U23954 (N_23954,N_14214,N_10230);
nand U23955 (N_23955,N_17419,N_18913);
nand U23956 (N_23956,N_14031,N_13769);
nor U23957 (N_23957,N_12840,N_15568);
nand U23958 (N_23958,N_12295,N_12605);
nand U23959 (N_23959,N_19887,N_19031);
and U23960 (N_23960,N_11706,N_10525);
or U23961 (N_23961,N_12748,N_12375);
nor U23962 (N_23962,N_12003,N_13281);
or U23963 (N_23963,N_14798,N_17640);
nand U23964 (N_23964,N_17621,N_14154);
or U23965 (N_23965,N_14390,N_11401);
and U23966 (N_23966,N_17213,N_11168);
xor U23967 (N_23967,N_11181,N_14148);
and U23968 (N_23968,N_10849,N_10580);
nand U23969 (N_23969,N_17482,N_11908);
nor U23970 (N_23970,N_18848,N_17866);
or U23971 (N_23971,N_19149,N_12897);
nor U23972 (N_23972,N_12580,N_18996);
and U23973 (N_23973,N_12755,N_18979);
nor U23974 (N_23974,N_16268,N_15234);
and U23975 (N_23975,N_16321,N_13314);
and U23976 (N_23976,N_18452,N_14410);
or U23977 (N_23977,N_19519,N_12396);
and U23978 (N_23978,N_11323,N_18160);
nor U23979 (N_23979,N_12378,N_12001);
nand U23980 (N_23980,N_19229,N_18137);
nor U23981 (N_23981,N_11655,N_12825);
nor U23982 (N_23982,N_12995,N_18716);
nand U23983 (N_23983,N_19547,N_18379);
nor U23984 (N_23984,N_14244,N_11808);
xnor U23985 (N_23985,N_10830,N_12569);
or U23986 (N_23986,N_15089,N_11716);
nand U23987 (N_23987,N_13102,N_16050);
nand U23988 (N_23988,N_10635,N_16598);
and U23989 (N_23989,N_14878,N_14723);
nor U23990 (N_23990,N_13588,N_19756);
xor U23991 (N_23991,N_13622,N_18953);
or U23992 (N_23992,N_12958,N_15389);
nand U23993 (N_23993,N_11559,N_12216);
nor U23994 (N_23994,N_16232,N_10303);
and U23995 (N_23995,N_11521,N_19604);
nor U23996 (N_23996,N_19646,N_10587);
nand U23997 (N_23997,N_10648,N_13869);
nor U23998 (N_23998,N_19605,N_11119);
and U23999 (N_23999,N_10515,N_18203);
and U24000 (N_24000,N_10013,N_10132);
and U24001 (N_24001,N_10621,N_17723);
and U24002 (N_24002,N_19987,N_11736);
nand U24003 (N_24003,N_15058,N_10597);
and U24004 (N_24004,N_15930,N_11729);
nand U24005 (N_24005,N_17146,N_19690);
nand U24006 (N_24006,N_18047,N_13184);
xor U24007 (N_24007,N_13805,N_10263);
or U24008 (N_24008,N_12827,N_19046);
and U24009 (N_24009,N_19932,N_17382);
nand U24010 (N_24010,N_17163,N_13979);
nand U24011 (N_24011,N_12739,N_14642);
and U24012 (N_24012,N_17051,N_17822);
or U24013 (N_24013,N_13168,N_15709);
or U24014 (N_24014,N_11730,N_19864);
nor U24015 (N_24015,N_14621,N_12131);
or U24016 (N_24016,N_16039,N_18259);
nand U24017 (N_24017,N_12844,N_10411);
nor U24018 (N_24018,N_13156,N_17077);
xor U24019 (N_24019,N_10955,N_11972);
nand U24020 (N_24020,N_12847,N_17377);
and U24021 (N_24021,N_18334,N_19807);
xor U24022 (N_24022,N_10960,N_18715);
nand U24023 (N_24023,N_17132,N_14489);
and U24024 (N_24024,N_16069,N_18645);
xnor U24025 (N_24025,N_14859,N_19780);
and U24026 (N_24026,N_11584,N_15413);
nor U24027 (N_24027,N_19439,N_10408);
nand U24028 (N_24028,N_13797,N_16945);
nor U24029 (N_24029,N_18165,N_19597);
nor U24030 (N_24030,N_11685,N_14910);
nor U24031 (N_24031,N_14759,N_10596);
and U24032 (N_24032,N_13206,N_10541);
or U24033 (N_24033,N_15952,N_11446);
and U24034 (N_24034,N_13031,N_19301);
or U24035 (N_24035,N_12849,N_19346);
or U24036 (N_24036,N_10516,N_18281);
nor U24037 (N_24037,N_14317,N_13952);
and U24038 (N_24038,N_18421,N_17141);
nand U24039 (N_24039,N_16423,N_17912);
xor U24040 (N_24040,N_16175,N_15233);
nand U24041 (N_24041,N_19017,N_14720);
nand U24042 (N_24042,N_15784,N_19490);
and U24043 (N_24043,N_17563,N_19763);
and U24044 (N_24044,N_15749,N_16558);
xor U24045 (N_24045,N_14865,N_17843);
and U24046 (N_24046,N_19160,N_14883);
nor U24047 (N_24047,N_16063,N_14440);
and U24048 (N_24048,N_14570,N_10144);
nor U24049 (N_24049,N_14880,N_16599);
or U24050 (N_24050,N_18584,N_16630);
and U24051 (N_24051,N_10845,N_19701);
and U24052 (N_24052,N_13078,N_17074);
nand U24053 (N_24053,N_16996,N_13304);
nor U24054 (N_24054,N_11547,N_14668);
xnor U24055 (N_24055,N_16656,N_12588);
nand U24056 (N_24056,N_10497,N_15872);
or U24057 (N_24057,N_16299,N_10342);
and U24058 (N_24058,N_11841,N_16440);
or U24059 (N_24059,N_12059,N_10915);
nand U24060 (N_24060,N_10820,N_15808);
nor U24061 (N_24061,N_17044,N_12654);
or U24062 (N_24062,N_10746,N_18445);
or U24063 (N_24063,N_11319,N_15835);
nor U24064 (N_24064,N_14943,N_11856);
and U24065 (N_24065,N_19206,N_13872);
nand U24066 (N_24066,N_13052,N_10936);
nor U24067 (N_24067,N_16618,N_17193);
and U24068 (N_24068,N_12963,N_15990);
or U24069 (N_24069,N_10453,N_11767);
or U24070 (N_24070,N_17869,N_14275);
or U24071 (N_24071,N_14818,N_18887);
nor U24072 (N_24072,N_18798,N_19151);
xnor U24073 (N_24073,N_16282,N_12713);
and U24074 (N_24074,N_18037,N_11173);
or U24075 (N_24075,N_12288,N_15528);
nor U24076 (N_24076,N_18430,N_13852);
and U24077 (N_24077,N_10286,N_12186);
nand U24078 (N_24078,N_13465,N_16949);
xnor U24079 (N_24079,N_19674,N_11444);
and U24080 (N_24080,N_13653,N_16898);
nand U24081 (N_24081,N_11938,N_16638);
xnor U24082 (N_24082,N_12028,N_18656);
xnor U24083 (N_24083,N_10631,N_13703);
nor U24084 (N_24084,N_15498,N_12507);
or U24085 (N_24085,N_13661,N_11460);
or U24086 (N_24086,N_14862,N_10488);
and U24087 (N_24087,N_19034,N_18503);
and U24088 (N_24088,N_15683,N_12327);
xor U24089 (N_24089,N_17022,N_16117);
or U24090 (N_24090,N_15486,N_12786);
or U24091 (N_24091,N_17390,N_15876);
nor U24092 (N_24092,N_15459,N_19360);
nand U24093 (N_24093,N_12408,N_12420);
nor U24094 (N_24094,N_12680,N_19753);
nand U24095 (N_24095,N_19437,N_18184);
xor U24096 (N_24096,N_17641,N_18644);
or U24097 (N_24097,N_13326,N_13664);
or U24098 (N_24098,N_17261,N_13919);
nand U24099 (N_24099,N_16276,N_17045);
nand U24100 (N_24100,N_19243,N_16881);
nor U24101 (N_24101,N_18049,N_16837);
xnor U24102 (N_24102,N_18377,N_16012);
or U24103 (N_24103,N_12426,N_11985);
or U24104 (N_24104,N_11503,N_17837);
nand U24105 (N_24105,N_13994,N_16305);
nand U24106 (N_24106,N_18906,N_19276);
nor U24107 (N_24107,N_14073,N_19513);
and U24108 (N_24108,N_13222,N_16353);
nor U24109 (N_24109,N_19810,N_10720);
xnor U24110 (N_24110,N_12836,N_11852);
nor U24111 (N_24111,N_16344,N_17694);
nor U24112 (N_24112,N_17424,N_14521);
xor U24113 (N_24113,N_12371,N_18018);
nand U24114 (N_24114,N_19446,N_19233);
and U24115 (N_24115,N_16534,N_12225);
and U24116 (N_24116,N_18627,N_19663);
nand U24117 (N_24117,N_11217,N_10529);
or U24118 (N_24118,N_13139,N_19049);
and U24119 (N_24119,N_10930,N_18526);
nor U24120 (N_24120,N_11108,N_19584);
nand U24121 (N_24121,N_19567,N_14443);
nand U24122 (N_24122,N_19241,N_15841);
or U24123 (N_24123,N_15076,N_17901);
nor U24124 (N_24124,N_14776,N_19059);
or U24125 (N_24125,N_17340,N_19406);
and U24126 (N_24126,N_14330,N_16210);
xnor U24127 (N_24127,N_12745,N_12148);
nand U24128 (N_24128,N_16026,N_13942);
xnor U24129 (N_24129,N_10460,N_12815);
xor U24130 (N_24130,N_16580,N_11131);
or U24131 (N_24131,N_15433,N_14813);
or U24132 (N_24132,N_12774,N_19143);
or U24133 (N_24133,N_16661,N_13034);
nand U24134 (N_24134,N_15225,N_15740);
xnor U24135 (N_24135,N_12848,N_14032);
or U24136 (N_24136,N_17323,N_12207);
and U24137 (N_24137,N_16668,N_13009);
and U24138 (N_24138,N_11341,N_10904);
and U24139 (N_24139,N_17362,N_17925);
nand U24140 (N_24140,N_11241,N_19836);
and U24141 (N_24141,N_15888,N_14989);
or U24142 (N_24142,N_11986,N_11640);
nor U24143 (N_24143,N_18177,N_18419);
xor U24144 (N_24144,N_13466,N_13001);
or U24145 (N_24145,N_16546,N_10223);
and U24146 (N_24146,N_16622,N_12643);
nor U24147 (N_24147,N_14885,N_15991);
or U24148 (N_24148,N_12824,N_16510);
nor U24149 (N_24149,N_14692,N_13904);
nand U24150 (N_24150,N_15303,N_19909);
or U24151 (N_24151,N_15306,N_19407);
and U24152 (N_24152,N_12688,N_17890);
and U24153 (N_24153,N_11809,N_13513);
and U24154 (N_24154,N_19033,N_19936);
nor U24155 (N_24155,N_15649,N_13061);
nor U24156 (N_24156,N_11400,N_11629);
nand U24157 (N_24157,N_12466,N_15453);
or U24158 (N_24158,N_11885,N_11512);
or U24159 (N_24159,N_15107,N_19089);
xor U24160 (N_24160,N_11633,N_14293);
nor U24161 (N_24161,N_11656,N_18232);
and U24162 (N_24162,N_19176,N_17457);
xor U24163 (N_24163,N_16818,N_14939);
nor U24164 (N_24164,N_10686,N_18156);
xor U24165 (N_24165,N_17423,N_19427);
nor U24166 (N_24166,N_18356,N_17420);
nor U24167 (N_24167,N_15553,N_13665);
or U24168 (N_24168,N_17642,N_15927);
nor U24169 (N_24169,N_14805,N_16986);
or U24170 (N_24170,N_12566,N_18651);
and U24171 (N_24171,N_12562,N_15120);
nor U24172 (N_24172,N_13276,N_18981);
or U24173 (N_24173,N_13313,N_12167);
or U24174 (N_24174,N_14306,N_12212);
and U24175 (N_24175,N_19244,N_10356);
nor U24176 (N_24176,N_10837,N_11337);
nand U24177 (N_24177,N_19565,N_15830);
or U24178 (N_24178,N_19536,N_12697);
xor U24179 (N_24179,N_17950,N_11968);
and U24180 (N_24180,N_13379,N_11518);
and U24181 (N_24181,N_19508,N_14556);
nor U24182 (N_24182,N_10947,N_19882);
xnor U24183 (N_24183,N_14732,N_12458);
nor U24184 (N_24184,N_15864,N_12669);
xor U24185 (N_24185,N_13060,N_19389);
nor U24186 (N_24186,N_18007,N_17907);
or U24187 (N_24187,N_11412,N_14445);
or U24188 (N_24188,N_11316,N_19942);
nor U24189 (N_24189,N_12277,N_18663);
nand U24190 (N_24190,N_12884,N_12382);
and U24191 (N_24191,N_13834,N_18817);
nand U24192 (N_24192,N_15348,N_10345);
nor U24193 (N_24193,N_12905,N_13208);
or U24194 (N_24194,N_15153,N_15232);
nand U24195 (N_24195,N_12546,N_17005);
or U24196 (N_24196,N_15268,N_16190);
or U24197 (N_24197,N_11451,N_10805);
nor U24198 (N_24198,N_10967,N_11828);
nor U24199 (N_24199,N_10679,N_14952);
and U24200 (N_24200,N_11011,N_16388);
nor U24201 (N_24201,N_14376,N_15357);
xnor U24202 (N_24202,N_18152,N_17886);
and U24203 (N_24203,N_11078,N_19702);
and U24204 (N_24204,N_11271,N_18097);
or U24205 (N_24205,N_18115,N_16973);
nand U24206 (N_24206,N_12057,N_12082);
and U24207 (N_24207,N_17026,N_19297);
and U24208 (N_24208,N_11126,N_17947);
nand U24209 (N_24209,N_19591,N_13026);
nor U24210 (N_24210,N_12425,N_11598);
nor U24211 (N_24211,N_17501,N_10951);
nand U24212 (N_24212,N_19552,N_17812);
or U24213 (N_24213,N_17265,N_10441);
or U24214 (N_24214,N_19252,N_13280);
nor U24215 (N_24215,N_13788,N_14007);
and U24216 (N_24216,N_15678,N_10523);
or U24217 (N_24217,N_13645,N_14235);
xnor U24218 (N_24218,N_10448,N_11187);
xnor U24219 (N_24219,N_19973,N_14618);
nor U24220 (N_24220,N_10398,N_15753);
and U24221 (N_24221,N_11883,N_19422);
or U24222 (N_24222,N_10522,N_11264);
or U24223 (N_24223,N_16731,N_12140);
nand U24224 (N_24224,N_11060,N_11882);
nand U24225 (N_24225,N_14252,N_14070);
nor U24226 (N_24226,N_18294,N_16625);
and U24227 (N_24227,N_12489,N_15004);
or U24228 (N_24228,N_10038,N_10395);
nor U24229 (N_24229,N_12056,N_12269);
or U24230 (N_24230,N_18472,N_18227);
nor U24231 (N_24231,N_18575,N_14120);
xnor U24232 (N_24232,N_13781,N_18106);
nand U24233 (N_24233,N_12975,N_14682);
xnor U24234 (N_24234,N_11801,N_10981);
and U24235 (N_24235,N_17916,N_17169);
or U24236 (N_24236,N_18487,N_18296);
nor U24237 (N_24237,N_17336,N_18357);
and U24238 (N_24238,N_17025,N_14377);
nor U24239 (N_24239,N_12637,N_12788);
nand U24240 (N_24240,N_15001,N_18728);
and U24241 (N_24241,N_13949,N_10892);
and U24242 (N_24242,N_14565,N_10598);
and U24243 (N_24243,N_17508,N_19175);
or U24244 (N_24244,N_14327,N_12742);
nor U24245 (N_24245,N_12265,N_11076);
or U24246 (N_24246,N_10359,N_16183);
and U24247 (N_24247,N_16278,N_18666);
nand U24248 (N_24248,N_14498,N_13676);
and U24249 (N_24249,N_15228,N_14771);
nor U24250 (N_24250,N_12012,N_19130);
and U24251 (N_24251,N_18406,N_18423);
nand U24252 (N_24252,N_10605,N_12163);
nor U24253 (N_24253,N_17605,N_12467);
nor U24254 (N_24254,N_11731,N_10964);
nand U24255 (N_24255,N_16036,N_15287);
and U24256 (N_24256,N_12660,N_14927);
and U24257 (N_24257,N_15333,N_11795);
or U24258 (N_24258,N_16266,N_11555);
xor U24259 (N_24259,N_12496,N_14793);
and U24260 (N_24260,N_19568,N_16348);
nand U24261 (N_24261,N_18928,N_13901);
and U24262 (N_24262,N_15937,N_11847);
and U24263 (N_24263,N_18742,N_17367);
nand U24264 (N_24264,N_18052,N_19576);
nand U24265 (N_24265,N_18904,N_14225);
or U24266 (N_24266,N_15932,N_12485);
and U24267 (N_24267,N_11208,N_12330);
nor U24268 (N_24268,N_14849,N_14628);
or U24269 (N_24269,N_15783,N_10863);
nor U24270 (N_24270,N_14033,N_13749);
nand U24271 (N_24271,N_19738,N_12246);
and U24272 (N_24272,N_17773,N_16804);
nand U24273 (N_24273,N_18878,N_17719);
and U24274 (N_24274,N_14380,N_17361);
nand U24275 (N_24275,N_14742,N_19491);
nor U24276 (N_24276,N_17909,N_12568);
or U24277 (N_24277,N_17868,N_15373);
and U24278 (N_24278,N_13270,N_13519);
and U24279 (N_24279,N_10544,N_10907);
and U24280 (N_24280,N_17452,N_10436);
or U24281 (N_24281,N_17542,N_13081);
xor U24282 (N_24282,N_19709,N_18263);
nand U24283 (N_24283,N_15536,N_15674);
and U24284 (N_24284,N_11513,N_10699);
xnor U24285 (N_24285,N_17318,N_10480);
nand U24286 (N_24286,N_15456,N_19319);
and U24287 (N_24287,N_11568,N_13603);
xor U24288 (N_24288,N_14982,N_13883);
xnor U24289 (N_24289,N_14077,N_13129);
or U24290 (N_24290,N_18731,N_14645);
xor U24291 (N_24291,N_13933,N_10841);
or U24292 (N_24292,N_11470,N_12372);
nor U24293 (N_24293,N_15032,N_13574);
or U24294 (N_24294,N_14749,N_19047);
or U24295 (N_24295,N_10179,N_15545);
and U24296 (N_24296,N_16146,N_13532);
and U24297 (N_24297,N_12543,N_11072);
and U24298 (N_24298,N_10430,N_19708);
or U24299 (N_24299,N_13059,N_17283);
nand U24300 (N_24300,N_17120,N_16619);
nand U24301 (N_24301,N_10317,N_18392);
nand U24302 (N_24302,N_19313,N_14016);
nand U24303 (N_24303,N_14913,N_12808);
nor U24304 (N_24304,N_10707,N_13879);
nor U24305 (N_24305,N_18418,N_11278);
xor U24306 (N_24306,N_16943,N_15314);
xor U24307 (N_24307,N_14510,N_13199);
nand U24308 (N_24308,N_17799,N_10085);
xor U24309 (N_24309,N_17204,N_11575);
xor U24310 (N_24310,N_13417,N_14663);
and U24311 (N_24311,N_14722,N_13619);
nand U24312 (N_24312,N_18929,N_19712);
nor U24313 (N_24313,N_11261,N_13123);
nand U24314 (N_24314,N_19958,N_14030);
or U24315 (N_24315,N_14745,N_13551);
or U24316 (N_24316,N_19473,N_17715);
xnor U24317 (N_24317,N_16081,N_12590);
or U24318 (N_24318,N_18262,N_17941);
nor U24319 (N_24319,N_12231,N_15325);
nor U24320 (N_24320,N_18494,N_10859);
nor U24321 (N_24321,N_18796,N_18556);
nor U24322 (N_24322,N_10322,N_10937);
and U24323 (N_24323,N_14018,N_14729);
nand U24324 (N_24324,N_17751,N_14294);
and U24325 (N_24325,N_16899,N_18247);
nor U24326 (N_24326,N_19275,N_16165);
or U24327 (N_24327,N_17999,N_17416);
nand U24328 (N_24328,N_11664,N_14889);
and U24329 (N_24329,N_14704,N_16306);
or U24330 (N_24330,N_17704,N_12104);
or U24331 (N_24331,N_12457,N_19183);
xnor U24332 (N_24332,N_18783,N_18750);
nand U24333 (N_24333,N_18333,N_14357);
nand U24334 (N_24334,N_10266,N_10856);
nand U24335 (N_24335,N_18486,N_13484);
or U24336 (N_24336,N_16017,N_13257);
and U24337 (N_24337,N_13583,N_11276);
or U24338 (N_24338,N_19762,N_15575);
or U24339 (N_24339,N_11367,N_16735);
or U24340 (N_24340,N_18416,N_19502);
nor U24341 (N_24341,N_12711,N_10365);
xor U24342 (N_24342,N_18433,N_15815);
xor U24343 (N_24343,N_13450,N_13526);
nor U24344 (N_24344,N_18699,N_19980);
nand U24345 (N_24345,N_18945,N_13010);
and U24346 (N_24346,N_14968,N_11909);
nand U24347 (N_24347,N_15200,N_17063);
xnor U24348 (N_24348,N_18405,N_18702);
nor U24349 (N_24349,N_10710,N_13369);
nand U24350 (N_24350,N_18592,N_10403);
or U24351 (N_24351,N_12559,N_18316);
nor U24352 (N_24352,N_10133,N_10289);
or U24353 (N_24353,N_11143,N_14059);
nand U24354 (N_24354,N_13800,N_14438);
or U24355 (N_24355,N_15965,N_15213);
xnor U24356 (N_24356,N_12804,N_17919);
and U24357 (N_24357,N_10853,N_17533);
or U24358 (N_24358,N_16857,N_19280);
nor U24359 (N_24359,N_10110,N_12990);
nor U24360 (N_24360,N_13411,N_17157);
nor U24361 (N_24361,N_19336,N_12611);
nand U24362 (N_24362,N_12359,N_14153);
nor U24363 (N_24363,N_17656,N_15061);
xor U24364 (N_24364,N_13991,N_11505);
and U24365 (N_24365,N_19851,N_17900);
nand U24366 (N_24366,N_17651,N_13638);
or U24367 (N_24367,N_18274,N_19609);
and U24368 (N_24368,N_14650,N_12552);
or U24369 (N_24369,N_18139,N_19398);
or U24370 (N_24370,N_11012,N_13735);
xor U24371 (N_24371,N_13970,N_12778);
xnor U24372 (N_24372,N_14662,N_12430);
and U24373 (N_24373,N_16336,N_18836);
and U24374 (N_24374,N_14525,N_11125);
nor U24375 (N_24375,N_15757,N_14107);
nor U24376 (N_24376,N_17574,N_16417);
and U24377 (N_24377,N_12809,N_11480);
and U24378 (N_24378,N_11225,N_10806);
nand U24379 (N_24379,N_14427,N_19710);
or U24380 (N_24380,N_16415,N_17634);
nor U24381 (N_24381,N_15250,N_16458);
or U24382 (N_24382,N_10389,N_11407);
or U24383 (N_24383,N_13039,N_11864);
and U24384 (N_24384,N_13377,N_16361);
and U24385 (N_24385,N_17995,N_14739);
and U24386 (N_24386,N_16730,N_10990);
xor U24387 (N_24387,N_14215,N_10879);
or U24388 (N_24388,N_18095,N_12040);
xor U24389 (N_24389,N_18873,N_16752);
nand U24390 (N_24390,N_16112,N_10800);
and U24391 (N_24391,N_16779,N_17898);
nand U24392 (N_24392,N_17409,N_10158);
xnor U24393 (N_24393,N_16442,N_18793);
nand U24394 (N_24394,N_18179,N_10056);
nor U24395 (N_24395,N_16607,N_10357);
and U24396 (N_24396,N_12889,N_16134);
or U24397 (N_24397,N_17360,N_18140);
and U24398 (N_24398,N_17210,N_18976);
and U24399 (N_24399,N_10734,N_12311);
and U24400 (N_24400,N_14206,N_16515);
or U24401 (N_24401,N_17138,N_19136);
nor U24402 (N_24402,N_14796,N_19593);
nor U24403 (N_24403,N_14071,N_12790);
and U24404 (N_24404,N_12197,N_16363);
nand U24405 (N_24405,N_17903,N_19666);
or U24406 (N_24406,N_12624,N_19461);
nor U24407 (N_24407,N_19464,N_14132);
nand U24408 (N_24408,N_12009,N_14097);
nor U24409 (N_24409,N_16594,N_14896);
and U24410 (N_24410,N_10694,N_16915);
nor U24411 (N_24411,N_17137,N_12296);
nor U24412 (N_24412,N_19961,N_16658);
or U24413 (N_24413,N_14361,N_17103);
and U24414 (N_24414,N_15840,N_12609);
and U24415 (N_24415,N_10684,N_12528);
or U24416 (N_24416,N_15093,N_17220);
and U24417 (N_24417,N_13830,N_15902);
nand U24418 (N_24418,N_19269,N_11157);
nand U24419 (N_24419,N_11524,N_10121);
nand U24420 (N_24420,N_17927,N_14108);
nor U24421 (N_24421,N_15197,N_13956);
and U24422 (N_24422,N_12850,N_14763);
nor U24423 (N_24423,N_13691,N_15894);
nor U24424 (N_24424,N_15595,N_11338);
and U24425 (N_24425,N_17058,N_14208);
nor U24426 (N_24426,N_14768,N_12301);
or U24427 (N_24427,N_12573,N_16317);
and U24428 (N_24428,N_13025,N_18372);
nor U24429 (N_24429,N_14877,N_12918);
nor U24430 (N_24430,N_19092,N_19813);
nand U24431 (N_24431,N_17517,N_16645);
and U24432 (N_24432,N_13640,N_17548);
and U24433 (N_24433,N_11884,N_16764);
nand U24434 (N_24434,N_17887,N_17279);
nor U24435 (N_24435,N_19667,N_16380);
nand U24436 (N_24436,N_15544,N_15903);
or U24437 (N_24437,N_16715,N_14644);
or U24438 (N_24438,N_19277,N_18558);
xnor U24439 (N_24439,N_19090,N_13657);
xnor U24440 (N_24440,N_19653,N_13282);
nand U24441 (N_24441,N_11161,N_17264);
nand U24442 (N_24442,N_16437,N_15048);
nor U24443 (N_24443,N_17153,N_12107);
and U24444 (N_24444,N_11837,N_19967);
nor U24445 (N_24445,N_17780,N_10983);
xor U24446 (N_24446,N_15635,N_11031);
or U24447 (N_24447,N_19230,N_10985);
and U24448 (N_24448,N_15951,N_14709);
nand U24449 (N_24449,N_13144,N_19544);
nor U24450 (N_24450,N_19636,N_13558);
and U24451 (N_24451,N_13013,N_10439);
or U24452 (N_24452,N_18252,N_10758);
nor U24453 (N_24453,N_17566,N_19994);
or U24454 (N_24454,N_19165,N_13566);
or U24455 (N_24455,N_18267,N_15497);
nand U24456 (N_24456,N_19601,N_19096);
nor U24457 (N_24457,N_16161,N_17622);
and U24458 (N_24458,N_17500,N_16342);
or U24459 (N_24459,N_15242,N_13460);
nor U24460 (N_24460,N_10669,N_19466);
or U24461 (N_24461,N_18858,N_17136);
nand U24462 (N_24462,N_12853,N_13875);
nor U24463 (N_24463,N_18801,N_19848);
nor U24464 (N_24464,N_12510,N_19772);
nor U24465 (N_24465,N_14223,N_16636);
nand U24466 (N_24466,N_13476,N_17603);
or U24467 (N_24467,N_12000,N_15525);
and U24468 (N_24468,N_15331,N_12614);
and U24469 (N_24469,N_16076,N_10878);
and U24470 (N_24470,N_11872,N_17879);
nor U24471 (N_24471,N_13616,N_12877);
nor U24472 (N_24472,N_16259,N_11118);
or U24473 (N_24473,N_17546,N_12759);
or U24474 (N_24474,N_18383,N_10323);
nand U24475 (N_24475,N_13481,N_18543);
or U24476 (N_24476,N_11544,N_16288);
nor U24477 (N_24477,N_18413,N_18235);
and U24478 (N_24478,N_16736,N_13178);
and U24479 (N_24479,N_18920,N_16068);
xor U24480 (N_24480,N_12097,N_17784);
or U24481 (N_24481,N_13831,N_15403);
nand U24482 (N_24482,N_15755,N_16387);
and U24483 (N_24483,N_11025,N_15744);
or U24484 (N_24484,N_15380,N_17328);
nor U24485 (N_24485,N_16862,N_13501);
nand U24486 (N_24486,N_12820,N_17667);
nand U24487 (N_24487,N_13446,N_17813);
or U24488 (N_24488,N_11237,N_13780);
or U24489 (N_24489,N_16319,N_14457);
or U24490 (N_24490,N_19896,N_10611);
nand U24491 (N_24491,N_10613,N_15408);
or U24492 (N_24492,N_19004,N_16946);
nand U24493 (N_24493,N_14797,N_10988);
nor U24494 (N_24494,N_18674,N_14062);
xor U24495 (N_24495,N_15877,N_11074);
xnor U24496 (N_24496,N_14402,N_13423);
nand U24497 (N_24497,N_19214,N_12437);
and U24498 (N_24498,N_16207,N_11639);
and U24499 (N_24499,N_14519,N_14448);
and U24500 (N_24500,N_13986,N_12522);
nor U24501 (N_24501,N_19541,N_13406);
nand U24502 (N_24502,N_17848,N_12631);
xor U24503 (N_24503,N_16480,N_16896);
and U24504 (N_24504,N_11595,N_10331);
nor U24505 (N_24505,N_16826,N_13118);
nand U24506 (N_24506,N_19673,N_15289);
nand U24507 (N_24507,N_13153,N_10404);
nor U24508 (N_24508,N_18046,N_13723);
nand U24509 (N_24509,N_12945,N_10153);
xnor U24510 (N_24510,N_18713,N_19083);
or U24511 (N_24511,N_18326,N_14593);
and U24512 (N_24512,N_16753,N_15448);
nor U24513 (N_24513,N_15051,N_16754);
nor U24514 (N_24514,N_13542,N_17229);
xor U24515 (N_24515,N_18660,N_11896);
nand U24516 (N_24516,N_17795,N_11484);
xnor U24517 (N_24517,N_11975,N_16037);
nand U24518 (N_24518,N_17343,N_11832);
and U24519 (N_24519,N_14450,N_18763);
xnor U24520 (N_24520,N_10927,N_10111);
nor U24521 (N_24521,N_12671,N_14917);
or U24522 (N_24522,N_19799,N_11782);
and U24523 (N_24523,N_11488,N_15482);
or U24524 (N_24524,N_18492,N_16096);
nand U24525 (N_24525,N_14217,N_15278);
nor U24526 (N_24526,N_14231,N_13575);
nand U24527 (N_24527,N_11295,N_10083);
and U24528 (N_24528,N_19647,N_18679);
nor U24529 (N_24529,N_18924,N_15029);
nand U24530 (N_24530,N_15530,N_17910);
and U24531 (N_24531,N_17842,N_14634);
and U24532 (N_24532,N_13853,N_17824);
or U24533 (N_24533,N_18524,N_14195);
xnor U24534 (N_24534,N_11233,N_16459);
nor U24535 (N_24535,N_17924,N_10103);
nand U24536 (N_24536,N_10644,N_10817);
nor U24537 (N_24537,N_18894,N_18272);
or U24538 (N_24538,N_13693,N_14853);
and U24539 (N_24539,N_14162,N_17050);
xor U24540 (N_24540,N_12917,N_12355);
and U24541 (N_24541,N_12585,N_16950);
and U24542 (N_24542,N_15741,N_18434);
or U24543 (N_24543,N_19187,N_18537);
nor U24544 (N_24544,N_19428,N_12213);
xor U24545 (N_24545,N_17363,N_12309);
nor U24546 (N_24546,N_12406,N_19705);
nor U24547 (N_24547,N_11127,N_14106);
nor U24548 (N_24548,N_14665,N_16478);
and U24549 (N_24549,N_10467,N_18824);
nor U24550 (N_24550,N_19440,N_13916);
and U24551 (N_24551,N_13596,N_13315);
nor U24552 (N_24552,N_11539,N_10226);
nand U24553 (N_24553,N_18845,N_15772);
and U24554 (N_24554,N_19231,N_13981);
nor U24555 (N_24555,N_17337,N_18266);
nand U24556 (N_24556,N_19016,N_10677);
nor U24557 (N_24557,N_16384,N_16965);
nand U24558 (N_24558,N_18264,N_16225);
or U24559 (N_24559,N_19497,N_19821);
nor U24560 (N_24560,N_17568,N_11388);
and U24561 (N_24561,N_19195,N_17684);
nand U24562 (N_24562,N_10569,N_14305);
or U24563 (N_24563,N_18550,N_17095);
and U24564 (N_24564,N_13508,N_17668);
nand U24565 (N_24565,N_11687,N_12239);
nor U24566 (N_24566,N_11494,N_19387);
nand U24567 (N_24567,N_18826,N_19220);
nor U24568 (N_24568,N_17441,N_10851);
nor U24569 (N_24569,N_18469,N_14054);
nand U24570 (N_24570,N_16888,N_11910);
nor U24571 (N_24571,N_14635,N_13878);
nor U24572 (N_24572,N_18458,N_19696);
nand U24573 (N_24573,N_10290,N_12970);
nand U24574 (N_24574,N_10413,N_15192);
nor U24575 (N_24575,N_15916,N_14452);
or U24576 (N_24576,N_12454,N_14378);
nor U24577 (N_24577,N_13233,N_10319);
nor U24578 (N_24578,N_15647,N_15185);
and U24579 (N_24579,N_12968,N_13989);
nand U24580 (N_24580,N_12648,N_13297);
nor U24581 (N_24581,N_14881,N_10774);
or U24582 (N_24582,N_10162,N_11660);
nand U24583 (N_24583,N_15834,N_12313);
xnor U24584 (N_24584,N_14241,N_13404);
xor U24585 (N_24585,N_10464,N_14752);
nor U24586 (N_24586,N_10921,N_15661);
xnor U24587 (N_24587,N_13119,N_16892);
nor U24588 (N_24588,N_10277,N_17786);
and U24589 (N_24589,N_16213,N_17998);
and U24590 (N_24590,N_15682,N_16153);
nor U24591 (N_24591,N_16028,N_12019);
nand U24592 (N_24592,N_12702,N_14248);
or U24593 (N_24593,N_17596,N_14269);
nor U24594 (N_24594,N_10087,N_14541);
or U24595 (N_24595,N_11424,N_13948);
or U24596 (N_24596,N_12757,N_12144);
nand U24597 (N_24597,N_13412,N_16808);
or U24598 (N_24598,N_15981,N_15462);
and U24599 (N_24599,N_11033,N_15788);
or U24600 (N_24600,N_16956,N_11361);
nor U24601 (N_24601,N_16586,N_15849);
nor U24602 (N_24602,N_11892,N_17530);
or U24603 (N_24603,N_16827,N_10093);
or U24604 (N_24604,N_10965,N_15964);
nor U24605 (N_24605,N_18480,N_19173);
nand U24606 (N_24606,N_11743,N_15126);
xor U24607 (N_24607,N_13296,N_11542);
nor U24608 (N_24608,N_15953,N_11339);
and U24609 (N_24609,N_13903,N_17149);
xnor U24610 (N_24610,N_12363,N_14760);
nor U24611 (N_24611,N_16836,N_15296);
nor U24612 (N_24612,N_13525,N_11646);
nor U24613 (N_24613,N_15777,N_17308);
nand U24614 (N_24614,N_19040,N_12829);
nor U24615 (N_24615,N_19503,N_16926);
xnor U24616 (N_24616,N_14736,N_18260);
or U24617 (N_24617,N_19257,N_19681);
nand U24618 (N_24618,N_14829,N_19796);
nand U24619 (N_24619,N_10175,N_11466);
nand U24620 (N_24620,N_18229,N_11462);
nand U24621 (N_24621,N_12484,N_10563);
nor U24622 (N_24622,N_17540,N_16991);
xor U24623 (N_24623,N_17809,N_17303);
nand U24624 (N_24624,N_10537,N_14211);
and U24625 (N_24625,N_13388,N_11283);
nor U24626 (N_24626,N_14684,N_16244);
xor U24627 (N_24627,N_12121,N_15066);
xor U24628 (N_24628,N_19337,N_19018);
nor U24629 (N_24629,N_16919,N_12538);
xor U24630 (N_24630,N_11950,N_14467);
nand U24631 (N_24631,N_19794,N_14708);
nand U24632 (N_24632,N_18686,N_19740);
nand U24633 (N_24633,N_16029,N_17860);
and U24634 (N_24634,N_15158,N_14432);
nor U24635 (N_24635,N_15928,N_15865);
or U24636 (N_24636,N_13553,N_12145);
or U24637 (N_24637,N_11744,N_12409);
or U24638 (N_24638,N_14028,N_10220);
xnor U24639 (N_24639,N_13389,N_17973);
and U24640 (N_24640,N_12720,N_15034);
nor U24641 (N_24641,N_18285,N_14002);
or U24642 (N_24642,N_18611,N_12344);
nor U24643 (N_24643,N_18447,N_17412);
and U24644 (N_24644,N_14061,N_17550);
nand U24645 (N_24645,N_14348,N_13598);
or U24646 (N_24646,N_13422,N_19613);
nand U24647 (N_24647,N_13701,N_19868);
xnor U24648 (N_24648,N_18387,N_19834);
xor U24649 (N_24649,N_15356,N_14057);
and U24650 (N_24650,N_17304,N_14458);
and U24651 (N_24651,N_11007,N_14058);
nor U24652 (N_24652,N_14419,N_19847);
or U24653 (N_24653,N_15559,N_14990);
or U24654 (N_24654,N_15038,N_18138);
nand U24655 (N_24655,N_16874,N_18512);
nor U24656 (N_24656,N_11658,N_14370);
xnor U24657 (N_24657,N_19029,N_10755);
nand U24658 (N_24658,N_11871,N_11533);
and U24659 (N_24659,N_16523,N_12183);
or U24660 (N_24660,N_11092,N_18770);
and U24661 (N_24661,N_12592,N_11793);
nor U24662 (N_24662,N_13223,N_19602);
or U24663 (N_24663,N_17731,N_10027);
nor U24664 (N_24664,N_18250,N_14245);
nor U24665 (N_24665,N_11889,N_10114);
and U24666 (N_24666,N_16395,N_18241);
nor U24667 (N_24667,N_12603,N_18151);
xor U24668 (N_24668,N_11842,N_16917);
nand U24669 (N_24669,N_11626,N_13309);
or U24670 (N_24670,N_15003,N_13939);
nand U24671 (N_24671,N_15941,N_16528);
xor U24672 (N_24672,N_14125,N_17931);
nor U24673 (N_24673,N_14310,N_18961);
or U24674 (N_24674,N_11417,N_17569);
nor U24675 (N_24675,N_19273,N_15693);
xnor U24676 (N_24676,N_10051,N_15824);
and U24677 (N_24677,N_13350,N_12793);
and U24678 (N_24678,N_17061,N_11628);
and U24679 (N_24679,N_14890,N_19201);
nand U24680 (N_24680,N_12883,N_10897);
or U24681 (N_24681,N_12634,N_17067);
and U24682 (N_24682,N_17008,N_16346);
xor U24683 (N_24683,N_17057,N_15826);
nand U24684 (N_24684,N_12967,N_16148);
nor U24685 (N_24685,N_14965,N_14384);
nand U24686 (N_24686,N_17728,N_15645);
nand U24687 (N_24687,N_12616,N_19730);
and U24688 (N_24688,N_15523,N_12571);
nor U24689 (N_24689,N_16931,N_17111);
or U24690 (N_24690,N_13428,N_10122);
nor U24691 (N_24691,N_10958,N_15583);
nand U24692 (N_24692,N_19770,N_11898);
or U24693 (N_24693,N_16041,N_19917);
or U24694 (N_24694,N_16455,N_13324);
nor U24695 (N_24695,N_19448,N_18889);
nor U24696 (N_24696,N_12936,N_14808);
xnor U24697 (N_24697,N_14674,N_19166);
or U24698 (N_24698,N_14794,N_15510);
xor U24699 (N_24699,N_17258,N_16356);
or U24700 (N_24700,N_15149,N_12004);
nor U24701 (N_24701,N_18161,N_19595);
or U24702 (N_24702,N_10843,N_12525);
nor U24703 (N_24703,N_19720,N_10315);
nor U24704 (N_24704,N_12589,N_15908);
or U24705 (N_24705,N_17288,N_18746);
and U24706 (N_24706,N_14394,N_11653);
or U24707 (N_24707,N_12199,N_15548);
or U24708 (N_24708,N_19694,N_17545);
nand U24709 (N_24709,N_18501,N_19162);
nor U24710 (N_24710,N_12334,N_18664);
nand U24711 (N_24711,N_18432,N_14343);
and U24712 (N_24712,N_16252,N_10492);
xnor U24713 (N_24713,N_14631,N_18220);
nor U24714 (N_24714,N_17123,N_19750);
xor U24715 (N_24715,N_14387,N_10422);
or U24716 (N_24716,N_11043,N_16358);
or U24717 (N_24717,N_10918,N_14700);
xor U24718 (N_24718,N_14912,N_18451);
nand U24719 (N_24719,N_17421,N_19950);
and U24720 (N_24720,N_19919,N_17444);
nand U24721 (N_24721,N_15305,N_19208);
nor U24722 (N_24722,N_10975,N_16031);
nand U24723 (N_24723,N_11325,N_14630);
nor U24724 (N_24724,N_13227,N_11169);
or U24725 (N_24725,N_13509,N_15188);
nand U24726 (N_24726,N_18048,N_10732);
nand U24727 (N_24727,N_15378,N_16548);
and U24728 (N_24728,N_13720,N_10283);
or U24729 (N_24729,N_16623,N_19965);
nand U24730 (N_24730,N_13819,N_17669);
nand U24731 (N_24731,N_12915,N_19356);
nor U24732 (N_24732,N_13163,N_10384);
xor U24733 (N_24733,N_17396,N_16410);
and U24734 (N_24734,N_17463,N_16884);
nor U24735 (N_24735,N_11347,N_10543);
nand U24736 (N_24736,N_13239,N_15754);
nand U24737 (N_24737,N_13607,N_18200);
and U24738 (N_24738,N_11474,N_12898);
and U24739 (N_24739,N_12851,N_13928);
and U24740 (N_24740,N_10555,N_18520);
and U24741 (N_24741,N_18841,N_17073);
or U24742 (N_24742,N_15982,N_10327);
nand U24743 (N_24743,N_13449,N_18094);
nor U24744 (N_24744,N_15685,N_12550);
or U24745 (N_24745,N_17653,N_13104);
nand U24746 (N_24746,N_10546,N_12303);
nand U24747 (N_24747,N_10876,N_18612);
or U24748 (N_24748,N_19889,N_19801);
and U24749 (N_24749,N_17713,N_19379);
and U24750 (N_24750,N_12627,N_13032);
nand U24751 (N_24751,N_17464,N_19084);
nand U24752 (N_24752,N_19873,N_17211);
or U24753 (N_24753,N_11603,N_10909);
nand U24754 (N_24754,N_11340,N_18723);
nor U24755 (N_24755,N_14000,N_17286);
and U24756 (N_24756,N_10246,N_19675);
nor U24757 (N_24757,N_19115,N_17807);
nor U24758 (N_24758,N_15446,N_16602);
or U24759 (N_24759,N_13452,N_11184);
nor U24760 (N_24760,N_10588,N_12499);
xor U24761 (N_24761,N_10456,N_15611);
or U24762 (N_24762,N_10025,N_16066);
or U24763 (N_24763,N_15891,N_14737);
or U24764 (N_24764,N_17305,N_18219);
nand U24765 (N_24765,N_14176,N_14928);
nand U24766 (N_24766,N_13764,N_14449);
and U24767 (N_24767,N_11610,N_10977);
or U24768 (N_24768,N_19721,N_18814);
nand U24769 (N_24769,N_10481,N_12453);
nor U24770 (N_24770,N_10198,N_15767);
or U24771 (N_24771,N_13495,N_17582);
xnor U24772 (N_24772,N_18366,N_11032);
xor U24773 (N_24773,N_14183,N_12266);
nand U24774 (N_24774,N_16635,N_16373);
and U24775 (N_24775,N_15450,N_14090);
and U24776 (N_24776,N_10418,N_19082);
and U24777 (N_24777,N_19267,N_10302);
nor U24778 (N_24778,N_10050,N_18157);
xnor U24779 (N_24779,N_14272,N_18832);
or U24780 (N_24780,N_17236,N_11567);
and U24781 (N_24781,N_16972,N_17368);
nor U24782 (N_24782,N_12051,N_16332);
xor U24783 (N_24783,N_12681,N_14585);
nand U24784 (N_24784,N_17609,N_11351);
nand U24785 (N_24785,N_14573,N_15111);
or U24786 (N_24786,N_14954,N_11654);
nor U24787 (N_24787,N_15016,N_19286);
nand U24788 (N_24788,N_10934,N_19291);
xnor U24789 (N_24789,N_18994,N_11982);
nand U24790 (N_24790,N_11888,N_12842);
nand U24791 (N_24791,N_18870,N_13162);
nor U24792 (N_24792,N_12761,N_18582);
or U24793 (N_24793,N_18672,N_18643);
nor U24794 (N_24794,N_16462,N_14012);
nor U24795 (N_24795,N_18667,N_13840);
and U24796 (N_24796,N_11426,N_15986);
nand U24797 (N_24797,N_18100,N_13339);
nor U24798 (N_24798,N_13547,N_14814);
nand U24799 (N_24799,N_14461,N_16057);
and U24800 (N_24800,N_19951,N_15598);
nand U24801 (N_24801,N_11681,N_19751);
or U24802 (N_24802,N_13159,N_19274);
nand U24803 (N_24803,N_13337,N_17231);
and U24804 (N_24804,N_11755,N_11980);
nand U24805 (N_24805,N_10745,N_14594);
nor U24806 (N_24806,N_16251,N_14826);
and U24807 (N_24807,N_14469,N_15517);
nor U24808 (N_24808,N_16309,N_13880);
or U24809 (N_24809,N_17101,N_19944);
and U24810 (N_24810,N_17549,N_15216);
or U24811 (N_24811,N_17608,N_12480);
xnor U24812 (N_24812,N_17321,N_16981);
and U24813 (N_24813,N_19477,N_11147);
and U24814 (N_24814,N_11789,N_14819);
or U24815 (N_24815,N_19559,N_15882);
or U24816 (N_24816,N_19831,N_13776);
and U24817 (N_24817,N_19430,N_10875);
nor U24818 (N_24818,N_14251,N_12424);
and U24819 (N_24819,N_13748,N_14192);
nand U24820 (N_24820,N_12854,N_17958);
xnor U24821 (N_24821,N_12072,N_11821);
nand U24822 (N_24822,N_13858,N_16324);
and U24823 (N_24823,N_14169,N_10554);
and U24824 (N_24824,N_15931,N_13802);
nor U24825 (N_24825,N_14129,N_18936);
nand U24826 (N_24826,N_18811,N_18394);
or U24827 (N_24827,N_17440,N_10127);
or U24828 (N_24828,N_14480,N_15852);
nand U24829 (N_24829,N_15414,N_19400);
or U24830 (N_24830,N_10643,N_10593);
xor U24831 (N_24831,N_14581,N_10812);
or U24832 (N_24832,N_19767,N_13759);
nor U24833 (N_24833,N_16273,N_16871);
nor U24834 (N_24834,N_15887,N_11529);
nand U24835 (N_24835,N_13992,N_16629);
nand U24836 (N_24836,N_18042,N_14278);
or U24837 (N_24837,N_11699,N_18940);
nand U24838 (N_24838,N_19055,N_13560);
or U24839 (N_24839,N_16476,N_18091);
or U24840 (N_24840,N_19097,N_12202);
nand U24841 (N_24841,N_11395,N_16486);
xnor U24842 (N_24842,N_16090,N_15473);
nand U24843 (N_24843,N_15975,N_19235);
nor U24844 (N_24844,N_11788,N_12440);
nand U24845 (N_24845,N_14891,N_14066);
nor U24846 (N_24846,N_10164,N_15398);
nor U24847 (N_24847,N_18515,N_17815);
or U24848 (N_24848,N_13256,N_15677);
xor U24849 (N_24849,N_11268,N_14640);
and U24850 (N_24850,N_19603,N_18777);
nand U24851 (N_24851,N_15361,N_10108);
nor U24852 (N_24852,N_17183,N_12556);
nand U24853 (N_24853,N_18711,N_16318);
xnor U24854 (N_24854,N_17121,N_14652);
and U24855 (N_24855,N_14227,N_19562);
and U24856 (N_24856,N_14242,N_14747);
nand U24857 (N_24857,N_16935,N_16126);
nor U24858 (N_24858,N_14416,N_11726);
or U24859 (N_24859,N_13055,N_16075);
and U24860 (N_24860,N_11570,N_14072);
or U24861 (N_24861,N_12987,N_16868);
nor U24862 (N_24862,N_15106,N_18112);
nor U24863 (N_24863,N_15976,N_18941);
nand U24864 (N_24864,N_12194,N_19835);
nor U24865 (N_24865,N_17181,N_17245);
nor U24866 (N_24866,N_16371,N_17484);
or U24867 (N_24867,N_11205,N_12402);
xnor U24868 (N_24868,N_17221,N_14778);
nand U24869 (N_24869,N_17672,N_18772);
nand U24870 (N_24870,N_14946,N_19739);
or U24871 (N_24871,N_14615,N_11703);
and U24872 (N_24872,N_14710,N_19205);
and U24873 (N_24873,N_17365,N_19450);
nand U24874 (N_24874,N_14582,N_13384);
or U24875 (N_24875,N_19044,N_15028);
nand U24876 (N_24876,N_19021,N_17933);
nand U24877 (N_24877,N_18309,N_13893);
nand U24878 (N_24878,N_14418,N_17701);
or U24879 (N_24879,N_11004,N_14595);
or U24880 (N_24880,N_12706,N_14393);
xor U24881 (N_24881,N_13613,N_11981);
and U24882 (N_24882,N_14355,N_18080);
nor U24883 (N_24883,N_10690,N_10328);
xnor U24884 (N_24884,N_15584,N_12245);
nand U24885 (N_24885,N_18872,N_13556);
nor U24886 (N_24886,N_10681,N_12459);
and U24887 (N_24887,N_14081,N_13340);
or U24888 (N_24888,N_11238,N_11440);
xor U24889 (N_24889,N_13220,N_10617);
nand U24890 (N_24890,N_15065,N_17789);
nor U24891 (N_24891,N_15643,N_13821);
xnor U24892 (N_24892,N_14600,N_16465);
and U24893 (N_24893,N_17492,N_10049);
xor U24894 (N_24894,N_12873,N_14738);
and U24895 (N_24895,N_17673,N_14746);
nor U24896 (N_24896,N_11523,N_11550);
nand U24897 (N_24897,N_17330,N_12356);
nand U24898 (N_24898,N_13927,N_18756);
or U24899 (N_24899,N_17495,N_11657);
nor U24900 (N_24900,N_13302,N_13478);
nand U24901 (N_24901,N_10693,N_17830);
nand U24902 (N_24902,N_18088,N_14289);
or U24903 (N_24903,N_15867,N_14171);
and U24904 (N_24904,N_10688,N_13008);
and U24905 (N_24905,N_12837,N_18144);
nand U24906 (N_24906,N_19804,N_10335);
nor U24907 (N_24907,N_18076,N_12639);
and U24908 (N_24908,N_18573,N_15270);
nor U24909 (N_24909,N_19451,N_14027);
and U24910 (N_24910,N_19986,N_17048);
or U24911 (N_24911,N_10376,N_10131);
and U24912 (N_24912,N_14874,N_10822);
and U24913 (N_24913,N_15075,N_15884);
and U24914 (N_24914,N_18538,N_14974);
xnor U24915 (N_24915,N_17934,N_17930);
nor U24916 (N_24916,N_14491,N_11486);
xor U24917 (N_24917,N_17498,N_14035);
and U24918 (N_24918,N_15514,N_18971);
or U24919 (N_24919,N_14118,N_16490);
and U24920 (N_24920,N_11686,N_18652);
or U24921 (N_24921,N_11284,N_10825);
and U24922 (N_24922,N_18336,N_12944);
or U24923 (N_24923,N_16136,N_15944);
nand U24924 (N_24924,N_10730,N_12153);
nor U24925 (N_24925,N_13771,N_10486);
and U24926 (N_24926,N_13363,N_18209);
or U24927 (N_24927,N_14339,N_14895);
xnor U24928 (N_24928,N_14157,N_19894);
or U24929 (N_24929,N_18962,N_15513);
nor U24930 (N_24930,N_14599,N_17594);
xor U24931 (N_24931,N_11823,N_15074);
nor U24932 (N_24932,N_12812,N_16498);
or U24933 (N_24933,N_18308,N_13174);
or U24934 (N_24934,N_10205,N_17544);
or U24935 (N_24935,N_14879,N_17923);
nor U24936 (N_24936,N_10009,N_14589);
and U24937 (N_24937,N_17895,N_18846);
nand U24938 (N_24938,N_13862,N_15656);
nor U24939 (N_24939,N_10279,N_19833);
or U24940 (N_24940,N_15349,N_17526);
nor U24941 (N_24941,N_15401,N_14715);
nor U24942 (N_24942,N_14906,N_14254);
xor U24943 (N_24943,N_13002,N_12092);
or U24944 (N_24944,N_11591,N_11951);
or U24945 (N_24945,N_10602,N_11450);
and U24946 (N_24946,N_10134,N_10532);
nor U24947 (N_24947,N_18744,N_13648);
or U24948 (N_24948,N_17473,N_16238);
nand U24949 (N_24949,N_16813,N_18450);
nor U24950 (N_24950,N_10249,N_15515);
nand U24951 (N_24951,N_11623,N_19158);
nor U24952 (N_24952,N_14020,N_12548);
nor U24953 (N_24953,N_16720,N_17217);
and U24954 (N_24954,N_15896,N_11759);
and U24955 (N_24955,N_11953,N_13617);
nor U24956 (N_24956,N_10139,N_13261);
nor U24957 (N_24957,N_13899,N_14091);
nor U24958 (N_24958,N_12752,N_12888);
and U24959 (N_24959,N_13792,N_11526);
and U24960 (N_24960,N_12768,N_11224);
and U24961 (N_24961,N_16693,N_10591);
nor U24962 (N_24962,N_16240,N_13642);
nor U24963 (N_24963,N_16897,N_11170);
nand U24964 (N_24964,N_12495,N_12777);
and U24965 (N_24965,N_17767,N_12304);
and U24966 (N_24966,N_11473,N_12261);
xnor U24967 (N_24967,N_16951,N_17619);
or U24968 (N_24968,N_14296,N_13005);
or U24969 (N_24969,N_12913,N_12065);
nor U24970 (N_24970,N_18706,N_14801);
or U24971 (N_24971,N_11770,N_10184);
or U24972 (N_24972,N_15178,N_16322);
nor U24973 (N_24973,N_14620,N_11958);
or U24974 (N_24974,N_16710,N_12312);
nand U24975 (N_24975,N_19634,N_19147);
and U24976 (N_24976,N_10054,N_16311);
nor U24977 (N_24977,N_15160,N_15116);
nand U24978 (N_24978,N_15201,N_14444);
nor U24979 (N_24979,N_13335,N_18506);
and U24980 (N_24980,N_16860,N_11611);
nand U24981 (N_24981,N_17921,N_17735);
and U24982 (N_24982,N_12341,N_19996);
or U24983 (N_24983,N_14095,N_13189);
and U24984 (N_24984,N_17002,N_17257);
nand U24985 (N_24985,N_16376,N_11727);
and U24986 (N_24986,N_15072,N_12215);
nand U24987 (N_24987,N_11602,N_16025);
or U24988 (N_24988,N_12405,N_14399);
xnor U24989 (N_24989,N_16262,N_19850);
nor U24990 (N_24990,N_11030,N_10170);
or U24991 (N_24991,N_15522,N_11002);
nand U24992 (N_24992,N_11357,N_18586);
nor U24993 (N_24993,N_11436,N_15786);
nor U24994 (N_24994,N_18412,N_19452);
nand U24995 (N_24995,N_13955,N_12650);
nand U24996 (N_24996,N_17491,N_18369);
and U24997 (N_24997,N_11083,N_12393);
or U24998 (N_24998,N_19974,N_15297);
and U24999 (N_24999,N_12956,N_10344);
or U25000 (N_25000,N_19216,N_11611);
and U25001 (N_25001,N_19378,N_16856);
and U25002 (N_25002,N_19647,N_11218);
nor U25003 (N_25003,N_11748,N_13145);
nor U25004 (N_25004,N_15761,N_19465);
or U25005 (N_25005,N_15317,N_11330);
or U25006 (N_25006,N_11559,N_10020);
nand U25007 (N_25007,N_17986,N_14489);
or U25008 (N_25008,N_17447,N_14672);
or U25009 (N_25009,N_15003,N_18417);
nand U25010 (N_25010,N_19682,N_11904);
nor U25011 (N_25011,N_13033,N_13550);
nand U25012 (N_25012,N_12710,N_13683);
nor U25013 (N_25013,N_17267,N_17774);
nor U25014 (N_25014,N_11923,N_11317);
nor U25015 (N_25015,N_15391,N_18939);
or U25016 (N_25016,N_10622,N_10080);
nor U25017 (N_25017,N_15457,N_14619);
or U25018 (N_25018,N_14131,N_11123);
nor U25019 (N_25019,N_19479,N_12138);
nand U25020 (N_25020,N_14357,N_19409);
nand U25021 (N_25021,N_19202,N_18785);
or U25022 (N_25022,N_12993,N_15221);
nor U25023 (N_25023,N_17789,N_14261);
nor U25024 (N_25024,N_11528,N_13237);
nand U25025 (N_25025,N_17762,N_12121);
and U25026 (N_25026,N_13340,N_14497);
or U25027 (N_25027,N_16355,N_18264);
or U25028 (N_25028,N_17451,N_19174);
and U25029 (N_25029,N_10694,N_15127);
and U25030 (N_25030,N_12042,N_18291);
nor U25031 (N_25031,N_15576,N_16467);
nand U25032 (N_25032,N_16649,N_10531);
nor U25033 (N_25033,N_11209,N_18673);
nor U25034 (N_25034,N_11100,N_14948);
nor U25035 (N_25035,N_14524,N_12929);
nor U25036 (N_25036,N_13603,N_17358);
or U25037 (N_25037,N_11871,N_14050);
or U25038 (N_25038,N_18301,N_16004);
and U25039 (N_25039,N_16511,N_12968);
nand U25040 (N_25040,N_11126,N_10500);
and U25041 (N_25041,N_17420,N_18720);
nor U25042 (N_25042,N_16357,N_11143);
nand U25043 (N_25043,N_11785,N_12585);
or U25044 (N_25044,N_16351,N_12092);
nor U25045 (N_25045,N_19280,N_17364);
xor U25046 (N_25046,N_19743,N_16113);
xor U25047 (N_25047,N_11990,N_17173);
and U25048 (N_25048,N_14871,N_11057);
nand U25049 (N_25049,N_18767,N_11160);
xnor U25050 (N_25050,N_10114,N_18075);
and U25051 (N_25051,N_19542,N_12992);
or U25052 (N_25052,N_11305,N_14987);
nand U25053 (N_25053,N_17021,N_18213);
nand U25054 (N_25054,N_19771,N_17168);
xor U25055 (N_25055,N_16084,N_16714);
nor U25056 (N_25056,N_19020,N_17784);
or U25057 (N_25057,N_14184,N_19491);
nand U25058 (N_25058,N_12470,N_16462);
nor U25059 (N_25059,N_16696,N_11904);
and U25060 (N_25060,N_12677,N_15597);
nand U25061 (N_25061,N_17380,N_16740);
nand U25062 (N_25062,N_17773,N_19306);
nand U25063 (N_25063,N_17540,N_17960);
and U25064 (N_25064,N_17188,N_10358);
nor U25065 (N_25065,N_11508,N_12326);
nand U25066 (N_25066,N_18337,N_14833);
or U25067 (N_25067,N_11693,N_15843);
nor U25068 (N_25068,N_12817,N_17404);
or U25069 (N_25069,N_16917,N_12242);
or U25070 (N_25070,N_12056,N_13230);
nor U25071 (N_25071,N_13954,N_10767);
and U25072 (N_25072,N_13534,N_18027);
nor U25073 (N_25073,N_17601,N_18831);
nand U25074 (N_25074,N_10688,N_19609);
and U25075 (N_25075,N_15540,N_10169);
xor U25076 (N_25076,N_18757,N_19186);
and U25077 (N_25077,N_19319,N_14395);
nand U25078 (N_25078,N_15602,N_12235);
nand U25079 (N_25079,N_11484,N_16870);
or U25080 (N_25080,N_11129,N_19617);
or U25081 (N_25081,N_13209,N_12116);
and U25082 (N_25082,N_13819,N_15153);
or U25083 (N_25083,N_15026,N_11999);
nor U25084 (N_25084,N_16276,N_14846);
and U25085 (N_25085,N_16231,N_18455);
or U25086 (N_25086,N_11021,N_15802);
and U25087 (N_25087,N_12984,N_14432);
or U25088 (N_25088,N_12210,N_18214);
nand U25089 (N_25089,N_18748,N_14181);
nor U25090 (N_25090,N_12959,N_12845);
and U25091 (N_25091,N_14179,N_17722);
nand U25092 (N_25092,N_11337,N_15981);
and U25093 (N_25093,N_11009,N_19210);
nor U25094 (N_25094,N_19354,N_12940);
or U25095 (N_25095,N_18481,N_11595);
nor U25096 (N_25096,N_16282,N_15007);
or U25097 (N_25097,N_14149,N_15589);
nor U25098 (N_25098,N_10018,N_12003);
nor U25099 (N_25099,N_16937,N_19896);
xor U25100 (N_25100,N_15439,N_11990);
xnor U25101 (N_25101,N_17496,N_13748);
and U25102 (N_25102,N_18612,N_11272);
or U25103 (N_25103,N_16472,N_13338);
or U25104 (N_25104,N_17039,N_10729);
nand U25105 (N_25105,N_19193,N_15985);
nand U25106 (N_25106,N_12542,N_15798);
nor U25107 (N_25107,N_11063,N_12319);
nand U25108 (N_25108,N_13778,N_19468);
nor U25109 (N_25109,N_16642,N_16372);
nand U25110 (N_25110,N_15810,N_18035);
xor U25111 (N_25111,N_15735,N_11652);
and U25112 (N_25112,N_19700,N_13814);
and U25113 (N_25113,N_18201,N_11170);
or U25114 (N_25114,N_14343,N_16568);
nor U25115 (N_25115,N_10403,N_15905);
xor U25116 (N_25116,N_13023,N_15533);
nor U25117 (N_25117,N_13219,N_16033);
or U25118 (N_25118,N_12729,N_14438);
nor U25119 (N_25119,N_10990,N_18929);
and U25120 (N_25120,N_13304,N_19124);
and U25121 (N_25121,N_12129,N_11166);
nor U25122 (N_25122,N_18285,N_16858);
or U25123 (N_25123,N_17724,N_13814);
nor U25124 (N_25124,N_19139,N_17700);
or U25125 (N_25125,N_13407,N_19036);
and U25126 (N_25126,N_13924,N_17599);
nand U25127 (N_25127,N_18455,N_19923);
nand U25128 (N_25128,N_11902,N_16677);
and U25129 (N_25129,N_18783,N_10516);
and U25130 (N_25130,N_19828,N_13284);
xnor U25131 (N_25131,N_13322,N_16942);
and U25132 (N_25132,N_18083,N_17339);
xor U25133 (N_25133,N_11752,N_12165);
or U25134 (N_25134,N_18787,N_10161);
or U25135 (N_25135,N_15828,N_19420);
and U25136 (N_25136,N_12242,N_14736);
nand U25137 (N_25137,N_14344,N_14518);
nand U25138 (N_25138,N_12373,N_12924);
xnor U25139 (N_25139,N_17863,N_17050);
and U25140 (N_25140,N_19889,N_17867);
nor U25141 (N_25141,N_14839,N_18975);
nor U25142 (N_25142,N_12831,N_16033);
or U25143 (N_25143,N_10458,N_15997);
and U25144 (N_25144,N_19086,N_11224);
nand U25145 (N_25145,N_14526,N_18285);
and U25146 (N_25146,N_15558,N_11786);
or U25147 (N_25147,N_15404,N_10505);
or U25148 (N_25148,N_16682,N_13893);
xor U25149 (N_25149,N_13872,N_13817);
xnor U25150 (N_25150,N_15358,N_13701);
or U25151 (N_25151,N_18173,N_17671);
and U25152 (N_25152,N_13653,N_19338);
or U25153 (N_25153,N_15497,N_19896);
or U25154 (N_25154,N_19461,N_14732);
or U25155 (N_25155,N_17465,N_15130);
and U25156 (N_25156,N_17986,N_19900);
nand U25157 (N_25157,N_11732,N_14818);
nor U25158 (N_25158,N_14391,N_12718);
nor U25159 (N_25159,N_10497,N_19998);
nor U25160 (N_25160,N_12789,N_12549);
or U25161 (N_25161,N_18619,N_10710);
nand U25162 (N_25162,N_13098,N_12697);
nor U25163 (N_25163,N_14209,N_17011);
or U25164 (N_25164,N_17126,N_11743);
nand U25165 (N_25165,N_19326,N_13231);
xor U25166 (N_25166,N_13674,N_10855);
and U25167 (N_25167,N_17081,N_18487);
and U25168 (N_25168,N_18365,N_14176);
nor U25169 (N_25169,N_15365,N_13639);
xnor U25170 (N_25170,N_13901,N_16083);
nand U25171 (N_25171,N_17141,N_17617);
nor U25172 (N_25172,N_11749,N_16339);
and U25173 (N_25173,N_14331,N_12898);
nor U25174 (N_25174,N_15086,N_17791);
nand U25175 (N_25175,N_12031,N_14817);
xnor U25176 (N_25176,N_18116,N_12626);
or U25177 (N_25177,N_14832,N_19907);
nor U25178 (N_25178,N_15035,N_16430);
nand U25179 (N_25179,N_10409,N_19170);
or U25180 (N_25180,N_17087,N_15847);
nand U25181 (N_25181,N_14055,N_13793);
xor U25182 (N_25182,N_14219,N_18993);
xnor U25183 (N_25183,N_12349,N_14818);
or U25184 (N_25184,N_10800,N_14722);
nand U25185 (N_25185,N_15202,N_13629);
nor U25186 (N_25186,N_12844,N_19546);
and U25187 (N_25187,N_15917,N_18651);
xor U25188 (N_25188,N_19397,N_17385);
or U25189 (N_25189,N_18789,N_16394);
and U25190 (N_25190,N_14442,N_19769);
and U25191 (N_25191,N_19131,N_12955);
and U25192 (N_25192,N_16643,N_11080);
nand U25193 (N_25193,N_13109,N_14169);
and U25194 (N_25194,N_18818,N_12370);
nor U25195 (N_25195,N_16957,N_15233);
and U25196 (N_25196,N_17842,N_17920);
nor U25197 (N_25197,N_10159,N_10403);
and U25198 (N_25198,N_18958,N_16618);
or U25199 (N_25199,N_19986,N_15022);
or U25200 (N_25200,N_12529,N_19475);
nor U25201 (N_25201,N_18381,N_19704);
nand U25202 (N_25202,N_17740,N_19882);
and U25203 (N_25203,N_18290,N_13319);
nor U25204 (N_25204,N_15686,N_12089);
nor U25205 (N_25205,N_17561,N_18077);
and U25206 (N_25206,N_10723,N_19294);
and U25207 (N_25207,N_18070,N_16344);
nand U25208 (N_25208,N_11263,N_17419);
nor U25209 (N_25209,N_13382,N_15822);
and U25210 (N_25210,N_16215,N_11912);
nor U25211 (N_25211,N_14045,N_12873);
xnor U25212 (N_25212,N_11769,N_15274);
or U25213 (N_25213,N_14175,N_13347);
or U25214 (N_25214,N_18532,N_18592);
and U25215 (N_25215,N_10637,N_15202);
and U25216 (N_25216,N_14701,N_19536);
or U25217 (N_25217,N_14656,N_18126);
nor U25218 (N_25218,N_18384,N_18895);
or U25219 (N_25219,N_11232,N_14073);
or U25220 (N_25220,N_13323,N_10867);
nand U25221 (N_25221,N_17853,N_10697);
and U25222 (N_25222,N_14295,N_13551);
nor U25223 (N_25223,N_18870,N_18419);
xor U25224 (N_25224,N_19250,N_18649);
and U25225 (N_25225,N_14120,N_11800);
nand U25226 (N_25226,N_16449,N_11940);
nand U25227 (N_25227,N_15966,N_19315);
xor U25228 (N_25228,N_11170,N_17242);
and U25229 (N_25229,N_13585,N_15580);
nand U25230 (N_25230,N_10624,N_10991);
nand U25231 (N_25231,N_14069,N_13501);
or U25232 (N_25232,N_17039,N_12940);
and U25233 (N_25233,N_12388,N_14513);
nor U25234 (N_25234,N_15059,N_12453);
nand U25235 (N_25235,N_12900,N_12183);
and U25236 (N_25236,N_18249,N_19212);
or U25237 (N_25237,N_18072,N_15030);
or U25238 (N_25238,N_11734,N_11963);
or U25239 (N_25239,N_18367,N_10558);
or U25240 (N_25240,N_19607,N_11587);
or U25241 (N_25241,N_19290,N_18212);
or U25242 (N_25242,N_12519,N_14930);
nor U25243 (N_25243,N_15388,N_19326);
and U25244 (N_25244,N_16300,N_17216);
nand U25245 (N_25245,N_10844,N_15820);
nand U25246 (N_25246,N_15239,N_14241);
nor U25247 (N_25247,N_15007,N_15168);
nand U25248 (N_25248,N_10174,N_17955);
nand U25249 (N_25249,N_10838,N_18512);
xor U25250 (N_25250,N_16161,N_10678);
and U25251 (N_25251,N_11819,N_16172);
xor U25252 (N_25252,N_17678,N_12685);
nor U25253 (N_25253,N_16748,N_16497);
and U25254 (N_25254,N_13179,N_14736);
nor U25255 (N_25255,N_16402,N_15614);
or U25256 (N_25256,N_14644,N_11198);
xor U25257 (N_25257,N_12654,N_11773);
nand U25258 (N_25258,N_18870,N_18731);
or U25259 (N_25259,N_18084,N_19456);
xnor U25260 (N_25260,N_18219,N_19137);
nand U25261 (N_25261,N_13839,N_13114);
and U25262 (N_25262,N_17249,N_14226);
nand U25263 (N_25263,N_13087,N_18902);
nand U25264 (N_25264,N_12814,N_12895);
nand U25265 (N_25265,N_14039,N_10745);
or U25266 (N_25266,N_16307,N_13421);
or U25267 (N_25267,N_17207,N_18581);
or U25268 (N_25268,N_12668,N_18929);
nor U25269 (N_25269,N_10417,N_17719);
nand U25270 (N_25270,N_19204,N_15759);
and U25271 (N_25271,N_18226,N_18407);
and U25272 (N_25272,N_16005,N_11297);
nor U25273 (N_25273,N_17508,N_18762);
or U25274 (N_25274,N_16924,N_10487);
or U25275 (N_25275,N_14392,N_17716);
nand U25276 (N_25276,N_12159,N_16212);
nor U25277 (N_25277,N_11730,N_11153);
and U25278 (N_25278,N_17483,N_18380);
or U25279 (N_25279,N_14016,N_12405);
or U25280 (N_25280,N_17042,N_11060);
xor U25281 (N_25281,N_16503,N_16587);
or U25282 (N_25282,N_11287,N_17590);
xnor U25283 (N_25283,N_14633,N_11265);
or U25284 (N_25284,N_17558,N_18558);
nor U25285 (N_25285,N_17708,N_13198);
nor U25286 (N_25286,N_14278,N_17928);
nor U25287 (N_25287,N_18079,N_19275);
and U25288 (N_25288,N_11214,N_14350);
or U25289 (N_25289,N_10704,N_15768);
nand U25290 (N_25290,N_13900,N_17102);
nand U25291 (N_25291,N_16332,N_17309);
or U25292 (N_25292,N_16056,N_12470);
and U25293 (N_25293,N_19986,N_14008);
nor U25294 (N_25294,N_16825,N_13938);
nor U25295 (N_25295,N_11074,N_16229);
or U25296 (N_25296,N_10362,N_11630);
and U25297 (N_25297,N_19867,N_11076);
and U25298 (N_25298,N_17941,N_16109);
nand U25299 (N_25299,N_11126,N_13987);
nor U25300 (N_25300,N_19190,N_18082);
or U25301 (N_25301,N_16105,N_13512);
or U25302 (N_25302,N_19439,N_14228);
nor U25303 (N_25303,N_18433,N_11025);
or U25304 (N_25304,N_18854,N_13527);
or U25305 (N_25305,N_18531,N_19734);
xnor U25306 (N_25306,N_12638,N_10784);
or U25307 (N_25307,N_15541,N_18724);
or U25308 (N_25308,N_12083,N_15506);
nor U25309 (N_25309,N_16067,N_13624);
and U25310 (N_25310,N_14989,N_17636);
or U25311 (N_25311,N_17297,N_19531);
or U25312 (N_25312,N_11183,N_12696);
or U25313 (N_25313,N_10845,N_19756);
nand U25314 (N_25314,N_11371,N_19290);
xor U25315 (N_25315,N_11704,N_13588);
and U25316 (N_25316,N_14924,N_11169);
nor U25317 (N_25317,N_18465,N_18574);
and U25318 (N_25318,N_12596,N_13901);
nor U25319 (N_25319,N_18061,N_10978);
and U25320 (N_25320,N_11137,N_17221);
and U25321 (N_25321,N_11677,N_16290);
nor U25322 (N_25322,N_19874,N_19529);
and U25323 (N_25323,N_12731,N_17484);
and U25324 (N_25324,N_10666,N_15257);
nor U25325 (N_25325,N_12779,N_15496);
or U25326 (N_25326,N_13890,N_16110);
and U25327 (N_25327,N_18913,N_16120);
or U25328 (N_25328,N_11309,N_14707);
or U25329 (N_25329,N_10124,N_15086);
nand U25330 (N_25330,N_17321,N_15468);
nor U25331 (N_25331,N_13295,N_11390);
nand U25332 (N_25332,N_17160,N_12177);
nand U25333 (N_25333,N_16558,N_19621);
nand U25334 (N_25334,N_14776,N_18778);
nor U25335 (N_25335,N_14706,N_15683);
nor U25336 (N_25336,N_16191,N_10815);
and U25337 (N_25337,N_14685,N_13121);
xnor U25338 (N_25338,N_18400,N_11236);
or U25339 (N_25339,N_16203,N_18068);
xor U25340 (N_25340,N_14382,N_12829);
nor U25341 (N_25341,N_18272,N_18730);
or U25342 (N_25342,N_19500,N_10784);
or U25343 (N_25343,N_15683,N_11420);
or U25344 (N_25344,N_10938,N_17291);
and U25345 (N_25345,N_17592,N_11759);
and U25346 (N_25346,N_18911,N_16101);
xor U25347 (N_25347,N_17297,N_18897);
nor U25348 (N_25348,N_13995,N_13927);
or U25349 (N_25349,N_14613,N_13843);
nand U25350 (N_25350,N_15171,N_17505);
nor U25351 (N_25351,N_14724,N_18226);
or U25352 (N_25352,N_14369,N_17564);
nand U25353 (N_25353,N_16502,N_17677);
nand U25354 (N_25354,N_19850,N_14574);
nand U25355 (N_25355,N_18178,N_19763);
nand U25356 (N_25356,N_18477,N_17934);
xor U25357 (N_25357,N_11814,N_10032);
and U25358 (N_25358,N_16078,N_11013);
and U25359 (N_25359,N_11933,N_16678);
nor U25360 (N_25360,N_15378,N_19063);
or U25361 (N_25361,N_11704,N_16893);
nor U25362 (N_25362,N_16936,N_14924);
and U25363 (N_25363,N_16729,N_11086);
nor U25364 (N_25364,N_15133,N_15587);
nor U25365 (N_25365,N_11833,N_19989);
or U25366 (N_25366,N_19340,N_14982);
and U25367 (N_25367,N_13340,N_17302);
nand U25368 (N_25368,N_19394,N_19288);
nand U25369 (N_25369,N_14393,N_19255);
nand U25370 (N_25370,N_12116,N_13975);
nand U25371 (N_25371,N_11509,N_19077);
or U25372 (N_25372,N_13668,N_16492);
or U25373 (N_25373,N_10217,N_15492);
nor U25374 (N_25374,N_17578,N_14381);
and U25375 (N_25375,N_16654,N_13319);
or U25376 (N_25376,N_12560,N_17672);
and U25377 (N_25377,N_17777,N_18506);
nor U25378 (N_25378,N_10970,N_12040);
nor U25379 (N_25379,N_19318,N_15629);
and U25380 (N_25380,N_11760,N_11495);
and U25381 (N_25381,N_16639,N_15903);
nand U25382 (N_25382,N_12876,N_18400);
nor U25383 (N_25383,N_14840,N_18383);
or U25384 (N_25384,N_12737,N_11108);
xor U25385 (N_25385,N_19614,N_18109);
nand U25386 (N_25386,N_18233,N_10819);
or U25387 (N_25387,N_15449,N_16812);
and U25388 (N_25388,N_11060,N_19227);
or U25389 (N_25389,N_15596,N_16711);
and U25390 (N_25390,N_14385,N_13906);
or U25391 (N_25391,N_17860,N_12154);
nor U25392 (N_25392,N_18028,N_16197);
nor U25393 (N_25393,N_14147,N_13669);
and U25394 (N_25394,N_11940,N_18978);
nand U25395 (N_25395,N_12200,N_13651);
and U25396 (N_25396,N_16445,N_15272);
nor U25397 (N_25397,N_13301,N_11747);
nand U25398 (N_25398,N_15664,N_18600);
nand U25399 (N_25399,N_13558,N_13213);
or U25400 (N_25400,N_10373,N_12515);
or U25401 (N_25401,N_17504,N_18999);
nor U25402 (N_25402,N_15151,N_14948);
nor U25403 (N_25403,N_15570,N_19792);
and U25404 (N_25404,N_19727,N_18564);
nand U25405 (N_25405,N_14057,N_14504);
nor U25406 (N_25406,N_16470,N_18121);
nand U25407 (N_25407,N_19149,N_16828);
and U25408 (N_25408,N_18339,N_17346);
nand U25409 (N_25409,N_17760,N_17412);
nand U25410 (N_25410,N_10868,N_12669);
nor U25411 (N_25411,N_10234,N_18037);
nor U25412 (N_25412,N_13750,N_14621);
or U25413 (N_25413,N_13554,N_14456);
and U25414 (N_25414,N_18010,N_16800);
nand U25415 (N_25415,N_16376,N_11821);
nand U25416 (N_25416,N_12461,N_18290);
and U25417 (N_25417,N_19064,N_13608);
nor U25418 (N_25418,N_13535,N_16734);
or U25419 (N_25419,N_16933,N_11066);
and U25420 (N_25420,N_12516,N_11577);
or U25421 (N_25421,N_19592,N_12557);
nand U25422 (N_25422,N_19289,N_17140);
nor U25423 (N_25423,N_17014,N_16577);
xnor U25424 (N_25424,N_15466,N_14256);
nor U25425 (N_25425,N_11029,N_15654);
xnor U25426 (N_25426,N_19007,N_18394);
nand U25427 (N_25427,N_19742,N_16652);
nand U25428 (N_25428,N_18670,N_12355);
and U25429 (N_25429,N_12304,N_10378);
and U25430 (N_25430,N_19086,N_15000);
or U25431 (N_25431,N_19515,N_16893);
nand U25432 (N_25432,N_10613,N_15090);
and U25433 (N_25433,N_17103,N_16778);
nand U25434 (N_25434,N_16526,N_15404);
nand U25435 (N_25435,N_14321,N_14134);
nand U25436 (N_25436,N_14772,N_19504);
nand U25437 (N_25437,N_12704,N_10335);
nand U25438 (N_25438,N_19853,N_11843);
or U25439 (N_25439,N_19253,N_18475);
xnor U25440 (N_25440,N_10965,N_13261);
nand U25441 (N_25441,N_13020,N_10410);
and U25442 (N_25442,N_10209,N_16675);
xor U25443 (N_25443,N_12119,N_13656);
xor U25444 (N_25444,N_12718,N_17420);
nand U25445 (N_25445,N_16868,N_16817);
or U25446 (N_25446,N_14224,N_14930);
or U25447 (N_25447,N_13189,N_12489);
and U25448 (N_25448,N_13049,N_18644);
xnor U25449 (N_25449,N_13833,N_19872);
nand U25450 (N_25450,N_17838,N_17466);
nand U25451 (N_25451,N_19459,N_18464);
and U25452 (N_25452,N_13071,N_16134);
or U25453 (N_25453,N_18247,N_13662);
xor U25454 (N_25454,N_19828,N_15443);
and U25455 (N_25455,N_13939,N_13480);
or U25456 (N_25456,N_14278,N_15433);
nor U25457 (N_25457,N_19466,N_16636);
or U25458 (N_25458,N_11111,N_19107);
or U25459 (N_25459,N_19011,N_18920);
and U25460 (N_25460,N_19072,N_11675);
or U25461 (N_25461,N_17467,N_10928);
nor U25462 (N_25462,N_12016,N_18662);
nor U25463 (N_25463,N_14323,N_13321);
xor U25464 (N_25464,N_16022,N_15758);
and U25465 (N_25465,N_15226,N_10993);
and U25466 (N_25466,N_10837,N_17653);
or U25467 (N_25467,N_11615,N_15944);
and U25468 (N_25468,N_15000,N_15316);
and U25469 (N_25469,N_16492,N_13661);
and U25470 (N_25470,N_13520,N_12520);
nand U25471 (N_25471,N_17263,N_19807);
and U25472 (N_25472,N_11313,N_17238);
nor U25473 (N_25473,N_12734,N_12716);
nor U25474 (N_25474,N_17615,N_15734);
and U25475 (N_25475,N_19425,N_12411);
nand U25476 (N_25476,N_10572,N_16623);
xnor U25477 (N_25477,N_14132,N_15098);
nor U25478 (N_25478,N_15686,N_11576);
nand U25479 (N_25479,N_12494,N_19465);
and U25480 (N_25480,N_19460,N_10087);
or U25481 (N_25481,N_17272,N_16049);
or U25482 (N_25482,N_12872,N_14070);
nor U25483 (N_25483,N_15938,N_18692);
nand U25484 (N_25484,N_10302,N_15188);
or U25485 (N_25485,N_16956,N_11143);
and U25486 (N_25486,N_15720,N_18618);
nand U25487 (N_25487,N_15592,N_18864);
or U25488 (N_25488,N_17739,N_16792);
nand U25489 (N_25489,N_17904,N_19934);
and U25490 (N_25490,N_14607,N_14361);
or U25491 (N_25491,N_15270,N_18682);
nor U25492 (N_25492,N_16226,N_14033);
and U25493 (N_25493,N_10835,N_12389);
and U25494 (N_25494,N_16598,N_10783);
nor U25495 (N_25495,N_18721,N_13701);
nand U25496 (N_25496,N_12492,N_14971);
nor U25497 (N_25497,N_10454,N_14297);
and U25498 (N_25498,N_17617,N_12987);
or U25499 (N_25499,N_13298,N_15577);
nor U25500 (N_25500,N_19217,N_13441);
or U25501 (N_25501,N_17594,N_10550);
nor U25502 (N_25502,N_12708,N_14242);
or U25503 (N_25503,N_18277,N_14487);
nand U25504 (N_25504,N_15564,N_17086);
nor U25505 (N_25505,N_18078,N_14827);
nand U25506 (N_25506,N_10214,N_15590);
or U25507 (N_25507,N_18969,N_12722);
nor U25508 (N_25508,N_10391,N_10040);
nand U25509 (N_25509,N_11367,N_15200);
or U25510 (N_25510,N_15821,N_15943);
or U25511 (N_25511,N_11494,N_18155);
or U25512 (N_25512,N_14158,N_17731);
nand U25513 (N_25513,N_16410,N_11440);
nand U25514 (N_25514,N_16662,N_13609);
and U25515 (N_25515,N_10674,N_13713);
nor U25516 (N_25516,N_10546,N_16343);
nand U25517 (N_25517,N_11600,N_18692);
or U25518 (N_25518,N_14237,N_14212);
nand U25519 (N_25519,N_15435,N_10571);
and U25520 (N_25520,N_13965,N_11727);
nand U25521 (N_25521,N_16021,N_11236);
or U25522 (N_25522,N_19347,N_11709);
and U25523 (N_25523,N_18452,N_12036);
xor U25524 (N_25524,N_16545,N_17542);
xor U25525 (N_25525,N_12064,N_17608);
or U25526 (N_25526,N_17561,N_17892);
or U25527 (N_25527,N_13280,N_10673);
and U25528 (N_25528,N_12772,N_19542);
nand U25529 (N_25529,N_13629,N_16264);
nor U25530 (N_25530,N_18175,N_19763);
nor U25531 (N_25531,N_18058,N_19765);
and U25532 (N_25532,N_15522,N_17592);
nor U25533 (N_25533,N_18706,N_11306);
nor U25534 (N_25534,N_12186,N_15607);
and U25535 (N_25535,N_17891,N_18368);
xnor U25536 (N_25536,N_18886,N_11651);
nor U25537 (N_25537,N_15569,N_19097);
and U25538 (N_25538,N_15207,N_14034);
or U25539 (N_25539,N_13009,N_15867);
or U25540 (N_25540,N_15004,N_17142);
or U25541 (N_25541,N_17817,N_16549);
xor U25542 (N_25542,N_16273,N_12374);
nand U25543 (N_25543,N_11344,N_17724);
nand U25544 (N_25544,N_14610,N_17568);
nand U25545 (N_25545,N_16525,N_13139);
nor U25546 (N_25546,N_11314,N_18068);
nand U25547 (N_25547,N_14863,N_15056);
nor U25548 (N_25548,N_16352,N_18886);
or U25549 (N_25549,N_10240,N_18849);
nor U25550 (N_25550,N_13102,N_17058);
nand U25551 (N_25551,N_15660,N_18071);
nand U25552 (N_25552,N_15024,N_12749);
nor U25553 (N_25553,N_10694,N_13761);
or U25554 (N_25554,N_18944,N_19949);
and U25555 (N_25555,N_10724,N_15899);
nand U25556 (N_25556,N_18090,N_15851);
and U25557 (N_25557,N_19077,N_19016);
and U25558 (N_25558,N_14490,N_12424);
nand U25559 (N_25559,N_13560,N_12582);
and U25560 (N_25560,N_14080,N_14374);
or U25561 (N_25561,N_14650,N_15467);
and U25562 (N_25562,N_12236,N_13102);
xnor U25563 (N_25563,N_13838,N_19162);
nor U25564 (N_25564,N_17848,N_10067);
or U25565 (N_25565,N_12145,N_17137);
or U25566 (N_25566,N_10903,N_15216);
nand U25567 (N_25567,N_10061,N_14824);
nor U25568 (N_25568,N_15947,N_11660);
xor U25569 (N_25569,N_18279,N_12053);
nand U25570 (N_25570,N_14020,N_16312);
or U25571 (N_25571,N_16737,N_19730);
and U25572 (N_25572,N_14462,N_18489);
nand U25573 (N_25573,N_17782,N_14639);
and U25574 (N_25574,N_10890,N_18978);
xnor U25575 (N_25575,N_12038,N_16024);
and U25576 (N_25576,N_16932,N_16237);
or U25577 (N_25577,N_17570,N_13098);
or U25578 (N_25578,N_15340,N_17378);
nor U25579 (N_25579,N_13449,N_15872);
xor U25580 (N_25580,N_10483,N_11269);
nand U25581 (N_25581,N_14496,N_10963);
and U25582 (N_25582,N_19700,N_19191);
nand U25583 (N_25583,N_10452,N_12906);
nor U25584 (N_25584,N_16647,N_12096);
and U25585 (N_25585,N_17370,N_10543);
nand U25586 (N_25586,N_18163,N_18491);
or U25587 (N_25587,N_19901,N_14561);
nor U25588 (N_25588,N_14410,N_17024);
xor U25589 (N_25589,N_16009,N_14221);
nand U25590 (N_25590,N_13012,N_17401);
nor U25591 (N_25591,N_12906,N_16181);
and U25592 (N_25592,N_17865,N_17378);
or U25593 (N_25593,N_13052,N_18653);
nor U25594 (N_25594,N_10710,N_10497);
nand U25595 (N_25595,N_14292,N_10544);
and U25596 (N_25596,N_15139,N_15803);
nand U25597 (N_25597,N_10781,N_17735);
nand U25598 (N_25598,N_10115,N_17285);
or U25599 (N_25599,N_13415,N_12492);
and U25600 (N_25600,N_10694,N_19962);
or U25601 (N_25601,N_12233,N_10444);
nand U25602 (N_25602,N_10651,N_17670);
and U25603 (N_25603,N_11932,N_14820);
nand U25604 (N_25604,N_18685,N_14588);
nor U25605 (N_25605,N_10326,N_16034);
or U25606 (N_25606,N_16094,N_17004);
or U25607 (N_25607,N_10688,N_10572);
nor U25608 (N_25608,N_18719,N_11620);
nor U25609 (N_25609,N_16394,N_11744);
or U25610 (N_25610,N_10193,N_16046);
nor U25611 (N_25611,N_12952,N_13555);
or U25612 (N_25612,N_15418,N_14250);
nand U25613 (N_25613,N_19268,N_18269);
or U25614 (N_25614,N_11665,N_12051);
nor U25615 (N_25615,N_18428,N_19221);
nor U25616 (N_25616,N_11408,N_14192);
and U25617 (N_25617,N_16363,N_11815);
nand U25618 (N_25618,N_15812,N_16847);
xnor U25619 (N_25619,N_10094,N_15332);
and U25620 (N_25620,N_15693,N_10028);
and U25621 (N_25621,N_19228,N_13514);
nand U25622 (N_25622,N_16663,N_12936);
or U25623 (N_25623,N_18830,N_16024);
nor U25624 (N_25624,N_12709,N_11456);
nor U25625 (N_25625,N_15033,N_18388);
nand U25626 (N_25626,N_11433,N_12797);
or U25627 (N_25627,N_10491,N_16510);
xor U25628 (N_25628,N_19923,N_17234);
and U25629 (N_25629,N_12709,N_12351);
nand U25630 (N_25630,N_13753,N_12125);
and U25631 (N_25631,N_10739,N_13066);
nor U25632 (N_25632,N_17939,N_19626);
or U25633 (N_25633,N_17026,N_12975);
nor U25634 (N_25634,N_15013,N_18861);
or U25635 (N_25635,N_10025,N_13900);
and U25636 (N_25636,N_11350,N_16908);
nor U25637 (N_25637,N_16775,N_16554);
nand U25638 (N_25638,N_17442,N_19735);
or U25639 (N_25639,N_14619,N_13461);
and U25640 (N_25640,N_10664,N_13462);
nor U25641 (N_25641,N_14814,N_12101);
nand U25642 (N_25642,N_19415,N_15033);
and U25643 (N_25643,N_18562,N_15387);
nand U25644 (N_25644,N_10373,N_10709);
or U25645 (N_25645,N_15026,N_16780);
xor U25646 (N_25646,N_18322,N_18902);
or U25647 (N_25647,N_16971,N_16424);
and U25648 (N_25648,N_12830,N_13144);
nor U25649 (N_25649,N_14026,N_11214);
nand U25650 (N_25650,N_11462,N_10865);
or U25651 (N_25651,N_10338,N_13440);
xor U25652 (N_25652,N_17406,N_14672);
nor U25653 (N_25653,N_11946,N_16974);
nand U25654 (N_25654,N_19326,N_19017);
or U25655 (N_25655,N_14293,N_16379);
and U25656 (N_25656,N_13592,N_15200);
xnor U25657 (N_25657,N_11024,N_18187);
xor U25658 (N_25658,N_19169,N_18153);
and U25659 (N_25659,N_17872,N_14751);
nor U25660 (N_25660,N_18200,N_12349);
or U25661 (N_25661,N_11155,N_17217);
xor U25662 (N_25662,N_12595,N_17262);
or U25663 (N_25663,N_11950,N_13356);
and U25664 (N_25664,N_12199,N_19573);
nand U25665 (N_25665,N_19809,N_16034);
and U25666 (N_25666,N_15357,N_11185);
and U25667 (N_25667,N_11424,N_18368);
or U25668 (N_25668,N_11610,N_17393);
nand U25669 (N_25669,N_19335,N_19043);
and U25670 (N_25670,N_14692,N_16173);
nor U25671 (N_25671,N_12662,N_18545);
or U25672 (N_25672,N_12114,N_18184);
nand U25673 (N_25673,N_14753,N_18507);
and U25674 (N_25674,N_17267,N_11152);
nand U25675 (N_25675,N_17026,N_10454);
or U25676 (N_25676,N_18818,N_14082);
nand U25677 (N_25677,N_16606,N_12690);
nor U25678 (N_25678,N_14158,N_14129);
nand U25679 (N_25679,N_19207,N_16282);
nor U25680 (N_25680,N_15023,N_15956);
and U25681 (N_25681,N_19591,N_16493);
and U25682 (N_25682,N_19660,N_19668);
and U25683 (N_25683,N_12186,N_13734);
nand U25684 (N_25684,N_17598,N_19905);
nand U25685 (N_25685,N_18956,N_17715);
and U25686 (N_25686,N_10833,N_17735);
nand U25687 (N_25687,N_15565,N_17259);
and U25688 (N_25688,N_16409,N_16621);
nand U25689 (N_25689,N_12163,N_13821);
nor U25690 (N_25690,N_18135,N_16351);
xnor U25691 (N_25691,N_19376,N_15357);
nor U25692 (N_25692,N_17839,N_14240);
nand U25693 (N_25693,N_15711,N_12650);
and U25694 (N_25694,N_19245,N_15402);
and U25695 (N_25695,N_15819,N_14364);
nor U25696 (N_25696,N_16913,N_18767);
or U25697 (N_25697,N_11745,N_10363);
or U25698 (N_25698,N_16910,N_14633);
xor U25699 (N_25699,N_11299,N_18658);
or U25700 (N_25700,N_13750,N_14865);
and U25701 (N_25701,N_12373,N_15953);
nand U25702 (N_25702,N_10040,N_19049);
nand U25703 (N_25703,N_14956,N_11127);
nor U25704 (N_25704,N_14095,N_12465);
nor U25705 (N_25705,N_13286,N_18778);
and U25706 (N_25706,N_12564,N_14270);
nand U25707 (N_25707,N_19311,N_11705);
xor U25708 (N_25708,N_14916,N_14083);
nand U25709 (N_25709,N_11471,N_14482);
nor U25710 (N_25710,N_18727,N_13688);
or U25711 (N_25711,N_19715,N_18585);
nand U25712 (N_25712,N_12881,N_14100);
nor U25713 (N_25713,N_11785,N_10506);
nor U25714 (N_25714,N_10113,N_12836);
and U25715 (N_25715,N_18263,N_10193);
nor U25716 (N_25716,N_18178,N_12721);
nand U25717 (N_25717,N_19291,N_11976);
or U25718 (N_25718,N_15029,N_18948);
nand U25719 (N_25719,N_10145,N_19205);
nor U25720 (N_25720,N_11419,N_15318);
nor U25721 (N_25721,N_17691,N_16486);
nand U25722 (N_25722,N_16023,N_13783);
nand U25723 (N_25723,N_12020,N_16890);
and U25724 (N_25724,N_17007,N_14320);
or U25725 (N_25725,N_19010,N_10439);
or U25726 (N_25726,N_15046,N_16747);
or U25727 (N_25727,N_11780,N_17028);
and U25728 (N_25728,N_11886,N_11865);
or U25729 (N_25729,N_19606,N_14626);
xnor U25730 (N_25730,N_11564,N_13246);
or U25731 (N_25731,N_11983,N_16049);
or U25732 (N_25732,N_17224,N_18537);
xnor U25733 (N_25733,N_11430,N_12688);
xnor U25734 (N_25734,N_17324,N_16238);
nor U25735 (N_25735,N_19534,N_19058);
nor U25736 (N_25736,N_10932,N_19308);
nor U25737 (N_25737,N_14705,N_13288);
and U25738 (N_25738,N_19909,N_15821);
and U25739 (N_25739,N_16155,N_11276);
nand U25740 (N_25740,N_10572,N_18220);
or U25741 (N_25741,N_14066,N_10895);
or U25742 (N_25742,N_15603,N_15098);
nor U25743 (N_25743,N_10562,N_10352);
nor U25744 (N_25744,N_19299,N_17391);
xnor U25745 (N_25745,N_13929,N_11408);
nand U25746 (N_25746,N_10112,N_10958);
and U25747 (N_25747,N_16965,N_10585);
nand U25748 (N_25748,N_17400,N_19936);
nor U25749 (N_25749,N_18603,N_14634);
xnor U25750 (N_25750,N_15874,N_15810);
and U25751 (N_25751,N_14124,N_12137);
and U25752 (N_25752,N_13805,N_18771);
xnor U25753 (N_25753,N_19706,N_14552);
nor U25754 (N_25754,N_16344,N_12619);
nand U25755 (N_25755,N_10122,N_13046);
nand U25756 (N_25756,N_16820,N_16986);
nor U25757 (N_25757,N_15316,N_12819);
nor U25758 (N_25758,N_14194,N_11174);
nor U25759 (N_25759,N_10002,N_18744);
xor U25760 (N_25760,N_13494,N_15010);
nand U25761 (N_25761,N_15929,N_15665);
nor U25762 (N_25762,N_18648,N_14049);
or U25763 (N_25763,N_17983,N_13095);
nor U25764 (N_25764,N_14488,N_18033);
nand U25765 (N_25765,N_15388,N_14215);
nand U25766 (N_25766,N_17881,N_11628);
and U25767 (N_25767,N_10270,N_15278);
or U25768 (N_25768,N_19990,N_17409);
and U25769 (N_25769,N_13400,N_12968);
nand U25770 (N_25770,N_12813,N_12092);
nor U25771 (N_25771,N_18709,N_16889);
nand U25772 (N_25772,N_15603,N_16581);
and U25773 (N_25773,N_18003,N_15024);
nor U25774 (N_25774,N_17685,N_19767);
and U25775 (N_25775,N_16754,N_10071);
and U25776 (N_25776,N_10915,N_17022);
or U25777 (N_25777,N_12515,N_17791);
nand U25778 (N_25778,N_10174,N_12902);
xor U25779 (N_25779,N_17531,N_10597);
and U25780 (N_25780,N_10349,N_10561);
xnor U25781 (N_25781,N_18517,N_13612);
nand U25782 (N_25782,N_13319,N_12880);
or U25783 (N_25783,N_17669,N_13129);
or U25784 (N_25784,N_16354,N_11999);
nor U25785 (N_25785,N_18478,N_11826);
nor U25786 (N_25786,N_11579,N_12635);
or U25787 (N_25787,N_18883,N_12795);
or U25788 (N_25788,N_13026,N_13609);
or U25789 (N_25789,N_11410,N_19229);
and U25790 (N_25790,N_12531,N_15488);
xor U25791 (N_25791,N_13293,N_14103);
or U25792 (N_25792,N_15603,N_14051);
nor U25793 (N_25793,N_15911,N_19558);
or U25794 (N_25794,N_10682,N_13582);
and U25795 (N_25795,N_11931,N_15580);
or U25796 (N_25796,N_11179,N_12021);
or U25797 (N_25797,N_19090,N_13140);
nand U25798 (N_25798,N_13498,N_11441);
and U25799 (N_25799,N_15367,N_15337);
xnor U25800 (N_25800,N_10528,N_12585);
and U25801 (N_25801,N_17109,N_10334);
and U25802 (N_25802,N_12819,N_19624);
and U25803 (N_25803,N_11740,N_18838);
nor U25804 (N_25804,N_14058,N_15793);
nand U25805 (N_25805,N_17646,N_16059);
and U25806 (N_25806,N_11422,N_15411);
nor U25807 (N_25807,N_13526,N_13501);
nand U25808 (N_25808,N_18628,N_11231);
and U25809 (N_25809,N_17827,N_10212);
nand U25810 (N_25810,N_15489,N_19996);
and U25811 (N_25811,N_18019,N_18624);
xnor U25812 (N_25812,N_15828,N_17135);
nor U25813 (N_25813,N_16428,N_17115);
nor U25814 (N_25814,N_16351,N_19613);
and U25815 (N_25815,N_15408,N_13199);
or U25816 (N_25816,N_19604,N_11990);
and U25817 (N_25817,N_11677,N_14984);
nor U25818 (N_25818,N_17695,N_14826);
and U25819 (N_25819,N_13430,N_11019);
nand U25820 (N_25820,N_15685,N_11914);
nand U25821 (N_25821,N_14785,N_11014);
nor U25822 (N_25822,N_19782,N_13007);
nor U25823 (N_25823,N_19993,N_11571);
nand U25824 (N_25824,N_12152,N_11623);
and U25825 (N_25825,N_19149,N_10448);
or U25826 (N_25826,N_10699,N_14128);
and U25827 (N_25827,N_14581,N_14585);
nand U25828 (N_25828,N_15662,N_18236);
nor U25829 (N_25829,N_16109,N_18810);
and U25830 (N_25830,N_13783,N_15933);
xnor U25831 (N_25831,N_10087,N_14911);
nand U25832 (N_25832,N_13573,N_12990);
nor U25833 (N_25833,N_12503,N_11436);
nand U25834 (N_25834,N_18469,N_12175);
nand U25835 (N_25835,N_13008,N_12369);
xor U25836 (N_25836,N_16438,N_13661);
and U25837 (N_25837,N_14120,N_15147);
nor U25838 (N_25838,N_18878,N_19231);
and U25839 (N_25839,N_15191,N_19742);
and U25840 (N_25840,N_15558,N_19930);
nand U25841 (N_25841,N_12877,N_15157);
or U25842 (N_25842,N_15654,N_16829);
nor U25843 (N_25843,N_12654,N_15596);
and U25844 (N_25844,N_18153,N_10234);
or U25845 (N_25845,N_13275,N_17437);
or U25846 (N_25846,N_17796,N_19245);
nand U25847 (N_25847,N_17873,N_18338);
nor U25848 (N_25848,N_15145,N_19230);
and U25849 (N_25849,N_13410,N_15526);
xnor U25850 (N_25850,N_17775,N_16726);
nand U25851 (N_25851,N_19725,N_14558);
and U25852 (N_25852,N_15282,N_19988);
nor U25853 (N_25853,N_12794,N_11596);
and U25854 (N_25854,N_10880,N_17170);
nand U25855 (N_25855,N_10927,N_18250);
and U25856 (N_25856,N_17289,N_18942);
nand U25857 (N_25857,N_16623,N_13217);
nand U25858 (N_25858,N_10715,N_15448);
or U25859 (N_25859,N_12465,N_16550);
nand U25860 (N_25860,N_13775,N_15300);
nand U25861 (N_25861,N_10582,N_12478);
or U25862 (N_25862,N_10682,N_18870);
and U25863 (N_25863,N_14369,N_14925);
and U25864 (N_25864,N_17171,N_14257);
nor U25865 (N_25865,N_15744,N_17802);
nor U25866 (N_25866,N_14121,N_11042);
nor U25867 (N_25867,N_14261,N_11324);
or U25868 (N_25868,N_17106,N_14255);
or U25869 (N_25869,N_18707,N_18943);
and U25870 (N_25870,N_16654,N_13223);
nand U25871 (N_25871,N_11956,N_16590);
and U25872 (N_25872,N_19382,N_18720);
nand U25873 (N_25873,N_15118,N_11599);
and U25874 (N_25874,N_15422,N_18294);
and U25875 (N_25875,N_16545,N_18195);
and U25876 (N_25876,N_12018,N_15556);
nand U25877 (N_25877,N_16674,N_19368);
or U25878 (N_25878,N_13827,N_13881);
or U25879 (N_25879,N_15899,N_15769);
and U25880 (N_25880,N_10036,N_13113);
nand U25881 (N_25881,N_14826,N_17006);
xor U25882 (N_25882,N_10425,N_11842);
and U25883 (N_25883,N_15583,N_12091);
nand U25884 (N_25884,N_18158,N_16480);
nand U25885 (N_25885,N_14975,N_13135);
nand U25886 (N_25886,N_11690,N_19129);
nand U25887 (N_25887,N_12177,N_18786);
nor U25888 (N_25888,N_12172,N_18334);
and U25889 (N_25889,N_10233,N_14351);
nand U25890 (N_25890,N_13457,N_12820);
nor U25891 (N_25891,N_16221,N_13549);
nand U25892 (N_25892,N_19382,N_18481);
nor U25893 (N_25893,N_12950,N_12806);
nor U25894 (N_25894,N_10547,N_10808);
xor U25895 (N_25895,N_10619,N_15723);
nand U25896 (N_25896,N_18941,N_18404);
xnor U25897 (N_25897,N_17441,N_16402);
or U25898 (N_25898,N_12312,N_12913);
xnor U25899 (N_25899,N_13971,N_15643);
or U25900 (N_25900,N_14074,N_17928);
nand U25901 (N_25901,N_12090,N_11820);
and U25902 (N_25902,N_16338,N_11054);
and U25903 (N_25903,N_12472,N_18179);
or U25904 (N_25904,N_12298,N_13881);
or U25905 (N_25905,N_14308,N_19551);
nand U25906 (N_25906,N_19573,N_12229);
xor U25907 (N_25907,N_19728,N_15057);
xor U25908 (N_25908,N_18088,N_11178);
and U25909 (N_25909,N_16058,N_15230);
nand U25910 (N_25910,N_14995,N_11194);
or U25911 (N_25911,N_11521,N_14773);
or U25912 (N_25912,N_16366,N_15995);
or U25913 (N_25913,N_19914,N_13462);
nand U25914 (N_25914,N_17923,N_17367);
and U25915 (N_25915,N_15327,N_11427);
nand U25916 (N_25916,N_18003,N_13158);
nor U25917 (N_25917,N_11653,N_15622);
nor U25918 (N_25918,N_18430,N_16284);
and U25919 (N_25919,N_16517,N_12357);
xor U25920 (N_25920,N_17860,N_12159);
nand U25921 (N_25921,N_12775,N_10420);
nor U25922 (N_25922,N_10282,N_17167);
and U25923 (N_25923,N_11768,N_19870);
or U25924 (N_25924,N_12260,N_12802);
nor U25925 (N_25925,N_19406,N_15988);
xnor U25926 (N_25926,N_12983,N_17446);
and U25927 (N_25927,N_14331,N_18739);
nand U25928 (N_25928,N_10044,N_15649);
and U25929 (N_25929,N_16041,N_12496);
xnor U25930 (N_25930,N_12202,N_19820);
or U25931 (N_25931,N_13050,N_18174);
or U25932 (N_25932,N_12170,N_18784);
nand U25933 (N_25933,N_18450,N_16537);
and U25934 (N_25934,N_16265,N_15899);
nor U25935 (N_25935,N_11358,N_16311);
nor U25936 (N_25936,N_15458,N_16518);
nand U25937 (N_25937,N_18370,N_12253);
nand U25938 (N_25938,N_10881,N_12710);
nand U25939 (N_25939,N_15973,N_12456);
nor U25940 (N_25940,N_14254,N_12804);
nor U25941 (N_25941,N_12301,N_10744);
nor U25942 (N_25942,N_10325,N_12462);
nand U25943 (N_25943,N_17505,N_12162);
or U25944 (N_25944,N_10668,N_15733);
and U25945 (N_25945,N_16814,N_11850);
or U25946 (N_25946,N_11299,N_14672);
nand U25947 (N_25947,N_11454,N_15017);
nor U25948 (N_25948,N_15105,N_11310);
or U25949 (N_25949,N_18310,N_19517);
xnor U25950 (N_25950,N_13559,N_17649);
xor U25951 (N_25951,N_12850,N_16232);
and U25952 (N_25952,N_13872,N_19040);
nor U25953 (N_25953,N_10265,N_12657);
and U25954 (N_25954,N_10171,N_17757);
xnor U25955 (N_25955,N_11269,N_19929);
xor U25956 (N_25956,N_15166,N_14651);
or U25957 (N_25957,N_10903,N_11589);
nand U25958 (N_25958,N_15430,N_13868);
and U25959 (N_25959,N_19818,N_12752);
and U25960 (N_25960,N_12886,N_17026);
nand U25961 (N_25961,N_17974,N_18800);
or U25962 (N_25962,N_18101,N_16783);
or U25963 (N_25963,N_17711,N_14460);
and U25964 (N_25964,N_19648,N_18688);
nor U25965 (N_25965,N_19302,N_10631);
nand U25966 (N_25966,N_10722,N_13082);
nor U25967 (N_25967,N_15450,N_18031);
and U25968 (N_25968,N_19718,N_11648);
and U25969 (N_25969,N_16901,N_15131);
xnor U25970 (N_25970,N_13723,N_13183);
or U25971 (N_25971,N_18965,N_10698);
nor U25972 (N_25972,N_12228,N_11731);
nor U25973 (N_25973,N_19744,N_14822);
xor U25974 (N_25974,N_17609,N_12312);
or U25975 (N_25975,N_19634,N_19556);
and U25976 (N_25976,N_14300,N_10917);
nand U25977 (N_25977,N_16047,N_12675);
or U25978 (N_25978,N_15570,N_17842);
and U25979 (N_25979,N_11652,N_10186);
or U25980 (N_25980,N_19967,N_12813);
nand U25981 (N_25981,N_15124,N_13831);
and U25982 (N_25982,N_18381,N_17546);
xor U25983 (N_25983,N_17527,N_17867);
and U25984 (N_25984,N_11722,N_12854);
xnor U25985 (N_25985,N_11063,N_18146);
nand U25986 (N_25986,N_13647,N_18491);
or U25987 (N_25987,N_16286,N_16797);
nor U25988 (N_25988,N_14793,N_15482);
nand U25989 (N_25989,N_13322,N_10111);
nor U25990 (N_25990,N_12963,N_12538);
nand U25991 (N_25991,N_10779,N_13052);
nand U25992 (N_25992,N_15763,N_15963);
nor U25993 (N_25993,N_17327,N_11412);
nand U25994 (N_25994,N_19875,N_18698);
nor U25995 (N_25995,N_11249,N_13609);
xor U25996 (N_25996,N_16890,N_11087);
nand U25997 (N_25997,N_15427,N_15168);
nand U25998 (N_25998,N_12022,N_10109);
or U25999 (N_25999,N_19569,N_17460);
nand U26000 (N_26000,N_12605,N_10570);
or U26001 (N_26001,N_16135,N_13830);
nor U26002 (N_26002,N_16209,N_14799);
nand U26003 (N_26003,N_19836,N_10252);
nand U26004 (N_26004,N_11035,N_18116);
or U26005 (N_26005,N_18610,N_15461);
and U26006 (N_26006,N_14282,N_11603);
and U26007 (N_26007,N_13433,N_10674);
nor U26008 (N_26008,N_12245,N_14956);
or U26009 (N_26009,N_15002,N_15111);
nor U26010 (N_26010,N_13836,N_12200);
or U26011 (N_26011,N_18926,N_14932);
nand U26012 (N_26012,N_12975,N_10653);
nor U26013 (N_26013,N_19392,N_12764);
and U26014 (N_26014,N_10921,N_18022);
nand U26015 (N_26015,N_16362,N_13313);
or U26016 (N_26016,N_15984,N_10858);
nand U26017 (N_26017,N_12223,N_13675);
nand U26018 (N_26018,N_17584,N_13016);
nand U26019 (N_26019,N_10823,N_19354);
nand U26020 (N_26020,N_17098,N_16457);
or U26021 (N_26021,N_13941,N_10137);
and U26022 (N_26022,N_19253,N_19992);
and U26023 (N_26023,N_14455,N_17247);
or U26024 (N_26024,N_14461,N_13898);
or U26025 (N_26025,N_10163,N_10159);
and U26026 (N_26026,N_19826,N_10183);
nand U26027 (N_26027,N_13473,N_11780);
nor U26028 (N_26028,N_19419,N_12622);
and U26029 (N_26029,N_19898,N_10715);
nand U26030 (N_26030,N_18350,N_17961);
nor U26031 (N_26031,N_15824,N_19054);
nand U26032 (N_26032,N_13543,N_15066);
nor U26033 (N_26033,N_18436,N_18103);
and U26034 (N_26034,N_17247,N_17941);
and U26035 (N_26035,N_17755,N_16354);
xnor U26036 (N_26036,N_19309,N_14974);
or U26037 (N_26037,N_18129,N_16142);
nand U26038 (N_26038,N_12388,N_19802);
nand U26039 (N_26039,N_15881,N_12245);
nor U26040 (N_26040,N_17230,N_12479);
nor U26041 (N_26041,N_12562,N_19844);
and U26042 (N_26042,N_12848,N_17431);
nand U26043 (N_26043,N_13501,N_14746);
or U26044 (N_26044,N_17625,N_17751);
nand U26045 (N_26045,N_13524,N_17288);
or U26046 (N_26046,N_15812,N_18289);
and U26047 (N_26047,N_12420,N_19217);
xnor U26048 (N_26048,N_11642,N_16666);
and U26049 (N_26049,N_19082,N_19347);
or U26050 (N_26050,N_14414,N_16377);
and U26051 (N_26051,N_16778,N_15725);
nand U26052 (N_26052,N_19187,N_10192);
and U26053 (N_26053,N_11438,N_19255);
nand U26054 (N_26054,N_17183,N_15692);
and U26055 (N_26055,N_17322,N_10648);
nand U26056 (N_26056,N_11872,N_14977);
xor U26057 (N_26057,N_17459,N_17363);
and U26058 (N_26058,N_12799,N_15344);
and U26059 (N_26059,N_10414,N_11286);
and U26060 (N_26060,N_18766,N_16750);
and U26061 (N_26061,N_15181,N_11291);
and U26062 (N_26062,N_15035,N_15236);
nor U26063 (N_26063,N_11390,N_13611);
nand U26064 (N_26064,N_17731,N_11355);
or U26065 (N_26065,N_16522,N_11923);
or U26066 (N_26066,N_11327,N_17498);
or U26067 (N_26067,N_17056,N_15062);
nor U26068 (N_26068,N_17372,N_15959);
nand U26069 (N_26069,N_14114,N_17077);
or U26070 (N_26070,N_17226,N_16009);
and U26071 (N_26071,N_10258,N_11867);
and U26072 (N_26072,N_13908,N_16529);
nand U26073 (N_26073,N_10440,N_15478);
xor U26074 (N_26074,N_12571,N_12194);
nand U26075 (N_26075,N_15380,N_18728);
and U26076 (N_26076,N_12979,N_11078);
nor U26077 (N_26077,N_10321,N_17203);
and U26078 (N_26078,N_14435,N_19331);
or U26079 (N_26079,N_13317,N_11199);
nand U26080 (N_26080,N_17588,N_10311);
nor U26081 (N_26081,N_19803,N_13066);
nand U26082 (N_26082,N_10042,N_11684);
xnor U26083 (N_26083,N_13434,N_12387);
xor U26084 (N_26084,N_11223,N_18957);
nand U26085 (N_26085,N_12856,N_16462);
or U26086 (N_26086,N_16928,N_15887);
nand U26087 (N_26087,N_13169,N_16532);
xor U26088 (N_26088,N_16428,N_16838);
or U26089 (N_26089,N_11281,N_12942);
nor U26090 (N_26090,N_12375,N_16635);
or U26091 (N_26091,N_15203,N_16689);
or U26092 (N_26092,N_16561,N_10891);
nand U26093 (N_26093,N_12510,N_10692);
nand U26094 (N_26094,N_10469,N_14525);
xnor U26095 (N_26095,N_14377,N_18897);
or U26096 (N_26096,N_18282,N_12324);
nor U26097 (N_26097,N_12168,N_18962);
or U26098 (N_26098,N_15840,N_18774);
or U26099 (N_26099,N_14528,N_19669);
nand U26100 (N_26100,N_11269,N_10476);
nand U26101 (N_26101,N_10355,N_13069);
or U26102 (N_26102,N_14851,N_15057);
nand U26103 (N_26103,N_17160,N_15579);
xnor U26104 (N_26104,N_16320,N_13889);
nor U26105 (N_26105,N_13966,N_15142);
xor U26106 (N_26106,N_15676,N_10911);
nand U26107 (N_26107,N_16752,N_15134);
or U26108 (N_26108,N_18707,N_19292);
and U26109 (N_26109,N_12994,N_16873);
or U26110 (N_26110,N_13226,N_13532);
nand U26111 (N_26111,N_16937,N_18700);
nand U26112 (N_26112,N_13518,N_16189);
nand U26113 (N_26113,N_13789,N_19074);
nand U26114 (N_26114,N_16247,N_18378);
and U26115 (N_26115,N_11726,N_10121);
xor U26116 (N_26116,N_15683,N_15861);
nor U26117 (N_26117,N_10572,N_12105);
nor U26118 (N_26118,N_18925,N_14694);
xor U26119 (N_26119,N_17660,N_14389);
and U26120 (N_26120,N_19516,N_14245);
nand U26121 (N_26121,N_15303,N_18820);
nand U26122 (N_26122,N_10370,N_15654);
xnor U26123 (N_26123,N_18181,N_11400);
or U26124 (N_26124,N_12202,N_18847);
xor U26125 (N_26125,N_15055,N_13858);
nor U26126 (N_26126,N_12421,N_12393);
or U26127 (N_26127,N_14729,N_17783);
nor U26128 (N_26128,N_16437,N_11878);
xnor U26129 (N_26129,N_13889,N_13006);
nor U26130 (N_26130,N_19091,N_16158);
nand U26131 (N_26131,N_17431,N_11243);
or U26132 (N_26132,N_18240,N_17460);
nor U26133 (N_26133,N_19242,N_10049);
nor U26134 (N_26134,N_14673,N_19002);
nor U26135 (N_26135,N_10052,N_15792);
nor U26136 (N_26136,N_16490,N_11193);
and U26137 (N_26137,N_13865,N_12978);
nor U26138 (N_26138,N_17753,N_12418);
xor U26139 (N_26139,N_15928,N_18562);
nand U26140 (N_26140,N_13172,N_10572);
nor U26141 (N_26141,N_13816,N_10853);
and U26142 (N_26142,N_11485,N_17084);
nand U26143 (N_26143,N_19193,N_11901);
or U26144 (N_26144,N_13474,N_18452);
nand U26145 (N_26145,N_11493,N_13389);
nor U26146 (N_26146,N_17540,N_17092);
nand U26147 (N_26147,N_19417,N_10971);
nor U26148 (N_26148,N_16186,N_10406);
and U26149 (N_26149,N_19624,N_14506);
or U26150 (N_26150,N_19403,N_16660);
and U26151 (N_26151,N_13046,N_19046);
and U26152 (N_26152,N_18885,N_18447);
and U26153 (N_26153,N_16657,N_12444);
xnor U26154 (N_26154,N_13692,N_14903);
nor U26155 (N_26155,N_16071,N_18442);
xnor U26156 (N_26156,N_13749,N_10938);
or U26157 (N_26157,N_16092,N_18013);
and U26158 (N_26158,N_14280,N_12239);
nand U26159 (N_26159,N_14435,N_13553);
or U26160 (N_26160,N_18031,N_10388);
nand U26161 (N_26161,N_19449,N_14681);
nor U26162 (N_26162,N_18180,N_14912);
nor U26163 (N_26163,N_18888,N_12702);
or U26164 (N_26164,N_13265,N_19490);
nor U26165 (N_26165,N_12028,N_17314);
nor U26166 (N_26166,N_19406,N_15720);
nand U26167 (N_26167,N_14535,N_14721);
or U26168 (N_26168,N_13898,N_12490);
and U26169 (N_26169,N_11257,N_14469);
and U26170 (N_26170,N_15859,N_13526);
and U26171 (N_26171,N_10989,N_19953);
xor U26172 (N_26172,N_12287,N_14895);
xor U26173 (N_26173,N_19197,N_14924);
nand U26174 (N_26174,N_11396,N_15130);
and U26175 (N_26175,N_17745,N_19337);
and U26176 (N_26176,N_13650,N_15878);
xnor U26177 (N_26177,N_10448,N_13988);
or U26178 (N_26178,N_16129,N_19625);
and U26179 (N_26179,N_15467,N_19645);
and U26180 (N_26180,N_16254,N_15675);
nor U26181 (N_26181,N_13189,N_18496);
nand U26182 (N_26182,N_17868,N_16346);
nor U26183 (N_26183,N_14320,N_11116);
xnor U26184 (N_26184,N_17671,N_10987);
xor U26185 (N_26185,N_14173,N_16780);
nand U26186 (N_26186,N_17617,N_12765);
nand U26187 (N_26187,N_17782,N_12821);
and U26188 (N_26188,N_10726,N_12964);
or U26189 (N_26189,N_15271,N_15398);
xor U26190 (N_26190,N_10740,N_11711);
nand U26191 (N_26191,N_15667,N_10836);
nor U26192 (N_26192,N_15900,N_11942);
or U26193 (N_26193,N_15242,N_13882);
nand U26194 (N_26194,N_19410,N_11250);
or U26195 (N_26195,N_10934,N_18672);
and U26196 (N_26196,N_15555,N_17473);
xor U26197 (N_26197,N_19513,N_14617);
and U26198 (N_26198,N_15130,N_16685);
nand U26199 (N_26199,N_18582,N_16825);
or U26200 (N_26200,N_10066,N_17493);
and U26201 (N_26201,N_12448,N_10986);
nand U26202 (N_26202,N_12206,N_19580);
nand U26203 (N_26203,N_17827,N_10830);
nand U26204 (N_26204,N_18420,N_14147);
nor U26205 (N_26205,N_12502,N_11351);
nand U26206 (N_26206,N_12192,N_18558);
and U26207 (N_26207,N_16942,N_12996);
and U26208 (N_26208,N_15935,N_15187);
and U26209 (N_26209,N_12261,N_19731);
nand U26210 (N_26210,N_15676,N_12824);
nor U26211 (N_26211,N_16861,N_10911);
and U26212 (N_26212,N_13402,N_10886);
nand U26213 (N_26213,N_10657,N_11584);
nor U26214 (N_26214,N_11349,N_12922);
or U26215 (N_26215,N_10664,N_18319);
or U26216 (N_26216,N_19724,N_13667);
or U26217 (N_26217,N_19268,N_16098);
nand U26218 (N_26218,N_11978,N_10305);
xor U26219 (N_26219,N_17439,N_17713);
and U26220 (N_26220,N_13527,N_11131);
and U26221 (N_26221,N_10877,N_13603);
and U26222 (N_26222,N_16675,N_10807);
nand U26223 (N_26223,N_17533,N_15069);
nor U26224 (N_26224,N_17550,N_12744);
nand U26225 (N_26225,N_16471,N_14684);
and U26226 (N_26226,N_18797,N_18394);
or U26227 (N_26227,N_13351,N_19087);
nand U26228 (N_26228,N_10478,N_17287);
nand U26229 (N_26229,N_15459,N_11481);
nand U26230 (N_26230,N_19227,N_11314);
or U26231 (N_26231,N_12847,N_17098);
nand U26232 (N_26232,N_18964,N_18338);
nand U26233 (N_26233,N_12523,N_10425);
or U26234 (N_26234,N_18138,N_12960);
nor U26235 (N_26235,N_14208,N_19859);
nand U26236 (N_26236,N_17420,N_17395);
and U26237 (N_26237,N_13269,N_12370);
or U26238 (N_26238,N_18089,N_14515);
or U26239 (N_26239,N_14828,N_12090);
nor U26240 (N_26240,N_18847,N_16199);
nor U26241 (N_26241,N_18181,N_10419);
or U26242 (N_26242,N_18631,N_17239);
and U26243 (N_26243,N_14091,N_10198);
nand U26244 (N_26244,N_14139,N_17986);
and U26245 (N_26245,N_14239,N_18262);
nor U26246 (N_26246,N_19275,N_14628);
or U26247 (N_26247,N_13649,N_10713);
xor U26248 (N_26248,N_15831,N_11433);
nor U26249 (N_26249,N_16099,N_12219);
and U26250 (N_26250,N_18747,N_17242);
nor U26251 (N_26251,N_10359,N_19620);
nor U26252 (N_26252,N_14323,N_11413);
or U26253 (N_26253,N_15114,N_15523);
or U26254 (N_26254,N_12323,N_16598);
or U26255 (N_26255,N_14376,N_11239);
or U26256 (N_26256,N_17795,N_19378);
and U26257 (N_26257,N_18846,N_16414);
nor U26258 (N_26258,N_18713,N_15605);
and U26259 (N_26259,N_10989,N_18713);
or U26260 (N_26260,N_12947,N_19046);
and U26261 (N_26261,N_14953,N_11792);
and U26262 (N_26262,N_12107,N_15737);
nor U26263 (N_26263,N_16888,N_19276);
nand U26264 (N_26264,N_15099,N_11045);
and U26265 (N_26265,N_14452,N_16562);
and U26266 (N_26266,N_17472,N_13667);
xnor U26267 (N_26267,N_15759,N_19166);
nand U26268 (N_26268,N_15870,N_11840);
nand U26269 (N_26269,N_15417,N_14247);
or U26270 (N_26270,N_19597,N_13046);
nor U26271 (N_26271,N_13501,N_18724);
and U26272 (N_26272,N_18453,N_19994);
or U26273 (N_26273,N_11240,N_13286);
or U26274 (N_26274,N_17291,N_18257);
xnor U26275 (N_26275,N_11599,N_10032);
nor U26276 (N_26276,N_14236,N_15741);
or U26277 (N_26277,N_14993,N_18491);
nand U26278 (N_26278,N_19704,N_19429);
nor U26279 (N_26279,N_16701,N_13789);
nor U26280 (N_26280,N_16747,N_19999);
or U26281 (N_26281,N_14869,N_14570);
or U26282 (N_26282,N_11356,N_19891);
xor U26283 (N_26283,N_16426,N_15526);
or U26284 (N_26284,N_17206,N_12213);
nor U26285 (N_26285,N_10771,N_12572);
nor U26286 (N_26286,N_13137,N_16308);
nand U26287 (N_26287,N_13861,N_17152);
or U26288 (N_26288,N_15310,N_10439);
or U26289 (N_26289,N_13968,N_15074);
and U26290 (N_26290,N_15033,N_13954);
and U26291 (N_26291,N_15725,N_12784);
nand U26292 (N_26292,N_15613,N_16570);
xnor U26293 (N_26293,N_12590,N_18034);
or U26294 (N_26294,N_17395,N_14222);
or U26295 (N_26295,N_15159,N_19455);
and U26296 (N_26296,N_12756,N_19670);
or U26297 (N_26297,N_13970,N_12038);
or U26298 (N_26298,N_18111,N_11797);
nor U26299 (N_26299,N_12848,N_12233);
nor U26300 (N_26300,N_18165,N_10426);
xor U26301 (N_26301,N_19877,N_18545);
and U26302 (N_26302,N_19677,N_12102);
or U26303 (N_26303,N_16698,N_17203);
or U26304 (N_26304,N_19043,N_11880);
nand U26305 (N_26305,N_19826,N_17309);
nand U26306 (N_26306,N_10228,N_17128);
nand U26307 (N_26307,N_16057,N_13959);
nor U26308 (N_26308,N_15285,N_15893);
or U26309 (N_26309,N_14538,N_14761);
or U26310 (N_26310,N_17186,N_15071);
nor U26311 (N_26311,N_12756,N_10629);
and U26312 (N_26312,N_15130,N_14125);
nand U26313 (N_26313,N_12743,N_14956);
nor U26314 (N_26314,N_15007,N_13896);
nor U26315 (N_26315,N_13436,N_15369);
nor U26316 (N_26316,N_10143,N_10835);
nor U26317 (N_26317,N_16005,N_10581);
nor U26318 (N_26318,N_14252,N_14679);
xnor U26319 (N_26319,N_11357,N_15545);
or U26320 (N_26320,N_11419,N_11197);
nor U26321 (N_26321,N_18410,N_18995);
nand U26322 (N_26322,N_16532,N_12995);
or U26323 (N_26323,N_11683,N_14107);
nor U26324 (N_26324,N_10070,N_19299);
or U26325 (N_26325,N_15528,N_14402);
xor U26326 (N_26326,N_19752,N_10172);
and U26327 (N_26327,N_15748,N_12948);
nor U26328 (N_26328,N_11188,N_11064);
nand U26329 (N_26329,N_19002,N_10727);
nand U26330 (N_26330,N_10697,N_12891);
nor U26331 (N_26331,N_11565,N_17814);
nor U26332 (N_26332,N_18607,N_18288);
nor U26333 (N_26333,N_19151,N_11215);
nand U26334 (N_26334,N_16734,N_19434);
and U26335 (N_26335,N_17118,N_18996);
xor U26336 (N_26336,N_13511,N_14515);
and U26337 (N_26337,N_13790,N_12822);
xnor U26338 (N_26338,N_13180,N_10574);
or U26339 (N_26339,N_12247,N_14094);
and U26340 (N_26340,N_12352,N_18029);
nand U26341 (N_26341,N_12624,N_12410);
xor U26342 (N_26342,N_13644,N_18628);
nand U26343 (N_26343,N_12980,N_18999);
and U26344 (N_26344,N_13424,N_17281);
nand U26345 (N_26345,N_18315,N_14855);
or U26346 (N_26346,N_14258,N_10436);
xnor U26347 (N_26347,N_13538,N_11281);
or U26348 (N_26348,N_13684,N_12344);
nand U26349 (N_26349,N_10833,N_14162);
and U26350 (N_26350,N_14199,N_15460);
and U26351 (N_26351,N_10651,N_14692);
nand U26352 (N_26352,N_15772,N_15094);
nand U26353 (N_26353,N_12558,N_19347);
and U26354 (N_26354,N_14450,N_11487);
xnor U26355 (N_26355,N_19735,N_18844);
or U26356 (N_26356,N_15899,N_13041);
xnor U26357 (N_26357,N_12730,N_10835);
nand U26358 (N_26358,N_17648,N_16324);
nor U26359 (N_26359,N_11237,N_15633);
and U26360 (N_26360,N_17658,N_13239);
nand U26361 (N_26361,N_17665,N_13314);
nand U26362 (N_26362,N_17168,N_13839);
nor U26363 (N_26363,N_15644,N_11650);
nand U26364 (N_26364,N_12432,N_15586);
or U26365 (N_26365,N_10803,N_12919);
xor U26366 (N_26366,N_19041,N_12074);
or U26367 (N_26367,N_12742,N_17397);
nor U26368 (N_26368,N_12662,N_17446);
nor U26369 (N_26369,N_17654,N_18574);
nor U26370 (N_26370,N_14709,N_14063);
and U26371 (N_26371,N_13078,N_12261);
and U26372 (N_26372,N_12157,N_12130);
and U26373 (N_26373,N_10853,N_19236);
and U26374 (N_26374,N_16070,N_15680);
or U26375 (N_26375,N_14733,N_18885);
and U26376 (N_26376,N_18117,N_10177);
nand U26377 (N_26377,N_19150,N_15571);
nor U26378 (N_26378,N_12666,N_12817);
nand U26379 (N_26379,N_14687,N_14856);
nor U26380 (N_26380,N_17393,N_13631);
and U26381 (N_26381,N_10749,N_17797);
xor U26382 (N_26382,N_15977,N_13804);
nor U26383 (N_26383,N_18527,N_19491);
and U26384 (N_26384,N_13190,N_14834);
or U26385 (N_26385,N_14877,N_15873);
or U26386 (N_26386,N_19451,N_18221);
or U26387 (N_26387,N_10129,N_15165);
nand U26388 (N_26388,N_13928,N_10832);
nor U26389 (N_26389,N_17731,N_15165);
xnor U26390 (N_26390,N_14890,N_17206);
or U26391 (N_26391,N_14490,N_11253);
xnor U26392 (N_26392,N_17583,N_11709);
or U26393 (N_26393,N_15990,N_18981);
and U26394 (N_26394,N_16556,N_17045);
and U26395 (N_26395,N_12157,N_18497);
nor U26396 (N_26396,N_14244,N_16819);
nand U26397 (N_26397,N_10276,N_11957);
or U26398 (N_26398,N_18314,N_17210);
nand U26399 (N_26399,N_16765,N_15635);
nand U26400 (N_26400,N_16529,N_16785);
nand U26401 (N_26401,N_12702,N_17652);
and U26402 (N_26402,N_16578,N_12827);
nand U26403 (N_26403,N_10607,N_12191);
and U26404 (N_26404,N_15257,N_15193);
or U26405 (N_26405,N_14095,N_14812);
and U26406 (N_26406,N_10329,N_11499);
or U26407 (N_26407,N_17919,N_14183);
nand U26408 (N_26408,N_12354,N_15090);
and U26409 (N_26409,N_19227,N_13266);
xnor U26410 (N_26410,N_17929,N_10988);
or U26411 (N_26411,N_16237,N_19178);
xor U26412 (N_26412,N_16080,N_18122);
xor U26413 (N_26413,N_12635,N_13633);
and U26414 (N_26414,N_19947,N_16921);
or U26415 (N_26415,N_14948,N_13946);
xnor U26416 (N_26416,N_14153,N_10858);
nand U26417 (N_26417,N_17233,N_13980);
or U26418 (N_26418,N_10709,N_11315);
nand U26419 (N_26419,N_11659,N_14854);
nand U26420 (N_26420,N_18573,N_11098);
nand U26421 (N_26421,N_11145,N_12598);
nor U26422 (N_26422,N_13761,N_18016);
nor U26423 (N_26423,N_10292,N_19622);
nor U26424 (N_26424,N_14500,N_18241);
xor U26425 (N_26425,N_18833,N_11391);
nand U26426 (N_26426,N_13872,N_14086);
and U26427 (N_26427,N_10736,N_12777);
or U26428 (N_26428,N_14229,N_12437);
and U26429 (N_26429,N_15441,N_13304);
nor U26430 (N_26430,N_19608,N_10757);
nand U26431 (N_26431,N_18942,N_18368);
xor U26432 (N_26432,N_18599,N_12000);
nand U26433 (N_26433,N_19306,N_14956);
or U26434 (N_26434,N_12959,N_17429);
nand U26435 (N_26435,N_10867,N_19969);
and U26436 (N_26436,N_18112,N_16445);
and U26437 (N_26437,N_16427,N_10743);
or U26438 (N_26438,N_12238,N_18671);
and U26439 (N_26439,N_13590,N_10016);
and U26440 (N_26440,N_11477,N_18097);
and U26441 (N_26441,N_17200,N_17501);
or U26442 (N_26442,N_13019,N_17778);
nand U26443 (N_26443,N_15816,N_14006);
and U26444 (N_26444,N_12564,N_10115);
and U26445 (N_26445,N_11370,N_14441);
xnor U26446 (N_26446,N_15923,N_19490);
or U26447 (N_26447,N_19565,N_11377);
and U26448 (N_26448,N_14419,N_18283);
xor U26449 (N_26449,N_13480,N_15376);
xnor U26450 (N_26450,N_18194,N_11260);
nand U26451 (N_26451,N_10440,N_12943);
or U26452 (N_26452,N_17250,N_10482);
nor U26453 (N_26453,N_19552,N_18454);
nand U26454 (N_26454,N_17234,N_14590);
or U26455 (N_26455,N_17925,N_10489);
or U26456 (N_26456,N_18520,N_17815);
or U26457 (N_26457,N_16230,N_11982);
nor U26458 (N_26458,N_16638,N_13459);
and U26459 (N_26459,N_18061,N_16026);
and U26460 (N_26460,N_15587,N_19088);
xnor U26461 (N_26461,N_16065,N_19894);
or U26462 (N_26462,N_19502,N_19393);
nor U26463 (N_26463,N_15525,N_19066);
nor U26464 (N_26464,N_18850,N_12665);
or U26465 (N_26465,N_18591,N_14101);
nor U26466 (N_26466,N_18410,N_16352);
or U26467 (N_26467,N_15973,N_12605);
or U26468 (N_26468,N_15302,N_15226);
nor U26469 (N_26469,N_10569,N_17172);
nor U26470 (N_26470,N_17118,N_19370);
and U26471 (N_26471,N_18000,N_18873);
or U26472 (N_26472,N_18844,N_12893);
xnor U26473 (N_26473,N_11863,N_12529);
and U26474 (N_26474,N_12153,N_19821);
and U26475 (N_26475,N_11888,N_14197);
nor U26476 (N_26476,N_18711,N_11226);
or U26477 (N_26477,N_17261,N_11224);
and U26478 (N_26478,N_13929,N_14014);
nand U26479 (N_26479,N_15769,N_18469);
or U26480 (N_26480,N_17239,N_15350);
nor U26481 (N_26481,N_16004,N_12716);
and U26482 (N_26482,N_14072,N_16686);
xor U26483 (N_26483,N_11432,N_15304);
nand U26484 (N_26484,N_10670,N_17175);
xor U26485 (N_26485,N_17400,N_19595);
and U26486 (N_26486,N_17691,N_18412);
nor U26487 (N_26487,N_13269,N_14563);
nor U26488 (N_26488,N_10359,N_18059);
nor U26489 (N_26489,N_16335,N_17394);
xnor U26490 (N_26490,N_18162,N_12359);
and U26491 (N_26491,N_16476,N_18274);
nor U26492 (N_26492,N_19954,N_17663);
nor U26493 (N_26493,N_15820,N_16555);
or U26494 (N_26494,N_19362,N_13417);
or U26495 (N_26495,N_12176,N_13737);
nor U26496 (N_26496,N_17206,N_13656);
nand U26497 (N_26497,N_12894,N_14221);
nand U26498 (N_26498,N_12060,N_16581);
and U26499 (N_26499,N_11302,N_18427);
xor U26500 (N_26500,N_18541,N_12726);
and U26501 (N_26501,N_15953,N_16745);
or U26502 (N_26502,N_19681,N_12343);
xnor U26503 (N_26503,N_18629,N_14434);
and U26504 (N_26504,N_19991,N_18633);
nor U26505 (N_26505,N_14104,N_12497);
xor U26506 (N_26506,N_11357,N_19334);
and U26507 (N_26507,N_11553,N_13458);
nand U26508 (N_26508,N_16650,N_11276);
nor U26509 (N_26509,N_14316,N_18595);
nand U26510 (N_26510,N_10896,N_16424);
nand U26511 (N_26511,N_11728,N_13881);
nor U26512 (N_26512,N_15926,N_10373);
nor U26513 (N_26513,N_15364,N_18105);
or U26514 (N_26514,N_13338,N_16438);
nand U26515 (N_26515,N_13446,N_17517);
nand U26516 (N_26516,N_14705,N_15727);
nand U26517 (N_26517,N_14284,N_12603);
and U26518 (N_26518,N_10891,N_19632);
xnor U26519 (N_26519,N_18990,N_12373);
and U26520 (N_26520,N_16228,N_10731);
nand U26521 (N_26521,N_13439,N_15760);
and U26522 (N_26522,N_19213,N_15746);
nand U26523 (N_26523,N_11498,N_14697);
nand U26524 (N_26524,N_14938,N_12198);
nor U26525 (N_26525,N_13397,N_10428);
nor U26526 (N_26526,N_11449,N_15973);
or U26527 (N_26527,N_12558,N_10021);
nand U26528 (N_26528,N_18933,N_18985);
nor U26529 (N_26529,N_18819,N_10612);
nor U26530 (N_26530,N_18290,N_10889);
nor U26531 (N_26531,N_12353,N_18408);
nand U26532 (N_26532,N_14453,N_11984);
nand U26533 (N_26533,N_12722,N_11114);
and U26534 (N_26534,N_17754,N_19503);
and U26535 (N_26535,N_15329,N_16059);
nor U26536 (N_26536,N_12264,N_18470);
and U26537 (N_26537,N_13869,N_14611);
or U26538 (N_26538,N_18772,N_14890);
or U26539 (N_26539,N_15482,N_19926);
and U26540 (N_26540,N_11096,N_16159);
nor U26541 (N_26541,N_18326,N_12235);
and U26542 (N_26542,N_19375,N_11927);
or U26543 (N_26543,N_16229,N_15899);
and U26544 (N_26544,N_11881,N_12754);
and U26545 (N_26545,N_12044,N_15072);
nand U26546 (N_26546,N_10465,N_14891);
nor U26547 (N_26547,N_13503,N_10708);
and U26548 (N_26548,N_19006,N_15100);
or U26549 (N_26549,N_13022,N_14283);
nor U26550 (N_26550,N_18881,N_13604);
nand U26551 (N_26551,N_19617,N_12174);
nand U26552 (N_26552,N_15737,N_13545);
nor U26553 (N_26553,N_10089,N_13452);
and U26554 (N_26554,N_11722,N_17073);
xor U26555 (N_26555,N_14497,N_16455);
or U26556 (N_26556,N_13528,N_15629);
nor U26557 (N_26557,N_17452,N_14976);
and U26558 (N_26558,N_11180,N_18318);
and U26559 (N_26559,N_17653,N_19867);
and U26560 (N_26560,N_15802,N_10016);
or U26561 (N_26561,N_14579,N_14256);
or U26562 (N_26562,N_11188,N_10349);
and U26563 (N_26563,N_13146,N_16542);
nor U26564 (N_26564,N_15455,N_19032);
or U26565 (N_26565,N_10158,N_19505);
nand U26566 (N_26566,N_16125,N_16637);
and U26567 (N_26567,N_19289,N_17106);
nand U26568 (N_26568,N_10548,N_18332);
or U26569 (N_26569,N_18350,N_12905);
nor U26570 (N_26570,N_16824,N_14980);
nor U26571 (N_26571,N_19586,N_10452);
and U26572 (N_26572,N_19457,N_10025);
or U26573 (N_26573,N_12973,N_12468);
or U26574 (N_26574,N_16410,N_15531);
or U26575 (N_26575,N_12420,N_11761);
nand U26576 (N_26576,N_15415,N_17592);
nor U26577 (N_26577,N_13727,N_17909);
and U26578 (N_26578,N_14727,N_11499);
nand U26579 (N_26579,N_15257,N_14652);
or U26580 (N_26580,N_16863,N_11631);
and U26581 (N_26581,N_14615,N_10645);
nor U26582 (N_26582,N_15497,N_10024);
nor U26583 (N_26583,N_10188,N_11193);
xor U26584 (N_26584,N_17253,N_18674);
nor U26585 (N_26585,N_13500,N_16782);
nor U26586 (N_26586,N_13661,N_13444);
nand U26587 (N_26587,N_18433,N_18794);
or U26588 (N_26588,N_12312,N_17086);
or U26589 (N_26589,N_14311,N_12973);
nand U26590 (N_26590,N_15944,N_13587);
and U26591 (N_26591,N_19037,N_15812);
nand U26592 (N_26592,N_18565,N_14813);
and U26593 (N_26593,N_13988,N_10100);
nand U26594 (N_26594,N_12418,N_19341);
nor U26595 (N_26595,N_18650,N_10773);
and U26596 (N_26596,N_19213,N_18592);
or U26597 (N_26597,N_19010,N_11309);
nand U26598 (N_26598,N_16209,N_13432);
and U26599 (N_26599,N_13624,N_14052);
nor U26600 (N_26600,N_11976,N_15777);
or U26601 (N_26601,N_19366,N_14522);
nand U26602 (N_26602,N_11702,N_17661);
nor U26603 (N_26603,N_15662,N_19442);
and U26604 (N_26604,N_10979,N_12588);
and U26605 (N_26605,N_12490,N_13063);
nand U26606 (N_26606,N_14221,N_13666);
and U26607 (N_26607,N_11599,N_19461);
nor U26608 (N_26608,N_10918,N_11989);
and U26609 (N_26609,N_19080,N_13524);
or U26610 (N_26610,N_13359,N_11611);
or U26611 (N_26611,N_12528,N_10839);
nand U26612 (N_26612,N_18984,N_14075);
and U26613 (N_26613,N_19840,N_16538);
and U26614 (N_26614,N_17466,N_17314);
or U26615 (N_26615,N_17748,N_17265);
or U26616 (N_26616,N_19296,N_16142);
nand U26617 (N_26617,N_12983,N_16051);
nor U26618 (N_26618,N_11428,N_19227);
nand U26619 (N_26619,N_12065,N_18670);
nand U26620 (N_26620,N_11194,N_17496);
nand U26621 (N_26621,N_10836,N_17576);
and U26622 (N_26622,N_13098,N_11014);
or U26623 (N_26623,N_15862,N_12567);
or U26624 (N_26624,N_10749,N_15191);
nor U26625 (N_26625,N_17578,N_16487);
and U26626 (N_26626,N_15700,N_15817);
and U26627 (N_26627,N_10828,N_18711);
nor U26628 (N_26628,N_10117,N_18587);
or U26629 (N_26629,N_12192,N_15888);
nor U26630 (N_26630,N_19076,N_16141);
or U26631 (N_26631,N_16391,N_16199);
and U26632 (N_26632,N_10886,N_17027);
nor U26633 (N_26633,N_18621,N_18246);
nor U26634 (N_26634,N_11389,N_15970);
or U26635 (N_26635,N_17898,N_12888);
nor U26636 (N_26636,N_19316,N_12654);
or U26637 (N_26637,N_19868,N_13800);
xnor U26638 (N_26638,N_17212,N_16521);
xnor U26639 (N_26639,N_18026,N_12242);
nor U26640 (N_26640,N_11076,N_16110);
xor U26641 (N_26641,N_13690,N_19723);
nor U26642 (N_26642,N_10226,N_10392);
or U26643 (N_26643,N_11006,N_11947);
or U26644 (N_26644,N_13606,N_18072);
or U26645 (N_26645,N_19133,N_13206);
nand U26646 (N_26646,N_13963,N_16574);
and U26647 (N_26647,N_19577,N_18681);
nor U26648 (N_26648,N_11574,N_14840);
and U26649 (N_26649,N_18981,N_19499);
xnor U26650 (N_26650,N_12560,N_19288);
xnor U26651 (N_26651,N_17162,N_11649);
nor U26652 (N_26652,N_17012,N_10631);
and U26653 (N_26653,N_18435,N_11227);
or U26654 (N_26654,N_14875,N_12342);
and U26655 (N_26655,N_12418,N_17435);
nand U26656 (N_26656,N_19916,N_12860);
or U26657 (N_26657,N_12296,N_10117);
and U26658 (N_26658,N_12662,N_15591);
xor U26659 (N_26659,N_10999,N_13254);
or U26660 (N_26660,N_18401,N_12574);
nand U26661 (N_26661,N_19157,N_13354);
nand U26662 (N_26662,N_14273,N_11424);
and U26663 (N_26663,N_10869,N_14067);
nor U26664 (N_26664,N_12148,N_11764);
nor U26665 (N_26665,N_16921,N_14899);
nor U26666 (N_26666,N_11919,N_17925);
and U26667 (N_26667,N_11693,N_14059);
nor U26668 (N_26668,N_18202,N_16064);
and U26669 (N_26669,N_13981,N_12583);
and U26670 (N_26670,N_18356,N_17165);
nand U26671 (N_26671,N_17433,N_18749);
or U26672 (N_26672,N_11583,N_12939);
nand U26673 (N_26673,N_10738,N_19403);
or U26674 (N_26674,N_16507,N_13313);
xor U26675 (N_26675,N_14147,N_10598);
nor U26676 (N_26676,N_14543,N_17173);
nor U26677 (N_26677,N_10183,N_19892);
or U26678 (N_26678,N_16043,N_11416);
and U26679 (N_26679,N_15571,N_13422);
nand U26680 (N_26680,N_16751,N_13754);
or U26681 (N_26681,N_19963,N_11452);
nor U26682 (N_26682,N_17475,N_12026);
or U26683 (N_26683,N_11845,N_14160);
or U26684 (N_26684,N_16448,N_18719);
or U26685 (N_26685,N_18677,N_18807);
xnor U26686 (N_26686,N_13990,N_12640);
nor U26687 (N_26687,N_12862,N_17409);
or U26688 (N_26688,N_14445,N_14870);
or U26689 (N_26689,N_17865,N_13752);
xor U26690 (N_26690,N_11893,N_10341);
nand U26691 (N_26691,N_11164,N_12319);
nor U26692 (N_26692,N_13199,N_17988);
nor U26693 (N_26693,N_12497,N_17903);
nor U26694 (N_26694,N_18351,N_16796);
nand U26695 (N_26695,N_12818,N_15761);
and U26696 (N_26696,N_17319,N_16566);
and U26697 (N_26697,N_10943,N_11628);
nor U26698 (N_26698,N_11732,N_16190);
nor U26699 (N_26699,N_12757,N_18982);
nand U26700 (N_26700,N_19713,N_12091);
nor U26701 (N_26701,N_14271,N_12722);
or U26702 (N_26702,N_17843,N_18033);
nor U26703 (N_26703,N_10415,N_16625);
nor U26704 (N_26704,N_18890,N_18431);
or U26705 (N_26705,N_14356,N_17788);
xnor U26706 (N_26706,N_19709,N_16524);
nor U26707 (N_26707,N_11268,N_19546);
nand U26708 (N_26708,N_14149,N_17778);
nor U26709 (N_26709,N_13464,N_16291);
and U26710 (N_26710,N_13767,N_14046);
nand U26711 (N_26711,N_14173,N_16312);
nor U26712 (N_26712,N_16596,N_19191);
or U26713 (N_26713,N_18145,N_17125);
nand U26714 (N_26714,N_16195,N_12989);
and U26715 (N_26715,N_11583,N_19886);
nor U26716 (N_26716,N_10398,N_11948);
and U26717 (N_26717,N_16905,N_15132);
or U26718 (N_26718,N_15620,N_11808);
nand U26719 (N_26719,N_14400,N_14308);
nor U26720 (N_26720,N_19536,N_11546);
or U26721 (N_26721,N_15291,N_12938);
or U26722 (N_26722,N_11428,N_13956);
and U26723 (N_26723,N_10488,N_10038);
xor U26724 (N_26724,N_19517,N_16537);
and U26725 (N_26725,N_17915,N_16516);
nor U26726 (N_26726,N_18720,N_17789);
nor U26727 (N_26727,N_14859,N_12927);
nand U26728 (N_26728,N_14870,N_18923);
nor U26729 (N_26729,N_14908,N_18526);
or U26730 (N_26730,N_19807,N_18370);
xor U26731 (N_26731,N_11539,N_12851);
or U26732 (N_26732,N_11228,N_19669);
xnor U26733 (N_26733,N_11018,N_10972);
and U26734 (N_26734,N_16778,N_11342);
and U26735 (N_26735,N_16146,N_12262);
and U26736 (N_26736,N_17821,N_11077);
nand U26737 (N_26737,N_15680,N_17108);
nand U26738 (N_26738,N_17194,N_18780);
nor U26739 (N_26739,N_14060,N_19501);
nand U26740 (N_26740,N_17842,N_19904);
or U26741 (N_26741,N_15361,N_10772);
xor U26742 (N_26742,N_10866,N_19334);
nor U26743 (N_26743,N_14234,N_10274);
and U26744 (N_26744,N_12438,N_12795);
xnor U26745 (N_26745,N_16197,N_12370);
or U26746 (N_26746,N_17222,N_10899);
nand U26747 (N_26747,N_18244,N_16030);
nand U26748 (N_26748,N_16031,N_17138);
or U26749 (N_26749,N_14169,N_14637);
nor U26750 (N_26750,N_11623,N_11474);
xnor U26751 (N_26751,N_17190,N_15108);
nor U26752 (N_26752,N_10368,N_14442);
and U26753 (N_26753,N_14844,N_11118);
nor U26754 (N_26754,N_16455,N_14163);
nand U26755 (N_26755,N_15219,N_11181);
nand U26756 (N_26756,N_19801,N_12215);
and U26757 (N_26757,N_18587,N_10851);
nor U26758 (N_26758,N_19503,N_17261);
nor U26759 (N_26759,N_15842,N_19409);
or U26760 (N_26760,N_11548,N_16534);
or U26761 (N_26761,N_14983,N_19932);
and U26762 (N_26762,N_14758,N_15361);
nand U26763 (N_26763,N_17924,N_10736);
and U26764 (N_26764,N_19776,N_11194);
nor U26765 (N_26765,N_17530,N_17305);
and U26766 (N_26766,N_14378,N_16872);
and U26767 (N_26767,N_16452,N_14200);
and U26768 (N_26768,N_14124,N_12665);
and U26769 (N_26769,N_18508,N_17186);
and U26770 (N_26770,N_12201,N_10939);
xor U26771 (N_26771,N_14946,N_17061);
xor U26772 (N_26772,N_10783,N_10092);
nor U26773 (N_26773,N_18015,N_11471);
and U26774 (N_26774,N_14825,N_12954);
nand U26775 (N_26775,N_12393,N_10688);
nand U26776 (N_26776,N_14990,N_17275);
nor U26777 (N_26777,N_18203,N_11943);
and U26778 (N_26778,N_19769,N_16913);
nor U26779 (N_26779,N_17752,N_15807);
or U26780 (N_26780,N_10291,N_15259);
nand U26781 (N_26781,N_12742,N_10989);
and U26782 (N_26782,N_11855,N_15619);
nor U26783 (N_26783,N_17132,N_11328);
nor U26784 (N_26784,N_11187,N_18090);
xnor U26785 (N_26785,N_15458,N_13849);
nor U26786 (N_26786,N_17563,N_16138);
and U26787 (N_26787,N_19560,N_15096);
and U26788 (N_26788,N_11542,N_17206);
and U26789 (N_26789,N_13805,N_13290);
or U26790 (N_26790,N_10498,N_13427);
and U26791 (N_26791,N_19028,N_14351);
nor U26792 (N_26792,N_12371,N_13085);
and U26793 (N_26793,N_13560,N_13127);
xor U26794 (N_26794,N_19674,N_15233);
nand U26795 (N_26795,N_15976,N_15538);
nand U26796 (N_26796,N_13416,N_14927);
and U26797 (N_26797,N_11382,N_12856);
and U26798 (N_26798,N_10026,N_15578);
and U26799 (N_26799,N_19531,N_11968);
nor U26800 (N_26800,N_13260,N_10728);
nand U26801 (N_26801,N_10309,N_19090);
xor U26802 (N_26802,N_16078,N_13421);
and U26803 (N_26803,N_19957,N_16978);
nor U26804 (N_26804,N_10981,N_11507);
and U26805 (N_26805,N_14190,N_11494);
and U26806 (N_26806,N_12941,N_14994);
nor U26807 (N_26807,N_10575,N_16448);
and U26808 (N_26808,N_12179,N_13201);
and U26809 (N_26809,N_12107,N_17880);
or U26810 (N_26810,N_15053,N_13090);
or U26811 (N_26811,N_18894,N_17589);
xnor U26812 (N_26812,N_10255,N_16360);
or U26813 (N_26813,N_11663,N_15929);
and U26814 (N_26814,N_11783,N_11004);
or U26815 (N_26815,N_12135,N_15399);
or U26816 (N_26816,N_18014,N_16411);
nor U26817 (N_26817,N_10425,N_17593);
nor U26818 (N_26818,N_19236,N_10674);
or U26819 (N_26819,N_16184,N_16224);
or U26820 (N_26820,N_14118,N_13355);
nand U26821 (N_26821,N_10349,N_18065);
xor U26822 (N_26822,N_14927,N_18228);
and U26823 (N_26823,N_18745,N_12351);
nor U26824 (N_26824,N_14428,N_17160);
nor U26825 (N_26825,N_18121,N_16869);
nand U26826 (N_26826,N_12298,N_16780);
nand U26827 (N_26827,N_14744,N_12945);
nand U26828 (N_26828,N_12950,N_19645);
nand U26829 (N_26829,N_15994,N_15201);
and U26830 (N_26830,N_14761,N_11027);
xor U26831 (N_26831,N_15341,N_10930);
nand U26832 (N_26832,N_13598,N_18706);
nor U26833 (N_26833,N_12566,N_18467);
xnor U26834 (N_26834,N_15229,N_11858);
nor U26835 (N_26835,N_18168,N_16710);
nand U26836 (N_26836,N_17581,N_14904);
nand U26837 (N_26837,N_15696,N_13560);
nand U26838 (N_26838,N_18564,N_19903);
or U26839 (N_26839,N_13648,N_15449);
or U26840 (N_26840,N_17911,N_14261);
or U26841 (N_26841,N_19023,N_19070);
nand U26842 (N_26842,N_19222,N_17559);
nor U26843 (N_26843,N_10258,N_18331);
or U26844 (N_26844,N_17403,N_18621);
nand U26845 (N_26845,N_10359,N_17568);
nor U26846 (N_26846,N_16622,N_18220);
and U26847 (N_26847,N_19245,N_12061);
and U26848 (N_26848,N_12317,N_12167);
or U26849 (N_26849,N_11938,N_17557);
xor U26850 (N_26850,N_19670,N_17909);
or U26851 (N_26851,N_17510,N_16288);
or U26852 (N_26852,N_15000,N_15633);
xnor U26853 (N_26853,N_10264,N_18036);
and U26854 (N_26854,N_10085,N_11551);
nor U26855 (N_26855,N_13685,N_11385);
or U26856 (N_26856,N_15325,N_12179);
or U26857 (N_26857,N_17584,N_18400);
nor U26858 (N_26858,N_14654,N_19681);
nor U26859 (N_26859,N_19938,N_10570);
nand U26860 (N_26860,N_19230,N_13016);
or U26861 (N_26861,N_18339,N_18135);
or U26862 (N_26862,N_10381,N_15426);
and U26863 (N_26863,N_15132,N_15838);
or U26864 (N_26864,N_17730,N_13927);
nor U26865 (N_26865,N_11644,N_12529);
nor U26866 (N_26866,N_14804,N_10325);
or U26867 (N_26867,N_14285,N_13445);
nor U26868 (N_26868,N_11853,N_11159);
and U26869 (N_26869,N_17241,N_17236);
nand U26870 (N_26870,N_13709,N_11009);
xnor U26871 (N_26871,N_18987,N_16121);
nand U26872 (N_26872,N_17475,N_13157);
or U26873 (N_26873,N_10106,N_14359);
nand U26874 (N_26874,N_15036,N_18454);
or U26875 (N_26875,N_18253,N_16224);
nor U26876 (N_26876,N_14797,N_11052);
nand U26877 (N_26877,N_17008,N_17907);
and U26878 (N_26878,N_16045,N_11528);
xnor U26879 (N_26879,N_19753,N_18823);
nor U26880 (N_26880,N_13014,N_16104);
or U26881 (N_26881,N_16059,N_11972);
xnor U26882 (N_26882,N_13573,N_11049);
or U26883 (N_26883,N_15532,N_10446);
nand U26884 (N_26884,N_17639,N_13623);
and U26885 (N_26885,N_11036,N_11758);
and U26886 (N_26886,N_10443,N_14652);
nand U26887 (N_26887,N_14642,N_10361);
nand U26888 (N_26888,N_19441,N_12378);
xor U26889 (N_26889,N_17607,N_10317);
or U26890 (N_26890,N_10213,N_12332);
nand U26891 (N_26891,N_16659,N_19097);
nand U26892 (N_26892,N_10438,N_18074);
or U26893 (N_26893,N_17259,N_19666);
or U26894 (N_26894,N_18350,N_16792);
or U26895 (N_26895,N_16864,N_12971);
and U26896 (N_26896,N_17219,N_18396);
or U26897 (N_26897,N_11731,N_19321);
and U26898 (N_26898,N_19794,N_16028);
nor U26899 (N_26899,N_12920,N_15470);
nor U26900 (N_26900,N_17391,N_19151);
and U26901 (N_26901,N_17806,N_14941);
nand U26902 (N_26902,N_17972,N_19947);
nor U26903 (N_26903,N_10524,N_10668);
and U26904 (N_26904,N_18509,N_14447);
or U26905 (N_26905,N_17128,N_15346);
nand U26906 (N_26906,N_19466,N_16327);
nand U26907 (N_26907,N_14510,N_11734);
nand U26908 (N_26908,N_17606,N_14899);
or U26909 (N_26909,N_13499,N_11690);
nor U26910 (N_26910,N_16130,N_14334);
xor U26911 (N_26911,N_16382,N_13894);
and U26912 (N_26912,N_10687,N_18382);
or U26913 (N_26913,N_15219,N_14145);
and U26914 (N_26914,N_18733,N_15674);
nand U26915 (N_26915,N_12827,N_17661);
nand U26916 (N_26916,N_10765,N_14993);
nand U26917 (N_26917,N_13791,N_15327);
or U26918 (N_26918,N_15996,N_16112);
nor U26919 (N_26919,N_17641,N_15597);
xor U26920 (N_26920,N_11764,N_19967);
nand U26921 (N_26921,N_10717,N_17278);
nor U26922 (N_26922,N_12351,N_18633);
nor U26923 (N_26923,N_17268,N_13409);
or U26924 (N_26924,N_10334,N_17077);
nor U26925 (N_26925,N_14026,N_17123);
or U26926 (N_26926,N_14725,N_13645);
nor U26927 (N_26927,N_19388,N_12318);
nor U26928 (N_26928,N_19487,N_10269);
and U26929 (N_26929,N_16747,N_16243);
nand U26930 (N_26930,N_17733,N_10685);
xnor U26931 (N_26931,N_10589,N_14508);
xnor U26932 (N_26932,N_14593,N_19999);
or U26933 (N_26933,N_17190,N_12858);
nand U26934 (N_26934,N_12124,N_10984);
and U26935 (N_26935,N_11900,N_16908);
nand U26936 (N_26936,N_18085,N_10764);
nor U26937 (N_26937,N_15768,N_13339);
nand U26938 (N_26938,N_15768,N_15136);
nor U26939 (N_26939,N_19691,N_12292);
or U26940 (N_26940,N_12096,N_16851);
nand U26941 (N_26941,N_17385,N_14836);
and U26942 (N_26942,N_18729,N_13678);
or U26943 (N_26943,N_15608,N_12552);
nand U26944 (N_26944,N_15335,N_17906);
nor U26945 (N_26945,N_18950,N_19445);
or U26946 (N_26946,N_19015,N_14752);
nand U26947 (N_26947,N_11433,N_15593);
nand U26948 (N_26948,N_11925,N_11374);
or U26949 (N_26949,N_18935,N_18686);
or U26950 (N_26950,N_16757,N_13008);
nand U26951 (N_26951,N_11885,N_15586);
or U26952 (N_26952,N_14268,N_13339);
nand U26953 (N_26953,N_14614,N_14343);
and U26954 (N_26954,N_19973,N_12967);
nor U26955 (N_26955,N_16888,N_15069);
xor U26956 (N_26956,N_18789,N_16767);
xnor U26957 (N_26957,N_12351,N_12634);
nor U26958 (N_26958,N_10381,N_12827);
nand U26959 (N_26959,N_13070,N_12924);
nor U26960 (N_26960,N_10987,N_18602);
and U26961 (N_26961,N_19360,N_11770);
or U26962 (N_26962,N_15345,N_18861);
nand U26963 (N_26963,N_16330,N_13326);
or U26964 (N_26964,N_13700,N_11958);
and U26965 (N_26965,N_17920,N_13713);
nor U26966 (N_26966,N_12795,N_14136);
and U26967 (N_26967,N_15217,N_18644);
or U26968 (N_26968,N_15873,N_12339);
and U26969 (N_26969,N_12527,N_16911);
or U26970 (N_26970,N_17130,N_19251);
nand U26971 (N_26971,N_11602,N_14980);
nor U26972 (N_26972,N_15043,N_10488);
and U26973 (N_26973,N_17124,N_13783);
or U26974 (N_26974,N_11985,N_16403);
and U26975 (N_26975,N_11573,N_19014);
or U26976 (N_26976,N_14354,N_12980);
nor U26977 (N_26977,N_10118,N_14062);
or U26978 (N_26978,N_19004,N_10936);
or U26979 (N_26979,N_18086,N_14010);
xnor U26980 (N_26980,N_18538,N_18726);
and U26981 (N_26981,N_17362,N_18630);
and U26982 (N_26982,N_12430,N_15893);
nand U26983 (N_26983,N_10390,N_16823);
and U26984 (N_26984,N_13505,N_17956);
nor U26985 (N_26985,N_12853,N_10083);
or U26986 (N_26986,N_19098,N_17468);
nand U26987 (N_26987,N_10016,N_19836);
nand U26988 (N_26988,N_10121,N_15427);
or U26989 (N_26989,N_19923,N_19243);
and U26990 (N_26990,N_19302,N_17894);
and U26991 (N_26991,N_10853,N_11171);
and U26992 (N_26992,N_10580,N_16390);
nand U26993 (N_26993,N_16786,N_18169);
nor U26994 (N_26994,N_16130,N_11421);
and U26995 (N_26995,N_11301,N_17585);
nor U26996 (N_26996,N_10520,N_11990);
nand U26997 (N_26997,N_16785,N_16548);
or U26998 (N_26998,N_18117,N_18550);
nor U26999 (N_26999,N_11436,N_12360);
nor U27000 (N_27000,N_18532,N_15515);
or U27001 (N_27001,N_13834,N_10879);
or U27002 (N_27002,N_12792,N_18035);
or U27003 (N_27003,N_10297,N_12901);
and U27004 (N_27004,N_10748,N_10190);
and U27005 (N_27005,N_14670,N_19513);
nand U27006 (N_27006,N_10343,N_15573);
nand U27007 (N_27007,N_12823,N_13939);
nand U27008 (N_27008,N_12874,N_10261);
nand U27009 (N_27009,N_12203,N_19899);
or U27010 (N_27010,N_15765,N_15768);
and U27011 (N_27011,N_14246,N_18266);
or U27012 (N_27012,N_15490,N_19669);
nand U27013 (N_27013,N_11124,N_19624);
or U27014 (N_27014,N_16065,N_15397);
nand U27015 (N_27015,N_15413,N_11108);
or U27016 (N_27016,N_11833,N_19517);
and U27017 (N_27017,N_19008,N_11017);
or U27018 (N_27018,N_17905,N_12303);
and U27019 (N_27019,N_13341,N_17159);
xnor U27020 (N_27020,N_17796,N_17310);
nand U27021 (N_27021,N_19415,N_17800);
or U27022 (N_27022,N_13195,N_15873);
nand U27023 (N_27023,N_17805,N_16047);
or U27024 (N_27024,N_10311,N_10656);
and U27025 (N_27025,N_19380,N_16035);
nor U27026 (N_27026,N_10041,N_13017);
nor U27027 (N_27027,N_17045,N_12928);
nor U27028 (N_27028,N_17984,N_15812);
nor U27029 (N_27029,N_13144,N_11856);
nor U27030 (N_27030,N_10921,N_18840);
nor U27031 (N_27031,N_11003,N_10589);
and U27032 (N_27032,N_15352,N_14567);
nand U27033 (N_27033,N_17925,N_13141);
nor U27034 (N_27034,N_16499,N_13595);
nand U27035 (N_27035,N_19876,N_11977);
nor U27036 (N_27036,N_11599,N_19071);
nand U27037 (N_27037,N_12980,N_19437);
nor U27038 (N_27038,N_13515,N_12183);
nand U27039 (N_27039,N_18708,N_19712);
and U27040 (N_27040,N_15537,N_16692);
or U27041 (N_27041,N_10783,N_13191);
and U27042 (N_27042,N_14994,N_18132);
and U27043 (N_27043,N_14135,N_19186);
and U27044 (N_27044,N_19801,N_12874);
nand U27045 (N_27045,N_11494,N_10752);
nor U27046 (N_27046,N_17088,N_11910);
nand U27047 (N_27047,N_10934,N_12719);
or U27048 (N_27048,N_19085,N_17628);
or U27049 (N_27049,N_16190,N_19442);
and U27050 (N_27050,N_10316,N_13594);
nand U27051 (N_27051,N_19439,N_18282);
nor U27052 (N_27052,N_12667,N_14052);
nand U27053 (N_27053,N_15414,N_17289);
nor U27054 (N_27054,N_16605,N_18393);
nand U27055 (N_27055,N_12770,N_14288);
or U27056 (N_27056,N_19863,N_11586);
and U27057 (N_27057,N_18971,N_17213);
and U27058 (N_27058,N_12438,N_17171);
or U27059 (N_27059,N_14842,N_14994);
nor U27060 (N_27060,N_15142,N_12134);
nand U27061 (N_27061,N_16342,N_16552);
nand U27062 (N_27062,N_15237,N_16937);
nor U27063 (N_27063,N_14813,N_14090);
and U27064 (N_27064,N_12671,N_11114);
nand U27065 (N_27065,N_16808,N_10129);
or U27066 (N_27066,N_16029,N_13589);
nand U27067 (N_27067,N_10337,N_10232);
nand U27068 (N_27068,N_14388,N_10549);
or U27069 (N_27069,N_10012,N_12792);
and U27070 (N_27070,N_16898,N_11949);
or U27071 (N_27071,N_19403,N_12264);
or U27072 (N_27072,N_12854,N_12699);
nand U27073 (N_27073,N_17389,N_10390);
nand U27074 (N_27074,N_10419,N_14612);
nor U27075 (N_27075,N_13568,N_15562);
nand U27076 (N_27076,N_15712,N_12928);
nand U27077 (N_27077,N_11419,N_16606);
and U27078 (N_27078,N_17227,N_11353);
nand U27079 (N_27079,N_19797,N_18566);
nor U27080 (N_27080,N_18483,N_12246);
xor U27081 (N_27081,N_19385,N_13878);
nor U27082 (N_27082,N_15361,N_10482);
nand U27083 (N_27083,N_10262,N_17150);
or U27084 (N_27084,N_16412,N_17718);
or U27085 (N_27085,N_16045,N_19566);
nand U27086 (N_27086,N_12268,N_18540);
nand U27087 (N_27087,N_17518,N_12390);
or U27088 (N_27088,N_18344,N_19259);
or U27089 (N_27089,N_18987,N_14287);
and U27090 (N_27090,N_17199,N_14536);
nor U27091 (N_27091,N_10032,N_14619);
and U27092 (N_27092,N_12998,N_16316);
xor U27093 (N_27093,N_12515,N_17690);
nor U27094 (N_27094,N_15246,N_15972);
or U27095 (N_27095,N_13322,N_11669);
xnor U27096 (N_27096,N_14197,N_17098);
or U27097 (N_27097,N_15089,N_14999);
and U27098 (N_27098,N_17910,N_11717);
nor U27099 (N_27099,N_14203,N_18466);
nand U27100 (N_27100,N_13957,N_17911);
nand U27101 (N_27101,N_16936,N_16183);
xnor U27102 (N_27102,N_15166,N_15815);
nand U27103 (N_27103,N_13429,N_16117);
nand U27104 (N_27104,N_11004,N_13270);
nand U27105 (N_27105,N_19682,N_13342);
xor U27106 (N_27106,N_19012,N_16939);
nand U27107 (N_27107,N_14084,N_14827);
nand U27108 (N_27108,N_11773,N_17650);
nand U27109 (N_27109,N_11443,N_15584);
and U27110 (N_27110,N_12790,N_16738);
nand U27111 (N_27111,N_18773,N_14083);
or U27112 (N_27112,N_18977,N_13868);
or U27113 (N_27113,N_11611,N_17515);
and U27114 (N_27114,N_14632,N_17165);
xor U27115 (N_27115,N_16908,N_19239);
nand U27116 (N_27116,N_15460,N_19182);
xor U27117 (N_27117,N_10788,N_14856);
or U27118 (N_27118,N_18006,N_18772);
xnor U27119 (N_27119,N_16523,N_17148);
nor U27120 (N_27120,N_13719,N_11687);
nand U27121 (N_27121,N_11167,N_10078);
or U27122 (N_27122,N_15456,N_19502);
nor U27123 (N_27123,N_13308,N_16877);
xnor U27124 (N_27124,N_16759,N_15165);
nor U27125 (N_27125,N_11617,N_16250);
nand U27126 (N_27126,N_13513,N_10134);
and U27127 (N_27127,N_17701,N_17927);
xnor U27128 (N_27128,N_14257,N_10309);
or U27129 (N_27129,N_15907,N_16601);
nor U27130 (N_27130,N_14025,N_19584);
nand U27131 (N_27131,N_19888,N_17790);
and U27132 (N_27132,N_14065,N_15245);
or U27133 (N_27133,N_12168,N_11228);
nor U27134 (N_27134,N_17856,N_10055);
and U27135 (N_27135,N_14137,N_14465);
nand U27136 (N_27136,N_14119,N_18103);
and U27137 (N_27137,N_18802,N_11175);
nor U27138 (N_27138,N_16226,N_12664);
nand U27139 (N_27139,N_16458,N_16582);
or U27140 (N_27140,N_13968,N_18668);
or U27141 (N_27141,N_14375,N_14415);
and U27142 (N_27142,N_18070,N_17036);
nand U27143 (N_27143,N_16506,N_15411);
or U27144 (N_27144,N_10165,N_13808);
or U27145 (N_27145,N_13951,N_19031);
or U27146 (N_27146,N_13324,N_17763);
or U27147 (N_27147,N_14394,N_12799);
or U27148 (N_27148,N_15905,N_17817);
nor U27149 (N_27149,N_11526,N_16383);
and U27150 (N_27150,N_13407,N_13842);
nor U27151 (N_27151,N_12189,N_11189);
nor U27152 (N_27152,N_19357,N_19081);
and U27153 (N_27153,N_15955,N_14882);
nor U27154 (N_27154,N_10903,N_11033);
or U27155 (N_27155,N_13807,N_13373);
nor U27156 (N_27156,N_15368,N_14076);
and U27157 (N_27157,N_13855,N_14207);
or U27158 (N_27158,N_14523,N_10677);
and U27159 (N_27159,N_13949,N_19039);
nor U27160 (N_27160,N_15896,N_10668);
or U27161 (N_27161,N_14509,N_17911);
xor U27162 (N_27162,N_16575,N_17109);
xnor U27163 (N_27163,N_13859,N_15673);
or U27164 (N_27164,N_11424,N_12317);
or U27165 (N_27165,N_15428,N_19999);
and U27166 (N_27166,N_13574,N_17685);
nand U27167 (N_27167,N_12198,N_17326);
nor U27168 (N_27168,N_13349,N_12145);
nand U27169 (N_27169,N_17069,N_12104);
or U27170 (N_27170,N_14762,N_11246);
nor U27171 (N_27171,N_16733,N_11770);
or U27172 (N_27172,N_18120,N_17470);
and U27173 (N_27173,N_11530,N_11200);
and U27174 (N_27174,N_14521,N_12189);
nor U27175 (N_27175,N_11366,N_14849);
and U27176 (N_27176,N_19585,N_13901);
nor U27177 (N_27177,N_13719,N_18132);
nor U27178 (N_27178,N_14716,N_16194);
or U27179 (N_27179,N_13460,N_11306);
nor U27180 (N_27180,N_11001,N_14420);
or U27181 (N_27181,N_11470,N_12811);
nor U27182 (N_27182,N_12039,N_19913);
or U27183 (N_27183,N_15031,N_15305);
and U27184 (N_27184,N_14861,N_19465);
and U27185 (N_27185,N_15406,N_19793);
nand U27186 (N_27186,N_17758,N_15847);
nand U27187 (N_27187,N_12027,N_19569);
nand U27188 (N_27188,N_19254,N_11599);
xor U27189 (N_27189,N_15697,N_16374);
or U27190 (N_27190,N_11182,N_12604);
and U27191 (N_27191,N_15705,N_13629);
nor U27192 (N_27192,N_18272,N_13522);
nand U27193 (N_27193,N_11343,N_18486);
nor U27194 (N_27194,N_13097,N_10423);
nand U27195 (N_27195,N_12124,N_11584);
or U27196 (N_27196,N_14919,N_14657);
nor U27197 (N_27197,N_17166,N_19876);
and U27198 (N_27198,N_11672,N_13499);
nor U27199 (N_27199,N_16654,N_13974);
nor U27200 (N_27200,N_19207,N_16027);
nand U27201 (N_27201,N_17478,N_15546);
nor U27202 (N_27202,N_17434,N_12570);
or U27203 (N_27203,N_18679,N_15870);
xor U27204 (N_27204,N_19705,N_15476);
xor U27205 (N_27205,N_12644,N_15490);
and U27206 (N_27206,N_19978,N_10652);
xor U27207 (N_27207,N_18279,N_17430);
nand U27208 (N_27208,N_11517,N_19536);
nand U27209 (N_27209,N_16246,N_12306);
or U27210 (N_27210,N_10967,N_13719);
and U27211 (N_27211,N_16707,N_12314);
nor U27212 (N_27212,N_11104,N_16251);
or U27213 (N_27213,N_12329,N_11206);
or U27214 (N_27214,N_15530,N_11375);
nand U27215 (N_27215,N_18476,N_10168);
nor U27216 (N_27216,N_15116,N_17160);
xor U27217 (N_27217,N_17987,N_15692);
nand U27218 (N_27218,N_13573,N_12447);
or U27219 (N_27219,N_16858,N_16975);
nor U27220 (N_27220,N_15867,N_14497);
nand U27221 (N_27221,N_19859,N_13900);
nand U27222 (N_27222,N_10158,N_16210);
nor U27223 (N_27223,N_15080,N_16026);
nor U27224 (N_27224,N_16268,N_12811);
and U27225 (N_27225,N_15363,N_16463);
or U27226 (N_27226,N_10787,N_11175);
nand U27227 (N_27227,N_12652,N_10347);
or U27228 (N_27228,N_15065,N_19527);
and U27229 (N_27229,N_10165,N_17639);
xor U27230 (N_27230,N_11863,N_12918);
xor U27231 (N_27231,N_15689,N_14088);
or U27232 (N_27232,N_18916,N_19451);
nor U27233 (N_27233,N_13731,N_12752);
xnor U27234 (N_27234,N_18612,N_17933);
or U27235 (N_27235,N_10559,N_15050);
and U27236 (N_27236,N_12797,N_19506);
nor U27237 (N_27237,N_13830,N_19000);
nor U27238 (N_27238,N_19347,N_12488);
or U27239 (N_27239,N_16855,N_18701);
or U27240 (N_27240,N_19086,N_14013);
nand U27241 (N_27241,N_15637,N_10138);
nand U27242 (N_27242,N_13947,N_18772);
or U27243 (N_27243,N_10027,N_18319);
or U27244 (N_27244,N_10048,N_15727);
nor U27245 (N_27245,N_10803,N_14210);
and U27246 (N_27246,N_13676,N_19341);
nor U27247 (N_27247,N_16202,N_16536);
nand U27248 (N_27248,N_16097,N_12974);
nor U27249 (N_27249,N_19515,N_11200);
and U27250 (N_27250,N_13771,N_16548);
and U27251 (N_27251,N_13595,N_17012);
and U27252 (N_27252,N_11437,N_18710);
and U27253 (N_27253,N_15477,N_17412);
nor U27254 (N_27254,N_17021,N_15167);
nand U27255 (N_27255,N_11864,N_17982);
or U27256 (N_27256,N_12289,N_12173);
or U27257 (N_27257,N_12516,N_10859);
and U27258 (N_27258,N_18642,N_18559);
and U27259 (N_27259,N_10677,N_10758);
and U27260 (N_27260,N_17755,N_15690);
or U27261 (N_27261,N_17347,N_10736);
xnor U27262 (N_27262,N_16829,N_19877);
nor U27263 (N_27263,N_14669,N_12618);
xnor U27264 (N_27264,N_16898,N_14511);
or U27265 (N_27265,N_14389,N_18081);
nand U27266 (N_27266,N_17200,N_19083);
nor U27267 (N_27267,N_18749,N_10921);
and U27268 (N_27268,N_15847,N_15640);
and U27269 (N_27269,N_17326,N_12834);
or U27270 (N_27270,N_18071,N_11798);
nand U27271 (N_27271,N_12648,N_19020);
nand U27272 (N_27272,N_11002,N_12061);
or U27273 (N_27273,N_14593,N_19234);
xor U27274 (N_27274,N_14633,N_19351);
or U27275 (N_27275,N_10150,N_17953);
and U27276 (N_27276,N_10349,N_13098);
or U27277 (N_27277,N_10865,N_18082);
nor U27278 (N_27278,N_16888,N_12038);
nor U27279 (N_27279,N_19213,N_17518);
nand U27280 (N_27280,N_18964,N_14956);
nand U27281 (N_27281,N_17822,N_14645);
or U27282 (N_27282,N_14063,N_17529);
nor U27283 (N_27283,N_12852,N_12083);
and U27284 (N_27284,N_15586,N_15019);
nand U27285 (N_27285,N_14947,N_16780);
or U27286 (N_27286,N_10397,N_17806);
and U27287 (N_27287,N_13954,N_17849);
and U27288 (N_27288,N_16037,N_16252);
nand U27289 (N_27289,N_12609,N_12906);
and U27290 (N_27290,N_19971,N_19450);
nor U27291 (N_27291,N_15045,N_15740);
or U27292 (N_27292,N_16003,N_12767);
nor U27293 (N_27293,N_11337,N_11251);
or U27294 (N_27294,N_13508,N_19409);
xnor U27295 (N_27295,N_13979,N_16523);
or U27296 (N_27296,N_17585,N_18610);
or U27297 (N_27297,N_15825,N_17723);
nand U27298 (N_27298,N_17046,N_19481);
and U27299 (N_27299,N_12673,N_19685);
nand U27300 (N_27300,N_10401,N_15922);
and U27301 (N_27301,N_16421,N_14690);
nor U27302 (N_27302,N_12263,N_14084);
or U27303 (N_27303,N_12181,N_14122);
nor U27304 (N_27304,N_17228,N_17685);
or U27305 (N_27305,N_14170,N_18922);
nor U27306 (N_27306,N_18265,N_11526);
nand U27307 (N_27307,N_12383,N_15533);
nor U27308 (N_27308,N_15789,N_14612);
and U27309 (N_27309,N_15910,N_19124);
and U27310 (N_27310,N_12497,N_15752);
nand U27311 (N_27311,N_17773,N_15074);
nor U27312 (N_27312,N_18729,N_18643);
and U27313 (N_27313,N_16399,N_18970);
nor U27314 (N_27314,N_13629,N_14354);
or U27315 (N_27315,N_11755,N_16294);
xor U27316 (N_27316,N_18617,N_18381);
and U27317 (N_27317,N_10417,N_15660);
or U27318 (N_27318,N_15569,N_15567);
nand U27319 (N_27319,N_13135,N_17746);
and U27320 (N_27320,N_19007,N_18361);
or U27321 (N_27321,N_13448,N_10677);
nor U27322 (N_27322,N_15985,N_12224);
nand U27323 (N_27323,N_10712,N_17267);
nand U27324 (N_27324,N_19026,N_11024);
and U27325 (N_27325,N_17281,N_10765);
nand U27326 (N_27326,N_18459,N_17611);
or U27327 (N_27327,N_12403,N_19127);
and U27328 (N_27328,N_17971,N_14580);
nor U27329 (N_27329,N_10520,N_15478);
or U27330 (N_27330,N_14438,N_18765);
xor U27331 (N_27331,N_12095,N_17968);
xor U27332 (N_27332,N_18175,N_15667);
xor U27333 (N_27333,N_16159,N_19782);
and U27334 (N_27334,N_12091,N_13279);
nor U27335 (N_27335,N_10813,N_10990);
nand U27336 (N_27336,N_11170,N_16338);
and U27337 (N_27337,N_13825,N_17979);
or U27338 (N_27338,N_13226,N_13157);
nand U27339 (N_27339,N_17631,N_16319);
and U27340 (N_27340,N_16770,N_14300);
nand U27341 (N_27341,N_10772,N_10762);
and U27342 (N_27342,N_12456,N_12877);
nor U27343 (N_27343,N_15897,N_18743);
and U27344 (N_27344,N_14884,N_11809);
or U27345 (N_27345,N_19441,N_14490);
and U27346 (N_27346,N_19074,N_19997);
nand U27347 (N_27347,N_11609,N_17999);
or U27348 (N_27348,N_19347,N_10398);
nor U27349 (N_27349,N_17571,N_10465);
nand U27350 (N_27350,N_17851,N_15517);
and U27351 (N_27351,N_13821,N_16812);
nor U27352 (N_27352,N_13910,N_13561);
and U27353 (N_27353,N_16842,N_14490);
or U27354 (N_27354,N_12832,N_18073);
nor U27355 (N_27355,N_14214,N_19096);
nor U27356 (N_27356,N_15159,N_19354);
nor U27357 (N_27357,N_11303,N_17431);
nand U27358 (N_27358,N_12537,N_11149);
nand U27359 (N_27359,N_11012,N_11187);
or U27360 (N_27360,N_13396,N_19663);
nor U27361 (N_27361,N_18690,N_17215);
or U27362 (N_27362,N_17877,N_12754);
xor U27363 (N_27363,N_15661,N_19099);
and U27364 (N_27364,N_11198,N_10145);
or U27365 (N_27365,N_16550,N_18448);
nand U27366 (N_27366,N_10224,N_13848);
or U27367 (N_27367,N_12436,N_11009);
nand U27368 (N_27368,N_11709,N_18102);
xor U27369 (N_27369,N_18402,N_17199);
and U27370 (N_27370,N_10483,N_15237);
and U27371 (N_27371,N_13121,N_14360);
and U27372 (N_27372,N_18830,N_15842);
nand U27373 (N_27373,N_15922,N_13790);
nor U27374 (N_27374,N_19138,N_12203);
or U27375 (N_27375,N_19497,N_10472);
nand U27376 (N_27376,N_11248,N_14332);
and U27377 (N_27377,N_13588,N_16821);
and U27378 (N_27378,N_10753,N_18430);
nand U27379 (N_27379,N_11823,N_19475);
nor U27380 (N_27380,N_10896,N_17115);
or U27381 (N_27381,N_14274,N_18109);
or U27382 (N_27382,N_17848,N_16019);
and U27383 (N_27383,N_16880,N_16801);
and U27384 (N_27384,N_10222,N_12107);
nand U27385 (N_27385,N_19994,N_17536);
nor U27386 (N_27386,N_13478,N_18467);
or U27387 (N_27387,N_16578,N_10020);
xor U27388 (N_27388,N_15117,N_18839);
nand U27389 (N_27389,N_16080,N_19086);
xor U27390 (N_27390,N_14123,N_16753);
or U27391 (N_27391,N_19240,N_10348);
nor U27392 (N_27392,N_11188,N_10282);
nor U27393 (N_27393,N_19250,N_10474);
nor U27394 (N_27394,N_10755,N_11675);
xnor U27395 (N_27395,N_15338,N_16604);
nand U27396 (N_27396,N_18951,N_19297);
or U27397 (N_27397,N_14842,N_10094);
and U27398 (N_27398,N_12579,N_10615);
or U27399 (N_27399,N_18762,N_12487);
nand U27400 (N_27400,N_11500,N_11367);
or U27401 (N_27401,N_13276,N_11716);
nand U27402 (N_27402,N_15478,N_12676);
or U27403 (N_27403,N_14039,N_18497);
nand U27404 (N_27404,N_17300,N_11314);
nor U27405 (N_27405,N_14150,N_14232);
nor U27406 (N_27406,N_18304,N_10907);
or U27407 (N_27407,N_17536,N_12946);
and U27408 (N_27408,N_17087,N_10704);
xnor U27409 (N_27409,N_14183,N_18048);
and U27410 (N_27410,N_18723,N_14584);
nand U27411 (N_27411,N_14787,N_19907);
and U27412 (N_27412,N_14656,N_10535);
nand U27413 (N_27413,N_15134,N_16847);
and U27414 (N_27414,N_13081,N_16417);
nor U27415 (N_27415,N_17712,N_12188);
nand U27416 (N_27416,N_18147,N_15133);
nor U27417 (N_27417,N_15735,N_11767);
nand U27418 (N_27418,N_11806,N_11775);
nand U27419 (N_27419,N_18279,N_19173);
and U27420 (N_27420,N_11628,N_11895);
nand U27421 (N_27421,N_12471,N_11380);
nand U27422 (N_27422,N_19277,N_13767);
and U27423 (N_27423,N_17059,N_14993);
nor U27424 (N_27424,N_12738,N_15092);
and U27425 (N_27425,N_18622,N_11394);
nand U27426 (N_27426,N_16869,N_16296);
nor U27427 (N_27427,N_14491,N_10105);
or U27428 (N_27428,N_10051,N_10426);
or U27429 (N_27429,N_13264,N_18862);
or U27430 (N_27430,N_12085,N_11524);
or U27431 (N_27431,N_18154,N_14116);
and U27432 (N_27432,N_17760,N_19348);
nand U27433 (N_27433,N_13113,N_11435);
xor U27434 (N_27434,N_12861,N_10219);
nand U27435 (N_27435,N_19891,N_10642);
or U27436 (N_27436,N_16102,N_11353);
nand U27437 (N_27437,N_15928,N_18193);
or U27438 (N_27438,N_16708,N_16263);
or U27439 (N_27439,N_15509,N_14805);
and U27440 (N_27440,N_18314,N_16302);
nor U27441 (N_27441,N_17052,N_16951);
and U27442 (N_27442,N_17467,N_10504);
nand U27443 (N_27443,N_14616,N_19806);
and U27444 (N_27444,N_16485,N_15873);
nand U27445 (N_27445,N_19605,N_15507);
xor U27446 (N_27446,N_15596,N_19497);
and U27447 (N_27447,N_13277,N_16139);
nor U27448 (N_27448,N_14189,N_10133);
and U27449 (N_27449,N_13238,N_12489);
nor U27450 (N_27450,N_16294,N_19155);
and U27451 (N_27451,N_18341,N_15866);
nor U27452 (N_27452,N_11591,N_13733);
or U27453 (N_27453,N_17939,N_14675);
or U27454 (N_27454,N_13225,N_17038);
nand U27455 (N_27455,N_18887,N_10013);
nand U27456 (N_27456,N_10471,N_15674);
and U27457 (N_27457,N_16268,N_18083);
and U27458 (N_27458,N_16644,N_18256);
or U27459 (N_27459,N_16665,N_11075);
or U27460 (N_27460,N_16233,N_15459);
nand U27461 (N_27461,N_18588,N_16588);
nor U27462 (N_27462,N_19042,N_15822);
nor U27463 (N_27463,N_12009,N_15719);
or U27464 (N_27464,N_16700,N_12079);
nand U27465 (N_27465,N_16170,N_12620);
xor U27466 (N_27466,N_19602,N_10452);
nor U27467 (N_27467,N_19588,N_19191);
nand U27468 (N_27468,N_15612,N_11713);
or U27469 (N_27469,N_11963,N_16030);
and U27470 (N_27470,N_18346,N_13203);
nand U27471 (N_27471,N_15161,N_18767);
nor U27472 (N_27472,N_12995,N_14696);
nand U27473 (N_27473,N_19647,N_17144);
or U27474 (N_27474,N_14936,N_19008);
nand U27475 (N_27475,N_14434,N_11308);
nor U27476 (N_27476,N_13625,N_14678);
nand U27477 (N_27477,N_17576,N_17267);
nor U27478 (N_27478,N_19873,N_12691);
and U27479 (N_27479,N_15874,N_15220);
xnor U27480 (N_27480,N_18101,N_13859);
nand U27481 (N_27481,N_16922,N_11213);
and U27482 (N_27482,N_16556,N_10580);
nor U27483 (N_27483,N_14006,N_18502);
and U27484 (N_27484,N_14709,N_10408);
nand U27485 (N_27485,N_10173,N_12181);
and U27486 (N_27486,N_19927,N_18310);
and U27487 (N_27487,N_16376,N_10520);
nand U27488 (N_27488,N_17575,N_10408);
nor U27489 (N_27489,N_14890,N_11222);
and U27490 (N_27490,N_17097,N_11624);
and U27491 (N_27491,N_11960,N_10414);
xor U27492 (N_27492,N_12192,N_17068);
nor U27493 (N_27493,N_16032,N_18975);
nor U27494 (N_27494,N_17476,N_12664);
and U27495 (N_27495,N_18576,N_11334);
or U27496 (N_27496,N_16597,N_16757);
nor U27497 (N_27497,N_13625,N_15566);
and U27498 (N_27498,N_11070,N_15988);
or U27499 (N_27499,N_15590,N_19557);
and U27500 (N_27500,N_14281,N_19978);
xor U27501 (N_27501,N_10852,N_13746);
or U27502 (N_27502,N_11736,N_12088);
or U27503 (N_27503,N_13135,N_12044);
nor U27504 (N_27504,N_10672,N_19725);
nor U27505 (N_27505,N_14141,N_14408);
xor U27506 (N_27506,N_18609,N_18073);
or U27507 (N_27507,N_15630,N_14809);
and U27508 (N_27508,N_18539,N_12725);
and U27509 (N_27509,N_18497,N_10639);
and U27510 (N_27510,N_17959,N_18329);
nand U27511 (N_27511,N_16448,N_13298);
nand U27512 (N_27512,N_19713,N_16426);
xnor U27513 (N_27513,N_15224,N_19113);
nand U27514 (N_27514,N_15644,N_16988);
nand U27515 (N_27515,N_12333,N_15644);
or U27516 (N_27516,N_11589,N_14353);
or U27517 (N_27517,N_18564,N_13099);
nor U27518 (N_27518,N_12392,N_13425);
and U27519 (N_27519,N_17437,N_19640);
and U27520 (N_27520,N_16062,N_15829);
nor U27521 (N_27521,N_14106,N_19172);
nand U27522 (N_27522,N_14705,N_19223);
and U27523 (N_27523,N_10046,N_13239);
nand U27524 (N_27524,N_11731,N_15656);
nand U27525 (N_27525,N_15591,N_12714);
and U27526 (N_27526,N_18997,N_16826);
and U27527 (N_27527,N_12404,N_11492);
xor U27528 (N_27528,N_15707,N_16624);
xnor U27529 (N_27529,N_17458,N_15253);
nand U27530 (N_27530,N_13270,N_17676);
nand U27531 (N_27531,N_18299,N_18538);
and U27532 (N_27532,N_13004,N_17449);
and U27533 (N_27533,N_15363,N_11827);
or U27534 (N_27534,N_14979,N_19936);
nand U27535 (N_27535,N_13008,N_15810);
or U27536 (N_27536,N_15901,N_16174);
and U27537 (N_27537,N_18977,N_13304);
nand U27538 (N_27538,N_17081,N_12608);
and U27539 (N_27539,N_14951,N_14916);
nor U27540 (N_27540,N_13545,N_18205);
xor U27541 (N_27541,N_18914,N_19272);
or U27542 (N_27542,N_17177,N_18730);
xnor U27543 (N_27543,N_11259,N_12290);
xnor U27544 (N_27544,N_18537,N_15858);
or U27545 (N_27545,N_17216,N_14900);
nand U27546 (N_27546,N_15932,N_18951);
and U27547 (N_27547,N_19418,N_16861);
or U27548 (N_27548,N_11629,N_16332);
or U27549 (N_27549,N_12690,N_11148);
nor U27550 (N_27550,N_18197,N_18018);
nor U27551 (N_27551,N_19036,N_15329);
nand U27552 (N_27552,N_19683,N_10977);
or U27553 (N_27553,N_11561,N_17473);
nor U27554 (N_27554,N_18809,N_17065);
and U27555 (N_27555,N_10774,N_12837);
nand U27556 (N_27556,N_18427,N_10983);
nor U27557 (N_27557,N_14649,N_11712);
or U27558 (N_27558,N_13423,N_13986);
nor U27559 (N_27559,N_13437,N_19972);
nand U27560 (N_27560,N_16470,N_11331);
nor U27561 (N_27561,N_12355,N_16815);
nor U27562 (N_27562,N_19254,N_19550);
or U27563 (N_27563,N_11887,N_18033);
and U27564 (N_27564,N_18055,N_18533);
or U27565 (N_27565,N_16552,N_11025);
or U27566 (N_27566,N_13080,N_12016);
and U27567 (N_27567,N_16087,N_18403);
xor U27568 (N_27568,N_19724,N_14265);
nor U27569 (N_27569,N_11483,N_14144);
and U27570 (N_27570,N_13350,N_17742);
and U27571 (N_27571,N_18662,N_18131);
nor U27572 (N_27572,N_11265,N_17646);
nor U27573 (N_27573,N_19864,N_12035);
nand U27574 (N_27574,N_13840,N_11325);
nand U27575 (N_27575,N_12394,N_10631);
and U27576 (N_27576,N_12665,N_13805);
nor U27577 (N_27577,N_14793,N_14374);
nor U27578 (N_27578,N_17869,N_12711);
and U27579 (N_27579,N_19816,N_11123);
nand U27580 (N_27580,N_11406,N_10728);
or U27581 (N_27581,N_18186,N_16030);
and U27582 (N_27582,N_11272,N_18620);
and U27583 (N_27583,N_18797,N_13765);
xor U27584 (N_27584,N_17237,N_16130);
xnor U27585 (N_27585,N_12716,N_16392);
and U27586 (N_27586,N_10793,N_13672);
nor U27587 (N_27587,N_14075,N_19768);
nor U27588 (N_27588,N_12548,N_18691);
and U27589 (N_27589,N_11702,N_13622);
nand U27590 (N_27590,N_19709,N_17859);
nand U27591 (N_27591,N_19957,N_16654);
nand U27592 (N_27592,N_18894,N_17934);
nor U27593 (N_27593,N_16967,N_17042);
nor U27594 (N_27594,N_12610,N_16142);
or U27595 (N_27595,N_11282,N_15932);
or U27596 (N_27596,N_17046,N_12951);
nor U27597 (N_27597,N_19669,N_17831);
nor U27598 (N_27598,N_11620,N_16826);
or U27599 (N_27599,N_11798,N_19471);
nor U27600 (N_27600,N_12969,N_19898);
nor U27601 (N_27601,N_15078,N_14175);
nand U27602 (N_27602,N_11356,N_19328);
or U27603 (N_27603,N_12373,N_13444);
and U27604 (N_27604,N_19935,N_10480);
and U27605 (N_27605,N_18338,N_14335);
and U27606 (N_27606,N_18315,N_13888);
and U27607 (N_27607,N_12058,N_10396);
or U27608 (N_27608,N_14248,N_14715);
nor U27609 (N_27609,N_14619,N_16684);
nand U27610 (N_27610,N_17157,N_18048);
nor U27611 (N_27611,N_14458,N_17974);
nand U27612 (N_27612,N_12665,N_10328);
nand U27613 (N_27613,N_14554,N_18745);
and U27614 (N_27614,N_12017,N_19339);
or U27615 (N_27615,N_12498,N_14746);
or U27616 (N_27616,N_14011,N_14428);
or U27617 (N_27617,N_18607,N_19042);
or U27618 (N_27618,N_18953,N_19385);
nand U27619 (N_27619,N_16337,N_11399);
xor U27620 (N_27620,N_14110,N_13632);
or U27621 (N_27621,N_16889,N_14248);
nor U27622 (N_27622,N_16194,N_14717);
or U27623 (N_27623,N_17408,N_19001);
or U27624 (N_27624,N_19006,N_13415);
nand U27625 (N_27625,N_15655,N_15105);
or U27626 (N_27626,N_12768,N_13051);
or U27627 (N_27627,N_13761,N_10709);
or U27628 (N_27628,N_13248,N_19692);
and U27629 (N_27629,N_12733,N_12365);
and U27630 (N_27630,N_13375,N_17547);
nor U27631 (N_27631,N_18799,N_14559);
nand U27632 (N_27632,N_18793,N_15542);
xnor U27633 (N_27633,N_13159,N_15631);
nor U27634 (N_27634,N_12622,N_15560);
xnor U27635 (N_27635,N_12041,N_17452);
nor U27636 (N_27636,N_13264,N_15494);
nor U27637 (N_27637,N_15196,N_19364);
nand U27638 (N_27638,N_15341,N_18479);
and U27639 (N_27639,N_17493,N_16100);
and U27640 (N_27640,N_15694,N_19531);
or U27641 (N_27641,N_18691,N_16761);
nand U27642 (N_27642,N_11075,N_10846);
or U27643 (N_27643,N_13427,N_18157);
and U27644 (N_27644,N_17498,N_10952);
and U27645 (N_27645,N_17620,N_15404);
and U27646 (N_27646,N_17779,N_17561);
or U27647 (N_27647,N_13349,N_16905);
xor U27648 (N_27648,N_12092,N_15012);
or U27649 (N_27649,N_15431,N_18520);
or U27650 (N_27650,N_12917,N_18102);
nor U27651 (N_27651,N_11353,N_14704);
nor U27652 (N_27652,N_18142,N_12668);
or U27653 (N_27653,N_15763,N_11029);
or U27654 (N_27654,N_13183,N_14653);
nand U27655 (N_27655,N_17351,N_10680);
or U27656 (N_27656,N_16691,N_12685);
nand U27657 (N_27657,N_19858,N_17956);
xnor U27658 (N_27658,N_13844,N_10522);
or U27659 (N_27659,N_19191,N_19702);
nand U27660 (N_27660,N_19513,N_15286);
or U27661 (N_27661,N_19578,N_16905);
nor U27662 (N_27662,N_17133,N_16008);
nor U27663 (N_27663,N_10309,N_10979);
or U27664 (N_27664,N_16561,N_16982);
xnor U27665 (N_27665,N_19472,N_16214);
and U27666 (N_27666,N_13589,N_15039);
and U27667 (N_27667,N_18998,N_18095);
nand U27668 (N_27668,N_12247,N_15650);
or U27669 (N_27669,N_13409,N_16222);
nand U27670 (N_27670,N_15077,N_18160);
and U27671 (N_27671,N_13273,N_12583);
xor U27672 (N_27672,N_14868,N_13948);
nand U27673 (N_27673,N_11333,N_12381);
and U27674 (N_27674,N_11109,N_16202);
nor U27675 (N_27675,N_13221,N_11748);
nand U27676 (N_27676,N_16894,N_16604);
nand U27677 (N_27677,N_18599,N_12821);
and U27678 (N_27678,N_18088,N_15781);
nand U27679 (N_27679,N_10142,N_11158);
xnor U27680 (N_27680,N_15869,N_12774);
nor U27681 (N_27681,N_11995,N_10230);
nor U27682 (N_27682,N_18581,N_11715);
or U27683 (N_27683,N_15460,N_14737);
nor U27684 (N_27684,N_13207,N_19534);
nor U27685 (N_27685,N_11282,N_17078);
nor U27686 (N_27686,N_11725,N_19585);
and U27687 (N_27687,N_10818,N_10836);
and U27688 (N_27688,N_18336,N_16526);
nand U27689 (N_27689,N_18718,N_14524);
nand U27690 (N_27690,N_10041,N_10067);
and U27691 (N_27691,N_17513,N_12658);
or U27692 (N_27692,N_10935,N_15054);
and U27693 (N_27693,N_18949,N_18021);
or U27694 (N_27694,N_17205,N_15446);
and U27695 (N_27695,N_17289,N_11274);
nand U27696 (N_27696,N_10643,N_19891);
and U27697 (N_27697,N_19474,N_15916);
and U27698 (N_27698,N_17151,N_14292);
nand U27699 (N_27699,N_14295,N_19060);
or U27700 (N_27700,N_18568,N_16137);
nand U27701 (N_27701,N_12818,N_10650);
and U27702 (N_27702,N_13134,N_15987);
and U27703 (N_27703,N_18371,N_13595);
and U27704 (N_27704,N_12498,N_10856);
and U27705 (N_27705,N_17414,N_10102);
nand U27706 (N_27706,N_13663,N_10173);
xor U27707 (N_27707,N_17771,N_18830);
or U27708 (N_27708,N_14247,N_16251);
nand U27709 (N_27709,N_18889,N_14109);
or U27710 (N_27710,N_11507,N_19554);
nor U27711 (N_27711,N_18071,N_14021);
and U27712 (N_27712,N_14137,N_12203);
nor U27713 (N_27713,N_12105,N_11626);
nand U27714 (N_27714,N_19301,N_12683);
or U27715 (N_27715,N_19826,N_11160);
and U27716 (N_27716,N_12871,N_18756);
and U27717 (N_27717,N_13442,N_15979);
and U27718 (N_27718,N_12785,N_13963);
nor U27719 (N_27719,N_11707,N_16946);
or U27720 (N_27720,N_15210,N_14169);
or U27721 (N_27721,N_18521,N_14883);
xor U27722 (N_27722,N_16522,N_17513);
nand U27723 (N_27723,N_11813,N_18035);
nor U27724 (N_27724,N_18167,N_19759);
xnor U27725 (N_27725,N_14619,N_18555);
xor U27726 (N_27726,N_10808,N_13393);
and U27727 (N_27727,N_11121,N_18582);
nand U27728 (N_27728,N_19172,N_10493);
nor U27729 (N_27729,N_16164,N_11781);
or U27730 (N_27730,N_11762,N_11775);
nand U27731 (N_27731,N_18518,N_17729);
and U27732 (N_27732,N_19958,N_10908);
or U27733 (N_27733,N_11697,N_18425);
nand U27734 (N_27734,N_12547,N_11732);
nand U27735 (N_27735,N_17041,N_11280);
nor U27736 (N_27736,N_15906,N_15534);
nand U27737 (N_27737,N_11342,N_18263);
nor U27738 (N_27738,N_15968,N_16258);
xor U27739 (N_27739,N_14621,N_14287);
nor U27740 (N_27740,N_12033,N_15196);
nand U27741 (N_27741,N_12247,N_13163);
nor U27742 (N_27742,N_15116,N_18618);
or U27743 (N_27743,N_13865,N_11535);
nand U27744 (N_27744,N_13303,N_13341);
nor U27745 (N_27745,N_19900,N_12563);
and U27746 (N_27746,N_19838,N_11560);
xor U27747 (N_27747,N_14600,N_12643);
nor U27748 (N_27748,N_12247,N_10240);
or U27749 (N_27749,N_19692,N_11426);
nor U27750 (N_27750,N_12135,N_13840);
or U27751 (N_27751,N_15533,N_11963);
or U27752 (N_27752,N_10799,N_12551);
nand U27753 (N_27753,N_11285,N_17556);
nand U27754 (N_27754,N_18063,N_16596);
and U27755 (N_27755,N_18201,N_11864);
nor U27756 (N_27756,N_17912,N_15235);
and U27757 (N_27757,N_14780,N_18451);
or U27758 (N_27758,N_11923,N_17524);
and U27759 (N_27759,N_15961,N_10567);
xnor U27760 (N_27760,N_19074,N_19533);
or U27761 (N_27761,N_11764,N_17843);
or U27762 (N_27762,N_15948,N_11522);
nor U27763 (N_27763,N_12373,N_16425);
or U27764 (N_27764,N_13537,N_16117);
nand U27765 (N_27765,N_19959,N_16119);
or U27766 (N_27766,N_19000,N_10193);
nor U27767 (N_27767,N_16746,N_15591);
or U27768 (N_27768,N_19708,N_12644);
or U27769 (N_27769,N_12785,N_11763);
or U27770 (N_27770,N_11261,N_18250);
nor U27771 (N_27771,N_16558,N_12435);
nand U27772 (N_27772,N_13319,N_15075);
xor U27773 (N_27773,N_11096,N_17523);
or U27774 (N_27774,N_17590,N_17909);
nor U27775 (N_27775,N_16160,N_14949);
and U27776 (N_27776,N_17100,N_17885);
or U27777 (N_27777,N_11600,N_14581);
or U27778 (N_27778,N_18248,N_16443);
and U27779 (N_27779,N_11709,N_18969);
or U27780 (N_27780,N_11937,N_12636);
nand U27781 (N_27781,N_17840,N_13605);
xor U27782 (N_27782,N_16895,N_10895);
and U27783 (N_27783,N_19531,N_19714);
nand U27784 (N_27784,N_15755,N_10464);
xor U27785 (N_27785,N_16418,N_14636);
nor U27786 (N_27786,N_18867,N_17364);
or U27787 (N_27787,N_15808,N_13742);
and U27788 (N_27788,N_12385,N_13588);
xnor U27789 (N_27789,N_10919,N_13880);
or U27790 (N_27790,N_12647,N_12147);
and U27791 (N_27791,N_17554,N_18836);
xor U27792 (N_27792,N_11817,N_14022);
or U27793 (N_27793,N_15280,N_12118);
and U27794 (N_27794,N_15941,N_13316);
and U27795 (N_27795,N_17524,N_19475);
or U27796 (N_27796,N_10935,N_15755);
nor U27797 (N_27797,N_19911,N_10854);
or U27798 (N_27798,N_19579,N_14940);
nand U27799 (N_27799,N_14322,N_18827);
and U27800 (N_27800,N_16839,N_10719);
nor U27801 (N_27801,N_19755,N_19598);
nor U27802 (N_27802,N_14960,N_14750);
and U27803 (N_27803,N_17055,N_13856);
or U27804 (N_27804,N_18588,N_13928);
nand U27805 (N_27805,N_17014,N_16271);
and U27806 (N_27806,N_15073,N_15406);
or U27807 (N_27807,N_19558,N_13812);
nand U27808 (N_27808,N_10898,N_18906);
nor U27809 (N_27809,N_14392,N_11336);
or U27810 (N_27810,N_15850,N_16678);
nor U27811 (N_27811,N_19502,N_19105);
and U27812 (N_27812,N_10259,N_14104);
or U27813 (N_27813,N_18059,N_15097);
nand U27814 (N_27814,N_12009,N_15902);
nand U27815 (N_27815,N_11745,N_13416);
nand U27816 (N_27816,N_10385,N_12911);
and U27817 (N_27817,N_13553,N_15599);
nor U27818 (N_27818,N_19143,N_12521);
nor U27819 (N_27819,N_13906,N_14448);
nor U27820 (N_27820,N_16689,N_14299);
or U27821 (N_27821,N_13011,N_10636);
or U27822 (N_27822,N_13316,N_11500);
and U27823 (N_27823,N_16579,N_17449);
nor U27824 (N_27824,N_12798,N_10155);
nand U27825 (N_27825,N_17435,N_12771);
or U27826 (N_27826,N_12995,N_15920);
nand U27827 (N_27827,N_12295,N_10531);
or U27828 (N_27828,N_15078,N_13811);
nand U27829 (N_27829,N_19734,N_18204);
nand U27830 (N_27830,N_14019,N_17481);
or U27831 (N_27831,N_10252,N_12364);
nand U27832 (N_27832,N_13178,N_10868);
and U27833 (N_27833,N_13568,N_14922);
nand U27834 (N_27834,N_17752,N_13019);
or U27835 (N_27835,N_14568,N_14599);
nor U27836 (N_27836,N_12813,N_17723);
xnor U27837 (N_27837,N_10196,N_15219);
and U27838 (N_27838,N_14631,N_11967);
nor U27839 (N_27839,N_12150,N_14832);
or U27840 (N_27840,N_10807,N_19472);
nand U27841 (N_27841,N_19091,N_18080);
xor U27842 (N_27842,N_11279,N_13099);
nand U27843 (N_27843,N_15293,N_13854);
and U27844 (N_27844,N_14050,N_15800);
xor U27845 (N_27845,N_12397,N_10584);
or U27846 (N_27846,N_14564,N_14580);
nor U27847 (N_27847,N_14204,N_19304);
and U27848 (N_27848,N_10010,N_15287);
nand U27849 (N_27849,N_19778,N_16994);
and U27850 (N_27850,N_18358,N_18649);
and U27851 (N_27851,N_19761,N_19161);
nand U27852 (N_27852,N_17587,N_19989);
nor U27853 (N_27853,N_13612,N_19176);
xor U27854 (N_27854,N_13229,N_12831);
and U27855 (N_27855,N_16858,N_13293);
nand U27856 (N_27856,N_13982,N_11891);
or U27857 (N_27857,N_18488,N_10005);
or U27858 (N_27858,N_12452,N_17257);
nand U27859 (N_27859,N_15762,N_11328);
and U27860 (N_27860,N_19238,N_19330);
or U27861 (N_27861,N_10801,N_15785);
and U27862 (N_27862,N_13132,N_19211);
nor U27863 (N_27863,N_19979,N_13571);
or U27864 (N_27864,N_13577,N_17410);
and U27865 (N_27865,N_16090,N_15919);
and U27866 (N_27866,N_19380,N_11864);
and U27867 (N_27867,N_11957,N_12663);
and U27868 (N_27868,N_11126,N_17914);
and U27869 (N_27869,N_11516,N_15933);
xor U27870 (N_27870,N_10092,N_19549);
nor U27871 (N_27871,N_10514,N_12014);
nor U27872 (N_27872,N_19809,N_13696);
nand U27873 (N_27873,N_16829,N_16137);
xnor U27874 (N_27874,N_10438,N_13073);
and U27875 (N_27875,N_17761,N_18993);
or U27876 (N_27876,N_14233,N_16309);
and U27877 (N_27877,N_17715,N_12266);
nand U27878 (N_27878,N_11172,N_10985);
and U27879 (N_27879,N_18481,N_14597);
or U27880 (N_27880,N_19058,N_12427);
nand U27881 (N_27881,N_12100,N_11518);
and U27882 (N_27882,N_16981,N_12702);
nor U27883 (N_27883,N_17553,N_14461);
nand U27884 (N_27884,N_11380,N_15435);
and U27885 (N_27885,N_17349,N_12736);
or U27886 (N_27886,N_19303,N_10615);
and U27887 (N_27887,N_10952,N_13454);
and U27888 (N_27888,N_15524,N_19820);
or U27889 (N_27889,N_11061,N_12456);
nand U27890 (N_27890,N_16929,N_17325);
nand U27891 (N_27891,N_11354,N_17147);
nor U27892 (N_27892,N_18091,N_17437);
nand U27893 (N_27893,N_19136,N_19974);
and U27894 (N_27894,N_15965,N_11099);
or U27895 (N_27895,N_17506,N_17137);
nor U27896 (N_27896,N_10216,N_18198);
xnor U27897 (N_27897,N_15801,N_12476);
nand U27898 (N_27898,N_14633,N_11130);
nand U27899 (N_27899,N_19121,N_12488);
xnor U27900 (N_27900,N_12417,N_17510);
xnor U27901 (N_27901,N_11306,N_15032);
nand U27902 (N_27902,N_17812,N_16197);
nand U27903 (N_27903,N_14833,N_15110);
nor U27904 (N_27904,N_14175,N_18687);
or U27905 (N_27905,N_16570,N_17612);
or U27906 (N_27906,N_10277,N_12478);
nand U27907 (N_27907,N_10135,N_18818);
or U27908 (N_27908,N_18553,N_14097);
and U27909 (N_27909,N_18251,N_15995);
nand U27910 (N_27910,N_15491,N_12035);
xnor U27911 (N_27911,N_19175,N_13841);
and U27912 (N_27912,N_15353,N_12596);
nor U27913 (N_27913,N_19100,N_17324);
or U27914 (N_27914,N_14948,N_18604);
or U27915 (N_27915,N_19265,N_15987);
or U27916 (N_27916,N_15345,N_18250);
nand U27917 (N_27917,N_15103,N_11500);
nor U27918 (N_27918,N_12451,N_19542);
and U27919 (N_27919,N_17715,N_12263);
and U27920 (N_27920,N_10350,N_15975);
nand U27921 (N_27921,N_11939,N_13155);
or U27922 (N_27922,N_12937,N_12204);
nand U27923 (N_27923,N_10200,N_18312);
or U27924 (N_27924,N_14512,N_19942);
nand U27925 (N_27925,N_17815,N_15037);
nand U27926 (N_27926,N_10110,N_12515);
and U27927 (N_27927,N_12593,N_14887);
nor U27928 (N_27928,N_10951,N_18831);
nand U27929 (N_27929,N_12963,N_14772);
or U27930 (N_27930,N_18118,N_13039);
nand U27931 (N_27931,N_14845,N_12693);
or U27932 (N_27932,N_18400,N_18097);
and U27933 (N_27933,N_15998,N_13890);
nor U27934 (N_27934,N_19143,N_11287);
xor U27935 (N_27935,N_19500,N_14996);
or U27936 (N_27936,N_12094,N_12890);
and U27937 (N_27937,N_16436,N_19797);
nand U27938 (N_27938,N_12068,N_15160);
and U27939 (N_27939,N_16706,N_14044);
or U27940 (N_27940,N_13041,N_14641);
nand U27941 (N_27941,N_17477,N_18065);
or U27942 (N_27942,N_10038,N_11050);
or U27943 (N_27943,N_11975,N_17026);
or U27944 (N_27944,N_14820,N_10578);
or U27945 (N_27945,N_14259,N_14592);
nor U27946 (N_27946,N_11030,N_11464);
xnor U27947 (N_27947,N_18232,N_10204);
and U27948 (N_27948,N_19482,N_16192);
nand U27949 (N_27949,N_14782,N_13909);
nor U27950 (N_27950,N_10224,N_14626);
nor U27951 (N_27951,N_12868,N_16922);
nand U27952 (N_27952,N_17949,N_19153);
or U27953 (N_27953,N_16203,N_15040);
and U27954 (N_27954,N_14559,N_10424);
and U27955 (N_27955,N_15129,N_15972);
and U27956 (N_27956,N_12657,N_16035);
and U27957 (N_27957,N_15654,N_15312);
and U27958 (N_27958,N_19106,N_10368);
or U27959 (N_27959,N_15632,N_17376);
or U27960 (N_27960,N_11024,N_16206);
or U27961 (N_27961,N_10441,N_13320);
nand U27962 (N_27962,N_18923,N_13736);
nor U27963 (N_27963,N_14922,N_10307);
or U27964 (N_27964,N_14627,N_11526);
and U27965 (N_27965,N_13783,N_17354);
xor U27966 (N_27966,N_14181,N_18275);
and U27967 (N_27967,N_19117,N_14240);
and U27968 (N_27968,N_15909,N_16370);
and U27969 (N_27969,N_13276,N_15481);
nand U27970 (N_27970,N_14916,N_15559);
nand U27971 (N_27971,N_17655,N_10660);
and U27972 (N_27972,N_17896,N_14708);
nand U27973 (N_27973,N_17980,N_11826);
or U27974 (N_27974,N_12130,N_19188);
nor U27975 (N_27975,N_15784,N_11159);
or U27976 (N_27976,N_11636,N_17680);
and U27977 (N_27977,N_10749,N_11662);
nand U27978 (N_27978,N_11534,N_11741);
nand U27979 (N_27979,N_10990,N_11148);
nor U27980 (N_27980,N_15846,N_11482);
xnor U27981 (N_27981,N_14642,N_14311);
and U27982 (N_27982,N_10200,N_16457);
nor U27983 (N_27983,N_19663,N_11639);
nor U27984 (N_27984,N_12138,N_18641);
and U27985 (N_27985,N_15630,N_19606);
and U27986 (N_27986,N_14413,N_13553);
nor U27987 (N_27987,N_15286,N_17646);
nand U27988 (N_27988,N_11926,N_14046);
nand U27989 (N_27989,N_16385,N_14229);
nor U27990 (N_27990,N_15889,N_10835);
xnor U27991 (N_27991,N_19733,N_16167);
nor U27992 (N_27992,N_19277,N_14910);
nand U27993 (N_27993,N_15378,N_10010);
nand U27994 (N_27994,N_11189,N_13742);
or U27995 (N_27995,N_12769,N_19564);
nor U27996 (N_27996,N_15939,N_16873);
nor U27997 (N_27997,N_10749,N_14473);
and U27998 (N_27998,N_13071,N_17001);
or U27999 (N_27999,N_13766,N_15470);
and U28000 (N_28000,N_19527,N_19145);
or U28001 (N_28001,N_11523,N_18757);
nor U28002 (N_28002,N_12132,N_12916);
nand U28003 (N_28003,N_14595,N_18513);
nor U28004 (N_28004,N_16308,N_13256);
or U28005 (N_28005,N_15420,N_15923);
nand U28006 (N_28006,N_17448,N_17770);
and U28007 (N_28007,N_16119,N_16844);
nand U28008 (N_28008,N_13455,N_17122);
and U28009 (N_28009,N_12181,N_19046);
or U28010 (N_28010,N_19637,N_15126);
nor U28011 (N_28011,N_10738,N_18707);
or U28012 (N_28012,N_11039,N_11115);
and U28013 (N_28013,N_16785,N_10764);
and U28014 (N_28014,N_18424,N_13993);
and U28015 (N_28015,N_17563,N_19052);
and U28016 (N_28016,N_16444,N_19681);
or U28017 (N_28017,N_10466,N_10901);
and U28018 (N_28018,N_18158,N_11853);
nand U28019 (N_28019,N_19067,N_11076);
or U28020 (N_28020,N_11817,N_14861);
nor U28021 (N_28021,N_19099,N_19351);
nand U28022 (N_28022,N_11940,N_14389);
nand U28023 (N_28023,N_18420,N_13633);
xnor U28024 (N_28024,N_13118,N_13026);
and U28025 (N_28025,N_19363,N_15747);
and U28026 (N_28026,N_18512,N_18062);
and U28027 (N_28027,N_18706,N_19658);
and U28028 (N_28028,N_12220,N_15332);
and U28029 (N_28029,N_11657,N_10723);
and U28030 (N_28030,N_11605,N_14456);
nand U28031 (N_28031,N_18481,N_11845);
nor U28032 (N_28032,N_18866,N_13800);
nor U28033 (N_28033,N_15157,N_19965);
nand U28034 (N_28034,N_12050,N_17296);
nor U28035 (N_28035,N_19373,N_19143);
or U28036 (N_28036,N_11129,N_12914);
xnor U28037 (N_28037,N_10340,N_17967);
nand U28038 (N_28038,N_12441,N_12836);
nand U28039 (N_28039,N_19440,N_11649);
nand U28040 (N_28040,N_19523,N_12190);
nor U28041 (N_28041,N_17813,N_13487);
nand U28042 (N_28042,N_14217,N_16004);
or U28043 (N_28043,N_10730,N_17242);
or U28044 (N_28044,N_17597,N_18699);
and U28045 (N_28045,N_14772,N_12115);
nand U28046 (N_28046,N_14114,N_16908);
xnor U28047 (N_28047,N_19566,N_14973);
and U28048 (N_28048,N_13478,N_10404);
and U28049 (N_28049,N_11762,N_18428);
nor U28050 (N_28050,N_10917,N_12208);
and U28051 (N_28051,N_11435,N_18907);
xnor U28052 (N_28052,N_12508,N_18636);
nand U28053 (N_28053,N_16440,N_17372);
nor U28054 (N_28054,N_18507,N_12889);
and U28055 (N_28055,N_11040,N_15263);
or U28056 (N_28056,N_11841,N_16315);
xor U28057 (N_28057,N_18191,N_19620);
and U28058 (N_28058,N_11795,N_18922);
nor U28059 (N_28059,N_19928,N_12130);
xnor U28060 (N_28060,N_18289,N_19318);
or U28061 (N_28061,N_18281,N_13123);
and U28062 (N_28062,N_15388,N_16381);
nand U28063 (N_28063,N_19601,N_11279);
and U28064 (N_28064,N_10272,N_10692);
nand U28065 (N_28065,N_11803,N_10039);
and U28066 (N_28066,N_11878,N_12380);
nand U28067 (N_28067,N_16242,N_13153);
nor U28068 (N_28068,N_19164,N_13062);
nand U28069 (N_28069,N_10775,N_17334);
and U28070 (N_28070,N_16300,N_14920);
nand U28071 (N_28071,N_15253,N_19417);
nand U28072 (N_28072,N_18110,N_13548);
or U28073 (N_28073,N_11091,N_12604);
and U28074 (N_28074,N_10084,N_16033);
nand U28075 (N_28075,N_13284,N_19323);
nor U28076 (N_28076,N_13540,N_14120);
nor U28077 (N_28077,N_12010,N_16674);
or U28078 (N_28078,N_10591,N_18100);
nand U28079 (N_28079,N_17354,N_18021);
or U28080 (N_28080,N_18435,N_18953);
or U28081 (N_28081,N_18835,N_18541);
nor U28082 (N_28082,N_12699,N_12565);
and U28083 (N_28083,N_14732,N_10791);
or U28084 (N_28084,N_14600,N_14753);
or U28085 (N_28085,N_13423,N_12950);
and U28086 (N_28086,N_19976,N_14799);
and U28087 (N_28087,N_19276,N_10139);
nor U28088 (N_28088,N_14373,N_13800);
or U28089 (N_28089,N_19988,N_10676);
and U28090 (N_28090,N_12358,N_19301);
and U28091 (N_28091,N_12577,N_19151);
nand U28092 (N_28092,N_11590,N_13277);
nand U28093 (N_28093,N_17768,N_11866);
nand U28094 (N_28094,N_12088,N_12651);
xor U28095 (N_28095,N_17660,N_14629);
nor U28096 (N_28096,N_11937,N_18304);
and U28097 (N_28097,N_19051,N_16745);
and U28098 (N_28098,N_14544,N_11570);
nand U28099 (N_28099,N_17885,N_16629);
nand U28100 (N_28100,N_10374,N_10323);
and U28101 (N_28101,N_10841,N_18521);
nor U28102 (N_28102,N_19556,N_19801);
and U28103 (N_28103,N_19910,N_19839);
nand U28104 (N_28104,N_11975,N_14032);
xnor U28105 (N_28105,N_16446,N_12803);
or U28106 (N_28106,N_17215,N_10323);
or U28107 (N_28107,N_17631,N_12312);
and U28108 (N_28108,N_13194,N_13383);
xnor U28109 (N_28109,N_17166,N_12101);
nor U28110 (N_28110,N_11927,N_10658);
or U28111 (N_28111,N_13372,N_18142);
and U28112 (N_28112,N_17537,N_13289);
nand U28113 (N_28113,N_14793,N_12452);
or U28114 (N_28114,N_16790,N_18515);
or U28115 (N_28115,N_11199,N_16938);
nand U28116 (N_28116,N_10951,N_17566);
nor U28117 (N_28117,N_15363,N_15368);
and U28118 (N_28118,N_11527,N_15146);
nor U28119 (N_28119,N_11942,N_10163);
nand U28120 (N_28120,N_19471,N_16599);
nand U28121 (N_28121,N_14118,N_10554);
nor U28122 (N_28122,N_13770,N_11771);
or U28123 (N_28123,N_10408,N_14077);
nor U28124 (N_28124,N_18059,N_15288);
nor U28125 (N_28125,N_10628,N_16247);
xor U28126 (N_28126,N_12256,N_15596);
nand U28127 (N_28127,N_12097,N_19048);
nor U28128 (N_28128,N_17224,N_13884);
or U28129 (N_28129,N_17962,N_13391);
or U28130 (N_28130,N_14332,N_15049);
nor U28131 (N_28131,N_13893,N_16082);
or U28132 (N_28132,N_18260,N_12288);
or U28133 (N_28133,N_19829,N_15256);
nand U28134 (N_28134,N_18438,N_16100);
and U28135 (N_28135,N_15162,N_15934);
or U28136 (N_28136,N_12098,N_19523);
nand U28137 (N_28137,N_12743,N_14100);
or U28138 (N_28138,N_13408,N_10616);
and U28139 (N_28139,N_16243,N_16569);
nand U28140 (N_28140,N_11447,N_17052);
nor U28141 (N_28141,N_16415,N_17912);
nand U28142 (N_28142,N_13135,N_14860);
and U28143 (N_28143,N_17910,N_18748);
xnor U28144 (N_28144,N_19398,N_14703);
or U28145 (N_28145,N_17507,N_19407);
and U28146 (N_28146,N_16929,N_19785);
nor U28147 (N_28147,N_15994,N_14734);
and U28148 (N_28148,N_12084,N_11199);
nand U28149 (N_28149,N_14071,N_10574);
nor U28150 (N_28150,N_17203,N_14765);
nor U28151 (N_28151,N_11956,N_13420);
nand U28152 (N_28152,N_10633,N_15453);
or U28153 (N_28153,N_18446,N_14736);
nor U28154 (N_28154,N_15708,N_15047);
and U28155 (N_28155,N_13756,N_16774);
and U28156 (N_28156,N_18031,N_12136);
nor U28157 (N_28157,N_12267,N_17919);
or U28158 (N_28158,N_11389,N_17986);
or U28159 (N_28159,N_18023,N_12377);
nand U28160 (N_28160,N_12118,N_11168);
and U28161 (N_28161,N_10174,N_12852);
xor U28162 (N_28162,N_11930,N_12444);
nor U28163 (N_28163,N_11065,N_11538);
nor U28164 (N_28164,N_18617,N_11213);
or U28165 (N_28165,N_13088,N_10898);
and U28166 (N_28166,N_10679,N_17983);
or U28167 (N_28167,N_13995,N_15641);
xnor U28168 (N_28168,N_10072,N_10764);
or U28169 (N_28169,N_16282,N_19385);
or U28170 (N_28170,N_15967,N_17394);
and U28171 (N_28171,N_10891,N_10853);
and U28172 (N_28172,N_13796,N_10862);
nand U28173 (N_28173,N_14734,N_17132);
xnor U28174 (N_28174,N_16987,N_11556);
nand U28175 (N_28175,N_18728,N_17278);
xor U28176 (N_28176,N_17543,N_18234);
or U28177 (N_28177,N_15612,N_19202);
nor U28178 (N_28178,N_13999,N_18805);
or U28179 (N_28179,N_11411,N_19894);
nor U28180 (N_28180,N_14239,N_17682);
and U28181 (N_28181,N_10081,N_13454);
and U28182 (N_28182,N_10619,N_16278);
and U28183 (N_28183,N_18980,N_17175);
nand U28184 (N_28184,N_19896,N_12840);
nor U28185 (N_28185,N_13196,N_16819);
and U28186 (N_28186,N_18379,N_15932);
and U28187 (N_28187,N_19482,N_17311);
nand U28188 (N_28188,N_15912,N_12193);
nor U28189 (N_28189,N_15724,N_15105);
nor U28190 (N_28190,N_12273,N_13210);
nor U28191 (N_28191,N_18812,N_15946);
or U28192 (N_28192,N_14821,N_17253);
nand U28193 (N_28193,N_19534,N_12293);
xor U28194 (N_28194,N_10533,N_11049);
and U28195 (N_28195,N_13695,N_19048);
nand U28196 (N_28196,N_17099,N_19240);
nand U28197 (N_28197,N_14586,N_13161);
nand U28198 (N_28198,N_12645,N_18582);
nor U28199 (N_28199,N_19903,N_15697);
and U28200 (N_28200,N_12110,N_14949);
or U28201 (N_28201,N_11674,N_19162);
or U28202 (N_28202,N_17527,N_12950);
or U28203 (N_28203,N_10389,N_13999);
nand U28204 (N_28204,N_17433,N_17770);
nor U28205 (N_28205,N_17526,N_16275);
nand U28206 (N_28206,N_17196,N_19520);
nor U28207 (N_28207,N_18805,N_11162);
and U28208 (N_28208,N_19208,N_16962);
nor U28209 (N_28209,N_17213,N_19537);
nor U28210 (N_28210,N_11523,N_19213);
nand U28211 (N_28211,N_10923,N_19004);
nor U28212 (N_28212,N_13247,N_19467);
xor U28213 (N_28213,N_16964,N_10899);
or U28214 (N_28214,N_16945,N_10629);
nor U28215 (N_28215,N_11188,N_15948);
or U28216 (N_28216,N_17456,N_15280);
or U28217 (N_28217,N_13269,N_10717);
nand U28218 (N_28218,N_12580,N_19028);
nand U28219 (N_28219,N_18018,N_16013);
nand U28220 (N_28220,N_16127,N_11898);
or U28221 (N_28221,N_17840,N_19866);
xor U28222 (N_28222,N_17884,N_16244);
nor U28223 (N_28223,N_10421,N_12189);
or U28224 (N_28224,N_18483,N_15869);
and U28225 (N_28225,N_16663,N_16516);
or U28226 (N_28226,N_15488,N_17887);
xnor U28227 (N_28227,N_18678,N_18666);
nand U28228 (N_28228,N_19113,N_11269);
nand U28229 (N_28229,N_15359,N_12674);
nor U28230 (N_28230,N_12165,N_18232);
or U28231 (N_28231,N_15368,N_11079);
nand U28232 (N_28232,N_11969,N_17870);
xor U28233 (N_28233,N_12462,N_16622);
nand U28234 (N_28234,N_17921,N_10939);
or U28235 (N_28235,N_12435,N_10573);
and U28236 (N_28236,N_19283,N_11552);
xnor U28237 (N_28237,N_13411,N_18814);
nand U28238 (N_28238,N_10340,N_18698);
nand U28239 (N_28239,N_10423,N_17370);
or U28240 (N_28240,N_14333,N_16739);
nand U28241 (N_28241,N_12822,N_14967);
nand U28242 (N_28242,N_13178,N_19142);
or U28243 (N_28243,N_10724,N_13251);
and U28244 (N_28244,N_11034,N_16248);
nand U28245 (N_28245,N_15775,N_13906);
xnor U28246 (N_28246,N_13501,N_11714);
xnor U28247 (N_28247,N_12856,N_17165);
nor U28248 (N_28248,N_13024,N_11331);
nor U28249 (N_28249,N_11821,N_19679);
and U28250 (N_28250,N_18470,N_15103);
nor U28251 (N_28251,N_10267,N_18686);
or U28252 (N_28252,N_12420,N_13993);
nand U28253 (N_28253,N_18958,N_16731);
xor U28254 (N_28254,N_19139,N_15768);
and U28255 (N_28255,N_11854,N_16759);
nand U28256 (N_28256,N_19776,N_18883);
nor U28257 (N_28257,N_11942,N_19228);
and U28258 (N_28258,N_18089,N_18698);
or U28259 (N_28259,N_16784,N_16848);
and U28260 (N_28260,N_11227,N_11287);
nand U28261 (N_28261,N_11026,N_10184);
nor U28262 (N_28262,N_13270,N_14004);
nor U28263 (N_28263,N_10839,N_14387);
nor U28264 (N_28264,N_16988,N_17528);
nor U28265 (N_28265,N_11462,N_12445);
and U28266 (N_28266,N_14798,N_13232);
nand U28267 (N_28267,N_12772,N_15560);
or U28268 (N_28268,N_10372,N_10645);
nor U28269 (N_28269,N_19214,N_14742);
nor U28270 (N_28270,N_11843,N_10484);
or U28271 (N_28271,N_12621,N_12243);
nand U28272 (N_28272,N_17977,N_11008);
nand U28273 (N_28273,N_16170,N_11829);
xor U28274 (N_28274,N_13073,N_17436);
and U28275 (N_28275,N_14194,N_17379);
and U28276 (N_28276,N_16070,N_19862);
and U28277 (N_28277,N_15556,N_17847);
or U28278 (N_28278,N_18520,N_16024);
nand U28279 (N_28279,N_10889,N_12677);
nand U28280 (N_28280,N_10359,N_15373);
or U28281 (N_28281,N_17918,N_17711);
and U28282 (N_28282,N_11222,N_15557);
nor U28283 (N_28283,N_19635,N_11836);
or U28284 (N_28284,N_12934,N_10668);
nor U28285 (N_28285,N_10064,N_18519);
and U28286 (N_28286,N_13150,N_18419);
nand U28287 (N_28287,N_10174,N_10547);
and U28288 (N_28288,N_12616,N_15851);
xor U28289 (N_28289,N_12320,N_14781);
nand U28290 (N_28290,N_18923,N_16415);
and U28291 (N_28291,N_19770,N_10660);
and U28292 (N_28292,N_17180,N_14838);
nand U28293 (N_28293,N_12192,N_10183);
and U28294 (N_28294,N_13727,N_19648);
nor U28295 (N_28295,N_12185,N_17167);
nor U28296 (N_28296,N_15247,N_18050);
nand U28297 (N_28297,N_12544,N_10339);
nor U28298 (N_28298,N_12421,N_18806);
nor U28299 (N_28299,N_18598,N_12122);
or U28300 (N_28300,N_10459,N_16171);
or U28301 (N_28301,N_11412,N_12175);
and U28302 (N_28302,N_19494,N_17649);
or U28303 (N_28303,N_12468,N_17507);
and U28304 (N_28304,N_18398,N_18371);
nand U28305 (N_28305,N_13965,N_15528);
or U28306 (N_28306,N_14985,N_10774);
nand U28307 (N_28307,N_11812,N_19392);
or U28308 (N_28308,N_11793,N_16940);
nor U28309 (N_28309,N_14111,N_12356);
nor U28310 (N_28310,N_12009,N_19898);
nor U28311 (N_28311,N_18871,N_17510);
and U28312 (N_28312,N_15746,N_18907);
or U28313 (N_28313,N_10320,N_13928);
xor U28314 (N_28314,N_19824,N_11852);
and U28315 (N_28315,N_14205,N_16457);
nand U28316 (N_28316,N_14743,N_13582);
nand U28317 (N_28317,N_14683,N_19764);
nor U28318 (N_28318,N_13248,N_19358);
or U28319 (N_28319,N_17762,N_13538);
nand U28320 (N_28320,N_18852,N_11991);
xnor U28321 (N_28321,N_11408,N_19592);
nand U28322 (N_28322,N_13338,N_17737);
and U28323 (N_28323,N_14753,N_13462);
or U28324 (N_28324,N_19764,N_18909);
and U28325 (N_28325,N_13996,N_18209);
or U28326 (N_28326,N_11248,N_15221);
xor U28327 (N_28327,N_12437,N_10954);
xnor U28328 (N_28328,N_14104,N_15271);
nand U28329 (N_28329,N_13153,N_10867);
nor U28330 (N_28330,N_13743,N_17206);
and U28331 (N_28331,N_15018,N_13515);
nand U28332 (N_28332,N_12988,N_17279);
nor U28333 (N_28333,N_10493,N_13667);
or U28334 (N_28334,N_14310,N_19216);
nand U28335 (N_28335,N_14211,N_18125);
and U28336 (N_28336,N_14910,N_10321);
nor U28337 (N_28337,N_17291,N_15873);
xor U28338 (N_28338,N_10763,N_14338);
and U28339 (N_28339,N_19387,N_13273);
nand U28340 (N_28340,N_15042,N_18965);
nor U28341 (N_28341,N_16392,N_15919);
and U28342 (N_28342,N_17412,N_13774);
nor U28343 (N_28343,N_19870,N_12626);
and U28344 (N_28344,N_14759,N_14985);
or U28345 (N_28345,N_16239,N_12132);
xor U28346 (N_28346,N_10727,N_16209);
and U28347 (N_28347,N_10881,N_10169);
or U28348 (N_28348,N_15848,N_15112);
nor U28349 (N_28349,N_18091,N_16809);
and U28350 (N_28350,N_11930,N_11310);
nor U28351 (N_28351,N_16836,N_13786);
xor U28352 (N_28352,N_16876,N_16062);
and U28353 (N_28353,N_13443,N_18377);
xnor U28354 (N_28354,N_15346,N_16084);
and U28355 (N_28355,N_19028,N_19894);
or U28356 (N_28356,N_13086,N_14486);
xor U28357 (N_28357,N_19758,N_12092);
nand U28358 (N_28358,N_16148,N_14987);
nor U28359 (N_28359,N_12109,N_12955);
or U28360 (N_28360,N_13555,N_18303);
xnor U28361 (N_28361,N_17415,N_13241);
or U28362 (N_28362,N_19577,N_15783);
nand U28363 (N_28363,N_17792,N_16150);
and U28364 (N_28364,N_16383,N_14852);
nand U28365 (N_28365,N_14442,N_17880);
nor U28366 (N_28366,N_14545,N_10145);
xor U28367 (N_28367,N_19556,N_13623);
xor U28368 (N_28368,N_10363,N_10099);
nand U28369 (N_28369,N_18922,N_15825);
or U28370 (N_28370,N_19776,N_18514);
nor U28371 (N_28371,N_19755,N_12444);
and U28372 (N_28372,N_19605,N_18764);
nand U28373 (N_28373,N_17837,N_11183);
and U28374 (N_28374,N_11977,N_19261);
or U28375 (N_28375,N_16854,N_12566);
nand U28376 (N_28376,N_13030,N_14552);
nand U28377 (N_28377,N_15342,N_16389);
or U28378 (N_28378,N_16180,N_10435);
and U28379 (N_28379,N_16313,N_12250);
nand U28380 (N_28380,N_17942,N_11459);
nor U28381 (N_28381,N_12188,N_17154);
or U28382 (N_28382,N_17300,N_11657);
or U28383 (N_28383,N_14562,N_16621);
or U28384 (N_28384,N_15916,N_16100);
nand U28385 (N_28385,N_19544,N_13393);
nand U28386 (N_28386,N_10253,N_10055);
nand U28387 (N_28387,N_14977,N_14282);
xnor U28388 (N_28388,N_10936,N_11979);
nor U28389 (N_28389,N_15000,N_13078);
nor U28390 (N_28390,N_17410,N_12128);
or U28391 (N_28391,N_19641,N_13803);
and U28392 (N_28392,N_17916,N_13545);
xnor U28393 (N_28393,N_14015,N_19763);
nand U28394 (N_28394,N_11009,N_15188);
nand U28395 (N_28395,N_17356,N_12973);
or U28396 (N_28396,N_18142,N_15517);
nor U28397 (N_28397,N_15208,N_14176);
nor U28398 (N_28398,N_14309,N_18812);
nor U28399 (N_28399,N_14945,N_16607);
nand U28400 (N_28400,N_14913,N_14163);
nand U28401 (N_28401,N_10696,N_14955);
nand U28402 (N_28402,N_11714,N_10100);
nor U28403 (N_28403,N_13169,N_19882);
nand U28404 (N_28404,N_15901,N_12690);
xor U28405 (N_28405,N_19219,N_13287);
and U28406 (N_28406,N_18411,N_18859);
or U28407 (N_28407,N_19493,N_11112);
nand U28408 (N_28408,N_17066,N_16654);
xor U28409 (N_28409,N_19468,N_17983);
or U28410 (N_28410,N_19221,N_13307);
and U28411 (N_28411,N_17392,N_15747);
or U28412 (N_28412,N_10964,N_13728);
or U28413 (N_28413,N_16237,N_11969);
xor U28414 (N_28414,N_10077,N_18561);
xnor U28415 (N_28415,N_19808,N_18734);
or U28416 (N_28416,N_10998,N_13427);
or U28417 (N_28417,N_15277,N_10677);
and U28418 (N_28418,N_12001,N_14434);
and U28419 (N_28419,N_18631,N_14149);
nand U28420 (N_28420,N_15897,N_19809);
and U28421 (N_28421,N_14120,N_15002);
nor U28422 (N_28422,N_18582,N_13008);
or U28423 (N_28423,N_15635,N_14229);
and U28424 (N_28424,N_11789,N_15124);
and U28425 (N_28425,N_17128,N_10122);
nor U28426 (N_28426,N_15279,N_11781);
xor U28427 (N_28427,N_14216,N_17929);
and U28428 (N_28428,N_14892,N_17359);
nand U28429 (N_28429,N_10608,N_10344);
nand U28430 (N_28430,N_18719,N_15847);
and U28431 (N_28431,N_16747,N_15062);
and U28432 (N_28432,N_15986,N_14386);
nor U28433 (N_28433,N_13499,N_16031);
nand U28434 (N_28434,N_14374,N_17929);
and U28435 (N_28435,N_11452,N_15509);
nor U28436 (N_28436,N_19938,N_18486);
nand U28437 (N_28437,N_14336,N_13929);
nor U28438 (N_28438,N_12358,N_15523);
nand U28439 (N_28439,N_19689,N_14717);
or U28440 (N_28440,N_18552,N_19711);
or U28441 (N_28441,N_15060,N_12005);
and U28442 (N_28442,N_12920,N_15351);
nand U28443 (N_28443,N_13736,N_19396);
nor U28444 (N_28444,N_12388,N_15941);
nand U28445 (N_28445,N_11159,N_11582);
nor U28446 (N_28446,N_14084,N_11123);
xor U28447 (N_28447,N_13702,N_14815);
and U28448 (N_28448,N_13293,N_11678);
xnor U28449 (N_28449,N_13535,N_15781);
or U28450 (N_28450,N_15954,N_15057);
and U28451 (N_28451,N_12775,N_12202);
nand U28452 (N_28452,N_18467,N_18810);
and U28453 (N_28453,N_16936,N_12839);
or U28454 (N_28454,N_12370,N_13365);
and U28455 (N_28455,N_16393,N_19716);
or U28456 (N_28456,N_15912,N_16093);
nor U28457 (N_28457,N_12529,N_11182);
xor U28458 (N_28458,N_14534,N_11401);
or U28459 (N_28459,N_17468,N_14079);
and U28460 (N_28460,N_16005,N_10281);
nor U28461 (N_28461,N_17936,N_11265);
or U28462 (N_28462,N_18668,N_17367);
or U28463 (N_28463,N_11708,N_17234);
nand U28464 (N_28464,N_19159,N_10169);
xor U28465 (N_28465,N_16716,N_19813);
nor U28466 (N_28466,N_18435,N_16539);
and U28467 (N_28467,N_12745,N_10839);
nor U28468 (N_28468,N_10123,N_12659);
and U28469 (N_28469,N_19426,N_19533);
or U28470 (N_28470,N_11602,N_13258);
nand U28471 (N_28471,N_11274,N_18578);
and U28472 (N_28472,N_19076,N_11744);
and U28473 (N_28473,N_10306,N_17789);
and U28474 (N_28474,N_11915,N_14094);
xnor U28475 (N_28475,N_12754,N_10250);
nand U28476 (N_28476,N_19320,N_11433);
or U28477 (N_28477,N_10266,N_15762);
nor U28478 (N_28478,N_14410,N_15966);
or U28479 (N_28479,N_11130,N_13920);
or U28480 (N_28480,N_11070,N_18787);
xnor U28481 (N_28481,N_13247,N_15873);
nand U28482 (N_28482,N_10524,N_12765);
and U28483 (N_28483,N_10507,N_16349);
and U28484 (N_28484,N_13189,N_19298);
nor U28485 (N_28485,N_15524,N_15542);
and U28486 (N_28486,N_15166,N_10571);
and U28487 (N_28487,N_19576,N_15230);
or U28488 (N_28488,N_17191,N_16737);
nand U28489 (N_28489,N_19262,N_18881);
and U28490 (N_28490,N_16069,N_15467);
or U28491 (N_28491,N_12846,N_12572);
nand U28492 (N_28492,N_13559,N_17292);
nand U28493 (N_28493,N_17590,N_16309);
nand U28494 (N_28494,N_13208,N_11830);
nand U28495 (N_28495,N_10837,N_17386);
and U28496 (N_28496,N_18906,N_16256);
and U28497 (N_28497,N_17034,N_16148);
nand U28498 (N_28498,N_19361,N_13514);
and U28499 (N_28499,N_12021,N_12472);
and U28500 (N_28500,N_10351,N_18628);
or U28501 (N_28501,N_13909,N_12076);
xor U28502 (N_28502,N_12013,N_12073);
and U28503 (N_28503,N_19874,N_16537);
nor U28504 (N_28504,N_10098,N_16974);
and U28505 (N_28505,N_18799,N_12998);
xor U28506 (N_28506,N_12286,N_12822);
xor U28507 (N_28507,N_19475,N_14868);
and U28508 (N_28508,N_10613,N_11477);
or U28509 (N_28509,N_15403,N_14000);
nor U28510 (N_28510,N_12899,N_13533);
nor U28511 (N_28511,N_14530,N_15008);
and U28512 (N_28512,N_12726,N_11414);
or U28513 (N_28513,N_11314,N_16095);
and U28514 (N_28514,N_11348,N_13072);
xor U28515 (N_28515,N_12626,N_18059);
and U28516 (N_28516,N_11995,N_13897);
nand U28517 (N_28517,N_10779,N_17793);
xor U28518 (N_28518,N_19509,N_19280);
xor U28519 (N_28519,N_16687,N_12701);
and U28520 (N_28520,N_15243,N_12984);
and U28521 (N_28521,N_12296,N_13215);
nor U28522 (N_28522,N_10189,N_13770);
nor U28523 (N_28523,N_16792,N_15562);
nand U28524 (N_28524,N_11503,N_16035);
nor U28525 (N_28525,N_14125,N_19391);
nand U28526 (N_28526,N_19566,N_15007);
and U28527 (N_28527,N_10404,N_14119);
nand U28528 (N_28528,N_11444,N_18612);
nand U28529 (N_28529,N_19416,N_12845);
nand U28530 (N_28530,N_12722,N_19007);
and U28531 (N_28531,N_14692,N_14157);
nor U28532 (N_28532,N_10648,N_10128);
or U28533 (N_28533,N_14593,N_17363);
nor U28534 (N_28534,N_16669,N_19692);
and U28535 (N_28535,N_13667,N_19011);
or U28536 (N_28536,N_14383,N_10415);
nor U28537 (N_28537,N_14251,N_13421);
nor U28538 (N_28538,N_14058,N_16972);
and U28539 (N_28539,N_14421,N_17189);
or U28540 (N_28540,N_16128,N_10787);
or U28541 (N_28541,N_11388,N_17765);
and U28542 (N_28542,N_14780,N_10884);
nand U28543 (N_28543,N_19270,N_18801);
nor U28544 (N_28544,N_14829,N_14186);
nor U28545 (N_28545,N_19089,N_18299);
or U28546 (N_28546,N_15709,N_12011);
nor U28547 (N_28547,N_12180,N_16492);
xor U28548 (N_28548,N_12522,N_11000);
nor U28549 (N_28549,N_13103,N_12595);
nand U28550 (N_28550,N_16437,N_13225);
xnor U28551 (N_28551,N_17495,N_15280);
or U28552 (N_28552,N_17751,N_17261);
xnor U28553 (N_28553,N_14478,N_17910);
or U28554 (N_28554,N_13395,N_18213);
xor U28555 (N_28555,N_19456,N_19268);
nor U28556 (N_28556,N_14472,N_15032);
or U28557 (N_28557,N_12058,N_10207);
nor U28558 (N_28558,N_18900,N_14224);
nor U28559 (N_28559,N_11038,N_13379);
or U28560 (N_28560,N_15984,N_10308);
and U28561 (N_28561,N_13852,N_18963);
or U28562 (N_28562,N_13179,N_14990);
xnor U28563 (N_28563,N_12371,N_17892);
nand U28564 (N_28564,N_11581,N_16454);
or U28565 (N_28565,N_19760,N_17051);
nand U28566 (N_28566,N_19424,N_11725);
nor U28567 (N_28567,N_15365,N_15394);
xnor U28568 (N_28568,N_12562,N_14238);
and U28569 (N_28569,N_12025,N_19810);
nand U28570 (N_28570,N_11515,N_14243);
and U28571 (N_28571,N_14983,N_12452);
or U28572 (N_28572,N_11521,N_12584);
nor U28573 (N_28573,N_19983,N_19350);
nor U28574 (N_28574,N_15078,N_17902);
nor U28575 (N_28575,N_19064,N_10551);
and U28576 (N_28576,N_17411,N_19723);
nand U28577 (N_28577,N_18521,N_10556);
nand U28578 (N_28578,N_10962,N_11974);
nand U28579 (N_28579,N_10442,N_15630);
nor U28580 (N_28580,N_12445,N_12606);
nand U28581 (N_28581,N_19076,N_18391);
or U28582 (N_28582,N_13827,N_18758);
and U28583 (N_28583,N_11733,N_15247);
nor U28584 (N_28584,N_13990,N_11010);
nand U28585 (N_28585,N_19565,N_13503);
nor U28586 (N_28586,N_18557,N_11722);
and U28587 (N_28587,N_16642,N_17302);
nor U28588 (N_28588,N_13682,N_15554);
nor U28589 (N_28589,N_12769,N_10728);
or U28590 (N_28590,N_12848,N_16073);
nor U28591 (N_28591,N_14985,N_19435);
and U28592 (N_28592,N_17377,N_16524);
xor U28593 (N_28593,N_12182,N_16012);
and U28594 (N_28594,N_10051,N_15916);
or U28595 (N_28595,N_18317,N_14047);
and U28596 (N_28596,N_12158,N_14310);
nor U28597 (N_28597,N_19837,N_16323);
or U28598 (N_28598,N_11898,N_19671);
nor U28599 (N_28599,N_10627,N_12494);
and U28600 (N_28600,N_17814,N_18870);
nand U28601 (N_28601,N_10145,N_10252);
and U28602 (N_28602,N_18653,N_15081);
or U28603 (N_28603,N_13383,N_18302);
or U28604 (N_28604,N_19021,N_13013);
and U28605 (N_28605,N_14559,N_11159);
and U28606 (N_28606,N_14316,N_11083);
or U28607 (N_28607,N_14660,N_10117);
and U28608 (N_28608,N_15325,N_12187);
nor U28609 (N_28609,N_13942,N_15187);
nand U28610 (N_28610,N_18148,N_18168);
nor U28611 (N_28611,N_12299,N_11808);
nand U28612 (N_28612,N_14189,N_10157);
and U28613 (N_28613,N_15999,N_18108);
nand U28614 (N_28614,N_19850,N_13814);
and U28615 (N_28615,N_13617,N_14802);
and U28616 (N_28616,N_11617,N_11401);
nand U28617 (N_28617,N_15953,N_18643);
or U28618 (N_28618,N_12864,N_15317);
xor U28619 (N_28619,N_15031,N_15075);
nand U28620 (N_28620,N_12315,N_14731);
nor U28621 (N_28621,N_10225,N_11311);
and U28622 (N_28622,N_14541,N_19526);
xor U28623 (N_28623,N_13262,N_19345);
xor U28624 (N_28624,N_17353,N_14516);
nand U28625 (N_28625,N_18442,N_15673);
nand U28626 (N_28626,N_16998,N_19501);
or U28627 (N_28627,N_15346,N_10337);
and U28628 (N_28628,N_18876,N_17109);
and U28629 (N_28629,N_15687,N_11738);
and U28630 (N_28630,N_11095,N_11578);
nand U28631 (N_28631,N_13974,N_15143);
nor U28632 (N_28632,N_12167,N_13128);
nor U28633 (N_28633,N_17796,N_13536);
nor U28634 (N_28634,N_17472,N_15942);
or U28635 (N_28635,N_14956,N_17465);
or U28636 (N_28636,N_16793,N_12304);
and U28637 (N_28637,N_12151,N_19137);
or U28638 (N_28638,N_13462,N_11666);
and U28639 (N_28639,N_14179,N_13004);
or U28640 (N_28640,N_15927,N_16938);
and U28641 (N_28641,N_18936,N_11802);
nand U28642 (N_28642,N_19985,N_17932);
and U28643 (N_28643,N_13189,N_10732);
and U28644 (N_28644,N_15579,N_12577);
nor U28645 (N_28645,N_13979,N_15466);
and U28646 (N_28646,N_11952,N_10766);
or U28647 (N_28647,N_16428,N_13102);
nand U28648 (N_28648,N_10316,N_10418);
and U28649 (N_28649,N_16285,N_19003);
and U28650 (N_28650,N_14645,N_10227);
nor U28651 (N_28651,N_16916,N_12499);
or U28652 (N_28652,N_14040,N_10513);
nor U28653 (N_28653,N_18707,N_18188);
and U28654 (N_28654,N_13889,N_15013);
xnor U28655 (N_28655,N_14033,N_18302);
and U28656 (N_28656,N_19317,N_18509);
nor U28657 (N_28657,N_18268,N_18431);
and U28658 (N_28658,N_15973,N_14096);
nor U28659 (N_28659,N_17752,N_10599);
nand U28660 (N_28660,N_15795,N_11166);
or U28661 (N_28661,N_10443,N_11707);
or U28662 (N_28662,N_10672,N_14162);
nor U28663 (N_28663,N_13064,N_16778);
or U28664 (N_28664,N_14273,N_17395);
nor U28665 (N_28665,N_12022,N_11664);
or U28666 (N_28666,N_19366,N_17690);
or U28667 (N_28667,N_13310,N_13573);
and U28668 (N_28668,N_14873,N_14998);
nand U28669 (N_28669,N_16741,N_12244);
and U28670 (N_28670,N_13675,N_13990);
or U28671 (N_28671,N_19544,N_11149);
nor U28672 (N_28672,N_19452,N_15932);
or U28673 (N_28673,N_12086,N_13560);
xnor U28674 (N_28674,N_15300,N_14241);
nor U28675 (N_28675,N_19180,N_16710);
nor U28676 (N_28676,N_15447,N_12514);
xor U28677 (N_28677,N_13584,N_17790);
nor U28678 (N_28678,N_19965,N_10888);
and U28679 (N_28679,N_13408,N_18470);
or U28680 (N_28680,N_17746,N_11855);
or U28681 (N_28681,N_13350,N_14536);
nor U28682 (N_28682,N_17175,N_19589);
and U28683 (N_28683,N_17051,N_16507);
and U28684 (N_28684,N_18818,N_12450);
or U28685 (N_28685,N_11276,N_10068);
or U28686 (N_28686,N_17296,N_16202);
and U28687 (N_28687,N_16863,N_15123);
or U28688 (N_28688,N_15656,N_19899);
or U28689 (N_28689,N_10078,N_16761);
nor U28690 (N_28690,N_16164,N_12358);
and U28691 (N_28691,N_13306,N_10963);
nand U28692 (N_28692,N_11908,N_19289);
nand U28693 (N_28693,N_16145,N_19083);
nand U28694 (N_28694,N_11505,N_18783);
and U28695 (N_28695,N_17559,N_14752);
or U28696 (N_28696,N_15363,N_14055);
and U28697 (N_28697,N_16100,N_11150);
nand U28698 (N_28698,N_18513,N_10039);
nor U28699 (N_28699,N_18406,N_11276);
nor U28700 (N_28700,N_17714,N_15234);
nor U28701 (N_28701,N_16097,N_17779);
and U28702 (N_28702,N_15130,N_14189);
xor U28703 (N_28703,N_12102,N_16027);
nand U28704 (N_28704,N_10433,N_18422);
nor U28705 (N_28705,N_15357,N_14010);
nand U28706 (N_28706,N_13141,N_13709);
nand U28707 (N_28707,N_12127,N_10505);
or U28708 (N_28708,N_11892,N_12114);
nor U28709 (N_28709,N_19970,N_15018);
nor U28710 (N_28710,N_13935,N_17428);
xor U28711 (N_28711,N_12970,N_15791);
nor U28712 (N_28712,N_12554,N_17732);
nand U28713 (N_28713,N_11665,N_15122);
and U28714 (N_28714,N_12868,N_18925);
xnor U28715 (N_28715,N_15661,N_10450);
nand U28716 (N_28716,N_10537,N_10964);
nor U28717 (N_28717,N_16722,N_18610);
xor U28718 (N_28718,N_13026,N_11934);
xnor U28719 (N_28719,N_16109,N_18640);
or U28720 (N_28720,N_14647,N_17234);
and U28721 (N_28721,N_17072,N_11364);
or U28722 (N_28722,N_14540,N_16759);
and U28723 (N_28723,N_17470,N_11513);
nand U28724 (N_28724,N_17272,N_12623);
and U28725 (N_28725,N_11132,N_17371);
nand U28726 (N_28726,N_12569,N_18192);
nor U28727 (N_28727,N_15147,N_12959);
and U28728 (N_28728,N_10989,N_11274);
or U28729 (N_28729,N_19794,N_11954);
nand U28730 (N_28730,N_12572,N_15962);
or U28731 (N_28731,N_18233,N_17464);
or U28732 (N_28732,N_11904,N_15313);
or U28733 (N_28733,N_14374,N_16782);
nand U28734 (N_28734,N_15299,N_19128);
nand U28735 (N_28735,N_12707,N_16827);
nand U28736 (N_28736,N_16125,N_12776);
or U28737 (N_28737,N_18591,N_16661);
nor U28738 (N_28738,N_17949,N_14506);
nor U28739 (N_28739,N_18954,N_14165);
and U28740 (N_28740,N_13597,N_15383);
and U28741 (N_28741,N_10107,N_15168);
nand U28742 (N_28742,N_12735,N_10510);
nor U28743 (N_28743,N_10189,N_15268);
and U28744 (N_28744,N_12809,N_14157);
nor U28745 (N_28745,N_12124,N_12647);
and U28746 (N_28746,N_16818,N_19395);
and U28747 (N_28747,N_19843,N_17337);
xor U28748 (N_28748,N_15573,N_14038);
xnor U28749 (N_28749,N_16183,N_14716);
nor U28750 (N_28750,N_13469,N_19857);
nand U28751 (N_28751,N_17750,N_14388);
and U28752 (N_28752,N_16840,N_13991);
nand U28753 (N_28753,N_10980,N_12398);
or U28754 (N_28754,N_18130,N_19663);
and U28755 (N_28755,N_12763,N_14197);
nand U28756 (N_28756,N_10944,N_12484);
nor U28757 (N_28757,N_12076,N_12753);
and U28758 (N_28758,N_19958,N_16149);
xor U28759 (N_28759,N_15317,N_19166);
and U28760 (N_28760,N_19356,N_16381);
nor U28761 (N_28761,N_11602,N_19614);
nor U28762 (N_28762,N_13063,N_16668);
or U28763 (N_28763,N_10231,N_14782);
or U28764 (N_28764,N_11848,N_12741);
nand U28765 (N_28765,N_11723,N_19096);
nand U28766 (N_28766,N_16128,N_14673);
or U28767 (N_28767,N_13018,N_10842);
or U28768 (N_28768,N_14766,N_17672);
nor U28769 (N_28769,N_19177,N_19615);
nor U28770 (N_28770,N_10523,N_17427);
nand U28771 (N_28771,N_11305,N_12503);
and U28772 (N_28772,N_15595,N_14204);
xor U28773 (N_28773,N_15819,N_13758);
and U28774 (N_28774,N_14706,N_10223);
and U28775 (N_28775,N_11321,N_11151);
nor U28776 (N_28776,N_10682,N_16162);
or U28777 (N_28777,N_17785,N_17543);
xnor U28778 (N_28778,N_10092,N_11010);
xnor U28779 (N_28779,N_11674,N_15648);
or U28780 (N_28780,N_19922,N_17226);
nand U28781 (N_28781,N_14176,N_18085);
or U28782 (N_28782,N_10545,N_15972);
nor U28783 (N_28783,N_13481,N_19041);
xnor U28784 (N_28784,N_13973,N_12462);
nor U28785 (N_28785,N_12177,N_17130);
nor U28786 (N_28786,N_12504,N_18744);
xnor U28787 (N_28787,N_13427,N_12423);
or U28788 (N_28788,N_14918,N_11812);
or U28789 (N_28789,N_16779,N_16656);
nor U28790 (N_28790,N_17339,N_12402);
and U28791 (N_28791,N_19715,N_10286);
and U28792 (N_28792,N_16112,N_14760);
nor U28793 (N_28793,N_13868,N_14675);
and U28794 (N_28794,N_11040,N_13829);
and U28795 (N_28795,N_16802,N_17581);
nand U28796 (N_28796,N_15671,N_15254);
and U28797 (N_28797,N_11661,N_15710);
nand U28798 (N_28798,N_12997,N_17498);
or U28799 (N_28799,N_13926,N_12460);
or U28800 (N_28800,N_14364,N_14535);
nand U28801 (N_28801,N_13063,N_18118);
and U28802 (N_28802,N_16035,N_19563);
nor U28803 (N_28803,N_15491,N_19834);
nand U28804 (N_28804,N_17203,N_15359);
or U28805 (N_28805,N_15477,N_14666);
or U28806 (N_28806,N_18140,N_13964);
nor U28807 (N_28807,N_12885,N_13924);
nor U28808 (N_28808,N_13617,N_19713);
and U28809 (N_28809,N_11980,N_13317);
nor U28810 (N_28810,N_13155,N_17013);
and U28811 (N_28811,N_11114,N_14459);
nand U28812 (N_28812,N_15395,N_10413);
and U28813 (N_28813,N_14362,N_18364);
nor U28814 (N_28814,N_19358,N_13924);
or U28815 (N_28815,N_12635,N_19815);
or U28816 (N_28816,N_16520,N_18174);
nand U28817 (N_28817,N_14761,N_19795);
nor U28818 (N_28818,N_12281,N_16352);
nand U28819 (N_28819,N_14584,N_11767);
or U28820 (N_28820,N_10711,N_10740);
or U28821 (N_28821,N_11605,N_18639);
nand U28822 (N_28822,N_12924,N_18929);
nor U28823 (N_28823,N_18754,N_18686);
and U28824 (N_28824,N_13685,N_15501);
and U28825 (N_28825,N_11514,N_10666);
or U28826 (N_28826,N_11483,N_11478);
or U28827 (N_28827,N_11372,N_18825);
nor U28828 (N_28828,N_19724,N_17749);
and U28829 (N_28829,N_14928,N_15399);
nor U28830 (N_28830,N_11884,N_16980);
or U28831 (N_28831,N_11148,N_16659);
xor U28832 (N_28832,N_17410,N_12164);
and U28833 (N_28833,N_18748,N_16705);
and U28834 (N_28834,N_12712,N_13688);
and U28835 (N_28835,N_15658,N_12382);
nand U28836 (N_28836,N_17157,N_13033);
nor U28837 (N_28837,N_11824,N_16398);
nand U28838 (N_28838,N_12804,N_16765);
nor U28839 (N_28839,N_14491,N_10872);
nor U28840 (N_28840,N_10371,N_15839);
nor U28841 (N_28841,N_18682,N_16875);
and U28842 (N_28842,N_15634,N_19288);
and U28843 (N_28843,N_13110,N_18571);
or U28844 (N_28844,N_16616,N_13525);
and U28845 (N_28845,N_10130,N_10891);
nor U28846 (N_28846,N_12613,N_16275);
nand U28847 (N_28847,N_18002,N_19437);
nor U28848 (N_28848,N_11441,N_19592);
or U28849 (N_28849,N_11240,N_11620);
or U28850 (N_28850,N_10264,N_16907);
or U28851 (N_28851,N_16859,N_14275);
xnor U28852 (N_28852,N_12438,N_13533);
or U28853 (N_28853,N_18555,N_19323);
or U28854 (N_28854,N_14163,N_19882);
nand U28855 (N_28855,N_17080,N_18328);
nor U28856 (N_28856,N_19299,N_15942);
and U28857 (N_28857,N_14814,N_16029);
or U28858 (N_28858,N_13264,N_10596);
and U28859 (N_28859,N_17006,N_12630);
xnor U28860 (N_28860,N_17115,N_17107);
or U28861 (N_28861,N_15520,N_19087);
nand U28862 (N_28862,N_10757,N_16457);
nor U28863 (N_28863,N_14929,N_11130);
and U28864 (N_28864,N_10938,N_17689);
and U28865 (N_28865,N_13830,N_14871);
or U28866 (N_28866,N_13766,N_10455);
nand U28867 (N_28867,N_18103,N_17782);
and U28868 (N_28868,N_11294,N_12112);
xor U28869 (N_28869,N_14038,N_10936);
and U28870 (N_28870,N_12650,N_16363);
or U28871 (N_28871,N_17950,N_15368);
and U28872 (N_28872,N_12910,N_15646);
or U28873 (N_28873,N_12952,N_17503);
or U28874 (N_28874,N_18906,N_11679);
and U28875 (N_28875,N_19690,N_18527);
and U28876 (N_28876,N_16459,N_14737);
or U28877 (N_28877,N_19365,N_10410);
and U28878 (N_28878,N_13044,N_17956);
nor U28879 (N_28879,N_12693,N_11740);
nor U28880 (N_28880,N_10281,N_14629);
nor U28881 (N_28881,N_19794,N_15560);
nor U28882 (N_28882,N_15972,N_19240);
xor U28883 (N_28883,N_10007,N_14725);
nand U28884 (N_28884,N_12108,N_10406);
xor U28885 (N_28885,N_14345,N_10661);
and U28886 (N_28886,N_16545,N_11299);
nand U28887 (N_28887,N_16172,N_14365);
nor U28888 (N_28888,N_14164,N_15071);
xnor U28889 (N_28889,N_15999,N_14176);
and U28890 (N_28890,N_14095,N_18408);
nand U28891 (N_28891,N_17960,N_10177);
and U28892 (N_28892,N_13514,N_14490);
nor U28893 (N_28893,N_15178,N_10109);
nand U28894 (N_28894,N_17229,N_16974);
or U28895 (N_28895,N_13728,N_10795);
and U28896 (N_28896,N_18362,N_12722);
nand U28897 (N_28897,N_10692,N_15058);
nand U28898 (N_28898,N_19066,N_11131);
or U28899 (N_28899,N_16518,N_13054);
or U28900 (N_28900,N_17780,N_17532);
nand U28901 (N_28901,N_13565,N_19937);
and U28902 (N_28902,N_14693,N_15776);
and U28903 (N_28903,N_11357,N_15920);
nor U28904 (N_28904,N_14502,N_11778);
nand U28905 (N_28905,N_18230,N_12478);
or U28906 (N_28906,N_18955,N_18258);
or U28907 (N_28907,N_10603,N_11101);
xnor U28908 (N_28908,N_12473,N_10874);
xnor U28909 (N_28909,N_15405,N_17435);
xor U28910 (N_28910,N_15080,N_16429);
xor U28911 (N_28911,N_10461,N_16643);
nand U28912 (N_28912,N_15456,N_13898);
or U28913 (N_28913,N_17250,N_16179);
or U28914 (N_28914,N_11671,N_14589);
nor U28915 (N_28915,N_16712,N_12387);
and U28916 (N_28916,N_16259,N_14761);
or U28917 (N_28917,N_18352,N_16833);
or U28918 (N_28918,N_13239,N_14356);
and U28919 (N_28919,N_14122,N_11713);
and U28920 (N_28920,N_17465,N_13313);
nand U28921 (N_28921,N_15102,N_18238);
or U28922 (N_28922,N_18722,N_17263);
nor U28923 (N_28923,N_12306,N_16714);
and U28924 (N_28924,N_11146,N_13910);
or U28925 (N_28925,N_15835,N_12833);
xnor U28926 (N_28926,N_19142,N_13717);
nand U28927 (N_28927,N_18776,N_17872);
nor U28928 (N_28928,N_19217,N_17538);
nand U28929 (N_28929,N_19107,N_16886);
nand U28930 (N_28930,N_18847,N_13338);
nand U28931 (N_28931,N_16551,N_12150);
and U28932 (N_28932,N_17462,N_15061);
nor U28933 (N_28933,N_15465,N_15128);
nor U28934 (N_28934,N_12116,N_10427);
nor U28935 (N_28935,N_14725,N_14680);
nand U28936 (N_28936,N_17754,N_13134);
and U28937 (N_28937,N_12732,N_19651);
or U28938 (N_28938,N_17857,N_14368);
nand U28939 (N_28939,N_16851,N_19237);
nand U28940 (N_28940,N_11141,N_13456);
nor U28941 (N_28941,N_15022,N_19305);
nand U28942 (N_28942,N_13896,N_16708);
or U28943 (N_28943,N_13680,N_14684);
nor U28944 (N_28944,N_11898,N_13984);
nor U28945 (N_28945,N_11431,N_16517);
nor U28946 (N_28946,N_18090,N_13082);
nand U28947 (N_28947,N_19895,N_18930);
xnor U28948 (N_28948,N_18035,N_15212);
and U28949 (N_28949,N_12956,N_13987);
and U28950 (N_28950,N_11674,N_19061);
xnor U28951 (N_28951,N_17865,N_13834);
xor U28952 (N_28952,N_11965,N_10370);
and U28953 (N_28953,N_15781,N_17769);
or U28954 (N_28954,N_16569,N_17305);
xnor U28955 (N_28955,N_11354,N_16872);
or U28956 (N_28956,N_19559,N_18354);
nand U28957 (N_28957,N_14687,N_18350);
or U28958 (N_28958,N_17389,N_16864);
and U28959 (N_28959,N_16095,N_15011);
or U28960 (N_28960,N_14154,N_19809);
nor U28961 (N_28961,N_12973,N_11567);
nor U28962 (N_28962,N_16450,N_11354);
or U28963 (N_28963,N_15046,N_18023);
nand U28964 (N_28964,N_17644,N_18031);
and U28965 (N_28965,N_13370,N_17343);
nand U28966 (N_28966,N_18574,N_15635);
nor U28967 (N_28967,N_10253,N_10597);
or U28968 (N_28968,N_15718,N_13863);
and U28969 (N_28969,N_13880,N_12518);
nor U28970 (N_28970,N_15262,N_18315);
and U28971 (N_28971,N_10840,N_11449);
nor U28972 (N_28972,N_15483,N_10858);
or U28973 (N_28973,N_18970,N_12323);
nor U28974 (N_28974,N_12956,N_17534);
nand U28975 (N_28975,N_14851,N_11031);
nand U28976 (N_28976,N_14752,N_19371);
nor U28977 (N_28977,N_12577,N_18926);
or U28978 (N_28978,N_10828,N_11198);
nand U28979 (N_28979,N_14725,N_11734);
nor U28980 (N_28980,N_15157,N_13057);
and U28981 (N_28981,N_14459,N_11880);
or U28982 (N_28982,N_13621,N_10512);
or U28983 (N_28983,N_13944,N_15379);
nor U28984 (N_28984,N_10540,N_16239);
or U28985 (N_28985,N_15165,N_14263);
nor U28986 (N_28986,N_15533,N_17965);
xnor U28987 (N_28987,N_19799,N_10985);
nor U28988 (N_28988,N_12691,N_14993);
nand U28989 (N_28989,N_16054,N_10428);
and U28990 (N_28990,N_10552,N_12605);
nor U28991 (N_28991,N_15071,N_12592);
or U28992 (N_28992,N_14961,N_18614);
or U28993 (N_28993,N_13738,N_13466);
or U28994 (N_28994,N_14079,N_18000);
xor U28995 (N_28995,N_16598,N_18316);
nand U28996 (N_28996,N_19128,N_12883);
and U28997 (N_28997,N_17715,N_17947);
or U28998 (N_28998,N_17640,N_11676);
and U28999 (N_28999,N_16859,N_19293);
nor U29000 (N_29000,N_19216,N_17010);
nand U29001 (N_29001,N_15176,N_16775);
nand U29002 (N_29002,N_10129,N_13647);
xnor U29003 (N_29003,N_17795,N_17212);
xor U29004 (N_29004,N_14838,N_15429);
nand U29005 (N_29005,N_17212,N_14708);
nor U29006 (N_29006,N_16692,N_19550);
or U29007 (N_29007,N_17504,N_16335);
nor U29008 (N_29008,N_18988,N_11199);
nor U29009 (N_29009,N_17945,N_15548);
and U29010 (N_29010,N_14777,N_16803);
and U29011 (N_29011,N_16416,N_19011);
or U29012 (N_29012,N_10798,N_10314);
xnor U29013 (N_29013,N_10245,N_19364);
and U29014 (N_29014,N_17682,N_16392);
nand U29015 (N_29015,N_19785,N_19931);
and U29016 (N_29016,N_13864,N_10186);
nand U29017 (N_29017,N_19549,N_17022);
nor U29018 (N_29018,N_13111,N_14640);
and U29019 (N_29019,N_16738,N_16599);
nand U29020 (N_29020,N_10422,N_19972);
and U29021 (N_29021,N_11338,N_13479);
nand U29022 (N_29022,N_15620,N_12119);
xnor U29023 (N_29023,N_16106,N_11657);
nor U29024 (N_29024,N_19909,N_11383);
xnor U29025 (N_29025,N_15759,N_14485);
nor U29026 (N_29026,N_17077,N_17913);
or U29027 (N_29027,N_10849,N_15785);
nor U29028 (N_29028,N_10387,N_19273);
and U29029 (N_29029,N_11284,N_15892);
and U29030 (N_29030,N_14670,N_12339);
nor U29031 (N_29031,N_10113,N_13023);
and U29032 (N_29032,N_15614,N_19925);
and U29033 (N_29033,N_16176,N_18615);
and U29034 (N_29034,N_10354,N_10394);
or U29035 (N_29035,N_18111,N_18327);
and U29036 (N_29036,N_12114,N_12305);
and U29037 (N_29037,N_10230,N_13877);
and U29038 (N_29038,N_11492,N_13587);
xnor U29039 (N_29039,N_11637,N_19667);
and U29040 (N_29040,N_16224,N_10275);
or U29041 (N_29041,N_11126,N_13931);
nand U29042 (N_29042,N_15378,N_19485);
nor U29043 (N_29043,N_18522,N_13526);
xor U29044 (N_29044,N_10533,N_18325);
xor U29045 (N_29045,N_14331,N_15842);
or U29046 (N_29046,N_12492,N_13349);
or U29047 (N_29047,N_17083,N_10217);
or U29048 (N_29048,N_12333,N_13824);
or U29049 (N_29049,N_13119,N_17821);
and U29050 (N_29050,N_15070,N_11170);
nand U29051 (N_29051,N_15220,N_19326);
nand U29052 (N_29052,N_16466,N_12084);
and U29053 (N_29053,N_19625,N_17421);
or U29054 (N_29054,N_11925,N_17147);
nand U29055 (N_29055,N_11684,N_15085);
and U29056 (N_29056,N_17265,N_14863);
or U29057 (N_29057,N_17460,N_14425);
nor U29058 (N_29058,N_11137,N_14017);
xor U29059 (N_29059,N_19109,N_10579);
nand U29060 (N_29060,N_17790,N_11455);
nand U29061 (N_29061,N_13206,N_16398);
nor U29062 (N_29062,N_10779,N_19623);
nand U29063 (N_29063,N_11186,N_19587);
nor U29064 (N_29064,N_13994,N_16906);
and U29065 (N_29065,N_15771,N_18556);
xnor U29066 (N_29066,N_18551,N_15589);
and U29067 (N_29067,N_17522,N_16976);
and U29068 (N_29068,N_18650,N_17910);
nor U29069 (N_29069,N_15681,N_17405);
or U29070 (N_29070,N_18829,N_16774);
nand U29071 (N_29071,N_19495,N_18685);
nor U29072 (N_29072,N_10686,N_13655);
or U29073 (N_29073,N_19012,N_12250);
and U29074 (N_29074,N_10443,N_14148);
nand U29075 (N_29075,N_13016,N_11281);
nor U29076 (N_29076,N_16466,N_16684);
or U29077 (N_29077,N_10951,N_13182);
and U29078 (N_29078,N_14877,N_17358);
and U29079 (N_29079,N_10923,N_10534);
nor U29080 (N_29080,N_10763,N_17036);
or U29081 (N_29081,N_14319,N_12865);
and U29082 (N_29082,N_18924,N_10273);
and U29083 (N_29083,N_16621,N_16394);
and U29084 (N_29084,N_15718,N_16096);
or U29085 (N_29085,N_18339,N_17986);
nor U29086 (N_29086,N_12025,N_11020);
nor U29087 (N_29087,N_11225,N_14483);
or U29088 (N_29088,N_15211,N_11242);
nand U29089 (N_29089,N_16254,N_11857);
nor U29090 (N_29090,N_18574,N_11659);
nor U29091 (N_29091,N_12803,N_17367);
and U29092 (N_29092,N_16938,N_13664);
nand U29093 (N_29093,N_14626,N_14099);
nor U29094 (N_29094,N_18215,N_15645);
or U29095 (N_29095,N_16808,N_14839);
nor U29096 (N_29096,N_12101,N_15875);
nand U29097 (N_29097,N_11792,N_19110);
nor U29098 (N_29098,N_17744,N_14682);
nor U29099 (N_29099,N_10761,N_12501);
nor U29100 (N_29100,N_18184,N_10065);
and U29101 (N_29101,N_12547,N_12984);
nor U29102 (N_29102,N_18871,N_15831);
or U29103 (N_29103,N_14706,N_11516);
nand U29104 (N_29104,N_14624,N_16604);
nor U29105 (N_29105,N_14149,N_14525);
nand U29106 (N_29106,N_11682,N_12025);
nand U29107 (N_29107,N_12085,N_17262);
or U29108 (N_29108,N_15498,N_17440);
nand U29109 (N_29109,N_15501,N_18132);
and U29110 (N_29110,N_14042,N_18945);
nand U29111 (N_29111,N_17360,N_14420);
nand U29112 (N_29112,N_10402,N_13391);
nand U29113 (N_29113,N_18938,N_15925);
nor U29114 (N_29114,N_12627,N_10447);
and U29115 (N_29115,N_10180,N_17523);
or U29116 (N_29116,N_11023,N_18044);
and U29117 (N_29117,N_15895,N_15567);
and U29118 (N_29118,N_13433,N_19269);
xnor U29119 (N_29119,N_13069,N_15793);
nor U29120 (N_29120,N_12037,N_17565);
and U29121 (N_29121,N_12343,N_19156);
and U29122 (N_29122,N_15271,N_12197);
or U29123 (N_29123,N_18809,N_13628);
and U29124 (N_29124,N_14064,N_19283);
and U29125 (N_29125,N_13277,N_10358);
and U29126 (N_29126,N_19659,N_10698);
nor U29127 (N_29127,N_18979,N_10543);
and U29128 (N_29128,N_19892,N_11446);
nor U29129 (N_29129,N_16224,N_14790);
nand U29130 (N_29130,N_13192,N_11082);
or U29131 (N_29131,N_13551,N_17083);
nor U29132 (N_29132,N_14964,N_11474);
nand U29133 (N_29133,N_10872,N_10731);
and U29134 (N_29134,N_14797,N_18197);
and U29135 (N_29135,N_12376,N_11655);
nand U29136 (N_29136,N_19744,N_12936);
nor U29137 (N_29137,N_14408,N_10321);
xor U29138 (N_29138,N_13508,N_13702);
and U29139 (N_29139,N_16018,N_18559);
nand U29140 (N_29140,N_19010,N_11918);
and U29141 (N_29141,N_12364,N_16650);
nand U29142 (N_29142,N_13838,N_11581);
nand U29143 (N_29143,N_17479,N_13265);
and U29144 (N_29144,N_16116,N_16388);
nand U29145 (N_29145,N_16042,N_12870);
and U29146 (N_29146,N_18055,N_12699);
nand U29147 (N_29147,N_17865,N_17572);
and U29148 (N_29148,N_17971,N_13385);
nor U29149 (N_29149,N_17236,N_17594);
and U29150 (N_29150,N_18249,N_10897);
or U29151 (N_29151,N_13100,N_11927);
and U29152 (N_29152,N_10078,N_14521);
nand U29153 (N_29153,N_16982,N_13359);
nand U29154 (N_29154,N_11607,N_18287);
xor U29155 (N_29155,N_15325,N_14750);
nor U29156 (N_29156,N_14141,N_17620);
nand U29157 (N_29157,N_19855,N_15431);
or U29158 (N_29158,N_15047,N_14688);
nand U29159 (N_29159,N_18908,N_11522);
and U29160 (N_29160,N_14478,N_13575);
and U29161 (N_29161,N_15790,N_18554);
xor U29162 (N_29162,N_11879,N_19121);
or U29163 (N_29163,N_14957,N_15872);
or U29164 (N_29164,N_12027,N_12928);
or U29165 (N_29165,N_16245,N_16855);
nor U29166 (N_29166,N_13723,N_14732);
nand U29167 (N_29167,N_18420,N_16938);
and U29168 (N_29168,N_19936,N_17513);
or U29169 (N_29169,N_11207,N_11720);
or U29170 (N_29170,N_11511,N_11768);
or U29171 (N_29171,N_16029,N_17636);
xor U29172 (N_29172,N_17730,N_19060);
nor U29173 (N_29173,N_12639,N_17774);
or U29174 (N_29174,N_11467,N_11571);
nor U29175 (N_29175,N_10019,N_12055);
xnor U29176 (N_29176,N_14036,N_16137);
or U29177 (N_29177,N_15065,N_18265);
or U29178 (N_29178,N_11333,N_11962);
nor U29179 (N_29179,N_15302,N_11309);
and U29180 (N_29180,N_11262,N_12494);
and U29181 (N_29181,N_12917,N_18602);
or U29182 (N_29182,N_10122,N_15242);
or U29183 (N_29183,N_16005,N_13108);
or U29184 (N_29184,N_17878,N_15144);
nor U29185 (N_29185,N_17686,N_14079);
nor U29186 (N_29186,N_10086,N_13351);
and U29187 (N_29187,N_16914,N_16139);
and U29188 (N_29188,N_19486,N_15705);
or U29189 (N_29189,N_11634,N_17986);
nand U29190 (N_29190,N_19832,N_17855);
and U29191 (N_29191,N_18433,N_18958);
and U29192 (N_29192,N_19510,N_19526);
and U29193 (N_29193,N_11923,N_13145);
nand U29194 (N_29194,N_15203,N_11486);
nor U29195 (N_29195,N_17495,N_15399);
nor U29196 (N_29196,N_19803,N_14464);
nand U29197 (N_29197,N_15146,N_13736);
nor U29198 (N_29198,N_12369,N_11003);
and U29199 (N_29199,N_11084,N_16717);
nand U29200 (N_29200,N_12955,N_18050);
nor U29201 (N_29201,N_18308,N_10771);
and U29202 (N_29202,N_18479,N_12123);
and U29203 (N_29203,N_18555,N_16578);
and U29204 (N_29204,N_18693,N_17775);
nor U29205 (N_29205,N_12707,N_13585);
or U29206 (N_29206,N_14542,N_16423);
nand U29207 (N_29207,N_11905,N_12467);
nor U29208 (N_29208,N_12145,N_12467);
xor U29209 (N_29209,N_15405,N_17639);
nor U29210 (N_29210,N_12588,N_13474);
or U29211 (N_29211,N_13374,N_18567);
and U29212 (N_29212,N_16203,N_17643);
nor U29213 (N_29213,N_10524,N_19341);
or U29214 (N_29214,N_16080,N_15285);
nor U29215 (N_29215,N_14708,N_19167);
xor U29216 (N_29216,N_10194,N_12667);
and U29217 (N_29217,N_17671,N_17674);
and U29218 (N_29218,N_17770,N_15743);
and U29219 (N_29219,N_19351,N_11545);
nand U29220 (N_29220,N_16486,N_12520);
and U29221 (N_29221,N_11919,N_14717);
nand U29222 (N_29222,N_18759,N_18090);
nand U29223 (N_29223,N_15927,N_16841);
nand U29224 (N_29224,N_19174,N_11149);
or U29225 (N_29225,N_11619,N_11369);
nand U29226 (N_29226,N_15466,N_19916);
xor U29227 (N_29227,N_16039,N_13633);
xor U29228 (N_29228,N_17718,N_18720);
nor U29229 (N_29229,N_12366,N_18215);
xor U29230 (N_29230,N_15369,N_10300);
and U29231 (N_29231,N_13002,N_19622);
or U29232 (N_29232,N_17222,N_16989);
nor U29233 (N_29233,N_10651,N_12104);
or U29234 (N_29234,N_11594,N_15160);
or U29235 (N_29235,N_17750,N_18633);
nor U29236 (N_29236,N_18725,N_16466);
or U29237 (N_29237,N_17911,N_15166);
nand U29238 (N_29238,N_11147,N_10766);
nor U29239 (N_29239,N_19923,N_18265);
nor U29240 (N_29240,N_19019,N_14004);
and U29241 (N_29241,N_13532,N_16851);
or U29242 (N_29242,N_17051,N_12068);
xor U29243 (N_29243,N_11260,N_11553);
or U29244 (N_29244,N_11644,N_13788);
nand U29245 (N_29245,N_10888,N_13112);
and U29246 (N_29246,N_12142,N_13713);
nand U29247 (N_29247,N_10537,N_10137);
and U29248 (N_29248,N_14796,N_16974);
nor U29249 (N_29249,N_14335,N_12449);
nand U29250 (N_29250,N_13752,N_12401);
nor U29251 (N_29251,N_10512,N_19476);
nor U29252 (N_29252,N_10533,N_11407);
nor U29253 (N_29253,N_10902,N_14378);
nor U29254 (N_29254,N_15714,N_12595);
xor U29255 (N_29255,N_10596,N_11897);
xor U29256 (N_29256,N_19559,N_10427);
and U29257 (N_29257,N_12809,N_14910);
xnor U29258 (N_29258,N_18379,N_13417);
nor U29259 (N_29259,N_14292,N_10448);
xor U29260 (N_29260,N_11396,N_12855);
and U29261 (N_29261,N_10669,N_19113);
and U29262 (N_29262,N_15081,N_13417);
and U29263 (N_29263,N_17606,N_11517);
nand U29264 (N_29264,N_15435,N_19299);
nor U29265 (N_29265,N_15935,N_16216);
and U29266 (N_29266,N_19306,N_12098);
and U29267 (N_29267,N_11477,N_19764);
xor U29268 (N_29268,N_18936,N_18236);
or U29269 (N_29269,N_18734,N_13957);
xnor U29270 (N_29270,N_13786,N_14486);
and U29271 (N_29271,N_12491,N_18518);
nand U29272 (N_29272,N_12155,N_16059);
nor U29273 (N_29273,N_18790,N_13516);
nor U29274 (N_29274,N_10580,N_17335);
nand U29275 (N_29275,N_14506,N_19171);
or U29276 (N_29276,N_16689,N_11031);
xor U29277 (N_29277,N_11195,N_14054);
nor U29278 (N_29278,N_15308,N_10830);
nor U29279 (N_29279,N_19156,N_18577);
and U29280 (N_29280,N_12829,N_16227);
nor U29281 (N_29281,N_12304,N_10062);
or U29282 (N_29282,N_17236,N_15347);
or U29283 (N_29283,N_15593,N_11306);
nand U29284 (N_29284,N_12177,N_16273);
nand U29285 (N_29285,N_19424,N_10483);
nand U29286 (N_29286,N_10133,N_13607);
xor U29287 (N_29287,N_18185,N_14643);
and U29288 (N_29288,N_15548,N_16619);
nor U29289 (N_29289,N_19905,N_18762);
nand U29290 (N_29290,N_18497,N_15854);
nand U29291 (N_29291,N_18833,N_11633);
nor U29292 (N_29292,N_16336,N_19877);
nor U29293 (N_29293,N_11778,N_17078);
xor U29294 (N_29294,N_14964,N_18479);
or U29295 (N_29295,N_11993,N_17415);
or U29296 (N_29296,N_17461,N_18533);
xor U29297 (N_29297,N_13619,N_18530);
nor U29298 (N_29298,N_13968,N_17858);
nor U29299 (N_29299,N_11569,N_19162);
xnor U29300 (N_29300,N_12930,N_10684);
nor U29301 (N_29301,N_14097,N_13590);
nand U29302 (N_29302,N_14534,N_18046);
or U29303 (N_29303,N_14246,N_15697);
or U29304 (N_29304,N_16318,N_11515);
and U29305 (N_29305,N_19771,N_13099);
nand U29306 (N_29306,N_16927,N_13056);
and U29307 (N_29307,N_15974,N_10961);
nor U29308 (N_29308,N_18109,N_10357);
nor U29309 (N_29309,N_11945,N_16029);
xnor U29310 (N_29310,N_19481,N_19871);
or U29311 (N_29311,N_15555,N_14640);
and U29312 (N_29312,N_19565,N_18459);
xor U29313 (N_29313,N_16227,N_18546);
nand U29314 (N_29314,N_15550,N_15386);
nand U29315 (N_29315,N_14453,N_14007);
or U29316 (N_29316,N_16836,N_19653);
or U29317 (N_29317,N_14753,N_11314);
and U29318 (N_29318,N_12848,N_15530);
and U29319 (N_29319,N_14959,N_12597);
nand U29320 (N_29320,N_16201,N_13500);
nand U29321 (N_29321,N_15004,N_18667);
xnor U29322 (N_29322,N_16214,N_17785);
or U29323 (N_29323,N_10473,N_10039);
and U29324 (N_29324,N_14822,N_12273);
and U29325 (N_29325,N_15781,N_16990);
nand U29326 (N_29326,N_16725,N_10635);
or U29327 (N_29327,N_14468,N_12444);
nand U29328 (N_29328,N_11566,N_18867);
nor U29329 (N_29329,N_13255,N_15062);
or U29330 (N_29330,N_18462,N_12734);
or U29331 (N_29331,N_16266,N_19790);
nand U29332 (N_29332,N_13993,N_19070);
and U29333 (N_29333,N_13831,N_10455);
or U29334 (N_29334,N_10672,N_15477);
or U29335 (N_29335,N_16047,N_18961);
xor U29336 (N_29336,N_12558,N_16555);
and U29337 (N_29337,N_18947,N_12374);
or U29338 (N_29338,N_13366,N_10088);
and U29339 (N_29339,N_15499,N_12419);
nor U29340 (N_29340,N_14790,N_17911);
nor U29341 (N_29341,N_19297,N_13441);
nand U29342 (N_29342,N_17526,N_15788);
nor U29343 (N_29343,N_12570,N_15449);
or U29344 (N_29344,N_15923,N_15854);
nor U29345 (N_29345,N_18029,N_15577);
nor U29346 (N_29346,N_10864,N_18104);
and U29347 (N_29347,N_16029,N_19391);
nand U29348 (N_29348,N_19965,N_17614);
nor U29349 (N_29349,N_12303,N_10652);
xor U29350 (N_29350,N_16369,N_11565);
xor U29351 (N_29351,N_17517,N_18793);
or U29352 (N_29352,N_11617,N_10248);
or U29353 (N_29353,N_14744,N_14920);
and U29354 (N_29354,N_17607,N_13075);
nor U29355 (N_29355,N_19584,N_14740);
nor U29356 (N_29356,N_11931,N_10817);
nor U29357 (N_29357,N_11242,N_16316);
nor U29358 (N_29358,N_18386,N_14678);
nand U29359 (N_29359,N_15697,N_14585);
xor U29360 (N_29360,N_13324,N_16330);
nor U29361 (N_29361,N_12809,N_14423);
xor U29362 (N_29362,N_18733,N_19119);
or U29363 (N_29363,N_12807,N_18088);
or U29364 (N_29364,N_14986,N_10876);
and U29365 (N_29365,N_13292,N_18863);
and U29366 (N_29366,N_18506,N_17338);
nand U29367 (N_29367,N_12113,N_19293);
or U29368 (N_29368,N_17221,N_18424);
nand U29369 (N_29369,N_16524,N_10596);
or U29370 (N_29370,N_15173,N_16316);
nor U29371 (N_29371,N_13365,N_18549);
nor U29372 (N_29372,N_15230,N_19323);
nand U29373 (N_29373,N_10397,N_16797);
nor U29374 (N_29374,N_12078,N_19311);
or U29375 (N_29375,N_12178,N_17556);
and U29376 (N_29376,N_17686,N_12796);
or U29377 (N_29377,N_12616,N_17025);
nand U29378 (N_29378,N_18325,N_17252);
xnor U29379 (N_29379,N_13955,N_11392);
or U29380 (N_29380,N_15765,N_11158);
nor U29381 (N_29381,N_19863,N_15110);
and U29382 (N_29382,N_16882,N_17694);
nand U29383 (N_29383,N_15118,N_12375);
nor U29384 (N_29384,N_13633,N_19948);
nor U29385 (N_29385,N_19052,N_10608);
xnor U29386 (N_29386,N_12767,N_17352);
or U29387 (N_29387,N_11437,N_10313);
or U29388 (N_29388,N_10321,N_13125);
or U29389 (N_29389,N_18589,N_12201);
and U29390 (N_29390,N_11499,N_17209);
nor U29391 (N_29391,N_14310,N_15393);
nor U29392 (N_29392,N_17097,N_18125);
nand U29393 (N_29393,N_16884,N_16302);
and U29394 (N_29394,N_10601,N_18547);
nand U29395 (N_29395,N_17322,N_18023);
nor U29396 (N_29396,N_18406,N_14453);
nand U29397 (N_29397,N_19748,N_19744);
nand U29398 (N_29398,N_16335,N_17808);
nand U29399 (N_29399,N_14215,N_13336);
nor U29400 (N_29400,N_14330,N_13008);
nand U29401 (N_29401,N_14117,N_10190);
nand U29402 (N_29402,N_14631,N_13485);
nand U29403 (N_29403,N_15684,N_13208);
nor U29404 (N_29404,N_17414,N_19165);
or U29405 (N_29405,N_15115,N_15178);
nand U29406 (N_29406,N_11890,N_19231);
and U29407 (N_29407,N_13490,N_13637);
nand U29408 (N_29408,N_18234,N_19278);
nor U29409 (N_29409,N_18309,N_15785);
or U29410 (N_29410,N_11054,N_17640);
or U29411 (N_29411,N_13845,N_15844);
and U29412 (N_29412,N_18101,N_13774);
or U29413 (N_29413,N_10667,N_14160);
and U29414 (N_29414,N_15708,N_14921);
xor U29415 (N_29415,N_11625,N_16514);
and U29416 (N_29416,N_14893,N_13486);
nand U29417 (N_29417,N_17765,N_10896);
nor U29418 (N_29418,N_16646,N_18749);
and U29419 (N_29419,N_11506,N_12232);
xor U29420 (N_29420,N_18200,N_10497);
or U29421 (N_29421,N_11052,N_17600);
nand U29422 (N_29422,N_16093,N_18851);
nand U29423 (N_29423,N_19642,N_15046);
xor U29424 (N_29424,N_14953,N_12737);
nand U29425 (N_29425,N_16504,N_12004);
nor U29426 (N_29426,N_14893,N_18206);
nor U29427 (N_29427,N_15307,N_11033);
and U29428 (N_29428,N_14714,N_18204);
nand U29429 (N_29429,N_10662,N_16035);
xor U29430 (N_29430,N_16380,N_10918);
or U29431 (N_29431,N_10192,N_11806);
nor U29432 (N_29432,N_19275,N_11138);
and U29433 (N_29433,N_17409,N_18381);
or U29434 (N_29434,N_11306,N_16401);
and U29435 (N_29435,N_13747,N_11263);
and U29436 (N_29436,N_19924,N_13704);
or U29437 (N_29437,N_15520,N_18659);
and U29438 (N_29438,N_16359,N_18676);
nand U29439 (N_29439,N_17461,N_15739);
xor U29440 (N_29440,N_19782,N_11019);
and U29441 (N_29441,N_17714,N_17898);
nor U29442 (N_29442,N_16374,N_19747);
nand U29443 (N_29443,N_18715,N_17031);
nand U29444 (N_29444,N_10084,N_13095);
nand U29445 (N_29445,N_10895,N_13451);
or U29446 (N_29446,N_16238,N_17759);
nand U29447 (N_29447,N_18980,N_19753);
nand U29448 (N_29448,N_19969,N_15722);
nand U29449 (N_29449,N_13039,N_16176);
nor U29450 (N_29450,N_15514,N_19609);
nor U29451 (N_29451,N_13294,N_12813);
nor U29452 (N_29452,N_17819,N_12255);
or U29453 (N_29453,N_17096,N_16919);
xnor U29454 (N_29454,N_13434,N_15303);
and U29455 (N_29455,N_10195,N_16494);
nor U29456 (N_29456,N_15922,N_11994);
or U29457 (N_29457,N_18380,N_18189);
or U29458 (N_29458,N_17455,N_16301);
nor U29459 (N_29459,N_12900,N_12613);
or U29460 (N_29460,N_16984,N_18294);
and U29461 (N_29461,N_15320,N_11823);
nand U29462 (N_29462,N_18417,N_18786);
xor U29463 (N_29463,N_11151,N_16919);
and U29464 (N_29464,N_14618,N_17410);
and U29465 (N_29465,N_16843,N_15695);
or U29466 (N_29466,N_13520,N_17670);
nor U29467 (N_29467,N_13649,N_14105);
or U29468 (N_29468,N_18548,N_18611);
and U29469 (N_29469,N_15473,N_18265);
xnor U29470 (N_29470,N_10487,N_15282);
or U29471 (N_29471,N_14875,N_14659);
or U29472 (N_29472,N_13542,N_16851);
nand U29473 (N_29473,N_11890,N_12676);
or U29474 (N_29474,N_19666,N_11148);
nor U29475 (N_29475,N_13359,N_13310);
and U29476 (N_29476,N_18282,N_11671);
nor U29477 (N_29477,N_14615,N_15917);
nor U29478 (N_29478,N_11928,N_14250);
nand U29479 (N_29479,N_16254,N_14067);
xor U29480 (N_29480,N_18174,N_16226);
and U29481 (N_29481,N_12080,N_16724);
nor U29482 (N_29482,N_17518,N_16049);
xnor U29483 (N_29483,N_19995,N_16513);
xnor U29484 (N_29484,N_15443,N_11037);
or U29485 (N_29485,N_11701,N_17634);
nor U29486 (N_29486,N_16524,N_17185);
or U29487 (N_29487,N_16809,N_15859);
nor U29488 (N_29488,N_19725,N_11250);
nand U29489 (N_29489,N_17686,N_12738);
nand U29490 (N_29490,N_11220,N_12867);
or U29491 (N_29491,N_17062,N_13033);
nor U29492 (N_29492,N_12464,N_17647);
and U29493 (N_29493,N_14668,N_17896);
xnor U29494 (N_29494,N_13078,N_10097);
nand U29495 (N_29495,N_19342,N_17997);
nor U29496 (N_29496,N_15053,N_11520);
xnor U29497 (N_29497,N_14117,N_19504);
or U29498 (N_29498,N_11590,N_14749);
or U29499 (N_29499,N_11906,N_14832);
or U29500 (N_29500,N_12426,N_16768);
nor U29501 (N_29501,N_14489,N_15972);
nor U29502 (N_29502,N_18415,N_13788);
and U29503 (N_29503,N_18291,N_18726);
or U29504 (N_29504,N_19336,N_12796);
or U29505 (N_29505,N_15899,N_13024);
and U29506 (N_29506,N_13890,N_18747);
or U29507 (N_29507,N_16828,N_11348);
nor U29508 (N_29508,N_19205,N_14065);
and U29509 (N_29509,N_12049,N_19750);
or U29510 (N_29510,N_19130,N_19810);
and U29511 (N_29511,N_19756,N_11144);
and U29512 (N_29512,N_11359,N_19327);
nand U29513 (N_29513,N_19832,N_17323);
nor U29514 (N_29514,N_14716,N_11142);
nor U29515 (N_29515,N_15069,N_13832);
and U29516 (N_29516,N_10505,N_13389);
and U29517 (N_29517,N_19730,N_15984);
and U29518 (N_29518,N_12553,N_19919);
nand U29519 (N_29519,N_14783,N_10195);
or U29520 (N_29520,N_10272,N_14203);
or U29521 (N_29521,N_16095,N_10924);
or U29522 (N_29522,N_10072,N_12496);
nor U29523 (N_29523,N_19240,N_18774);
or U29524 (N_29524,N_15027,N_13721);
nor U29525 (N_29525,N_17248,N_16212);
nand U29526 (N_29526,N_19396,N_11200);
or U29527 (N_29527,N_19067,N_14611);
or U29528 (N_29528,N_13394,N_12385);
or U29529 (N_29529,N_12773,N_11415);
and U29530 (N_29530,N_15267,N_15100);
and U29531 (N_29531,N_16136,N_13518);
xnor U29532 (N_29532,N_14705,N_17109);
nor U29533 (N_29533,N_19095,N_14724);
xor U29534 (N_29534,N_16905,N_17052);
and U29535 (N_29535,N_12353,N_14613);
nor U29536 (N_29536,N_17212,N_17046);
nor U29537 (N_29537,N_15610,N_15695);
or U29538 (N_29538,N_15336,N_19184);
nor U29539 (N_29539,N_11212,N_11440);
nand U29540 (N_29540,N_17946,N_17624);
nor U29541 (N_29541,N_13215,N_18667);
xnor U29542 (N_29542,N_15660,N_17690);
xor U29543 (N_29543,N_13262,N_18113);
nor U29544 (N_29544,N_16152,N_18525);
nand U29545 (N_29545,N_19321,N_10948);
xor U29546 (N_29546,N_11635,N_11954);
nor U29547 (N_29547,N_17092,N_13187);
xor U29548 (N_29548,N_17492,N_12315);
or U29549 (N_29549,N_12354,N_11936);
and U29550 (N_29550,N_16810,N_13313);
nand U29551 (N_29551,N_17272,N_12418);
nand U29552 (N_29552,N_18692,N_11493);
and U29553 (N_29553,N_11080,N_16620);
nor U29554 (N_29554,N_19801,N_12199);
nor U29555 (N_29555,N_15901,N_17581);
xnor U29556 (N_29556,N_16018,N_14658);
and U29557 (N_29557,N_15876,N_13032);
or U29558 (N_29558,N_11208,N_16877);
or U29559 (N_29559,N_13622,N_18072);
nand U29560 (N_29560,N_15746,N_11435);
nor U29561 (N_29561,N_15444,N_13254);
or U29562 (N_29562,N_16722,N_14463);
and U29563 (N_29563,N_18254,N_16778);
or U29564 (N_29564,N_12307,N_17103);
nor U29565 (N_29565,N_18344,N_16084);
or U29566 (N_29566,N_10341,N_14705);
and U29567 (N_29567,N_14723,N_13797);
nand U29568 (N_29568,N_17793,N_15920);
nor U29569 (N_29569,N_16359,N_16236);
nand U29570 (N_29570,N_12474,N_16360);
and U29571 (N_29571,N_15462,N_18520);
nand U29572 (N_29572,N_10707,N_13396);
nor U29573 (N_29573,N_15653,N_14174);
nor U29574 (N_29574,N_16686,N_17006);
or U29575 (N_29575,N_17772,N_13930);
xor U29576 (N_29576,N_19521,N_19296);
nand U29577 (N_29577,N_11471,N_10584);
and U29578 (N_29578,N_19331,N_14416);
and U29579 (N_29579,N_14472,N_11203);
nand U29580 (N_29580,N_15481,N_10712);
nand U29581 (N_29581,N_19327,N_16953);
or U29582 (N_29582,N_13807,N_19013);
nand U29583 (N_29583,N_16212,N_12172);
nand U29584 (N_29584,N_15086,N_13687);
nand U29585 (N_29585,N_18641,N_14010);
nor U29586 (N_29586,N_15482,N_10873);
or U29587 (N_29587,N_17772,N_19099);
xor U29588 (N_29588,N_14341,N_11254);
and U29589 (N_29589,N_19551,N_15651);
nor U29590 (N_29590,N_10996,N_18717);
and U29591 (N_29591,N_16556,N_14666);
or U29592 (N_29592,N_17899,N_16873);
and U29593 (N_29593,N_19750,N_18352);
nor U29594 (N_29594,N_14567,N_14797);
and U29595 (N_29595,N_10923,N_13833);
nor U29596 (N_29596,N_15774,N_18513);
xor U29597 (N_29597,N_13489,N_16772);
and U29598 (N_29598,N_14183,N_16983);
nor U29599 (N_29599,N_11697,N_10217);
and U29600 (N_29600,N_18248,N_14378);
nor U29601 (N_29601,N_17616,N_15142);
nor U29602 (N_29602,N_10488,N_12800);
nor U29603 (N_29603,N_12717,N_14392);
nor U29604 (N_29604,N_12184,N_16633);
and U29605 (N_29605,N_13175,N_14947);
nor U29606 (N_29606,N_11625,N_18879);
and U29607 (N_29607,N_19695,N_14054);
and U29608 (N_29608,N_13875,N_18266);
nor U29609 (N_29609,N_16422,N_16019);
or U29610 (N_29610,N_19691,N_12505);
nand U29611 (N_29611,N_13399,N_13336);
xnor U29612 (N_29612,N_19208,N_10328);
or U29613 (N_29613,N_14018,N_16415);
nor U29614 (N_29614,N_10484,N_12002);
and U29615 (N_29615,N_15921,N_11918);
nor U29616 (N_29616,N_18999,N_11805);
nor U29617 (N_29617,N_14791,N_11450);
xnor U29618 (N_29618,N_10926,N_10787);
or U29619 (N_29619,N_16374,N_14379);
xor U29620 (N_29620,N_12690,N_16325);
nor U29621 (N_29621,N_14866,N_15569);
and U29622 (N_29622,N_14514,N_10464);
and U29623 (N_29623,N_14422,N_18964);
or U29624 (N_29624,N_14126,N_18166);
xnor U29625 (N_29625,N_10328,N_14372);
xnor U29626 (N_29626,N_12384,N_14022);
nor U29627 (N_29627,N_19108,N_11277);
or U29628 (N_29628,N_15030,N_10058);
nor U29629 (N_29629,N_17947,N_16353);
nor U29630 (N_29630,N_17521,N_13127);
nand U29631 (N_29631,N_19421,N_16648);
nand U29632 (N_29632,N_19775,N_15595);
and U29633 (N_29633,N_13653,N_15203);
and U29634 (N_29634,N_19812,N_12920);
or U29635 (N_29635,N_16023,N_16373);
or U29636 (N_29636,N_11422,N_15633);
or U29637 (N_29637,N_17710,N_14305);
nand U29638 (N_29638,N_18349,N_14060);
or U29639 (N_29639,N_10590,N_13807);
nor U29640 (N_29640,N_11095,N_11153);
nand U29641 (N_29641,N_14575,N_10045);
and U29642 (N_29642,N_10626,N_16665);
xor U29643 (N_29643,N_13976,N_17483);
and U29644 (N_29644,N_14294,N_14923);
and U29645 (N_29645,N_18578,N_10293);
nand U29646 (N_29646,N_19758,N_12851);
xnor U29647 (N_29647,N_17456,N_13026);
or U29648 (N_29648,N_11768,N_17058);
nor U29649 (N_29649,N_17346,N_19549);
or U29650 (N_29650,N_14080,N_16585);
nand U29651 (N_29651,N_13644,N_14294);
xor U29652 (N_29652,N_18705,N_11747);
nor U29653 (N_29653,N_15154,N_17011);
or U29654 (N_29654,N_12352,N_10452);
nand U29655 (N_29655,N_13532,N_10024);
and U29656 (N_29656,N_11182,N_17540);
and U29657 (N_29657,N_14958,N_17832);
nor U29658 (N_29658,N_12469,N_14073);
and U29659 (N_29659,N_14634,N_12022);
or U29660 (N_29660,N_11349,N_12947);
or U29661 (N_29661,N_17761,N_16377);
or U29662 (N_29662,N_19494,N_14948);
nand U29663 (N_29663,N_11732,N_19870);
or U29664 (N_29664,N_18411,N_11309);
and U29665 (N_29665,N_14294,N_15144);
and U29666 (N_29666,N_19570,N_19941);
and U29667 (N_29667,N_19544,N_15506);
nor U29668 (N_29668,N_18780,N_12862);
nand U29669 (N_29669,N_11519,N_11731);
nor U29670 (N_29670,N_15363,N_11648);
and U29671 (N_29671,N_15554,N_10294);
and U29672 (N_29672,N_14021,N_13597);
or U29673 (N_29673,N_15089,N_11588);
and U29674 (N_29674,N_17919,N_12073);
and U29675 (N_29675,N_14698,N_18491);
or U29676 (N_29676,N_18542,N_16358);
nor U29677 (N_29677,N_16567,N_17306);
nand U29678 (N_29678,N_14100,N_10827);
and U29679 (N_29679,N_19005,N_18791);
and U29680 (N_29680,N_10142,N_11974);
and U29681 (N_29681,N_11050,N_15325);
nand U29682 (N_29682,N_13702,N_13147);
nor U29683 (N_29683,N_12471,N_16943);
or U29684 (N_29684,N_10433,N_10345);
nor U29685 (N_29685,N_18268,N_14272);
nor U29686 (N_29686,N_10579,N_19236);
nor U29687 (N_29687,N_13327,N_15386);
nand U29688 (N_29688,N_17363,N_16153);
nand U29689 (N_29689,N_19766,N_12988);
nand U29690 (N_29690,N_11001,N_18299);
or U29691 (N_29691,N_19131,N_18183);
nand U29692 (N_29692,N_14177,N_10773);
nor U29693 (N_29693,N_12479,N_14781);
nor U29694 (N_29694,N_11763,N_17311);
nor U29695 (N_29695,N_12158,N_12935);
xor U29696 (N_29696,N_14940,N_11843);
nor U29697 (N_29697,N_11147,N_16341);
and U29698 (N_29698,N_19290,N_17451);
xnor U29699 (N_29699,N_11528,N_17854);
or U29700 (N_29700,N_17527,N_18832);
and U29701 (N_29701,N_10907,N_15640);
or U29702 (N_29702,N_16858,N_14621);
and U29703 (N_29703,N_10040,N_14764);
nand U29704 (N_29704,N_10785,N_15187);
nand U29705 (N_29705,N_16523,N_15058);
and U29706 (N_29706,N_10569,N_17518);
xor U29707 (N_29707,N_12513,N_16768);
nand U29708 (N_29708,N_18396,N_13191);
nor U29709 (N_29709,N_17383,N_16067);
and U29710 (N_29710,N_11628,N_11100);
and U29711 (N_29711,N_13342,N_15300);
and U29712 (N_29712,N_14187,N_17422);
nand U29713 (N_29713,N_11881,N_17857);
and U29714 (N_29714,N_16458,N_18584);
nor U29715 (N_29715,N_16009,N_11201);
or U29716 (N_29716,N_16495,N_17278);
nor U29717 (N_29717,N_13875,N_17127);
and U29718 (N_29718,N_10461,N_13327);
nand U29719 (N_29719,N_14012,N_17585);
or U29720 (N_29720,N_18432,N_16944);
xor U29721 (N_29721,N_12626,N_17311);
nand U29722 (N_29722,N_15577,N_13129);
xor U29723 (N_29723,N_10797,N_10743);
nand U29724 (N_29724,N_12776,N_13738);
nor U29725 (N_29725,N_11110,N_16048);
nor U29726 (N_29726,N_19653,N_14317);
or U29727 (N_29727,N_16940,N_12129);
and U29728 (N_29728,N_12948,N_13107);
nand U29729 (N_29729,N_18095,N_13457);
and U29730 (N_29730,N_16717,N_19740);
nand U29731 (N_29731,N_14894,N_10544);
and U29732 (N_29732,N_11471,N_19820);
nand U29733 (N_29733,N_17296,N_16394);
nor U29734 (N_29734,N_13226,N_14656);
nand U29735 (N_29735,N_19936,N_15402);
nor U29736 (N_29736,N_11671,N_16320);
nor U29737 (N_29737,N_10001,N_18559);
nand U29738 (N_29738,N_13028,N_15333);
xnor U29739 (N_29739,N_12618,N_11940);
nand U29740 (N_29740,N_12842,N_15324);
or U29741 (N_29741,N_18712,N_16330);
xor U29742 (N_29742,N_15997,N_11524);
or U29743 (N_29743,N_14888,N_13812);
nor U29744 (N_29744,N_13344,N_17934);
or U29745 (N_29745,N_12047,N_12732);
and U29746 (N_29746,N_12456,N_16719);
nor U29747 (N_29747,N_19333,N_14362);
or U29748 (N_29748,N_15100,N_11880);
or U29749 (N_29749,N_16863,N_17088);
nor U29750 (N_29750,N_10086,N_15672);
and U29751 (N_29751,N_11068,N_15399);
or U29752 (N_29752,N_18560,N_14211);
or U29753 (N_29753,N_16390,N_18621);
nor U29754 (N_29754,N_18976,N_15575);
nor U29755 (N_29755,N_17197,N_13414);
nor U29756 (N_29756,N_13007,N_12201);
nor U29757 (N_29757,N_15239,N_11639);
nand U29758 (N_29758,N_17064,N_18057);
nor U29759 (N_29759,N_16572,N_16075);
nor U29760 (N_29760,N_15715,N_18725);
nand U29761 (N_29761,N_11082,N_10692);
or U29762 (N_29762,N_15299,N_19759);
nand U29763 (N_29763,N_15061,N_11610);
or U29764 (N_29764,N_15291,N_17224);
or U29765 (N_29765,N_19683,N_18108);
nor U29766 (N_29766,N_11044,N_11066);
or U29767 (N_29767,N_12284,N_18833);
and U29768 (N_29768,N_17160,N_10371);
or U29769 (N_29769,N_15395,N_10258);
xor U29770 (N_29770,N_13269,N_12779);
and U29771 (N_29771,N_17368,N_14323);
xor U29772 (N_29772,N_13914,N_12531);
nand U29773 (N_29773,N_16438,N_17726);
nand U29774 (N_29774,N_16060,N_13654);
xor U29775 (N_29775,N_10126,N_15721);
or U29776 (N_29776,N_18729,N_16267);
and U29777 (N_29777,N_13027,N_18832);
or U29778 (N_29778,N_16339,N_19890);
nand U29779 (N_29779,N_18189,N_13541);
nor U29780 (N_29780,N_13719,N_17453);
xor U29781 (N_29781,N_18853,N_15836);
and U29782 (N_29782,N_11994,N_18183);
nand U29783 (N_29783,N_15667,N_14676);
nand U29784 (N_29784,N_18586,N_17330);
nor U29785 (N_29785,N_12565,N_13104);
and U29786 (N_29786,N_18075,N_10157);
and U29787 (N_29787,N_10716,N_17800);
or U29788 (N_29788,N_17488,N_17697);
nor U29789 (N_29789,N_17607,N_16182);
nand U29790 (N_29790,N_18983,N_16714);
nor U29791 (N_29791,N_14929,N_18790);
nand U29792 (N_29792,N_18865,N_11582);
nor U29793 (N_29793,N_17681,N_10216);
and U29794 (N_29794,N_13415,N_13897);
and U29795 (N_29795,N_13953,N_12126);
nand U29796 (N_29796,N_10642,N_14049);
and U29797 (N_29797,N_19405,N_14597);
nand U29798 (N_29798,N_15582,N_11923);
or U29799 (N_29799,N_13464,N_19287);
xnor U29800 (N_29800,N_19996,N_16058);
nand U29801 (N_29801,N_14155,N_19488);
nand U29802 (N_29802,N_16335,N_14025);
xor U29803 (N_29803,N_10902,N_19745);
nor U29804 (N_29804,N_10056,N_16299);
nand U29805 (N_29805,N_16772,N_18630);
and U29806 (N_29806,N_18015,N_19352);
nor U29807 (N_29807,N_10606,N_10170);
xnor U29808 (N_29808,N_15822,N_10223);
and U29809 (N_29809,N_19798,N_15004);
xor U29810 (N_29810,N_16050,N_15309);
xnor U29811 (N_29811,N_10157,N_11316);
or U29812 (N_29812,N_16499,N_18073);
nor U29813 (N_29813,N_12410,N_14489);
nand U29814 (N_29814,N_16815,N_18275);
nand U29815 (N_29815,N_15261,N_19604);
and U29816 (N_29816,N_10361,N_12277);
nor U29817 (N_29817,N_15609,N_12304);
and U29818 (N_29818,N_12544,N_14873);
nor U29819 (N_29819,N_15412,N_18148);
and U29820 (N_29820,N_19105,N_16804);
nand U29821 (N_29821,N_10564,N_11815);
and U29822 (N_29822,N_19999,N_10058);
nand U29823 (N_29823,N_14086,N_11894);
or U29824 (N_29824,N_17190,N_17718);
nand U29825 (N_29825,N_18621,N_11115);
or U29826 (N_29826,N_18251,N_13277);
xor U29827 (N_29827,N_19473,N_17949);
nor U29828 (N_29828,N_16696,N_12265);
or U29829 (N_29829,N_16898,N_19968);
and U29830 (N_29830,N_16212,N_17893);
nor U29831 (N_29831,N_12732,N_10335);
nand U29832 (N_29832,N_15881,N_16813);
or U29833 (N_29833,N_19348,N_11142);
nor U29834 (N_29834,N_19588,N_12878);
nand U29835 (N_29835,N_12307,N_15334);
and U29836 (N_29836,N_11705,N_15390);
or U29837 (N_29837,N_17755,N_13989);
nand U29838 (N_29838,N_14547,N_14072);
nand U29839 (N_29839,N_18111,N_11663);
and U29840 (N_29840,N_15336,N_14842);
and U29841 (N_29841,N_10322,N_19837);
nand U29842 (N_29842,N_18401,N_13483);
and U29843 (N_29843,N_11561,N_13019);
nor U29844 (N_29844,N_18416,N_15674);
and U29845 (N_29845,N_17392,N_13542);
or U29846 (N_29846,N_13384,N_10526);
and U29847 (N_29847,N_10400,N_19300);
and U29848 (N_29848,N_13981,N_16543);
xor U29849 (N_29849,N_12499,N_14569);
or U29850 (N_29850,N_16079,N_12794);
and U29851 (N_29851,N_10795,N_18880);
and U29852 (N_29852,N_11405,N_12957);
nor U29853 (N_29853,N_16072,N_15967);
nand U29854 (N_29854,N_14592,N_18998);
or U29855 (N_29855,N_11691,N_19888);
xor U29856 (N_29856,N_13849,N_14396);
nand U29857 (N_29857,N_18792,N_17780);
or U29858 (N_29858,N_17169,N_14191);
nor U29859 (N_29859,N_11065,N_14159);
nand U29860 (N_29860,N_11829,N_11713);
nand U29861 (N_29861,N_16874,N_14454);
or U29862 (N_29862,N_15210,N_18522);
or U29863 (N_29863,N_13613,N_18875);
and U29864 (N_29864,N_13403,N_14381);
and U29865 (N_29865,N_15154,N_14997);
or U29866 (N_29866,N_19914,N_11835);
nor U29867 (N_29867,N_15738,N_13922);
and U29868 (N_29868,N_13038,N_19961);
xnor U29869 (N_29869,N_13456,N_10691);
nor U29870 (N_29870,N_10891,N_11373);
xor U29871 (N_29871,N_10723,N_10513);
nand U29872 (N_29872,N_14674,N_12077);
or U29873 (N_29873,N_15508,N_10912);
nor U29874 (N_29874,N_10569,N_17972);
nor U29875 (N_29875,N_13710,N_10581);
nand U29876 (N_29876,N_12187,N_17132);
nand U29877 (N_29877,N_16619,N_17562);
and U29878 (N_29878,N_14816,N_12040);
or U29879 (N_29879,N_14224,N_11694);
nand U29880 (N_29880,N_10072,N_17693);
or U29881 (N_29881,N_11659,N_11904);
nand U29882 (N_29882,N_14426,N_12531);
nor U29883 (N_29883,N_19354,N_12162);
and U29884 (N_29884,N_18360,N_11080);
nand U29885 (N_29885,N_14039,N_19704);
xnor U29886 (N_29886,N_11115,N_16700);
and U29887 (N_29887,N_17896,N_12023);
nor U29888 (N_29888,N_13863,N_12825);
or U29889 (N_29889,N_19708,N_13541);
nand U29890 (N_29890,N_17716,N_10624);
and U29891 (N_29891,N_16254,N_17381);
and U29892 (N_29892,N_17375,N_15696);
or U29893 (N_29893,N_17850,N_10251);
nor U29894 (N_29894,N_15694,N_18635);
nand U29895 (N_29895,N_10588,N_14388);
nor U29896 (N_29896,N_18988,N_13623);
xor U29897 (N_29897,N_12090,N_18992);
xor U29898 (N_29898,N_15710,N_12478);
xnor U29899 (N_29899,N_15810,N_13256);
and U29900 (N_29900,N_13403,N_15297);
nand U29901 (N_29901,N_15521,N_16997);
and U29902 (N_29902,N_11019,N_13596);
or U29903 (N_29903,N_14439,N_14553);
and U29904 (N_29904,N_13710,N_16449);
and U29905 (N_29905,N_10288,N_18228);
and U29906 (N_29906,N_18679,N_16761);
or U29907 (N_29907,N_16089,N_10806);
or U29908 (N_29908,N_15783,N_15332);
nand U29909 (N_29909,N_15142,N_13538);
nor U29910 (N_29910,N_16931,N_18318);
nand U29911 (N_29911,N_19544,N_14913);
nor U29912 (N_29912,N_16382,N_19276);
nor U29913 (N_29913,N_14869,N_14899);
xnor U29914 (N_29914,N_10841,N_15581);
xnor U29915 (N_29915,N_16587,N_13931);
nand U29916 (N_29916,N_14529,N_14311);
or U29917 (N_29917,N_15547,N_15108);
or U29918 (N_29918,N_10017,N_13833);
nor U29919 (N_29919,N_18234,N_10209);
nor U29920 (N_29920,N_11226,N_18760);
xnor U29921 (N_29921,N_15425,N_14501);
nor U29922 (N_29922,N_11952,N_17302);
or U29923 (N_29923,N_17916,N_12351);
nand U29924 (N_29924,N_18544,N_16512);
nor U29925 (N_29925,N_18892,N_14247);
or U29926 (N_29926,N_18705,N_15981);
and U29927 (N_29927,N_19212,N_17819);
or U29928 (N_29928,N_14222,N_15770);
nand U29929 (N_29929,N_11939,N_17065);
and U29930 (N_29930,N_10388,N_15422);
xor U29931 (N_29931,N_15607,N_14715);
xor U29932 (N_29932,N_16649,N_15556);
nor U29933 (N_29933,N_17300,N_11587);
nor U29934 (N_29934,N_18135,N_16119);
nand U29935 (N_29935,N_10834,N_14047);
nor U29936 (N_29936,N_13815,N_12670);
and U29937 (N_29937,N_11373,N_13148);
or U29938 (N_29938,N_19605,N_10485);
and U29939 (N_29939,N_10298,N_11071);
and U29940 (N_29940,N_16039,N_14998);
nand U29941 (N_29941,N_16984,N_16545);
or U29942 (N_29942,N_14748,N_14503);
nand U29943 (N_29943,N_10342,N_11935);
and U29944 (N_29944,N_10885,N_10126);
xnor U29945 (N_29945,N_10265,N_12564);
or U29946 (N_29946,N_10953,N_17929);
nor U29947 (N_29947,N_13545,N_10054);
and U29948 (N_29948,N_12528,N_15540);
nor U29949 (N_29949,N_19704,N_12359);
and U29950 (N_29950,N_18039,N_15074);
nand U29951 (N_29951,N_17412,N_16993);
nor U29952 (N_29952,N_12779,N_14983);
and U29953 (N_29953,N_16638,N_15134);
nor U29954 (N_29954,N_12611,N_12622);
and U29955 (N_29955,N_11527,N_15832);
nand U29956 (N_29956,N_14882,N_14801);
nand U29957 (N_29957,N_19904,N_15768);
or U29958 (N_29958,N_10385,N_11439);
nor U29959 (N_29959,N_10717,N_10538);
nand U29960 (N_29960,N_17949,N_14287);
and U29961 (N_29961,N_15700,N_11827);
nor U29962 (N_29962,N_10381,N_10026);
nand U29963 (N_29963,N_17234,N_11134);
or U29964 (N_29964,N_11084,N_14923);
nand U29965 (N_29965,N_10269,N_13907);
nand U29966 (N_29966,N_11731,N_11849);
nor U29967 (N_29967,N_17839,N_17152);
nand U29968 (N_29968,N_14795,N_15599);
nor U29969 (N_29969,N_12413,N_10253);
and U29970 (N_29970,N_18757,N_19960);
and U29971 (N_29971,N_12065,N_14675);
and U29972 (N_29972,N_10163,N_18830);
nand U29973 (N_29973,N_16783,N_15009);
nand U29974 (N_29974,N_14004,N_10634);
and U29975 (N_29975,N_15629,N_19675);
and U29976 (N_29976,N_10074,N_19185);
nand U29977 (N_29977,N_17496,N_19579);
nand U29978 (N_29978,N_17974,N_15021);
or U29979 (N_29979,N_12821,N_15895);
nor U29980 (N_29980,N_12964,N_11095);
xnor U29981 (N_29981,N_14206,N_13928);
nor U29982 (N_29982,N_13084,N_10408);
or U29983 (N_29983,N_19452,N_13465);
nor U29984 (N_29984,N_19458,N_12425);
or U29985 (N_29985,N_17868,N_13119);
nor U29986 (N_29986,N_15370,N_18882);
or U29987 (N_29987,N_14845,N_16108);
and U29988 (N_29988,N_18623,N_19088);
nor U29989 (N_29989,N_11640,N_18883);
and U29990 (N_29990,N_16537,N_13359);
and U29991 (N_29991,N_19744,N_11081);
and U29992 (N_29992,N_12100,N_11907);
nand U29993 (N_29993,N_11117,N_19033);
and U29994 (N_29994,N_17999,N_17409);
and U29995 (N_29995,N_14036,N_13151);
xor U29996 (N_29996,N_16107,N_15826);
nand U29997 (N_29997,N_17031,N_15050);
nor U29998 (N_29998,N_13612,N_11383);
nor U29999 (N_29999,N_19128,N_17963);
nand U30000 (N_30000,N_22033,N_20858);
or U30001 (N_30001,N_22132,N_22782);
or U30002 (N_30002,N_24365,N_23993);
or U30003 (N_30003,N_27088,N_26749);
or U30004 (N_30004,N_29511,N_21039);
xor U30005 (N_30005,N_25325,N_20140);
nand U30006 (N_30006,N_26733,N_20658);
nand U30007 (N_30007,N_23495,N_22669);
nand U30008 (N_30008,N_27866,N_28407);
nand U30009 (N_30009,N_21441,N_21467);
and U30010 (N_30010,N_21384,N_28097);
or U30011 (N_30011,N_25808,N_25644);
and U30012 (N_30012,N_23003,N_20973);
or U30013 (N_30013,N_26321,N_24510);
xnor U30014 (N_30014,N_28439,N_21472);
and U30015 (N_30015,N_25460,N_25503);
nor U30016 (N_30016,N_27851,N_22888);
and U30017 (N_30017,N_25729,N_21959);
nand U30018 (N_30018,N_24835,N_21923);
nor U30019 (N_30019,N_22849,N_22030);
nand U30020 (N_30020,N_29115,N_28771);
xnor U30021 (N_30021,N_26647,N_23490);
nor U30022 (N_30022,N_29648,N_21122);
nor U30023 (N_30023,N_22490,N_28377);
nor U30024 (N_30024,N_21527,N_20726);
xnor U30025 (N_30025,N_22929,N_28085);
or U30026 (N_30026,N_27638,N_21437);
and U30027 (N_30027,N_22122,N_29484);
or U30028 (N_30028,N_23920,N_23481);
and U30029 (N_30029,N_25650,N_29688);
nor U30030 (N_30030,N_26718,N_24973);
or U30031 (N_30031,N_29033,N_27634);
nand U30032 (N_30032,N_24666,N_21982);
or U30033 (N_30033,N_27691,N_22433);
and U30034 (N_30034,N_24946,N_20917);
or U30035 (N_30035,N_29908,N_29582);
or U30036 (N_30036,N_27723,N_28864);
nor U30037 (N_30037,N_26947,N_26966);
or U30038 (N_30038,N_22439,N_23008);
nor U30039 (N_30039,N_26461,N_20539);
or U30040 (N_30040,N_27533,N_25712);
xnor U30041 (N_30041,N_21872,N_26286);
or U30042 (N_30042,N_29683,N_23581);
nor U30043 (N_30043,N_20297,N_21880);
nor U30044 (N_30044,N_20408,N_20629);
nand U30045 (N_30045,N_23916,N_27079);
or U30046 (N_30046,N_22947,N_21623);
nor U30047 (N_30047,N_26005,N_20284);
or U30048 (N_30048,N_23099,N_29021);
or U30049 (N_30049,N_24026,N_23299);
nor U30050 (N_30050,N_22593,N_21821);
and U30051 (N_30051,N_24176,N_23111);
and U30052 (N_30052,N_21108,N_22142);
or U30053 (N_30053,N_26208,N_25666);
nor U30054 (N_30054,N_21973,N_29491);
or U30055 (N_30055,N_23087,N_29264);
nor U30056 (N_30056,N_23990,N_22316);
and U30057 (N_30057,N_24538,N_24439);
nor U30058 (N_30058,N_21838,N_27952);
and U30059 (N_30059,N_24185,N_23749);
and U30060 (N_30060,N_25851,N_24484);
and U30061 (N_30061,N_20871,N_20526);
xnor U30062 (N_30062,N_29451,N_25701);
and U30063 (N_30063,N_27190,N_28489);
and U30064 (N_30064,N_29707,N_22774);
nand U30065 (N_30065,N_28357,N_29913);
nor U30066 (N_30066,N_28106,N_29882);
nor U30067 (N_30067,N_29637,N_24713);
and U30068 (N_30068,N_25233,N_20243);
nor U30069 (N_30069,N_23665,N_24002);
xnor U30070 (N_30070,N_27432,N_22060);
nor U30071 (N_30071,N_22743,N_21805);
and U30072 (N_30072,N_21845,N_27782);
nor U30073 (N_30073,N_29110,N_22044);
nand U30074 (N_30074,N_28276,N_25497);
or U30075 (N_30075,N_22797,N_26405);
nor U30076 (N_30076,N_29804,N_25065);
or U30077 (N_30077,N_23283,N_26398);
or U30078 (N_30078,N_26883,N_28075);
nor U30079 (N_30079,N_23694,N_20427);
nand U30080 (N_30080,N_25525,N_27383);
or U30081 (N_30081,N_26373,N_26061);
nor U30082 (N_30082,N_22816,N_20435);
or U30083 (N_30083,N_24663,N_29011);
nand U30084 (N_30084,N_24469,N_21575);
nor U30085 (N_30085,N_26701,N_24989);
or U30086 (N_30086,N_22135,N_24281);
nor U30087 (N_30087,N_29124,N_23122);
nor U30088 (N_30088,N_20781,N_24130);
nor U30089 (N_30089,N_27564,N_25394);
nand U30090 (N_30090,N_25379,N_21248);
and U30091 (N_30091,N_22498,N_27548);
nor U30092 (N_30092,N_21731,N_21702);
and U30093 (N_30093,N_20759,N_20684);
xor U30094 (N_30094,N_27076,N_20316);
nor U30095 (N_30095,N_28229,N_22120);
nor U30096 (N_30096,N_26618,N_23478);
nand U30097 (N_30097,N_25002,N_27673);
nor U30098 (N_30098,N_21770,N_29029);
nand U30099 (N_30099,N_22228,N_25723);
or U30100 (N_30100,N_23801,N_25377);
and U30101 (N_30101,N_26785,N_26201);
or U30102 (N_30102,N_24191,N_26519);
or U30103 (N_30103,N_28495,N_29714);
and U30104 (N_30104,N_28277,N_25541);
or U30105 (N_30105,N_23459,N_26536);
nor U30106 (N_30106,N_24341,N_21092);
and U30107 (N_30107,N_29500,N_23373);
nand U30108 (N_30108,N_20402,N_29221);
nor U30109 (N_30109,N_21135,N_25324);
nor U30110 (N_30110,N_25090,N_25979);
nand U30111 (N_30111,N_21809,N_20456);
nand U30112 (N_30112,N_23187,N_29784);
and U30113 (N_30113,N_29171,N_27276);
and U30114 (N_30114,N_27238,N_25019);
nor U30115 (N_30115,N_21190,N_21130);
nor U30116 (N_30116,N_21921,N_23966);
nor U30117 (N_30117,N_22821,N_23304);
and U30118 (N_30118,N_20974,N_28023);
or U30119 (N_30119,N_24244,N_27012);
nor U30120 (N_30120,N_23416,N_24422);
and U30121 (N_30121,N_29699,N_28126);
and U30122 (N_30122,N_27081,N_24159);
and U30123 (N_30123,N_25321,N_21667);
and U30124 (N_30124,N_24058,N_28271);
nor U30125 (N_30125,N_20665,N_28831);
and U30126 (N_30126,N_29860,N_29969);
nor U30127 (N_30127,N_29348,N_27797);
or U30128 (N_30128,N_27311,N_20621);
nand U30129 (N_30129,N_20116,N_26620);
or U30130 (N_30130,N_25473,N_21440);
or U30131 (N_30131,N_26724,N_21278);
xor U30132 (N_30132,N_27570,N_26251);
nor U30133 (N_30133,N_21019,N_29539);
or U30134 (N_30134,N_23190,N_24459);
or U30135 (N_30135,N_20851,N_29712);
nand U30136 (N_30136,N_27559,N_20880);
or U30137 (N_30137,N_22602,N_25048);
xor U30138 (N_30138,N_20487,N_26206);
xnor U30139 (N_30139,N_24918,N_23599);
or U30140 (N_30140,N_26556,N_25353);
or U30141 (N_30141,N_22104,N_21879);
nor U30142 (N_30142,N_25208,N_25357);
nand U30143 (N_30143,N_26220,N_26554);
and U30144 (N_30144,N_27579,N_27931);
and U30145 (N_30145,N_28070,N_23663);
and U30146 (N_30146,N_26154,N_29287);
or U30147 (N_30147,N_24719,N_23396);
xor U30148 (N_30148,N_23433,N_22221);
xor U30149 (N_30149,N_25501,N_21744);
nor U30150 (N_30150,N_21313,N_20843);
and U30151 (N_30151,N_20511,N_24115);
xor U30152 (N_30152,N_29122,N_29662);
or U30153 (N_30153,N_20475,N_25249);
nand U30154 (N_30154,N_21300,N_26514);
nand U30155 (N_30155,N_22628,N_22497);
nor U30156 (N_30156,N_29106,N_22327);
or U30157 (N_30157,N_23005,N_20497);
and U30158 (N_30158,N_20139,N_20033);
nor U30159 (N_30159,N_27343,N_25575);
xor U30160 (N_30160,N_25934,N_22858);
or U30161 (N_30161,N_22031,N_27742);
nor U30162 (N_30162,N_23561,N_25752);
nand U30163 (N_30163,N_21392,N_20868);
and U30164 (N_30164,N_28122,N_29663);
nor U30165 (N_30165,N_21670,N_25197);
or U30166 (N_30166,N_23704,N_23114);
and U30167 (N_30167,N_22538,N_26122);
and U30168 (N_30168,N_21065,N_21624);
or U30169 (N_30169,N_20407,N_27889);
and U30170 (N_30170,N_22253,N_21598);
nand U30171 (N_30171,N_29706,N_20030);
nand U30172 (N_30172,N_26503,N_23148);
nand U30173 (N_30173,N_22304,N_24850);
nor U30174 (N_30174,N_24517,N_22420);
and U30175 (N_30175,N_23783,N_25075);
and U30176 (N_30176,N_28713,N_23204);
nand U30177 (N_30177,N_23149,N_29709);
or U30178 (N_30178,N_24304,N_22807);
nand U30179 (N_30179,N_25602,N_25969);
or U30180 (N_30180,N_24386,N_22360);
or U30181 (N_30181,N_23234,N_22454);
xor U30182 (N_30182,N_27899,N_20058);
and U30183 (N_30183,N_29204,N_24692);
or U30184 (N_30184,N_25856,N_24683);
and U30185 (N_30185,N_21884,N_21329);
and U30186 (N_30186,N_21727,N_26330);
xnor U30187 (N_30187,N_28565,N_22097);
nand U30188 (N_30188,N_22921,N_21853);
xnor U30189 (N_30189,N_27593,N_25632);
nand U30190 (N_30190,N_24527,N_28644);
xor U30191 (N_30191,N_28472,N_28453);
nor U30192 (N_30192,N_21317,N_20300);
nand U30193 (N_30193,N_21170,N_26680);
and U30194 (N_30194,N_27733,N_28561);
and U30195 (N_30195,N_24198,N_27926);
nand U30196 (N_30196,N_25058,N_26541);
and U30197 (N_30197,N_24774,N_27323);
and U30198 (N_30198,N_22941,N_26234);
xor U30199 (N_30199,N_20281,N_29226);
and U30200 (N_30200,N_27933,N_21179);
or U30201 (N_30201,N_22185,N_20031);
or U30202 (N_30202,N_26786,N_27769);
nand U30203 (N_30203,N_22173,N_28185);
and U30204 (N_30204,N_27685,N_29392);
nand U30205 (N_30205,N_29595,N_21126);
nand U30206 (N_30206,N_29280,N_22007);
nand U30207 (N_30207,N_28485,N_26432);
nor U30208 (N_30208,N_24875,N_24845);
and U30209 (N_30209,N_26690,N_22488);
xnor U30210 (N_30210,N_28571,N_21298);
and U30211 (N_30211,N_25868,N_29194);
or U30212 (N_30212,N_28873,N_27761);
nor U30213 (N_30213,N_27770,N_20661);
nand U30214 (N_30214,N_26027,N_25192);
xor U30215 (N_30215,N_25014,N_25757);
nand U30216 (N_30216,N_29135,N_22883);
or U30217 (N_30217,N_24591,N_28088);
and U30218 (N_30218,N_24912,N_22512);
and U30219 (N_30219,N_29812,N_25830);
and U30220 (N_30220,N_24633,N_27752);
nand U30221 (N_30221,N_23430,N_20592);
nor U30222 (N_30222,N_20500,N_28691);
nand U30223 (N_30223,N_23246,N_20131);
nand U30224 (N_30224,N_25457,N_27523);
or U30225 (N_30225,N_20046,N_26813);
nand U30226 (N_30226,N_29968,N_29018);
and U30227 (N_30227,N_21209,N_27253);
and U30228 (N_30228,N_23411,N_22051);
and U30229 (N_30229,N_20888,N_23914);
and U30230 (N_30230,N_28090,N_28076);
nor U30231 (N_30231,N_22974,N_23588);
xnor U30232 (N_30232,N_24747,N_22103);
or U30233 (N_30233,N_29019,N_23476);
nor U30234 (N_30234,N_20869,N_25446);
nor U30235 (N_30235,N_25173,N_22091);
nor U30236 (N_30236,N_26305,N_23985);
or U30237 (N_30237,N_23102,N_29156);
xnor U30238 (N_30238,N_22499,N_23155);
and U30239 (N_30239,N_25433,N_29726);
or U30240 (N_30240,N_22267,N_24024);
nor U30241 (N_30241,N_23844,N_25623);
or U30242 (N_30242,N_25329,N_25283);
nand U30243 (N_30243,N_22540,N_22922);
nand U30244 (N_30244,N_23516,N_20146);
nor U30245 (N_30245,N_28342,N_26320);
and U30246 (N_30246,N_21568,N_21421);
and U30247 (N_30247,N_21798,N_27743);
nand U30248 (N_30248,N_28012,N_23718);
or U30249 (N_30249,N_20036,N_20115);
or U30250 (N_30250,N_25733,N_21952);
and U30251 (N_30251,N_28436,N_27610);
xor U30252 (N_30252,N_27053,N_21611);
and U30253 (N_30253,N_25322,N_21000);
nand U30254 (N_30254,N_27505,N_21625);
nor U30255 (N_30255,N_20686,N_26625);
or U30256 (N_30256,N_20999,N_24947);
nor U30257 (N_30257,N_29079,N_20688);
nand U30258 (N_30258,N_27994,N_20735);
nand U30259 (N_30259,N_27671,N_20787);
nor U30260 (N_30260,N_20133,N_24980);
or U30261 (N_30261,N_25782,N_25056);
nor U30262 (N_30262,N_23793,N_20950);
or U30263 (N_30263,N_26545,N_21752);
nand U30264 (N_30264,N_24150,N_20225);
nor U30265 (N_30265,N_24920,N_23260);
and U30266 (N_30266,N_25144,N_26230);
and U30267 (N_30267,N_25680,N_28886);
and U30268 (N_30268,N_27167,N_23787);
xnor U30269 (N_30269,N_28518,N_25371);
nand U30270 (N_30270,N_28036,N_24300);
nand U30271 (N_30271,N_25892,N_21022);
and U30272 (N_30272,N_23037,N_25532);
or U30273 (N_30273,N_27915,N_29049);
or U30274 (N_30274,N_29689,N_27474);
or U30275 (N_30275,N_29176,N_20605);
nor U30276 (N_30276,N_20675,N_21653);
xor U30277 (N_30277,N_28467,N_23021);
or U30278 (N_30278,N_29530,N_23058);
and U30279 (N_30279,N_25311,N_24294);
or U30280 (N_30280,N_23466,N_20863);
or U30281 (N_30281,N_26147,N_24228);
nand U30282 (N_30282,N_26851,N_27821);
nand U30283 (N_30283,N_23737,N_23059);
or U30284 (N_30284,N_21438,N_28511);
nor U30285 (N_30285,N_20985,N_27052);
xnor U30286 (N_30286,N_25376,N_22409);
nor U30287 (N_30287,N_25147,N_22308);
or U30288 (N_30288,N_22002,N_24631);
or U30289 (N_30289,N_26210,N_25124);
and U30290 (N_30290,N_27524,N_23168);
and U30291 (N_30291,N_23189,N_27541);
and U30292 (N_30292,N_29549,N_24498);
or U30293 (N_30293,N_23865,N_26946);
or U30294 (N_30294,N_23975,N_20259);
nand U30295 (N_30295,N_23429,N_24627);
nor U30296 (N_30296,N_22994,N_28067);
nand U30297 (N_30297,N_29416,N_26306);
nor U30298 (N_30298,N_22978,N_25230);
nand U30299 (N_30299,N_27278,N_23469);
or U30300 (N_30300,N_27200,N_28093);
xor U30301 (N_30301,N_24212,N_22694);
or U30302 (N_30302,N_28029,N_23837);
nor U30303 (N_30303,N_24158,N_21825);
nor U30304 (N_30304,N_28005,N_28159);
nand U30305 (N_30305,N_28345,N_29134);
and U30306 (N_30306,N_22618,N_22930);
nand U30307 (N_30307,N_21127,N_29561);
xnor U30308 (N_30308,N_26716,N_24789);
nor U30309 (N_30309,N_27577,N_23949);
nor U30310 (N_30310,N_23514,N_28618);
and U30311 (N_30311,N_25698,N_28323);
nand U30312 (N_30312,N_22814,N_28336);
nor U30313 (N_30313,N_24908,N_22070);
and U30314 (N_30314,N_20531,N_23223);
nand U30315 (N_30315,N_28679,N_21009);
and U30316 (N_30316,N_21276,N_21328);
or U30317 (N_30317,N_29618,N_25565);
and U30318 (N_30318,N_23981,N_25450);
nand U30319 (N_30319,N_23047,N_24731);
nor U30320 (N_30320,N_21174,N_23662);
xor U30321 (N_30321,N_29685,N_25605);
and U30322 (N_30322,N_20378,N_20965);
nor U30323 (N_30323,N_27969,N_22845);
nor U30324 (N_30324,N_22015,N_21206);
nand U30325 (N_30325,N_25801,N_23198);
nand U30326 (N_30326,N_23841,N_24334);
nor U30327 (N_30327,N_22478,N_21269);
nor U30328 (N_30328,N_24271,N_29395);
nor U30329 (N_30329,N_23517,N_21931);
nor U30330 (N_30330,N_29380,N_23670);
xor U30331 (N_30331,N_27690,N_23642);
nor U30332 (N_30332,N_22961,N_22714);
and U30333 (N_30333,N_23144,N_23651);
nand U30334 (N_30334,N_28955,N_26173);
or U30335 (N_30335,N_21609,N_26617);
nor U30336 (N_30336,N_22565,N_26875);
or U30337 (N_30337,N_24240,N_23504);
nand U30338 (N_30338,N_29369,N_26916);
nor U30339 (N_30339,N_21338,N_20295);
nor U30340 (N_30340,N_20020,N_25703);
nor U30341 (N_30341,N_20749,N_26792);
xor U30342 (N_30342,N_26940,N_24133);
nand U30343 (N_30343,N_26582,N_27701);
nor U30344 (N_30344,N_25118,N_25063);
and U30345 (N_30345,N_21337,N_22806);
and U30346 (N_30346,N_26521,N_21492);
nand U30347 (N_30347,N_20625,N_26138);
or U30348 (N_30348,N_28598,N_24406);
nand U30349 (N_30349,N_23986,N_25076);
xnor U30350 (N_30350,N_22434,N_27407);
nor U30351 (N_30351,N_22213,N_26354);
or U30352 (N_30352,N_25242,N_23751);
nor U30353 (N_30353,N_27737,N_26042);
and U30354 (N_30354,N_26463,N_20745);
or U30355 (N_30355,N_26911,N_22134);
and U30356 (N_30356,N_21383,N_29281);
nand U30357 (N_30357,N_29386,N_20877);
and U30358 (N_30358,N_23220,N_29796);
and U30359 (N_30359,N_25248,N_21998);
and U30360 (N_30360,N_27083,N_24356);
or U30361 (N_30361,N_27639,N_21267);
nor U30362 (N_30362,N_28230,N_23525);
nand U30363 (N_30363,N_20632,N_22966);
or U30364 (N_30364,N_20035,N_23281);
or U30365 (N_30365,N_28554,N_27852);
nand U30366 (N_30366,N_25445,N_27504);
nor U30367 (N_30367,N_27038,N_24557);
and U30368 (N_30368,N_23842,N_25171);
nand U30369 (N_30369,N_27153,N_27551);
and U30370 (N_30370,N_26585,N_23073);
or U30371 (N_30371,N_22178,N_29232);
nor U30372 (N_30372,N_23507,N_27672);
and U30373 (N_30373,N_26259,N_21914);
xnor U30374 (N_30374,N_25668,N_22069);
and U30375 (N_30375,N_28652,N_23460);
nor U30376 (N_30376,N_25217,N_28290);
nand U30377 (N_30377,N_21684,N_26957);
nor U30378 (N_30378,N_23773,N_21435);
nor U30379 (N_30379,N_21698,N_21720);
or U30380 (N_30380,N_28900,N_27886);
or U30381 (N_30381,N_21377,N_29446);
and U30382 (N_30382,N_29360,N_28242);
nor U30383 (N_30383,N_23544,N_24087);
nor U30384 (N_30384,N_29301,N_20064);
xor U30385 (N_30385,N_24938,N_28057);
nor U30386 (N_30386,N_21528,N_26632);
xnor U30387 (N_30387,N_26179,N_27808);
nor U30388 (N_30388,N_27684,N_24025);
xor U30389 (N_30389,N_26668,N_22662);
nor U30390 (N_30390,N_28113,N_21478);
and U30391 (N_30391,N_22681,N_29946);
nor U30392 (N_30392,N_24607,N_25026);
and U30393 (N_30393,N_22296,N_26692);
nor U30394 (N_30394,N_21846,N_20060);
or U30395 (N_30395,N_23337,N_29872);
or U30396 (N_30396,N_25461,N_29282);
and U30397 (N_30397,N_21169,N_21415);
nor U30398 (N_30398,N_26930,N_25443);
or U30399 (N_30399,N_24923,N_24592);
and U30400 (N_30400,N_20341,N_27956);
nor U30401 (N_30401,N_21318,N_28260);
and U30402 (N_30402,N_24044,N_23484);
xnor U30403 (N_30403,N_27357,N_20450);
nor U30404 (N_30404,N_20163,N_28809);
nor U30405 (N_30405,N_23943,N_25347);
and U30406 (N_30406,N_23730,N_27015);
or U30407 (N_30407,N_24497,N_24114);
xnor U30408 (N_30408,N_21036,N_24028);
and U30409 (N_30409,N_20900,N_26999);
and U30410 (N_30410,N_20233,N_28974);
and U30411 (N_30411,N_29246,N_20845);
nand U30412 (N_30412,N_28199,N_20522);
and U30413 (N_30413,N_27439,N_26638);
and U30414 (N_30414,N_20956,N_24284);
or U30415 (N_30415,N_24526,N_28209);
nor U30416 (N_30416,N_23926,N_25990);
nor U30417 (N_30417,N_20200,N_28137);
and U30418 (N_30418,N_22812,N_26741);
nor U30419 (N_30419,N_24362,N_26948);
and U30420 (N_30420,N_28545,N_28662);
xnor U30421 (N_30421,N_21149,N_21602);
and U30422 (N_30422,N_25114,N_27929);
or U30423 (N_30423,N_20441,N_26708);
and U30424 (N_30424,N_20876,N_27301);
nand U30425 (N_30425,N_26133,N_25308);
nor U30426 (N_30426,N_22429,N_26057);
nor U30427 (N_30427,N_26856,N_28218);
xnor U30428 (N_30428,N_28066,N_22016);
and U30429 (N_30429,N_20345,N_22995);
nor U30430 (N_30430,N_28812,N_29117);
or U30431 (N_30431,N_23859,N_20360);
or U30432 (N_30432,N_26293,N_24858);
xnor U30433 (N_30433,N_20028,N_21807);
nand U30434 (N_30434,N_22037,N_21689);
and U30435 (N_30435,N_28615,N_23358);
and U30436 (N_30436,N_27068,N_28469);
nand U30437 (N_30437,N_22475,N_26177);
nand U30438 (N_30438,N_26796,N_28578);
xor U30439 (N_30439,N_21388,N_21719);
nor U30440 (N_30440,N_20042,N_24937);
and U30441 (N_30441,N_20377,N_22281);
nand U30442 (N_30442,N_23634,N_27689);
nor U30443 (N_30443,N_29774,N_23454);
or U30444 (N_30444,N_20488,N_28604);
and U30445 (N_30445,N_24675,N_20125);
nand U30446 (N_30446,N_20611,N_28896);
nor U30447 (N_30447,N_24934,N_29202);
or U30448 (N_30448,N_25995,N_25642);
or U30449 (N_30449,N_23638,N_21399);
nand U30450 (N_30450,N_29701,N_21412);
or U30451 (N_30451,N_25012,N_25126);
or U30452 (N_30452,N_23597,N_24475);
or U30453 (N_30453,N_26236,N_26593);
or U30454 (N_30454,N_20918,N_28632);
nand U30455 (N_30455,N_29223,N_23848);
nand U30456 (N_30456,N_21980,N_27388);
or U30457 (N_30457,N_22098,N_28350);
or U30458 (N_30458,N_28333,N_25653);
nor U30459 (N_30459,N_27268,N_29564);
and U30460 (N_30460,N_20422,N_22321);
or U30461 (N_30461,N_23060,N_28026);
and U30462 (N_30462,N_29729,N_26216);
nor U30463 (N_30463,N_25032,N_29108);
or U30464 (N_30464,N_21722,N_27507);
and U30465 (N_30465,N_28614,N_25290);
and U30466 (N_30466,N_20874,N_27798);
or U30467 (N_30467,N_21852,N_20706);
or U30468 (N_30468,N_28019,N_22043);
xnor U30469 (N_30469,N_29922,N_20148);
and U30470 (N_30470,N_21355,N_21911);
nor U30471 (N_30471,N_29728,N_20136);
nand U30472 (N_30472,N_29455,N_20144);
xor U30473 (N_30473,N_25767,N_25133);
nor U30474 (N_30474,N_28686,N_25552);
nor U30475 (N_30475,N_27807,N_26377);
or U30476 (N_30476,N_23885,N_20338);
nand U30477 (N_30477,N_24690,N_20461);
nor U30478 (N_30478,N_22052,N_24561);
or U30479 (N_30479,N_23320,N_23790);
nand U30480 (N_30480,N_28786,N_22075);
and U30481 (N_30481,N_27018,N_25388);
nand U30482 (N_30482,N_28160,N_29353);
and U30483 (N_30483,N_21981,N_22309);
or U30484 (N_30484,N_20301,N_27718);
nand U30485 (N_30485,N_29507,N_24518);
or U30486 (N_30486,N_25987,N_27874);
and U30487 (N_30487,N_20196,N_21005);
nor U30488 (N_30488,N_27376,N_22742);
or U30489 (N_30489,N_23064,N_24337);
nand U30490 (N_30490,N_27172,N_26355);
xnor U30491 (N_30491,N_22829,N_24846);
nand U30492 (N_30492,N_28825,N_24739);
xnor U30493 (N_30493,N_29616,N_22735);
xor U30494 (N_30494,N_20052,N_20510);
xor U30495 (N_30495,N_28658,N_23566);
or U30496 (N_30496,N_24291,N_22148);
or U30497 (N_30497,N_21491,N_28585);
and U30498 (N_30498,N_21735,N_27982);
and U30499 (N_30499,N_21090,N_24219);
and U30500 (N_30500,N_26637,N_21908);
or U30501 (N_30501,N_29790,N_27308);
nor U30502 (N_30502,N_27193,N_25909);
and U30503 (N_30503,N_24791,N_22278);
xnor U30504 (N_30504,N_20633,N_26097);
xor U30505 (N_30505,N_24837,N_23854);
nand U30506 (N_30506,N_28528,N_22456);
nor U30507 (N_30507,N_21746,N_21094);
and U30508 (N_30508,N_20697,N_23184);
nor U30509 (N_30509,N_26642,N_29420);
or U30510 (N_30510,N_25905,N_25508);
nor U30511 (N_30511,N_21817,N_20969);
and U30512 (N_30512,N_29635,N_20289);
and U30513 (N_30513,N_25458,N_25366);
xor U30514 (N_30514,N_29001,N_23777);
or U30515 (N_30515,N_29004,N_26979);
and U30516 (N_30516,N_25559,N_22196);
and U30517 (N_30517,N_28071,N_29944);
or U30518 (N_30518,N_28870,N_21538);
or U30519 (N_30519,N_29863,N_21458);
nor U30520 (N_30520,N_28884,N_21968);
or U30521 (N_30521,N_23456,N_23887);
or U30522 (N_30522,N_24221,N_26890);
nand U30523 (N_30523,N_21232,N_29240);
and U30524 (N_30524,N_22979,N_20241);
or U30525 (N_30525,N_29972,N_23824);
nand U30526 (N_30526,N_20175,N_22305);
nor U30527 (N_30527,N_23622,N_23094);
nand U30528 (N_30528,N_22057,N_23397);
nand U30529 (N_30529,N_26719,N_29158);
nand U30530 (N_30530,N_20979,N_25500);
nand U30531 (N_30531,N_22382,N_23860);
nand U30532 (N_30532,N_22237,N_25005);
nor U30533 (N_30533,N_26287,N_29390);
nor U30534 (N_30534,N_29572,N_27983);
or U30535 (N_30535,N_21042,N_20966);
nor U30536 (N_30536,N_25589,N_21289);
nand U30537 (N_30537,N_26886,N_24905);
nand U30538 (N_30538,N_29184,N_20504);
nand U30539 (N_30539,N_22559,N_23011);
and U30540 (N_30540,N_28581,N_26760);
and U30541 (N_30541,N_21603,N_20569);
nor U30542 (N_30542,N_23221,N_29649);
xor U30543 (N_30543,N_20654,N_25378);
or U30544 (N_30544,N_29192,N_28452);
nor U30545 (N_30545,N_23479,N_20127);
nand U30546 (N_30546,N_24400,N_24828);
or U30547 (N_30547,N_27865,N_28972);
and U30548 (N_30548,N_24571,N_29235);
nor U30549 (N_30549,N_21109,N_24339);
or U30550 (N_30550,N_25510,N_27848);
or U30551 (N_30551,N_29418,N_27884);
nand U30552 (N_30552,N_28858,N_25434);
nor U30553 (N_30553,N_28438,N_21453);
or U30554 (N_30554,N_27061,N_21301);
nor U30555 (N_30555,N_20564,N_26568);
or U30556 (N_30556,N_27783,N_25906);
or U30557 (N_30557,N_28282,N_26508);
xor U30558 (N_30558,N_22383,N_23224);
and U30559 (N_30559,N_28646,N_23624);
nand U30560 (N_30560,N_29073,N_20315);
nor U30561 (N_30561,N_22218,N_23667);
or U30562 (N_30562,N_23427,N_29198);
or U30563 (N_30563,N_21940,N_21083);
and U30564 (N_30564,N_22398,N_23354);
nor U30565 (N_30565,N_22254,N_20914);
or U30566 (N_30566,N_25582,N_27666);
nor U30567 (N_30567,N_20169,N_27904);
and U30568 (N_30568,N_29414,N_28714);
and U30569 (N_30569,N_26022,N_22076);
and U30570 (N_30570,N_22526,N_28053);
and U30571 (N_30571,N_29771,N_28153);
and U30572 (N_30572,N_26976,N_28400);
or U30573 (N_30573,N_27342,N_28551);
nor U30574 (N_30574,N_24384,N_28688);
and U30575 (N_30575,N_26766,N_23513);
nor U30576 (N_30576,N_24906,N_22917);
and U30577 (N_30577,N_29768,N_20172);
or U30578 (N_30578,N_24354,N_29075);
xnor U30579 (N_30579,N_28621,N_20587);
nand U30580 (N_30580,N_29288,N_24105);
nor U30581 (N_30581,N_27799,N_21664);
xor U30582 (N_30582,N_28981,N_20687);
nand U30583 (N_30583,N_20394,N_23276);
nand U30584 (N_30584,N_20774,N_23652);
nor U30585 (N_30585,N_20419,N_22337);
and U30586 (N_30586,N_28429,N_28587);
or U30587 (N_30587,N_24245,N_24137);
nor U30588 (N_30588,N_24042,N_20643);
nor U30589 (N_30589,N_27173,N_27912);
nand U30590 (N_30590,N_24143,N_28569);
nand U30591 (N_30591,N_25982,N_25512);
or U30592 (N_30592,N_24216,N_24095);
or U30593 (N_30593,N_22598,N_24573);
nor U30594 (N_30594,N_20810,N_25989);
xnor U30595 (N_30595,N_22533,N_26590);
or U30596 (N_30596,N_22422,N_23036);
and U30597 (N_30597,N_24964,N_26839);
and U30598 (N_30598,N_20051,N_23802);
nand U30599 (N_30599,N_27314,N_28902);
or U30600 (N_30600,N_23820,N_20232);
nand U30601 (N_30601,N_23425,N_23017);
and U30602 (N_30602,N_21525,N_22046);
nor U30603 (N_30603,N_29673,N_28146);
nor U30604 (N_30604,N_21520,N_23421);
nand U30605 (N_30605,N_27377,N_23760);
nor U30606 (N_30606,N_22428,N_20722);
or U30607 (N_30607,N_26880,N_20124);
nand U30608 (N_30608,N_22323,N_20262);
and U30609 (N_30609,N_23488,N_29323);
and U30610 (N_30610,N_25626,N_23308);
and U30611 (N_30611,N_28953,N_29779);
and U30612 (N_30612,N_28501,N_27037);
nand U30613 (N_30613,N_20350,N_20549);
nor U30614 (N_30614,N_23267,N_27247);
and U30615 (N_30615,N_20111,N_29208);
nor U30616 (N_30616,N_29026,N_20708);
nand U30617 (N_30617,N_28856,N_24998);
xnor U30618 (N_30618,N_26700,N_27463);
nor U30619 (N_30619,N_25097,N_23141);
nor U30620 (N_30620,N_28839,N_22352);
nor U30621 (N_30621,N_23810,N_26973);
nand U30622 (N_30622,N_20393,N_29841);
or U30623 (N_30623,N_28092,N_21284);
and U30624 (N_30624,N_25556,N_28187);
nor U30625 (N_30625,N_22953,N_24121);
nand U30626 (N_30626,N_26337,N_28634);
and U30627 (N_30627,N_29636,N_27197);
xnor U30628 (N_30628,N_20476,N_21599);
nor U30629 (N_30629,N_23159,N_29587);
nor U30630 (N_30630,N_27386,N_22472);
or U30631 (N_30631,N_22039,N_29087);
or U30632 (N_30632,N_27885,N_28142);
nor U30633 (N_30633,N_20299,N_24694);
nand U30634 (N_30634,N_22312,N_21617);
or U30635 (N_30635,N_22642,N_25842);
nor U30636 (N_30636,N_21678,N_25518);
xor U30637 (N_30637,N_25361,N_24306);
and U30638 (N_30638,N_27034,N_24703);
or U30639 (N_30639,N_26084,N_20835);
nand U30640 (N_30640,N_28083,N_21444);
xnor U30641 (N_30641,N_23194,N_22163);
or U30642 (N_30642,N_22728,N_20177);
and U30643 (N_30643,N_20126,N_22701);
and U30644 (N_30644,N_22692,N_22564);
and U30645 (N_30645,N_29123,N_22509);
or U30646 (N_30646,N_25146,N_29383);
and U30647 (N_30647,N_29499,N_23365);
and U30648 (N_30648,N_22443,N_28540);
or U30649 (N_30649,N_23762,N_24909);
and U30650 (N_30650,N_22931,N_29449);
or U30651 (N_30651,N_23560,N_26836);
nor U30652 (N_30652,N_26540,N_25432);
and U30653 (N_30653,N_26721,N_20024);
and U30654 (N_30654,N_29849,N_22578);
or U30655 (N_30655,N_28784,N_27767);
and U30656 (N_30656,N_29210,N_22610);
nand U30657 (N_30657,N_21052,N_27219);
nor U30658 (N_30658,N_24124,N_24237);
or U30659 (N_30659,N_29265,N_25574);
nor U30660 (N_30660,N_29909,N_22734);
nor U30661 (N_30661,N_26365,N_26729);
and U30662 (N_30662,N_20964,N_29438);
and U30663 (N_30663,N_24532,N_20724);
and U30664 (N_30664,N_27814,N_20376);
or U30665 (N_30665,N_24761,N_21953);
or U30666 (N_30666,N_26093,N_22479);
nor U30667 (N_30667,N_22333,N_25628);
nor U30668 (N_30668,N_20802,N_27753);
and U30669 (N_30669,N_22048,N_20844);
or U30670 (N_30670,N_29935,N_26551);
nand U30671 (N_30671,N_26933,N_22566);
nor U30672 (N_30672,N_29296,N_23845);
or U30673 (N_30673,N_23615,N_23817);
and U30674 (N_30674,N_25619,N_24548);
or U30675 (N_30675,N_23867,N_21069);
nor U30676 (N_30676,N_20915,N_24986);
nand U30677 (N_30677,N_20946,N_24039);
and U30678 (N_30678,N_25490,N_21710);
nand U30679 (N_30679,N_28810,N_23775);
nand U30680 (N_30680,N_23991,N_28394);
or U30681 (N_30681,N_21342,N_24578);
xor U30682 (N_30682,N_29109,N_23134);
nand U30683 (N_30683,N_22675,N_20269);
nand U30684 (N_30684,N_23066,N_21027);
nand U30685 (N_30685,N_26914,N_23195);
and U30686 (N_30686,N_24740,N_25207);
nand U30687 (N_30687,N_28267,N_26548);
nor U30688 (N_30688,N_22049,N_23092);
and U30689 (N_30689,N_20572,N_29469);
and U30690 (N_30690,N_29938,N_26095);
nand U30691 (N_30691,N_20403,N_22311);
or U30692 (N_30692,N_21986,N_24073);
or U30693 (N_30693,N_28049,N_26338);
and U30694 (N_30694,N_25326,N_25346);
nand U30695 (N_30695,N_20249,N_24056);
xnor U30696 (N_30696,N_27201,N_22293);
or U30697 (N_30697,N_21563,N_28968);
xnor U30698 (N_30698,N_24301,N_29057);
nand U30699 (N_30699,N_22794,N_27999);
nand U30700 (N_30700,N_20426,N_20566);
nand U30701 (N_30701,N_23536,N_23126);
xnor U30702 (N_30702,N_22487,N_22084);
nor U30703 (N_30703,N_24891,N_29289);
or U30704 (N_30704,N_20603,N_28648);
or U30705 (N_30705,N_21693,N_24307);
nand U30706 (N_30706,N_26421,N_21081);
nor U30707 (N_30707,N_25119,N_27351);
or U30708 (N_30708,N_28434,N_22303);
and U30709 (N_30709,N_29660,N_20546);
nor U30710 (N_30710,N_28109,N_21322);
and U30711 (N_30711,N_27095,N_26105);
or U30712 (N_30712,N_20608,N_26524);
and U30713 (N_30713,N_26663,N_21331);
xnor U30714 (N_30714,N_21059,N_20123);
and U30715 (N_30715,N_22128,N_23927);
or U30716 (N_30716,N_23346,N_21714);
and U30717 (N_30717,N_28560,N_27073);
or U30718 (N_30718,N_22866,N_22081);
and U30719 (N_30719,N_26868,N_27744);
or U30720 (N_30720,N_24021,N_20361);
nand U30721 (N_30721,N_23984,N_21704);
xor U30722 (N_30722,N_23909,N_26557);
and U30723 (N_30723,N_26192,N_21955);
nand U30724 (N_30724,N_21787,N_27184);
or U30725 (N_30725,N_26431,N_26623);
and U30726 (N_30726,N_20597,N_29245);
nor U30727 (N_30727,N_23782,N_23910);
nor U30728 (N_30728,N_29437,N_25468);
or U30729 (N_30729,N_28441,N_26314);
nand U30730 (N_30730,N_23872,N_21512);
and U30731 (N_30731,N_23687,N_28965);
or U30732 (N_30732,N_24336,N_26858);
nand U30733 (N_30733,N_26202,N_20857);
nand U30734 (N_30734,N_24751,N_26991);
nand U30735 (N_30735,N_20814,N_26838);
nor U30736 (N_30736,N_21503,N_22581);
nor U30737 (N_30737,N_21448,N_27657);
or U30738 (N_30738,N_29382,N_22880);
nand U30739 (N_30739,N_28944,N_26804);
nand U30740 (N_30740,N_23121,N_26400);
xor U30741 (N_30741,N_23110,N_24141);
nor U30742 (N_30742,N_27109,N_27536);
nand U30743 (N_30743,N_28178,N_28958);
nor U30744 (N_30744,N_20324,N_26255);
and U30745 (N_30745,N_28584,N_23950);
nand U30746 (N_30746,N_20460,N_25220);
and U30747 (N_30747,N_28620,N_21198);
and U30748 (N_30748,N_23171,N_27511);
or U30749 (N_30749,N_21359,N_24057);
nand U30750 (N_30750,N_28206,N_24147);
nor U30751 (N_30751,N_28617,N_26263);
nor U30752 (N_30752,N_23746,N_28383);
nand U30753 (N_30753,N_22968,N_29315);
or U30754 (N_30754,N_25101,N_27224);
xor U30755 (N_30755,N_21294,N_24474);
nand U30756 (N_30756,N_27204,N_24070);
xor U30757 (N_30757,N_28003,N_20548);
and U30758 (N_30758,N_20006,N_25138);
or U30759 (N_30759,N_25478,N_26423);
or U30760 (N_30760,N_26789,N_20507);
or U30761 (N_30761,N_25211,N_20304);
and U30762 (N_30762,N_26126,N_26261);
or U30763 (N_30763,N_22702,N_28301);
nor U30764 (N_30764,N_29760,N_21551);
nor U30765 (N_30765,N_24785,N_27539);
and U30766 (N_30766,N_26592,N_20178);
and U30767 (N_30767,N_28788,N_23226);
and U30768 (N_30768,N_24876,N_21935);
nand U30769 (N_30769,N_28231,N_25925);
and U30770 (N_30770,N_28132,N_22773);
and U30771 (N_30771,N_23961,N_21202);
and U30772 (N_30772,N_27146,N_22234);
nand U30773 (N_30773,N_26457,N_25768);
and U30774 (N_30774,N_29995,N_20444);
and U30775 (N_30775,N_24620,N_29069);
and U30776 (N_30776,N_23446,N_22706);
nor U30777 (N_30777,N_27367,N_28622);
or U30778 (N_30778,N_23410,N_28709);
nand U30779 (N_30779,N_22596,N_29834);
xor U30780 (N_30780,N_22575,N_21066);
nor U30781 (N_30781,N_26443,N_26504);
and U30782 (N_30782,N_21712,N_25880);
or U30783 (N_30783,N_27936,N_22508);
nor U30784 (N_30784,N_24749,N_23083);
nand U30785 (N_30785,N_25234,N_23306);
and U30786 (N_30786,N_26020,N_26727);
nor U30787 (N_30787,N_27082,N_27928);
xnor U30788 (N_30788,N_23177,N_25890);
and U30789 (N_30789,N_22291,N_23163);
or U30790 (N_30790,N_28890,N_26934);
or U30791 (N_30791,N_29187,N_29270);
or U30792 (N_30792,N_28311,N_29698);
xnor U30793 (N_30793,N_21594,N_23214);
and U30794 (N_30794,N_26834,N_27307);
xor U30795 (N_30795,N_22284,N_23115);
and U30796 (N_30796,N_20737,N_21569);
nand U30797 (N_30797,N_28826,N_24849);
nor U30798 (N_30798,N_22678,N_25788);
or U30799 (N_30799,N_21147,N_20971);
nand U30800 (N_30800,N_29593,N_25600);
and U30801 (N_30801,N_23273,N_26372);
nor U30802 (N_30802,N_27725,N_29754);
nand U30803 (N_30803,N_24187,N_29592);
nor U30804 (N_30804,N_23103,N_20474);
or U30805 (N_30805,N_27820,N_25339);
xor U30806 (N_30806,N_24801,N_23357);
and U30807 (N_30807,N_20272,N_26748);
or U30808 (N_30808,N_23592,N_21420);
nor U30809 (N_30809,N_26090,N_22403);
or U30810 (N_30810,N_28931,N_20720);
and U30811 (N_30811,N_29681,N_26738);
nor U30812 (N_30812,N_20071,N_29818);
xor U30813 (N_30813,N_28659,N_29118);
and U30814 (N_30814,N_20852,N_20162);
nand U30815 (N_30815,N_24211,N_24559);
or U30816 (N_30816,N_25709,N_22242);
or U30817 (N_30817,N_26417,N_26073);
or U30818 (N_30818,N_25627,N_27606);
or U30819 (N_30819,N_23200,N_28424);
and U30820 (N_30820,N_24951,N_24890);
xnor U30821 (N_30821,N_25863,N_28149);
nor U30822 (N_30822,N_26712,N_25465);
and U30823 (N_30823,N_26248,N_29676);
and U30824 (N_30824,N_21271,N_27498);
or U30825 (N_30825,N_20208,N_27496);
or U30826 (N_30826,N_25304,N_29816);
and U30827 (N_30827,N_24092,N_21246);
nand U30828 (N_30828,N_25686,N_20121);
nor U30829 (N_30829,N_28050,N_26019);
nor U30830 (N_30830,N_25776,N_29581);
nand U30831 (N_30831,N_28951,N_23840);
nand U30832 (N_30832,N_28514,N_28715);
nor U30833 (N_30833,N_23828,N_24558);
and U30834 (N_30834,N_25155,N_23575);
or U30835 (N_30835,N_24967,N_28851);
xor U30836 (N_30836,N_21785,N_24186);
nand U30837 (N_30837,N_20239,N_29553);
nand U30838 (N_30838,N_21734,N_20655);
or U30839 (N_30839,N_20025,N_27678);
or U30840 (N_30840,N_26188,N_27787);
and U30841 (N_30841,N_25195,N_26903);
nor U30842 (N_30842,N_21049,N_28364);
nand U30843 (N_30843,N_25313,N_20860);
and U30844 (N_30844,N_20391,N_26531);
nand U30845 (N_30845,N_24396,N_20619);
nor U30846 (N_30846,N_22059,N_20769);
or U30847 (N_30847,N_23952,N_25400);
nor U30848 (N_30848,N_23573,N_24312);
nor U30849 (N_30849,N_26175,N_24324);
nand U30850 (N_30850,N_29538,N_26580);
or U30851 (N_30851,N_22166,N_26752);
nand U30852 (N_30852,N_25262,N_25568);
nand U30853 (N_30853,N_23105,N_20477);
nor U30854 (N_30854,N_21247,N_24671);
nand U30855 (N_30855,N_27574,N_26035);
nor U30856 (N_30856,N_24075,N_20365);
and U30857 (N_30857,N_23133,N_27958);
nand U30858 (N_30858,N_24618,N_21215);
nand U30859 (N_30859,N_23179,N_25099);
or U30860 (N_30860,N_21031,N_22956);
nor U30861 (N_30861,N_29642,N_22342);
or U30862 (N_30862,N_28737,N_21419);
and U30863 (N_30863,N_20490,N_22340);
and U30864 (N_30864,N_28318,N_27009);
nor U30865 (N_30865,N_20945,N_27422);
nand U30866 (N_30866,N_23641,N_26028);
xnor U30867 (N_30867,N_28431,N_24711);
nor U30868 (N_30868,N_24200,N_20878);
nand U30869 (N_30869,N_20418,N_24169);
xor U30870 (N_30870,N_20088,N_28440);
nor U30871 (N_30871,N_25779,N_28665);
xor U30872 (N_30872,N_27179,N_21876);
xnor U30873 (N_30873,N_22001,N_22310);
and U30874 (N_30874,N_20809,N_27861);
nor U30875 (N_30875,N_24493,N_25104);
nor U30876 (N_30876,N_24762,N_21151);
nand U30877 (N_30877,N_25135,N_21501);
nand U30878 (N_30878,N_26351,N_27084);
or U30879 (N_30879,N_21699,N_24471);
or U30880 (N_30880,N_27245,N_20323);
nor U30881 (N_30881,N_21369,N_26871);
and U30882 (N_30882,N_27028,N_29411);
or U30883 (N_30883,N_25122,N_29653);
and U30884 (N_30884,N_20423,N_23533);
xnor U30885 (N_30885,N_25564,N_21427);
xnor U30886 (N_30886,N_28447,N_24537);
nand U30887 (N_30887,N_26972,N_26231);
nor U30888 (N_30888,N_24033,N_27236);
or U30889 (N_30889,N_20358,N_24374);
nor U30890 (N_30890,N_24639,N_25435);
nand U30891 (N_30891,N_27775,N_22574);
or U30892 (N_30892,N_22359,N_26656);
and U30893 (N_30893,N_23255,N_28124);
nand U30894 (N_30894,N_20838,N_29269);
nand U30895 (N_30895,N_29629,N_24257);
or U30896 (N_30896,N_24014,N_23039);
nand U30897 (N_30897,N_27414,N_27385);
and U30898 (N_30898,N_29040,N_21570);
and U30899 (N_30899,N_27542,N_27140);
and U30900 (N_30900,N_26807,N_22899);
xor U30901 (N_30901,N_20707,N_23932);
or U30902 (N_30902,N_24360,N_21068);
nor U30903 (N_30903,N_25720,N_26132);
xnor U30904 (N_30904,N_27182,N_27227);
or U30905 (N_30905,N_24959,N_24418);
nand U30906 (N_30906,N_28293,N_24246);
nor U30907 (N_30907,N_27024,N_24582);
nor U30908 (N_30908,N_20812,N_28265);
and U30909 (N_30909,N_22946,N_21110);
nor U30910 (N_30910,N_25591,N_21034);
nor U30911 (N_30911,N_23537,N_29641);
or U30912 (N_30912,N_27875,N_26949);
and U30913 (N_30913,N_27604,N_20113);
xor U30914 (N_30914,N_20823,N_24672);
or U30915 (N_30915,N_23464,N_24079);
or U30916 (N_30916,N_27532,N_29624);
nand U30917 (N_30917,N_29141,N_23690);
nor U30918 (N_30918,N_21893,N_23169);
or U30919 (N_30919,N_25921,N_29738);
nor U30920 (N_30920,N_25036,N_23855);
nand U30921 (N_30921,N_28411,N_23296);
nand U30922 (N_30922,N_26467,N_21079);
and U30923 (N_30923,N_23473,N_26281);
xor U30924 (N_30924,N_23322,N_22935);
nand U30925 (N_30925,N_26731,N_20557);
nor U30926 (N_30926,N_26960,N_26869);
nor U30927 (N_30927,N_25265,N_22521);
and U30928 (N_30928,N_28408,N_26017);
nor U30929 (N_30929,N_29667,N_29419);
or U30930 (N_30930,N_25431,N_27789);
nor U30931 (N_30931,N_27431,N_27086);
and U30932 (N_30932,N_26412,N_22511);
and U30933 (N_30933,N_22273,N_27100);
or U30934 (N_30934,N_26247,N_29195);
nor U30935 (N_30935,N_27217,N_29548);
or U30936 (N_30936,N_24894,N_23602);
xor U30937 (N_30937,N_29948,N_25513);
or U30938 (N_30938,N_25245,N_24903);
or U30939 (N_30939,N_25930,N_23388);
and U30940 (N_30940,N_26673,N_29168);
nor U30941 (N_30941,N_27615,N_27720);
or U30942 (N_30942,N_24164,N_27007);
and U30943 (N_30943,N_21372,N_25344);
or U30944 (N_30944,N_21368,N_26781);
or U30945 (N_30945,N_29675,N_20218);
nor U30946 (N_30946,N_28544,N_26535);
nor U30947 (N_30947,N_21145,N_20637);
and U30948 (N_30948,N_28517,N_24231);
nand U30949 (N_30949,N_25035,N_23995);
and U30950 (N_30950,N_23362,N_27191);
nand U30951 (N_30951,N_26151,N_28924);
nand U30952 (N_30952,N_27880,N_24078);
nand U30953 (N_30953,N_29577,N_29879);
nor U30954 (N_30954,N_20347,N_25810);
nor U30955 (N_30955,N_20059,N_22412);
or U30956 (N_30956,N_29436,N_26588);
nor U30957 (N_30957,N_21469,N_20839);
nand U30958 (N_30958,N_25089,N_22640);
or U30959 (N_30959,N_27136,N_23455);
or U30960 (N_30960,N_22061,N_29058);
or U30961 (N_30961,N_22920,N_22250);
nor U30962 (N_30962,N_26756,N_23574);
or U30963 (N_30963,N_20583,N_24146);
nand U30964 (N_30964,N_28711,N_29725);
or U30965 (N_30965,N_21239,N_22345);
and U30966 (N_30966,N_25561,N_29481);
nor U30967 (N_30967,N_28645,N_20228);
nand U30968 (N_30968,N_25639,N_25018);
nor U30969 (N_30969,N_21201,N_29810);
nor U30970 (N_30970,N_22471,N_26433);
xor U30971 (N_30971,N_21183,N_23384);
nor U30972 (N_30972,N_22373,N_26840);
nor U30973 (N_30973,N_26189,N_20580);
and U30974 (N_30974,N_26885,N_29785);
nor U30975 (N_30975,N_24995,N_27644);
and U30976 (N_30976,N_24411,N_26139);
nor U30977 (N_30977,N_23165,N_25350);
nor U30978 (N_30978,N_23637,N_23607);
nand U30979 (N_30979,N_22064,N_26407);
nor U30980 (N_30980,N_29031,N_26492);
nor U30981 (N_30981,N_26603,N_26598);
nor U30982 (N_30982,N_23029,N_26747);
or U30983 (N_30983,N_23571,N_28846);
nand U30984 (N_30984,N_29772,N_22525);
xor U30985 (N_30985,N_28428,N_23901);
and U30986 (N_30986,N_29305,N_24824);
nand U30987 (N_30987,N_24261,N_27472);
nor U30988 (N_30988,N_27460,N_20449);
and U30989 (N_30989,N_22820,N_29666);
or U30990 (N_30990,N_21474,N_25815);
nor U30991 (N_30991,N_28163,N_23118);
nor U30992 (N_30992,N_20240,N_29522);
nand U30993 (N_30993,N_21873,N_29166);
nand U30994 (N_30994,N_26549,N_29800);
nor U30995 (N_30995,N_24520,N_21218);
xor U30996 (N_30996,N_22183,N_26195);
nand U30997 (N_30997,N_25907,N_20387);
and U30998 (N_30998,N_27171,N_25953);
and U30999 (N_30999,N_27501,N_20409);
xnor U31000 (N_31000,N_29610,N_21812);
or U31001 (N_31001,N_24725,N_26128);
nor U31002 (N_31002,N_25023,N_22767);
nor U31003 (N_31003,N_28374,N_26468);
nor U31004 (N_31004,N_23568,N_27141);
and U31005 (N_31005,N_22215,N_20188);
or U31006 (N_31006,N_20932,N_27556);
nand U31007 (N_31007,N_29131,N_26112);
nor U31008 (N_31008,N_28479,N_27647);
and U31009 (N_31009,N_23655,N_27954);
nor U31010 (N_31010,N_28200,N_28207);
nor U31011 (N_31011,N_28998,N_21966);
or U31012 (N_31012,N_20889,N_26476);
xor U31013 (N_31013,N_24709,N_20122);
and U31014 (N_31014,N_22346,N_21308);
or U31015 (N_31015,N_20586,N_22362);
or U31016 (N_31016,N_23052,N_28165);
or U31017 (N_31017,N_27274,N_29625);
nor U31018 (N_31018,N_21951,N_27842);
xor U31019 (N_31019,N_28123,N_21402);
nor U31020 (N_31020,N_28069,N_21690);
nor U31021 (N_31021,N_21775,N_24165);
nand U31022 (N_31022,N_24258,N_21422);
nor U31023 (N_31023,N_24566,N_21793);
nor U31024 (N_31024,N_20217,N_21275);
and U31025 (N_31025,N_27202,N_23679);
and U31026 (N_31026,N_22609,N_24329);
xor U31027 (N_31027,N_24794,N_21738);
and U31028 (N_31028,N_20796,N_29189);
nor U31029 (N_31029,N_27627,N_28926);
xnor U31030 (N_31030,N_21242,N_28952);
nor U31031 (N_31031,N_26870,N_23123);
nand U31032 (N_31032,N_21767,N_25044);
nor U31033 (N_31033,N_22195,N_28060);
nand U31034 (N_31034,N_24741,N_26021);
nand U31035 (N_31035,N_28324,N_25852);
or U31036 (N_31036,N_22591,N_20887);
or U31037 (N_31037,N_22017,N_29514);
nand U31038 (N_31038,N_22704,N_23424);
nand U31039 (N_31039,N_27260,N_28256);
or U31040 (N_31040,N_24173,N_20606);
or U31041 (N_31041,N_29316,N_26671);
and U31042 (N_31042,N_28180,N_21801);
nor U31043 (N_31043,N_27145,N_22054);
or U31044 (N_31044,N_28975,N_27748);
nor U31045 (N_31045,N_28666,N_29344);
or U31046 (N_31046,N_24929,N_24320);
or U31047 (N_31047,N_20540,N_22087);
nor U31048 (N_31048,N_26483,N_23252);
nand U31049 (N_31049,N_26466,N_24834);
or U31050 (N_31050,N_22665,N_20489);
and U31051 (N_31051,N_27231,N_26703);
and U31052 (N_31052,N_22747,N_27643);
or U31053 (N_31053,N_21302,N_21470);
or U31054 (N_31054,N_26728,N_22758);
and U31055 (N_31055,N_25393,N_27724);
and U31056 (N_31056,N_24206,N_20336);
or U31057 (N_31057,N_29034,N_26169);
or U31058 (N_31058,N_20885,N_25681);
nor U31059 (N_31059,N_23471,N_25143);
nand U31060 (N_31060,N_24088,N_22977);
nand U31061 (N_31061,N_20008,N_21828);
nand U31062 (N_31062,N_21552,N_27466);
and U31063 (N_31063,N_25928,N_23228);
and U31064 (N_31064,N_23185,N_22203);
xnor U31065 (N_31065,N_25548,N_21804);
or U31066 (N_31066,N_23501,N_27813);
or U31067 (N_31067,N_29953,N_22026);
nand U31068 (N_31068,N_27216,N_29337);
nor U31069 (N_31069,N_26576,N_26264);
xor U31070 (N_31070,N_29474,N_28466);
and U31071 (N_31071,N_29475,N_25505);
nand U31072 (N_31072,N_24842,N_27180);
or U31073 (N_31073,N_21637,N_20790);
or U31074 (N_31074,N_24770,N_26196);
nand U31075 (N_31075,N_28152,N_24564);
or U31076 (N_31076,N_21395,N_28903);
xor U31077 (N_31077,N_28313,N_23765);
or U31078 (N_31078,N_21214,N_26977);
nor U31079 (N_31079,N_26058,N_23772);
and U31080 (N_31080,N_28988,N_21379);
nor U31081 (N_31081,N_22414,N_28219);
nor U31082 (N_31082,N_24992,N_23548);
or U31083 (N_31083,N_28882,N_23321);
nand U31084 (N_31084,N_25162,N_24224);
and U31085 (N_31085,N_22838,N_22184);
nor U31086 (N_31086,N_28169,N_24054);
or U31087 (N_31087,N_29801,N_23776);
or U31088 (N_31088,N_29104,N_28533);
nor U31089 (N_31089,N_25085,N_29143);
nor U31090 (N_31090,N_28556,N_27118);
nor U31091 (N_31091,N_29971,N_23742);
and U31092 (N_31092,N_28987,N_27375);
nor U31093 (N_31093,N_22229,N_28920);
and U31094 (N_31094,N_29797,N_29980);
xor U31095 (N_31095,N_29487,N_21933);
nor U31096 (N_31096,N_29161,N_24182);
or U31097 (N_31097,N_20829,N_20556);
nand U31098 (N_31098,N_21683,N_24830);
and U31099 (N_31099,N_25537,N_22868);
nor U31100 (N_31100,N_22551,N_27477);
or U31101 (N_31101,N_22784,N_29188);
and U31102 (N_31102,N_27970,N_21133);
and U31103 (N_31103,N_29952,N_21963);
nand U31104 (N_31104,N_21479,N_20762);
or U31105 (N_31105,N_26000,N_22862);
nand U31106 (N_31106,N_21325,N_24234);
and U31107 (N_31107,N_22276,N_21316);
xnor U31108 (N_31108,N_23946,N_26814);
xor U31109 (N_31109,N_29893,N_26391);
nand U31110 (N_31110,N_22171,N_25226);
or U31111 (N_31111,N_26904,N_29486);
nand U31112 (N_31112,N_25915,N_27636);
nor U31113 (N_31113,N_21632,N_22056);
nand U31114 (N_31114,N_20650,N_27358);
and U31115 (N_31115,N_25456,N_21647);
nor U31116 (N_31116,N_26742,N_28416);
or U31117 (N_31117,N_27006,N_21404);
xor U31118 (N_31118,N_25877,N_25115);
nand U31119 (N_31119,N_25421,N_21696);
nor U31120 (N_31120,N_28457,N_20237);
or U31121 (N_31121,N_28588,N_25178);
xor U31122 (N_31122,N_27249,N_27675);
or U31123 (N_31123,N_20811,N_20996);
nand U31124 (N_31124,N_25787,N_24482);
or U31125 (N_31125,N_22965,N_22502);
and U31126 (N_31126,N_26002,N_24798);
nor U31127 (N_31127,N_26788,N_20710);
and U31128 (N_31128,N_23119,N_24669);
nor U31129 (N_31129,N_28167,N_25992);
and U31130 (N_31130,N_25783,N_29578);
and U31131 (N_31131,N_26101,N_28683);
or U31132 (N_31132,N_23895,N_29452);
nand U31133 (N_31133,N_27930,N_28935);
nor U31134 (N_31134,N_27995,N_20265);
or U31135 (N_31135,N_27014,N_22432);
xor U31136 (N_31136,N_25444,N_28861);
nor U31137 (N_31137,N_22230,N_29989);
or U31138 (N_31138,N_22967,N_29693);
or U31139 (N_31139,N_26777,N_25679);
or U31140 (N_31140,N_29717,N_22445);
and U31141 (N_31141,N_27483,N_20988);
nor U31142 (N_31142,N_29792,N_25422);
and U31143 (N_31143,N_21922,N_23458);
and U31144 (N_31144,N_28234,N_26791);
nor U31145 (N_31145,N_20000,N_23034);
or U31146 (N_31146,N_29200,N_22599);
or U31147 (N_31147,N_22850,N_25486);
nor U31148 (N_31148,N_24641,N_22269);
and U31149 (N_31149,N_23502,N_28158);
nor U31150 (N_31150,N_23724,N_28605);
and U31151 (N_31151,N_22164,N_22170);
nor U31152 (N_31152,N_21091,N_28162);
xnor U31153 (N_31153,N_20260,N_27419);
nand U31154 (N_31154,N_27949,N_22626);
or U31155 (N_31155,N_29429,N_21969);
nand U31156 (N_31156,N_20590,N_20993);
and U31157 (N_31157,N_24494,N_28390);
nand U31158 (N_31158,N_27021,N_29111);
nand U31159 (N_31159,N_22198,N_21137);
nand U31160 (N_31160,N_26378,N_26484);
nor U31161 (N_31161,N_29990,N_28705);
and U31162 (N_31162,N_20613,N_27519);
and U31163 (N_31163,N_23880,N_25331);
nand U31164 (N_31164,N_25107,N_24601);
and U31165 (N_31165,N_22126,N_28929);
nor U31166 (N_31166,N_27139,N_29626);
and U31167 (N_31167,N_22460,N_26250);
nand U31168 (N_31168,N_29271,N_21296);
nor U31169 (N_31169,N_28914,N_22725);
xnor U31170 (N_31170,N_28895,N_29129);
nor U31171 (N_31171,N_20026,N_26328);
or U31172 (N_31172,N_26127,N_26806);
nor U31173 (N_31173,N_29236,N_20043);
and U31174 (N_31174,N_22960,N_22464);
xor U31175 (N_31175,N_29857,N_20738);
nor U31176 (N_31176,N_23091,N_22238);
nand U31177 (N_31177,N_23347,N_29276);
and U31178 (N_31178,N_26121,N_26994);
or U31179 (N_31179,N_24859,N_27903);
or U31180 (N_31180,N_28770,N_23004);
nand U31181 (N_31181,N_22417,N_28954);
nand U31182 (N_31182,N_23564,N_27461);
or U31183 (N_31183,N_22133,N_21917);
and U31184 (N_31184,N_23056,N_22027);
nand U31185 (N_31185,N_24285,N_28899);
or U31186 (N_31186,N_24933,N_24008);
and U31187 (N_31187,N_23385,N_24464);
nor U31188 (N_31188,N_20909,N_22851);
or U31189 (N_31189,N_27927,N_25081);
nor U31190 (N_31190,N_22576,N_22466);
xnor U31191 (N_31191,N_27036,N_22292);
and U31192 (N_31192,N_28639,N_29970);
nor U31193 (N_31193,N_28589,N_23958);
nand U31194 (N_31194,N_28435,N_28979);
or U31195 (N_31195,N_26778,N_22631);
xnor U31196 (N_31196,N_21582,N_25132);
and U31197 (N_31197,N_22688,N_27162);
nor U31198 (N_31198,N_27177,N_28048);
xor U31199 (N_31199,N_25898,N_26300);
nor U31200 (N_31200,N_22650,N_29840);
xor U31201 (N_31201,N_28372,N_27452);
and U31202 (N_31202,N_25887,N_26954);
nor U31203 (N_31203,N_22641,N_28650);
or U31204 (N_31204,N_29228,N_23355);
nand U31205 (N_31205,N_29844,N_26500);
and U31206 (N_31206,N_20676,N_26874);
xnor U31207 (N_31207,N_25280,N_28649);
or U31208 (N_31208,N_29763,N_29749);
nor U31209 (N_31209,N_26619,N_25706);
nor U31210 (N_31210,N_28398,N_21273);
nor U31211 (N_31211,N_28512,N_25790);
nand U31212 (N_31212,N_27340,N_21652);
and U31213 (N_31213,N_21434,N_20425);
and U31214 (N_31214,N_21695,N_26381);
or U31215 (N_31215,N_25713,N_20202);
nor U31216 (N_31216,N_28800,N_27900);
nand U31217 (N_31217,N_28121,N_20601);
and U31218 (N_31218,N_20355,N_24428);
nor U31219 (N_31219,N_27706,N_20266);
nand U31220 (N_31220,N_29273,N_20777);
and U31221 (N_31221,N_29183,N_21633);
xor U31222 (N_31222,N_28470,N_26427);
nor U31223 (N_31223,N_27213,N_29777);
or U31224 (N_31224,N_27434,N_28254);
nand U31225 (N_31225,N_23407,N_21341);
xnor U31226 (N_31226,N_25106,N_22891);
or U31227 (N_31227,N_27441,N_25380);
or U31228 (N_31228,N_29949,N_28493);
nor U31229 (N_31229,N_28058,N_24867);
nor U31230 (N_31230,N_29252,N_29460);
or U31231 (N_31231,N_28698,N_26415);
nand U31232 (N_31232,N_26944,N_20782);
and U31233 (N_31233,N_23231,N_29157);
and U31234 (N_31234,N_20747,N_20150);
or U31235 (N_31235,N_29185,N_25306);
nor U31236 (N_31236,N_26505,N_21187);
nor U31237 (N_31237,N_24925,N_28303);
and U31238 (N_31238,N_27791,N_24436);
nor U31239 (N_31239,N_22144,N_26087);
and U31240 (N_31240,N_21573,N_23201);
nand U31241 (N_31241,N_22252,N_22062);
nor U31242 (N_31242,N_27746,N_24599);
or U31243 (N_31243,N_27945,N_28680);
and U31244 (N_31244,N_26083,N_26029);
xnor U31245 (N_31245,N_21168,N_23303);
or U31246 (N_31246,N_29775,N_20892);
or U31247 (N_31247,N_29755,N_27896);
nand U31248 (N_31248,N_23311,N_22938);
or U31249 (N_31249,N_22394,N_25370);
or U31250 (N_31250,N_24431,N_20773);
xnor U31251 (N_31251,N_21837,N_27233);
or U31252 (N_31252,N_26928,N_27475);
or U31253 (N_31253,N_28515,N_21312);
nand U31254 (N_31254,N_21548,N_22727);
and U31255 (N_31255,N_20311,N_23856);
or U31256 (N_31256,N_21976,N_29408);
or U31257 (N_31257,N_27867,N_27825);
and U31258 (N_31258,N_24962,N_24038);
or U31259 (N_31259,N_24412,N_29095);
nor U31260 (N_31260,N_25873,N_26406);
nor U31261 (N_31261,N_26537,N_20589);
nor U31262 (N_31262,N_26995,N_26734);
or U31263 (N_31263,N_27208,N_22290);
xor U31264 (N_31264,N_25609,N_22623);
xor U31265 (N_31265,N_25127,N_29410);
nand U31266 (N_31266,N_20011,N_20766);
or U31267 (N_31267,N_20415,N_27594);
nor U31268 (N_31268,N_26226,N_29509);
or U31269 (N_31269,N_28692,N_29942);
xnor U31270 (N_31270,N_25663,N_24433);
nand U31271 (N_31271,N_28212,N_24635);
or U31272 (N_31272,N_23104,N_24945);
nor U31273 (N_31273,N_29164,N_23720);
nand U31274 (N_31274,N_26984,N_28264);
nor U31275 (N_31275,N_21178,N_24775);
nor U31276 (N_31276,N_23428,N_27658);
or U31277 (N_31277,N_27870,N_29598);
or U31278 (N_31278,N_20751,N_28960);
nand U31279 (N_31279,N_29547,N_23711);
or U31280 (N_31280,N_25389,N_29661);
and U31281 (N_31281,N_25901,N_22830);
and U31282 (N_31282,N_26864,N_23562);
and U31283 (N_31283,N_28796,N_20972);
xnor U31284 (N_31284,N_25540,N_28384);
xor U31285 (N_31285,N_27039,N_26826);
and U31286 (N_31286,N_23590,N_21771);
xor U31287 (N_31287,N_27629,N_25152);
or U31288 (N_31288,N_21724,N_29517);
nor U31289 (N_31289,N_25576,N_27425);
nor U31290 (N_31290,N_27334,N_29910);
or U31291 (N_31291,N_27792,N_25977);
and U31292 (N_31292,N_26653,N_29378);
nand U31293 (N_31293,N_26759,N_21191);
nor U31294 (N_31294,N_24082,N_24139);
or U31295 (N_31295,N_27152,N_26023);
nand U31296 (N_31296,N_21989,N_25521);
nor U31297 (N_31297,N_26135,N_22670);
nor U31298 (N_31298,N_22313,N_21197);
nand U31299 (N_31299,N_25166,N_26888);
and U31300 (N_31300,N_21115,N_29278);
nand U31301 (N_31301,N_21063,N_28747);
nor U31302 (N_31302,N_26496,N_24112);
nor U31303 (N_31303,N_23948,N_29798);
xor U31304 (N_31304,N_28933,N_20752);
and U31305 (N_31305,N_25824,N_21773);
or U31306 (N_31306,N_29734,N_25677);
and U31307 (N_31307,N_23172,N_20096);
and U31308 (N_31308,N_24881,N_23457);
and U31309 (N_31309,N_28190,N_22823);
and U31310 (N_31310,N_26790,N_29015);
nand U31311 (N_31311,N_25399,N_21459);
and U31312 (N_31312,N_25480,N_27174);
nor U31313 (N_31313,N_24784,N_27586);
and U31314 (N_31314,N_28676,N_23569);
xnor U31315 (N_31315,N_22435,N_24948);
nand U31316 (N_31316,N_21204,N_27796);
nor U31317 (N_31317,N_21895,N_27714);
xor U31318 (N_31318,N_27151,N_25429);
nor U31319 (N_31319,N_24479,N_29823);
or U31320 (N_31320,N_23379,N_27924);
and U31321 (N_31321,N_29350,N_29691);
nand U31322 (N_31322,N_23339,N_24783);
nor U31323 (N_31323,N_23862,N_26212);
and U31324 (N_31324,N_28657,N_21748);
and U31325 (N_31325,N_25330,N_22996);
or U31326 (N_31326,N_21740,N_23601);
or U31327 (N_31327,N_24235,N_20238);
and U31328 (N_31328,N_20923,N_29926);
and U31329 (N_31329,N_28247,N_22542);
nor U31330 (N_31330,N_27859,N_24803);
nor U31331 (N_31331,N_28494,N_24247);
or U31332 (N_31332,N_20783,N_20628);
or U31333 (N_31333,N_28404,N_27154);
nor U31334 (N_31334,N_24145,N_23277);
or U31335 (N_31335,N_20532,N_26704);
nor U31336 (N_31336,N_26026,N_27553);
and U31337 (N_31337,N_21984,N_26694);
nand U31338 (N_31338,N_25535,N_22577);
xnor U31339 (N_31339,N_25368,N_23868);
nor U31340 (N_31340,N_28308,N_26016);
or U31341 (N_31341,N_26031,N_25288);
nor U31342 (N_31342,N_20662,N_20010);
and U31343 (N_31343,N_26379,N_29826);
or U31344 (N_31344,N_22295,N_25976);
or U31345 (N_31345,N_23796,N_24215);
or U31346 (N_31346,N_20094,N_23697);
nor U31347 (N_31347,N_23905,N_28450);
or U31348 (N_31348,N_29588,N_25342);
nor U31349 (N_31349,N_29631,N_25775);
nand U31350 (N_31350,N_28086,N_24587);
nand U31351 (N_31351,N_26303,N_23904);
nor U31352 (N_31352,N_28464,N_25491);
and U31353 (N_31353,N_28888,N_25763);
nand U31354 (N_31354,N_20114,N_22018);
nand U31355 (N_31355,N_22558,N_27113);
xor U31356 (N_31356,N_25738,N_20922);
or U31357 (N_31357,N_26900,N_24195);
nor U31358 (N_31358,N_29654,N_27520);
and U31359 (N_31359,N_21291,N_24766);
and U31360 (N_31360,N_27850,N_28463);
and U31361 (N_31361,N_24328,N_24287);
nand U31362 (N_31362,N_27901,N_24027);
and U31363 (N_31363,N_28174,N_27106);
and U31364 (N_31364,N_24302,N_22951);
nand U31365 (N_31365,N_28287,N_24481);
xor U31366 (N_31366,N_22870,N_28334);
nor U31367 (N_31367,N_24346,N_28459);
xnor U31368 (N_31368,N_23314,N_25294);
and U31369 (N_31369,N_22155,N_25045);
nor U31370 (N_31370,N_29512,N_26660);
and U31371 (N_31371,N_20327,N_28566);
nand U31372 (N_31372,N_22981,N_25669);
nand U31373 (N_31373,N_26512,N_24610);
nand U31374 (N_31374,N_28750,N_25693);
or U31375 (N_31375,N_28672,N_24492);
and U31376 (N_31376,N_29250,N_25033);
and U31377 (N_31377,N_20807,N_21185);
or U31378 (N_31378,N_20244,N_23890);
or U31379 (N_31379,N_22325,N_26676);
nand U31380 (N_31380,N_28358,N_21515);
or U31381 (N_31381,N_27755,N_22397);
nand U31382 (N_31382,N_28171,N_27838);
xnor U31383 (N_31383,N_27327,N_22483);
and U31384 (N_31384,N_29056,N_29711);
and U31385 (N_31385,N_25100,N_27469);
and U31386 (N_31386,N_27232,N_20373);
nor U31387 (N_31387,N_24325,N_28415);
xor U31388 (N_31388,N_20975,N_22881);
nor U31389 (N_31389,N_21796,N_26867);
or U31390 (N_31390,N_26410,N_21307);
nor U31391 (N_31391,N_23584,N_25238);
nor U31392 (N_31392,N_25791,N_27864);
nand U31393 (N_31393,N_29304,N_20104);
nand U31394 (N_31394,N_25398,N_22954);
and U31395 (N_31395,N_20561,N_21047);
and U31396 (N_31396,N_27719,N_21506);
nor U31397 (N_31397,N_25647,N_21819);
and U31398 (N_31398,N_28403,N_20184);
nand U31399 (N_31399,N_22154,N_28458);
nor U31400 (N_31400,N_26342,N_22606);
xnor U31401 (N_31401,N_23757,N_21886);
or U31402 (N_31402,N_29417,N_27563);
xor U31403 (N_31403,N_28572,N_27618);
or U31404 (N_31404,N_23979,N_25522);
nand U31405 (N_31405,N_24055,N_27528);
xor U31406 (N_31406,N_25038,N_23188);
or U31407 (N_31407,N_23218,N_26893);
nor U31408 (N_31408,N_25066,N_20210);
and U31409 (N_31409,N_21892,N_25168);
and U31410 (N_31410,N_25754,N_21958);
xor U31411 (N_31411,N_21255,N_28863);
or U31412 (N_31412,N_21662,N_23098);
nor U31413 (N_31413,N_22074,N_25629);
nand U31414 (N_31414,N_21175,N_24351);
xnor U31415 (N_31415,N_28930,N_22527);
xor U31416 (N_31416,N_28696,N_23026);
and U31417 (N_31417,N_29478,N_28995);
and U31418 (N_31418,N_29133,N_26156);
and U31419 (N_31419,N_29457,N_20968);
and U31420 (N_31420,N_20053,N_23482);
nand U31421 (N_31421,N_29096,N_20446);
nor U31422 (N_31422,N_22202,N_21165);
xnor U31423 (N_31423,N_22000,N_25275);
and U31424 (N_31424,N_23630,N_22217);
and U31425 (N_31425,N_28432,N_24500);
and U31426 (N_31426,N_24676,N_20742);
nand U31427 (N_31427,N_20453,N_26399);
or U31428 (N_31428,N_28456,N_20192);
nand U31429 (N_31429,N_29895,N_28848);
or U31430 (N_31430,N_25314,N_28213);
nand U31431 (N_31431,N_20062,N_23217);
or U31432 (N_31432,N_22753,N_21557);
and U31433 (N_31433,N_29045,N_27246);
or U31434 (N_31434,N_29247,N_25908);
and U31435 (N_31435,N_20145,N_24621);
nor U31436 (N_31436,N_25807,N_28044);
and U31437 (N_31437,N_22241,N_25203);
or U31438 (N_31438,N_22162,N_29687);
and U31439 (N_31439,N_22469,N_20520);
xnor U31440 (N_31440,N_24443,N_28909);
nand U31441 (N_31441,N_29017,N_20516);
or U31442 (N_31442,N_21389,N_21675);
and U31443 (N_31443,N_20414,N_26635);
xor U31444 (N_31444,N_29646,N_21207);
and U31445 (N_31445,N_24399,N_28623);
nor U31446 (N_31446,N_25615,N_25672);
nor U31447 (N_31447,N_26100,N_27161);
and U31448 (N_31448,N_21407,N_20741);
nand U31449 (N_31449,N_23595,N_26360);
nand U31450 (N_31450,N_27001,N_27549);
nand U31451 (N_31451,N_29992,N_22560);
nand U31452 (N_31452,N_22554,N_20732);
or U31453 (N_31453,N_22211,N_24619);
and U31454 (N_31454,N_25293,N_25159);
nand U31455 (N_31455,N_24708,N_24413);
and U31456 (N_31456,N_21848,N_20936);
and U31457 (N_31457,N_21716,N_29459);
or U31458 (N_31458,N_24533,N_25654);
or U31459 (N_31459,N_29954,N_22503);
and U31460 (N_31460,N_21018,N_24726);
nand U31461 (N_31461,N_21162,N_23618);
nand U31462 (N_31462,N_21559,N_26699);
or U31463 (N_31463,N_27043,N_20070);
or U31464 (N_31464,N_28654,N_27802);
or U31465 (N_31465,N_29492,N_29867);
xor U31466 (N_31466,N_20925,N_21336);
nand U31467 (N_31467,N_23439,N_20931);
or U31468 (N_31468,N_24654,N_29368);
or U31469 (N_31469,N_25762,N_20746);
xor U31470 (N_31470,N_20939,N_23955);
nor U31471 (N_31471,N_22347,N_22989);
nand U31472 (N_31472,N_26739,N_22193);
nor U31473 (N_31473,N_27026,N_27824);
and U31474 (N_31474,N_24873,N_22733);
nor U31475 (N_31475,N_29476,N_27582);
xnor U31476 (N_31476,N_27362,N_21733);
or U31477 (N_31477,N_28262,N_28412);
nand U31478 (N_31478,N_29050,N_29958);
nor U31479 (N_31479,N_26561,N_23063);
nand U31480 (N_31480,N_20380,N_26763);
nand U31481 (N_31481,N_26800,N_23735);
and U31482 (N_31482,N_26367,N_25263);
or U31483 (N_31483,N_21189,N_24273);
nor U31484 (N_31484,N_24895,N_26905);
nand U31485 (N_31485,N_22013,N_21161);
nor U31486 (N_31486,N_21596,N_28887);
and U31487 (N_31487,N_21056,N_29851);
and U31488 (N_31488,N_26658,N_28215);
or U31489 (N_31489,N_24832,N_25658);
and U31490 (N_31490,N_29431,N_27305);
or U31491 (N_31491,N_21152,N_25209);
and U31492 (N_31492,N_25648,N_25817);
nand U31493 (N_31493,N_28790,N_21494);
and U31494 (N_31494,N_26767,N_21844);
nand U31495 (N_31495,N_23589,N_24018);
and U31496 (N_31496,N_22109,N_20330);
or U31497 (N_31497,N_20627,N_25538);
and U31498 (N_31498,N_29591,N_23792);
nand U31499 (N_31499,N_25667,N_27503);
nand U31500 (N_31500,N_27710,N_21726);
xor U31501 (N_31501,N_26968,N_24887);
or U31502 (N_31502,N_24266,N_28253);
xnor U31503 (N_31503,N_27361,N_22399);
or U31504 (N_31504,N_23924,N_29853);
and U31505 (N_31505,N_28539,N_20518);
or U31506 (N_31506,N_20357,N_28077);
and U31507 (N_31507,N_27398,N_27919);
nand U31508 (N_31508,N_24160,N_29358);
and U31509 (N_31509,N_20002,N_25483);
nor U31510 (N_31510,N_24194,N_24942);
xnor U31511 (N_31511,N_28575,N_26103);
and U31512 (N_31512,N_29907,N_24685);
xnor U31513 (N_31513,N_28719,N_29153);
nor U31514 (N_31514,N_20370,N_24119);
and U31515 (N_31515,N_26717,N_28599);
or U31516 (N_31516,N_25319,N_24135);
nand U31517 (N_31517,N_27406,N_23753);
and U31518 (N_31518,N_27664,N_26438);
nor U31519 (N_31519,N_24052,N_25549);
nand U31520 (N_31520,N_21715,N_25881);
or U31521 (N_31521,N_21350,N_27192);
nor U31522 (N_31522,N_29097,N_22699);
and U31523 (N_31523,N_26134,N_20502);
or U31524 (N_31524,N_20170,N_24333);
nor U31525 (N_31525,N_28721,N_24321);
nor U31526 (N_31526,N_24642,N_23931);
and U31527 (N_31527,N_25514,N_26520);
nor U31528 (N_31528,N_24331,N_28602);
or U31529 (N_31529,N_28678,N_27025);
and U31530 (N_31530,N_28042,N_21097);
or U31531 (N_31531,N_28808,N_22705);
and U31532 (N_31532,N_27317,N_29898);
nor U31533 (N_31533,N_29053,N_24252);
and U31534 (N_31534,N_23280,N_27905);
or U31535 (N_31535,N_28760,N_27041);
or U31536 (N_31536,N_24453,N_28706);
nor U31537 (N_31537,N_27700,N_27620);
or U31538 (N_31538,N_20575,N_25536);
nor U31539 (N_31539,N_26564,N_25383);
nor U31540 (N_31540,N_20356,N_24370);
nand U31541 (N_31541,N_29939,N_29335);
nor U31542 (N_31542,N_24990,N_22025);
xor U31543 (N_31543,N_28319,N_25160);
or U31544 (N_31544,N_27602,N_22603);
nand U31545 (N_31545,N_22107,N_26771);
xor U31546 (N_31546,N_28135,N_24743);
and U31547 (N_31547,N_25942,N_20947);
nor U31548 (N_31548,N_27070,N_23750);
nand U31549 (N_31549,N_20165,N_26185);
nor U31550 (N_31550,N_26346,N_27312);
nor U31551 (N_31551,N_26935,N_23522);
and U31552 (N_31552,N_28052,N_29950);
or U31553 (N_31553,N_23922,N_20614);
and U31554 (N_31554,N_24546,N_21153);
nand U31555 (N_31555,N_28590,N_23336);
xor U31556 (N_31556,N_28119,N_29242);
xor U31557 (N_31557,N_29257,N_25167);
nor U31558 (N_31558,N_21983,N_21885);
nor U31559 (N_31559,N_22117,N_28347);
and U31560 (N_31560,N_24065,N_26160);
or U31561 (N_31561,N_25606,N_22885);
nor U31562 (N_31562,N_25812,N_23831);
nor U31563 (N_31563,N_25617,N_21026);
nor U31564 (N_31564,N_29846,N_21971);
or U31565 (N_31565,N_27833,N_22101);
or U31566 (N_31566,N_21862,N_23398);
xor U31567 (N_31567,N_29892,N_20084);
nor U31568 (N_31568,N_21992,N_29767);
and U31569 (N_31569,N_22401,N_25904);
nand U31570 (N_31570,N_28131,N_28967);
nor U31571 (N_31571,N_28673,N_27271);
or U31572 (N_31572,N_29443,N_25305);
and U31573 (N_31573,N_23291,N_29811);
xor U31574 (N_31574,N_25918,N_22073);
nand U31575 (N_31575,N_27252,N_20995);
and U31576 (N_31576,N_26794,N_27938);
nor U31577 (N_31577,N_27321,N_20032);
and U31578 (N_31578,N_26912,N_25944);
nand U31579 (N_31579,N_22042,N_22355);
xor U31580 (N_31580,N_23147,N_29679);
and U31581 (N_31581,N_24796,N_20542);
nor U31582 (N_31582,N_20158,N_26547);
xnor U31583 (N_31583,N_21580,N_21924);
nand U31584 (N_31584,N_28577,N_29332);
and U31585 (N_31585,N_24534,N_23727);
nand U31586 (N_31586,N_29988,N_26879);
and U31587 (N_31587,N_28798,N_24340);
nor U31588 (N_31588,N_23010,N_29012);
and U31589 (N_31589,N_20711,N_26408);
xor U31590 (N_31590,N_20799,N_23677);
or U31591 (N_31591,N_20527,N_24916);
and U31592 (N_31592,N_25003,N_24667);
or U31593 (N_31593,N_25759,N_26627);
and U31594 (N_31594,N_26820,N_20333);
nor U31595 (N_31595,N_26298,N_23524);
xnor U31596 (N_31596,N_25069,N_20108);
xnor U31597 (N_31597,N_27378,N_28143);
nand U31598 (N_31598,N_21087,N_25030);
and U31599 (N_31599,N_28580,N_26555);
xnor U31600 (N_31600,N_25334,N_26477);
nand U31601 (N_31601,N_26318,N_23402);
and U31602 (N_31602,N_25010,N_23328);
xor U31603 (N_31603,N_21199,N_24109);
and U31604 (N_31604,N_23095,N_26243);
nor U31605 (N_31605,N_24572,N_22671);
or U31606 (N_31606,N_28946,N_20896);
or U31607 (N_31607,N_26958,N_24265);
or U31608 (N_31608,N_28284,N_21413);
and U31609 (N_31609,N_27370,N_21403);
or U31610 (N_31610,N_29843,N_26822);
nand U31611 (N_31611,N_23508,N_22065);
or U31612 (N_31612,N_21171,N_26362);
nand U31613 (N_31613,N_27868,N_25037);
nor U31614 (N_31614,N_22009,N_26595);
nor U31615 (N_31615,N_28941,N_27509);
or U31616 (N_31616,N_24636,N_22277);
nand U31617 (N_31617,N_23789,N_23146);
nand U31618 (N_31618,N_20335,N_25029);
and U31619 (N_31619,N_21676,N_25229);
xnor U31620 (N_31620,N_23100,N_23743);
or U31621 (N_31621,N_23487,N_22684);
xor U31622 (N_31622,N_24733,N_21112);
and U31623 (N_31623,N_22811,N_23449);
nor U31624 (N_31624,N_22677,N_25530);
nor U31625 (N_31625,N_28997,N_20466);
and U31626 (N_31626,N_25015,N_22136);
or U31627 (N_31627,N_26736,N_23930);
nor U31628 (N_31628,N_28221,N_20180);
and U31629 (N_31629,N_29599,N_29354);
nand U31630 (N_31630,N_23295,N_24506);
nor U31631 (N_31631,N_28117,N_20433);
nor U31632 (N_31632,N_20997,N_23717);
and U31633 (N_31633,N_29984,N_24468);
nor U31634 (N_31634,N_21521,N_24499);
or U31635 (N_31635,N_25052,N_27732);
or U31636 (N_31636,N_28370,N_21964);
nor U31637 (N_31637,N_21405,N_25778);
or U31638 (N_31638,N_26711,N_26665);
nand U31639 (N_31639,N_21305,N_26831);
nor U31640 (N_31640,N_29404,N_29786);
and U31641 (N_31641,N_23646,N_29448);
or U31642 (N_31642,N_25341,N_26726);
or U31643 (N_31643,N_23839,N_24103);
or U31644 (N_31644,N_23499,N_28516);
or U31645 (N_31645,N_20156,N_26527);
nor U31646 (N_31646,N_27941,N_23976);
and U31647 (N_31647,N_29934,N_27984);
or U31648 (N_31648,N_27235,N_26285);
nor U31649 (N_31649,N_25809,N_26142);
and U31650 (N_31650,N_27877,N_22837);
or U31651 (N_31651,N_24031,N_27320);
nor U31652 (N_31652,N_24866,N_23247);
nand U31653 (N_31653,N_27126,N_20495);
nand U31654 (N_31654,N_22539,N_23412);
nor U31655 (N_31655,N_25973,N_27985);
nand U31656 (N_31656,N_29861,N_25891);
or U31657 (N_31657,N_29314,N_27476);
nor U31658 (N_31658,N_23675,N_28118);
nand U31659 (N_31659,N_21718,N_20727);
or U31660 (N_31660,N_28852,N_26333);
or U31661 (N_31661,N_26927,N_23836);
or U31662 (N_31662,N_28420,N_20907);
nand U31663 (N_31663,N_22801,N_21610);
or U31664 (N_31664,N_26848,N_23625);
and U31665 (N_31665,N_27243,N_23691);
nor U31666 (N_31666,N_25092,N_26323);
nor U31667 (N_31667,N_28758,N_28837);
xor U31668 (N_31668,N_21881,N_22517);
and U31669 (N_31669,N_21148,N_28054);
and U31670 (N_31670,N_20544,N_28214);
or U31671 (N_31671,N_23823,N_23298);
nand U31672 (N_31672,N_21060,N_25367);
nand U31673 (N_31673,N_28147,N_23462);
or U31674 (N_31674,N_23024,N_23018);
or U31675 (N_31675,N_21590,N_27846);
or U31676 (N_31676,N_20641,N_26352);
or U31677 (N_31677,N_26667,N_24658);
nand U31678 (N_31678,N_26844,N_28862);
nand U31679 (N_31679,N_20800,N_22740);
or U31680 (N_31680,N_26530,N_23241);
and U31681 (N_31681,N_22561,N_25751);
and U31682 (N_31682,N_25736,N_27815);
or U31683 (N_31683,N_24802,N_21562);
or U31684 (N_31684,N_29130,N_29152);
and U31685 (N_31685,N_25727,N_22872);
nor U31686 (N_31686,N_27267,N_27115);
nand U31687 (N_31687,N_29889,N_23330);
nand U31688 (N_31688,N_29686,N_26409);
xor U31689 (N_31689,N_27486,N_22111);
and U31690 (N_31690,N_22860,N_23386);
and U31691 (N_31691,N_27119,N_23392);
or U31692 (N_31692,N_29773,N_20712);
or U31693 (N_31693,N_27294,N_23209);
or U31694 (N_31694,N_24950,N_22600);
xnor U31695 (N_31695,N_27906,N_22515);
nor U31696 (N_31696,N_29866,N_25312);
and U31697 (N_31697,N_23376,N_27360);
nand U31698 (N_31698,N_26326,N_25692);
nor U31699 (N_31699,N_20666,N_23049);
nor U31700 (N_31700,N_28136,N_25316);
or U31701 (N_31701,N_27567,N_22813);
or U31702 (N_31702,N_27659,N_29835);
or U31703 (N_31703,N_27785,N_23798);
nor U31704 (N_31704,N_29868,N_22915);
and U31705 (N_31705,N_28035,N_28226);
and U31706 (N_31706,N_23414,N_23434);
and U31707 (N_31707,N_29979,N_22607);
or U31708 (N_31708,N_25121,N_22188);
and U31709 (N_31709,N_23954,N_21280);
nor U31710 (N_31710,N_25922,N_20744);
xnor U31711 (N_31711,N_24847,N_20579);
or U31712 (N_31712,N_25865,N_27072);
or U31713 (N_31713,N_21803,N_24917);
and U31714 (N_31714,N_25201,N_24456);
nand U31715 (N_31715,N_26054,N_21103);
xor U31716 (N_31716,N_28748,N_25804);
or U31717 (N_31717,N_26475,N_29757);
and U31718 (N_31718,N_23874,N_29920);
or U31719 (N_31719,N_28611,N_23644);
and U31720 (N_31720,N_21823,N_26437);
nor U31721 (N_31721,N_21745,N_27467);
nor U31722 (N_31722,N_29201,N_29870);
nand U31723 (N_31723,N_26150,N_20992);
or U31724 (N_31724,N_21685,N_26370);
and U31725 (N_31725,N_26553,N_26723);
and U31726 (N_31726,N_28196,N_28956);
and U31727 (N_31727,N_21531,N_29461);
or U31728 (N_31728,N_20760,N_26908);
or U31729 (N_31729,N_26714,N_20642);
and U31730 (N_31730,N_24131,N_23970);
xor U31731 (N_31731,N_26546,N_23413);
and U31732 (N_31732,N_27166,N_24332);
nor U31733 (N_31733,N_23813,N_29070);
or U31734 (N_31734,N_23164,N_26163);
or U31735 (N_31735,N_28455,N_27064);
xnor U31736 (N_31736,N_21545,N_26919);
nor U31737 (N_31737,N_27458,N_23668);
and U31738 (N_31738,N_27451,N_24735);
nor U31739 (N_31739,N_29025,N_23660);
nor U31740 (N_31740,N_24843,N_26621);
nor U31741 (N_31741,N_27698,N_24782);
nor U31742 (N_31742,N_21987,N_23702);
nor U31743 (N_31743,N_29409,N_20944);
nand U31744 (N_31744,N_27296,N_22514);
nand U31745 (N_31745,N_27750,N_23997);
or U31746 (N_31746,N_21345,N_27581);
nand U31747 (N_31747,N_29744,N_26276);
nand U31748 (N_31748,N_20147,N_29864);
or U31749 (N_31749,N_25406,N_25405);
nor U31750 (N_31750,N_23186,N_22438);
nand U31751 (N_31751,N_21385,N_27527);
xnor U31752 (N_31752,N_21340,N_29313);
nand U31753 (N_31753,N_26244,N_29220);
or U31754 (N_31754,N_28964,N_26581);
or U31755 (N_31755,N_29923,N_28156);
and U31756 (N_31756,N_28519,N_20097);
nand U31757 (N_31757,N_24812,N_29510);
nand U31758 (N_31758,N_25276,N_27387);
nor U31759 (N_31759,N_27045,N_20805);
nor U31760 (N_31760,N_27715,N_21565);
nor U31761 (N_31761,N_22729,N_25832);
and U31762 (N_31762,N_28637,N_24577);
and U31763 (N_31763,N_24067,N_20534);
nand U31764 (N_31764,N_20573,N_25495);
nand U31765 (N_31765,N_29445,N_22306);
nor U31766 (N_31766,N_26386,N_24897);
nand U31767 (N_31767,N_21732,N_23062);
nor U31768 (N_31768,N_26162,N_20836);
nor U31769 (N_31769,N_24375,N_24437);
or U31770 (N_31770,N_27512,N_22952);
xor U31771 (N_31771,N_23556,N_21999);
nand U31772 (N_31772,N_27078,N_23623);
nor U31773 (N_31773,N_29356,N_27279);
nor U31774 (N_31774,N_20018,N_28389);
nand U31775 (N_31775,N_21781,N_29583);
or U31776 (N_31776,N_29978,N_21995);
nand U31777 (N_31777,N_28272,N_28834);
nor U31778 (N_31778,N_28022,N_28969);
and U31779 (N_31779,N_28193,N_29559);
or U31780 (N_31780,N_21038,N_25837);
and U31781 (N_31781,N_24462,N_29859);
or U31782 (N_31782,N_21820,N_28179);
nor U31783 (N_31783,N_25645,N_23081);
xor U31784 (N_31784,N_22776,N_23310);
or U31785 (N_31785,N_26115,N_24047);
xor U31786 (N_31786,N_24170,N_29197);
xor U31787 (N_31787,N_23755,N_20709);
and U31788 (N_31788,N_20680,N_22380);
nor U31789 (N_31789,N_23626,N_24229);
and U31790 (N_31790,N_27102,N_26937);
or U31791 (N_31791,N_24310,N_29912);
or U31792 (N_31792,N_23605,N_26832);
and U31793 (N_31793,N_28173,N_20065);
nand U31794 (N_31794,N_22674,N_27326);
and U31795 (N_31795,N_20622,N_28186);
or U31796 (N_31796,N_25527,N_23197);
nor U31797 (N_31797,N_29074,N_21994);
or U31798 (N_31798,N_24153,N_21875);
and U31799 (N_31799,N_29612,N_29027);
xnor U31800 (N_31800,N_23778,N_21343);
or U31801 (N_31801,N_26532,N_26571);
nor U31802 (N_31802,N_25597,N_27297);
nor U31803 (N_31803,N_24010,N_29545);
xor U31804 (N_31804,N_23701,N_26072);
or U31805 (N_31805,N_24448,N_21480);
and U31806 (N_31806,N_28849,N_22697);
nor U31807 (N_31807,N_22258,N_20310);
and U31808 (N_31808,N_24383,N_28898);
nor U31809 (N_31809,N_23250,N_22861);
and U31810 (N_31810,N_27729,N_28091);
nand U31811 (N_31811,N_28104,N_23233);
or U31812 (N_31812,N_29916,N_23811);
nand U31813 (N_31813,N_27830,N_24022);
and U31814 (N_31814,N_28791,N_23419);
xnor U31815 (N_31815,N_26237,N_26644);
nand U31816 (N_31816,N_25593,N_26672);
nand U31817 (N_31817,N_25952,N_26458);
and U31818 (N_31818,N_25061,N_20728);
or U31819 (N_31819,N_24295,N_23210);
nor U31820 (N_31820,N_21362,N_21524);
or U31821 (N_31821,N_23086,N_25531);
nor U31822 (N_31822,N_20862,N_29932);
nand U31823 (N_31823,N_25261,N_26071);
and U31824 (N_31824,N_23465,N_27013);
nand U31825 (N_31825,N_24487,N_27674);
or U31826 (N_31826,N_20498,N_22192);
and U31827 (N_31827,N_28859,N_24638);
and U31828 (N_31828,N_26990,N_28068);
nor U31829 (N_31829,N_23917,N_29665);
and U31830 (N_31830,N_21490,N_25237);
nor U31831 (N_31831,N_20990,N_26918);
or U31832 (N_31832,N_26359,N_26283);
and U31833 (N_31833,N_24129,N_25279);
or U31834 (N_31834,N_27298,N_26626);
nor U31835 (N_31835,N_26784,N_28497);
nand U31836 (N_31836,N_20904,N_23736);
and U31837 (N_31837,N_21244,N_21500);
nor U31838 (N_31838,N_20736,N_27380);
or U31839 (N_31839,N_21516,N_26262);
xor U31840 (N_31840,N_22381,N_21542);
or U31841 (N_31841,N_22748,N_27228);
and U31842 (N_31842,N_22661,N_22406);
and U31843 (N_31843,N_23272,N_24326);
or U31844 (N_31844,N_21282,N_24196);
and U31845 (N_31845,N_24076,N_22932);
or U31846 (N_31846,N_20182,N_25869);
and U31847 (N_31847,N_26252,N_24971);
or U31848 (N_31848,N_27531,N_24704);
or U31849 (N_31849,N_27508,N_24012);
xnor U31850 (N_31850,N_28999,N_25479);
nand U31851 (N_31851,N_25857,N_25678);
or U31852 (N_31852,N_29783,N_21634);
nor U31853 (N_31853,N_28732,N_28875);
or U31854 (N_31854,N_22392,N_28546);
nor U31855 (N_31855,N_20279,N_23229);
nand U31856 (N_31856,N_26899,N_29212);
xor U31857 (N_31857,N_25927,N_28326);
nand U31858 (N_31858,N_28354,N_28248);
nand U31859 (N_31859,N_29336,N_28502);
and U31860 (N_31860,N_26172,N_27449);
nand U31861 (N_31861,N_24656,N_21320);
or U31862 (N_31862,N_28529,N_27225);
or U31863 (N_31863,N_23781,N_27660);
xnor U31864 (N_31864,N_21358,N_27879);
nor U31865 (N_31865,N_22685,N_20927);
nor U31866 (N_31866,N_21035,N_25292);
nand U31867 (N_31867,N_27840,N_24712);
nor U31868 (N_31868,N_22893,N_20926);
and U31869 (N_31869,N_28488,N_24397);
nor U31870 (N_31870,N_29037,N_24208);
nand U31871 (N_31871,N_29359,N_24253);
or U31872 (N_31872,N_21547,N_22660);
nor U31873 (N_31873,N_22079,N_28806);
xor U31874 (N_31874,N_27059,N_25789);
or U31875 (N_31875,N_27576,N_20776);
or U31876 (N_31876,N_28916,N_25102);
nor U31877 (N_31877,N_21398,N_22904);
nor U31878 (N_31878,N_26324,N_24650);
nor U31879 (N_31879,N_22572,N_29458);
and U31880 (N_31880,N_24949,N_27416);
or U31881 (N_31881,N_23360,N_22288);
and U31882 (N_31882,N_26099,N_28982);
and U31883 (N_31883,N_25493,N_24579);
or U31884 (N_31884,N_27967,N_26964);
nor U31885 (N_31885,N_20313,N_23816);
or U31886 (N_31886,N_24851,N_25438);
xnor U31887 (N_31887,N_23382,N_24096);
nor U31888 (N_31888,N_23175,N_24004);
or U31889 (N_31889,N_29051,N_26273);
nor U31890 (N_31890,N_26012,N_29975);
or U31891 (N_31891,N_29036,N_21333);
nor U31892 (N_31892,N_23818,N_22738);
nor U31893 (N_31893,N_23593,N_24415);
nor U31894 (N_31894,N_27908,N_29371);
nand U31895 (N_31895,N_29085,N_28534);
nand U31896 (N_31896,N_27603,N_21243);
or U31897 (N_31897,N_20792,N_26539);
nor U31898 (N_31898,N_23555,N_28297);
xor U31899 (N_31899,N_22386,N_24342);
or U31900 (N_31900,N_23326,N_24472);
and U31901 (N_31901,N_20958,N_28315);
and U31902 (N_31902,N_23334,N_28703);
and U31903 (N_31903,N_25006,N_27888);
or U31904 (N_31904,N_20366,N_21279);
nand U31905 (N_31905,N_22505,N_21857);
nand U31906 (N_31906,N_27667,N_24807);
nand U31907 (N_31907,N_21436,N_29263);
or U31908 (N_31908,N_22962,N_25180);
or U31909 (N_31909,N_26579,N_25428);
or U31910 (N_31910,N_25489,N_20034);
nand U31911 (N_31911,N_29604,N_26383);
nand U31912 (N_31912,N_27290,N_21240);
nor U31913 (N_31913,N_28211,N_26420);
or U31914 (N_31914,N_29746,N_26062);
nor U31915 (N_31915,N_25295,N_23552);
or U31916 (N_31916,N_25773,N_23290);
nor U31917 (N_31917,N_22969,N_20318);
nor U31918 (N_31918,N_20873,N_21074);
and U31919 (N_31919,N_27669,N_25264);
nand U31920 (N_31920,N_25109,N_20372);
and U31921 (N_31921,N_25640,N_23639);
nor U31922 (N_31922,N_24943,N_21077);
and U31923 (N_31923,N_25784,N_26036);
and U31924 (N_31924,N_22040,N_20112);
and U31925 (N_31925,N_22550,N_22792);
and U31926 (N_31926,N_26850,N_21075);
or U31927 (N_31927,N_23846,N_24800);
and U31928 (N_31928,N_25725,N_26166);
nand U31929 (N_31929,N_25210,N_26450);
xnor U31930 (N_31930,N_25662,N_27734);
or U31931 (N_31931,N_25095,N_22846);
and U31932 (N_31932,N_28733,N_23725);
nand U31933 (N_31933,N_26340,N_27240);
nor U31934 (N_31934,N_24282,N_28296);
or U31935 (N_31935,N_27069,N_22709);
and U31936 (N_31936,N_21967,N_23006);
nand U31937 (N_31937,N_26203,N_23227);
nor U31938 (N_31938,N_29077,N_25882);
nor U31939 (N_31939,N_29234,N_23391);
nand U31940 (N_31940,N_22876,N_23305);
and U31941 (N_31941,N_22919,N_20743);
and U31942 (N_31942,N_28302,N_23852);
and U31943 (N_31943,N_20808,N_29838);
xor U31944 (N_31944,N_25963,N_26921);
or U31945 (N_31945,N_29782,N_20567);
or U31946 (N_31946,N_28295,N_26801);
nand U31947 (N_31947,N_23506,N_29126);
or U31948 (N_31948,N_29536,N_22159);
or U31949 (N_31949,N_23945,N_25186);
and U31950 (N_31950,N_27731,N_24090);
nand U31951 (N_31951,N_20168,N_21783);
nand U31952 (N_31952,N_28681,N_20984);
xnor U31953 (N_31953,N_28317,N_27816);
nor U31954 (N_31954,N_26963,N_29585);
or U31955 (N_31955,N_28824,N_26861);
nand U31956 (N_31956,N_22950,N_21449);
nand U31957 (N_31957,N_28328,N_22894);
nand U31958 (N_31958,N_21041,N_29825);
or U31959 (N_31959,N_27538,N_23587);
and U31960 (N_31960,N_23535,N_24034);
nand U31961 (N_31961,N_27557,N_24043);
nor U31962 (N_31962,N_22092,N_26102);
nor U31963 (N_31963,N_26159,N_21157);
xor U31964 (N_31964,N_28170,N_23287);
nor U31965 (N_31965,N_24322,N_26397);
nand U31966 (N_31966,N_26896,N_28208);
nor U31967 (N_31967,N_27029,N_21608);
xnor U31968 (N_31968,N_20186,N_20331);
and U31969 (N_31969,N_25236,N_27641);
or U31970 (N_31970,N_28773,N_22047);
nand U31971 (N_31971,N_26929,N_27338);
and U31972 (N_31972,N_21373,N_21482);
and U31973 (N_31973,N_29918,N_26757);
and U31974 (N_31974,N_20519,N_28735);
nand U31975 (N_31975,N_26606,N_20242);
nor U31976 (N_31976,N_21033,N_24529);
nand U31977 (N_31977,N_27341,N_22363);
and U31978 (N_31978,N_29317,N_23857);
and U31979 (N_31979,N_28978,N_23208);
nor U31980 (N_31980,N_22271,N_26357);
nand U31981 (N_31981,N_25199,N_20791);
and U31982 (N_31982,N_29325,N_26211);
nand U31983 (N_31983,N_27649,N_24489);
and U31984 (N_31984,N_21454,N_24293);
nor U31985 (N_31985,N_29567,N_23825);
and U31986 (N_31986,N_23591,N_27521);
nor U31987 (N_31987,N_24759,N_24773);
nor U31988 (N_31988,N_27911,N_24817);
or U31989 (N_31989,N_26223,N_27625);
xor U31990 (N_31990,N_20793,N_28592);
nand U31991 (N_31991,N_23786,N_22842);
and U31992 (N_31992,N_28777,N_22579);
and U31993 (N_31993,N_25553,N_28375);
xor U31994 (N_31994,N_21576,N_23875);
or U31995 (N_31995,N_28002,N_26153);
and U31996 (N_31996,N_24806,N_29320);
nor U31997 (N_31997,N_20517,N_23401);
nand U31998 (N_31998,N_24746,N_25874);
and U31999 (N_31999,N_20881,N_26854);
nor U32000 (N_32000,N_22336,N_20685);
nor U32001 (N_32001,N_23084,N_20093);
and U32002 (N_32002,N_21618,N_25980);
or U32003 (N_32003,N_23154,N_21627);
nand U32004 (N_32004,N_22205,N_26497);
nor U32005 (N_32005,N_26827,N_21739);
nor U32006 (N_32006,N_27423,N_25695);
nand U32007 (N_32007,N_23450,N_21292);
nand U32008 (N_32008,N_23025,N_20831);
or U32009 (N_32009,N_24602,N_26272);
or U32010 (N_32010,N_23767,N_29319);
or U32011 (N_32011,N_22948,N_27804);
nand U32012 (N_32012,N_28094,N_23057);
and U32013 (N_32013,N_24432,N_26970);
nand U32014 (N_32014,N_27259,N_29065);
and U32015 (N_32015,N_24871,N_24292);
and U32016 (N_32016,N_25413,N_21615);
or U32017 (N_32017,N_26209,N_27947);
and U32018 (N_32018,N_28718,N_29160);
or U32019 (N_32019,N_27514,N_26375);
or U32020 (N_32020,N_28191,N_29793);
nand U32021 (N_32021,N_25938,N_21540);
nor U32022 (N_32022,N_24189,N_20286);
nand U32023 (N_32023,N_20014,N_22197);
xnor U32024 (N_32024,N_22652,N_26088);
nor U32025 (N_32025,N_20756,N_27281);
xnor U32026 (N_32026,N_23937,N_28168);
nor U32027 (N_32027,N_23090,N_22477);
or U32028 (N_32028,N_24454,N_20344);
nand U32029 (N_32029,N_26174,N_23143);
and U32030 (N_32030,N_23436,N_28582);
nor U32031 (N_32031,N_26892,N_28478);
nand U32032 (N_32032,N_25633,N_23124);
or U32033 (N_32033,N_24305,N_24496);
and U32034 (N_32034,N_25189,N_20307);
or U32035 (N_32035,N_25177,N_20464);
or U32036 (N_32036,N_24316,N_29982);
xnor U32037 (N_32037,N_28557,N_29937);
nor U32038 (N_32038,N_22255,N_21705);
nand U32039 (N_32039,N_21339,N_21203);
nand U32040 (N_32040,N_28108,N_23973);
or U32041 (N_32041,N_27990,N_24222);
and U32042 (N_32042,N_28228,N_24254);
xnor U32043 (N_32043,N_22020,N_20703);
and U32044 (N_32044,N_22864,N_27155);
nor U32045 (N_32045,N_27187,N_24840);
and U32046 (N_32046,N_27212,N_29936);
nor U32047 (N_32047,N_25327,N_20713);
and U32048 (N_32048,N_26059,N_21925);
xor U32049 (N_32049,N_25277,N_24398);
nand U32050 (N_32050,N_22395,N_28936);
nor U32051 (N_32051,N_20599,N_24994);
nand U32052 (N_32052,N_23120,N_26033);
or U32053 (N_32053,N_29684,N_22257);
or U32054 (N_32054,N_21533,N_23546);
or U32055 (N_32055,N_23486,N_20505);
and U32056 (N_32056,N_20875,N_27809);
nor U32057 (N_32057,N_28661,N_29742);
nor U32058 (N_32058,N_24879,N_26402);
nor U32059 (N_32059,N_25499,N_29178);
nand U32060 (N_32060,N_24914,N_26304);
nand U32061 (N_32061,N_23538,N_23977);
or U32062 (N_32062,N_26693,N_24576);
and U32063 (N_32063,N_29533,N_29103);
nand U32064 (N_32064,N_24597,N_23978);
nor U32065 (N_32065,N_22522,N_26215);
nor U32066 (N_32066,N_28841,N_25569);
or U32067 (N_32067,N_21577,N_21393);
nand U32068 (N_32068,N_28503,N_23960);
or U32069 (N_32069,N_27727,N_26390);
and U32070 (N_32070,N_28947,N_27612);
nor U32071 (N_32071,N_26307,N_24857);
and U32072 (N_32072,N_26198,N_21008);
or U32073 (N_32073,N_23729,N_25766);
nor U32074 (N_32074,N_29703,N_23230);
xnor U32075 (N_32075,N_24700,N_29865);
xor U32076 (N_32076,N_23364,N_24734);
nand U32077 (N_32077,N_26633,N_24061);
nand U32078 (N_32078,N_20595,N_26943);
or U32079 (N_32079,N_28369,N_22180);
nor U32080 (N_32080,N_28477,N_29423);
and U32081 (N_32081,N_24997,N_27272);
nand U32082 (N_32082,N_22518,N_24684);
xor U32083 (N_32083,N_29809,N_23666);
nor U32084 (N_32084,N_28576,N_27124);
nand U32085 (N_32085,N_28655,N_27210);
or U32086 (N_32086,N_24205,N_27206);
and U32087 (N_32087,N_28312,N_29175);
nor U32088 (N_32088,N_29523,N_20813);
xor U32089 (N_32089,N_27003,N_24720);
or U32090 (N_32090,N_22595,N_20187);
nand U32091 (N_32091,N_20693,N_29960);
or U32092 (N_32092,N_29243,N_26648);
xor U32093 (N_32093,N_28027,N_20445);
or U32094 (N_32094,N_20645,N_21263);
or U32095 (N_32095,N_26161,N_26371);
and U32096 (N_32096,N_25960,N_21657);
and U32097 (N_32097,N_29550,N_25631);
nor U32098 (N_32098,N_25562,N_27275);
and U32099 (N_32099,N_28148,N_24763);
and U32100 (N_32100,N_24068,N_24507);
xor U32101 (N_32101,N_23150,N_22693);
xnor U32102 (N_32102,N_25878,N_27270);
nor U32103 (N_32103,N_29718,N_27670);
and U32104 (N_32104,N_23116,N_26811);
and U32105 (N_32105,N_20049,N_29248);
and U32106 (N_32106,N_24764,N_27091);
or U32107 (N_32107,N_20038,N_28465);
nand U32108 (N_32108,N_25355,N_23088);
and U32109 (N_32109,N_26824,N_28129);
nand U32110 (N_32110,N_24089,N_22492);
or U32111 (N_32111,N_29396,N_29674);
nand U32112 (N_32112,N_21606,N_25737);
nand U32113 (N_32113,N_26584,N_23547);
or U32114 (N_32114,N_24445,N_29310);
or U32115 (N_32115,N_23301,N_20576);
nand U32116 (N_32116,N_23863,N_22099);
or U32117 (N_32117,N_20933,N_20463);
nor U32118 (N_32118,N_23151,N_27716);
nand U32119 (N_32119,N_21016,N_22302);
or U32120 (N_32120,N_26753,N_21777);
nor U32121 (N_32121,N_25854,N_29761);
or U32122 (N_32122,N_28781,N_22646);
or U32123 (N_32123,N_28366,N_23534);
nand U32124 (N_32124,N_25418,N_22372);
and U32125 (N_32125,N_26897,N_22275);
or U32126 (N_32126,N_20367,N_24268);
xnor U32127 (N_32127,N_27143,N_28797);
nor U32128 (N_32128,N_23794,N_28854);
or U32129 (N_32129,N_28904,N_25655);
xnor U32130 (N_32130,N_24080,N_27887);
nand U32131 (N_32131,N_29704,N_28351);
and U32132 (N_32132,N_28881,N_25349);
nand U32133 (N_32133,N_20639,N_20638);
nor U32134 (N_32134,N_24359,N_22072);
nor U32135 (N_32135,N_27996,N_28154);
and U32136 (N_32136,N_23511,N_20678);
and U32137 (N_32137,N_21076,N_24015);
nand U32138 (N_32138,N_25962,N_24614);
xnor U32139 (N_32139,N_26053,N_23125);
nand U32140 (N_32140,N_24530,N_22024);
xor U32141 (N_32141,N_24535,N_25704);
and U32142 (N_32142,N_29740,N_22021);
xnor U32143 (N_32143,N_27499,N_22407);
nor U32144 (N_32144,N_20472,N_25084);
or U32145 (N_32145,N_20577,N_29563);
or U32146 (N_32146,N_27261,N_20825);
nor U32147 (N_32147,N_20970,N_28498);
and U32148 (N_32148,N_21184,N_27635);
nand U32149 (N_32149,N_28258,N_20551);
and U32150 (N_32150,N_24180,N_28600);
and U32151 (N_32151,N_21910,N_21975);
nand U32152 (N_32152,N_28817,N_28343);
nand U32153 (N_32153,N_23074,N_29633);
or U32154 (N_32154,N_21487,N_29824);
nand U32155 (N_32155,N_24808,N_20151);
and U32156 (N_32156,N_23161,N_20943);
and U32157 (N_32157,N_29605,N_29532);
nor U32158 (N_32158,N_24624,N_21361);
and U32159 (N_32159,N_29083,N_25949);
and U32160 (N_32160,N_26601,N_22783);
or U32161 (N_32161,N_22800,N_29239);
xnor U32162 (N_32162,N_25971,N_24203);
nor U32163 (N_32163,N_25567,N_26007);
nor U32164 (N_32164,N_21304,N_21566);
or U32165 (N_32165,N_25860,N_28004);
and U32166 (N_32166,N_25028,N_20523);
nand U32167 (N_32167,N_24603,N_26018);
nor U32168 (N_32168,N_24077,N_24364);
or U32169 (N_32169,N_22910,N_29144);
nand U32170 (N_32170,N_20412,N_26452);
or U32171 (N_32171,N_27817,N_27258);
and U32172 (N_32172,N_26639,N_24434);
and U32173 (N_32173,N_24927,N_23567);
and U32174 (N_32174,N_22106,N_22597);
xor U32175 (N_32175,N_21006,N_21682);
nor U32176 (N_32176,N_25224,N_25760);
nor U32177 (N_32177,N_20291,N_20916);
or U32178 (N_32178,N_21326,N_21138);
nand U32179 (N_32179,N_27354,N_21549);
nor U32180 (N_32180,N_24063,N_21443);
and U32181 (N_32181,N_27619,N_25850);
or U32182 (N_32182,N_29850,N_29341);
nand U32183 (N_32183,N_23352,N_29020);
or U32184 (N_32184,N_28996,N_25463);
and U32185 (N_32185,N_28273,N_26941);
or U32186 (N_32186,N_27957,N_27890);
and U32187 (N_32187,N_21816,N_27781);
or U32188 (N_32188,N_21297,N_22041);
and U32189 (N_32189,N_22719,N_29032);
nor U32190 (N_32190,N_29405,N_26932);
nor U32191 (N_32191,N_27178,N_27033);
or U32192 (N_32192,N_24707,N_28716);
nand U32193 (N_32193,N_25993,N_21430);
or U32194 (N_32194,N_21370,N_28769);
nand U32195 (N_32195,N_21360,N_24839);
nand U32196 (N_32196,N_22095,N_25673);
nor U32197 (N_32197,N_26254,N_26056);
or U32198 (N_32198,N_23131,N_21965);
and U32199 (N_32199,N_20317,N_29615);
and U32200 (N_32200,N_27611,N_29259);
or U32201 (N_32201,N_25042,N_26222);
nor U32202 (N_32202,N_22343,N_23485);
or U32203 (N_32203,N_29116,N_20287);
and U32204 (N_32204,N_21433,N_21763);
nand U32205 (N_32205,N_28244,N_24754);
nor U32206 (N_32206,N_25426,N_25384);
nor U32207 (N_32207,N_23541,N_22945);
and U32208 (N_32208,N_24598,N_26454);
xnor U32209 (N_32209,N_27571,N_28008);
xor U32210 (N_32210,N_26513,N_21589);
and U32211 (N_32211,N_24102,N_22270);
and U32212 (N_32212,N_29389,N_27016);
or U32213 (N_32213,N_20303,N_28490);
nor U32214 (N_32214,N_23809,N_29177);
nand U32215 (N_32215,N_25214,N_29000);
nor U32216 (N_32216,N_24318,N_27424);
and U32217 (N_32217,N_20465,N_24404);
nand U32218 (N_32218,N_26998,N_29425);
and U32219 (N_32219,N_23256,N_23616);
or U32220 (N_32220,N_28868,N_21579);
nor U32221 (N_32221,N_21903,N_28172);
or U32222 (N_32222,N_24385,N_22879);
and U32223 (N_32223,N_23643,N_24485);
nand U32224 (N_32224,N_29447,N_25861);
or U32225 (N_32225,N_25813,N_20095);
nor U32226 (N_32226,N_25253,N_24745);
nor U32227 (N_32227,N_20903,N_26341);
or U32228 (N_32228,N_28821,N_29132);
nand U32229 (N_32229,N_22421,N_25043);
xnor U32230 (N_32230,N_27623,N_28980);
or U32231 (N_32231,N_27600,N_22718);
nor U32232 (N_32232,N_21100,N_28310);
or U32233 (N_32233,N_21765,N_22711);
xnor U32234 (N_32234,N_25579,N_25745);
and U32235 (N_32235,N_23338,N_28047);
and U32236 (N_32236,N_25577,N_29608);
nor U32237 (N_32237,N_22153,N_25130);
nor U32238 (N_32238,N_28177,N_28684);
and U32239 (N_32239,N_25983,N_27717);
and U32240 (N_32240,N_20142,N_22068);
or U32241 (N_32241,N_25572,N_24424);
or U32242 (N_32242,N_25459,N_20134);
and U32243 (N_32243,N_27793,N_20755);
nor U32244 (N_32244,N_21290,N_20092);
or U32245 (N_32245,N_27404,N_24860);
xor U32246 (N_32246,N_24555,N_23543);
or U32247 (N_32247,N_21347,N_26275);
and U32248 (N_32248,N_28710,N_29307);
nor U32249 (N_32249,N_23881,N_28096);
or U32250 (N_32250,N_22077,N_24567);
or U32251 (N_32251,N_28362,N_27244);
and U32252 (N_32252,N_27910,N_21972);
nand U32253 (N_32253,N_28869,N_29381);
or U32254 (N_32254,N_20246,N_24006);
nor U32255 (N_32255,N_25716,N_26118);
nor U32256 (N_32256,N_29638,N_27650);
and U32257 (N_32257,N_22486,N_24314);
nand U32258 (N_32258,N_29613,N_27482);
nand U32259 (N_32259,N_20898,N_28240);
nand U32260 (N_32260,N_24243,N_24822);
or U32261 (N_32261,N_28164,N_22976);
nand U32262 (N_32262,N_27127,N_20257);
nand U32263 (N_32263,N_20623,N_21104);
or U32264 (N_32264,N_25472,N_24106);
nand U32265 (N_32265,N_22934,N_22587);
and U32266 (N_32266,N_22647,N_23302);
and U32267 (N_32267,N_29279,N_25900);
and U32268 (N_32268,N_27598,N_20942);
nand U32269 (N_32269,N_25318,N_23882);
xnor U32270 (N_32270,N_29643,N_25041);
or U32271 (N_32271,N_29862,N_25395);
and U32272 (N_32272,N_21554,N_22730);
nor U32273 (N_32273,N_27616,N_20438);
nor U32274 (N_32274,N_25410,N_26445);
xnor U32275 (N_32275,N_28727,N_20227);
nor U32276 (N_32276,N_21365,N_27379);
or U32277 (N_32277,N_20149,N_29142);
and U32278 (N_32278,N_25409,N_25821);
nand U32279 (N_32279,N_28779,N_24981);
nand U32280 (N_32280,N_20397,N_21671);
nand U32281 (N_32281,N_23453,N_23265);
and U32282 (N_32282,N_29659,N_22571);
or U32283 (N_32283,N_25652,N_20848);
or U32284 (N_32284,N_21530,N_27624);
nor U32285 (N_32285,N_21250,N_29055);
nor U32286 (N_32286,N_26003,N_26725);
nand U32287 (N_32287,N_22405,N_28281);
and U32288 (N_32288,N_28339,N_27494);
nand U32289 (N_32289,N_22789,N_22624);
and U32290 (N_32290,N_28906,N_21697);
and U32291 (N_32291,N_24134,N_20690);
and U32292 (N_32292,N_26624,N_26876);
or U32293 (N_32293,N_23674,N_24378);
or U32294 (N_32294,N_29750,N_25222);
nand U32295 (N_32295,N_24421,N_20075);
and U32296 (N_32296,N_25826,N_29655);
nand U32297 (N_32297,N_26332,N_20354);
nand U32298 (N_32298,N_26574,N_21620);
xor U32299 (N_32299,N_22256,N_21703);
nor U32300 (N_32300,N_28883,N_20986);
nor U32301 (N_32301,N_26282,N_24380);
nand U32302 (N_32302,N_24585,N_23040);
and U32303 (N_32303,N_29565,N_27062);
nor U32304 (N_32304,N_27648,N_25691);
or U32305 (N_32305,N_24660,N_28405);
or U32306 (N_32306,N_26884,N_26043);
and U32307 (N_32307,N_28547,N_27203);
or U32308 (N_32308,N_27988,N_21093);
nor U32309 (N_32309,N_20668,N_26945);
nand U32310 (N_32310,N_26502,N_26894);
nand U32311 (N_32311,N_24861,N_26040);
and U32312 (N_32312,N_21123,N_23549);
or U32313 (N_32313,N_20321,N_27019);
nand U32314 (N_32314,N_27211,N_21397);
nor U32315 (N_32315,N_27510,N_23897);
or U32316 (N_32316,N_22165,N_28316);
or U32317 (N_32317,N_23669,N_20664);
nand U32318 (N_32318,N_24190,N_23205);
and U32319 (N_32319,N_23673,N_27333);
nor U32320 (N_32320,N_22389,N_20998);
nand U32321 (N_32321,N_25416,N_27337);
nor U32322 (N_32322,N_27111,N_25281);
or U32323 (N_32323,N_26325,N_25112);
or U32324 (N_32324,N_23676,N_24347);
or U32325 (N_32325,N_23996,N_24823);
nand U32326 (N_32326,N_24525,N_20312);
nand U32327 (N_32327,N_20013,N_25988);
or U32328 (N_32328,N_20560,N_24682);
or U32329 (N_32329,N_24596,N_24889);
nor U32330 (N_32330,N_22993,N_28263);
or U32331 (N_32331,N_22297,N_22992);
nor U32332 (N_32332,N_29113,N_25711);
nor U32333 (N_32333,N_22531,N_22843);
nand U32334 (N_32334,N_25958,N_25057);
nor U32335 (N_32335,N_21264,N_28629);
or U32336 (N_32336,N_24540,N_29400);
and U32337 (N_32337,N_22790,N_22683);
and U32338 (N_32338,N_22611,N_20381);
xnor U32339 (N_32339,N_22029,N_25872);
nor U32340 (N_32340,N_20362,N_21904);
nor U32341 (N_32341,N_27017,N_24335);
nand U32342 (N_32342,N_25297,N_26184);
and U32343 (N_32343,N_20129,N_23733);
nor U32344 (N_32344,N_27408,N_28633);
nand U32345 (N_32345,N_27738,N_24193);
nand U32346 (N_32346,N_24792,N_23876);
nand U32347 (N_32347,N_21181,N_23324);
nand U32348 (N_32348,N_25656,N_23892);
nor U32349 (N_32349,N_24864,N_24367);
nand U32350 (N_32350,N_22745,N_28830);
or U32351 (N_32351,N_22328,N_27403);
or U32352 (N_32352,N_25462,N_23769);
xnor U32353 (N_32353,N_26471,N_20962);
nand U32354 (N_32354,N_29531,N_25948);
and U32355 (N_32355,N_25302,N_26041);
and U32356 (N_32356,N_24752,N_27826);
nor U32357 (N_32357,N_21830,N_28270);
and U32358 (N_32358,N_20021,N_26435);
nand U32359 (N_32359,N_22376,N_26566);
and U32360 (N_32360,N_20384,N_26809);
and U32361 (N_32361,N_22339,N_28386);
nor U32362 (N_32362,N_22447,N_21518);
and U32363 (N_32363,N_26239,N_29139);
or U32364 (N_32364,N_29105,N_26114);
and U32365 (N_32365,N_21024,N_24821);
and U32366 (N_32366,N_28745,N_22639);
or U32367 (N_32367,N_24118,N_20479);
and U32368 (N_32368,N_26982,N_21134);
or U32369 (N_32369,N_21656,N_25206);
nor U32370 (N_32370,N_28994,N_22493);
nand U32371 (N_32371,N_22124,N_28198);
and U32372 (N_32372,N_28496,N_20209);
or U32373 (N_32373,N_28009,N_20388);
and U32374 (N_32374,N_20274,N_23557);
nor U32375 (N_32375,N_28504,N_27552);
nor U32376 (N_32376,N_27951,N_22717);
xnor U32377 (N_32377,N_25792,N_25957);
or U32378 (N_32378,N_25943,N_21124);
and U32379 (N_32379,N_22385,N_23166);
nand U32380 (N_32380,N_22653,N_24003);
and U32381 (N_32381,N_24662,N_25517);
and U32382 (N_32382,N_24391,N_23496);
nand U32383 (N_32383,N_25223,N_27712);
nand U32384 (N_32384,N_24392,N_20068);
nand U32385 (N_32385,N_21367,N_21498);
and U32386 (N_32386,N_29415,N_29721);
xor U32387 (N_32387,N_28957,N_24317);
and U32388 (N_32388,N_20763,N_28250);
or U32389 (N_32389,N_24071,N_29627);
nor U32390 (N_32390,N_22012,N_28815);
or U32391 (N_32391,N_29462,N_25239);
or U32392 (N_32392,N_22379,N_25637);
and U32393 (N_32393,N_20004,N_27488);
nand U32394 (N_32394,N_29312,N_27522);
nand U32395 (N_32395,N_26110,N_27662);
or U32396 (N_32396,N_25017,N_21641);
xor U32397 (N_32397,N_24091,N_29125);
nand U32398 (N_32398,N_26301,N_27592);
or U32399 (N_32399,N_21376,N_28765);
nor U32400 (N_32400,N_26473,N_26744);
nand U32401 (N_32401,N_26186,N_26345);
xor U32402 (N_32402,N_26769,N_26082);
and U32403 (N_32403,N_26221,N_25424);
or U32404 (N_32404,N_23035,N_21150);
and U32405 (N_32405,N_23489,N_23680);
or U32406 (N_32406,N_25726,N_22484);
or U32407 (N_32407,N_22474,N_24758);
or U32408 (N_32408,N_25219,N_22654);
and U32409 (N_32409,N_23259,N_24410);
nor U32410 (N_32410,N_20481,N_27446);
nand U32411 (N_32411,N_27568,N_21098);
and U32412 (N_32412,N_27042,N_24514);
or U32413 (N_32413,N_22506,N_23583);
or U32414 (N_32414,N_20750,N_23366);
nand U32415 (N_32415,N_26837,N_25351);
nand U32416 (N_32416,N_27350,N_25798);
xnor U32417 (N_32417,N_28728,N_24626);
or U32418 (N_32418,N_20340,N_24611);
or U32419 (N_32419,N_24788,N_29009);
nand U32420 (N_32420,N_21423,N_25542);
nand U32421 (N_32421,N_27543,N_20636);
nor U32422 (N_32422,N_24117,N_23586);
or U32423 (N_32423,N_26523,N_23829);
nand U32424 (N_32424,N_27125,N_20154);
and U32425 (N_32425,N_25769,N_23710);
and U32426 (N_32426,N_20159,N_20837);
nand U32427 (N_32427,N_26238,N_27464);
nor U32428 (N_32428,N_22361,N_28460);
xor U32429 (N_32429,N_24911,N_22905);
or U32430 (N_32430,N_20081,N_27950);
nor U32431 (N_32431,N_26339,N_27087);
and U32432 (N_32432,N_25111,N_26989);
or U32433 (N_32433,N_20795,N_21309);
or U32434 (N_32434,N_29303,N_20276);
and U32435 (N_32435,N_27726,N_26516);
and U32436 (N_32436,N_20057,N_24705);
nand U32437 (N_32437,N_27565,N_24450);
nor U32438 (N_32438,N_23317,N_26349);
and U32439 (N_32439,N_27129,N_28799);
nand U32440 (N_32440,N_22023,N_23572);
nand U32441 (N_32441,N_26952,N_21020);
nor U32442 (N_32442,N_27032,N_28795);
nor U32443 (N_32443,N_21241,N_20565);
nand U32444 (N_32444,N_27426,N_20768);
nand U32445 (N_32445,N_22696,N_28125);
nand U32446 (N_32446,N_29574,N_20905);
nor U32447 (N_32447,N_23715,N_29664);
and U32448 (N_32448,N_28241,N_23158);
or U32449 (N_32449,N_28630,N_24848);
xnor U32450 (N_32450,N_25011,N_24730);
or U32451 (N_32451,N_21425,N_27844);
nand U32452 (N_32452,N_26846,N_26604);
xnor U32453 (N_32453,N_21567,N_26609);
or U32454 (N_32454,N_21446,N_27049);
nor U32455 (N_32455,N_27128,N_22116);
nor U32456 (N_32456,N_20827,N_22441);
xnor U32457 (N_32457,N_21571,N_21344);
nor U32458 (N_32458,N_28874,N_28140);
nand U32459 (N_32459,N_22391,N_24171);
or U32460 (N_32460,N_29596,N_27544);
nor U32461 (N_32461,N_23182,N_22835);
nand U32462 (N_32462,N_21526,N_25859);
or U32463 (N_32463,N_27396,N_22470);
nor U32464 (N_32464,N_29528,N_21916);
or U32465 (N_32465,N_21646,N_26559);
xor U32466 (N_32466,N_20594,N_23853);
nand U32467 (N_32467,N_28827,N_24438);
nor U32468 (N_32468,N_20570,N_28243);
xor U32469 (N_32469,N_20529,N_28612);
and U32470 (N_32470,N_20452,N_25705);
or U32471 (N_32471,N_26207,N_22034);
or U32472 (N_32472,N_20547,N_23821);
nand U32473 (N_32473,N_29739,N_29454);
and U32474 (N_32474,N_21894,N_24361);
and U32475 (N_32475,N_28116,N_27968);
nand U32476 (N_32476,N_24123,N_28878);
nor U32477 (N_32477,N_24615,N_22712);
nand U32478 (N_32478,N_28419,N_24046);
nor U32479 (N_32479,N_28832,N_25985);
nor U32480 (N_32480,N_27589,N_25047);
nor U32481 (N_32481,N_27389,N_28382);
nor U32482 (N_32482,N_24116,N_25610);
or U32483 (N_32483,N_26774,N_20714);
or U32484 (N_32484,N_23399,N_23167);
nand U32485 (N_32485,N_25730,N_26538);
and U32486 (N_32486,N_26171,N_27020);
and U32487 (N_32487,N_24539,N_26253);
xor U32488 (N_32488,N_22769,N_29412);
nor U32489 (N_32489,N_23176,N_29927);
and U32490 (N_32490,N_26768,N_23196);
and U32491 (N_32491,N_24795,N_22315);
nand U32492 (N_32492,N_29489,N_27444);
or U32493 (N_32493,N_22971,N_27288);
nor U32494 (N_32494,N_25193,N_26046);
nand U32495 (N_32495,N_26424,N_22853);
nor U32496 (N_32496,N_25657,N_28061);
nand U32497 (N_32497,N_25772,N_28766);
nand U32498 (N_32498,N_26049,N_26628);
and U32499 (N_32499,N_25903,N_21167);
nor U32500 (N_32500,N_23606,N_20674);
nor U32501 (N_32501,N_28963,N_24505);
nand U32502 (N_32502,N_28261,N_26533);
and U32503 (N_32503,N_27071,N_24262);
nor U32504 (N_32504,N_26482,N_21119);
nor U32505 (N_32505,N_23093,N_21788);
and U32506 (N_32506,N_23393,N_29467);
nor U32507 (N_32507,N_28725,N_22320);
nor U32508 (N_32508,N_22283,N_23286);
nand U32509 (N_32509,N_26143,N_27104);
or U32510 (N_32510,N_25919,N_26065);
or U32511 (N_32511,N_28607,N_25961);
nand U32512 (N_32512,N_24956,N_21544);
or U32513 (N_32513,N_20954,N_22570);
or U32514 (N_32514,N_20176,N_29991);
and U32515 (N_32515,N_25475,N_22298);
nor U32516 (N_32516,N_27646,N_21334);
nor U32517 (N_32517,N_29854,N_24132);
xor U32518 (N_32518,N_29433,N_23238);
and U32519 (N_32519,N_20692,N_21348);
nor U32520 (N_32520,N_27097,N_26980);
and U32521 (N_32521,N_25825,N_22553);
nor U32522 (N_32522,N_22700,N_29261);
or U32523 (N_32523,N_23497,N_24826);
and U32524 (N_32524,N_21017,N_21899);
or U32525 (N_32525,N_24655,N_25266);
or U32526 (N_32526,N_22629,N_24155);
nor U32527 (N_32527,N_25758,N_21909);
nor U32528 (N_32528,N_27622,N_29140);
nand U32529 (N_32529,N_25385,N_27336);
or U32530 (N_32530,N_22161,N_20120);
nand U32531 (N_32531,N_20247,N_20850);
and U32532 (N_32532,N_23784,N_21426);
nand U32533 (N_32533,N_24377,N_22446);
nand U32534 (N_32534,N_29473,N_29286);
or U32535 (N_32535,N_25749,N_28772);
or U32536 (N_32536,N_23405,N_25481);
nand U32537 (N_32537,N_23192,N_20138);
or U32538 (N_32538,N_27526,N_29190);
nand U32539 (N_32539,N_22005,N_20485);
and U32540 (N_32540,N_23953,N_26797);
nor U32541 (N_32541,N_27057,N_24556);
xnor U32542 (N_32542,N_20041,N_22608);
nor U32543 (N_32543,N_27077,N_29504);
or U32544 (N_32544,N_24476,N_23369);
nor U32545 (N_32545,N_22110,N_21679);
and U32546 (N_32546,N_23492,N_21160);
xnor U32547 (N_32547,N_22787,N_22390);
xnor U32548 (N_32548,N_28268,N_20657);
nand U32549 (N_32549,N_21095,N_21451);
nor U32550 (N_32550,N_23723,N_27944);
nor U32551 (N_32551,N_26599,N_23046);
nand U32552 (N_32552,N_26289,N_25423);
nor U32553 (N_32553,N_28739,N_29534);
or U32554 (N_32554,N_23577,N_25071);
or U32555 (N_32555,N_21970,N_24072);
nand U32556 (N_32556,N_26394,N_26961);
nor U32557 (N_32557,N_23808,N_25103);
nor U32558 (N_32558,N_29090,N_24423);
nand U32559 (N_32559,N_23445,N_28842);
nor U32560 (N_32560,N_25715,N_22708);
nand U32561 (N_32561,N_23375,N_28065);
or U32562 (N_32562,N_21511,N_25732);
nand U32563 (N_32563,N_22886,N_23826);
xor U32564 (N_32564,N_27325,N_26529);
nor U32565 (N_32565,N_24809,N_20901);
nor U32566 (N_32566,N_23503,N_24697);
or U32567 (N_32567,N_26155,N_25068);
and U32568 (N_32568,N_25072,N_28409);
nand U32569 (N_32569,N_26060,N_28192);
xor U32570 (N_32570,N_27369,N_22329);
and U32571 (N_32571,N_27355,N_25834);
and U32572 (N_32572,N_20864,N_21311);
or U32573 (N_32573,N_27344,N_28668);
nand U32574 (N_32574,N_28320,N_21672);
xnor U32575 (N_32575,N_20699,N_25059);
or U32576 (N_32576,N_26416,N_21792);
and U32577 (N_32577,N_25062,N_22408);
and U32578 (N_32578,N_29847,N_23526);
and U32579 (N_32579,N_26456,N_24605);
nor U32580 (N_32580,N_22759,N_24928);
or U32581 (N_32581,N_24926,N_28385);
or U32582 (N_32582,N_21164,N_28017);
or U32583 (N_32583,N_27116,N_26451);
and U32584 (N_32584,N_25139,N_27961);
nand U32585 (N_32585,N_28225,N_25286);
nor U32586 (N_32586,N_27749,N_28062);
nand U32587 (N_32587,N_23528,N_23877);
nor U32588 (N_32588,N_22448,N_29805);
nand U32589 (N_32589,N_25849,N_25184);
nor U32590 (N_32590,N_27853,N_22764);
or U32591 (N_32591,N_26802,N_24483);
or U32592 (N_32592,N_23279,N_27175);
nor U32593 (N_32593,N_26819,N_29769);
nand U32594 (N_32594,N_29828,N_20538);
nor U32595 (N_32595,N_22841,N_26442);
nor U32596 (N_32596,N_25300,N_20185);
nor U32597 (N_32597,N_22982,N_22957);
nor U32598 (N_32598,N_26448,N_24987);
or U32599 (N_32599,N_24163,N_25607);
nor U32600 (N_32600,N_20189,N_28445);
nand U32601 (N_32601,N_21941,N_24972);
nor U32602 (N_32602,N_25117,N_25805);
or U32603 (N_32603,N_20630,N_23191);
nand U32604 (N_32604,N_23264,N_22332);
nand U32605 (N_32605,N_21655,N_21943);
or U32606 (N_32606,N_29930,N_29639);
nand U32607 (N_32607,N_21766,N_21226);
nor U32608 (N_32608,N_27721,N_20525);
nor U32609 (N_32609,N_24776,N_21497);
or U32610 (N_32610,N_20929,N_21266);
nor U32611 (N_32611,N_25885,N_20258);
nand U32612 (N_32612,N_21356,N_23292);
nor U32613 (N_32613,N_27688,N_23268);
and U32614 (N_32614,N_28227,N_22703);
nor U32615 (N_32615,N_24154,N_28736);
and U32616 (N_32616,N_22854,N_23934);
nor U32617 (N_32617,N_26480,N_26829);
or U32618 (N_32618,N_26887,N_25232);
and U32619 (N_32619,N_21229,N_27366);
nor U32620 (N_32620,N_21410,N_21213);
or U32621 (N_32621,N_20283,N_27035);
and U32622 (N_32622,N_22751,N_25836);
and U32623 (N_32623,N_27194,N_23878);
nand U32624 (N_32624,N_26038,N_20715);
nor U32625 (N_32625,N_22695,N_28656);
or U32626 (N_32626,N_28195,N_26335);
nor U32627 (N_32627,N_24698,N_20467);
nor U32628 (N_32628,N_28989,N_25939);
nand U32629 (N_32629,N_27435,N_27223);
nor U32630 (N_32630,N_22370,N_24670);
and U32631 (N_32631,N_20328,N_29791);
or U32632 (N_32632,N_25488,N_25051);
or U32633 (N_32633,N_26745,N_20351);
nor U32634 (N_32634,N_20346,N_27847);
nand U32635 (N_32635,N_28783,N_25328);
nor U32636 (N_32636,N_22191,N_28045);
and U32637 (N_32637,N_22066,N_26646);
nor U32638 (N_32638,N_20870,N_24829);
xnor U32639 (N_32639,N_21463,N_22822);
nand U32640 (N_32640,N_25194,N_24757);
or U32641 (N_32641,N_22424,N_25021);
xnor U32642 (N_32642,N_29732,N_21182);
or U32643 (N_32643,N_22528,N_26577);
nand U32644 (N_32644,N_22844,N_20949);
xnor U32645 (N_32645,N_21028,N_27702);
or U32646 (N_32646,N_25717,N_24651);
and U32647 (N_32647,N_20226,N_20417);
xor U32648 (N_32648,N_24108,N_29501);
or U32649 (N_32649,N_24202,N_25554);
xnor U32650 (N_32650,N_25603,N_28107);
and U32651 (N_32651,N_26279,N_26776);
and U32652 (N_32652,N_25829,N_28734);
and U32653 (N_32653,N_22771,N_23089);
or U32654 (N_32654,N_22895,N_27803);
nor U32655 (N_32655,N_21272,N_26368);
nand U32656 (N_32656,N_26130,N_20528);
nand U32657 (N_32657,N_27998,N_25271);
nor U32658 (N_32658,N_22168,N_23967);
nand U32659 (N_32659,N_28421,N_29505);
nand U32660 (N_32660,N_25621,N_28912);
and U32661 (N_32661,N_26891,N_29145);
nand U32662 (N_32662,N_24278,N_25125);
nor U32663 (N_32663,N_27894,N_22274);
nand U32664 (N_32664,N_23353,N_27655);
or U32665 (N_32665,N_24138,N_29634);
nand U32666 (N_32666,N_25689,N_21156);
nand U32667 (N_32667,N_26889,N_25001);
or U32668 (N_32668,N_28291,N_20902);
and U32669 (N_32669,N_23350,N_29999);
and U32670 (N_32670,N_29326,N_28866);
or U32671 (N_32671,N_25862,N_21378);
and U32672 (N_32672,N_29814,N_25190);
nor U32673 (N_32673,N_25034,N_23193);
nor U32674 (N_32674,N_20644,N_20473);
or U32675 (N_32675,N_27418,N_25391);
nor U32676 (N_32676,N_20436,N_24486);
nor U32677 (N_32677,N_25550,N_22557);
nand U32678 (N_32678,N_24659,N_24214);
and U32679 (N_32679,N_29609,N_22713);
xor U32680 (N_32680,N_24000,N_29071);
and U32681 (N_32681,N_24648,N_21535);
nor U32682 (N_32682,N_25185,N_20023);
nand U32683 (N_32683,N_27264,N_20492);
and U32684 (N_32684,N_26441,N_20928);
nor U32685 (N_32685,N_23832,N_26032);
nand U32686 (N_32686,N_22916,N_24345);
xor U32687 (N_32687,N_20961,N_23249);
nor U32688 (N_32688,N_27105,N_29736);
or U32689 (N_32689,N_25373,N_27918);
or U32690 (N_32690,N_29628,N_21687);
nand U32691 (N_32691,N_23764,N_20392);
and U32692 (N_32692,N_20588,N_20764);
and U32693 (N_32693,N_25710,N_29078);
xor U32694 (N_32694,N_29541,N_27138);
and U32695 (N_32695,N_25956,N_29488);
xnor U32696 (N_32696,N_24509,N_28222);
nor U32697 (N_32697,N_23838,N_23551);
or U32698 (N_32698,N_20983,N_21578);
or U32699 (N_32699,N_20245,N_28606);
xor U32700 (N_32700,N_20994,N_23728);
xor U32701 (N_32701,N_23461,N_20689);
nor U32702 (N_32702,N_21101,N_22053);
xnor U32703 (N_32703,N_25307,N_23758);
nor U32704 (N_32704,N_29924,N_23893);
nor U32705 (N_32705,N_27633,N_28811);
nor U32706 (N_32706,N_28437,N_20775);
nand U32707 (N_32707,N_26008,N_24313);
nor U32708 (N_32708,N_22423,N_29060);
or U32709 (N_32709,N_22637,N_28922);
nor U32710 (N_32710,N_26654,N_29165);
xor U32711 (N_32711,N_25966,N_27159);
or U32712 (N_32712,N_25372,N_24748);
nand U32713 (N_32713,N_22239,N_22088);
and U32714 (N_32714,N_27630,N_25670);
nand U32715 (N_32715,N_29503,N_29003);
nand U32716 (N_32716,N_21043,N_23900);
nor U32717 (N_32717,N_25598,N_21680);
nand U32718 (N_32718,N_20364,N_28039);
nor U32719 (N_32719,N_29996,N_24035);
nor U32720 (N_32720,N_26158,N_21131);
nand U32721 (N_32721,N_27836,N_26655);
nand U32722 (N_32722,N_25439,N_23705);
nand U32723 (N_32723,N_20399,N_27428);
or U32724 (N_32724,N_27390,N_28508);
nor U32725 (N_32725,N_26735,N_25897);
nor U32726 (N_32726,N_23377,N_29668);
nand U32727 (N_32727,N_29249,N_28283);
and U32728 (N_32728,N_29778,N_28555);
xnor U32729 (N_32729,N_27993,N_29876);
and U32730 (N_32730,N_29434,N_28275);
nand U32731 (N_32731,N_25587,N_22925);
or U32732 (N_32732,N_28426,N_26706);
nor U32733 (N_32733,N_24041,N_29225);
nor U32734 (N_32734,N_22524,N_27683);
or U32735 (N_32735,N_29873,N_23400);
nor U32736 (N_32736,N_22761,N_21725);
xor U32737 (N_32737,N_21001,N_25296);
nand U32738 (N_32738,N_20842,N_28643);
nand U32739 (N_32739,N_28865,N_21583);
nand U32740 (N_32740,N_27433,N_21824);
or U32741 (N_32741,N_21913,N_28252);
and U32742 (N_32742,N_20785,N_20934);
or U32743 (N_32743,N_27920,N_22093);
or U32744 (N_32744,N_29169,N_23258);
xor U32745 (N_32745,N_24898,N_23510);
nand U32746 (N_32746,N_20219,N_20911);
or U32747 (N_32747,N_22958,N_23519);
nand U32748 (N_32748,N_24127,N_26852);
nand U32749 (N_32749,N_24941,N_27881);
nand U32750 (N_32750,N_22358,N_29061);
nor U32751 (N_32751,N_28867,N_28966);
or U32752 (N_32752,N_22436,N_24177);
and U32753 (N_32753,N_23372,N_20771);
and U32754 (N_32754,N_28422,N_24965);
or U32755 (N_32755,N_26205,N_24750);
nand U32756 (N_32756,N_27085,N_23235);
xor U32757 (N_32757,N_29856,N_22612);
xor U32758 (N_32758,N_28141,N_29887);
and U32759 (N_32759,N_25091,N_21295);
or U32760 (N_32760,N_24811,N_23833);
or U32761 (N_32761,N_28699,N_23349);
and U32762 (N_32762,N_29199,N_21651);
nor U32763 (N_32763,N_26384,N_29789);
nand U32764 (N_32764,N_25182,N_20432);
nor U32765 (N_32765,N_26067,N_23180);
and U32766 (N_32766,N_27979,N_24330);
nand U32767 (N_32767,N_23356,N_24255);
xor U32768 (N_32768,N_23071,N_21481);
nor U32769 (N_32769,N_21380,N_21555);
nand U32770 (N_32770,N_22573,N_24288);
nand U32771 (N_32771,N_29562,N_26241);
and U32772 (N_32772,N_22248,N_26847);
nand U32773 (N_32773,N_21366,N_24363);
xor U32774 (N_32774,N_23617,N_29136);
xor U32775 (N_32775,N_28959,N_25936);
nor U32776 (N_32776,N_25917,N_22220);
or U32777 (N_32777,N_20471,N_26233);
and U32778 (N_32778,N_20293,N_20369);
nor U32779 (N_32779,N_21849,N_20080);
nor U32780 (N_32780,N_25013,N_26047);
nand U32781 (N_32781,N_26878,N_24545);
and U32782 (N_32782,N_22763,N_25188);
nand U32783 (N_32783,N_21957,N_23452);
nor U32784 (N_32784,N_24049,N_20334);
and U32785 (N_32785,N_27573,N_28891);
or U32786 (N_32786,N_27289,N_21915);
nor U32787 (N_32787,N_24279,N_23470);
nor U32788 (N_32788,N_29346,N_21281);
nand U32789 (N_32789,N_22887,N_27709);
nand U32790 (N_32790,N_25910,N_23956);
or U32791 (N_32791,N_29815,N_26509);
and U32792 (N_32792,N_22754,N_25951);
nand U32793 (N_32793,N_24023,N_22354);
nand U32794 (N_32794,N_25975,N_28847);
xor U32795 (N_32795,N_29391,N_22160);
and U32796 (N_32796,N_22353,N_27092);
or U32797 (N_32797,N_24066,N_20229);
xnor U32798 (N_32798,N_27786,N_20440);
nor U32799 (N_32799,N_23799,N_21258);
or U32800 (N_32800,N_21795,N_25415);
nor U32801 (N_32801,N_21200,N_28073);
xnor U32802 (N_32802,N_25212,N_28669);
or U32803 (N_32803,N_27965,N_28749);
or U32804 (N_32804,N_29657,N_23117);
and U32805 (N_32805,N_28740,N_27942);
or U32806 (N_32806,N_20040,N_23576);
nor U32807 (N_32807,N_25070,N_21708);
nand U32808 (N_32808,N_28280,N_23378);
nand U32809 (N_32809,N_22082,N_28462);
or U32810 (N_32810,N_29945,N_28338);
or U32811 (N_32811,N_23132,N_29881);
nor U32812 (N_32812,N_21855,N_24297);
and U32813 (N_32813,N_22516,N_24120);
nand U32814 (N_32814,N_22933,N_22975);
xor U32815 (N_32815,N_25515,N_29933);
and U32816 (N_32816,N_29138,N_25039);
nand U32817 (N_32817,N_23686,N_21919);
nand U32818 (N_32818,N_28756,N_27722);
and U32819 (N_32819,N_25840,N_21044);
nand U32820 (N_32820,N_28110,N_26353);
nand U32821 (N_32821,N_26113,N_26329);
or U32822 (N_32822,N_29506,N_27759);
nand U32823 (N_32823,N_24250,N_24081);
nand U32824 (N_32824,N_27220,N_25298);
xnor U32825 (N_32825,N_25020,N_27677);
nand U32826 (N_32826,N_20048,N_28694);
nor U32827 (N_32827,N_26881,N_26629);
nor U32828 (N_32828,N_21628,N_23333);
or U32829 (N_32829,N_23579,N_24665);
or U32830 (N_32830,N_26670,N_26988);
nor U32831 (N_32831,N_27917,N_27023);
nand U32832 (N_32832,N_28940,N_23418);
and U32833 (N_32833,N_26469,N_23431);
nand U32834 (N_32834,N_29299,N_29450);
xnor U32835 (N_32835,N_20861,N_27609);
nor U32836 (N_32836,N_28755,N_21723);
nand U32837 (N_32837,N_26534,N_20405);
and U32838 (N_32838,N_25464,N_25272);
xor U32839 (N_32839,N_24465,N_20483);
xnor U32840 (N_32840,N_22788,N_28246);
nand U32841 (N_32841,N_24550,N_20734);
nor U32842 (N_32842,N_21694,N_27986);
or U32843 (N_32843,N_29154,N_22201);
and U32844 (N_32844,N_28603,N_25858);
nor U32845 (N_32845,N_23957,N_24416);
nand U32846 (N_32846,N_28329,N_20581);
and U32847 (N_32847,N_25447,N_27676);
nand U32848 (N_32848,N_22828,N_25375);
and U32849 (N_32849,N_27399,N_20819);
and U32850 (N_32850,N_21140,N_29230);
nor U32851 (N_32851,N_24549,N_23341);
nand U32852 (N_32852,N_26141,N_23570);
xor U32853 (N_32853,N_21850,N_20846);
xnor U32854 (N_32854,N_29670,N_24093);
nor U32855 (N_32855,N_29680,N_22937);
or U32856 (N_32856,N_28901,N_22462);
nor U32857 (N_32857,N_23515,N_25998);
and U32858 (N_32858,N_22536,N_25414);
or U32859 (N_32859,N_24030,N_23156);
xnor U32860 (N_32860,N_25348,N_29277);
nor U32861 (N_32861,N_23170,N_26664);
nand U32862 (N_32862,N_29570,N_20078);
xor U32863 (N_32863,N_24148,N_28574);
nand U32864 (N_32864,N_27322,N_22425);
and U32865 (N_32865,N_23390,N_22757);
nor U32866 (N_32866,N_28278,N_22485);
nor U32867 (N_32867,N_21499,N_26079);
nand U32868 (N_32868,N_26915,N_29720);
nand U32869 (N_32869,N_26511,N_22791);
and U32870 (N_32870,N_28722,N_23293);
or U32871 (N_32871,N_23944,N_27960);
nand U32872 (N_32872,N_28203,N_27645);
xnor U32873 (N_32873,N_28157,N_29502);
nand U32874 (N_32874,N_23545,N_25735);
nand U32875 (N_32875,N_28396,N_28274);
and U32876 (N_32876,N_28885,N_22746);
or U32877 (N_32877,N_25991,N_29088);
nand U32878 (N_32878,N_26269,N_22690);
nand U32879 (N_32879,N_23633,N_21116);
nand U32880 (N_32880,N_21871,N_24521);
nor U32881 (N_32881,N_24263,N_22589);
and U32882 (N_32882,N_29370,N_24315);
nor U32883 (N_32883,N_29943,N_23278);
and U32884 (N_32884,N_25899,N_29880);
or U32885 (N_32885,N_24944,N_22548);
nand U32886 (N_32886,N_22613,N_28423);
and U32887 (N_32887,N_20396,N_28471);
or U32888 (N_32888,N_27183,N_23033);
or U32889 (N_32889,N_27250,N_24647);
nand U32890 (N_32890,N_29928,N_29059);
or U32891 (N_32891,N_21483,N_25455);
or U32892 (N_32892,N_26290,N_24863);
nand U32893 (N_32893,N_24100,N_21543);
nor U32894 (N_32894,N_23849,N_23936);
and U32895 (N_32895,N_20309,N_21669);
or U32896 (N_32896,N_23604,N_27257);
nor U32897 (N_32897,N_23243,N_29268);
nor U32898 (N_32898,N_24157,N_26985);
nand U32899 (N_32899,N_21245,N_29203);
xnor U32900 (N_32900,N_28475,N_29258);
nor U32901 (N_32901,N_22365,N_22212);
or U32902 (N_32902,N_29601,N_29521);
nor U32903 (N_32903,N_23898,N_26315);
nor U32904 (N_32904,N_29602,N_24368);
nand U32905 (N_32905,N_23031,N_26746);
and U32906 (N_32906,N_21774,N_20086);
nor U32907 (N_32907,N_20600,N_21141);
or U32908 (N_32908,N_20130,N_26608);
nor U32909 (N_32909,N_27546,N_20794);
nor U32910 (N_32910,N_24932,N_28636);
and U32911 (N_32911,N_27263,N_22630);
and U32912 (N_32912,N_24402,N_26652);
nand U32913 (N_32913,N_26816,N_27022);
or U32914 (N_32914,N_29554,N_26713);
nor U32915 (N_32915,N_26462,N_22627);
xor U32916 (N_32916,N_28363,N_22848);
nor U32917 (N_32917,N_29052,N_22226);
nand U32918 (N_32918,N_23408,N_21605);
or U32919 (N_32919,N_29852,N_26204);
nor U32920 (N_32920,N_21485,N_24695);
and U32921 (N_32921,N_21462,N_23696);
nor U32922 (N_32922,N_27148,N_28349);
and U32923 (N_32923,N_27897,N_21129);
nand U32924 (N_32924,N_20015,N_22491);
nand U32925 (N_32925,N_28774,N_24531);
or U32926 (N_32926,N_24429,N_27493);
or U32927 (N_32927,N_27661,N_27417);
nand U32928 (N_32928,N_26481,N_21613);
nor U32929 (N_32929,N_29878,N_29318);
nand U32930 (N_32930,N_24902,N_26754);
nand U32931 (N_32931,N_25659,N_28376);
or U32932 (N_32932,N_23129,N_21907);
xnor U32933 (N_32933,N_20359,N_20788);
nor U32934 (N_32934,N_28991,N_27971);
nand U32935 (N_32935,N_22552,N_29993);
xnor U32936 (N_32936,N_25614,N_28820);
and U32937 (N_32937,N_21691,N_28778);
and U32938 (N_32938,N_20824,N_20953);
nor U32939 (N_32939,N_21810,N_29855);
nand U32940 (N_32940,N_20478,N_28031);
nor U32941 (N_32941,N_27991,N_29216);
or U32942 (N_32942,N_22344,N_20157);
nand U32943 (N_32943,N_26740,N_29839);
or U32944 (N_32944,N_24488,N_26849);
and U32945 (N_32945,N_28818,N_25883);
and U32946 (N_32946,N_27812,N_29007);
and U32947 (N_32947,N_29929,N_20199);
xor U32948 (N_32948,N_23494,N_21616);
and U32949 (N_32949,N_29753,N_28853);
nand U32950 (N_32950,N_28015,N_28001);
nor U32951 (N_32951,N_22984,N_23908);
or U32952 (N_32952,N_25382,N_20886);
nor U32953 (N_32953,N_22786,N_28828);
or U32954 (N_32954,N_20610,N_20339);
nor U32955 (N_32955,N_26808,N_27668);
and U32956 (N_32956,N_25843,N_29874);
nor U32957 (N_32957,N_22590,N_20509);
nand U32958 (N_32958,N_28414,N_29376);
or U32959 (N_32959,N_23432,N_26803);
nor U32960 (N_32960,N_20302,N_25761);
nand U32961 (N_32961,N_20866,N_20385);
xnor U32962 (N_32962,N_26218,N_21237);
or U32963 (N_32963,N_27490,N_24816);
nor U32964 (N_32964,N_21158,N_28183);
nor U32965 (N_32965,N_28365,N_20550);
and U32966 (N_32966,N_20016,N_22543);
and U32967 (N_32967,N_26770,N_26793);
nand U32968 (N_32968,N_29998,N_24319);
xor U32969 (N_32969,N_25129,N_27051);
nand U32970 (N_32970,N_23483,N_22585);
and U32971 (N_32971,N_23683,N_28690);
nor U32972 (N_32972,N_26070,N_22468);
nand U32973 (N_32973,N_25965,N_27402);
or U32974 (N_32974,N_28166,N_20119);
xor U32975 (N_32975,N_25477,N_28353);
nor U32976 (N_32976,N_23061,N_23627);
or U32977 (N_32977,N_26570,N_29652);
nand U32978 (N_32978,N_25317,N_27382);
nor U32979 (N_32979,N_20618,N_26009);
xor U32980 (N_32980,N_24204,N_21581);
nand U32981 (N_32981,N_21707,N_27462);
and U32982 (N_32982,N_25050,N_25970);
or U32983 (N_32983,N_28204,N_29295);
nor U32984 (N_32984,N_24984,N_26974);
and U32985 (N_32985,N_25696,N_23609);
nand U32986 (N_32986,N_25240,N_23814);
or U32987 (N_32987,N_22071,N_27805);
nand U32988 (N_32988,N_28764,N_25174);
or U32989 (N_32989,N_25660,N_28913);
and U32990 (N_32990,N_23275,N_27854);
xnor U32991 (N_32991,N_27381,N_25974);
and U32992 (N_32992,N_20679,N_29580);
nand U32993 (N_32993,N_20952,N_24952);
and U32994 (N_32994,N_28860,N_28663);
nand U32995 (N_32995,N_23248,N_24382);
nor U32996 (N_32996,N_24466,N_29886);
nand U32997 (N_32997,N_23174,N_27843);
or U32998 (N_32998,N_20022,N_22476);
or U32999 (N_32999,N_24444,N_27909);
nor U33000 (N_33000,N_20195,N_29808);
or U33001 (N_33001,N_22455,N_27835);
xnor U33002 (N_33002,N_21155,N_22808);
and U33003 (N_33003,N_27489,N_23498);
or U33004 (N_33004,N_27708,N_26235);
or U33005 (N_33005,N_26560,N_24226);
and U33006 (N_33006,N_24417,N_28074);
xnor U33007 (N_33007,N_29393,N_20921);
and U33008 (N_33008,N_22562,N_29959);
and U33009 (N_33009,N_26662,N_26773);
or U33010 (N_33010,N_29394,N_24677);
nand U33011 (N_33011,N_24020,N_27760);
nor U33012 (N_33012,N_23345,N_28087);
nor U33013 (N_33013,N_20152,N_20982);
or U33014 (N_33014,N_26550,N_22825);
and U33015 (N_33015,N_25427,N_22182);
nor U33016 (N_33016,N_26213,N_25387);
and U33017 (N_33017,N_24563,N_20005);
xnor U33018 (N_33018,N_29300,N_28161);
and U33019 (N_33019,N_26649,N_21658);
nand U33020 (N_33020,N_24233,N_27764);
nand U33021 (N_33021,N_26048,N_25120);
xor U33022 (N_33022,N_27757,N_25740);
and U33023 (N_33023,N_24815,N_28081);
or U33024 (N_33024,N_21639,N_23236);
nor U33025 (N_33025,N_21400,N_24940);
nand U33026 (N_33026,N_25401,N_24630);
nor U33027 (N_33027,N_28845,N_29513);
nand U33028 (N_33028,N_29758,N_24737);
nor U33029 (N_33029,N_25278,N_23441);
nand U33030 (N_33030,N_22115,N_25846);
xnor U33031 (N_33031,N_22580,N_26657);
xor U33032 (N_33032,N_29651,N_27976);
nor U33033 (N_33033,N_20801,N_22659);
nand U33034 (N_33034,N_29672,N_22649);
nor U33035 (N_33035,N_27790,N_21050);
nand U33036 (N_33036,N_24353,N_29903);
or U33037 (N_33037,N_29422,N_25254);
or U33038 (N_33038,N_24606,N_27215);
and U33039 (N_33039,N_23512,N_28970);
and U33040 (N_33040,N_22251,N_27766);
nand U33041 (N_33041,N_26181,N_28693);
xor U33042 (N_33042,N_22918,N_28759);
nand U33043 (N_33043,N_25638,N_28064);
nand U33044 (N_33044,N_23096,N_26270);
or U33045 (N_33045,N_26228,N_23244);
nand U33046 (N_33046,N_20820,N_24586);
xor U33047 (N_33047,N_25454,N_21889);
and U33048 (N_33048,N_23135,N_22224);
nand U33049 (N_33049,N_22826,N_23307);
and U33050 (N_33050,N_27163,N_29921);
nor U33051 (N_33051,N_22911,N_24921);
nand U33052 (N_33052,N_25096,N_29594);
and U33053 (N_33053,N_23902,N_25016);
or U33054 (N_33054,N_29751,N_28237);
or U33055 (N_33055,N_28992,N_29911);
or U33056 (N_33056,N_25507,N_23998);
nor U33057 (N_33057,N_25218,N_22294);
nand U33058 (N_33058,N_20319,N_23207);
nor U33059 (N_33059,N_23271,N_24239);
or U33060 (N_33060,N_20584,N_21826);
nand U33061 (N_33061,N_24086,N_20106);
nor U33062 (N_33062,N_25156,N_22884);
nor U33063 (N_33063,N_29745,N_29526);
nand U33064 (N_33064,N_26651,N_24005);
nor U33065 (N_33065,N_24999,N_27169);
and U33066 (N_33066,N_29527,N_24629);
xor U33067 (N_33067,N_27977,N_26460);
nand U33068 (N_33068,N_22731,N_21778);
and U33069 (N_33069,N_22010,N_21408);
nor U33070 (N_33070,N_24681,N_21468);
nor U33071 (N_33071,N_20920,N_27696);
nand U33072 (N_33072,N_27966,N_22067);
and U33073 (N_33073,N_29432,N_23928);
or U33074 (N_33074,N_29524,N_23315);
nor U33075 (N_33075,N_22810,N_20730);
nand U33076 (N_33076,N_23242,N_28182);
nor U33077 (N_33077,N_22400,N_27487);
and U33078 (N_33078,N_20691,N_27096);
and U33079 (N_33079,N_21346,N_28314);
xnor U33080 (N_33080,N_26895,N_24595);
xor U33081 (N_33081,N_29180,N_20268);
nand U33082 (N_33082,N_20895,N_29568);
and U33083 (N_33083,N_25374,N_28543);
or U33084 (N_33084,N_23251,N_22437);
nand U33085 (N_33085,N_29748,N_22119);
nor U33086 (N_33086,N_21132,N_22882);
nand U33087 (N_33087,N_25777,N_26877);
nand U33088 (N_33088,N_25524,N_20987);
or U33089 (N_33089,N_20007,N_20640);
nand U33090 (N_33090,N_24575,N_24059);
nand U33091 (N_33091,N_24357,N_29357);
nand U33092 (N_33092,N_25196,N_25025);
nand U33093 (N_33093,N_21293,N_25161);
nand U33094 (N_33094,N_26543,N_26395);
xor U33095 (N_33095,N_29696,N_26780);
nor U33096 (N_33096,N_26182,N_24820);
nor U33097 (N_33097,N_28356,N_29191);
nand U33098 (N_33098,N_25799,N_24554);
xor U33099 (N_33099,N_29022,N_25893);
xor U33100 (N_33100,N_24755,N_24508);
xor U33101 (N_33101,N_26853,N_25580);
nand U33102 (N_33102,N_28631,N_29167);
nor U33103 (N_33103,N_20231,N_21747);
xnor U33104 (N_33104,N_21477,N_27832);
nor U33105 (N_33105,N_28918,N_29028);
xnor U33106 (N_33106,N_23042,N_26925);
and U33107 (N_33107,N_23152,N_27391);
nand U33108 (N_33108,N_25093,N_29644);
nand U33109 (N_33109,N_27221,N_22744);
xnor U33110 (N_33110,N_25806,N_28150);
nor U33111 (N_33111,N_22260,N_26705);
xor U33112 (N_33112,N_20484,N_28597);
nand U33113 (N_33113,N_24872,N_25364);
nand U33114 (N_33114,N_24107,N_26265);
nor U33115 (N_33115,N_29820,N_28624);
nand U33116 (N_33116,N_27373,N_28591);
nor U33117 (N_33117,N_24350,N_20480);
or U33118 (N_33118,N_26616,N_24878);
or U33119 (N_33119,N_20700,N_21832);
or U33120 (N_33120,N_28536,N_24358);
nand U33121 (N_33121,N_27266,N_29831);
and U33122 (N_33122,N_25116,N_29173);
nor U33123 (N_33123,N_23779,N_29211);
and U33124 (N_33124,N_27705,N_24661);
and U33125 (N_33125,N_24825,N_26109);
or U33126 (N_33126,N_27654,N_21591);
or U33127 (N_33127,N_24435,N_25309);
nand U33128 (N_33128,N_24053,N_22535);
or U33129 (N_33129,N_29120,N_22158);
nand U33130 (N_33130,N_22672,N_29650);
xnor U33131 (N_33131,N_27248,N_25476);
nand U33132 (N_33132,N_22190,N_28753);
or U33133 (N_33133,N_29002,N_27309);
nand U33134 (N_33134,N_26055,N_29858);
nand U33135 (N_33135,N_26170,N_24344);
nor U33136 (N_33136,N_28738,N_26956);
or U33137 (N_33137,N_28492,N_25722);
xnor U33138 (N_33138,N_25539,N_29322);
and U33139 (N_33139,N_20223,N_23285);
and U33140 (N_33140,N_20515,N_23051);
and U33141 (N_33141,N_28893,N_25419);
or U33142 (N_33142,N_25794,N_22634);
and U33143 (N_33143,N_20428,N_28388);
nor U33144 (N_33144,N_20981,N_21741);
and U33145 (N_33145,N_20039,N_23759);
nor U33146 (N_33146,N_23559,N_28145);
xnor U33147 (N_33147,N_25999,N_21285);
or U33148 (N_33148,N_20957,N_27420);
nor U33149 (N_33149,N_22644,N_23344);
or U33150 (N_33150,N_25402,N_27554);
nor U33151 (N_33151,N_23791,N_27315);
nor U33152 (N_33152,N_20179,N_22223);
or U33153 (N_33153,N_27913,N_23594);
and U33154 (N_33154,N_25336,N_27656);
nand U33155 (N_33155,N_28100,N_27651);
nand U33156 (N_33156,N_28499,N_25818);
or U33157 (N_33157,N_23600,N_21071);
and U33158 (N_33158,N_21860,N_24870);
and U33159 (N_33159,N_22636,N_27479);
nor U33160 (N_33160,N_22322,N_21584);
nor U33161 (N_33161,N_26277,N_24604);
and U33162 (N_33162,N_22901,N_23550);
or U33163 (N_33163,N_23219,N_21867);
or U33164 (N_33164,N_22927,N_28013);
nor U33165 (N_33165,N_28804,N_28807);
or U33166 (N_33166,N_20213,N_21084);
or U33167 (N_33167,N_23879,N_25707);
nor U33168 (N_33168,N_25545,N_25616);
and U33169 (N_33169,N_25684,N_27492);
and U33170 (N_33170,N_28647,N_24710);
xor U33171 (N_33171,N_27306,N_20055);
or U33172 (N_33172,N_27872,N_26782);
or U33173 (N_33173,N_21737,N_23222);
nand U33174 (N_33174,N_25412,N_28542);
nand U33175 (N_33175,N_26104,N_29584);
or U33176 (N_33176,N_22411,N_20009);
nor U33177 (N_33177,N_23019,N_21755);
nand U33178 (N_33178,N_23883,N_26975);
nand U33179 (N_33179,N_20275,N_27590);
nand U33180 (N_33180,N_29086,N_27122);
nand U33181 (N_33181,N_24218,N_22986);
and U33182 (N_33182,N_27818,N_20164);
or U33183 (N_33183,N_20779,N_25151);
nand U33184 (N_33184,N_28762,N_26376);
or U33185 (N_33185,N_27513,N_26267);
and U33186 (N_33186,N_25080,N_25596);
or U33187 (N_33187,N_25941,N_21642);
xor U33188 (N_33188,N_23319,N_24880);
or U33189 (N_33189,N_29349,N_27368);
and U33190 (N_33190,N_29917,N_29515);
nand U33191 (N_33191,N_26123,N_24248);
nor U33192 (N_33192,N_28220,N_28742);
and U33193 (N_33193,N_21840,N_25618);
nand U33194 (N_33194,N_29759,N_26860);
and U33195 (N_33195,N_23474,N_20325);
and U33196 (N_33196,N_27345,N_26939);
nor U33197 (N_33197,N_21352,N_23822);
or U33198 (N_33198,N_28344,N_23754);
or U33199 (N_33199,N_21089,N_29023);
or U33200 (N_33200,N_29544,N_27427);
or U33201 (N_33201,N_28473,N_24862);
and U33202 (N_33202,N_20913,N_27285);
or U33203 (N_33203,N_25586,N_21382);
and U33204 (N_33204,N_24504,N_27293);
nand U33205 (N_33205,N_24805,N_25396);
nand U33206 (N_33206,N_29700,N_23843);
or U33207 (N_33207,N_20285,N_26587);
xnor U33208 (N_33208,N_22413,N_20696);
or U33209 (N_33209,N_26678,N_25494);
nor U33210 (N_33210,N_21529,N_23974);
nand U33211 (N_33211,N_20254,N_24409);
nor U33212 (N_33212,N_26393,N_26015);
xnor U33213 (N_33213,N_20856,N_27637);
nor U33214 (N_33214,N_25498,N_21125);
nand U33215 (N_33215,N_20206,N_23580);
xnor U33216 (N_33216,N_21686,N_23389);
and U33217 (N_33217,N_20818,N_24051);
nand U33218 (N_33218,N_29566,N_21937);
xor U33219 (N_33219,N_21504,N_28986);
nor U33220 (N_33220,N_22529,N_25274);
nand U33221 (N_33221,N_21743,N_27008);
xnor U33222 (N_33222,N_26487,N_27287);
and U33223 (N_33223,N_27302,N_28950);
and U33224 (N_33224,N_22549,N_26779);
and U33225 (N_33225,N_20626,N_28224);
or U33226 (N_33226,N_24753,N_22125);
xnor U33227 (N_33227,N_28726,N_29149);
xor U33228 (N_33228,N_26446,N_26922);
or U33229 (N_33229,N_29006,N_21259);
nand U33230 (N_33230,N_20767,N_21701);
nor U33231 (N_33231,N_27330,N_28704);
and U33232 (N_33232,N_23719,N_28708);
and U33233 (N_33233,N_29788,N_22998);
xor U33234 (N_33234,N_24420,N_24868);
or U33235 (N_33235,N_26331,N_29869);
or U33236 (N_33236,N_26425,N_25879);
xor U33237 (N_33237,N_27123,N_29787);
or U33238 (N_33238,N_28563,N_28348);
and U33239 (N_33239,N_22544,N_20733);
and U33240 (N_33240,N_26069,N_20930);
or U33241 (N_33241,N_24664,N_24303);
xnor U33242 (N_33242,N_26080,N_21946);
or U33243 (N_33243,N_21890,N_22286);
nand U33244 (N_33244,N_24767,N_25643);
nor U33245 (N_33245,N_21948,N_22839);
nand U33246 (N_33246,N_27780,N_29611);
nand U33247 (N_33247,N_23539,N_23700);
nand U33248 (N_33248,N_29715,N_28911);
nor U33249 (N_33249,N_23013,N_26157);
nand U33250 (N_33250,N_28480,N_25984);
nand U33251 (N_33251,N_20012,N_26495);
or U33252 (N_33252,N_24907,N_20695);
nor U33253 (N_33253,N_21688,N_24037);
or U33254 (N_33254,N_27601,N_24644);
nor U33255 (N_33255,N_26229,N_22105);
xor U33256 (N_33256,N_24623,N_22805);
nand U33257 (N_33257,N_22169,N_29213);
xor U33258 (N_33258,N_26227,N_21509);
nand U33259 (N_33259,N_23695,N_22227);
nor U33260 (N_33260,N_23312,N_21363);
or U33261 (N_33261,N_22616,N_23022);
nor U33262 (N_33262,N_23714,N_29084);
and U33263 (N_33263,N_22167,N_22085);
nand U33264 (N_33264,N_28948,N_25533);
nand U33265 (N_33265,N_26686,N_29366);
or U33266 (N_33266,N_23212,N_24569);
nand U33267 (N_33267,N_29439,N_25771);
nor U33268 (N_33268,N_27089,N_27328);
nand U33269 (N_33269,N_28971,N_20421);
and U33270 (N_33270,N_28491,N_27823);
nor U33271 (N_33271,N_24125,N_29076);
nor U33272 (N_33272,N_21829,N_24447);
or U33273 (N_33273,N_25511,N_20620);
or U33274 (N_33274,N_20398,N_28032);
and U33275 (N_33275,N_22086,N_24935);
and U33276 (N_33276,N_26051,N_28505);
and U33277 (N_33277,N_28586,N_23596);
nand U33278 (N_33278,N_25543,N_21120);
nor U33279 (N_33279,N_24457,N_22556);
or U33280 (N_33280,N_24512,N_25811);
xnor U33281 (N_33281,N_24286,N_24403);
and U33282 (N_33282,N_27614,N_25200);
and U33283 (N_33283,N_26403,N_29623);
and U33284 (N_33284,N_28932,N_24588);
xor U33285 (N_33285,N_26817,N_20612);
nand U33286 (N_33286,N_23613,N_21962);
nor U33287 (N_33287,N_28084,N_26552);
nand U33288 (N_33288,N_25911,N_22809);
and U33289 (N_33289,N_24813,N_28731);
nand U33290 (N_33290,N_24062,N_26292);
nor U33291 (N_33291,N_24797,N_24970);
nand U33292 (N_33292,N_26092,N_27558);
nand U33293 (N_33293,N_21107,N_22679);
or U33294 (N_33294,N_23873,N_22131);
or U33295 (N_33295,N_23706,N_24179);
and U33296 (N_33296,N_27447,N_24772);
nand U33297 (N_33297,N_27331,N_24836);
nor U33298 (N_33298,N_28550,N_22856);
or U33299 (N_33299,N_29496,N_21870);
nor U33300 (N_33300,N_21768,N_20704);
nand U33301 (N_33301,N_24855,N_22225);
nor U33302 (N_33302,N_22127,N_24674);
and U33303 (N_33303,N_23866,N_26517);
and U33304 (N_33304,N_23130,N_25204);
nand U33305 (N_33305,N_24064,N_22896);
or U33306 (N_33306,N_20804,N_23313);
nor U33307 (N_33307,N_23542,N_27580);
or U33308 (N_33308,N_23108,N_25408);
xnor U33309 (N_33309,N_21205,N_24111);
nand U33310 (N_33310,N_27893,N_25087);
and U33311 (N_33311,N_20847,N_23263);
nand U33312 (N_33312,N_24589,N_25055);
xnor U33313 (N_33313,N_28285,N_20201);
nand U33314 (N_33314,N_23325,N_21288);
nand U33315 (N_33315,N_25131,N_29830);
nand U33316 (N_33316,N_22873,N_21836);
nor U33317 (N_33317,N_25267,N_20085);
nor U33318 (N_33318,N_24373,N_22594);
xnor U33319 (N_33319,N_28043,N_20977);
xnor U33320 (N_33320,N_21396,N_20797);
nor U33321 (N_33321,N_20069,N_28201);
xnor U33322 (N_33322,N_21764,N_28558);
nor U33323 (N_33323,N_23907,N_21985);
nand U33324 (N_33324,N_20448,N_26014);
or U33325 (N_33325,N_24372,N_27561);
and U33326 (N_33326,N_20072,N_23199);
nand U33327 (N_33327,N_25690,N_20821);
or U33328 (N_33328,N_20248,N_22368);
nand U33329 (N_33329,N_27607,N_21631);
xnor U33330 (N_33330,N_27455,N_22006);
nor U33331 (N_33331,N_24966,N_21508);
nor U33332 (N_33332,N_24379,N_28819);
or U33333 (N_33333,N_22997,N_22341);
or U33334 (N_33334,N_20375,N_28829);
and U33335 (N_33335,N_21761,N_22489);
nand U33336 (N_33336,N_21668,N_28332);
xor U33337 (N_33337,N_28299,N_28889);
nand U33338 (N_33338,N_28938,N_26418);
nand U33339 (N_33339,N_24977,N_25641);
or U33340 (N_33340,N_25492,N_21128);
nor U33341 (N_33341,N_27827,N_20019);
or U33342 (N_33342,N_29174,N_21230);
nor U33343 (N_33343,N_27324,N_26440);
nand U33344 (N_33344,N_25920,N_25487);
xnor U33345 (N_33345,N_26119,N_21750);
nor U33346 (N_33346,N_25150,N_28425);
nand U33347 (N_33347,N_22716,N_24199);
and U33348 (N_33348,N_20294,N_28835);
xnor U33349 (N_33349,N_21144,N_27849);
and U33350 (N_33350,N_21938,N_22356);
nand U33351 (N_33351,N_22635,N_25157);
or U33352 (N_33352,N_29334,N_28594);
xnor U33353 (N_33353,N_29497,N_23351);
nor U33354 (N_33354,N_20056,N_29888);
or U33355 (N_33355,N_22768,N_26828);
nor U33356 (N_33356,N_23162,N_29361);
nor U33357 (N_33357,N_29466,N_27765);
xor U33358 (N_33358,N_26347,N_25864);
or U33359 (N_33359,N_26630,N_29426);
and U33360 (N_33360,N_24366,N_27692);
and U33361 (N_33361,N_29964,N_23443);
and U33362 (N_33362,N_28642,N_25315);
nor U33363 (N_33363,N_21939,N_23553);
or U33364 (N_33364,N_21877,N_25259);
nand U33365 (N_33365,N_27963,N_29362);
and U33366 (N_33366,N_24714,N_21221);
nor U33367 (N_33367,N_25354,N_21086);
nand U33368 (N_33368,N_25523,N_25978);
xnor U33369 (N_33369,N_24172,N_27440);
or U33370 (N_33370,N_25924,N_24547);
nand U33371 (N_33371,N_24275,N_27283);
or U33372 (N_33372,N_28568,N_29363);
nand U33373 (N_33373,N_21314,N_21471);
or U33374 (N_33374,N_22906,N_29671);
and U33375 (N_33375,N_22189,N_22545);
xnor U33376 (N_33376,N_25895,N_20001);
xnor U33377 (N_33377,N_24883,N_23632);
or U33378 (N_33378,N_26992,N_26180);
nor U33379 (N_33379,N_29977,N_24854);
nor U33380 (N_33380,N_25123,N_28919);
and U33381 (N_33381,N_21808,N_23554);
xor U33382 (N_33382,N_27882,N_25743);
nor U33383 (N_33383,N_20003,N_23007);
or U33384 (N_33384,N_25411,N_22495);
and U33385 (N_33385,N_22604,N_25664);
and U33386 (N_33386,N_29046,N_26025);
or U33387 (N_33387,N_22214,N_22875);
nand U33388 (N_33388,N_22114,N_28016);
nand U33389 (N_33389,N_22004,N_29713);
nor U33390 (N_33390,N_22970,N_29347);
nor U33391 (N_33391,N_23636,N_28962);
xnor U33392 (N_33392,N_21447,N_22501);
and U33393 (N_33393,N_24779,N_26597);
or U33394 (N_33394,N_23894,N_27801);
nand U33395 (N_33395,N_21742,N_23664);
and U33396 (N_33396,N_27584,N_23713);
nor U33397 (N_33397,N_24101,N_21717);
nor U33398 (N_33398,N_26001,N_20533);
or U33399 (N_33399,N_21592,N_28524);
nor U33400 (N_33400,N_29338,N_22619);
and U33401 (N_33401,N_26583,N_27778);
and U33402 (N_33402,N_24600,N_22990);
or U33403 (N_33403,N_22393,N_28610);
xnor U33404 (N_33404,N_26125,N_27763);
xor U33405 (N_33405,N_25929,N_28942);
nand U33406 (N_33406,N_22324,N_27883);
xor U33407 (N_33407,N_20091,N_20815);
and U33408 (N_33408,N_20222,N_27117);
and U33409 (N_33409,N_26430,N_23225);
nor U33410 (N_33410,N_24838,N_22080);
nand U33411 (N_33411,N_27170,N_24289);
xor U33412 (N_33412,N_21096,N_22890);
and U33413 (N_33413,N_20099,N_23518);
nor U33414 (N_33414,N_29579,N_20221);
or U33415 (N_33415,N_21216,N_25699);
nor U33416 (N_33416,N_21882,N_21173);
nand U33417 (N_33417,N_24381,N_22307);
and U33418 (N_33418,N_29162,N_22720);
and U33419 (N_33419,N_29297,N_22179);
or U33420 (N_33420,N_22964,N_22620);
or U33421 (N_33421,N_28451,N_28822);
nor U33422 (N_33422,N_23216,N_26951);
and U33423 (N_33423,N_21188,N_28289);
or U33424 (N_33424,N_26485,N_22187);
nor U33425 (N_33425,N_25583,N_20721);
and U33426 (N_33426,N_24084,N_28570);
nor U33427 (N_33427,N_20951,N_28011);
nand U33428 (N_33428,N_20562,N_28522);
or U33429 (N_33429,N_29885,N_24819);
or U33430 (N_33430,N_23257,N_21947);
xor U33431 (N_33431,N_24480,N_22204);
xor U33432 (N_33432,N_29224,N_26190);
xnor U33433 (N_33433,N_29100,N_29589);
and U33434 (N_33434,N_27313,N_29267);
nand U33435 (N_33435,N_21721,N_22722);
and U33436 (N_33436,N_27112,N_23565);
or U33437 (N_33437,N_21622,N_22664);
or U33438 (N_33438,N_29375,N_21813);
nand U33439 (N_33439,N_26486,N_23178);
and U33440 (N_33440,N_26387,N_29367);
or U33441 (N_33441,N_21310,N_28034);
nand U33442 (N_33442,N_28037,N_25728);
or U33443 (N_33443,N_28368,N_27411);
xor U33444 (N_33444,N_25425,N_27234);
or U33445 (N_33445,N_24590,N_28233);
nor U33446 (N_33446,N_26146,N_27495);
or U33447 (N_33447,N_24442,N_23722);
xnor U33448 (N_33448,N_26607,N_22019);
nand U33449 (N_33449,N_28855,N_29495);
or U33450 (N_33450,N_27058,N_29603);
nor U33451 (N_33451,N_24050,N_24473);
nor U33452 (N_33452,N_27149,N_25649);
nand U33453 (N_33453,N_27754,N_24553);
nand U33454 (N_33454,N_28144,N_22102);
nand U33455 (N_33455,N_27934,N_24011);
nand U33456 (N_33456,N_24769,N_21956);
and U33457 (N_33457,N_21630,N_24574);
nand U33458 (N_33458,N_28288,N_21561);
nor U33459 (N_33459,N_22583,N_29098);
or U33460 (N_33460,N_29196,N_20615);
nand U33461 (N_33461,N_29833,N_24634);
xor U33462 (N_33462,N_26695,N_29597);
or U33463 (N_33463,N_22300,N_26702);
nor U33464 (N_33464,N_27226,N_20128);
or U33465 (N_33465,N_26772,N_20054);
nand U33466 (N_33466,N_23112,N_26013);
nor U33467 (N_33467,N_29776,N_29215);
or U33468 (N_33468,N_20171,N_22050);
or U33469 (N_33469,N_25137,N_28392);
xnor U33470 (N_33470,N_26350,N_26841);
nand U33471 (N_33471,N_24979,N_28330);
and U33472 (N_33472,N_27359,N_24673);
and U33473 (N_33473,N_24786,N_27413);
xor U33474 (N_33474,N_21465,N_23128);
or U33475 (N_33475,N_29905,N_23739);
nor U33476 (N_33476,N_26611,N_20865);
nor U33477 (N_33477,N_27196,N_29387);
nand U33478 (N_33478,N_25996,N_25241);
nand U33479 (N_33479,N_25931,N_27384);
and U33480 (N_33480,N_28018,N_27478);
nand U33481 (N_33481,N_21493,N_28251);
nand U33482 (N_33482,N_28341,N_21057);
nand U33483 (N_33483,N_24724,N_28321);
nand U33484 (N_33484,N_26426,N_27735);
or U33485 (N_33485,N_29403,N_26296);
nor U33486 (N_33486,N_23681,N_24727);
and U33487 (N_33487,N_22605,N_22987);
and U33488 (N_33488,N_20224,N_29435);
or U33489 (N_33489,N_28814,N_24613);
and U33490 (N_33490,N_23289,N_20976);
nand U33491 (N_33491,N_23731,N_29262);
nand U33492 (N_33492,N_24110,N_28102);
nor U33493 (N_33493,N_27955,N_28101);
and U33494 (N_33494,N_20216,N_25839);
and U33495 (N_33495,N_24978,N_26356);
or U33496 (N_33496,N_28530,N_26096);
and U33497 (N_33497,N_25437,N_26907);
nand U33498 (N_33498,N_25994,N_23653);
and U33499 (N_33499,N_27992,N_23254);
xor U33500 (N_33500,N_25153,N_25268);
xnor U33501 (N_33501,N_27299,N_26863);
nand U33502 (N_33502,N_29456,N_25338);
and U33503 (N_33503,N_24543,N_29727);
xnor U33504 (N_33504,N_28130,N_23774);
nand U33505 (N_33505,N_25563,N_22766);
nor U33506 (N_33506,N_29962,N_26291);
and U33507 (N_33507,N_28239,N_21037);
nor U33508 (N_33508,N_25968,N_22874);
nor U33509 (N_33509,N_24649,N_23520);
and U33510 (N_33510,N_27599,N_20082);
nand U33511 (N_33511,N_20989,N_24643);
nor U33512 (N_33512,N_21929,N_22473);
or U33513 (N_33513,N_21023,N_22349);
xor U33514 (N_33514,N_28780,N_21088);
and U33515 (N_33515,N_25225,N_21595);
or U33516 (N_33516,N_23009,N_21760);
and U33517 (N_33517,N_25430,N_24458);
nor U33518 (N_33518,N_25630,N_27547);
or U33519 (N_33519,N_29351,N_22338);
nor U33520 (N_33520,N_29560,N_29708);
nor U33521 (N_33521,N_25145,N_26364);
nor U33522 (N_33522,N_29883,N_20037);
and U33523 (N_33523,N_29896,N_29352);
and U33524 (N_33524,N_26319,N_22186);
nor U33525 (N_33525,N_26242,N_27943);
nor U33526 (N_33526,N_23771,N_27436);
or U33527 (N_33527,N_29441,N_24996);
or U33528 (N_33528,N_24960,N_24975);
or U33529 (N_33529,N_29427,N_23463);
nand U33530 (N_33530,N_22656,N_25889);
nor U33531 (N_33531,N_26835,N_21078);
nor U33532 (N_33532,N_21386,N_29063);
nor U33533 (N_33533,N_23915,N_27347);
or U33534 (N_33534,N_25827,N_27772);
or U33535 (N_33535,N_24827,N_20879);
and U33536 (N_33536,N_27962,N_23598);
nand U33537 (N_33537,N_23015,N_23097);
or U33538 (N_33538,N_27066,N_27114);
xnor U33539 (N_33539,N_28509,N_29182);
and U33540 (N_33540,N_25719,N_21934);
and U33541 (N_33541,N_29829,N_20656);
and U33542 (N_33542,N_27751,N_27132);
nand U33543 (N_33543,N_25179,N_21303);
nor U33544 (N_33544,N_24343,N_28552);
xor U33545 (N_33545,N_26193,N_21142);
or U33546 (N_33546,N_23610,N_29682);
or U33547 (N_33547,N_21253,N_21374);
and U33548 (N_33548,N_20314,N_26499);
nand U33549 (N_33549,N_24503,N_27107);
nor U33550 (N_33550,N_27189,N_26783);
nand U33551 (N_33551,N_25337,N_21105);
and U33552 (N_33552,N_20308,N_28030);
and U33553 (N_33553,N_23886,N_29342);
nor U33554 (N_33554,N_26902,N_27304);
xor U33555 (N_33555,N_27199,N_28188);
or U33556 (N_33556,N_20191,N_24976);
and U33557 (N_33557,N_22500,N_20512);
and U33558 (N_33558,N_29101,N_29656);
or U33559 (N_33559,N_26453,N_24298);
nand U33560 (N_33560,N_21601,N_25291);
nor U33561 (N_33561,N_24701,N_23316);
or U33562 (N_33562,N_21064,N_29094);
nand U33563 (N_33563,N_24756,N_22366);
nor U33564 (N_33564,N_24083,N_28235);
nand U33565 (N_33565,N_29963,N_26622);
xor U33566 (N_33566,N_24888,N_25972);
nor U33567 (N_33567,N_22878,N_27663);
nand U33568 (N_33568,N_25608,N_25079);
and U33569 (N_33569,N_28249,N_29890);
nor U33570 (N_33570,N_28079,N_22374);
and U33571 (N_33571,N_22149,N_22780);
nor U33572 (N_33572,N_28127,N_21621);
and U33573 (N_33573,N_24048,N_25369);
xor U33574 (N_33574,N_29632,N_25359);
xnor U33575 (N_33575,N_26086,N_24210);
nand U33576 (N_33576,N_20322,N_23444);
and U33577 (N_33577,N_23631,N_22867);
nand U33578 (N_33578,N_26573,N_24270);
xor U33579 (N_33579,N_22442,N_25216);
nand U33580 (N_33580,N_27205,N_21432);
or U33581 (N_33581,N_21476,N_23269);
and U33582 (N_33582,N_21062,N_21928);
nand U33583 (N_33583,N_29622,N_28700);
or U33584 (N_33584,N_23608,N_25169);
and U33585 (N_33585,N_20220,N_29690);
nand U33586 (N_33586,N_21274,N_22319);
or U33587 (N_33587,N_25471,N_28194);
or U33588 (N_33588,N_20137,N_23712);
or U33589 (N_33589,N_25054,N_26317);
and U33590 (N_33590,N_26563,N_20290);
or U33591 (N_33591,N_23851,N_28907);
and U33592 (N_33592,N_29151,N_21560);
or U33593 (N_33593,N_24593,N_28298);
and U33594 (N_33594,N_26674,N_27776);
and U33595 (N_33595,N_21040,N_26268);
nand U33596 (N_33596,N_28641,N_26906);
nor U33597 (N_33597,N_22877,N_28695);
nor U33598 (N_33598,N_20167,N_22249);
nor U33599 (N_33599,N_26572,N_22375);
nand U33600 (N_33600,N_25555,N_20659);
xor U33601 (N_33601,N_29372,N_28744);
or U33602 (N_33602,N_21864,N_24408);
and U33603 (N_33603,N_27895,N_28596);
and U33604 (N_33604,N_23671,N_29766);
nand U33605 (N_33605,N_29569,N_26312);
nor U33606 (N_33606,N_25822,N_27255);
nand U33607 (N_33607,N_24910,N_20758);
and U33608 (N_33608,N_28651,N_22739);
or U33609 (N_33609,N_22402,N_29600);
xnor U33610 (N_33610,N_26063,N_21926);
nor U33611 (N_33611,N_29067,N_25301);
or U33612 (N_33612,N_23933,N_22765);
and U33613 (N_33613,N_22582,N_29817);
nor U33614 (N_33614,N_22482,N_25671);
or U33615 (N_33615,N_25547,N_29068);
or U33616 (N_33616,N_25896,N_23232);
and U33617 (N_33617,N_28483,N_24149);
nor U33618 (N_33618,N_24122,N_28535);
nand U33619 (N_33619,N_21729,N_22113);
nor U33620 (N_33620,N_24717,N_26643);
or U33621 (N_33621,N_22617,N_20029);
nand U33622 (N_33622,N_24274,N_24013);
nand U33623 (N_33623,N_20459,N_25287);
nand U33624 (N_33624,N_25940,N_27686);
and U33625 (N_33625,N_25485,N_26137);
nand U33626 (N_33626,N_26037,N_23620);
nand U33627 (N_33627,N_23437,N_20826);
or U33628 (N_33628,N_24961,N_26078);
or U33629 (N_33629,N_29875,N_23935);
or U33630 (N_33630,N_28993,N_23332);
and U33631 (N_33631,N_21757,N_26506);
nand U33632 (N_33632,N_26825,N_24188);
and U33633 (N_33633,N_20937,N_26923);
nand U33634 (N_33634,N_23395,N_27356);
and U33635 (N_33635,N_24478,N_22936);
xor U33636 (N_33636,N_21574,N_20559);
nand U33637 (N_33637,N_21650,N_26640);
nand U33638 (N_33638,N_29493,N_24387);
xnor U33639 (N_33639,N_22266,N_28255);
nand U33640 (N_33640,N_20772,N_25947);
nand U33641 (N_33641,N_23628,N_21030);
xor U33642 (N_33642,N_20468,N_26688);
and U33643 (N_33643,N_22687,N_20194);
xnor U33644 (N_33644,N_28410,N_28245);
and U33645 (N_33645,N_29645,N_25566);
nor U33646 (N_33646,N_22143,N_25746);
xnor U33647 (N_33647,N_28894,N_27506);
and U33648 (N_33648,N_20083,N_28418);
nand U33649 (N_33649,N_20672,N_21869);
and U33650 (N_33650,N_26634,N_24209);
and U33651 (N_33651,N_25845,N_21762);
and U33652 (N_33652,N_20822,N_27207);
or U33653 (N_33653,N_22983,N_25935);
nand U33654 (N_33654,N_26798,N_24594);
nor U33655 (N_33655,N_24524,N_27262);
and U33656 (N_33656,N_21638,N_21139);
or U33657 (N_33657,N_29044,N_28236);
nor U33658 (N_33658,N_22208,N_27711);
nor U33659 (N_33659,N_27005,N_28674);
and U33660 (N_33660,N_28836,N_20404);
or U33661 (N_33661,N_27806,N_23423);
nor U33662 (N_33662,N_24348,N_28660);
xor U33663 (N_33663,N_26842,N_24777);
or U33664 (N_33664,N_23138,N_25516);
and U33665 (N_33665,N_23079,N_24477);
or U33666 (N_33666,N_26715,N_24455);
or U33667 (N_33667,N_27442,N_22279);
or U33668 (N_33668,N_26909,N_24542);
or U33669 (N_33669,N_22534,N_21118);
and U33670 (N_33670,N_24936,N_20143);
and U33671 (N_33671,N_25244,N_26145);
and U33672 (N_33672,N_25634,N_21572);
nor U33673 (N_33673,N_26120,N_24277);
and U33674 (N_33674,N_22673,N_22145);
and U33675 (N_33675,N_22959,N_28115);
nand U33676 (N_33676,N_28059,N_23563);
nor U33677 (N_33677,N_25841,N_26528);
or U33678 (N_33678,N_26525,N_28640);
nor U33679 (N_33679,N_27429,N_20050);
nor U33680 (N_33680,N_26363,N_21604);
nand U33681 (N_33681,N_28266,N_26478);
or U33682 (N_33682,N_23044,N_28601);
and U33683 (N_33683,N_27353,N_21332);
and U33684 (N_33684,N_22999,N_25008);
nor U33685 (N_33685,N_25363,N_26683);
nand U33686 (N_33686,N_23527,N_25077);
nor U33687 (N_33687,N_24040,N_20673);
or U33688 (N_33688,N_28877,N_24653);
nand U33689 (N_33689,N_20967,N_25913);
and U33690 (N_33690,N_21021,N_29558);
or U33691 (N_33691,N_27740,N_28670);
nor U33692 (N_33692,N_23072,N_26258);
nand U33693 (N_33693,N_28337,N_23721);
nor U33694 (N_33694,N_21800,N_28454);
nand U33695 (N_33695,N_21401,N_28359);
and U33696 (N_33696,N_22003,N_21661);
or U33697 (N_33697,N_27131,N_27265);
and U33698 (N_33698,N_24519,N_26168);
nor U33699 (N_33699,N_29292,N_21861);
nor U33700 (N_33700,N_23069,N_27098);
nor U33701 (N_33701,N_26129,N_23500);
or U33702 (N_33702,N_23693,N_21456);
or U33703 (N_33703,N_28443,N_25345);
and U33704 (N_33704,N_22371,N_29072);
or U33705 (N_33705,N_20183,N_28038);
and U33706 (N_33706,N_29398,N_28294);
or U33707 (N_33707,N_21854,N_29092);
or U33708 (N_33708,N_22721,N_24799);
or U33709 (N_33709,N_26225,N_25397);
nand U33710 (N_33710,N_27628,N_25835);
or U33711 (N_33711,N_23348,N_24924);
and U33712 (N_33712,N_27922,N_24113);
and U33713 (N_33713,N_22176,N_27762);
nor U33714 (N_33714,N_25202,N_21514);
xnor U33715 (N_33715,N_23380,N_20251);
nand U33716 (N_33716,N_25451,N_27374);
or U33717 (N_33717,N_29241,N_24230);
nand U33718 (N_33718,N_27535,N_22889);
nor U33719 (N_33719,N_23621,N_26901);
and U33720 (N_33720,N_22686,N_20607);
nand U33721 (N_33721,N_29575,N_27237);
and U33722 (N_33722,N_27695,N_22151);
nor U33723 (N_33723,N_22175,N_22523);
and U33724 (N_33724,N_21930,N_23938);
and U33725 (N_33725,N_26510,N_25067);
nor U33726 (N_33726,N_29047,N_29743);
nand U33727 (N_33727,N_24192,N_26762);
or U33728 (N_33728,N_29617,N_25526);
nand U33729 (N_33729,N_24452,N_29465);
xnor U33730 (N_33730,N_26659,N_20955);
or U33731 (N_33731,N_21002,N_21863);
or U33732 (N_33732,N_20935,N_27135);
nand U33733 (N_33733,N_22625,N_26313);
nor U33734 (N_33734,N_21799,N_22752);
nor U33735 (N_33735,N_22541,N_28532);
and U33736 (N_33736,N_26310,N_23139);
or U33737 (N_33737,N_23107,N_29941);
nand U33738 (N_33738,N_25914,N_22177);
and U33739 (N_33739,N_25599,N_22691);
or U33740 (N_33740,N_21700,N_29274);
xor U33741 (N_33741,N_26950,N_23640);
and U33742 (N_33742,N_20524,N_27284);
xnor U33743 (N_33743,N_28720,N_24584);
xnor U33744 (N_33744,N_26066,N_26034);
and U33745 (N_33745,N_27857,N_22387);
nor U33746 (N_33746,N_20443,N_27777);
and U33747 (N_33747,N_25828,N_26470);
xor U33748 (N_33748,N_27394,N_20288);
and U33749 (N_33749,N_24900,N_27856);
or U33750 (N_33750,N_29193,N_27572);
xor U33751 (N_33751,N_23142,N_26224);
and U33752 (N_33752,N_25959,N_26064);
nand U33753 (N_33753,N_21177,N_20203);
nor U33754 (N_33754,N_22236,N_27470);
nor U33755 (N_33755,N_21891,N_28176);
and U33756 (N_33756,N_23869,N_22240);
and U33757 (N_33757,N_23888,N_21154);
and U33758 (N_33758,N_21797,N_24742);
nand U33759 (N_33759,N_21431,N_25933);
nand U33760 (N_33760,N_28105,N_22900);
or U33761 (N_33761,N_27795,N_26526);
or U33762 (N_33762,N_21014,N_26004);
nand U33763 (N_33763,N_22123,N_28805);
nand U33764 (N_33764,N_25520,N_25007);
nand U33765 (N_33765,N_23795,N_20499);
nand U33766 (N_33766,N_20349,N_28723);
nor U33767 (N_33767,N_20027,N_20205);
and U33768 (N_33768,N_22923,N_21659);
nor U33769 (N_33769,N_25916,N_25964);
nor U33770 (N_33770,N_25243,N_23288);
and U33771 (N_33771,N_27346,N_22817);
or U33772 (N_33772,N_21032,N_21254);
and U33773 (N_33773,N_28616,N_23884);
and U33774 (N_33774,N_21306,N_20617);
nand U33775 (N_33775,N_21391,N_27150);
and U33776 (N_33776,N_25098,N_25747);
nor U33777 (N_33777,N_26459,N_20585);
xnor U33778 (N_33778,N_23475,N_23045);
nor U33779 (N_33779,N_27055,N_22137);
xor U33780 (N_33780,N_28677,N_21143);
or U33781 (N_33781,N_24349,N_20255);
and U33782 (N_33782,N_28840,N_21993);
nand U33783 (N_33783,N_22737,N_27050);
nand U33784 (N_33784,N_26959,N_29490);
nand U33785 (N_33785,N_23415,N_29148);
or U33786 (N_33786,N_26873,N_23747);
and U33787 (N_33787,N_26614,N_22798);
nor U33788 (N_33788,N_21827,N_25853);
nand U33789 (N_33789,N_21635,N_27566);
nor U33790 (N_33790,N_21888,N_29494);
nor U33791 (N_33791,N_28507,N_26334);
nand U33792 (N_33792,N_22530,N_23109);
and U33793 (N_33793,N_28526,N_26249);
nor U33794 (N_33794,N_25588,N_25392);
nor U33795 (N_33795,N_28391,N_28730);
nand U33796 (N_33796,N_21225,N_29764);
or U33797 (N_33797,N_26490,N_25187);
nand U33798 (N_33798,N_28833,N_29756);
nor U33799 (N_33799,N_21464,N_23140);
xnor U33800 (N_33800,N_26567,N_21666);
or U33801 (N_33801,N_21072,N_24678);
and U33802 (N_33802,N_23331,N_21261);
nand U33803 (N_33803,N_25573,N_27617);
and U33804 (N_33804,N_23076,N_22465);
nand U33805 (N_33805,N_25624,N_20496);
xor U33806 (N_33806,N_29373,N_23678);
and U33807 (N_33807,N_24451,N_26758);
nand U33808 (N_33808,N_29795,N_20554);
or U33809 (N_33809,N_26089,N_25466);
and U33810 (N_33810,N_21818,N_25718);
xnor U33811 (N_33811,N_23493,N_27121);
or U33812 (N_33812,N_26920,N_23899);
nand U33813 (N_33813,N_21219,N_23342);
or U33814 (N_33814,N_21067,N_24915);
nand U33815 (N_33815,N_24280,N_27295);
xor U33816 (N_33816,N_24716,N_28743);
and U33817 (N_33817,N_20731,N_25612);
and U33818 (N_33818,N_27596,N_29275);
nand U33819 (N_33819,N_25176,N_22427);
or U33820 (N_33820,N_28120,N_25870);
nand U33821 (N_33821,N_26085,N_22335);
and U33822 (N_33822,N_22156,N_24128);
nand U33823 (N_33823,N_20173,N_21648);
and U33824 (N_33824,N_21629,N_20834);
or U33825 (N_33825,N_21194,N_21319);
nand U33826 (N_33826,N_21858,N_26967);
xor U33827 (N_33827,N_27348,N_20906);
and U33828 (N_33828,N_25997,N_25333);
nor U33829 (N_33829,N_21010,N_20671);
or U33830 (N_33830,N_25335,N_29324);
or U33831 (N_33831,N_23137,N_25558);
nand U33832 (N_33832,N_24841,N_25604);
and U33833 (N_33833,N_25228,N_24608);
and U33834 (N_33834,N_28205,N_28754);
and U33835 (N_33835,N_26165,N_22261);
xnor U33836 (N_33836,N_23911,N_26765);
nor U33837 (N_33837,N_21851,N_21553);
or U33838 (N_33838,N_29093,N_20648);
or U33839 (N_33839,N_25482,N_28792);
nor U33840 (N_33840,N_22680,N_28541);
or U33841 (N_33841,N_28006,N_24470);
and U33842 (N_33842,N_27728,N_20991);
or U33843 (N_33843,N_22263,N_21587);
nor U33844 (N_33844,N_22318,N_21082);
nor U33845 (N_33845,N_29678,N_27067);
nor U33846 (N_33846,N_25529,N_29498);
and U33847 (N_33847,N_22096,N_28619);
nand U33848 (N_33848,N_21099,N_28921);
nand U33849 (N_33849,N_26214,N_22235);
nand U33850 (N_33850,N_26636,N_21180);
nand U33851 (N_33851,N_23530,N_22444);
and U33852 (N_33852,N_28990,N_25820);
nor U33853 (N_33853,N_22206,N_26444);
xnor U33854 (N_33854,N_27443,N_24781);
nor U33855 (N_33855,N_29677,N_26117);
and U33856 (N_33856,N_22496,N_25560);
nor U33857 (N_33857,N_29238,N_29842);
xnor U33858 (N_33858,N_26787,N_23028);
and U33859 (N_33859,N_28776,N_29529);
nor U33860 (N_33860,N_29121,N_27736);
nor U33861 (N_33861,N_26810,N_23409);
nor U33862 (N_33862,N_27907,N_23491);
and U33863 (N_33863,N_22461,N_20919);
nor U33864 (N_33864,N_27400,N_20959);
and U33865 (N_33865,N_29520,N_29931);
xnor U33866 (N_33866,N_27438,N_23505);
nor U33867 (N_33867,N_21222,N_28724);
nand U33868 (N_33868,N_27745,N_20667);
and U33869 (N_33869,N_24541,N_20067);
and U33870 (N_33870,N_26696,N_28803);
nand U33871 (N_33871,N_21550,N_27046);
or U33872 (N_33872,N_29170,N_28151);
or U33873 (N_33873,N_25474,N_20978);
nor U33874 (N_33874,N_21654,N_21991);
and U33875 (N_33875,N_26612,N_23016);
and U33876 (N_33876,N_23659,N_29453);
or U33877 (N_33877,N_25257,N_23053);
and U33878 (N_33878,N_24491,N_26821);
and U33879 (N_33879,N_20698,N_24388);
nor U33880 (N_33880,N_26050,N_24609);
nand U33881 (N_33881,N_29222,N_25734);
or U33882 (N_33882,N_29253,N_20778);
or U33883 (N_33883,N_27209,N_23923);
or U33884 (N_33884,N_24389,N_25685);
nand U33885 (N_33885,N_20753,N_20780);
or U33886 (N_33886,N_25250,N_25902);
and U33887 (N_33887,N_24885,N_26862);
xnor U33888 (N_33888,N_21961,N_23442);
or U33889 (N_33889,N_24151,N_23812);
and U33890 (N_33890,N_25356,N_28080);
xnor U33891 (N_33891,N_22840,N_25546);
or U33892 (N_33892,N_22715,N_20867);
nand U33893 (N_33893,N_22796,N_22847);
and U33894 (N_33894,N_25867,N_24581);
and U33895 (N_33895,N_24939,N_29997);
xnor U33896 (N_33896,N_21834,N_23785);
nor U33897 (N_33897,N_25148,N_27120);
xor U33898 (N_33898,N_21085,N_22449);
or U33899 (N_33899,N_24856,N_22781);
nor U33900 (N_33900,N_27133,N_26422);
or U33901 (N_33901,N_23698,N_22222);
nand U33902 (N_33902,N_23422,N_28794);
nand U33903 (N_33903,N_24522,N_29802);
or U33904 (N_33904,N_29091,N_20416);
or U33905 (N_33905,N_27054,N_22209);
or U33906 (N_33906,N_21517,N_23770);
xor U33907 (N_33907,N_29477,N_25252);
nor U33908 (N_33908,N_28638,N_27871);
and U33909 (N_33909,N_20400,N_21780);
or U33910 (N_33910,N_25198,N_20563);
and U33911 (N_33911,N_28752,N_22367);
nand U33912 (N_33912,N_24617,N_23661);
or U33913 (N_33913,N_21534,N_21046);
and U33914 (N_33914,N_23962,N_21172);
nor U33915 (N_33915,N_22949,N_22513);
nand U33916 (N_33916,N_29384,N_28876);
or U33917 (N_33917,N_22621,N_23645);
nand U33918 (N_33918,N_25110,N_23688);
and U33919 (N_33919,N_27101,N_29546);
nor U33920 (N_33920,N_23999,N_23467);
or U33921 (N_33921,N_21473,N_21806);
and U33922 (N_33922,N_27047,N_25950);
and U33923 (N_33923,N_28635,N_20596);
nor U33924 (N_33924,N_28112,N_29340);
nor U33925 (N_33925,N_26413,N_22233);
nand U33926 (N_33926,N_20161,N_23075);
and U33927 (N_33927,N_28729,N_27921);
nor U33928 (N_33928,N_28352,N_21776);
or U33929 (N_33929,N_24029,N_29480);
nand U33930 (N_33930,N_24892,N_28653);
nor U33931 (N_33931,N_28564,N_29537);
and U33932 (N_33932,N_21523,N_23383);
and U33933 (N_33933,N_26955,N_25876);
and U33934 (N_33934,N_20602,N_22736);
xnor U33935 (N_33935,N_25744,N_25721);
or U33936 (N_33936,N_20718,N_23085);
or U33937 (N_33937,N_27405,N_25086);
or U33938 (N_33938,N_25440,N_27681);
xnor U33939 (N_33939,N_27652,N_22108);
or U33940 (N_33940,N_29013,N_27640);
nand U33941 (N_33941,N_29794,N_29005);
nand U33942 (N_33942,N_25584,N_22089);
nand U33943 (N_33943,N_27090,N_29089);
nor U33944 (N_33944,N_28761,N_20624);
nor U33945 (N_33945,N_22836,N_23861);
or U33946 (N_33946,N_27892,N_29321);
nor U33947 (N_33947,N_22265,N_24311);
nand U33948 (N_33948,N_28905,N_26075);
nand U33949 (N_33949,N_21556,N_26107);
xor U33950 (N_33950,N_27044,N_21782);
or U33951 (N_33951,N_29906,N_29284);
nor U33952 (N_33952,N_26732,N_28007);
or U33953 (N_33953,N_20118,N_22914);
nand U33954 (N_33954,N_26685,N_25060);
or U33955 (N_33955,N_24696,N_22772);
nand U33956 (N_33956,N_28671,N_25780);
xnor U33957 (N_33957,N_29327,N_25256);
and U33958 (N_33958,N_22638,N_27707);
nand U33959 (N_33959,N_23532,N_23585);
or U33960 (N_33960,N_21495,N_21357);
nor U33961 (N_33961,N_24516,N_24242);
or U33962 (N_33962,N_28917,N_23847);
xnor U33963 (N_33963,N_21842,N_20859);
nand U33964 (N_33964,N_24283,N_26682);
and U33965 (N_33965,N_22723,N_24877);
and U33966 (N_33966,N_28346,N_27002);
or U33967 (N_33967,N_22378,N_24628);
nand U33968 (N_33968,N_29107,N_28399);
or U33969 (N_33969,N_23738,N_28379);
nand U33970 (N_33970,N_27788,N_29030);
or U33971 (N_33971,N_27318,N_20798);
nor U33972 (N_33972,N_27773,N_29891);
and U33973 (N_33973,N_28915,N_27393);
or U33974 (N_33974,N_26684,N_22568);
and U33975 (N_33975,N_22282,N_27741);
nand U33976 (N_33976,N_26479,N_20941);
xnor U33977 (N_33977,N_21460,N_25731);
xnor U33978 (N_33978,N_29723,N_23708);
and U33979 (N_33979,N_26522,N_22364);
nand U33980 (N_33980,N_27550,N_28843);
and U33981 (N_33981,N_20482,N_28801);
or U33982 (N_33982,N_25258,N_27855);
nor U33983 (N_33983,N_21196,N_25024);
or U33984 (N_33984,N_20368,N_22537);
nor U33985 (N_33985,N_21121,N_22038);
and U33986 (N_33986,N_23989,N_22762);
or U33987 (N_33987,N_23438,N_23440);
and U33988 (N_33988,N_29227,N_28685);
or U33989 (N_33989,N_25848,N_26465);
and U33990 (N_33990,N_27329,N_22749);
nor U33991 (N_33991,N_22289,N_20960);
nand U33992 (N_33992,N_29048,N_27587);
xor U33993 (N_33993,N_20278,N_21649);
or U33994 (N_33994,N_23870,N_21486);
or U33995 (N_33995,N_20651,N_23082);
nand U33996 (N_33996,N_29741,N_24689);
nand U33997 (N_33997,N_20250,N_24430);
nand U33998 (N_33998,N_23077,N_22147);
and U33999 (N_33999,N_27902,N_26194);
xnor U34000 (N_34000,N_23740,N_24913);
nand U34001 (N_34001,N_27181,N_20493);
and U34002 (N_34002,N_23734,N_29430);
nor U34003 (N_34003,N_26278,N_25886);
nor U34004 (N_34004,N_29981,N_20558);
or U34005 (N_34005,N_25875,N_21003);
xnor U34006 (N_34006,N_20442,N_23448);
and U34007 (N_34007,N_29309,N_27953);
or U34008 (N_34008,N_23656,N_29542);
xnor U34009 (N_34009,N_27811,N_26697);
nor U34010 (N_34010,N_25362,N_24166);
and U34011 (N_34011,N_25764,N_20855);
nand U34012 (N_34012,N_24267,N_29957);
and U34013 (N_34013,N_26833,N_25303);
nor U34014 (N_34014,N_29955,N_27030);
and U34015 (N_34015,N_29780,N_21887);
nor U34016 (N_34016,N_24793,N_28095);
and U34017 (N_34017,N_21252,N_20910);
and U34018 (N_34018,N_25449,N_23183);
nor U34019 (N_34019,N_27575,N_28775);
nor U34020 (N_34020,N_28687,N_22028);
or U34021 (N_34021,N_27099,N_22200);
or U34022 (N_34022,N_22118,N_28189);
or U34023 (N_34023,N_24256,N_21055);
nor U34024 (N_34024,N_24060,N_22262);
nand U34025 (N_34025,N_22963,N_22510);
or U34026 (N_34026,N_21558,N_26578);
nand U34027 (N_34027,N_24963,N_20830);
and U34028 (N_34028,N_23078,N_22824);
or U34029 (N_34029,N_22314,N_25509);
nand U34030 (N_34030,N_21371,N_28976);
nand U34031 (N_34031,N_26631,N_28785);
and U34032 (N_34032,N_29482,N_29293);
and U34033 (N_34033,N_21224,N_22259);
xnor U34034 (N_34034,N_22667,N_29724);
nand U34035 (N_34035,N_21593,N_21287);
nor U34036 (N_34036,N_26575,N_27578);
or U34037 (N_34037,N_24738,N_29483);
or U34038 (N_34038,N_21906,N_26591);
or U34039 (N_34039,N_28908,N_20211);
nor U34040 (N_34040,N_25702,N_29413);
nor U34041 (N_34041,N_20552,N_28782);
nor U34042 (N_34042,N_24771,N_25255);
nand U34043 (N_34043,N_28549,N_27878);
or U34044 (N_34044,N_25651,N_24657);
or U34045 (N_34045,N_20256,N_25803);
or U34046 (N_34046,N_26710,N_29619);
nand U34047 (N_34047,N_25932,N_22892);
and U34048 (N_34048,N_22940,N_26491);
or U34049 (N_34049,N_24988,N_21607);
or U34050 (N_34050,N_29899,N_22129);
and U34051 (N_34051,N_25765,N_26488);
nand U34052 (N_34052,N_27363,N_23447);
and U34053 (N_34053,N_26823,N_20719);
or U34054 (N_34054,N_21234,N_22078);
xor U34055 (N_34055,N_20198,N_22760);
nor U34056 (N_34056,N_21349,N_26815);
nor U34057 (N_34057,N_29008,N_20132);
xor U34058 (N_34058,N_21409,N_20616);
nor U34059 (N_34059,N_29329,N_21461);
nor U34060 (N_34060,N_23913,N_25078);
nand U34061 (N_34061,N_28021,N_27040);
xor U34062 (N_34062,N_29555,N_29229);
nand U34063 (N_34063,N_25009,N_24958);
and U34064 (N_34064,N_29535,N_20748);
nor U34065 (N_34065,N_29099,N_25452);
or U34066 (N_34066,N_26965,N_24787);
or U34067 (N_34067,N_28175,N_27134);
xor U34068 (N_34068,N_26515,N_28378);
or U34069 (N_34069,N_27537,N_21054);
or U34070 (N_34070,N_23929,N_26855);
nand U34071 (N_34071,N_27591,N_24646);
nand U34072 (N_34072,N_23672,N_21814);
nor U34073 (N_34073,N_24241,N_29900);
nand U34074 (N_34074,N_20264,N_21439);
and U34075 (N_34075,N_22857,N_29552);
or U34076 (N_34076,N_21663,N_26308);
nand U34077 (N_34077,N_22651,N_29915);
nand U34078 (N_34078,N_23106,N_28939);
or U34079 (N_34079,N_22803,N_27837);
and U34080 (N_34080,N_25064,N_22827);
nand U34081 (N_34081,N_20631,N_21452);
xnor U34082 (N_34082,N_27515,N_21390);
nand U34083 (N_34083,N_28712,N_27822);
or U34084 (N_34084,N_25323,N_21416);
or U34085 (N_34085,N_24227,N_20568);
nor U34086 (N_34086,N_27286,N_26288);
or U34087 (N_34087,N_26144,N_24901);
nand U34088 (N_34088,N_28573,N_26309);
nor U34089 (N_34089,N_20320,N_22615);
nand U34090 (N_34090,N_22384,N_22100);
nor U34091 (N_34091,N_27239,N_27093);
nand U34092 (N_34092,N_26542,N_25986);
nor U34093 (N_34093,N_21751,N_25755);
nor U34094 (N_34094,N_20948,N_24544);
and U34095 (N_34095,N_24168,N_29244);
nand U34096 (N_34096,N_22907,N_27445);
or U34097 (N_34097,N_25484,N_21868);
nor U34098 (N_34098,N_27110,N_22396);
or U34099 (N_34099,N_20816,N_22245);
nor U34100 (N_34100,N_29822,N_28476);
nor U34101 (N_34101,N_24213,N_21960);
xnor U34102 (N_34102,N_23529,N_25816);
nand U34103 (N_34103,N_20063,N_28056);
and U34104 (N_34104,N_29039,N_27157);
and U34105 (N_34105,N_22804,N_23359);
nand U34106 (N_34106,N_20280,N_20100);
nor U34107 (N_34107,N_20413,N_27987);
and U34108 (N_34108,N_21769,N_20739);
or U34109 (N_34109,N_24232,N_25448);
and U34110 (N_34110,N_20725,N_23274);
and U34111 (N_34111,N_23153,N_27485);
and U34112 (N_34112,N_23318,N_20754);
or U34113 (N_34113,N_25661,N_23202);
or U34114 (N_34114,N_20458,N_24352);
nand U34115 (N_34115,N_21897,N_29904);
and U34116 (N_34116,N_21186,N_21713);
and U34117 (N_34117,N_28393,N_26931);
xor U34118 (N_34118,N_26257,N_25866);
and U34119 (N_34119,N_25436,N_23363);
nor U34120 (N_34120,N_28768,N_21645);
nor U34121 (N_34121,N_21220,N_23181);
xor U34122 (N_34122,N_27273,N_26191);
nor U34123 (N_34123,N_26284,N_22415);
and U34124 (N_34124,N_25742,N_24427);
nor U34125 (N_34125,N_29333,N_26562);
xnor U34126 (N_34126,N_24390,N_23245);
nand U34127 (N_34127,N_26830,N_21865);
nor U34128 (N_34128,N_21327,N_21114);
nand U34129 (N_34129,N_20296,N_25270);
and U34130 (N_34130,N_26197,N_24019);
nand U34131 (N_34131,N_22121,N_23896);
and U34132 (N_34132,N_20501,N_25046);
nand U34133 (N_34133,N_22458,N_23988);
or U34134 (N_34134,N_26558,N_25227);
or U34135 (N_34135,N_20439,N_29172);
and U34136 (N_34136,N_24308,N_20508);
nor U34137 (N_34137,N_29206,N_28072);
or U34138 (N_34138,N_29471,N_20833);
nand U34139 (N_34139,N_22633,N_25613);
or U34140 (N_34140,N_22463,N_21417);
nor U34141 (N_34141,N_22903,N_26913);
or U34142 (N_34142,N_28961,N_26953);
nand U34143 (N_34143,N_28279,N_28286);
nand U34144 (N_34144,N_25128,N_29967);
and U34145 (N_34145,N_27932,N_25795);
and U34146 (N_34146,N_20236,N_27534);
xor U34147 (N_34147,N_22666,N_26419);
and U34148 (N_34148,N_28327,N_28816);
and U34149 (N_34149,N_25404,N_21429);
and U34150 (N_34150,N_25420,N_27626);
nor U34151 (N_34151,N_28548,N_23800);
and U34152 (N_34152,N_25136,N_28269);
or U34153 (N_34153,N_24732,N_28449);
and U34154 (N_34154,N_28945,N_21335);
or U34155 (N_34155,N_23038,N_27680);
nor U34156 (N_34156,N_26260,N_26030);
nand U34157 (N_34157,N_26641,N_21537);
xnor U34158 (N_34158,N_28381,N_28128);
xnor U34159 (N_34159,N_24502,N_21315);
nor U34160 (N_34160,N_26200,N_22231);
nand U34161 (N_34161,N_28689,N_26348);
nor U34162 (N_34162,N_21510,N_23426);
nand U34163 (N_34163,N_20431,N_25831);
nand U34164 (N_34164,N_24440,N_28482);
nor U34165 (N_34165,N_25800,N_22172);
nand U34166 (N_34166,N_29735,N_20683);
nand U34167 (N_34167,N_22174,N_25797);
nand U34168 (N_34168,N_26971,N_29207);
or U34169 (N_34169,N_25284,N_28500);
nand U34170 (N_34170,N_20541,N_24167);
nor U34171 (N_34171,N_20045,N_24551);
nand U34172 (N_34172,N_25694,N_24679);
or U34173 (N_34173,N_26687,N_24174);
and U34174 (N_34174,N_28531,N_21113);
or U34175 (N_34175,N_28746,N_22450);
nand U34176 (N_34176,N_23068,N_22588);
nor U34177 (N_34177,N_29186,N_26044);
or U34178 (N_34178,N_21754,N_26382);
xnor U34179 (N_34179,N_27784,N_25094);
nand U34180 (N_34180,N_27819,N_23420);
nor U34181 (N_34181,N_23983,N_25871);
or U34182 (N_34182,N_27845,N_26081);
and U34183 (N_34183,N_23965,N_22756);
xnor U34184 (N_34184,N_27074,N_29054);
and U34185 (N_34185,N_20494,N_21249);
nor U34186 (N_34186,N_20215,N_21692);
or U34187 (N_34187,N_29035,N_20849);
or U34188 (N_34188,N_26489,N_25142);
nor U34189 (N_34189,N_23054,N_21466);
and U34190 (N_34190,N_25496,N_26447);
nand U34191 (N_34191,N_26681,N_27319);
or U34192 (N_34192,N_29127,N_25004);
nand U34193 (N_34193,N_20389,N_27679);
and U34194 (N_34194,N_27682,N_26039);
or U34195 (N_34195,N_27779,N_20530);
and U34196 (N_34196,N_25912,N_26707);
nor U34197 (N_34197,N_21166,N_28446);
xnor U34198 (N_34198,N_22152,N_26720);
nand U34199 (N_34199,N_24760,N_27176);
and U34200 (N_34200,N_22453,N_23815);
or U34201 (N_34201,N_27103,N_29695);
and U34202 (N_34202,N_26297,N_27468);
nor U34203 (N_34203,N_21507,N_20420);
nor U34204 (N_34204,N_22726,N_22063);
or U34205 (N_34205,N_21238,N_20897);
nor U34206 (N_34206,N_25946,N_23582);
and U34207 (N_34207,N_20938,N_27583);
and U34208 (N_34208,N_29897,N_24007);
nor U34209 (N_34209,N_24446,N_24299);
or U34210 (N_34210,N_20379,N_21286);
xor U34211 (N_34211,N_28028,N_28367);
nor U34212 (N_34212,N_25403,N_20090);
nor U34213 (N_34213,N_26761,N_23827);
nor U34214 (N_34214,N_22698,N_20646);
xnor U34215 (N_34215,N_25049,N_27004);
and U34216 (N_34216,N_28595,N_27502);
xor U34217 (N_34217,N_22410,N_29813);
nand U34218 (N_34218,N_20789,N_24276);
and U34219 (N_34219,N_28430,N_22035);
or U34220 (N_34220,N_28608,N_21619);
nand U34221 (N_34221,N_29799,N_29119);
and U34222 (N_34222,N_26111,N_28098);
or U34223 (N_34223,N_28380,N_22388);
nor U34224 (N_34224,N_20386,N_22755);
nor U34225 (N_34225,N_23451,N_25687);
or U34226 (N_34226,N_29010,N_27303);
and U34227 (N_34227,N_24161,N_28844);
or U34228 (N_34228,N_29256,N_28309);
nand U34229 (N_34229,N_25739,N_20882);
nand U34230 (N_34230,N_29752,N_20103);
xnor U34231 (N_34231,N_24290,N_27768);
and U34232 (N_34232,N_23113,N_26131);
nor U34233 (N_34233,N_20924,N_23969);
xor U34234 (N_34234,N_25134,N_24501);
nand U34235 (N_34235,N_24393,N_23921);
nand U34236 (N_34236,N_24016,N_24699);
xnor U34237 (N_34237,N_27465,N_29306);
nand U34238 (N_34238,N_22317,N_25022);
nand U34239 (N_34239,N_20899,N_29951);
xor U34240 (N_34240,N_20451,N_21007);
xnor U34241 (N_34241,N_24968,N_29128);
or U34242 (N_34242,N_21730,N_22973);
or U34243 (N_34243,N_21442,N_23367);
or U34244 (N_34244,N_25611,N_24974);
nor U34245 (N_34245,N_26343,N_26136);
or U34246 (N_34246,N_26294,N_29747);
nand U34247 (N_34247,N_29669,N_24414);
and U34248 (N_34248,N_26764,N_20521);
nor U34249 (N_34249,N_24152,N_24259);
or U34250 (N_34250,N_27699,N_21227);
and U34251 (N_34251,N_28442,N_29871);
or U34252 (N_34252,N_23266,N_20207);
xnor U34253 (N_34253,N_23239,N_27218);
or U34254 (N_34254,N_26199,N_28202);
and U34255 (N_34255,N_26615,N_21564);
nor U34256 (N_34256,N_20716,N_22045);
or U34257 (N_34257,N_22815,N_23649);
and U34258 (N_34258,N_29940,N_25332);
nor U34259 (N_34259,N_21847,N_28468);
or U34260 (N_34260,N_20230,N_25040);
xor U34261 (N_34261,N_20670,N_28103);
or U34262 (N_34262,N_26388,N_26187);
and U34263 (N_34263,N_27158,N_27080);
or U34264 (N_34264,N_29976,N_29311);
and U34265 (N_34265,N_27229,N_29137);
or U34266 (N_34266,N_23635,N_23685);
and U34267 (N_34267,N_27254,N_29266);
and U34268 (N_34268,N_21212,N_29556);
and U34269 (N_34269,N_28138,N_29987);
nor U34270 (N_34270,N_20234,N_25246);
nand U34271 (N_34271,N_20098,N_24126);
and U34272 (N_34272,N_22689,N_22299);
nand U34273 (N_34273,N_26429,N_20102);
nand U34274 (N_34274,N_27831,N_21048);
and U34275 (N_34275,N_22150,N_27456);
and U34276 (N_34276,N_21228,N_23619);
or U34277 (N_34277,N_22972,N_21736);
or U34278 (N_34278,N_20253,N_22912);
nand U34279 (N_34279,N_25557,N_29543);
and U34280 (N_34280,N_26589,N_23766);
nor U34281 (N_34281,N_22793,N_23658);
nand U34282 (N_34282,N_24142,N_23925);
and U34283 (N_34283,N_20430,N_29576);
nand U34284 (N_34284,N_26750,N_22898);
nand U34285 (N_34285,N_26737,N_26743);
and U34286 (N_34286,N_28525,N_21324);
and U34287 (N_34287,N_29218,N_29894);
nand U34288 (N_34288,N_21944,N_27997);
or U34289 (N_34289,N_24691,N_24790);
and U34290 (N_34290,N_28892,N_23012);
xor U34291 (N_34291,N_28306,N_23048);
and U34292 (N_34292,N_23173,N_23270);
nor U34293 (N_34293,N_26565,N_22083);
and U34294 (N_34294,N_24814,N_28983);
nor U34295 (N_34295,N_22980,N_25453);
and U34296 (N_34296,N_24612,N_22601);
xnor U34297 (N_34297,N_29255,N_25945);
xor U34298 (N_34298,N_27560,N_27421);
or U34299 (N_34299,N_22897,N_26183);
nand U34300 (N_34300,N_24570,N_27365);
nor U34301 (N_34301,N_26843,N_23803);
nand U34302 (N_34302,N_26596,N_23807);
xor U34303 (N_34303,N_20273,N_21950);
xnor U34304 (N_34304,N_26569,N_29710);
nor U34305 (N_34305,N_21949,N_23157);
or U34306 (N_34306,N_22244,N_28217);
nand U34307 (N_34307,N_26926,N_26178);
or U34308 (N_34308,N_22926,N_29082);
or U34309 (N_34309,N_26148,N_20166);
nand U34310 (N_34310,N_21484,N_20074);
or U34311 (N_34311,N_20872,N_26689);
and U34312 (N_34312,N_20077,N_20105);
nor U34313 (N_34313,N_23647,N_21004);
xor U34314 (N_34314,N_20963,N_28474);
xor U34315 (N_34315,N_21898,N_27409);
nor U34316 (N_34316,N_29719,N_28089);
or U34317 (N_34317,N_21208,N_23480);
nand U34318 (N_34318,N_21070,N_20406);
or U34319 (N_34319,N_20757,N_25697);
nor U34320 (N_34320,N_22268,N_21588);
nor U34321 (N_34321,N_23939,N_27300);
nand U34322 (N_34322,N_20342,N_25683);
xnor U34323 (N_34323,N_28055,N_25954);
nand U34324 (N_34324,N_26709,N_20893);
and U34325 (N_34325,N_25923,N_29343);
or U34326 (N_34326,N_23889,N_21061);
nor U34327 (N_34327,N_23982,N_25149);
and U34328 (N_34328,N_25158,N_22991);
or U34329 (N_34329,N_24236,N_27794);
or U34330 (N_34330,N_28014,N_21270);
and U34331 (N_34331,N_28197,N_20828);
xor U34332 (N_34332,N_22732,N_26439);
xor U34333 (N_34333,N_21111,N_27349);
and U34334 (N_34334,N_28051,N_27130);
and U34335 (N_34335,N_24536,N_28872);
or U34336 (N_34336,N_23300,N_29630);
or U34337 (N_34337,N_29290,N_26866);
nand U34338 (N_34338,N_26691,N_29694);
nor U34339 (N_34339,N_22567,N_21758);
and U34340 (N_34340,N_20390,N_26812);
and U34341 (N_34341,N_28486,N_29159);
and U34342 (N_34342,N_20047,N_26865);
or U34343 (N_34343,N_27310,N_24680);
nor U34344 (N_34344,N_22452,N_22855);
and U34345 (N_34345,N_21597,N_23394);
nor U34346 (N_34346,N_29388,N_22369);
and U34347 (N_34347,N_26256,N_21878);
and U34348 (N_34348,N_23578,N_25205);
nand U34349 (N_34349,N_27063,N_24687);
nor U34350 (N_34350,N_23000,N_26077);
or U34351 (N_34351,N_24702,N_21299);
or U34352 (N_34352,N_25665,N_29365);
nor U34353 (N_34353,N_27898,N_21457);
nand U34354 (N_34354,N_28910,N_23309);
nand U34355 (N_34355,N_28181,N_23629);
or U34356 (N_34356,N_28793,N_26374);
nand U34357 (N_34357,N_26751,N_24094);
nand U34358 (N_34358,N_27160,N_20536);
nor U34359 (N_34359,N_24338,N_29845);
nor U34360 (N_34360,N_24982,N_22913);
and U34361 (N_34361,N_29877,N_22440);
or U34362 (N_34362,N_25467,N_26978);
nor U34363 (N_34363,N_22909,N_25000);
nor U34364 (N_34364,N_29947,N_24405);
nor U34365 (N_34365,N_23043,N_25213);
nand U34366 (N_34366,N_29428,N_26266);
or U34367 (N_34367,N_20135,N_25750);
nand U34368 (N_34368,N_29364,N_23752);
and U34369 (N_34369,N_21387,N_29716);
or U34370 (N_34370,N_25601,N_21519);
or U34371 (N_34371,N_21013,N_28937);
and U34372 (N_34372,N_27364,N_28510);
xor U34373 (N_34373,N_26076,N_23603);
and U34374 (N_34374,N_21260,N_22663);
nor U34375 (N_34375,N_20061,N_25802);
nor U34376 (N_34376,N_24085,N_22614);
nand U34377 (N_34377,N_27974,N_20261);
or U34378 (N_34378,N_20437,N_25053);
nor U34379 (N_34379,N_20660,N_24804);
nor U34380 (N_34380,N_24736,N_29345);
or U34381 (N_34381,N_22008,N_22431);
nand U34382 (N_34382,N_29986,N_23261);
or U34383 (N_34383,N_27448,N_20653);
nand U34384 (N_34384,N_28307,N_28139);
nor U34385 (N_34385,N_26962,N_22219);
nand U34386 (N_34386,N_20649,N_28850);
nor U34387 (N_34387,N_28763,N_28025);
nand U34388 (N_34388,N_20429,N_22331);
xor U34389 (N_34389,N_26140,N_24074);
and U34390 (N_34390,N_28579,N_22194);
nand U34391 (N_34391,N_24371,N_22481);
and U34392 (N_34392,N_28259,N_23744);
nand U34393 (N_34393,N_22532,N_21445);
and U34394 (N_34394,N_23521,N_27642);
or U34395 (N_34395,N_26385,N_21883);
nand U34396 (N_34396,N_26245,N_25814);
nand U34397 (N_34397,N_26401,N_25407);
or U34398 (N_34398,N_27562,N_24144);
nor U34399 (N_34399,N_29399,N_29956);
or U34400 (N_34400,N_21025,N_20723);
or U34401 (N_34401,N_20663,N_21257);
or U34402 (N_34402,N_23067,N_24425);
nand U34403 (N_34403,N_26805,N_27834);
and U34404 (N_34404,N_27703,N_23788);
nor U34405 (N_34405,N_24865,N_21424);
nor U34406 (N_34406,N_22750,N_28667);
or U34407 (N_34407,N_22301,N_21364);
nand U34408 (N_34408,N_27800,N_21835);
or U34409 (N_34409,N_23732,N_28977);
nor U34410 (N_34410,N_28406,N_23797);
or U34411 (N_34411,N_22908,N_23941);
nand U34412 (N_34412,N_25140,N_27144);
or U34413 (N_34413,N_26280,N_26464);
xnor U34414 (N_34414,N_28562,N_25688);
xor U34415 (N_34415,N_21677,N_28238);
nor U34416 (N_34416,N_26316,N_20447);
nand U34417 (N_34417,N_29401,N_29062);
nand U34418 (N_34418,N_27747,N_22592);
or U34419 (N_34419,N_20884,N_27277);
and U34420 (N_34420,N_24309,N_24426);
or U34421 (N_34421,N_29374,N_23942);
or U34422 (N_34422,N_22985,N_29421);
and U34423 (N_34423,N_29251,N_26986);
or U34424 (N_34424,N_25282,N_24207);
xnor U34425 (N_34425,N_26369,N_20181);
and U34426 (N_34426,N_23830,N_27980);
or U34427 (N_34427,N_21231,N_22334);
nand U34428 (N_34428,N_27280,N_22655);
nor U34429 (N_34429,N_22955,N_24264);
or U34430 (N_34430,N_26845,N_27975);
nor U34431 (N_34431,N_24884,N_29781);
nand U34432 (N_34432,N_28033,N_23055);
xnor U34433 (N_34433,N_21711,N_27165);
or U34434 (N_34434,N_20705,N_23834);
or U34435 (N_34435,N_25285,N_21709);
and U34436 (N_34436,N_24780,N_29181);
xnor U34437 (N_34437,N_25855,N_25786);
and U34438 (N_34438,N_24136,N_29821);
and U34439 (N_34439,N_23211,N_28520);
and U34440 (N_34440,N_29730,N_23468);
nor U34441 (N_34441,N_24583,N_21539);
nor U34442 (N_34442,N_29214,N_23080);
and U34443 (N_34443,N_26396,N_20277);
xnor U34444 (N_34444,N_21794,N_22852);
or U34445 (N_34445,N_26010,N_27529);
or U34446 (N_34446,N_29038,N_25504);
nand U34447 (N_34447,N_23145,N_29146);
or U34448 (N_34448,N_27739,N_20784);
or U34449 (N_34449,N_21268,N_22818);
or U34450 (N_34450,N_22802,N_29607);
nor U34451 (N_34451,N_28553,N_23477);
nand U34452 (N_34452,N_23682,N_26098);
and U34453 (N_34453,N_24969,N_22032);
xnor U34454 (N_34454,N_26404,N_20883);
or U34455 (N_34455,N_21706,N_29807);
nor U34456 (N_34456,N_21997,N_20197);
and U34457 (N_34457,N_26795,N_25154);
nand U34458 (N_34458,N_25590,N_20470);
or U34459 (N_34459,N_24515,N_23654);
nand U34460 (N_34460,N_23558,N_25365);
and U34461 (N_34461,N_23136,N_21978);
nor U34462 (N_34462,N_27251,N_25502);
or U34463 (N_34463,N_23994,N_27869);
or U34464 (N_34464,N_21784,N_28300);
and U34465 (N_34465,N_27164,N_26669);
xnor U34466 (N_34466,N_23804,N_28099);
nand U34467 (N_34467,N_28427,N_26898);
or U34468 (N_34468,N_20270,N_24369);
and U34469 (N_34469,N_29803,N_26344);
nand U34470 (N_34470,N_23335,N_23343);
and U34471 (N_34471,N_27168,N_24565);
nand U34472 (N_34472,N_25519,N_26434);
and U34473 (N_34473,N_22799,N_21323);
nor U34474 (N_34474,N_25417,N_28527);
xnor U34475 (N_34475,N_27410,N_21541);
nor U34476 (N_34476,N_21918,N_25756);
and U34477 (N_34477,N_27500,N_29150);
nor U34478 (N_34478,N_21351,N_23906);
nor U34479 (N_34479,N_28401,N_27048);
and U34480 (N_34480,N_29254,N_20740);
and U34481 (N_34481,N_21756,N_28340);
and U34482 (N_34482,N_20087,N_25823);
nand U34483 (N_34483,N_24810,N_28625);
nand U34484 (N_34484,N_25113,N_25847);
nand U34485 (N_34485,N_28078,N_25088);
nor U34486 (N_34486,N_24768,N_20841);
nor U34487 (N_34487,N_27613,N_21636);
and U34488 (N_34488,N_23964,N_24401);
or U34489 (N_34489,N_20101,N_22775);
or U34490 (N_34490,N_27497,N_21505);
nor U34491 (N_34491,N_24886,N_26164);
or U34492 (N_34492,N_27937,N_21277);
or U34493 (N_34493,N_21979,N_23959);
or U34494 (N_34494,N_26358,N_26006);
and U34495 (N_34495,N_20271,N_22404);
and U34496 (N_34496,N_25741,N_24178);
nor U34497 (N_34497,N_20455,N_27415);
nand U34498 (N_34498,N_23919,N_29064);
xnor U34499 (N_34499,N_28360,N_23381);
and U34500 (N_34500,N_26936,N_25753);
and U34501 (N_34501,N_21475,N_21977);
nor U34502 (N_34502,N_20348,N_24323);
or U34503 (N_34503,N_21896,N_20571);
nand U34504 (N_34504,N_29702,N_24251);
nand U34505 (N_34505,N_23756,N_22036);
nand U34506 (N_34506,N_20890,N_22351);
nand U34507 (N_34507,N_25844,N_29081);
or U34508 (N_34508,N_21945,N_28024);
or U34509 (N_34509,N_25581,N_22348);
or U34510 (N_34510,N_21942,N_29463);
and U34511 (N_34511,N_27000,N_23041);
and U34512 (N_34512,N_29994,N_24449);
nor U34513 (N_34513,N_25551,N_29272);
and U34514 (N_34514,N_23297,N_24162);
or U34515 (N_34515,N_28767,N_21159);
nor U34516 (N_34516,N_27031,N_27839);
nand U34517 (N_34517,N_25165,N_27525);
and U34518 (N_34518,N_20252,N_26336);
or U34519 (N_34519,N_23963,N_23689);
nand U34520 (N_34520,N_29302,N_24523);
nand U34521 (N_34521,N_23871,N_27517);
or U34522 (N_34522,N_24327,N_29339);
or U34523 (N_34523,N_25635,N_24175);
or U34524 (N_34524,N_23707,N_20578);
or U34525 (N_34525,N_24220,N_28304);
nand U34526 (N_34526,N_27186,N_21406);
nor U34527 (N_34527,N_24622,N_22207);
nor U34528 (N_34528,N_27605,N_21674);
or U34529 (N_34529,N_26987,N_28223);
nor U34530 (N_34530,N_27959,N_25833);
or U34531 (N_34531,N_26052,N_25955);
and U34532 (N_34532,N_24744,N_26610);
nand U34533 (N_34533,N_26799,N_28292);
and U34534 (N_34534,N_26074,N_22139);
and U34535 (N_34535,N_29219,N_20669);
nor U34536 (N_34536,N_22507,N_26602);
nor U34537 (N_34537,N_24296,N_26996);
xnor U34538 (N_34538,N_27147,N_24580);
or U34539 (N_34539,N_27471,N_27858);
xor U34540 (N_34540,N_24874,N_26872);
nand U34541 (N_34541,N_27241,N_29472);
or U34542 (N_34542,N_20729,N_29540);
or U34543 (N_34543,N_28593,N_24197);
xor U34544 (N_34544,N_27392,N_22658);
xor U34545 (N_34545,N_20535,N_23329);
nand U34546 (N_34546,N_26666,N_27756);
nor U34547 (N_34547,N_22022,N_24407);
nand U34548 (N_34548,N_27430,N_28010);
nor U34549 (N_34549,N_21815,N_20383);
nor U34550 (N_34550,N_20160,N_24668);
or U34551 (N_34551,N_23284,N_26271);
and U34552 (N_34552,N_28973,N_20107);
xnor U34553 (N_34553,N_24954,N_21859);
and U34554 (N_34554,N_20486,N_25595);
or U34555 (N_34555,N_20537,N_23819);
and U34556 (N_34556,N_21450,N_27437);
and U34557 (N_34557,N_24355,N_24461);
xnor U34558 (N_34558,N_24899,N_20840);
nand U34559 (N_34559,N_27094,N_22519);
and U34560 (N_34560,N_24140,N_25141);
nand U34561 (N_34561,N_20717,N_20891);
or U34562 (N_34562,N_29765,N_21489);
nand U34563 (N_34563,N_23523,N_24560);
and U34564 (N_34564,N_28538,N_21513);
nor U34565 (N_34565,N_20353,N_21193);
nand U34566 (N_34566,N_23648,N_21936);
nor U34567 (N_34567,N_21586,N_22943);
and U34568 (N_34568,N_22014,N_23030);
and U34569 (N_34569,N_29397,N_28789);
nand U34570 (N_34570,N_23761,N_28675);
and U34571 (N_34571,N_23404,N_28751);
nand U34572 (N_34572,N_22418,N_28361);
nor U34573 (N_34573,N_24099,N_24552);
nor U34574 (N_34574,N_20337,N_28433);
and U34575 (N_34575,N_24184,N_25074);
nand U34576 (N_34576,N_26274,N_27453);
nand U34577 (N_34577,N_23903,N_22130);
or U34578 (N_34578,N_29479,N_25571);
nand U34579 (N_34579,N_22643,N_23509);
nor U34580 (N_34580,N_26981,N_23127);
xor U34581 (N_34581,N_24441,N_22859);
nor U34582 (N_34582,N_22632,N_25676);
nand U34583 (N_34583,N_27027,N_29424);
or U34584 (N_34584,N_24919,N_28857);
nand U34585 (N_34585,N_23240,N_28628);
nor U34586 (N_34586,N_21496,N_26217);
or U34587 (N_34587,N_28567,N_22377);
nor U34588 (N_34588,N_21753,N_29837);
nor U34589 (N_34589,N_23160,N_21330);
or U34590 (N_34590,N_21192,N_22710);
nor U34591 (N_34591,N_20395,N_22138);
and U34592 (N_34592,N_22430,N_29518);
nand U34593 (N_34593,N_24833,N_23912);
or U34594 (N_34594,N_27412,N_26414);
or U34595 (N_34595,N_24181,N_23684);
nand U34596 (N_34596,N_26594,N_29217);
and U34597 (N_34597,N_22146,N_20371);
or U34598 (N_34598,N_27011,N_29440);
or U34599 (N_34599,N_26116,N_23403);
and U34600 (N_34600,N_29385,N_27972);
or U34601 (N_34601,N_21414,N_27450);
nor U34602 (N_34602,N_24463,N_22232);
nand U34603 (N_34603,N_25682,N_22584);
nor U34604 (N_34604,N_27230,N_27860);
nor U34605 (N_34605,N_28114,N_20434);
nor U34606 (N_34606,N_26679,N_27108);
nor U34607 (N_34607,N_22157,N_23980);
nor U34608 (N_34608,N_29308,N_25622);
nor U34609 (N_34609,N_27545,N_27060);
nand U34610 (N_34610,N_27978,N_20382);
and U34611 (N_34611,N_23699,N_27697);
and U34612 (N_34612,N_27242,N_20089);
and U34613 (N_34613,N_27946,N_25781);
or U34614 (N_34614,N_22668,N_25215);
nand U34615 (N_34615,N_20329,N_20282);
nand U34616 (N_34616,N_29884,N_20363);
or U34617 (N_34617,N_22094,N_24931);
nor U34618 (N_34618,N_21394,N_27075);
or U34619 (N_34619,N_25636,N_20109);
nand U34620 (N_34620,N_27758,N_20770);
nand U34621 (N_34621,N_23070,N_24017);
nand U34622 (N_34622,N_22140,N_25340);
and U34623 (N_34623,N_28880,N_29557);
or U34624 (N_34624,N_21163,N_23472);
nor U34625 (N_34625,N_25231,N_27862);
or U34626 (N_34626,N_25894,N_21665);
nand U34627 (N_34627,N_28985,N_20681);
nor U34628 (N_34628,N_20582,N_21866);
or U34629 (N_34629,N_24688,N_27480);
nor U34630 (N_34630,N_23726,N_22865);
nor U34631 (N_34631,N_29114,N_25675);
nand U34632 (N_34632,N_20553,N_29016);
or U34633 (N_34633,N_21996,N_22777);
xnor U34634 (N_34634,N_20292,N_28041);
or U34635 (N_34635,N_29112,N_26983);
or U34636 (N_34636,N_20677,N_25544);
and U34637 (N_34637,N_20204,N_21786);
nor U34638 (N_34638,N_20079,N_28387);
nand U34639 (N_34639,N_25073,N_29965);
and U34640 (N_34640,N_24778,N_24249);
nand U34641 (N_34641,N_24156,N_22199);
nor U34642 (N_34642,N_24637,N_22264);
nand U34643 (N_34643,N_21058,N_28682);
or U34644 (N_34644,N_28481,N_24098);
nor U34645 (N_34645,N_28506,N_20598);
nor U34646 (N_34646,N_29444,N_23215);
or U34647 (N_34647,N_28925,N_23014);
and U34648 (N_34648,N_23940,N_24625);
and U34649 (N_34649,N_24183,N_28335);
and U34650 (N_34650,N_25181,N_27925);
xnor U34651 (N_34651,N_20153,N_22555);
or U34652 (N_34652,N_29692,N_22419);
or U34653 (N_34653,N_28949,N_28395);
nand U34654 (N_34654,N_22011,N_27481);
or U34655 (N_34655,N_24045,N_22869);
or U34656 (N_34656,N_27222,N_22819);
or U34657 (N_34657,N_26152,N_22326);
nand U34658 (N_34658,N_29919,N_26091);
or U34659 (N_34659,N_24032,N_28757);
nor U34660 (N_34660,N_22285,N_21927);
or U34661 (N_34661,N_26518,N_26124);
or U34662 (N_34662,N_23971,N_24983);
xor U34663 (N_34663,N_26997,N_24104);
or U34664 (N_34664,N_29291,N_22770);
nor U34665 (N_34665,N_22457,N_27459);
nor U34666 (N_34666,N_29586,N_26924);
or U34667 (N_34667,N_23206,N_29260);
nand U34668 (N_34668,N_28133,N_24395);
nor U34669 (N_34669,N_28355,N_27195);
nand U34670 (N_34670,N_24729,N_28461);
nor U34671 (N_34671,N_29620,N_25714);
nor U34672 (N_34672,N_26882,N_27891);
nor U34673 (N_34673,N_24869,N_27352);
and U34674 (N_34674,N_20854,N_24922);
and U34675 (N_34675,N_29606,N_24693);
or U34676 (N_34676,N_27771,N_29573);
nand U34677 (N_34677,N_26917,N_28802);
and U34678 (N_34678,N_26859,N_27631);
and U34679 (N_34679,N_28184,N_22622);
nor U34680 (N_34680,N_23614,N_21210);
or U34681 (N_34681,N_22547,N_26361);
nor U34682 (N_34682,N_23972,N_22504);
and U34683 (N_34683,N_21626,N_23716);
or U34684 (N_34684,N_26507,N_21051);
xnor U34685 (N_34685,N_26755,N_27269);
or U34686 (N_34686,N_20545,N_20853);
or U34687 (N_34687,N_24722,N_25310);
nor U34688 (N_34688,N_28697,N_21900);
nor U34689 (N_34689,N_20513,N_20652);
or U34690 (N_34690,N_21236,N_28897);
nand U34691 (N_34691,N_23417,N_27876);
or U34692 (N_34692,N_24223,N_25888);
nand U34693 (N_34693,N_21233,N_22480);
and U34694 (N_34694,N_27973,N_21779);
nand U34695 (N_34695,N_28232,N_21901);
and U34696 (N_34696,N_28257,N_21673);
and U34697 (N_34697,N_23101,N_22863);
nor U34698 (N_34698,N_22451,N_26938);
nand U34699 (N_34699,N_29551,N_20609);
and U34700 (N_34700,N_29231,N_24238);
or U34701 (N_34701,N_29516,N_24721);
xor U34702 (N_34702,N_26327,N_24955);
or U34703 (N_34703,N_25170,N_25442);
nor U34704 (N_34704,N_27841,N_24419);
and U34705 (N_34705,N_28879,N_26494);
or U34706 (N_34706,N_27632,N_24568);
or U34707 (N_34707,N_27137,N_28537);
nor U34708 (N_34708,N_21029,N_27687);
nor U34709 (N_34709,N_23703,N_25235);
nand U34710 (N_34710,N_28928,N_20457);
and U34711 (N_34711,N_23001,N_20694);
xnor U34712 (N_34712,N_22563,N_27339);
or U34713 (N_34713,N_20193,N_26389);
nor U34714 (N_34714,N_22682,N_25646);
and U34715 (N_34715,N_20647,N_29377);
nor U34716 (N_34716,N_21614,N_22426);
nor U34717 (N_34717,N_21146,N_29966);
nor U34718 (N_34718,N_25967,N_22928);
xnor U34719 (N_34719,N_22779,N_22924);
nor U34720 (N_34720,N_23805,N_21822);
nand U34721 (N_34721,N_22357,N_21223);
nor U34722 (N_34722,N_20155,N_29066);
and U34723 (N_34723,N_29406,N_21600);
nor U34724 (N_34724,N_22494,N_24715);
nand U34725 (N_34725,N_25838,N_24818);
nor U34726 (N_34726,N_20401,N_21833);
nor U34727 (N_34727,N_29402,N_20908);
and U34728 (N_34728,N_21802,N_20980);
and U34729 (N_34729,N_25108,N_20806);
or U34730 (N_34730,N_28155,N_23371);
nor U34731 (N_34731,N_23612,N_24831);
xor U34732 (N_34732,N_29914,N_25981);
and U34733 (N_34733,N_23531,N_23951);
or U34734 (N_34734,N_25534,N_28444);
nor U34735 (N_34735,N_20267,N_25343);
nand U34736 (N_34736,N_23282,N_23435);
and U34737 (N_34737,N_25105,N_23002);
nand U34738 (N_34738,N_21932,N_28210);
nand U34739 (N_34739,N_29647,N_24562);
xor U34740 (N_34740,N_27693,N_28000);
nor U34741 (N_34741,N_24260,N_22741);
and U34742 (N_34742,N_27530,N_25819);
xor U34743 (N_34743,N_24985,N_25172);
nand U34744 (N_34744,N_22707,N_27156);
and U34745 (N_34745,N_20174,N_25620);
and U34746 (N_34746,N_22834,N_26942);
xor U34747 (N_34747,N_23891,N_23213);
nor U34748 (N_34748,N_29485,N_26818);
xnor U34749 (N_34749,N_26730,N_21856);
nor U34750 (N_34750,N_26176,N_21811);
xor U34751 (N_34751,N_27939,N_26775);
nor U34752 (N_34752,N_29819,N_27518);
and U34753 (N_34753,N_20117,N_28484);
and U34754 (N_34754,N_20514,N_29508);
or U34755 (N_34755,N_28583,N_25247);
or U34756 (N_34756,N_23741,N_24269);
and U34757 (N_34757,N_20765,N_21728);
nor U34758 (N_34758,N_25269,N_20326);
nor U34759 (N_34759,N_23947,N_23850);
nand U34760 (N_34760,N_28063,N_20306);
and U34761 (N_34761,N_29468,N_22272);
xnor U34762 (N_34762,N_20263,N_29294);
nor U34763 (N_34763,N_29733,N_29179);
nand U34764 (N_34764,N_29163,N_22832);
and U34765 (N_34765,N_20543,N_27372);
and U34766 (N_34766,N_28626,N_23709);
and U34767 (N_34767,N_22657,N_29379);
and U34768 (N_34768,N_23763,N_27491);
nor U34769 (N_34769,N_24728,N_20332);
nand U34770 (N_34770,N_29985,N_28046);
or U34771 (N_34771,N_22831,N_26380);
nand U34772 (N_34772,N_24036,N_29621);
nor U34773 (N_34773,N_21073,N_21375);
nor U34774 (N_34774,N_20604,N_20491);
nand U34775 (N_34775,N_28373,N_24376);
and U34776 (N_34776,N_24953,N_28707);
and U34777 (N_34777,N_25785,N_26106);
nand U34778 (N_34778,N_28813,N_29614);
xor U34779 (N_34779,N_23768,N_22141);
nor U34780 (N_34780,N_29407,N_29737);
nor U34781 (N_34781,N_27873,N_28111);
or U34782 (N_34782,N_21256,N_28934);
nor U34783 (N_34783,N_28325,N_25320);
nor U34784 (N_34784,N_25469,N_29442);
nor U34785 (N_34785,N_27484,N_23323);
nand U34786 (N_34786,N_22280,N_27454);
nand U34787 (N_34787,N_26698,N_23650);
and U34788 (N_34788,N_23968,N_28322);
nand U34789 (N_34789,N_24490,N_27214);
nand U34790 (N_34790,N_21321,N_20593);
or U34791 (N_34791,N_25221,N_21905);
nand U34792 (N_34792,N_21418,N_28487);
and U34793 (N_34793,N_25506,N_24528);
xnor U34794 (N_34794,N_29283,N_23387);
or U34795 (N_34795,N_20462,N_22795);
or U34796 (N_34796,N_27395,N_25027);
nand U34797 (N_34797,N_22778,N_24511);
nor U34798 (N_34798,N_21265,N_22988);
or U34799 (N_34799,N_29974,N_21353);
and U34800 (N_34800,N_20410,N_24069);
or U34801 (N_34801,N_21644,N_28984);
nand U34802 (N_34802,N_28082,N_27371);
and U34803 (N_34803,N_20190,N_22090);
or U34804 (N_34804,N_29762,N_21012);
and U34805 (N_34805,N_25175,N_21643);
or U34806 (N_34806,N_26045,N_25793);
and U34807 (N_34807,N_24853,N_28397);
nand U34808 (N_34808,N_27010,N_26650);
nand U34809 (N_34809,N_23374,N_25360);
nor U34810 (N_34810,N_22942,N_26677);
xor U34811 (N_34811,N_27713,N_26449);
nand U34812 (N_34812,N_21912,N_25748);
nor U34813 (N_34813,N_21011,N_25926);
and U34814 (N_34814,N_28402,N_27056);
or U34815 (N_34815,N_21488,N_23987);
and U34816 (N_34816,N_29836,N_29827);
xor U34817 (N_34817,N_26024,N_26366);
or U34818 (N_34818,N_24495,N_28927);
or U34819 (N_34819,N_23748,N_26605);
or U34820 (N_34820,N_21411,N_24844);
nand U34821 (N_34821,N_24991,N_22586);
xor U34822 (N_34822,N_29722,N_26857);
nor U34823 (N_34823,N_27401,N_22902);
and U34824 (N_34824,N_27989,N_22467);
or U34825 (N_34825,N_21428,N_25163);
or U34826 (N_34826,N_28627,N_20591);
or U34827 (N_34827,N_20073,N_21522);
nand U34828 (N_34828,N_20374,N_27665);
nand U34829 (N_34829,N_21988,N_28609);
and U34830 (N_34830,N_22676,N_22210);
or U34831 (N_34831,N_24993,N_26411);
xor U34832 (N_34832,N_29983,N_20555);
xor U34833 (N_34833,N_20076,N_21536);
or U34834 (N_34834,N_26613,N_21789);
xnor U34835 (N_34835,N_26474,N_23020);
nor U34836 (N_34836,N_23657,N_21354);
nor U34837 (N_34837,N_27981,N_23806);
or U34838 (N_34838,N_29285,N_22058);
nor U34839 (N_34839,N_21841,N_23237);
nand U34840 (N_34840,N_22871,N_20212);
or U34841 (N_34841,N_22055,N_21681);
nand U34842 (N_34842,N_28134,N_24632);
or U34843 (N_34843,N_29014,N_24718);
nand U34844 (N_34844,N_26149,N_20214);
nand U34845 (N_34845,N_25381,N_27256);
or U34846 (N_34846,N_28413,N_25625);
nor U34847 (N_34847,N_23692,N_21585);
or U34848 (N_34848,N_26645,N_26232);
nand U34849 (N_34849,N_29525,N_29470);
and U34850 (N_34850,N_25191,N_27292);
nor U34851 (N_34851,N_22246,N_23050);
nand U34852 (N_34852,N_27597,N_28331);
or U34853 (N_34853,N_28020,N_25390);
and U34854 (N_34854,N_23253,N_27595);
xor U34855 (N_34855,N_21612,N_21532);
xor U34856 (N_34856,N_29658,N_27964);
or U34857 (N_34857,N_27142,N_25770);
or U34858 (N_34858,N_21954,N_25700);
nand U34859 (N_34859,N_28923,N_21772);
or U34860 (N_34860,N_29519,N_21839);
nor U34861 (N_34861,N_24957,N_21102);
nor U34862 (N_34862,N_20503,N_24904);
xnor U34863 (N_34863,N_24460,N_28702);
nand U34864 (N_34864,N_22546,N_28871);
or U34865 (N_34865,N_27457,N_26094);
or U34866 (N_34866,N_28417,N_24645);
and U34867 (N_34867,N_25251,N_20574);
and U34868 (N_34868,N_22939,N_25708);
and U34869 (N_34869,N_25289,N_21502);
nand U34870 (N_34870,N_20506,N_29731);
nand U34871 (N_34871,N_27935,N_26455);
nor U34872 (N_34872,N_26428,N_21843);
or U34873 (N_34873,N_21874,N_27332);
and U34874 (N_34874,N_24652,N_27940);
nor U34875 (N_34875,N_29705,N_26302);
and U34876 (N_34876,N_28513,N_24686);
nor U34877 (N_34877,N_29590,N_23540);
nand U34878 (N_34878,N_23992,N_25937);
or U34879 (N_34879,N_21262,N_20066);
and U34880 (N_34880,N_28943,N_20634);
and U34881 (N_34881,N_29233,N_27316);
and U34882 (N_34882,N_20017,N_26675);
or U34883 (N_34883,N_21455,N_24272);
and U34884 (N_34884,N_28559,N_23340);
nand U34885 (N_34885,N_23023,N_22645);
xnor U34886 (N_34886,N_28741,N_24930);
nor U34887 (N_34887,N_20352,N_29041);
and U34888 (N_34888,N_20702,N_24467);
nand U34889 (N_34889,N_20235,N_28613);
and U34890 (N_34890,N_29331,N_29147);
nor U34891 (N_34891,N_29640,N_20298);
xnor U34892 (N_34892,N_28717,N_26722);
or U34893 (N_34893,N_23294,N_26011);
nand U34894 (N_34894,N_26167,N_23835);
nor U34895 (N_34895,N_20940,N_20110);
nand U34896 (N_34896,N_28216,N_27810);
or U34897 (N_34897,N_29806,N_26501);
nand U34898 (N_34898,N_24765,N_24723);
and U34899 (N_34899,N_23361,N_25528);
nand U34900 (N_34900,N_25183,N_27185);
and U34901 (N_34901,N_23032,N_29770);
nor U34902 (N_34902,N_20761,N_27829);
nor U34903 (N_34903,N_20454,N_21136);
nand U34904 (N_34904,N_26068,N_29209);
or U34905 (N_34905,N_24097,N_26910);
or U34906 (N_34906,N_22330,N_27065);
or U34907 (N_34907,N_29571,N_23327);
nand U34908 (N_34908,N_24394,N_24616);
nor U34909 (N_34909,N_23611,N_28040);
nor U34910 (N_34910,N_26436,N_29355);
xor U34911 (N_34911,N_25164,N_24217);
and U34912 (N_34912,N_27188,N_25578);
and U34913 (N_34913,N_21749,N_26493);
xnor U34914 (N_34914,N_22350,N_26544);
nor U34915 (N_34915,N_29848,N_28838);
nor U34916 (N_34916,N_21759,N_25352);
or U34917 (N_34917,N_20786,N_23918);
nor U34918 (N_34918,N_25031,N_23027);
or U34919 (N_34919,N_27621,N_29330);
nor U34920 (N_34920,N_22243,N_27282);
or U34921 (N_34921,N_29961,N_26392);
and U34922 (N_34922,N_21640,N_25796);
and U34923 (N_34923,N_24896,N_21211);
and U34924 (N_34924,N_29328,N_27916);
xnor U34925 (N_34925,N_24009,N_29024);
and U34926 (N_34926,N_25299,N_21045);
nand U34927 (N_34927,N_20469,N_22648);
or U34928 (N_34928,N_26219,N_21920);
or U34929 (N_34929,N_21117,N_25570);
and U34930 (N_34930,N_21660,N_29832);
and U34931 (N_34931,N_20817,N_25592);
nor U34932 (N_34932,N_27923,N_27516);
nor U34933 (N_34933,N_27653,N_21053);
or U34934 (N_34934,N_27291,N_22416);
nand U34935 (N_34935,N_26108,N_22833);
nand U34936 (N_34936,N_20682,N_27828);
or U34937 (N_34937,N_25083,N_29205);
nand U34938 (N_34938,N_25386,N_27335);
nand U34939 (N_34939,N_23864,N_21015);
and U34940 (N_34940,N_29155,N_21080);
nand U34941 (N_34941,N_21195,N_20411);
or U34942 (N_34942,N_21902,N_21217);
or U34943 (N_34943,N_25585,N_28305);
nand U34944 (N_34944,N_22569,N_22785);
nor U34945 (N_34945,N_25470,N_27694);
xor U34946 (N_34946,N_29298,N_26299);
and U34947 (N_34947,N_23262,N_20044);
nor U34948 (N_34948,N_26295,N_22944);
nor U34949 (N_34949,N_22287,N_24513);
nand U34950 (N_34950,N_22216,N_25774);
nand U34951 (N_34951,N_21283,N_27863);
nand U34952 (N_34952,N_29102,N_29925);
nor U34953 (N_34953,N_29080,N_23858);
or U34954 (N_34954,N_26969,N_26322);
or U34955 (N_34955,N_21235,N_25441);
nor U34956 (N_34956,N_24225,N_25082);
and U34957 (N_34957,N_22459,N_25358);
nand U34958 (N_34958,N_24640,N_24706);
or U34959 (N_34959,N_24852,N_29237);
nand U34960 (N_34960,N_27948,N_20701);
or U34961 (N_34961,N_29043,N_28823);
nor U34962 (N_34962,N_27198,N_27914);
nor U34963 (N_34963,N_21831,N_26498);
xor U34964 (N_34964,N_24201,N_27555);
nor U34965 (N_34965,N_22247,N_23370);
nand U34966 (N_34966,N_25273,N_21546);
nand U34967 (N_34967,N_21791,N_21790);
and U34968 (N_34968,N_22520,N_23203);
or U34969 (N_34969,N_21974,N_27585);
nor U34970 (N_34970,N_20343,N_25724);
nand U34971 (N_34971,N_26993,N_25674);
or U34972 (N_34972,N_28701,N_22112);
or U34973 (N_34973,N_27473,N_29973);
or U34974 (N_34974,N_22724,N_29697);
nor U34975 (N_34975,N_23406,N_20832);
and U34976 (N_34976,N_29464,N_27540);
or U34977 (N_34977,N_26586,N_26472);
or U34978 (N_34978,N_29042,N_26246);
or U34979 (N_34979,N_27704,N_25594);
nor U34980 (N_34980,N_20912,N_24893);
and U34981 (N_34981,N_27588,N_27397);
and U34982 (N_34982,N_20305,N_23745);
and U34983 (N_34983,N_21106,N_28521);
nor U34984 (N_34984,N_21251,N_22181);
xnor U34985 (N_34985,N_23065,N_26311);
nor U34986 (N_34986,N_28448,N_24001);
and U34987 (N_34987,N_27569,N_29901);
and U34988 (N_34988,N_21990,N_28787);
xor U34989 (N_34989,N_25260,N_27774);
xnor U34990 (N_34990,N_20894,N_28523);
nand U34991 (N_34991,N_26600,N_20803);
or U34992 (N_34992,N_29902,N_25884);
nand U34993 (N_34993,N_23780,N_28664);
nand U34994 (N_34994,N_20635,N_26661);
nor U34995 (N_34995,N_21176,N_20141);
nor U34996 (N_34996,N_20424,N_27608);
nand U34997 (N_34997,N_26240,N_28371);
nor U34998 (N_34998,N_21381,N_27730);
or U34999 (N_34999,N_23368,N_24882);
or U35000 (N_35000,N_28450,N_24424);
nand U35001 (N_35001,N_25014,N_20393);
nand U35002 (N_35002,N_29014,N_20590);
nor U35003 (N_35003,N_23262,N_25575);
nand U35004 (N_35004,N_24971,N_26778);
nand U35005 (N_35005,N_20169,N_20776);
nand U35006 (N_35006,N_26556,N_25018);
and U35007 (N_35007,N_29928,N_21840);
or U35008 (N_35008,N_27011,N_25091);
or U35009 (N_35009,N_28757,N_25933);
nor U35010 (N_35010,N_28092,N_27135);
and U35011 (N_35011,N_29944,N_25587);
or U35012 (N_35012,N_24056,N_22799);
or U35013 (N_35013,N_26678,N_21141);
nand U35014 (N_35014,N_23746,N_22816);
nand U35015 (N_35015,N_23953,N_29563);
nor U35016 (N_35016,N_23286,N_23546);
or U35017 (N_35017,N_25769,N_25923);
and U35018 (N_35018,N_26725,N_28641);
and U35019 (N_35019,N_24502,N_23713);
nor U35020 (N_35020,N_27075,N_28832);
nand U35021 (N_35021,N_20406,N_23202);
nand U35022 (N_35022,N_26585,N_20642);
nor U35023 (N_35023,N_24542,N_28039);
nand U35024 (N_35024,N_22125,N_29806);
or U35025 (N_35025,N_22227,N_22286);
nor U35026 (N_35026,N_27331,N_24309);
or U35027 (N_35027,N_28446,N_28730);
and U35028 (N_35028,N_23556,N_25425);
xor U35029 (N_35029,N_24017,N_26074);
or U35030 (N_35030,N_29556,N_22486);
nand U35031 (N_35031,N_22779,N_26980);
or U35032 (N_35032,N_23480,N_22446);
and U35033 (N_35033,N_22737,N_27959);
xor U35034 (N_35034,N_22669,N_28466);
or U35035 (N_35035,N_23463,N_23464);
nor U35036 (N_35036,N_23591,N_27992);
and U35037 (N_35037,N_20931,N_26328);
nand U35038 (N_35038,N_25029,N_23511);
nor U35039 (N_35039,N_25023,N_20220);
nor U35040 (N_35040,N_21939,N_21535);
and U35041 (N_35041,N_26274,N_26412);
xor U35042 (N_35042,N_22605,N_25712);
and U35043 (N_35043,N_26107,N_24879);
or U35044 (N_35044,N_20728,N_24808);
xor U35045 (N_35045,N_28809,N_26876);
and U35046 (N_35046,N_25179,N_23382);
or U35047 (N_35047,N_24462,N_23029);
nor U35048 (N_35048,N_24740,N_29957);
or U35049 (N_35049,N_25485,N_21293);
nand U35050 (N_35050,N_25399,N_20779);
nand U35051 (N_35051,N_20900,N_21701);
nor U35052 (N_35052,N_28637,N_26302);
xnor U35053 (N_35053,N_20764,N_23907);
xnor U35054 (N_35054,N_27849,N_25973);
or U35055 (N_35055,N_21184,N_20512);
xor U35056 (N_35056,N_24675,N_21331);
and U35057 (N_35057,N_26805,N_21280);
and U35058 (N_35058,N_28265,N_21521);
and U35059 (N_35059,N_22811,N_26341);
xor U35060 (N_35060,N_28088,N_24509);
nor U35061 (N_35061,N_28346,N_24584);
and U35062 (N_35062,N_25875,N_22737);
and U35063 (N_35063,N_24867,N_24719);
and U35064 (N_35064,N_27717,N_29295);
or U35065 (N_35065,N_25401,N_25753);
nor U35066 (N_35066,N_27066,N_26973);
nor U35067 (N_35067,N_20156,N_22876);
nand U35068 (N_35068,N_25786,N_20227);
nor U35069 (N_35069,N_21290,N_21577);
nor U35070 (N_35070,N_21891,N_29301);
xor U35071 (N_35071,N_22028,N_27838);
or U35072 (N_35072,N_21184,N_27552);
and U35073 (N_35073,N_28212,N_21231);
or U35074 (N_35074,N_25559,N_27163);
nand U35075 (N_35075,N_28150,N_20101);
or U35076 (N_35076,N_27608,N_20447);
nor U35077 (N_35077,N_27397,N_28455);
nor U35078 (N_35078,N_24136,N_21389);
nand U35079 (N_35079,N_23985,N_29043);
and U35080 (N_35080,N_20367,N_22093);
xor U35081 (N_35081,N_23423,N_21428);
or U35082 (N_35082,N_23314,N_29914);
and U35083 (N_35083,N_27650,N_23437);
and U35084 (N_35084,N_28965,N_23739);
or U35085 (N_35085,N_21182,N_23097);
or U35086 (N_35086,N_28463,N_23627);
nor U35087 (N_35087,N_25510,N_21811);
nor U35088 (N_35088,N_25042,N_20662);
nor U35089 (N_35089,N_29016,N_22611);
nor U35090 (N_35090,N_25310,N_26629);
or U35091 (N_35091,N_21446,N_27249);
nand U35092 (N_35092,N_21330,N_21084);
nor U35093 (N_35093,N_29588,N_28349);
xnor U35094 (N_35094,N_20647,N_22071);
nor U35095 (N_35095,N_27707,N_23471);
and U35096 (N_35096,N_25838,N_25883);
nand U35097 (N_35097,N_29630,N_24304);
nor U35098 (N_35098,N_26343,N_25280);
nor U35099 (N_35099,N_27128,N_20300);
nand U35100 (N_35100,N_29918,N_20237);
or U35101 (N_35101,N_24356,N_23207);
or U35102 (N_35102,N_20689,N_25722);
and U35103 (N_35103,N_24893,N_27014);
and U35104 (N_35104,N_24856,N_23319);
xor U35105 (N_35105,N_20197,N_23218);
nand U35106 (N_35106,N_23043,N_29080);
nand U35107 (N_35107,N_23868,N_29740);
nand U35108 (N_35108,N_21588,N_22357);
and U35109 (N_35109,N_23640,N_28769);
xor U35110 (N_35110,N_28014,N_21281);
nor U35111 (N_35111,N_25507,N_29601);
and U35112 (N_35112,N_28772,N_25549);
xnor U35113 (N_35113,N_29826,N_27984);
nor U35114 (N_35114,N_29208,N_22096);
and U35115 (N_35115,N_24303,N_28057);
nor U35116 (N_35116,N_27510,N_25308);
and U35117 (N_35117,N_22659,N_21327);
nor U35118 (N_35118,N_27490,N_20462);
nand U35119 (N_35119,N_25884,N_29207);
nand U35120 (N_35120,N_22183,N_25759);
nand U35121 (N_35121,N_25285,N_29498);
or U35122 (N_35122,N_24464,N_22089);
or U35123 (N_35123,N_23703,N_29736);
nand U35124 (N_35124,N_24666,N_27780);
and U35125 (N_35125,N_26243,N_26009);
and U35126 (N_35126,N_24844,N_27437);
nor U35127 (N_35127,N_23281,N_20644);
nor U35128 (N_35128,N_28659,N_27971);
nor U35129 (N_35129,N_29580,N_26898);
or U35130 (N_35130,N_27918,N_27880);
xnor U35131 (N_35131,N_28015,N_24059);
nand U35132 (N_35132,N_25954,N_27035);
nor U35133 (N_35133,N_23230,N_21221);
nand U35134 (N_35134,N_26440,N_22173);
xor U35135 (N_35135,N_29337,N_25569);
or U35136 (N_35136,N_24014,N_25011);
nand U35137 (N_35137,N_21115,N_26697);
xor U35138 (N_35138,N_22972,N_21322);
and U35139 (N_35139,N_20088,N_21723);
nand U35140 (N_35140,N_27242,N_26103);
nor U35141 (N_35141,N_29023,N_29365);
xnor U35142 (N_35142,N_21688,N_23952);
xnor U35143 (N_35143,N_23601,N_25421);
and U35144 (N_35144,N_27719,N_28144);
nand U35145 (N_35145,N_27683,N_25859);
and U35146 (N_35146,N_26901,N_20842);
or U35147 (N_35147,N_24693,N_26692);
nand U35148 (N_35148,N_25479,N_21752);
nand U35149 (N_35149,N_20973,N_22721);
and U35150 (N_35150,N_23077,N_28731);
nor U35151 (N_35151,N_28904,N_28653);
or U35152 (N_35152,N_21544,N_25806);
nor U35153 (N_35153,N_24202,N_29351);
and U35154 (N_35154,N_23272,N_27055);
nor U35155 (N_35155,N_20646,N_21702);
xnor U35156 (N_35156,N_29390,N_27102);
nor U35157 (N_35157,N_23272,N_29200);
and U35158 (N_35158,N_23581,N_23201);
nand U35159 (N_35159,N_28155,N_27727);
or U35160 (N_35160,N_26077,N_22203);
and U35161 (N_35161,N_28463,N_26018);
and U35162 (N_35162,N_29223,N_29010);
or U35163 (N_35163,N_29350,N_20722);
and U35164 (N_35164,N_23714,N_26161);
nor U35165 (N_35165,N_20585,N_28471);
or U35166 (N_35166,N_24702,N_24693);
nor U35167 (N_35167,N_28754,N_20144);
or U35168 (N_35168,N_29835,N_26612);
or U35169 (N_35169,N_23055,N_21990);
nand U35170 (N_35170,N_23717,N_24108);
nor U35171 (N_35171,N_26210,N_28973);
or U35172 (N_35172,N_25765,N_26375);
or U35173 (N_35173,N_27030,N_28779);
nand U35174 (N_35174,N_26267,N_22504);
nor U35175 (N_35175,N_26021,N_25170);
xnor U35176 (N_35176,N_22593,N_22552);
nand U35177 (N_35177,N_24218,N_21707);
nand U35178 (N_35178,N_20520,N_28700);
or U35179 (N_35179,N_23726,N_23120);
xor U35180 (N_35180,N_25768,N_24732);
or U35181 (N_35181,N_20491,N_29944);
xnor U35182 (N_35182,N_28162,N_27692);
nor U35183 (N_35183,N_24295,N_23570);
nand U35184 (N_35184,N_25122,N_26947);
and U35185 (N_35185,N_26282,N_28732);
and U35186 (N_35186,N_24499,N_26278);
xor U35187 (N_35187,N_26829,N_25348);
nand U35188 (N_35188,N_23959,N_25898);
nor U35189 (N_35189,N_24823,N_21303);
and U35190 (N_35190,N_22762,N_29976);
xnor U35191 (N_35191,N_23528,N_22047);
or U35192 (N_35192,N_22609,N_26648);
and U35193 (N_35193,N_20958,N_27457);
nand U35194 (N_35194,N_20479,N_20829);
and U35195 (N_35195,N_21985,N_22445);
nor U35196 (N_35196,N_21181,N_21714);
nand U35197 (N_35197,N_28561,N_24144);
nand U35198 (N_35198,N_21729,N_20187);
nand U35199 (N_35199,N_23906,N_25023);
nand U35200 (N_35200,N_27283,N_27417);
nor U35201 (N_35201,N_21270,N_29602);
nand U35202 (N_35202,N_23072,N_23887);
and U35203 (N_35203,N_28969,N_25421);
and U35204 (N_35204,N_21580,N_29050);
nor U35205 (N_35205,N_20207,N_20163);
or U35206 (N_35206,N_23284,N_24646);
or U35207 (N_35207,N_21778,N_21608);
nor U35208 (N_35208,N_21432,N_29677);
xnor U35209 (N_35209,N_23683,N_20416);
or U35210 (N_35210,N_29698,N_20677);
nand U35211 (N_35211,N_28945,N_29572);
nand U35212 (N_35212,N_24310,N_28128);
or U35213 (N_35213,N_24816,N_25252);
nand U35214 (N_35214,N_29175,N_26039);
and U35215 (N_35215,N_27634,N_20396);
and U35216 (N_35216,N_20736,N_28074);
and U35217 (N_35217,N_25298,N_28584);
nand U35218 (N_35218,N_21400,N_29887);
nand U35219 (N_35219,N_24442,N_20588);
nand U35220 (N_35220,N_22506,N_28724);
and U35221 (N_35221,N_25687,N_26351);
nand U35222 (N_35222,N_27779,N_27141);
or U35223 (N_35223,N_28783,N_23774);
xnor U35224 (N_35224,N_25138,N_21252);
and U35225 (N_35225,N_28147,N_21470);
and U35226 (N_35226,N_25887,N_22460);
or U35227 (N_35227,N_24505,N_28189);
or U35228 (N_35228,N_21744,N_28544);
nor U35229 (N_35229,N_26010,N_27959);
nor U35230 (N_35230,N_23150,N_21503);
or U35231 (N_35231,N_24526,N_22513);
nand U35232 (N_35232,N_21152,N_22687);
xor U35233 (N_35233,N_29976,N_20940);
and U35234 (N_35234,N_21442,N_27571);
nand U35235 (N_35235,N_29459,N_26416);
nand U35236 (N_35236,N_26733,N_23543);
nand U35237 (N_35237,N_20635,N_29810);
or U35238 (N_35238,N_25325,N_20298);
and U35239 (N_35239,N_21849,N_22800);
and U35240 (N_35240,N_25663,N_28570);
nand U35241 (N_35241,N_22195,N_22250);
nand U35242 (N_35242,N_21527,N_25517);
and U35243 (N_35243,N_26457,N_20013);
xnor U35244 (N_35244,N_21203,N_25382);
nor U35245 (N_35245,N_22637,N_29721);
and U35246 (N_35246,N_29188,N_21263);
or U35247 (N_35247,N_28021,N_21979);
and U35248 (N_35248,N_27878,N_23036);
xnor U35249 (N_35249,N_26990,N_20286);
and U35250 (N_35250,N_22148,N_25560);
nor U35251 (N_35251,N_22663,N_25753);
xor U35252 (N_35252,N_20115,N_25784);
nor U35253 (N_35253,N_27690,N_21693);
nand U35254 (N_35254,N_27126,N_22552);
nand U35255 (N_35255,N_28075,N_23722);
and U35256 (N_35256,N_26556,N_25963);
xnor U35257 (N_35257,N_29893,N_27214);
nor U35258 (N_35258,N_20041,N_27377);
nand U35259 (N_35259,N_25122,N_28691);
and U35260 (N_35260,N_26890,N_20881);
nor U35261 (N_35261,N_23481,N_25142);
or U35262 (N_35262,N_29289,N_24366);
and U35263 (N_35263,N_24547,N_29781);
xor U35264 (N_35264,N_25700,N_20096);
and U35265 (N_35265,N_23695,N_27802);
or U35266 (N_35266,N_20338,N_24477);
nor U35267 (N_35267,N_29224,N_25508);
and U35268 (N_35268,N_21548,N_24261);
xor U35269 (N_35269,N_28918,N_24603);
or U35270 (N_35270,N_29912,N_27390);
xor U35271 (N_35271,N_29650,N_20762);
nand U35272 (N_35272,N_21051,N_24300);
and U35273 (N_35273,N_24919,N_22394);
nand U35274 (N_35274,N_22177,N_28669);
and U35275 (N_35275,N_24803,N_27956);
nor U35276 (N_35276,N_29884,N_29239);
or U35277 (N_35277,N_22668,N_23737);
nor U35278 (N_35278,N_26563,N_21700);
and U35279 (N_35279,N_23517,N_28537);
nand U35280 (N_35280,N_29156,N_29209);
nor U35281 (N_35281,N_24871,N_23361);
nor U35282 (N_35282,N_27912,N_27260);
nand U35283 (N_35283,N_23954,N_24774);
nor U35284 (N_35284,N_26849,N_24237);
and U35285 (N_35285,N_25001,N_26280);
nand U35286 (N_35286,N_25157,N_26885);
xor U35287 (N_35287,N_23370,N_26998);
xnor U35288 (N_35288,N_26385,N_20150);
xor U35289 (N_35289,N_24146,N_21790);
and U35290 (N_35290,N_27100,N_25078);
and U35291 (N_35291,N_22315,N_29179);
or U35292 (N_35292,N_20155,N_26950);
and U35293 (N_35293,N_24858,N_29546);
nor U35294 (N_35294,N_26473,N_28579);
or U35295 (N_35295,N_28837,N_20969);
or U35296 (N_35296,N_29182,N_20424);
or U35297 (N_35297,N_24880,N_27632);
or U35298 (N_35298,N_21006,N_23052);
nand U35299 (N_35299,N_20720,N_25402);
nor U35300 (N_35300,N_24216,N_28964);
and U35301 (N_35301,N_26277,N_23604);
or U35302 (N_35302,N_24176,N_21302);
and U35303 (N_35303,N_25850,N_26859);
nor U35304 (N_35304,N_21342,N_26879);
nor U35305 (N_35305,N_21786,N_29918);
nand U35306 (N_35306,N_21702,N_20892);
nor U35307 (N_35307,N_24988,N_21652);
nor U35308 (N_35308,N_27994,N_29164);
and U35309 (N_35309,N_25551,N_29073);
or U35310 (N_35310,N_24132,N_23235);
or U35311 (N_35311,N_23202,N_21188);
nor U35312 (N_35312,N_24175,N_22722);
nand U35313 (N_35313,N_28527,N_25367);
or U35314 (N_35314,N_21064,N_28858);
nand U35315 (N_35315,N_29331,N_26427);
nand U35316 (N_35316,N_27379,N_29093);
or U35317 (N_35317,N_26541,N_20430);
nor U35318 (N_35318,N_25728,N_26276);
nor U35319 (N_35319,N_27049,N_21329);
nand U35320 (N_35320,N_24340,N_22702);
or U35321 (N_35321,N_22422,N_29405);
or U35322 (N_35322,N_20618,N_23170);
nor U35323 (N_35323,N_26710,N_29066);
nand U35324 (N_35324,N_22518,N_23401);
nor U35325 (N_35325,N_29119,N_27244);
nor U35326 (N_35326,N_22675,N_29051);
nand U35327 (N_35327,N_24464,N_20140);
or U35328 (N_35328,N_24905,N_22942);
nor U35329 (N_35329,N_22887,N_23990);
nand U35330 (N_35330,N_25660,N_24089);
nand U35331 (N_35331,N_24752,N_26975);
xnor U35332 (N_35332,N_23505,N_26907);
nand U35333 (N_35333,N_29311,N_29602);
nor U35334 (N_35334,N_25025,N_27750);
or U35335 (N_35335,N_29442,N_29874);
or U35336 (N_35336,N_27948,N_28888);
nand U35337 (N_35337,N_23399,N_27822);
or U35338 (N_35338,N_20877,N_21857);
and U35339 (N_35339,N_20320,N_21267);
nand U35340 (N_35340,N_25409,N_28966);
and U35341 (N_35341,N_22749,N_27564);
and U35342 (N_35342,N_27243,N_21910);
nand U35343 (N_35343,N_26265,N_26800);
or U35344 (N_35344,N_28671,N_27075);
xnor U35345 (N_35345,N_24470,N_26597);
or U35346 (N_35346,N_20438,N_23614);
nor U35347 (N_35347,N_28853,N_26884);
nor U35348 (N_35348,N_25425,N_23125);
nor U35349 (N_35349,N_24357,N_25445);
and U35350 (N_35350,N_23149,N_22376);
nand U35351 (N_35351,N_24171,N_25081);
or U35352 (N_35352,N_28058,N_25130);
and U35353 (N_35353,N_23060,N_22218);
or U35354 (N_35354,N_26991,N_24144);
nand U35355 (N_35355,N_26361,N_26923);
and U35356 (N_35356,N_26140,N_27031);
nand U35357 (N_35357,N_21083,N_27022);
or U35358 (N_35358,N_21459,N_28486);
nand U35359 (N_35359,N_23559,N_20130);
and U35360 (N_35360,N_26381,N_20270);
nor U35361 (N_35361,N_28595,N_23829);
and U35362 (N_35362,N_22976,N_26784);
nand U35363 (N_35363,N_25171,N_29719);
and U35364 (N_35364,N_25343,N_21432);
and U35365 (N_35365,N_27193,N_21021);
nand U35366 (N_35366,N_21532,N_23539);
nand U35367 (N_35367,N_24025,N_26584);
nand U35368 (N_35368,N_22534,N_29360);
or U35369 (N_35369,N_23569,N_24894);
or U35370 (N_35370,N_27494,N_25430);
nor U35371 (N_35371,N_29988,N_25609);
or U35372 (N_35372,N_25493,N_26265);
nor U35373 (N_35373,N_20469,N_26620);
nor U35374 (N_35374,N_29522,N_23047);
and U35375 (N_35375,N_23148,N_29121);
or U35376 (N_35376,N_27836,N_21446);
or U35377 (N_35377,N_28488,N_28409);
nor U35378 (N_35378,N_29870,N_25137);
or U35379 (N_35379,N_29384,N_28604);
nand U35380 (N_35380,N_23631,N_24773);
nand U35381 (N_35381,N_23105,N_21157);
nor U35382 (N_35382,N_29327,N_20574);
or U35383 (N_35383,N_22782,N_28009);
xnor U35384 (N_35384,N_21101,N_29309);
nand U35385 (N_35385,N_28408,N_21569);
xor U35386 (N_35386,N_21564,N_26633);
and U35387 (N_35387,N_27167,N_22001);
and U35388 (N_35388,N_25541,N_24185);
xnor U35389 (N_35389,N_26863,N_25950);
or U35390 (N_35390,N_21722,N_29402);
and U35391 (N_35391,N_26918,N_22773);
nor U35392 (N_35392,N_29876,N_22156);
nor U35393 (N_35393,N_23941,N_22481);
nor U35394 (N_35394,N_22599,N_23268);
nand U35395 (N_35395,N_28101,N_23372);
nor U35396 (N_35396,N_26558,N_26286);
nor U35397 (N_35397,N_24897,N_22234);
nor U35398 (N_35398,N_22293,N_26621);
or U35399 (N_35399,N_24592,N_21553);
or U35400 (N_35400,N_25588,N_26262);
nand U35401 (N_35401,N_23849,N_29021);
xnor U35402 (N_35402,N_22653,N_22493);
nand U35403 (N_35403,N_25332,N_23397);
and U35404 (N_35404,N_25588,N_29154);
nor U35405 (N_35405,N_26953,N_23782);
nand U35406 (N_35406,N_20372,N_22900);
nor U35407 (N_35407,N_26737,N_29756);
nor U35408 (N_35408,N_29186,N_23613);
or U35409 (N_35409,N_21831,N_20465);
xor U35410 (N_35410,N_27619,N_21739);
nor U35411 (N_35411,N_28379,N_27031);
nand U35412 (N_35412,N_22645,N_24887);
and U35413 (N_35413,N_26626,N_23263);
and U35414 (N_35414,N_23783,N_29443);
and U35415 (N_35415,N_27656,N_28669);
and U35416 (N_35416,N_26433,N_25035);
and U35417 (N_35417,N_26348,N_20077);
nand U35418 (N_35418,N_28170,N_25305);
nand U35419 (N_35419,N_21924,N_22316);
nand U35420 (N_35420,N_28620,N_21392);
or U35421 (N_35421,N_29698,N_20668);
xnor U35422 (N_35422,N_27664,N_26436);
nand U35423 (N_35423,N_29960,N_27653);
xor U35424 (N_35424,N_21322,N_24861);
nand U35425 (N_35425,N_20048,N_22179);
or U35426 (N_35426,N_29706,N_23461);
nor U35427 (N_35427,N_24402,N_24599);
nor U35428 (N_35428,N_21776,N_29398);
or U35429 (N_35429,N_25146,N_25491);
nand U35430 (N_35430,N_21602,N_27069);
or U35431 (N_35431,N_20491,N_26366);
nor U35432 (N_35432,N_22163,N_28708);
or U35433 (N_35433,N_23918,N_26147);
xnor U35434 (N_35434,N_29061,N_23240);
and U35435 (N_35435,N_24412,N_28343);
xor U35436 (N_35436,N_25403,N_27811);
and U35437 (N_35437,N_21654,N_29911);
or U35438 (N_35438,N_25578,N_29330);
nand U35439 (N_35439,N_20457,N_25218);
nor U35440 (N_35440,N_21193,N_25017);
or U35441 (N_35441,N_22449,N_28124);
or U35442 (N_35442,N_25094,N_21729);
and U35443 (N_35443,N_28963,N_27744);
or U35444 (N_35444,N_24970,N_20754);
nor U35445 (N_35445,N_29453,N_28371);
xor U35446 (N_35446,N_27860,N_21243);
and U35447 (N_35447,N_24123,N_27827);
or U35448 (N_35448,N_29531,N_29780);
and U35449 (N_35449,N_28155,N_28254);
nor U35450 (N_35450,N_28421,N_21854);
nor U35451 (N_35451,N_26430,N_21447);
xor U35452 (N_35452,N_24082,N_26828);
and U35453 (N_35453,N_21352,N_22452);
nand U35454 (N_35454,N_24835,N_20728);
xor U35455 (N_35455,N_29848,N_26425);
and U35456 (N_35456,N_26255,N_21683);
or U35457 (N_35457,N_29251,N_26990);
or U35458 (N_35458,N_25236,N_28459);
or U35459 (N_35459,N_25482,N_24192);
or U35460 (N_35460,N_23136,N_22131);
and U35461 (N_35461,N_28708,N_26847);
or U35462 (N_35462,N_29038,N_27390);
nor U35463 (N_35463,N_23741,N_26376);
or U35464 (N_35464,N_23834,N_21367);
nor U35465 (N_35465,N_20482,N_21672);
nand U35466 (N_35466,N_28257,N_21770);
and U35467 (N_35467,N_23509,N_28409);
and U35468 (N_35468,N_23436,N_21671);
and U35469 (N_35469,N_25279,N_27066);
nand U35470 (N_35470,N_20380,N_29692);
nand U35471 (N_35471,N_24769,N_22883);
and U35472 (N_35472,N_24138,N_21284);
or U35473 (N_35473,N_24269,N_24387);
or U35474 (N_35474,N_24825,N_26874);
or U35475 (N_35475,N_24217,N_29517);
xor U35476 (N_35476,N_29338,N_22144);
or U35477 (N_35477,N_23423,N_26401);
nand U35478 (N_35478,N_24718,N_24414);
and U35479 (N_35479,N_26507,N_25315);
and U35480 (N_35480,N_26986,N_27710);
nand U35481 (N_35481,N_26303,N_24901);
nand U35482 (N_35482,N_24271,N_26559);
or U35483 (N_35483,N_25079,N_23064);
or U35484 (N_35484,N_28499,N_22829);
and U35485 (N_35485,N_24171,N_29920);
or U35486 (N_35486,N_23104,N_29748);
nand U35487 (N_35487,N_26794,N_28636);
nor U35488 (N_35488,N_21192,N_23853);
xor U35489 (N_35489,N_22008,N_21973);
nand U35490 (N_35490,N_20152,N_27448);
nor U35491 (N_35491,N_20855,N_26618);
nor U35492 (N_35492,N_28492,N_23806);
nand U35493 (N_35493,N_22918,N_21620);
nor U35494 (N_35494,N_29858,N_27708);
or U35495 (N_35495,N_20917,N_20503);
nand U35496 (N_35496,N_27246,N_24960);
xnor U35497 (N_35497,N_21828,N_23768);
or U35498 (N_35498,N_21457,N_23859);
or U35499 (N_35499,N_27939,N_21935);
or U35500 (N_35500,N_22810,N_27707);
or U35501 (N_35501,N_20005,N_28126);
nand U35502 (N_35502,N_26260,N_27831);
nand U35503 (N_35503,N_22581,N_26383);
or U35504 (N_35504,N_22470,N_26618);
and U35505 (N_35505,N_23327,N_25443);
nand U35506 (N_35506,N_29598,N_28358);
and U35507 (N_35507,N_27575,N_28461);
or U35508 (N_35508,N_27232,N_26763);
nand U35509 (N_35509,N_28652,N_22048);
xor U35510 (N_35510,N_20587,N_29103);
nor U35511 (N_35511,N_28640,N_21056);
and U35512 (N_35512,N_23550,N_27033);
or U35513 (N_35513,N_28919,N_27061);
nor U35514 (N_35514,N_26872,N_23589);
and U35515 (N_35515,N_26489,N_23890);
and U35516 (N_35516,N_24249,N_20652);
or U35517 (N_35517,N_20523,N_28062);
nand U35518 (N_35518,N_22339,N_22433);
nor U35519 (N_35519,N_24419,N_26180);
and U35520 (N_35520,N_28616,N_25855);
nand U35521 (N_35521,N_26206,N_21791);
and U35522 (N_35522,N_26299,N_20758);
xor U35523 (N_35523,N_20885,N_24776);
nor U35524 (N_35524,N_26950,N_22882);
nand U35525 (N_35525,N_29546,N_25540);
or U35526 (N_35526,N_27071,N_28324);
nor U35527 (N_35527,N_20317,N_24511);
nand U35528 (N_35528,N_22760,N_29536);
and U35529 (N_35529,N_22086,N_26314);
or U35530 (N_35530,N_24088,N_26933);
nor U35531 (N_35531,N_27462,N_29375);
nand U35532 (N_35532,N_22156,N_26782);
nor U35533 (N_35533,N_29542,N_28160);
xor U35534 (N_35534,N_25469,N_24877);
and U35535 (N_35535,N_28214,N_28373);
or U35536 (N_35536,N_26203,N_21535);
nor U35537 (N_35537,N_20993,N_29853);
or U35538 (N_35538,N_29704,N_26540);
nand U35539 (N_35539,N_24365,N_22766);
nor U35540 (N_35540,N_24725,N_29923);
nor U35541 (N_35541,N_29647,N_20555);
or U35542 (N_35542,N_29596,N_21825);
or U35543 (N_35543,N_25961,N_26686);
nand U35544 (N_35544,N_24146,N_26070);
and U35545 (N_35545,N_24932,N_25799);
and U35546 (N_35546,N_24760,N_29333);
or U35547 (N_35547,N_23478,N_23440);
nor U35548 (N_35548,N_26152,N_21856);
or U35549 (N_35549,N_23223,N_21933);
nand U35550 (N_35550,N_29214,N_25638);
and U35551 (N_35551,N_20006,N_27090);
nand U35552 (N_35552,N_28228,N_26598);
nor U35553 (N_35553,N_27599,N_25851);
or U35554 (N_35554,N_25873,N_22011);
nor U35555 (N_35555,N_27535,N_21029);
nand U35556 (N_35556,N_27247,N_23443);
nand U35557 (N_35557,N_24101,N_24068);
nor U35558 (N_35558,N_26315,N_22706);
or U35559 (N_35559,N_24735,N_24905);
xor U35560 (N_35560,N_26484,N_21389);
xnor U35561 (N_35561,N_24083,N_29573);
nor U35562 (N_35562,N_24413,N_24799);
nand U35563 (N_35563,N_26543,N_29274);
xnor U35564 (N_35564,N_22371,N_20505);
and U35565 (N_35565,N_24631,N_27421);
nand U35566 (N_35566,N_27266,N_29799);
nor U35567 (N_35567,N_24919,N_27312);
and U35568 (N_35568,N_27778,N_20892);
and U35569 (N_35569,N_21999,N_23524);
or U35570 (N_35570,N_24971,N_28249);
nand U35571 (N_35571,N_20818,N_25972);
and U35572 (N_35572,N_23183,N_28059);
or U35573 (N_35573,N_27604,N_27837);
nand U35574 (N_35574,N_25721,N_28063);
nand U35575 (N_35575,N_26735,N_28414);
nor U35576 (N_35576,N_27860,N_20450);
nor U35577 (N_35577,N_27645,N_29344);
xor U35578 (N_35578,N_23974,N_21272);
xor U35579 (N_35579,N_27766,N_24312);
or U35580 (N_35580,N_26226,N_23754);
xnor U35581 (N_35581,N_29210,N_24004);
or U35582 (N_35582,N_21058,N_26453);
nand U35583 (N_35583,N_20515,N_29212);
or U35584 (N_35584,N_28137,N_22620);
nor U35585 (N_35585,N_29033,N_23212);
and U35586 (N_35586,N_23306,N_25200);
or U35587 (N_35587,N_23639,N_22682);
or U35588 (N_35588,N_26865,N_25138);
xor U35589 (N_35589,N_27779,N_20976);
and U35590 (N_35590,N_21971,N_20137);
nand U35591 (N_35591,N_29183,N_27524);
nand U35592 (N_35592,N_20466,N_23471);
or U35593 (N_35593,N_20850,N_20212);
nand U35594 (N_35594,N_24028,N_27862);
and U35595 (N_35595,N_21277,N_28381);
nor U35596 (N_35596,N_22084,N_28799);
nand U35597 (N_35597,N_27035,N_23710);
and U35598 (N_35598,N_22033,N_23067);
or U35599 (N_35599,N_27556,N_21987);
or U35600 (N_35600,N_20568,N_27324);
and U35601 (N_35601,N_27892,N_24778);
nor U35602 (N_35602,N_24658,N_29976);
nand U35603 (N_35603,N_21637,N_25680);
nor U35604 (N_35604,N_20099,N_22412);
nand U35605 (N_35605,N_23642,N_22332);
and U35606 (N_35606,N_26052,N_27567);
nand U35607 (N_35607,N_25260,N_22113);
nor U35608 (N_35608,N_28768,N_28878);
nor U35609 (N_35609,N_25207,N_22207);
nand U35610 (N_35610,N_20201,N_25224);
nor U35611 (N_35611,N_20504,N_29301);
nand U35612 (N_35612,N_28080,N_29221);
xor U35613 (N_35613,N_22880,N_27900);
or U35614 (N_35614,N_25105,N_27588);
xnor U35615 (N_35615,N_27806,N_23683);
or U35616 (N_35616,N_27537,N_27226);
and U35617 (N_35617,N_27707,N_28678);
and U35618 (N_35618,N_20257,N_27890);
nand U35619 (N_35619,N_21498,N_29981);
nor U35620 (N_35620,N_28385,N_25581);
and U35621 (N_35621,N_22341,N_22986);
nand U35622 (N_35622,N_29182,N_21112);
nand U35623 (N_35623,N_20248,N_24749);
nor U35624 (N_35624,N_23895,N_28694);
nand U35625 (N_35625,N_28308,N_24731);
and U35626 (N_35626,N_24844,N_24489);
xnor U35627 (N_35627,N_28845,N_28344);
nor U35628 (N_35628,N_23239,N_23440);
or U35629 (N_35629,N_23876,N_25605);
nor U35630 (N_35630,N_29045,N_23670);
nand U35631 (N_35631,N_23671,N_29256);
nand U35632 (N_35632,N_21462,N_28091);
and U35633 (N_35633,N_20392,N_25322);
or U35634 (N_35634,N_28684,N_26185);
nor U35635 (N_35635,N_22995,N_29320);
or U35636 (N_35636,N_28064,N_27853);
nor U35637 (N_35637,N_25166,N_27635);
nand U35638 (N_35638,N_21160,N_23349);
nand U35639 (N_35639,N_28479,N_20180);
and U35640 (N_35640,N_26183,N_25414);
nand U35641 (N_35641,N_25627,N_25540);
nand U35642 (N_35642,N_24680,N_20725);
nand U35643 (N_35643,N_28162,N_24025);
or U35644 (N_35644,N_22494,N_23140);
and U35645 (N_35645,N_23526,N_23225);
and U35646 (N_35646,N_21422,N_25372);
nand U35647 (N_35647,N_29313,N_28421);
or U35648 (N_35648,N_26272,N_26495);
and U35649 (N_35649,N_27079,N_29528);
and U35650 (N_35650,N_22040,N_27491);
nand U35651 (N_35651,N_21397,N_26574);
xor U35652 (N_35652,N_24136,N_29035);
xnor U35653 (N_35653,N_26375,N_21962);
and U35654 (N_35654,N_22287,N_22474);
and U35655 (N_35655,N_22223,N_27789);
nand U35656 (N_35656,N_26578,N_20761);
nand U35657 (N_35657,N_23815,N_22834);
nand U35658 (N_35658,N_21230,N_26848);
nand U35659 (N_35659,N_26490,N_27635);
nor U35660 (N_35660,N_28922,N_24330);
and U35661 (N_35661,N_21354,N_22601);
and U35662 (N_35662,N_26234,N_26207);
nand U35663 (N_35663,N_28509,N_28261);
or U35664 (N_35664,N_21957,N_25229);
nand U35665 (N_35665,N_25347,N_27102);
and U35666 (N_35666,N_23685,N_25789);
xnor U35667 (N_35667,N_27522,N_27747);
nand U35668 (N_35668,N_20153,N_26781);
nand U35669 (N_35669,N_27517,N_22076);
or U35670 (N_35670,N_21018,N_25129);
or U35671 (N_35671,N_20622,N_20791);
or U35672 (N_35672,N_25295,N_28734);
or U35673 (N_35673,N_23983,N_27090);
xnor U35674 (N_35674,N_27659,N_26235);
nand U35675 (N_35675,N_28504,N_28086);
nor U35676 (N_35676,N_25610,N_26374);
nor U35677 (N_35677,N_22519,N_26040);
nand U35678 (N_35678,N_26068,N_22919);
xnor U35679 (N_35679,N_20081,N_20523);
or U35680 (N_35680,N_24041,N_28767);
nor U35681 (N_35681,N_29040,N_27812);
and U35682 (N_35682,N_25592,N_24671);
or U35683 (N_35683,N_23908,N_25130);
nor U35684 (N_35684,N_21990,N_29418);
nor U35685 (N_35685,N_28969,N_23156);
xor U35686 (N_35686,N_22270,N_22210);
nor U35687 (N_35687,N_27612,N_27487);
or U35688 (N_35688,N_27845,N_27661);
and U35689 (N_35689,N_23075,N_25790);
nor U35690 (N_35690,N_27287,N_23665);
or U35691 (N_35691,N_25771,N_20415);
and U35692 (N_35692,N_21244,N_27817);
nor U35693 (N_35693,N_29361,N_25923);
xnor U35694 (N_35694,N_27557,N_25711);
nor U35695 (N_35695,N_26930,N_22235);
nor U35696 (N_35696,N_20856,N_22919);
or U35697 (N_35697,N_25131,N_28238);
nor U35698 (N_35698,N_25345,N_25228);
and U35699 (N_35699,N_26058,N_22759);
and U35700 (N_35700,N_25224,N_29609);
and U35701 (N_35701,N_23441,N_23258);
nor U35702 (N_35702,N_26424,N_26882);
xnor U35703 (N_35703,N_25792,N_26101);
xor U35704 (N_35704,N_25784,N_22122);
nand U35705 (N_35705,N_22059,N_26753);
nand U35706 (N_35706,N_25246,N_27980);
or U35707 (N_35707,N_29761,N_29168);
and U35708 (N_35708,N_22170,N_21810);
and U35709 (N_35709,N_26028,N_29814);
or U35710 (N_35710,N_26651,N_27934);
xnor U35711 (N_35711,N_24584,N_23505);
nand U35712 (N_35712,N_20360,N_27026);
nor U35713 (N_35713,N_21559,N_25046);
nand U35714 (N_35714,N_29143,N_25190);
and U35715 (N_35715,N_26186,N_21062);
xnor U35716 (N_35716,N_29551,N_25390);
nand U35717 (N_35717,N_25174,N_25565);
and U35718 (N_35718,N_23812,N_23766);
and U35719 (N_35719,N_28753,N_23423);
nor U35720 (N_35720,N_26410,N_20129);
nand U35721 (N_35721,N_26498,N_29416);
or U35722 (N_35722,N_25755,N_28531);
nor U35723 (N_35723,N_29110,N_21088);
xnor U35724 (N_35724,N_26669,N_21471);
or U35725 (N_35725,N_22244,N_25853);
xor U35726 (N_35726,N_25463,N_23079);
and U35727 (N_35727,N_29406,N_24038);
nand U35728 (N_35728,N_20661,N_27575);
or U35729 (N_35729,N_20440,N_25313);
and U35730 (N_35730,N_27973,N_23911);
or U35731 (N_35731,N_20580,N_20532);
nand U35732 (N_35732,N_29305,N_22770);
nor U35733 (N_35733,N_24765,N_22623);
and U35734 (N_35734,N_27590,N_23650);
nor U35735 (N_35735,N_26239,N_25108);
nand U35736 (N_35736,N_29990,N_24180);
or U35737 (N_35737,N_28949,N_24001);
and U35738 (N_35738,N_27036,N_20915);
or U35739 (N_35739,N_25749,N_27996);
or U35740 (N_35740,N_22985,N_24426);
xnor U35741 (N_35741,N_28206,N_23386);
xnor U35742 (N_35742,N_24106,N_24843);
nor U35743 (N_35743,N_29543,N_23993);
or U35744 (N_35744,N_20259,N_26341);
nor U35745 (N_35745,N_20400,N_23036);
xnor U35746 (N_35746,N_20573,N_29492);
xor U35747 (N_35747,N_23065,N_27017);
and U35748 (N_35748,N_23750,N_26242);
xor U35749 (N_35749,N_26293,N_21043);
and U35750 (N_35750,N_21814,N_29798);
nand U35751 (N_35751,N_29477,N_26284);
and U35752 (N_35752,N_26579,N_29166);
nor U35753 (N_35753,N_26699,N_29336);
nor U35754 (N_35754,N_27610,N_28923);
or U35755 (N_35755,N_25718,N_21746);
nand U35756 (N_35756,N_20662,N_26968);
or U35757 (N_35757,N_27573,N_26815);
nor U35758 (N_35758,N_23999,N_29682);
or U35759 (N_35759,N_21198,N_25973);
or U35760 (N_35760,N_28888,N_20066);
or U35761 (N_35761,N_21167,N_29805);
nand U35762 (N_35762,N_29342,N_21752);
nor U35763 (N_35763,N_29936,N_28474);
and U35764 (N_35764,N_22265,N_24051);
nor U35765 (N_35765,N_24364,N_20156);
nand U35766 (N_35766,N_22668,N_24502);
or U35767 (N_35767,N_20443,N_23885);
nor U35768 (N_35768,N_21236,N_20058);
and U35769 (N_35769,N_28173,N_29549);
nor U35770 (N_35770,N_25048,N_21533);
nand U35771 (N_35771,N_28689,N_22011);
or U35772 (N_35772,N_29686,N_25650);
xnor U35773 (N_35773,N_28379,N_25378);
xnor U35774 (N_35774,N_24407,N_21813);
nand U35775 (N_35775,N_23698,N_21937);
and U35776 (N_35776,N_23779,N_27259);
nand U35777 (N_35777,N_23015,N_25222);
nor U35778 (N_35778,N_27819,N_26922);
nand U35779 (N_35779,N_22104,N_28748);
xor U35780 (N_35780,N_27544,N_21282);
nor U35781 (N_35781,N_28661,N_21053);
xor U35782 (N_35782,N_27572,N_21170);
or U35783 (N_35783,N_21823,N_28729);
nand U35784 (N_35784,N_24606,N_29058);
nor U35785 (N_35785,N_23441,N_28746);
nand U35786 (N_35786,N_21197,N_20369);
or U35787 (N_35787,N_27946,N_27134);
nor U35788 (N_35788,N_28636,N_26490);
xor U35789 (N_35789,N_22912,N_23419);
nor U35790 (N_35790,N_23756,N_27018);
and U35791 (N_35791,N_20509,N_25823);
nor U35792 (N_35792,N_28820,N_22608);
nor U35793 (N_35793,N_27986,N_21393);
nor U35794 (N_35794,N_26009,N_26745);
nor U35795 (N_35795,N_23357,N_20744);
and U35796 (N_35796,N_26502,N_27427);
xor U35797 (N_35797,N_22243,N_27635);
or U35798 (N_35798,N_27879,N_21931);
nand U35799 (N_35799,N_28152,N_20778);
and U35800 (N_35800,N_27034,N_20498);
nor U35801 (N_35801,N_22366,N_28399);
and U35802 (N_35802,N_24834,N_27085);
or U35803 (N_35803,N_28389,N_26370);
nand U35804 (N_35804,N_21894,N_24808);
nor U35805 (N_35805,N_29192,N_27099);
and U35806 (N_35806,N_29894,N_21241);
or U35807 (N_35807,N_22589,N_21816);
nor U35808 (N_35808,N_21461,N_25534);
and U35809 (N_35809,N_20252,N_21823);
nor U35810 (N_35810,N_28818,N_21006);
xnor U35811 (N_35811,N_20652,N_25103);
xor U35812 (N_35812,N_20008,N_27468);
nor U35813 (N_35813,N_27289,N_23888);
nand U35814 (N_35814,N_27239,N_21421);
nand U35815 (N_35815,N_25864,N_24435);
and U35816 (N_35816,N_22387,N_29696);
nor U35817 (N_35817,N_20934,N_29006);
nor U35818 (N_35818,N_29564,N_26499);
or U35819 (N_35819,N_24201,N_24398);
nand U35820 (N_35820,N_28240,N_22781);
nor U35821 (N_35821,N_21671,N_23254);
and U35822 (N_35822,N_25755,N_21500);
nand U35823 (N_35823,N_29595,N_25666);
nor U35824 (N_35824,N_20367,N_23155);
xor U35825 (N_35825,N_29050,N_20590);
and U35826 (N_35826,N_23272,N_22237);
or U35827 (N_35827,N_25031,N_28013);
and U35828 (N_35828,N_21793,N_26437);
nand U35829 (N_35829,N_25239,N_28778);
xor U35830 (N_35830,N_27123,N_26890);
or U35831 (N_35831,N_29084,N_23579);
and U35832 (N_35832,N_23552,N_28721);
xor U35833 (N_35833,N_20538,N_24944);
nand U35834 (N_35834,N_25072,N_21221);
and U35835 (N_35835,N_20860,N_24999);
nor U35836 (N_35836,N_26564,N_26313);
or U35837 (N_35837,N_26746,N_26872);
and U35838 (N_35838,N_27210,N_21565);
nor U35839 (N_35839,N_20044,N_24432);
nand U35840 (N_35840,N_23100,N_27067);
nand U35841 (N_35841,N_24448,N_23711);
nand U35842 (N_35842,N_24136,N_27406);
and U35843 (N_35843,N_21494,N_26449);
or U35844 (N_35844,N_21798,N_24137);
nand U35845 (N_35845,N_29638,N_26904);
nor U35846 (N_35846,N_28634,N_23037);
nand U35847 (N_35847,N_24401,N_29607);
xor U35848 (N_35848,N_27213,N_25025);
or U35849 (N_35849,N_26560,N_28175);
nand U35850 (N_35850,N_29799,N_29599);
or U35851 (N_35851,N_28484,N_29402);
nor U35852 (N_35852,N_20164,N_25698);
nand U35853 (N_35853,N_23995,N_25034);
and U35854 (N_35854,N_25497,N_25194);
nand U35855 (N_35855,N_24950,N_26515);
and U35856 (N_35856,N_23034,N_23759);
or U35857 (N_35857,N_22132,N_29245);
and U35858 (N_35858,N_27579,N_26203);
and U35859 (N_35859,N_27825,N_29128);
or U35860 (N_35860,N_26607,N_28440);
or U35861 (N_35861,N_26793,N_23962);
nand U35862 (N_35862,N_29203,N_25337);
or U35863 (N_35863,N_28540,N_29380);
xor U35864 (N_35864,N_24584,N_21768);
or U35865 (N_35865,N_27637,N_26631);
nand U35866 (N_35866,N_29188,N_21379);
xor U35867 (N_35867,N_23600,N_28608);
nand U35868 (N_35868,N_21799,N_27581);
or U35869 (N_35869,N_28147,N_27661);
and U35870 (N_35870,N_21529,N_26566);
nor U35871 (N_35871,N_21962,N_24757);
and U35872 (N_35872,N_29942,N_23326);
nor U35873 (N_35873,N_29250,N_22758);
or U35874 (N_35874,N_27396,N_25079);
nand U35875 (N_35875,N_28237,N_20031);
or U35876 (N_35876,N_23918,N_20281);
nand U35877 (N_35877,N_26337,N_20314);
xor U35878 (N_35878,N_29650,N_23773);
nor U35879 (N_35879,N_20907,N_22907);
nor U35880 (N_35880,N_28718,N_25090);
or U35881 (N_35881,N_22518,N_26752);
or U35882 (N_35882,N_29381,N_29466);
or U35883 (N_35883,N_23034,N_23742);
nor U35884 (N_35884,N_29182,N_26010);
or U35885 (N_35885,N_25261,N_28261);
nand U35886 (N_35886,N_23050,N_24093);
or U35887 (N_35887,N_21134,N_23129);
nand U35888 (N_35888,N_29310,N_25388);
and U35889 (N_35889,N_20201,N_23448);
nand U35890 (N_35890,N_21817,N_28698);
nor U35891 (N_35891,N_29523,N_26325);
nor U35892 (N_35892,N_21251,N_20453);
or U35893 (N_35893,N_29550,N_23119);
nand U35894 (N_35894,N_29861,N_25279);
or U35895 (N_35895,N_26878,N_24176);
or U35896 (N_35896,N_25419,N_27547);
nand U35897 (N_35897,N_20669,N_20704);
nor U35898 (N_35898,N_25224,N_23794);
and U35899 (N_35899,N_25396,N_21359);
nand U35900 (N_35900,N_25797,N_20042);
nand U35901 (N_35901,N_29111,N_28250);
nor U35902 (N_35902,N_28742,N_24312);
nand U35903 (N_35903,N_29764,N_27873);
and U35904 (N_35904,N_24725,N_29797);
nand U35905 (N_35905,N_24382,N_22805);
nor U35906 (N_35906,N_21630,N_22611);
nand U35907 (N_35907,N_22923,N_22286);
xor U35908 (N_35908,N_23390,N_28544);
or U35909 (N_35909,N_21574,N_29818);
or U35910 (N_35910,N_22039,N_28868);
nand U35911 (N_35911,N_28366,N_22288);
nor U35912 (N_35912,N_28356,N_24102);
and U35913 (N_35913,N_28057,N_22560);
nand U35914 (N_35914,N_25345,N_26729);
nor U35915 (N_35915,N_25788,N_21903);
and U35916 (N_35916,N_21883,N_26614);
nand U35917 (N_35917,N_20166,N_29041);
or U35918 (N_35918,N_27493,N_24609);
nor U35919 (N_35919,N_29768,N_20573);
and U35920 (N_35920,N_20031,N_20673);
nor U35921 (N_35921,N_20707,N_22506);
and U35922 (N_35922,N_28265,N_20829);
and U35923 (N_35923,N_23719,N_29399);
nor U35924 (N_35924,N_25496,N_23111);
nand U35925 (N_35925,N_24960,N_29794);
nor U35926 (N_35926,N_29714,N_20797);
nand U35927 (N_35927,N_22584,N_28957);
nor U35928 (N_35928,N_27834,N_29204);
xor U35929 (N_35929,N_28179,N_23449);
nor U35930 (N_35930,N_20191,N_22970);
nand U35931 (N_35931,N_22538,N_24229);
nand U35932 (N_35932,N_24534,N_28461);
nand U35933 (N_35933,N_29293,N_29822);
or U35934 (N_35934,N_20998,N_21202);
nand U35935 (N_35935,N_27675,N_25070);
nand U35936 (N_35936,N_20787,N_23305);
nand U35937 (N_35937,N_23476,N_20594);
nor U35938 (N_35938,N_24121,N_28780);
xnor U35939 (N_35939,N_27785,N_28239);
nor U35940 (N_35940,N_28406,N_24079);
xor U35941 (N_35941,N_20804,N_21256);
nor U35942 (N_35942,N_29832,N_21295);
nor U35943 (N_35943,N_26244,N_26868);
or U35944 (N_35944,N_28975,N_23485);
and U35945 (N_35945,N_21511,N_20021);
nand U35946 (N_35946,N_28550,N_21967);
and U35947 (N_35947,N_27518,N_22823);
nor U35948 (N_35948,N_22138,N_25020);
nor U35949 (N_35949,N_29076,N_22147);
or U35950 (N_35950,N_20921,N_20113);
nor U35951 (N_35951,N_21837,N_29621);
or U35952 (N_35952,N_27739,N_26704);
nand U35953 (N_35953,N_26379,N_25157);
nor U35954 (N_35954,N_29713,N_23913);
nand U35955 (N_35955,N_27560,N_25388);
and U35956 (N_35956,N_22439,N_25947);
and U35957 (N_35957,N_20464,N_24905);
and U35958 (N_35958,N_26833,N_20258);
nor U35959 (N_35959,N_22386,N_20060);
and U35960 (N_35960,N_23927,N_20199);
nand U35961 (N_35961,N_20831,N_21619);
xnor U35962 (N_35962,N_25522,N_22511);
nor U35963 (N_35963,N_28459,N_28254);
nand U35964 (N_35964,N_28427,N_21070);
nor U35965 (N_35965,N_23034,N_24673);
or U35966 (N_35966,N_22794,N_27620);
and U35967 (N_35967,N_22695,N_21342);
and U35968 (N_35968,N_28382,N_21537);
nand U35969 (N_35969,N_27090,N_28048);
or U35970 (N_35970,N_25335,N_23523);
nand U35971 (N_35971,N_29894,N_22679);
and U35972 (N_35972,N_29042,N_23545);
and U35973 (N_35973,N_20062,N_27025);
nand U35974 (N_35974,N_28981,N_21292);
nand U35975 (N_35975,N_28959,N_28018);
or U35976 (N_35976,N_26164,N_29480);
nand U35977 (N_35977,N_24318,N_27658);
nand U35978 (N_35978,N_24118,N_29479);
or U35979 (N_35979,N_25352,N_25773);
or U35980 (N_35980,N_29326,N_25469);
nor U35981 (N_35981,N_24466,N_20805);
nor U35982 (N_35982,N_24398,N_28161);
nand U35983 (N_35983,N_20437,N_23359);
nand U35984 (N_35984,N_26899,N_23064);
nor U35985 (N_35985,N_25661,N_23226);
or U35986 (N_35986,N_20940,N_26044);
or U35987 (N_35987,N_22208,N_25097);
nor U35988 (N_35988,N_20031,N_28901);
or U35989 (N_35989,N_28751,N_21033);
xnor U35990 (N_35990,N_20038,N_21183);
nand U35991 (N_35991,N_23211,N_24821);
and U35992 (N_35992,N_25535,N_20103);
or U35993 (N_35993,N_21189,N_26611);
nor U35994 (N_35994,N_28674,N_24280);
nand U35995 (N_35995,N_26486,N_23157);
or U35996 (N_35996,N_27540,N_24369);
or U35997 (N_35997,N_23368,N_20910);
nand U35998 (N_35998,N_29321,N_23797);
nand U35999 (N_35999,N_29090,N_29119);
nand U36000 (N_36000,N_21777,N_25727);
nor U36001 (N_36001,N_24122,N_20009);
nand U36002 (N_36002,N_26330,N_20845);
or U36003 (N_36003,N_20861,N_20764);
nor U36004 (N_36004,N_24335,N_28740);
and U36005 (N_36005,N_23076,N_23724);
nand U36006 (N_36006,N_23139,N_22774);
nor U36007 (N_36007,N_26409,N_26495);
xor U36008 (N_36008,N_20525,N_26144);
xnor U36009 (N_36009,N_24831,N_25299);
and U36010 (N_36010,N_20927,N_23509);
and U36011 (N_36011,N_27820,N_24509);
nor U36012 (N_36012,N_22956,N_20818);
nand U36013 (N_36013,N_26580,N_27796);
nor U36014 (N_36014,N_29784,N_24262);
xnor U36015 (N_36015,N_20101,N_25157);
xnor U36016 (N_36016,N_28247,N_27812);
nor U36017 (N_36017,N_20347,N_23085);
or U36018 (N_36018,N_20876,N_27086);
and U36019 (N_36019,N_20919,N_27978);
nor U36020 (N_36020,N_25427,N_27680);
or U36021 (N_36021,N_25649,N_27036);
nor U36022 (N_36022,N_28713,N_28254);
nor U36023 (N_36023,N_22485,N_29273);
and U36024 (N_36024,N_29981,N_25179);
and U36025 (N_36025,N_22492,N_28501);
nand U36026 (N_36026,N_29554,N_29888);
nand U36027 (N_36027,N_21669,N_28382);
nor U36028 (N_36028,N_21458,N_23766);
or U36029 (N_36029,N_21527,N_20974);
nor U36030 (N_36030,N_28565,N_20721);
and U36031 (N_36031,N_23338,N_20358);
and U36032 (N_36032,N_29876,N_28487);
and U36033 (N_36033,N_26866,N_24235);
nor U36034 (N_36034,N_24630,N_21868);
or U36035 (N_36035,N_28224,N_27914);
and U36036 (N_36036,N_24129,N_23527);
and U36037 (N_36037,N_28309,N_28159);
or U36038 (N_36038,N_25222,N_27402);
nand U36039 (N_36039,N_26835,N_27260);
xor U36040 (N_36040,N_26289,N_27952);
and U36041 (N_36041,N_24100,N_26132);
and U36042 (N_36042,N_21295,N_25260);
nand U36043 (N_36043,N_24644,N_29752);
nand U36044 (N_36044,N_22142,N_26650);
or U36045 (N_36045,N_25416,N_22374);
nand U36046 (N_36046,N_22430,N_28284);
nor U36047 (N_36047,N_28592,N_27443);
or U36048 (N_36048,N_25786,N_23312);
nor U36049 (N_36049,N_21860,N_26994);
and U36050 (N_36050,N_28026,N_23345);
and U36051 (N_36051,N_28785,N_29035);
and U36052 (N_36052,N_21965,N_21913);
nor U36053 (N_36053,N_24448,N_22953);
or U36054 (N_36054,N_22070,N_23632);
nand U36055 (N_36055,N_21861,N_23724);
xor U36056 (N_36056,N_24796,N_27617);
nor U36057 (N_36057,N_20157,N_23606);
nor U36058 (N_36058,N_25479,N_25416);
nor U36059 (N_36059,N_24040,N_26387);
or U36060 (N_36060,N_28754,N_25128);
nand U36061 (N_36061,N_27586,N_23060);
nand U36062 (N_36062,N_25238,N_24530);
or U36063 (N_36063,N_25660,N_29580);
and U36064 (N_36064,N_25076,N_29138);
nand U36065 (N_36065,N_21497,N_25118);
nor U36066 (N_36066,N_25282,N_25813);
and U36067 (N_36067,N_21882,N_23812);
nor U36068 (N_36068,N_20732,N_29286);
nand U36069 (N_36069,N_20057,N_28308);
and U36070 (N_36070,N_20944,N_23028);
nand U36071 (N_36071,N_24547,N_20146);
and U36072 (N_36072,N_22484,N_25812);
or U36073 (N_36073,N_23487,N_21381);
and U36074 (N_36074,N_29709,N_29462);
nor U36075 (N_36075,N_22696,N_26421);
or U36076 (N_36076,N_21724,N_24434);
nor U36077 (N_36077,N_20352,N_27752);
nand U36078 (N_36078,N_28399,N_23764);
or U36079 (N_36079,N_28879,N_21549);
nand U36080 (N_36080,N_24894,N_23085);
and U36081 (N_36081,N_20341,N_27069);
nor U36082 (N_36082,N_22336,N_23583);
and U36083 (N_36083,N_23830,N_22418);
nand U36084 (N_36084,N_25041,N_29051);
nor U36085 (N_36085,N_23561,N_20826);
and U36086 (N_36086,N_28729,N_25382);
and U36087 (N_36087,N_29690,N_20273);
or U36088 (N_36088,N_26078,N_22802);
nor U36089 (N_36089,N_29641,N_26632);
nand U36090 (N_36090,N_21161,N_20645);
or U36091 (N_36091,N_25338,N_22714);
and U36092 (N_36092,N_29636,N_20819);
nor U36093 (N_36093,N_24968,N_27174);
nor U36094 (N_36094,N_26532,N_23912);
nor U36095 (N_36095,N_28624,N_29035);
or U36096 (N_36096,N_27963,N_28620);
nor U36097 (N_36097,N_22780,N_26028);
or U36098 (N_36098,N_23365,N_24272);
or U36099 (N_36099,N_20249,N_26566);
or U36100 (N_36100,N_25810,N_23364);
nand U36101 (N_36101,N_29289,N_20408);
nand U36102 (N_36102,N_27496,N_20447);
or U36103 (N_36103,N_22957,N_24548);
or U36104 (N_36104,N_25048,N_28702);
or U36105 (N_36105,N_25502,N_25285);
xnor U36106 (N_36106,N_23144,N_25791);
and U36107 (N_36107,N_25947,N_25731);
nand U36108 (N_36108,N_29181,N_26022);
or U36109 (N_36109,N_25208,N_27240);
nor U36110 (N_36110,N_29175,N_22438);
or U36111 (N_36111,N_24667,N_29639);
xor U36112 (N_36112,N_20101,N_26588);
and U36113 (N_36113,N_21024,N_24416);
nor U36114 (N_36114,N_28733,N_27965);
xnor U36115 (N_36115,N_28464,N_27490);
nand U36116 (N_36116,N_21262,N_22548);
nor U36117 (N_36117,N_23990,N_27605);
or U36118 (N_36118,N_27373,N_20741);
nand U36119 (N_36119,N_24849,N_23285);
xnor U36120 (N_36120,N_25999,N_26221);
nor U36121 (N_36121,N_26237,N_21448);
nor U36122 (N_36122,N_25659,N_25966);
nor U36123 (N_36123,N_21130,N_23324);
and U36124 (N_36124,N_20117,N_22252);
and U36125 (N_36125,N_22117,N_29436);
and U36126 (N_36126,N_27691,N_20161);
or U36127 (N_36127,N_24814,N_21972);
nor U36128 (N_36128,N_29230,N_21079);
and U36129 (N_36129,N_28813,N_24118);
and U36130 (N_36130,N_26892,N_29049);
nor U36131 (N_36131,N_20430,N_22161);
nor U36132 (N_36132,N_22744,N_28024);
or U36133 (N_36133,N_20188,N_29660);
nand U36134 (N_36134,N_24816,N_29068);
nor U36135 (N_36135,N_28741,N_22831);
xnor U36136 (N_36136,N_22929,N_28053);
nor U36137 (N_36137,N_27433,N_20852);
nand U36138 (N_36138,N_26687,N_22678);
nor U36139 (N_36139,N_22166,N_29395);
nor U36140 (N_36140,N_25624,N_27165);
nand U36141 (N_36141,N_25118,N_20399);
nor U36142 (N_36142,N_29933,N_20000);
xor U36143 (N_36143,N_24600,N_27905);
nand U36144 (N_36144,N_20774,N_20732);
xnor U36145 (N_36145,N_28248,N_24054);
xor U36146 (N_36146,N_26511,N_20692);
or U36147 (N_36147,N_25368,N_22567);
nand U36148 (N_36148,N_27776,N_24092);
nor U36149 (N_36149,N_20110,N_28550);
and U36150 (N_36150,N_28729,N_22113);
or U36151 (N_36151,N_26813,N_21729);
xor U36152 (N_36152,N_25675,N_24078);
nand U36153 (N_36153,N_22163,N_20318);
xor U36154 (N_36154,N_25653,N_26878);
nand U36155 (N_36155,N_24724,N_29007);
or U36156 (N_36156,N_21522,N_22156);
nor U36157 (N_36157,N_25594,N_27931);
xor U36158 (N_36158,N_28174,N_22820);
nor U36159 (N_36159,N_22914,N_28412);
xor U36160 (N_36160,N_20027,N_24313);
or U36161 (N_36161,N_25908,N_22509);
and U36162 (N_36162,N_24426,N_21498);
nor U36163 (N_36163,N_22125,N_20205);
nor U36164 (N_36164,N_25915,N_29712);
or U36165 (N_36165,N_22001,N_23589);
nand U36166 (N_36166,N_21562,N_20948);
or U36167 (N_36167,N_26090,N_20321);
or U36168 (N_36168,N_21612,N_21003);
nand U36169 (N_36169,N_22276,N_29904);
or U36170 (N_36170,N_25507,N_23872);
nand U36171 (N_36171,N_29060,N_26529);
nand U36172 (N_36172,N_24540,N_21926);
and U36173 (N_36173,N_24045,N_21378);
or U36174 (N_36174,N_21067,N_28344);
nand U36175 (N_36175,N_23515,N_26422);
nand U36176 (N_36176,N_25885,N_27312);
and U36177 (N_36177,N_29467,N_28007);
and U36178 (N_36178,N_20356,N_26655);
nand U36179 (N_36179,N_26707,N_25526);
or U36180 (N_36180,N_27227,N_25490);
or U36181 (N_36181,N_22438,N_22762);
nor U36182 (N_36182,N_28586,N_25998);
nor U36183 (N_36183,N_21150,N_28679);
or U36184 (N_36184,N_25877,N_27170);
or U36185 (N_36185,N_21279,N_28669);
nor U36186 (N_36186,N_23474,N_23697);
xor U36187 (N_36187,N_29608,N_28472);
nand U36188 (N_36188,N_28153,N_23439);
nand U36189 (N_36189,N_21780,N_26069);
nor U36190 (N_36190,N_28186,N_29777);
nand U36191 (N_36191,N_27775,N_23297);
nor U36192 (N_36192,N_28224,N_21227);
or U36193 (N_36193,N_20164,N_26974);
nor U36194 (N_36194,N_20461,N_28872);
nor U36195 (N_36195,N_24336,N_26577);
and U36196 (N_36196,N_27830,N_20251);
or U36197 (N_36197,N_29646,N_26110);
nor U36198 (N_36198,N_20315,N_21482);
and U36199 (N_36199,N_25269,N_25672);
and U36200 (N_36200,N_28432,N_24536);
and U36201 (N_36201,N_29108,N_27743);
nand U36202 (N_36202,N_25883,N_21196);
nor U36203 (N_36203,N_26674,N_25701);
and U36204 (N_36204,N_26388,N_20631);
and U36205 (N_36205,N_27219,N_23743);
xor U36206 (N_36206,N_24840,N_26596);
xnor U36207 (N_36207,N_26444,N_28967);
or U36208 (N_36208,N_25090,N_22270);
or U36209 (N_36209,N_23227,N_23306);
and U36210 (N_36210,N_26074,N_28834);
or U36211 (N_36211,N_22922,N_29228);
nand U36212 (N_36212,N_28510,N_28727);
or U36213 (N_36213,N_26349,N_29146);
nand U36214 (N_36214,N_21819,N_28787);
or U36215 (N_36215,N_26519,N_27170);
nand U36216 (N_36216,N_21779,N_20927);
or U36217 (N_36217,N_23835,N_29380);
nor U36218 (N_36218,N_27187,N_29804);
nor U36219 (N_36219,N_27436,N_25092);
nand U36220 (N_36220,N_28390,N_25921);
and U36221 (N_36221,N_21572,N_26786);
and U36222 (N_36222,N_28601,N_21971);
nand U36223 (N_36223,N_22881,N_29060);
xor U36224 (N_36224,N_28189,N_22747);
nand U36225 (N_36225,N_23316,N_27123);
nand U36226 (N_36226,N_26741,N_20831);
nor U36227 (N_36227,N_21749,N_21340);
and U36228 (N_36228,N_22996,N_22894);
nor U36229 (N_36229,N_25511,N_26658);
and U36230 (N_36230,N_20727,N_26965);
and U36231 (N_36231,N_25582,N_23678);
or U36232 (N_36232,N_24467,N_27152);
xor U36233 (N_36233,N_27717,N_28529);
and U36234 (N_36234,N_20736,N_25754);
or U36235 (N_36235,N_26359,N_26802);
nand U36236 (N_36236,N_20715,N_28290);
and U36237 (N_36237,N_20854,N_24237);
nor U36238 (N_36238,N_25420,N_22103);
or U36239 (N_36239,N_22048,N_24309);
xor U36240 (N_36240,N_28265,N_27675);
and U36241 (N_36241,N_20577,N_25988);
nand U36242 (N_36242,N_27685,N_22901);
nand U36243 (N_36243,N_27283,N_27694);
or U36244 (N_36244,N_25398,N_27809);
and U36245 (N_36245,N_28154,N_27656);
xnor U36246 (N_36246,N_21685,N_27261);
and U36247 (N_36247,N_21901,N_28899);
xor U36248 (N_36248,N_26744,N_27742);
xor U36249 (N_36249,N_23748,N_20576);
and U36250 (N_36250,N_21535,N_25906);
and U36251 (N_36251,N_27749,N_29311);
and U36252 (N_36252,N_21360,N_28338);
nand U36253 (N_36253,N_29378,N_25096);
nor U36254 (N_36254,N_26966,N_20678);
and U36255 (N_36255,N_27213,N_24420);
or U36256 (N_36256,N_27431,N_27122);
nor U36257 (N_36257,N_27350,N_26345);
and U36258 (N_36258,N_29817,N_25122);
or U36259 (N_36259,N_29329,N_25109);
xnor U36260 (N_36260,N_25184,N_28543);
nand U36261 (N_36261,N_23744,N_20943);
nand U36262 (N_36262,N_29378,N_29334);
and U36263 (N_36263,N_24290,N_29650);
or U36264 (N_36264,N_22220,N_26594);
nand U36265 (N_36265,N_26917,N_27581);
nand U36266 (N_36266,N_26881,N_23213);
and U36267 (N_36267,N_26923,N_27131);
and U36268 (N_36268,N_24864,N_29916);
nand U36269 (N_36269,N_22607,N_22160);
nor U36270 (N_36270,N_24443,N_21569);
and U36271 (N_36271,N_28716,N_29697);
nand U36272 (N_36272,N_24998,N_25603);
nor U36273 (N_36273,N_26335,N_26676);
or U36274 (N_36274,N_26842,N_20520);
or U36275 (N_36275,N_22172,N_23309);
nor U36276 (N_36276,N_21257,N_21194);
xor U36277 (N_36277,N_24181,N_24315);
nand U36278 (N_36278,N_22527,N_25629);
nand U36279 (N_36279,N_27047,N_20276);
nor U36280 (N_36280,N_22524,N_28296);
xnor U36281 (N_36281,N_21810,N_26700);
nand U36282 (N_36282,N_21333,N_27008);
and U36283 (N_36283,N_21816,N_23202);
nor U36284 (N_36284,N_29334,N_20533);
or U36285 (N_36285,N_22207,N_21605);
nand U36286 (N_36286,N_29384,N_22288);
and U36287 (N_36287,N_20309,N_20851);
or U36288 (N_36288,N_29935,N_20830);
xor U36289 (N_36289,N_20202,N_24918);
or U36290 (N_36290,N_21990,N_28142);
nor U36291 (N_36291,N_23665,N_25791);
xnor U36292 (N_36292,N_21783,N_24443);
nand U36293 (N_36293,N_26910,N_21130);
nand U36294 (N_36294,N_26721,N_28542);
or U36295 (N_36295,N_25658,N_29164);
or U36296 (N_36296,N_25923,N_20439);
nand U36297 (N_36297,N_25418,N_29530);
nand U36298 (N_36298,N_23865,N_23416);
nor U36299 (N_36299,N_20441,N_26901);
xnor U36300 (N_36300,N_27845,N_21731);
and U36301 (N_36301,N_24797,N_23472);
xor U36302 (N_36302,N_28300,N_21998);
or U36303 (N_36303,N_22983,N_22698);
nand U36304 (N_36304,N_29235,N_23327);
and U36305 (N_36305,N_22654,N_29654);
or U36306 (N_36306,N_24213,N_27027);
nand U36307 (N_36307,N_24619,N_23753);
or U36308 (N_36308,N_21298,N_25692);
nand U36309 (N_36309,N_29293,N_21385);
or U36310 (N_36310,N_24612,N_23455);
and U36311 (N_36311,N_27040,N_23731);
nand U36312 (N_36312,N_20715,N_28532);
or U36313 (N_36313,N_23285,N_29654);
nor U36314 (N_36314,N_24674,N_23569);
or U36315 (N_36315,N_23309,N_26077);
nand U36316 (N_36316,N_27729,N_25191);
xnor U36317 (N_36317,N_20500,N_25835);
and U36318 (N_36318,N_27430,N_29211);
and U36319 (N_36319,N_29142,N_22708);
nand U36320 (N_36320,N_25818,N_20044);
or U36321 (N_36321,N_25547,N_24424);
or U36322 (N_36322,N_22292,N_25279);
nand U36323 (N_36323,N_24040,N_21587);
and U36324 (N_36324,N_25539,N_21392);
nand U36325 (N_36325,N_25433,N_25217);
xnor U36326 (N_36326,N_29314,N_22889);
nor U36327 (N_36327,N_23623,N_27908);
or U36328 (N_36328,N_25642,N_27873);
nor U36329 (N_36329,N_24124,N_26710);
nor U36330 (N_36330,N_29484,N_29807);
nand U36331 (N_36331,N_26708,N_26652);
nand U36332 (N_36332,N_24935,N_24447);
nor U36333 (N_36333,N_28049,N_23567);
and U36334 (N_36334,N_21139,N_20847);
or U36335 (N_36335,N_20958,N_21128);
and U36336 (N_36336,N_21046,N_21141);
nor U36337 (N_36337,N_29953,N_27700);
and U36338 (N_36338,N_23848,N_28803);
and U36339 (N_36339,N_28677,N_24215);
or U36340 (N_36340,N_20991,N_29173);
nand U36341 (N_36341,N_20105,N_29965);
nand U36342 (N_36342,N_22726,N_27484);
nand U36343 (N_36343,N_25650,N_27002);
or U36344 (N_36344,N_22084,N_20608);
and U36345 (N_36345,N_21732,N_23549);
nand U36346 (N_36346,N_22299,N_23215);
or U36347 (N_36347,N_28084,N_21775);
nand U36348 (N_36348,N_29987,N_23451);
or U36349 (N_36349,N_21877,N_24860);
or U36350 (N_36350,N_21294,N_29347);
and U36351 (N_36351,N_24307,N_27032);
xor U36352 (N_36352,N_28925,N_26868);
nor U36353 (N_36353,N_26858,N_26428);
nor U36354 (N_36354,N_24028,N_24086);
or U36355 (N_36355,N_23340,N_24096);
nor U36356 (N_36356,N_22440,N_24449);
and U36357 (N_36357,N_27944,N_24980);
nand U36358 (N_36358,N_24033,N_22047);
nand U36359 (N_36359,N_29815,N_20744);
xnor U36360 (N_36360,N_21661,N_29922);
or U36361 (N_36361,N_21824,N_22373);
xnor U36362 (N_36362,N_24582,N_29185);
xnor U36363 (N_36363,N_20909,N_27551);
or U36364 (N_36364,N_21838,N_27594);
and U36365 (N_36365,N_27273,N_23238);
nand U36366 (N_36366,N_29893,N_26844);
nor U36367 (N_36367,N_25765,N_29363);
or U36368 (N_36368,N_28650,N_24510);
or U36369 (N_36369,N_29455,N_29203);
or U36370 (N_36370,N_28692,N_22294);
nand U36371 (N_36371,N_24866,N_20930);
or U36372 (N_36372,N_29143,N_20074);
or U36373 (N_36373,N_24005,N_22331);
nor U36374 (N_36374,N_29210,N_28389);
nor U36375 (N_36375,N_22284,N_26168);
or U36376 (N_36376,N_22807,N_27655);
and U36377 (N_36377,N_24099,N_28131);
or U36378 (N_36378,N_27485,N_24044);
or U36379 (N_36379,N_28770,N_26998);
or U36380 (N_36380,N_26816,N_20405);
nand U36381 (N_36381,N_24310,N_21716);
and U36382 (N_36382,N_27957,N_22669);
and U36383 (N_36383,N_24605,N_29851);
or U36384 (N_36384,N_28392,N_23047);
nand U36385 (N_36385,N_24218,N_29016);
nand U36386 (N_36386,N_25868,N_26662);
nor U36387 (N_36387,N_22056,N_20439);
nor U36388 (N_36388,N_25910,N_21376);
or U36389 (N_36389,N_26808,N_26041);
nor U36390 (N_36390,N_20213,N_24487);
nand U36391 (N_36391,N_21555,N_22037);
nor U36392 (N_36392,N_22470,N_22368);
or U36393 (N_36393,N_26799,N_28148);
and U36394 (N_36394,N_20419,N_26593);
nand U36395 (N_36395,N_23738,N_28719);
nand U36396 (N_36396,N_20592,N_27171);
and U36397 (N_36397,N_24819,N_28237);
nand U36398 (N_36398,N_21011,N_25138);
nand U36399 (N_36399,N_25590,N_28678);
or U36400 (N_36400,N_24499,N_24985);
xnor U36401 (N_36401,N_21804,N_20108);
or U36402 (N_36402,N_27988,N_27890);
nor U36403 (N_36403,N_28667,N_26737);
and U36404 (N_36404,N_21970,N_23642);
nor U36405 (N_36405,N_27271,N_25025);
nor U36406 (N_36406,N_28002,N_21403);
nand U36407 (N_36407,N_25942,N_29316);
nor U36408 (N_36408,N_27166,N_20400);
or U36409 (N_36409,N_23651,N_24497);
and U36410 (N_36410,N_28220,N_24009);
xnor U36411 (N_36411,N_25236,N_24069);
or U36412 (N_36412,N_21301,N_21780);
nand U36413 (N_36413,N_21289,N_27359);
nor U36414 (N_36414,N_20703,N_25494);
xor U36415 (N_36415,N_21451,N_24371);
or U36416 (N_36416,N_29309,N_23540);
or U36417 (N_36417,N_20066,N_29815);
nor U36418 (N_36418,N_25736,N_27896);
and U36419 (N_36419,N_29701,N_23982);
and U36420 (N_36420,N_28884,N_21180);
or U36421 (N_36421,N_29847,N_23635);
and U36422 (N_36422,N_27026,N_26668);
and U36423 (N_36423,N_22351,N_21381);
nor U36424 (N_36424,N_29431,N_21493);
and U36425 (N_36425,N_25899,N_24501);
nor U36426 (N_36426,N_25958,N_27087);
nand U36427 (N_36427,N_24623,N_29228);
and U36428 (N_36428,N_26512,N_24591);
or U36429 (N_36429,N_24353,N_29608);
nor U36430 (N_36430,N_20458,N_26756);
and U36431 (N_36431,N_25522,N_29930);
nand U36432 (N_36432,N_23075,N_25842);
and U36433 (N_36433,N_22264,N_26182);
nand U36434 (N_36434,N_20594,N_24165);
or U36435 (N_36435,N_24119,N_27177);
and U36436 (N_36436,N_26315,N_25539);
or U36437 (N_36437,N_28607,N_22855);
nand U36438 (N_36438,N_24497,N_22275);
and U36439 (N_36439,N_21025,N_25095);
nand U36440 (N_36440,N_25825,N_28414);
or U36441 (N_36441,N_23521,N_25688);
or U36442 (N_36442,N_28845,N_26901);
nor U36443 (N_36443,N_21904,N_28818);
xor U36444 (N_36444,N_28169,N_21260);
nor U36445 (N_36445,N_26933,N_28598);
or U36446 (N_36446,N_25961,N_20614);
and U36447 (N_36447,N_23069,N_26488);
and U36448 (N_36448,N_24131,N_20810);
and U36449 (N_36449,N_20490,N_28700);
and U36450 (N_36450,N_22255,N_27535);
and U36451 (N_36451,N_29213,N_28223);
nor U36452 (N_36452,N_28882,N_26065);
xnor U36453 (N_36453,N_21507,N_27163);
or U36454 (N_36454,N_29114,N_29129);
or U36455 (N_36455,N_24973,N_20849);
or U36456 (N_36456,N_24640,N_23272);
nand U36457 (N_36457,N_25952,N_28989);
xnor U36458 (N_36458,N_29653,N_27205);
or U36459 (N_36459,N_25118,N_28016);
xor U36460 (N_36460,N_22022,N_27392);
and U36461 (N_36461,N_27923,N_26592);
or U36462 (N_36462,N_27877,N_27317);
or U36463 (N_36463,N_26796,N_21125);
or U36464 (N_36464,N_29803,N_20753);
or U36465 (N_36465,N_25202,N_26888);
nand U36466 (N_36466,N_26987,N_26774);
or U36467 (N_36467,N_23066,N_26541);
xnor U36468 (N_36468,N_27068,N_21310);
nand U36469 (N_36469,N_26844,N_26945);
and U36470 (N_36470,N_27148,N_24640);
nor U36471 (N_36471,N_29681,N_26755);
and U36472 (N_36472,N_21365,N_27605);
and U36473 (N_36473,N_28068,N_22392);
or U36474 (N_36474,N_24395,N_23874);
nor U36475 (N_36475,N_28521,N_20337);
and U36476 (N_36476,N_22904,N_26847);
or U36477 (N_36477,N_23925,N_20759);
nand U36478 (N_36478,N_25635,N_22498);
nand U36479 (N_36479,N_24640,N_27825);
xor U36480 (N_36480,N_22195,N_28293);
and U36481 (N_36481,N_29958,N_26843);
nor U36482 (N_36482,N_22033,N_23201);
nor U36483 (N_36483,N_20813,N_29247);
and U36484 (N_36484,N_24986,N_25966);
nor U36485 (N_36485,N_25928,N_20561);
nor U36486 (N_36486,N_24212,N_21959);
nand U36487 (N_36487,N_25444,N_24145);
or U36488 (N_36488,N_23372,N_29583);
and U36489 (N_36489,N_23772,N_29652);
and U36490 (N_36490,N_20699,N_29991);
and U36491 (N_36491,N_29804,N_28010);
nor U36492 (N_36492,N_20369,N_22712);
nand U36493 (N_36493,N_28839,N_22777);
nor U36494 (N_36494,N_24490,N_26623);
nand U36495 (N_36495,N_21212,N_26248);
or U36496 (N_36496,N_25510,N_26056);
nand U36497 (N_36497,N_22879,N_21168);
or U36498 (N_36498,N_29412,N_23008);
nand U36499 (N_36499,N_24932,N_26593);
and U36500 (N_36500,N_23898,N_27572);
nand U36501 (N_36501,N_29655,N_28547);
or U36502 (N_36502,N_25404,N_27542);
nor U36503 (N_36503,N_28134,N_22762);
nand U36504 (N_36504,N_20763,N_21080);
nand U36505 (N_36505,N_26704,N_24829);
nand U36506 (N_36506,N_26394,N_27786);
or U36507 (N_36507,N_29034,N_24749);
nor U36508 (N_36508,N_22713,N_21346);
nor U36509 (N_36509,N_24076,N_29229);
or U36510 (N_36510,N_27755,N_20218);
or U36511 (N_36511,N_23810,N_26792);
and U36512 (N_36512,N_25586,N_22607);
or U36513 (N_36513,N_24262,N_27912);
and U36514 (N_36514,N_25620,N_23228);
and U36515 (N_36515,N_20006,N_25567);
or U36516 (N_36516,N_27746,N_22474);
nand U36517 (N_36517,N_20560,N_21023);
nand U36518 (N_36518,N_25249,N_21921);
nor U36519 (N_36519,N_26089,N_25634);
or U36520 (N_36520,N_29932,N_22290);
and U36521 (N_36521,N_20227,N_29594);
and U36522 (N_36522,N_26271,N_25289);
nand U36523 (N_36523,N_26745,N_22906);
or U36524 (N_36524,N_23680,N_22866);
and U36525 (N_36525,N_25880,N_25505);
xor U36526 (N_36526,N_22978,N_27590);
and U36527 (N_36527,N_20806,N_29995);
nor U36528 (N_36528,N_28594,N_24442);
xnor U36529 (N_36529,N_23263,N_29283);
nand U36530 (N_36530,N_29590,N_22809);
nor U36531 (N_36531,N_26626,N_24195);
or U36532 (N_36532,N_25178,N_27286);
nor U36533 (N_36533,N_24768,N_26383);
nor U36534 (N_36534,N_24618,N_26896);
nor U36535 (N_36535,N_21089,N_25236);
nand U36536 (N_36536,N_20191,N_23640);
and U36537 (N_36537,N_24125,N_23947);
and U36538 (N_36538,N_25494,N_21464);
xnor U36539 (N_36539,N_27275,N_28973);
nand U36540 (N_36540,N_25790,N_26380);
and U36541 (N_36541,N_24531,N_26671);
or U36542 (N_36542,N_26726,N_23612);
nor U36543 (N_36543,N_26847,N_21912);
and U36544 (N_36544,N_22548,N_21020);
or U36545 (N_36545,N_26874,N_20050);
nand U36546 (N_36546,N_22072,N_25677);
nor U36547 (N_36547,N_27086,N_25559);
nor U36548 (N_36548,N_25302,N_28913);
or U36549 (N_36549,N_20525,N_29987);
and U36550 (N_36550,N_23827,N_28904);
nand U36551 (N_36551,N_25770,N_29561);
nand U36552 (N_36552,N_21882,N_21023);
nor U36553 (N_36553,N_27471,N_29464);
nand U36554 (N_36554,N_21529,N_28708);
nand U36555 (N_36555,N_26844,N_29471);
nand U36556 (N_36556,N_23405,N_24129);
nand U36557 (N_36557,N_21708,N_26763);
and U36558 (N_36558,N_25632,N_29687);
or U36559 (N_36559,N_27908,N_24079);
and U36560 (N_36560,N_20559,N_22677);
nand U36561 (N_36561,N_29299,N_20612);
nand U36562 (N_36562,N_21530,N_22349);
and U36563 (N_36563,N_26608,N_29829);
and U36564 (N_36564,N_20763,N_20407);
xor U36565 (N_36565,N_27779,N_26226);
xor U36566 (N_36566,N_27233,N_28843);
nand U36567 (N_36567,N_21174,N_25160);
nor U36568 (N_36568,N_25817,N_27233);
nand U36569 (N_36569,N_21153,N_22689);
nor U36570 (N_36570,N_23249,N_25989);
or U36571 (N_36571,N_23455,N_20990);
or U36572 (N_36572,N_24271,N_28530);
and U36573 (N_36573,N_23671,N_21700);
xor U36574 (N_36574,N_27016,N_25765);
nor U36575 (N_36575,N_28379,N_22037);
nand U36576 (N_36576,N_25532,N_22838);
xor U36577 (N_36577,N_23321,N_23087);
or U36578 (N_36578,N_25974,N_25363);
xnor U36579 (N_36579,N_23470,N_25786);
nor U36580 (N_36580,N_23689,N_29215);
nor U36581 (N_36581,N_27199,N_26801);
nor U36582 (N_36582,N_20212,N_24808);
or U36583 (N_36583,N_25426,N_29888);
nand U36584 (N_36584,N_26275,N_24886);
nand U36585 (N_36585,N_21183,N_20356);
and U36586 (N_36586,N_26135,N_24794);
or U36587 (N_36587,N_23316,N_29238);
or U36588 (N_36588,N_25337,N_22131);
or U36589 (N_36589,N_21958,N_21539);
nand U36590 (N_36590,N_21439,N_29719);
nand U36591 (N_36591,N_28943,N_24891);
nand U36592 (N_36592,N_21731,N_24018);
nand U36593 (N_36593,N_22896,N_22059);
xor U36594 (N_36594,N_23120,N_22647);
or U36595 (N_36595,N_28107,N_21996);
and U36596 (N_36596,N_23294,N_27013);
nand U36597 (N_36597,N_28358,N_21339);
nor U36598 (N_36598,N_21667,N_24782);
nand U36599 (N_36599,N_25359,N_27354);
nor U36600 (N_36600,N_20651,N_22627);
and U36601 (N_36601,N_22009,N_24551);
nor U36602 (N_36602,N_29423,N_29805);
and U36603 (N_36603,N_26704,N_20248);
or U36604 (N_36604,N_29280,N_25958);
nor U36605 (N_36605,N_25775,N_28792);
xnor U36606 (N_36606,N_23264,N_25161);
nor U36607 (N_36607,N_22584,N_24687);
xor U36608 (N_36608,N_29492,N_22353);
nor U36609 (N_36609,N_26414,N_27867);
xor U36610 (N_36610,N_28555,N_29382);
and U36611 (N_36611,N_28445,N_21528);
or U36612 (N_36612,N_25344,N_26746);
nand U36613 (N_36613,N_20686,N_22269);
nand U36614 (N_36614,N_20574,N_26023);
nand U36615 (N_36615,N_29506,N_22561);
nand U36616 (N_36616,N_22756,N_29307);
and U36617 (N_36617,N_24553,N_25373);
nand U36618 (N_36618,N_20874,N_22914);
nand U36619 (N_36619,N_22023,N_24678);
xnor U36620 (N_36620,N_23585,N_21085);
nand U36621 (N_36621,N_27403,N_26209);
nand U36622 (N_36622,N_27650,N_21522);
nand U36623 (N_36623,N_27567,N_24390);
or U36624 (N_36624,N_25406,N_22903);
or U36625 (N_36625,N_29910,N_27987);
nor U36626 (N_36626,N_20658,N_24101);
and U36627 (N_36627,N_20069,N_24840);
nand U36628 (N_36628,N_20655,N_28984);
nand U36629 (N_36629,N_29136,N_29257);
or U36630 (N_36630,N_20754,N_26556);
nor U36631 (N_36631,N_21485,N_27474);
and U36632 (N_36632,N_29120,N_22296);
nor U36633 (N_36633,N_28195,N_29606);
nor U36634 (N_36634,N_21153,N_29484);
and U36635 (N_36635,N_27836,N_21250);
nand U36636 (N_36636,N_21705,N_26163);
nor U36637 (N_36637,N_28813,N_24471);
nor U36638 (N_36638,N_27655,N_20128);
nand U36639 (N_36639,N_24915,N_25217);
nand U36640 (N_36640,N_22509,N_21367);
or U36641 (N_36641,N_27899,N_29721);
nand U36642 (N_36642,N_27903,N_28458);
or U36643 (N_36643,N_21869,N_21406);
nand U36644 (N_36644,N_21226,N_29642);
or U36645 (N_36645,N_29495,N_23473);
nor U36646 (N_36646,N_20591,N_25316);
and U36647 (N_36647,N_25477,N_26336);
nand U36648 (N_36648,N_25064,N_21117);
nor U36649 (N_36649,N_27686,N_20091);
xor U36650 (N_36650,N_27247,N_21053);
or U36651 (N_36651,N_22458,N_25411);
nor U36652 (N_36652,N_28050,N_27341);
nand U36653 (N_36653,N_25083,N_24859);
and U36654 (N_36654,N_25603,N_29472);
or U36655 (N_36655,N_27298,N_23925);
nand U36656 (N_36656,N_20187,N_21523);
and U36657 (N_36657,N_24982,N_23650);
or U36658 (N_36658,N_22947,N_27055);
nand U36659 (N_36659,N_26428,N_25345);
or U36660 (N_36660,N_28463,N_21100);
nor U36661 (N_36661,N_23570,N_28395);
and U36662 (N_36662,N_27575,N_24361);
or U36663 (N_36663,N_20118,N_20021);
nand U36664 (N_36664,N_28626,N_25605);
nor U36665 (N_36665,N_26670,N_22178);
or U36666 (N_36666,N_24956,N_27446);
nand U36667 (N_36667,N_26346,N_27781);
xor U36668 (N_36668,N_26646,N_28361);
xnor U36669 (N_36669,N_27721,N_20150);
nor U36670 (N_36670,N_22306,N_28003);
nor U36671 (N_36671,N_28492,N_26839);
xor U36672 (N_36672,N_25919,N_26516);
and U36673 (N_36673,N_27470,N_26990);
and U36674 (N_36674,N_25760,N_27689);
nor U36675 (N_36675,N_27922,N_23920);
nor U36676 (N_36676,N_25852,N_29773);
xnor U36677 (N_36677,N_29402,N_26206);
and U36678 (N_36678,N_21600,N_25434);
and U36679 (N_36679,N_28912,N_22041);
or U36680 (N_36680,N_25935,N_27545);
and U36681 (N_36681,N_24533,N_28405);
or U36682 (N_36682,N_24492,N_24153);
nand U36683 (N_36683,N_28397,N_22717);
or U36684 (N_36684,N_29959,N_20243);
and U36685 (N_36685,N_27217,N_23866);
nor U36686 (N_36686,N_27342,N_22467);
or U36687 (N_36687,N_20740,N_21192);
or U36688 (N_36688,N_26583,N_22270);
nor U36689 (N_36689,N_23748,N_28583);
nand U36690 (N_36690,N_23703,N_29455);
xor U36691 (N_36691,N_23244,N_20973);
xor U36692 (N_36692,N_21452,N_28924);
nor U36693 (N_36693,N_21512,N_20258);
nor U36694 (N_36694,N_21090,N_27147);
nor U36695 (N_36695,N_26578,N_20823);
nor U36696 (N_36696,N_26750,N_29794);
nor U36697 (N_36697,N_22485,N_26481);
nand U36698 (N_36698,N_27964,N_28873);
and U36699 (N_36699,N_27429,N_21211);
nand U36700 (N_36700,N_25519,N_28192);
xnor U36701 (N_36701,N_25873,N_28111);
nor U36702 (N_36702,N_24311,N_23254);
nor U36703 (N_36703,N_24027,N_26275);
nand U36704 (N_36704,N_23642,N_29236);
nand U36705 (N_36705,N_22080,N_29453);
or U36706 (N_36706,N_25166,N_24011);
or U36707 (N_36707,N_29811,N_25101);
nand U36708 (N_36708,N_22925,N_20534);
nand U36709 (N_36709,N_26449,N_20872);
xnor U36710 (N_36710,N_21693,N_22847);
or U36711 (N_36711,N_21125,N_21191);
nand U36712 (N_36712,N_25411,N_20286);
and U36713 (N_36713,N_27514,N_29448);
nand U36714 (N_36714,N_25182,N_29912);
nand U36715 (N_36715,N_24403,N_29735);
or U36716 (N_36716,N_25439,N_27874);
xor U36717 (N_36717,N_20644,N_26731);
nand U36718 (N_36718,N_29367,N_25227);
or U36719 (N_36719,N_28093,N_23408);
nand U36720 (N_36720,N_29128,N_26948);
or U36721 (N_36721,N_20398,N_20151);
or U36722 (N_36722,N_26868,N_21297);
nand U36723 (N_36723,N_25274,N_23451);
or U36724 (N_36724,N_27354,N_21674);
nand U36725 (N_36725,N_23554,N_28276);
nand U36726 (N_36726,N_29162,N_21864);
and U36727 (N_36727,N_24672,N_29093);
and U36728 (N_36728,N_21910,N_21879);
or U36729 (N_36729,N_27145,N_27702);
and U36730 (N_36730,N_27547,N_22157);
xor U36731 (N_36731,N_28505,N_23781);
nor U36732 (N_36732,N_25622,N_29012);
or U36733 (N_36733,N_22934,N_23815);
nand U36734 (N_36734,N_26020,N_21489);
nor U36735 (N_36735,N_23836,N_22434);
nand U36736 (N_36736,N_23572,N_26134);
xnor U36737 (N_36737,N_22892,N_20406);
nor U36738 (N_36738,N_26307,N_24574);
xnor U36739 (N_36739,N_28741,N_27711);
or U36740 (N_36740,N_29915,N_24613);
or U36741 (N_36741,N_27676,N_29847);
nand U36742 (N_36742,N_25219,N_24051);
or U36743 (N_36743,N_20458,N_27513);
nand U36744 (N_36744,N_22611,N_25155);
nand U36745 (N_36745,N_27826,N_23858);
and U36746 (N_36746,N_24257,N_23335);
or U36747 (N_36747,N_23987,N_26052);
or U36748 (N_36748,N_27440,N_22254);
nand U36749 (N_36749,N_24405,N_27032);
or U36750 (N_36750,N_24803,N_25862);
and U36751 (N_36751,N_22157,N_23954);
nor U36752 (N_36752,N_26885,N_25288);
or U36753 (N_36753,N_23604,N_21121);
nor U36754 (N_36754,N_26510,N_23482);
and U36755 (N_36755,N_25921,N_23684);
or U36756 (N_36756,N_28356,N_28949);
and U36757 (N_36757,N_23473,N_25633);
and U36758 (N_36758,N_23086,N_24141);
or U36759 (N_36759,N_25793,N_24463);
nor U36760 (N_36760,N_22706,N_29818);
and U36761 (N_36761,N_21564,N_29621);
or U36762 (N_36762,N_26101,N_25484);
nor U36763 (N_36763,N_21103,N_28620);
nor U36764 (N_36764,N_23685,N_24512);
and U36765 (N_36765,N_21486,N_25991);
or U36766 (N_36766,N_28703,N_29092);
and U36767 (N_36767,N_22738,N_20081);
or U36768 (N_36768,N_20010,N_28113);
or U36769 (N_36769,N_20141,N_23401);
and U36770 (N_36770,N_23503,N_20842);
nor U36771 (N_36771,N_28135,N_21153);
or U36772 (N_36772,N_24549,N_23560);
nand U36773 (N_36773,N_23122,N_29465);
and U36774 (N_36774,N_27883,N_29363);
xor U36775 (N_36775,N_24935,N_23301);
and U36776 (N_36776,N_21331,N_29658);
nand U36777 (N_36777,N_24064,N_20844);
nor U36778 (N_36778,N_28206,N_23477);
nand U36779 (N_36779,N_24441,N_26731);
nor U36780 (N_36780,N_29758,N_28780);
and U36781 (N_36781,N_22061,N_24508);
and U36782 (N_36782,N_28027,N_23826);
xnor U36783 (N_36783,N_20065,N_28151);
and U36784 (N_36784,N_23977,N_28701);
nor U36785 (N_36785,N_24666,N_20229);
nand U36786 (N_36786,N_20722,N_23376);
and U36787 (N_36787,N_27994,N_26279);
nor U36788 (N_36788,N_22313,N_25124);
and U36789 (N_36789,N_21220,N_26027);
nand U36790 (N_36790,N_21464,N_22279);
nand U36791 (N_36791,N_22113,N_23654);
nand U36792 (N_36792,N_27560,N_27069);
nand U36793 (N_36793,N_24184,N_24653);
xnor U36794 (N_36794,N_25344,N_22008);
nor U36795 (N_36795,N_23103,N_29942);
nor U36796 (N_36796,N_20192,N_20982);
and U36797 (N_36797,N_27817,N_27631);
nor U36798 (N_36798,N_26340,N_26552);
nand U36799 (N_36799,N_20284,N_28445);
or U36800 (N_36800,N_22662,N_23400);
nand U36801 (N_36801,N_22603,N_22433);
nand U36802 (N_36802,N_21097,N_28826);
or U36803 (N_36803,N_20002,N_25761);
and U36804 (N_36804,N_24677,N_28933);
nor U36805 (N_36805,N_29727,N_28031);
nor U36806 (N_36806,N_27430,N_25726);
nand U36807 (N_36807,N_28835,N_26536);
and U36808 (N_36808,N_24584,N_20212);
or U36809 (N_36809,N_24230,N_27838);
or U36810 (N_36810,N_28490,N_21273);
and U36811 (N_36811,N_20091,N_29812);
and U36812 (N_36812,N_24266,N_29413);
nor U36813 (N_36813,N_23885,N_29018);
or U36814 (N_36814,N_22432,N_27277);
xor U36815 (N_36815,N_25829,N_21084);
nand U36816 (N_36816,N_23889,N_27489);
nand U36817 (N_36817,N_23827,N_20588);
and U36818 (N_36818,N_24900,N_22227);
or U36819 (N_36819,N_28630,N_23996);
or U36820 (N_36820,N_21014,N_22023);
and U36821 (N_36821,N_21244,N_28101);
or U36822 (N_36822,N_28073,N_29330);
nand U36823 (N_36823,N_28331,N_28586);
nor U36824 (N_36824,N_24786,N_20392);
and U36825 (N_36825,N_21506,N_29820);
nor U36826 (N_36826,N_26898,N_29961);
and U36827 (N_36827,N_20229,N_23681);
or U36828 (N_36828,N_20092,N_27246);
xnor U36829 (N_36829,N_25049,N_22634);
nand U36830 (N_36830,N_25987,N_23768);
nand U36831 (N_36831,N_22850,N_26221);
nor U36832 (N_36832,N_21978,N_28588);
nor U36833 (N_36833,N_22828,N_21660);
nor U36834 (N_36834,N_24659,N_25193);
nor U36835 (N_36835,N_24040,N_26595);
nor U36836 (N_36836,N_29436,N_22952);
nand U36837 (N_36837,N_24134,N_25667);
nand U36838 (N_36838,N_29362,N_24038);
or U36839 (N_36839,N_27946,N_29910);
nor U36840 (N_36840,N_20947,N_20977);
xnor U36841 (N_36841,N_25718,N_29796);
nand U36842 (N_36842,N_24918,N_25102);
nor U36843 (N_36843,N_25156,N_24264);
nand U36844 (N_36844,N_21190,N_26099);
nor U36845 (N_36845,N_23170,N_20397);
or U36846 (N_36846,N_20719,N_27510);
or U36847 (N_36847,N_25980,N_26790);
or U36848 (N_36848,N_29025,N_22444);
nand U36849 (N_36849,N_22925,N_27815);
nor U36850 (N_36850,N_27774,N_25151);
and U36851 (N_36851,N_22993,N_23205);
nand U36852 (N_36852,N_29396,N_25507);
and U36853 (N_36853,N_21267,N_23658);
nor U36854 (N_36854,N_23935,N_20749);
nor U36855 (N_36855,N_23913,N_22374);
xnor U36856 (N_36856,N_26331,N_22133);
and U36857 (N_36857,N_27157,N_23912);
nor U36858 (N_36858,N_25067,N_24995);
nand U36859 (N_36859,N_26042,N_25990);
nor U36860 (N_36860,N_27988,N_22504);
and U36861 (N_36861,N_27301,N_24190);
and U36862 (N_36862,N_27472,N_20971);
nand U36863 (N_36863,N_25042,N_23726);
nand U36864 (N_36864,N_24840,N_25113);
and U36865 (N_36865,N_25869,N_23183);
and U36866 (N_36866,N_21023,N_25709);
nand U36867 (N_36867,N_21812,N_26582);
nand U36868 (N_36868,N_24542,N_26505);
or U36869 (N_36869,N_20935,N_20545);
nand U36870 (N_36870,N_25709,N_23143);
or U36871 (N_36871,N_21697,N_22192);
or U36872 (N_36872,N_20397,N_26134);
nor U36873 (N_36873,N_22392,N_20643);
and U36874 (N_36874,N_20406,N_29421);
nor U36875 (N_36875,N_23698,N_29081);
and U36876 (N_36876,N_23978,N_29205);
nand U36877 (N_36877,N_26204,N_25862);
or U36878 (N_36878,N_21503,N_26869);
or U36879 (N_36879,N_24165,N_25882);
xor U36880 (N_36880,N_23734,N_20628);
nor U36881 (N_36881,N_24646,N_28232);
nor U36882 (N_36882,N_28103,N_26143);
or U36883 (N_36883,N_21569,N_26804);
or U36884 (N_36884,N_28918,N_27997);
or U36885 (N_36885,N_29891,N_23179);
and U36886 (N_36886,N_27034,N_27811);
nand U36887 (N_36887,N_21445,N_23475);
and U36888 (N_36888,N_22721,N_24129);
nor U36889 (N_36889,N_29096,N_28236);
and U36890 (N_36890,N_22160,N_21837);
or U36891 (N_36891,N_23201,N_22931);
or U36892 (N_36892,N_25598,N_25025);
nand U36893 (N_36893,N_23453,N_23340);
nand U36894 (N_36894,N_26060,N_21256);
and U36895 (N_36895,N_26366,N_28879);
nand U36896 (N_36896,N_29527,N_26692);
nor U36897 (N_36897,N_20923,N_20524);
and U36898 (N_36898,N_20434,N_21502);
nor U36899 (N_36899,N_22284,N_24891);
or U36900 (N_36900,N_29693,N_20109);
and U36901 (N_36901,N_20404,N_22335);
and U36902 (N_36902,N_22987,N_24585);
and U36903 (N_36903,N_29896,N_23799);
nand U36904 (N_36904,N_29583,N_21026);
nand U36905 (N_36905,N_22789,N_21901);
and U36906 (N_36906,N_25068,N_21033);
or U36907 (N_36907,N_29445,N_24915);
nand U36908 (N_36908,N_20247,N_24148);
nand U36909 (N_36909,N_27987,N_21537);
nand U36910 (N_36910,N_25444,N_26335);
nand U36911 (N_36911,N_22643,N_22830);
nor U36912 (N_36912,N_26207,N_21642);
and U36913 (N_36913,N_24767,N_21808);
or U36914 (N_36914,N_21641,N_25117);
nand U36915 (N_36915,N_24341,N_23328);
nand U36916 (N_36916,N_26006,N_20585);
or U36917 (N_36917,N_24142,N_29976);
nor U36918 (N_36918,N_23017,N_22777);
nand U36919 (N_36919,N_23808,N_28526);
xor U36920 (N_36920,N_23375,N_27843);
or U36921 (N_36921,N_24727,N_29466);
or U36922 (N_36922,N_29256,N_21700);
xnor U36923 (N_36923,N_23114,N_25609);
nor U36924 (N_36924,N_29134,N_28139);
xnor U36925 (N_36925,N_21922,N_26455);
nor U36926 (N_36926,N_21061,N_28461);
and U36927 (N_36927,N_26965,N_24167);
nand U36928 (N_36928,N_22062,N_26265);
and U36929 (N_36929,N_27635,N_27156);
nor U36930 (N_36930,N_21108,N_22810);
or U36931 (N_36931,N_23102,N_22790);
or U36932 (N_36932,N_23855,N_24487);
nand U36933 (N_36933,N_20025,N_21290);
nand U36934 (N_36934,N_23416,N_20817);
and U36935 (N_36935,N_23359,N_23096);
nand U36936 (N_36936,N_28179,N_25116);
and U36937 (N_36937,N_29818,N_26932);
nand U36938 (N_36938,N_28423,N_23397);
or U36939 (N_36939,N_29673,N_27985);
or U36940 (N_36940,N_27642,N_21157);
or U36941 (N_36941,N_29500,N_24356);
or U36942 (N_36942,N_29736,N_25764);
nor U36943 (N_36943,N_24628,N_24149);
and U36944 (N_36944,N_24217,N_23849);
or U36945 (N_36945,N_25112,N_28695);
and U36946 (N_36946,N_24103,N_29874);
or U36947 (N_36947,N_29934,N_23982);
nand U36948 (N_36948,N_21059,N_25291);
xnor U36949 (N_36949,N_20662,N_29598);
and U36950 (N_36950,N_27052,N_20248);
nor U36951 (N_36951,N_21917,N_23328);
or U36952 (N_36952,N_24112,N_28437);
nor U36953 (N_36953,N_24767,N_21733);
and U36954 (N_36954,N_26518,N_22931);
or U36955 (N_36955,N_23046,N_27223);
and U36956 (N_36956,N_20418,N_24587);
nor U36957 (N_36957,N_21738,N_23824);
nand U36958 (N_36958,N_21724,N_22839);
or U36959 (N_36959,N_20845,N_27846);
and U36960 (N_36960,N_28916,N_27904);
and U36961 (N_36961,N_27529,N_28376);
nor U36962 (N_36962,N_20894,N_20512);
and U36963 (N_36963,N_23833,N_22007);
and U36964 (N_36964,N_25639,N_24005);
nand U36965 (N_36965,N_25058,N_29266);
and U36966 (N_36966,N_27407,N_21029);
or U36967 (N_36967,N_21930,N_24878);
or U36968 (N_36968,N_22583,N_27140);
nor U36969 (N_36969,N_28747,N_21274);
nand U36970 (N_36970,N_28060,N_25432);
and U36971 (N_36971,N_22844,N_26696);
xnor U36972 (N_36972,N_20793,N_23302);
nor U36973 (N_36973,N_23970,N_22476);
or U36974 (N_36974,N_23078,N_21297);
nor U36975 (N_36975,N_26936,N_22142);
or U36976 (N_36976,N_27864,N_27914);
and U36977 (N_36977,N_23940,N_22195);
nand U36978 (N_36978,N_27724,N_28343);
nand U36979 (N_36979,N_23683,N_24962);
nor U36980 (N_36980,N_21595,N_25278);
or U36981 (N_36981,N_20414,N_20741);
and U36982 (N_36982,N_22317,N_27507);
nor U36983 (N_36983,N_27983,N_25975);
or U36984 (N_36984,N_26858,N_25003);
xnor U36985 (N_36985,N_23573,N_24326);
or U36986 (N_36986,N_23741,N_21905);
and U36987 (N_36987,N_21354,N_26777);
nor U36988 (N_36988,N_23777,N_25548);
or U36989 (N_36989,N_22958,N_21669);
or U36990 (N_36990,N_28716,N_23624);
or U36991 (N_36991,N_27037,N_26508);
nand U36992 (N_36992,N_26093,N_21740);
nand U36993 (N_36993,N_23087,N_26231);
nand U36994 (N_36994,N_29025,N_28342);
nor U36995 (N_36995,N_21496,N_24846);
xnor U36996 (N_36996,N_22137,N_21407);
nor U36997 (N_36997,N_29879,N_20351);
or U36998 (N_36998,N_26527,N_20900);
or U36999 (N_36999,N_24764,N_21237);
and U37000 (N_37000,N_27205,N_26895);
nand U37001 (N_37001,N_26295,N_27106);
or U37002 (N_37002,N_26769,N_26499);
and U37003 (N_37003,N_26862,N_20382);
or U37004 (N_37004,N_20905,N_29634);
xnor U37005 (N_37005,N_23134,N_27673);
nand U37006 (N_37006,N_26636,N_25879);
and U37007 (N_37007,N_20624,N_23213);
nand U37008 (N_37008,N_27267,N_29541);
and U37009 (N_37009,N_22537,N_25959);
or U37010 (N_37010,N_27562,N_24431);
or U37011 (N_37011,N_20707,N_25798);
nor U37012 (N_37012,N_27503,N_29596);
or U37013 (N_37013,N_29892,N_29415);
or U37014 (N_37014,N_25329,N_24811);
nor U37015 (N_37015,N_24401,N_28620);
or U37016 (N_37016,N_26946,N_22847);
nor U37017 (N_37017,N_28392,N_28333);
nand U37018 (N_37018,N_27164,N_25358);
or U37019 (N_37019,N_21047,N_24249);
or U37020 (N_37020,N_25949,N_24039);
nand U37021 (N_37021,N_24291,N_24284);
and U37022 (N_37022,N_29005,N_22919);
nand U37023 (N_37023,N_21144,N_27158);
and U37024 (N_37024,N_21666,N_21829);
nand U37025 (N_37025,N_28270,N_28831);
xor U37026 (N_37026,N_20268,N_22638);
nand U37027 (N_37027,N_28046,N_26677);
or U37028 (N_37028,N_24708,N_29917);
nor U37029 (N_37029,N_24424,N_20303);
and U37030 (N_37030,N_27501,N_20028);
xnor U37031 (N_37031,N_25876,N_28228);
and U37032 (N_37032,N_22008,N_23511);
and U37033 (N_37033,N_26569,N_27931);
and U37034 (N_37034,N_25817,N_22029);
nand U37035 (N_37035,N_25542,N_25533);
or U37036 (N_37036,N_29591,N_25011);
or U37037 (N_37037,N_25123,N_27693);
nand U37038 (N_37038,N_20827,N_24915);
and U37039 (N_37039,N_26459,N_20723);
nor U37040 (N_37040,N_20741,N_21799);
or U37041 (N_37041,N_26962,N_28906);
nor U37042 (N_37042,N_23643,N_22137);
xnor U37043 (N_37043,N_26280,N_22018);
or U37044 (N_37044,N_26642,N_22964);
or U37045 (N_37045,N_28969,N_24642);
or U37046 (N_37046,N_26395,N_28284);
or U37047 (N_37047,N_25301,N_23865);
nor U37048 (N_37048,N_21726,N_29129);
or U37049 (N_37049,N_26115,N_22467);
xor U37050 (N_37050,N_26667,N_22918);
and U37051 (N_37051,N_22404,N_25991);
xnor U37052 (N_37052,N_21500,N_24390);
nand U37053 (N_37053,N_26973,N_29182);
nand U37054 (N_37054,N_25177,N_20192);
or U37055 (N_37055,N_29387,N_24939);
and U37056 (N_37056,N_20800,N_25050);
nor U37057 (N_37057,N_25696,N_26115);
nand U37058 (N_37058,N_29120,N_29618);
nor U37059 (N_37059,N_20515,N_23769);
xor U37060 (N_37060,N_29745,N_25416);
nand U37061 (N_37061,N_25345,N_20555);
or U37062 (N_37062,N_21006,N_25604);
nand U37063 (N_37063,N_20006,N_24613);
and U37064 (N_37064,N_23407,N_29883);
and U37065 (N_37065,N_20715,N_27793);
nand U37066 (N_37066,N_23639,N_26994);
and U37067 (N_37067,N_21562,N_25638);
nand U37068 (N_37068,N_27304,N_25841);
xor U37069 (N_37069,N_21749,N_20910);
or U37070 (N_37070,N_21436,N_27907);
and U37071 (N_37071,N_21714,N_27640);
or U37072 (N_37072,N_20291,N_28993);
nor U37073 (N_37073,N_22349,N_23136);
nor U37074 (N_37074,N_21765,N_25580);
nand U37075 (N_37075,N_22768,N_20724);
xor U37076 (N_37076,N_28439,N_27776);
nand U37077 (N_37077,N_27399,N_25677);
or U37078 (N_37078,N_20140,N_21234);
or U37079 (N_37079,N_29669,N_21371);
xnor U37080 (N_37080,N_21869,N_21771);
or U37081 (N_37081,N_22490,N_26702);
nor U37082 (N_37082,N_25341,N_24761);
or U37083 (N_37083,N_24510,N_29402);
nor U37084 (N_37084,N_26475,N_23800);
xnor U37085 (N_37085,N_29415,N_29199);
nor U37086 (N_37086,N_21996,N_21852);
nor U37087 (N_37087,N_24404,N_24467);
nand U37088 (N_37088,N_28464,N_26775);
nor U37089 (N_37089,N_24903,N_22701);
nand U37090 (N_37090,N_20468,N_23442);
or U37091 (N_37091,N_26578,N_26654);
or U37092 (N_37092,N_20295,N_20315);
and U37093 (N_37093,N_27299,N_26795);
and U37094 (N_37094,N_21742,N_28480);
and U37095 (N_37095,N_24689,N_20949);
or U37096 (N_37096,N_26966,N_28945);
nand U37097 (N_37097,N_21281,N_21876);
nand U37098 (N_37098,N_24772,N_25729);
nand U37099 (N_37099,N_23635,N_20893);
nor U37100 (N_37100,N_27233,N_24645);
and U37101 (N_37101,N_22635,N_21825);
and U37102 (N_37102,N_25162,N_29623);
nand U37103 (N_37103,N_27445,N_22591);
nor U37104 (N_37104,N_21528,N_20233);
and U37105 (N_37105,N_25845,N_21359);
nor U37106 (N_37106,N_24355,N_22591);
and U37107 (N_37107,N_23130,N_22115);
and U37108 (N_37108,N_20290,N_26718);
nor U37109 (N_37109,N_26414,N_21528);
or U37110 (N_37110,N_27955,N_24531);
or U37111 (N_37111,N_22996,N_23642);
nor U37112 (N_37112,N_24482,N_27648);
and U37113 (N_37113,N_28595,N_25260);
nand U37114 (N_37114,N_28807,N_25117);
and U37115 (N_37115,N_29144,N_26882);
nor U37116 (N_37116,N_21671,N_20908);
or U37117 (N_37117,N_25441,N_24303);
or U37118 (N_37118,N_22179,N_29760);
nor U37119 (N_37119,N_20017,N_22469);
and U37120 (N_37120,N_29299,N_25291);
nand U37121 (N_37121,N_20147,N_20105);
nor U37122 (N_37122,N_24570,N_24477);
nor U37123 (N_37123,N_24865,N_25487);
xnor U37124 (N_37124,N_21320,N_28766);
nor U37125 (N_37125,N_22103,N_21708);
or U37126 (N_37126,N_20135,N_25767);
and U37127 (N_37127,N_27583,N_20003);
nand U37128 (N_37128,N_24610,N_28967);
and U37129 (N_37129,N_29768,N_29334);
nand U37130 (N_37130,N_25614,N_29037);
and U37131 (N_37131,N_29015,N_25119);
xor U37132 (N_37132,N_22798,N_22749);
or U37133 (N_37133,N_25301,N_20854);
nand U37134 (N_37134,N_27645,N_29048);
nor U37135 (N_37135,N_24067,N_21836);
and U37136 (N_37136,N_21900,N_22673);
nand U37137 (N_37137,N_22335,N_22169);
and U37138 (N_37138,N_20615,N_25612);
and U37139 (N_37139,N_24811,N_28766);
or U37140 (N_37140,N_29814,N_23150);
or U37141 (N_37141,N_25814,N_23324);
or U37142 (N_37142,N_27598,N_23715);
or U37143 (N_37143,N_23790,N_23206);
or U37144 (N_37144,N_27532,N_26637);
and U37145 (N_37145,N_25483,N_29195);
and U37146 (N_37146,N_27146,N_28632);
nor U37147 (N_37147,N_22544,N_22508);
nor U37148 (N_37148,N_28388,N_26954);
nand U37149 (N_37149,N_20367,N_27950);
or U37150 (N_37150,N_25544,N_22322);
nand U37151 (N_37151,N_23208,N_20146);
nor U37152 (N_37152,N_29139,N_20479);
nand U37153 (N_37153,N_29952,N_24182);
or U37154 (N_37154,N_29381,N_21263);
and U37155 (N_37155,N_25072,N_26759);
nor U37156 (N_37156,N_25774,N_23989);
or U37157 (N_37157,N_28036,N_24099);
nand U37158 (N_37158,N_28368,N_26684);
and U37159 (N_37159,N_29746,N_21290);
and U37160 (N_37160,N_25565,N_27187);
and U37161 (N_37161,N_20798,N_22046);
xor U37162 (N_37162,N_29809,N_25416);
nor U37163 (N_37163,N_26626,N_20396);
nand U37164 (N_37164,N_20098,N_28819);
nand U37165 (N_37165,N_21488,N_27098);
nor U37166 (N_37166,N_25335,N_26696);
nor U37167 (N_37167,N_21298,N_27053);
nand U37168 (N_37168,N_22459,N_29173);
nor U37169 (N_37169,N_26674,N_21569);
nor U37170 (N_37170,N_27035,N_29017);
nor U37171 (N_37171,N_25018,N_21358);
nand U37172 (N_37172,N_29228,N_27660);
nand U37173 (N_37173,N_25693,N_25610);
xnor U37174 (N_37174,N_28207,N_23815);
and U37175 (N_37175,N_24624,N_24552);
nor U37176 (N_37176,N_28582,N_29532);
nor U37177 (N_37177,N_22262,N_22532);
nor U37178 (N_37178,N_24341,N_29034);
and U37179 (N_37179,N_26386,N_20641);
nor U37180 (N_37180,N_20941,N_29018);
nand U37181 (N_37181,N_24303,N_29679);
or U37182 (N_37182,N_20102,N_29580);
and U37183 (N_37183,N_25227,N_23156);
or U37184 (N_37184,N_24977,N_28518);
xnor U37185 (N_37185,N_26960,N_29313);
and U37186 (N_37186,N_28156,N_24800);
and U37187 (N_37187,N_29651,N_22896);
and U37188 (N_37188,N_28762,N_26582);
nand U37189 (N_37189,N_28200,N_24691);
nor U37190 (N_37190,N_26161,N_26503);
nand U37191 (N_37191,N_27597,N_23668);
nand U37192 (N_37192,N_24591,N_21154);
xor U37193 (N_37193,N_24809,N_23305);
and U37194 (N_37194,N_21469,N_21708);
nor U37195 (N_37195,N_23382,N_20751);
or U37196 (N_37196,N_29609,N_25613);
xnor U37197 (N_37197,N_26696,N_21704);
nor U37198 (N_37198,N_27554,N_22233);
nor U37199 (N_37199,N_26684,N_28639);
or U37200 (N_37200,N_29494,N_23749);
xor U37201 (N_37201,N_29200,N_26769);
nor U37202 (N_37202,N_25075,N_24849);
nand U37203 (N_37203,N_25384,N_23858);
or U37204 (N_37204,N_26152,N_23497);
and U37205 (N_37205,N_29182,N_23830);
and U37206 (N_37206,N_25009,N_20552);
or U37207 (N_37207,N_22286,N_22527);
nor U37208 (N_37208,N_21787,N_21637);
nand U37209 (N_37209,N_21753,N_23359);
or U37210 (N_37210,N_29928,N_25538);
xor U37211 (N_37211,N_27823,N_22168);
or U37212 (N_37212,N_24319,N_21480);
nand U37213 (N_37213,N_24317,N_29140);
or U37214 (N_37214,N_20587,N_27207);
or U37215 (N_37215,N_27717,N_28541);
xor U37216 (N_37216,N_25582,N_21140);
or U37217 (N_37217,N_23266,N_22248);
nor U37218 (N_37218,N_25101,N_21743);
nand U37219 (N_37219,N_21448,N_26128);
nor U37220 (N_37220,N_25575,N_29983);
or U37221 (N_37221,N_29850,N_26503);
nand U37222 (N_37222,N_24855,N_21031);
nand U37223 (N_37223,N_21875,N_25681);
or U37224 (N_37224,N_20330,N_29450);
or U37225 (N_37225,N_20433,N_28425);
xnor U37226 (N_37226,N_21412,N_27570);
nand U37227 (N_37227,N_26736,N_24680);
or U37228 (N_37228,N_25354,N_29191);
nor U37229 (N_37229,N_23978,N_29519);
or U37230 (N_37230,N_28518,N_29295);
nor U37231 (N_37231,N_22024,N_28395);
or U37232 (N_37232,N_28193,N_21770);
nand U37233 (N_37233,N_24046,N_24806);
or U37234 (N_37234,N_27944,N_26687);
and U37235 (N_37235,N_22747,N_27302);
or U37236 (N_37236,N_20420,N_23808);
or U37237 (N_37237,N_28476,N_28405);
nor U37238 (N_37238,N_21722,N_25610);
nor U37239 (N_37239,N_27432,N_29871);
or U37240 (N_37240,N_24602,N_25796);
nor U37241 (N_37241,N_25797,N_24527);
nand U37242 (N_37242,N_25867,N_25486);
or U37243 (N_37243,N_29783,N_24131);
nand U37244 (N_37244,N_20045,N_21943);
and U37245 (N_37245,N_23032,N_24372);
nand U37246 (N_37246,N_28179,N_20977);
nor U37247 (N_37247,N_23445,N_29486);
nand U37248 (N_37248,N_27545,N_22481);
nor U37249 (N_37249,N_20704,N_23214);
xnor U37250 (N_37250,N_21630,N_23149);
xnor U37251 (N_37251,N_24179,N_26021);
nor U37252 (N_37252,N_21907,N_25749);
nand U37253 (N_37253,N_21208,N_20830);
and U37254 (N_37254,N_22648,N_28760);
nand U37255 (N_37255,N_20693,N_29898);
nor U37256 (N_37256,N_22601,N_27854);
nand U37257 (N_37257,N_26794,N_27530);
or U37258 (N_37258,N_29280,N_24567);
nor U37259 (N_37259,N_23695,N_20798);
or U37260 (N_37260,N_21911,N_23451);
or U37261 (N_37261,N_24135,N_26973);
or U37262 (N_37262,N_20162,N_24095);
nor U37263 (N_37263,N_20310,N_25893);
and U37264 (N_37264,N_24100,N_27166);
nor U37265 (N_37265,N_21730,N_25606);
or U37266 (N_37266,N_22186,N_20445);
nor U37267 (N_37267,N_26763,N_24931);
or U37268 (N_37268,N_20846,N_20594);
and U37269 (N_37269,N_26515,N_23680);
nor U37270 (N_37270,N_28484,N_25984);
nand U37271 (N_37271,N_27944,N_22539);
xor U37272 (N_37272,N_23013,N_23272);
or U37273 (N_37273,N_21467,N_23534);
nor U37274 (N_37274,N_27646,N_24178);
xor U37275 (N_37275,N_27669,N_20637);
nand U37276 (N_37276,N_22865,N_28701);
nand U37277 (N_37277,N_20773,N_22780);
nor U37278 (N_37278,N_23183,N_28952);
or U37279 (N_37279,N_25674,N_25995);
xnor U37280 (N_37280,N_27574,N_29903);
nor U37281 (N_37281,N_29616,N_20683);
nor U37282 (N_37282,N_21635,N_29756);
or U37283 (N_37283,N_27391,N_29897);
or U37284 (N_37284,N_23874,N_22002);
and U37285 (N_37285,N_22876,N_21637);
nand U37286 (N_37286,N_21910,N_26029);
or U37287 (N_37287,N_24035,N_27737);
nor U37288 (N_37288,N_20971,N_23492);
or U37289 (N_37289,N_21517,N_27155);
and U37290 (N_37290,N_24601,N_26768);
or U37291 (N_37291,N_23045,N_26994);
nor U37292 (N_37292,N_28234,N_28270);
nor U37293 (N_37293,N_21349,N_21232);
and U37294 (N_37294,N_22812,N_22851);
nand U37295 (N_37295,N_29129,N_24259);
or U37296 (N_37296,N_21495,N_26052);
nand U37297 (N_37297,N_26152,N_23821);
or U37298 (N_37298,N_20926,N_27421);
or U37299 (N_37299,N_22910,N_28454);
xor U37300 (N_37300,N_20887,N_21602);
nand U37301 (N_37301,N_24866,N_23501);
or U37302 (N_37302,N_20242,N_25907);
nor U37303 (N_37303,N_28431,N_29682);
and U37304 (N_37304,N_28985,N_26409);
and U37305 (N_37305,N_27959,N_22310);
nor U37306 (N_37306,N_21247,N_21301);
and U37307 (N_37307,N_23478,N_24761);
and U37308 (N_37308,N_26025,N_26825);
nand U37309 (N_37309,N_20944,N_28926);
nor U37310 (N_37310,N_20187,N_24909);
or U37311 (N_37311,N_23964,N_25353);
nor U37312 (N_37312,N_23360,N_23723);
or U37313 (N_37313,N_20118,N_26588);
or U37314 (N_37314,N_29509,N_29837);
nand U37315 (N_37315,N_20519,N_27301);
and U37316 (N_37316,N_21876,N_28504);
xnor U37317 (N_37317,N_20516,N_20631);
nand U37318 (N_37318,N_23850,N_24271);
nand U37319 (N_37319,N_26372,N_27297);
and U37320 (N_37320,N_27519,N_21293);
xor U37321 (N_37321,N_25426,N_26273);
nor U37322 (N_37322,N_26387,N_24694);
or U37323 (N_37323,N_27275,N_23623);
and U37324 (N_37324,N_23141,N_23312);
nor U37325 (N_37325,N_29157,N_26679);
nand U37326 (N_37326,N_28217,N_28942);
and U37327 (N_37327,N_28066,N_27529);
or U37328 (N_37328,N_23543,N_23467);
and U37329 (N_37329,N_25140,N_29674);
and U37330 (N_37330,N_26743,N_28573);
nor U37331 (N_37331,N_23039,N_22182);
and U37332 (N_37332,N_29516,N_23868);
nand U37333 (N_37333,N_24836,N_28643);
nand U37334 (N_37334,N_29090,N_21701);
and U37335 (N_37335,N_28867,N_25536);
xor U37336 (N_37336,N_25990,N_25841);
and U37337 (N_37337,N_21930,N_24054);
xnor U37338 (N_37338,N_29350,N_21165);
nor U37339 (N_37339,N_22652,N_27591);
and U37340 (N_37340,N_20324,N_27655);
xnor U37341 (N_37341,N_28731,N_29779);
and U37342 (N_37342,N_24628,N_29180);
nor U37343 (N_37343,N_27148,N_20643);
nor U37344 (N_37344,N_24226,N_20695);
nor U37345 (N_37345,N_21894,N_25791);
and U37346 (N_37346,N_25126,N_26492);
nand U37347 (N_37347,N_28137,N_27336);
nor U37348 (N_37348,N_27878,N_23742);
or U37349 (N_37349,N_29768,N_25859);
nor U37350 (N_37350,N_23870,N_28548);
nor U37351 (N_37351,N_24931,N_27579);
and U37352 (N_37352,N_23604,N_22666);
nor U37353 (N_37353,N_29332,N_21036);
and U37354 (N_37354,N_24688,N_27127);
nand U37355 (N_37355,N_24388,N_20191);
nand U37356 (N_37356,N_25255,N_22988);
nor U37357 (N_37357,N_27643,N_26508);
or U37358 (N_37358,N_27520,N_25658);
nand U37359 (N_37359,N_26734,N_28556);
and U37360 (N_37360,N_28927,N_22269);
nand U37361 (N_37361,N_23312,N_26967);
nor U37362 (N_37362,N_27822,N_21838);
nand U37363 (N_37363,N_25634,N_26226);
nand U37364 (N_37364,N_22529,N_26574);
nor U37365 (N_37365,N_23194,N_26892);
nor U37366 (N_37366,N_29949,N_21044);
or U37367 (N_37367,N_20312,N_21875);
nor U37368 (N_37368,N_21466,N_27312);
and U37369 (N_37369,N_22087,N_29828);
and U37370 (N_37370,N_24288,N_26371);
nand U37371 (N_37371,N_29184,N_20972);
and U37372 (N_37372,N_23320,N_27879);
or U37373 (N_37373,N_28221,N_21609);
nor U37374 (N_37374,N_29934,N_24577);
xor U37375 (N_37375,N_21114,N_23011);
nor U37376 (N_37376,N_24632,N_22596);
nand U37377 (N_37377,N_24339,N_24831);
or U37378 (N_37378,N_20860,N_20388);
nand U37379 (N_37379,N_27325,N_20146);
xor U37380 (N_37380,N_26215,N_21279);
or U37381 (N_37381,N_21353,N_20484);
nor U37382 (N_37382,N_22646,N_20848);
nand U37383 (N_37383,N_29735,N_25945);
xnor U37384 (N_37384,N_23245,N_23229);
and U37385 (N_37385,N_23276,N_20624);
and U37386 (N_37386,N_28130,N_27860);
or U37387 (N_37387,N_25630,N_21508);
or U37388 (N_37388,N_23759,N_23780);
nor U37389 (N_37389,N_21525,N_29644);
xor U37390 (N_37390,N_21056,N_22428);
and U37391 (N_37391,N_25011,N_20587);
or U37392 (N_37392,N_23633,N_28120);
nor U37393 (N_37393,N_29377,N_20074);
nand U37394 (N_37394,N_21799,N_24022);
nor U37395 (N_37395,N_24865,N_26302);
nor U37396 (N_37396,N_29149,N_27802);
and U37397 (N_37397,N_25211,N_25400);
xnor U37398 (N_37398,N_24848,N_23199);
nand U37399 (N_37399,N_21935,N_29724);
or U37400 (N_37400,N_24382,N_25247);
and U37401 (N_37401,N_22684,N_27949);
nor U37402 (N_37402,N_24628,N_24734);
nor U37403 (N_37403,N_29663,N_22725);
or U37404 (N_37404,N_22247,N_27563);
or U37405 (N_37405,N_25716,N_21637);
or U37406 (N_37406,N_24031,N_23443);
nor U37407 (N_37407,N_29346,N_21548);
and U37408 (N_37408,N_29443,N_29278);
and U37409 (N_37409,N_24700,N_23497);
nor U37410 (N_37410,N_29716,N_22645);
xnor U37411 (N_37411,N_28802,N_20365);
or U37412 (N_37412,N_26903,N_22391);
nor U37413 (N_37413,N_22026,N_24141);
or U37414 (N_37414,N_27632,N_23457);
or U37415 (N_37415,N_25507,N_25980);
and U37416 (N_37416,N_24622,N_22329);
or U37417 (N_37417,N_25706,N_22107);
or U37418 (N_37418,N_26148,N_25352);
nor U37419 (N_37419,N_25820,N_20628);
and U37420 (N_37420,N_23620,N_22001);
or U37421 (N_37421,N_21620,N_20682);
nor U37422 (N_37422,N_23323,N_20444);
nand U37423 (N_37423,N_25703,N_25539);
and U37424 (N_37424,N_24605,N_21395);
and U37425 (N_37425,N_22001,N_28447);
or U37426 (N_37426,N_25675,N_29953);
and U37427 (N_37427,N_25675,N_25471);
nor U37428 (N_37428,N_25029,N_28579);
xnor U37429 (N_37429,N_28659,N_22185);
or U37430 (N_37430,N_25392,N_23800);
and U37431 (N_37431,N_24416,N_24920);
nor U37432 (N_37432,N_29168,N_28131);
nand U37433 (N_37433,N_26486,N_21704);
nand U37434 (N_37434,N_20303,N_21499);
nor U37435 (N_37435,N_27157,N_24617);
and U37436 (N_37436,N_28083,N_23429);
nand U37437 (N_37437,N_29133,N_25187);
xor U37438 (N_37438,N_21280,N_23736);
nand U37439 (N_37439,N_29134,N_29664);
or U37440 (N_37440,N_24307,N_27311);
and U37441 (N_37441,N_26562,N_28795);
and U37442 (N_37442,N_25123,N_26741);
nor U37443 (N_37443,N_26954,N_25579);
nand U37444 (N_37444,N_21460,N_29741);
or U37445 (N_37445,N_23807,N_26619);
nand U37446 (N_37446,N_29545,N_21147);
xor U37447 (N_37447,N_24281,N_21579);
and U37448 (N_37448,N_27635,N_24347);
nor U37449 (N_37449,N_20282,N_21581);
nand U37450 (N_37450,N_26650,N_28580);
and U37451 (N_37451,N_23963,N_24782);
or U37452 (N_37452,N_20535,N_27367);
nand U37453 (N_37453,N_20184,N_20557);
nand U37454 (N_37454,N_28314,N_25196);
or U37455 (N_37455,N_29764,N_25366);
and U37456 (N_37456,N_24654,N_21298);
and U37457 (N_37457,N_23456,N_22011);
and U37458 (N_37458,N_29547,N_24672);
nand U37459 (N_37459,N_26150,N_22597);
nand U37460 (N_37460,N_26953,N_28197);
nand U37461 (N_37461,N_22152,N_22739);
nor U37462 (N_37462,N_27952,N_22744);
and U37463 (N_37463,N_23421,N_21805);
nor U37464 (N_37464,N_27764,N_20195);
or U37465 (N_37465,N_27084,N_21943);
and U37466 (N_37466,N_28192,N_21617);
nand U37467 (N_37467,N_25315,N_29397);
nor U37468 (N_37468,N_23700,N_27629);
nand U37469 (N_37469,N_27276,N_28036);
or U37470 (N_37470,N_26726,N_23322);
nor U37471 (N_37471,N_28790,N_20850);
nor U37472 (N_37472,N_24158,N_23299);
and U37473 (N_37473,N_22952,N_28687);
nand U37474 (N_37474,N_24262,N_20121);
nor U37475 (N_37475,N_29652,N_20697);
nand U37476 (N_37476,N_26271,N_23332);
nand U37477 (N_37477,N_21504,N_20412);
or U37478 (N_37478,N_29655,N_26947);
xnor U37479 (N_37479,N_27190,N_29017);
nor U37480 (N_37480,N_25746,N_23074);
and U37481 (N_37481,N_26157,N_27078);
nand U37482 (N_37482,N_21568,N_24914);
or U37483 (N_37483,N_20643,N_20825);
or U37484 (N_37484,N_25338,N_22783);
xor U37485 (N_37485,N_20411,N_22282);
nor U37486 (N_37486,N_27832,N_28212);
nand U37487 (N_37487,N_20736,N_24134);
nor U37488 (N_37488,N_22272,N_22023);
nor U37489 (N_37489,N_29502,N_21510);
and U37490 (N_37490,N_28936,N_22344);
xor U37491 (N_37491,N_24764,N_26674);
nor U37492 (N_37492,N_28807,N_22594);
or U37493 (N_37493,N_25617,N_27970);
nor U37494 (N_37494,N_23023,N_20865);
or U37495 (N_37495,N_25407,N_24777);
or U37496 (N_37496,N_26655,N_25746);
nand U37497 (N_37497,N_25480,N_20977);
xnor U37498 (N_37498,N_28438,N_20156);
nor U37499 (N_37499,N_26238,N_20872);
and U37500 (N_37500,N_24913,N_28049);
and U37501 (N_37501,N_23729,N_29318);
and U37502 (N_37502,N_23846,N_21437);
and U37503 (N_37503,N_25200,N_20589);
or U37504 (N_37504,N_29200,N_29918);
nor U37505 (N_37505,N_24907,N_28136);
nor U37506 (N_37506,N_24958,N_26508);
nor U37507 (N_37507,N_20205,N_23722);
or U37508 (N_37508,N_23623,N_22544);
xor U37509 (N_37509,N_28060,N_25679);
and U37510 (N_37510,N_22774,N_23550);
and U37511 (N_37511,N_23205,N_26756);
nor U37512 (N_37512,N_21218,N_25833);
nand U37513 (N_37513,N_29273,N_29697);
and U37514 (N_37514,N_20676,N_27729);
nor U37515 (N_37515,N_22311,N_28033);
nor U37516 (N_37516,N_25626,N_27661);
and U37517 (N_37517,N_25864,N_23788);
xnor U37518 (N_37518,N_23905,N_24725);
nand U37519 (N_37519,N_24952,N_22402);
nor U37520 (N_37520,N_26875,N_20723);
or U37521 (N_37521,N_28193,N_24796);
nor U37522 (N_37522,N_23908,N_28685);
nor U37523 (N_37523,N_21476,N_26745);
or U37524 (N_37524,N_24669,N_25035);
or U37525 (N_37525,N_20014,N_22916);
and U37526 (N_37526,N_21497,N_26003);
or U37527 (N_37527,N_29874,N_23001);
and U37528 (N_37528,N_25165,N_28762);
nand U37529 (N_37529,N_29171,N_27171);
or U37530 (N_37530,N_26329,N_24635);
nor U37531 (N_37531,N_22181,N_29253);
and U37532 (N_37532,N_24882,N_25499);
nand U37533 (N_37533,N_28315,N_20094);
and U37534 (N_37534,N_23732,N_23628);
nor U37535 (N_37535,N_21877,N_23201);
nor U37536 (N_37536,N_26151,N_25976);
and U37537 (N_37537,N_24584,N_21631);
and U37538 (N_37538,N_22868,N_22530);
nor U37539 (N_37539,N_22657,N_28300);
or U37540 (N_37540,N_20964,N_20715);
xor U37541 (N_37541,N_29457,N_29399);
nand U37542 (N_37542,N_29256,N_28012);
and U37543 (N_37543,N_26443,N_24834);
and U37544 (N_37544,N_26226,N_24921);
nor U37545 (N_37545,N_25412,N_25772);
or U37546 (N_37546,N_23121,N_20177);
or U37547 (N_37547,N_20147,N_23868);
and U37548 (N_37548,N_25342,N_24308);
and U37549 (N_37549,N_28707,N_21492);
nor U37550 (N_37550,N_22815,N_21438);
nor U37551 (N_37551,N_23517,N_25760);
or U37552 (N_37552,N_25310,N_21295);
nand U37553 (N_37553,N_20658,N_27534);
xnor U37554 (N_37554,N_23507,N_28316);
and U37555 (N_37555,N_29399,N_29039);
nand U37556 (N_37556,N_26583,N_26776);
nor U37557 (N_37557,N_22766,N_23394);
nand U37558 (N_37558,N_20957,N_28677);
or U37559 (N_37559,N_28182,N_27606);
or U37560 (N_37560,N_28188,N_20960);
xor U37561 (N_37561,N_26384,N_27580);
and U37562 (N_37562,N_29342,N_29005);
nor U37563 (N_37563,N_29744,N_27911);
or U37564 (N_37564,N_22587,N_21006);
or U37565 (N_37565,N_23622,N_23022);
and U37566 (N_37566,N_26177,N_23366);
nand U37567 (N_37567,N_24070,N_24733);
and U37568 (N_37568,N_27027,N_21287);
xnor U37569 (N_37569,N_27552,N_22419);
or U37570 (N_37570,N_25079,N_22454);
or U37571 (N_37571,N_28191,N_27822);
nand U37572 (N_37572,N_20378,N_23285);
nand U37573 (N_37573,N_20776,N_27773);
nor U37574 (N_37574,N_22588,N_25424);
or U37575 (N_37575,N_29842,N_27438);
nand U37576 (N_37576,N_24487,N_28744);
or U37577 (N_37577,N_21677,N_23925);
and U37578 (N_37578,N_24806,N_28470);
nor U37579 (N_37579,N_22152,N_28845);
and U37580 (N_37580,N_20598,N_24631);
nor U37581 (N_37581,N_23176,N_26291);
or U37582 (N_37582,N_22964,N_20407);
nor U37583 (N_37583,N_21484,N_27559);
or U37584 (N_37584,N_20223,N_27872);
or U37585 (N_37585,N_24294,N_28656);
nand U37586 (N_37586,N_22992,N_23608);
and U37587 (N_37587,N_29055,N_29217);
nand U37588 (N_37588,N_28422,N_24977);
nor U37589 (N_37589,N_25653,N_25263);
nor U37590 (N_37590,N_20418,N_24489);
nand U37591 (N_37591,N_27886,N_26199);
nand U37592 (N_37592,N_28074,N_28081);
nand U37593 (N_37593,N_23426,N_20293);
nor U37594 (N_37594,N_24116,N_27637);
or U37595 (N_37595,N_20492,N_20969);
nor U37596 (N_37596,N_24837,N_21613);
or U37597 (N_37597,N_24995,N_20331);
and U37598 (N_37598,N_29633,N_26516);
nor U37599 (N_37599,N_20693,N_25736);
or U37600 (N_37600,N_29154,N_25865);
or U37601 (N_37601,N_23979,N_22672);
and U37602 (N_37602,N_24899,N_22205);
and U37603 (N_37603,N_24860,N_28665);
and U37604 (N_37604,N_23178,N_27924);
and U37605 (N_37605,N_22230,N_26492);
or U37606 (N_37606,N_21590,N_28272);
and U37607 (N_37607,N_29720,N_25001);
nor U37608 (N_37608,N_20146,N_25261);
nand U37609 (N_37609,N_22637,N_25597);
and U37610 (N_37610,N_20331,N_25878);
or U37611 (N_37611,N_22251,N_28095);
xnor U37612 (N_37612,N_23849,N_26347);
and U37613 (N_37613,N_25518,N_29194);
nor U37614 (N_37614,N_25259,N_26266);
xnor U37615 (N_37615,N_28900,N_28945);
or U37616 (N_37616,N_28220,N_27111);
nand U37617 (N_37617,N_21340,N_20648);
and U37618 (N_37618,N_25816,N_28396);
or U37619 (N_37619,N_21075,N_24899);
nand U37620 (N_37620,N_21490,N_26194);
or U37621 (N_37621,N_24167,N_25543);
nor U37622 (N_37622,N_24327,N_28944);
nand U37623 (N_37623,N_20142,N_24736);
nor U37624 (N_37624,N_27451,N_20729);
or U37625 (N_37625,N_22185,N_21507);
nand U37626 (N_37626,N_29886,N_23540);
xnor U37627 (N_37627,N_25330,N_24889);
nand U37628 (N_37628,N_21931,N_20246);
nand U37629 (N_37629,N_22079,N_20647);
and U37630 (N_37630,N_20683,N_20831);
nor U37631 (N_37631,N_25835,N_28778);
or U37632 (N_37632,N_22872,N_22552);
nand U37633 (N_37633,N_22537,N_27935);
and U37634 (N_37634,N_24323,N_27049);
or U37635 (N_37635,N_20051,N_21912);
xnor U37636 (N_37636,N_28685,N_23373);
nor U37637 (N_37637,N_20687,N_23908);
and U37638 (N_37638,N_28993,N_21003);
nor U37639 (N_37639,N_21748,N_21036);
nand U37640 (N_37640,N_24348,N_29427);
or U37641 (N_37641,N_28271,N_28809);
nand U37642 (N_37642,N_22954,N_26365);
and U37643 (N_37643,N_27730,N_27678);
or U37644 (N_37644,N_20052,N_24119);
nor U37645 (N_37645,N_21818,N_25214);
or U37646 (N_37646,N_21840,N_26942);
or U37647 (N_37647,N_24096,N_27475);
xor U37648 (N_37648,N_27969,N_23839);
nand U37649 (N_37649,N_26954,N_21597);
and U37650 (N_37650,N_23164,N_25537);
or U37651 (N_37651,N_29821,N_22344);
nor U37652 (N_37652,N_20768,N_21325);
nor U37653 (N_37653,N_23284,N_21602);
nand U37654 (N_37654,N_28370,N_23510);
nor U37655 (N_37655,N_21742,N_26267);
and U37656 (N_37656,N_25376,N_28125);
nand U37657 (N_37657,N_20292,N_20785);
or U37658 (N_37658,N_23940,N_23796);
nand U37659 (N_37659,N_21187,N_27413);
nand U37660 (N_37660,N_26131,N_25562);
and U37661 (N_37661,N_22435,N_27859);
and U37662 (N_37662,N_21272,N_26819);
or U37663 (N_37663,N_25673,N_21886);
or U37664 (N_37664,N_20247,N_25758);
or U37665 (N_37665,N_27180,N_22563);
nand U37666 (N_37666,N_22481,N_26924);
nand U37667 (N_37667,N_28919,N_25381);
nor U37668 (N_37668,N_27327,N_25266);
nor U37669 (N_37669,N_27447,N_28525);
and U37670 (N_37670,N_29202,N_24589);
and U37671 (N_37671,N_24325,N_24154);
and U37672 (N_37672,N_26872,N_20145);
and U37673 (N_37673,N_28765,N_28219);
and U37674 (N_37674,N_27523,N_25022);
and U37675 (N_37675,N_23952,N_20043);
or U37676 (N_37676,N_22704,N_28263);
or U37677 (N_37677,N_23695,N_22526);
and U37678 (N_37678,N_24728,N_26475);
nand U37679 (N_37679,N_23880,N_24385);
xnor U37680 (N_37680,N_29999,N_27823);
and U37681 (N_37681,N_24276,N_21311);
or U37682 (N_37682,N_28679,N_27489);
and U37683 (N_37683,N_27188,N_24769);
nor U37684 (N_37684,N_28103,N_29093);
and U37685 (N_37685,N_28593,N_20324);
or U37686 (N_37686,N_26418,N_20289);
or U37687 (N_37687,N_24809,N_21709);
nand U37688 (N_37688,N_24427,N_23042);
and U37689 (N_37689,N_23476,N_28885);
nor U37690 (N_37690,N_29212,N_22885);
or U37691 (N_37691,N_29451,N_24316);
or U37692 (N_37692,N_28816,N_26823);
and U37693 (N_37693,N_24772,N_23880);
nor U37694 (N_37694,N_24277,N_26422);
and U37695 (N_37695,N_20579,N_29855);
nand U37696 (N_37696,N_20658,N_20593);
nor U37697 (N_37697,N_22072,N_28266);
nor U37698 (N_37698,N_29352,N_22700);
or U37699 (N_37699,N_24311,N_26317);
and U37700 (N_37700,N_28081,N_26112);
or U37701 (N_37701,N_22704,N_23427);
nand U37702 (N_37702,N_24434,N_24282);
or U37703 (N_37703,N_25269,N_22590);
and U37704 (N_37704,N_20635,N_24153);
nor U37705 (N_37705,N_22041,N_26818);
nor U37706 (N_37706,N_22038,N_23659);
or U37707 (N_37707,N_22758,N_26555);
or U37708 (N_37708,N_27455,N_24798);
xnor U37709 (N_37709,N_26576,N_20479);
and U37710 (N_37710,N_20277,N_25541);
nor U37711 (N_37711,N_27733,N_25728);
and U37712 (N_37712,N_26880,N_20330);
nor U37713 (N_37713,N_23073,N_24456);
xnor U37714 (N_37714,N_21423,N_20719);
or U37715 (N_37715,N_24024,N_25129);
or U37716 (N_37716,N_23675,N_23619);
and U37717 (N_37717,N_26966,N_26324);
or U37718 (N_37718,N_20032,N_28561);
or U37719 (N_37719,N_27140,N_24665);
nand U37720 (N_37720,N_24947,N_27858);
or U37721 (N_37721,N_24091,N_27969);
or U37722 (N_37722,N_23942,N_24161);
nand U37723 (N_37723,N_23850,N_22295);
nor U37724 (N_37724,N_25550,N_23415);
and U37725 (N_37725,N_28543,N_24070);
or U37726 (N_37726,N_25868,N_24342);
or U37727 (N_37727,N_27177,N_29535);
or U37728 (N_37728,N_26884,N_21577);
nand U37729 (N_37729,N_24756,N_24688);
or U37730 (N_37730,N_22613,N_24155);
xor U37731 (N_37731,N_23393,N_21442);
nand U37732 (N_37732,N_25976,N_28859);
nor U37733 (N_37733,N_22692,N_26392);
nor U37734 (N_37734,N_24410,N_23844);
and U37735 (N_37735,N_26957,N_22179);
and U37736 (N_37736,N_29071,N_29184);
xnor U37737 (N_37737,N_20089,N_23952);
nand U37738 (N_37738,N_20342,N_29936);
nor U37739 (N_37739,N_21818,N_20598);
and U37740 (N_37740,N_27025,N_28311);
or U37741 (N_37741,N_22494,N_24655);
nand U37742 (N_37742,N_22579,N_28281);
xor U37743 (N_37743,N_21844,N_28901);
xnor U37744 (N_37744,N_24822,N_27151);
xnor U37745 (N_37745,N_25117,N_22753);
nand U37746 (N_37746,N_23243,N_27136);
xnor U37747 (N_37747,N_29690,N_20258);
nor U37748 (N_37748,N_26129,N_29861);
nor U37749 (N_37749,N_29248,N_26095);
nand U37750 (N_37750,N_26987,N_29716);
and U37751 (N_37751,N_20278,N_24000);
or U37752 (N_37752,N_29072,N_28563);
nand U37753 (N_37753,N_29601,N_21068);
or U37754 (N_37754,N_28990,N_28084);
or U37755 (N_37755,N_27205,N_22682);
xnor U37756 (N_37756,N_26398,N_28816);
xnor U37757 (N_37757,N_26935,N_20650);
or U37758 (N_37758,N_20810,N_28734);
or U37759 (N_37759,N_21510,N_22173);
nand U37760 (N_37760,N_27145,N_21955);
nand U37761 (N_37761,N_26582,N_29629);
nor U37762 (N_37762,N_20860,N_25953);
and U37763 (N_37763,N_25341,N_21185);
or U37764 (N_37764,N_27368,N_23730);
or U37765 (N_37765,N_28314,N_21073);
nand U37766 (N_37766,N_25083,N_23209);
nand U37767 (N_37767,N_22708,N_27630);
xor U37768 (N_37768,N_20814,N_22510);
or U37769 (N_37769,N_28341,N_27954);
nand U37770 (N_37770,N_28964,N_27581);
and U37771 (N_37771,N_26827,N_23739);
or U37772 (N_37772,N_28438,N_26064);
nor U37773 (N_37773,N_24723,N_29968);
and U37774 (N_37774,N_24785,N_20729);
xor U37775 (N_37775,N_22172,N_21245);
nor U37776 (N_37776,N_26062,N_25383);
nand U37777 (N_37777,N_29243,N_24122);
or U37778 (N_37778,N_20973,N_26026);
or U37779 (N_37779,N_20401,N_23712);
or U37780 (N_37780,N_26081,N_23897);
nor U37781 (N_37781,N_25661,N_28386);
and U37782 (N_37782,N_23850,N_21476);
and U37783 (N_37783,N_20382,N_26188);
and U37784 (N_37784,N_21554,N_26039);
or U37785 (N_37785,N_29711,N_20179);
xnor U37786 (N_37786,N_22029,N_21340);
and U37787 (N_37787,N_21215,N_22459);
xor U37788 (N_37788,N_21433,N_28963);
nor U37789 (N_37789,N_20639,N_23131);
nor U37790 (N_37790,N_26086,N_24466);
and U37791 (N_37791,N_21821,N_21783);
nand U37792 (N_37792,N_24119,N_26445);
nor U37793 (N_37793,N_27486,N_25440);
and U37794 (N_37794,N_28995,N_27041);
nand U37795 (N_37795,N_28551,N_26362);
and U37796 (N_37796,N_24058,N_26676);
nand U37797 (N_37797,N_25720,N_24755);
nand U37798 (N_37798,N_21321,N_25791);
nand U37799 (N_37799,N_28572,N_27680);
nand U37800 (N_37800,N_23111,N_22300);
xnor U37801 (N_37801,N_26290,N_20501);
nand U37802 (N_37802,N_21648,N_22763);
nand U37803 (N_37803,N_23713,N_21556);
and U37804 (N_37804,N_21641,N_24199);
or U37805 (N_37805,N_21607,N_22045);
nor U37806 (N_37806,N_24416,N_20446);
and U37807 (N_37807,N_25089,N_20335);
or U37808 (N_37808,N_28996,N_21633);
or U37809 (N_37809,N_29597,N_26192);
nor U37810 (N_37810,N_27829,N_27505);
nor U37811 (N_37811,N_29890,N_23568);
nand U37812 (N_37812,N_22953,N_28745);
or U37813 (N_37813,N_26121,N_23441);
and U37814 (N_37814,N_20607,N_25662);
and U37815 (N_37815,N_28256,N_24958);
and U37816 (N_37816,N_28859,N_21262);
or U37817 (N_37817,N_24024,N_22138);
xor U37818 (N_37818,N_22103,N_21677);
or U37819 (N_37819,N_21105,N_28779);
nor U37820 (N_37820,N_26943,N_25952);
nor U37821 (N_37821,N_27210,N_25433);
and U37822 (N_37822,N_27987,N_21388);
nand U37823 (N_37823,N_27711,N_27737);
xnor U37824 (N_37824,N_20976,N_23641);
nor U37825 (N_37825,N_24361,N_26379);
xor U37826 (N_37826,N_27559,N_26628);
nand U37827 (N_37827,N_27738,N_21841);
nor U37828 (N_37828,N_28012,N_23114);
and U37829 (N_37829,N_27123,N_20072);
and U37830 (N_37830,N_25098,N_27139);
nor U37831 (N_37831,N_21061,N_21682);
nor U37832 (N_37832,N_28501,N_21629);
or U37833 (N_37833,N_20806,N_20326);
or U37834 (N_37834,N_26268,N_27534);
or U37835 (N_37835,N_25113,N_25599);
nor U37836 (N_37836,N_27572,N_26817);
and U37837 (N_37837,N_20938,N_23894);
and U37838 (N_37838,N_20044,N_29757);
xor U37839 (N_37839,N_24000,N_22490);
xor U37840 (N_37840,N_21101,N_27284);
nand U37841 (N_37841,N_28557,N_20605);
nor U37842 (N_37842,N_22642,N_20241);
and U37843 (N_37843,N_26499,N_26134);
xor U37844 (N_37844,N_28609,N_25144);
and U37845 (N_37845,N_24075,N_21451);
or U37846 (N_37846,N_24075,N_24526);
and U37847 (N_37847,N_27062,N_21369);
xor U37848 (N_37848,N_22180,N_23581);
or U37849 (N_37849,N_22988,N_20600);
nand U37850 (N_37850,N_26598,N_26018);
nor U37851 (N_37851,N_21561,N_23276);
nor U37852 (N_37852,N_28431,N_29512);
and U37853 (N_37853,N_27634,N_28725);
nand U37854 (N_37854,N_24721,N_26975);
and U37855 (N_37855,N_27002,N_20763);
nand U37856 (N_37856,N_25529,N_22859);
and U37857 (N_37857,N_20378,N_20757);
and U37858 (N_37858,N_21074,N_29099);
and U37859 (N_37859,N_23015,N_28593);
nor U37860 (N_37860,N_23939,N_20438);
and U37861 (N_37861,N_22155,N_24466);
nor U37862 (N_37862,N_21172,N_24869);
xnor U37863 (N_37863,N_25877,N_23436);
or U37864 (N_37864,N_23256,N_28678);
nand U37865 (N_37865,N_25981,N_24629);
nor U37866 (N_37866,N_22308,N_23452);
nor U37867 (N_37867,N_20878,N_22010);
nand U37868 (N_37868,N_26369,N_28534);
or U37869 (N_37869,N_23351,N_24148);
and U37870 (N_37870,N_22999,N_28859);
and U37871 (N_37871,N_21540,N_27164);
or U37872 (N_37872,N_21838,N_21872);
nand U37873 (N_37873,N_28613,N_21686);
nand U37874 (N_37874,N_28735,N_21644);
nor U37875 (N_37875,N_29809,N_21467);
and U37876 (N_37876,N_20588,N_26549);
xnor U37877 (N_37877,N_24773,N_29570);
or U37878 (N_37878,N_24253,N_22597);
nand U37879 (N_37879,N_24302,N_29786);
nor U37880 (N_37880,N_28159,N_29665);
xnor U37881 (N_37881,N_20029,N_27121);
or U37882 (N_37882,N_26817,N_26984);
nor U37883 (N_37883,N_21200,N_22329);
nor U37884 (N_37884,N_22208,N_23327);
and U37885 (N_37885,N_25924,N_29254);
nand U37886 (N_37886,N_20798,N_27987);
or U37887 (N_37887,N_26917,N_21539);
nand U37888 (N_37888,N_28249,N_26234);
nor U37889 (N_37889,N_28466,N_21561);
nand U37890 (N_37890,N_23130,N_27570);
or U37891 (N_37891,N_23990,N_29824);
or U37892 (N_37892,N_22544,N_28206);
or U37893 (N_37893,N_29631,N_29401);
nor U37894 (N_37894,N_25894,N_29164);
or U37895 (N_37895,N_23482,N_20677);
or U37896 (N_37896,N_28897,N_26519);
or U37897 (N_37897,N_23071,N_23601);
xnor U37898 (N_37898,N_26601,N_27625);
nand U37899 (N_37899,N_20369,N_23122);
xor U37900 (N_37900,N_25239,N_20181);
nor U37901 (N_37901,N_27110,N_22669);
and U37902 (N_37902,N_22323,N_23191);
xor U37903 (N_37903,N_26398,N_25524);
nor U37904 (N_37904,N_21424,N_26169);
or U37905 (N_37905,N_25637,N_27492);
nor U37906 (N_37906,N_20529,N_22060);
xor U37907 (N_37907,N_21562,N_22718);
nand U37908 (N_37908,N_26027,N_22196);
and U37909 (N_37909,N_25914,N_23552);
nand U37910 (N_37910,N_29411,N_29040);
xnor U37911 (N_37911,N_24978,N_26973);
or U37912 (N_37912,N_21791,N_29686);
nor U37913 (N_37913,N_28604,N_20613);
nor U37914 (N_37914,N_20225,N_29792);
nand U37915 (N_37915,N_29828,N_25202);
xnor U37916 (N_37916,N_23811,N_23852);
nor U37917 (N_37917,N_23892,N_26135);
nor U37918 (N_37918,N_20775,N_22830);
nand U37919 (N_37919,N_23077,N_20166);
nor U37920 (N_37920,N_21208,N_28360);
nand U37921 (N_37921,N_27468,N_22623);
nor U37922 (N_37922,N_27077,N_27997);
nand U37923 (N_37923,N_25322,N_26124);
nand U37924 (N_37924,N_29727,N_26099);
nor U37925 (N_37925,N_26561,N_20093);
or U37926 (N_37926,N_26300,N_26089);
nor U37927 (N_37927,N_22113,N_20814);
and U37928 (N_37928,N_22416,N_22474);
or U37929 (N_37929,N_28127,N_20235);
or U37930 (N_37930,N_24118,N_28737);
or U37931 (N_37931,N_26248,N_28532);
and U37932 (N_37932,N_29276,N_20452);
nand U37933 (N_37933,N_20103,N_26966);
and U37934 (N_37934,N_28011,N_25960);
or U37935 (N_37935,N_21433,N_20731);
and U37936 (N_37936,N_29624,N_29805);
xor U37937 (N_37937,N_27376,N_22621);
and U37938 (N_37938,N_22047,N_25572);
and U37939 (N_37939,N_29036,N_22402);
nor U37940 (N_37940,N_27184,N_20084);
or U37941 (N_37941,N_22021,N_26824);
or U37942 (N_37942,N_24838,N_24665);
or U37943 (N_37943,N_27779,N_22638);
or U37944 (N_37944,N_24968,N_20383);
or U37945 (N_37945,N_27602,N_23559);
and U37946 (N_37946,N_24073,N_29404);
nor U37947 (N_37947,N_28596,N_21618);
nand U37948 (N_37948,N_24530,N_25143);
nor U37949 (N_37949,N_20028,N_20216);
nor U37950 (N_37950,N_22251,N_25034);
nor U37951 (N_37951,N_28278,N_28363);
or U37952 (N_37952,N_28700,N_29193);
nor U37953 (N_37953,N_29556,N_21367);
or U37954 (N_37954,N_23545,N_22489);
and U37955 (N_37955,N_26653,N_22554);
xnor U37956 (N_37956,N_26080,N_23664);
nand U37957 (N_37957,N_21507,N_26150);
nand U37958 (N_37958,N_21999,N_22674);
xor U37959 (N_37959,N_20208,N_25674);
or U37960 (N_37960,N_28126,N_28647);
and U37961 (N_37961,N_22975,N_27618);
nand U37962 (N_37962,N_29473,N_20940);
nand U37963 (N_37963,N_28329,N_29756);
nor U37964 (N_37964,N_22266,N_21178);
nor U37965 (N_37965,N_21247,N_24909);
xnor U37966 (N_37966,N_26791,N_22918);
or U37967 (N_37967,N_22684,N_24768);
xor U37968 (N_37968,N_24544,N_20240);
nor U37969 (N_37969,N_29863,N_22177);
nor U37970 (N_37970,N_27098,N_21072);
or U37971 (N_37971,N_29583,N_24897);
nor U37972 (N_37972,N_21223,N_24170);
and U37973 (N_37973,N_27909,N_22042);
or U37974 (N_37974,N_22871,N_25624);
nor U37975 (N_37975,N_26658,N_27291);
or U37976 (N_37976,N_24529,N_25288);
and U37977 (N_37977,N_22921,N_28960);
and U37978 (N_37978,N_27952,N_21700);
nor U37979 (N_37979,N_25502,N_27192);
or U37980 (N_37980,N_26231,N_24639);
and U37981 (N_37981,N_29079,N_28335);
or U37982 (N_37982,N_25898,N_28918);
or U37983 (N_37983,N_22475,N_22464);
xnor U37984 (N_37984,N_26823,N_23289);
nor U37985 (N_37985,N_20570,N_21653);
and U37986 (N_37986,N_28034,N_28133);
and U37987 (N_37987,N_28086,N_27236);
and U37988 (N_37988,N_24897,N_21940);
xnor U37989 (N_37989,N_29143,N_22075);
nor U37990 (N_37990,N_25882,N_20348);
xor U37991 (N_37991,N_26888,N_22297);
and U37992 (N_37992,N_27080,N_20039);
nor U37993 (N_37993,N_27145,N_24587);
nand U37994 (N_37994,N_25698,N_24689);
nor U37995 (N_37995,N_24969,N_21617);
nand U37996 (N_37996,N_21803,N_20945);
nor U37997 (N_37997,N_26129,N_22863);
xor U37998 (N_37998,N_27848,N_23664);
xor U37999 (N_37999,N_23739,N_25715);
nor U38000 (N_38000,N_25928,N_25654);
nor U38001 (N_38001,N_21322,N_23591);
xor U38002 (N_38002,N_20640,N_21346);
nor U38003 (N_38003,N_24377,N_21488);
nor U38004 (N_38004,N_27655,N_28835);
or U38005 (N_38005,N_24940,N_25184);
and U38006 (N_38006,N_24314,N_27011);
or U38007 (N_38007,N_26641,N_26116);
nand U38008 (N_38008,N_21728,N_28636);
nor U38009 (N_38009,N_29485,N_29869);
and U38010 (N_38010,N_29758,N_21393);
and U38011 (N_38011,N_27257,N_26091);
or U38012 (N_38012,N_21938,N_20466);
or U38013 (N_38013,N_20224,N_26395);
or U38014 (N_38014,N_21672,N_21567);
xor U38015 (N_38015,N_20032,N_29650);
nor U38016 (N_38016,N_20452,N_21716);
and U38017 (N_38017,N_28937,N_26987);
nand U38018 (N_38018,N_23998,N_26769);
and U38019 (N_38019,N_20749,N_21731);
nand U38020 (N_38020,N_24695,N_28036);
nand U38021 (N_38021,N_28773,N_21568);
nor U38022 (N_38022,N_29289,N_29798);
nor U38023 (N_38023,N_25925,N_26356);
nand U38024 (N_38024,N_26870,N_26088);
nor U38025 (N_38025,N_26670,N_28110);
nor U38026 (N_38026,N_24858,N_25603);
xnor U38027 (N_38027,N_24330,N_25317);
nand U38028 (N_38028,N_21740,N_25804);
and U38029 (N_38029,N_22522,N_29352);
nand U38030 (N_38030,N_26308,N_20223);
and U38031 (N_38031,N_21473,N_21896);
and U38032 (N_38032,N_20855,N_28475);
or U38033 (N_38033,N_20603,N_28282);
nand U38034 (N_38034,N_27291,N_20871);
nor U38035 (N_38035,N_24431,N_29425);
or U38036 (N_38036,N_25999,N_27712);
nand U38037 (N_38037,N_26678,N_27417);
nor U38038 (N_38038,N_24973,N_26362);
nor U38039 (N_38039,N_27572,N_29026);
and U38040 (N_38040,N_28752,N_22175);
and U38041 (N_38041,N_20505,N_28195);
and U38042 (N_38042,N_29413,N_27237);
or U38043 (N_38043,N_22748,N_24873);
nor U38044 (N_38044,N_21567,N_22231);
or U38045 (N_38045,N_27797,N_22393);
nand U38046 (N_38046,N_29525,N_27979);
xor U38047 (N_38047,N_23204,N_26729);
or U38048 (N_38048,N_21661,N_27108);
nor U38049 (N_38049,N_22342,N_23422);
nor U38050 (N_38050,N_21354,N_28401);
nor U38051 (N_38051,N_24825,N_25731);
xor U38052 (N_38052,N_23408,N_21579);
nor U38053 (N_38053,N_26920,N_26107);
and U38054 (N_38054,N_24508,N_24125);
nor U38055 (N_38055,N_21950,N_29938);
nor U38056 (N_38056,N_26997,N_24809);
or U38057 (N_38057,N_21890,N_26412);
and U38058 (N_38058,N_20380,N_26708);
xor U38059 (N_38059,N_28883,N_21094);
nand U38060 (N_38060,N_26546,N_29419);
nand U38061 (N_38061,N_26259,N_29725);
and U38062 (N_38062,N_25391,N_26767);
and U38063 (N_38063,N_20095,N_21909);
xnor U38064 (N_38064,N_26712,N_20000);
nand U38065 (N_38065,N_29268,N_20488);
xnor U38066 (N_38066,N_25639,N_26613);
and U38067 (N_38067,N_24218,N_28481);
or U38068 (N_38068,N_21192,N_20785);
nand U38069 (N_38069,N_24089,N_23957);
or U38070 (N_38070,N_22838,N_29522);
or U38071 (N_38071,N_27186,N_22964);
or U38072 (N_38072,N_24611,N_23325);
nor U38073 (N_38073,N_24209,N_26388);
nor U38074 (N_38074,N_26433,N_28449);
nor U38075 (N_38075,N_22569,N_26037);
nand U38076 (N_38076,N_21820,N_22147);
xor U38077 (N_38077,N_28566,N_28817);
nand U38078 (N_38078,N_23226,N_21486);
or U38079 (N_38079,N_28716,N_24664);
and U38080 (N_38080,N_28055,N_25591);
and U38081 (N_38081,N_20486,N_20889);
nand U38082 (N_38082,N_29546,N_24737);
and U38083 (N_38083,N_26963,N_20633);
and U38084 (N_38084,N_20308,N_22598);
xor U38085 (N_38085,N_20335,N_22646);
and U38086 (N_38086,N_21483,N_26240);
xnor U38087 (N_38087,N_27764,N_26227);
xnor U38088 (N_38088,N_24576,N_21094);
or U38089 (N_38089,N_27764,N_22325);
or U38090 (N_38090,N_26013,N_28758);
nor U38091 (N_38091,N_25099,N_22032);
or U38092 (N_38092,N_22312,N_21895);
xnor U38093 (N_38093,N_28958,N_26234);
nor U38094 (N_38094,N_29407,N_20591);
nand U38095 (N_38095,N_23733,N_21491);
and U38096 (N_38096,N_29221,N_26319);
nor U38097 (N_38097,N_20559,N_28870);
or U38098 (N_38098,N_25580,N_29349);
xnor U38099 (N_38099,N_29843,N_25924);
nor U38100 (N_38100,N_29315,N_24346);
nand U38101 (N_38101,N_24632,N_24309);
xnor U38102 (N_38102,N_24884,N_20877);
or U38103 (N_38103,N_20799,N_24551);
nand U38104 (N_38104,N_24222,N_22229);
nand U38105 (N_38105,N_25664,N_28396);
or U38106 (N_38106,N_25251,N_27946);
nand U38107 (N_38107,N_28195,N_24811);
nor U38108 (N_38108,N_26188,N_20502);
and U38109 (N_38109,N_27333,N_22641);
nor U38110 (N_38110,N_25350,N_26129);
or U38111 (N_38111,N_21214,N_24165);
and U38112 (N_38112,N_26364,N_22199);
xor U38113 (N_38113,N_20568,N_20710);
or U38114 (N_38114,N_27980,N_20648);
nand U38115 (N_38115,N_23710,N_20180);
xor U38116 (N_38116,N_26687,N_20445);
or U38117 (N_38117,N_26475,N_22826);
nor U38118 (N_38118,N_25067,N_22739);
nor U38119 (N_38119,N_28240,N_25013);
or U38120 (N_38120,N_28401,N_21220);
nand U38121 (N_38121,N_26131,N_23311);
and U38122 (N_38122,N_25060,N_22701);
or U38123 (N_38123,N_28313,N_26233);
nor U38124 (N_38124,N_27096,N_22640);
and U38125 (N_38125,N_26628,N_24063);
nand U38126 (N_38126,N_24919,N_22590);
xor U38127 (N_38127,N_20196,N_25290);
xnor U38128 (N_38128,N_20539,N_20999);
and U38129 (N_38129,N_22587,N_22542);
nor U38130 (N_38130,N_24469,N_25024);
or U38131 (N_38131,N_27097,N_24191);
nor U38132 (N_38132,N_25278,N_26453);
or U38133 (N_38133,N_26658,N_27608);
xor U38134 (N_38134,N_24378,N_29582);
and U38135 (N_38135,N_28502,N_25128);
nand U38136 (N_38136,N_20472,N_25718);
nand U38137 (N_38137,N_21249,N_28101);
and U38138 (N_38138,N_29224,N_29868);
nor U38139 (N_38139,N_29777,N_23396);
and U38140 (N_38140,N_20744,N_24894);
xnor U38141 (N_38141,N_25417,N_28720);
nor U38142 (N_38142,N_23709,N_22286);
or U38143 (N_38143,N_22895,N_29258);
xnor U38144 (N_38144,N_25364,N_27669);
and U38145 (N_38145,N_20246,N_24681);
nand U38146 (N_38146,N_24015,N_25153);
nand U38147 (N_38147,N_23606,N_20873);
and U38148 (N_38148,N_24349,N_28107);
or U38149 (N_38149,N_20357,N_23921);
nand U38150 (N_38150,N_29600,N_26448);
xor U38151 (N_38151,N_23499,N_23254);
and U38152 (N_38152,N_29504,N_29302);
xor U38153 (N_38153,N_23200,N_24231);
nand U38154 (N_38154,N_28858,N_27306);
nor U38155 (N_38155,N_26850,N_24200);
nor U38156 (N_38156,N_21235,N_23239);
nand U38157 (N_38157,N_20546,N_27609);
nand U38158 (N_38158,N_26627,N_23805);
nand U38159 (N_38159,N_25070,N_20152);
and U38160 (N_38160,N_27490,N_27007);
nand U38161 (N_38161,N_24990,N_23370);
xnor U38162 (N_38162,N_26593,N_28406);
xor U38163 (N_38163,N_24798,N_27341);
xnor U38164 (N_38164,N_20969,N_23924);
nand U38165 (N_38165,N_26184,N_29570);
and U38166 (N_38166,N_26138,N_28406);
or U38167 (N_38167,N_25373,N_24304);
nor U38168 (N_38168,N_22963,N_23100);
and U38169 (N_38169,N_20082,N_26318);
nand U38170 (N_38170,N_23559,N_27376);
or U38171 (N_38171,N_26591,N_26976);
and U38172 (N_38172,N_25814,N_24713);
and U38173 (N_38173,N_20355,N_23609);
and U38174 (N_38174,N_29814,N_23940);
nand U38175 (N_38175,N_23698,N_27762);
nand U38176 (N_38176,N_20790,N_21002);
nor U38177 (N_38177,N_27522,N_25489);
nor U38178 (N_38178,N_24749,N_23628);
nand U38179 (N_38179,N_27274,N_21801);
xor U38180 (N_38180,N_29657,N_22885);
and U38181 (N_38181,N_28116,N_22700);
nor U38182 (N_38182,N_20841,N_22422);
nor U38183 (N_38183,N_20793,N_28849);
and U38184 (N_38184,N_21690,N_22223);
or U38185 (N_38185,N_21979,N_28916);
or U38186 (N_38186,N_28934,N_20457);
nor U38187 (N_38187,N_21154,N_27300);
or U38188 (N_38188,N_20379,N_28599);
or U38189 (N_38189,N_24595,N_28521);
and U38190 (N_38190,N_24056,N_20661);
nand U38191 (N_38191,N_25914,N_29816);
or U38192 (N_38192,N_20023,N_27424);
or U38193 (N_38193,N_27146,N_27490);
nand U38194 (N_38194,N_23695,N_24130);
or U38195 (N_38195,N_29121,N_24102);
nand U38196 (N_38196,N_26813,N_29824);
and U38197 (N_38197,N_23528,N_20966);
nand U38198 (N_38198,N_29482,N_24057);
or U38199 (N_38199,N_27681,N_26448);
nor U38200 (N_38200,N_20449,N_21872);
nor U38201 (N_38201,N_21373,N_26387);
nand U38202 (N_38202,N_21336,N_25342);
nand U38203 (N_38203,N_24463,N_24916);
nor U38204 (N_38204,N_29752,N_21444);
nand U38205 (N_38205,N_29632,N_25299);
nor U38206 (N_38206,N_26452,N_29035);
nand U38207 (N_38207,N_29335,N_26789);
and U38208 (N_38208,N_24750,N_27105);
and U38209 (N_38209,N_23170,N_23503);
and U38210 (N_38210,N_21122,N_25994);
and U38211 (N_38211,N_23416,N_23054);
xor U38212 (N_38212,N_20669,N_26210);
or U38213 (N_38213,N_26993,N_27490);
or U38214 (N_38214,N_28022,N_21571);
or U38215 (N_38215,N_21200,N_29048);
and U38216 (N_38216,N_29073,N_25455);
nand U38217 (N_38217,N_23353,N_22233);
nand U38218 (N_38218,N_25639,N_29377);
nor U38219 (N_38219,N_26415,N_20978);
nor U38220 (N_38220,N_25033,N_23027);
or U38221 (N_38221,N_27538,N_29820);
or U38222 (N_38222,N_25938,N_23438);
and U38223 (N_38223,N_26567,N_27055);
nor U38224 (N_38224,N_26949,N_24731);
xor U38225 (N_38225,N_23142,N_28450);
nand U38226 (N_38226,N_20132,N_27700);
nor U38227 (N_38227,N_27610,N_20305);
nand U38228 (N_38228,N_23342,N_28782);
and U38229 (N_38229,N_25174,N_26543);
and U38230 (N_38230,N_21695,N_28238);
nand U38231 (N_38231,N_28781,N_21167);
nor U38232 (N_38232,N_26176,N_20550);
nor U38233 (N_38233,N_26715,N_20990);
and U38234 (N_38234,N_23715,N_21716);
xnor U38235 (N_38235,N_24010,N_24074);
and U38236 (N_38236,N_25976,N_27711);
or U38237 (N_38237,N_26078,N_25053);
nor U38238 (N_38238,N_25258,N_25056);
nor U38239 (N_38239,N_29116,N_24860);
and U38240 (N_38240,N_28349,N_21474);
or U38241 (N_38241,N_26023,N_22126);
and U38242 (N_38242,N_26127,N_28501);
and U38243 (N_38243,N_23497,N_29893);
nand U38244 (N_38244,N_21548,N_23082);
or U38245 (N_38245,N_26236,N_23008);
nand U38246 (N_38246,N_23742,N_22537);
nor U38247 (N_38247,N_25636,N_25256);
nand U38248 (N_38248,N_25959,N_23966);
nand U38249 (N_38249,N_29096,N_25111);
or U38250 (N_38250,N_28155,N_26740);
and U38251 (N_38251,N_20758,N_28218);
or U38252 (N_38252,N_29530,N_23793);
and U38253 (N_38253,N_27195,N_25566);
xnor U38254 (N_38254,N_20453,N_20456);
or U38255 (N_38255,N_21749,N_28472);
nand U38256 (N_38256,N_23702,N_29547);
xnor U38257 (N_38257,N_23702,N_22787);
nor U38258 (N_38258,N_27573,N_23036);
nand U38259 (N_38259,N_28999,N_28638);
or U38260 (N_38260,N_26416,N_21159);
and U38261 (N_38261,N_23983,N_26413);
or U38262 (N_38262,N_26831,N_29839);
nor U38263 (N_38263,N_24252,N_23144);
xor U38264 (N_38264,N_28287,N_25620);
and U38265 (N_38265,N_25281,N_28862);
xnor U38266 (N_38266,N_25945,N_26078);
and U38267 (N_38267,N_28261,N_24023);
or U38268 (N_38268,N_22524,N_23551);
nor U38269 (N_38269,N_25760,N_27139);
nor U38270 (N_38270,N_29891,N_21426);
or U38271 (N_38271,N_29030,N_27329);
nand U38272 (N_38272,N_26171,N_28852);
nor U38273 (N_38273,N_23587,N_29528);
nand U38274 (N_38274,N_24924,N_22688);
nor U38275 (N_38275,N_24846,N_27273);
and U38276 (N_38276,N_27176,N_28840);
and U38277 (N_38277,N_21572,N_27223);
or U38278 (N_38278,N_28373,N_28182);
nor U38279 (N_38279,N_25455,N_20536);
xor U38280 (N_38280,N_26235,N_20111);
nand U38281 (N_38281,N_28845,N_27572);
or U38282 (N_38282,N_21167,N_22805);
nand U38283 (N_38283,N_27581,N_23246);
or U38284 (N_38284,N_26778,N_27214);
or U38285 (N_38285,N_26886,N_22053);
or U38286 (N_38286,N_28915,N_23157);
and U38287 (N_38287,N_25427,N_29315);
nor U38288 (N_38288,N_23996,N_29984);
nand U38289 (N_38289,N_23456,N_27286);
or U38290 (N_38290,N_26009,N_27329);
or U38291 (N_38291,N_20614,N_23094);
nand U38292 (N_38292,N_27642,N_28706);
nor U38293 (N_38293,N_25571,N_27659);
and U38294 (N_38294,N_22033,N_22116);
and U38295 (N_38295,N_25890,N_24273);
or U38296 (N_38296,N_26410,N_24034);
or U38297 (N_38297,N_28005,N_21759);
or U38298 (N_38298,N_23038,N_25875);
nor U38299 (N_38299,N_27930,N_27583);
or U38300 (N_38300,N_20868,N_21480);
xor U38301 (N_38301,N_27221,N_26983);
and U38302 (N_38302,N_26071,N_23846);
xor U38303 (N_38303,N_26634,N_20132);
nand U38304 (N_38304,N_28985,N_28142);
and U38305 (N_38305,N_28297,N_26079);
nor U38306 (N_38306,N_21451,N_20510);
and U38307 (N_38307,N_21034,N_22645);
or U38308 (N_38308,N_22494,N_29201);
or U38309 (N_38309,N_24636,N_24027);
and U38310 (N_38310,N_24343,N_27914);
or U38311 (N_38311,N_26702,N_24458);
nor U38312 (N_38312,N_29977,N_20262);
or U38313 (N_38313,N_28207,N_27570);
and U38314 (N_38314,N_20518,N_20751);
nand U38315 (N_38315,N_25620,N_27768);
nand U38316 (N_38316,N_20788,N_28754);
or U38317 (N_38317,N_20914,N_25880);
and U38318 (N_38318,N_21219,N_21801);
or U38319 (N_38319,N_29465,N_23957);
xor U38320 (N_38320,N_29450,N_26652);
nor U38321 (N_38321,N_24008,N_22397);
nand U38322 (N_38322,N_20819,N_27078);
nand U38323 (N_38323,N_26500,N_28629);
xor U38324 (N_38324,N_20642,N_26769);
and U38325 (N_38325,N_29902,N_25415);
nand U38326 (N_38326,N_21123,N_29247);
nand U38327 (N_38327,N_29630,N_22433);
or U38328 (N_38328,N_21201,N_22157);
nor U38329 (N_38329,N_20696,N_23828);
nand U38330 (N_38330,N_28291,N_27758);
or U38331 (N_38331,N_22146,N_22613);
and U38332 (N_38332,N_23658,N_28617);
or U38333 (N_38333,N_29706,N_22200);
and U38334 (N_38334,N_29229,N_20371);
nand U38335 (N_38335,N_26731,N_23523);
nand U38336 (N_38336,N_26108,N_20054);
nand U38337 (N_38337,N_24859,N_25756);
xnor U38338 (N_38338,N_28548,N_28980);
or U38339 (N_38339,N_23370,N_27035);
and U38340 (N_38340,N_23139,N_23820);
nand U38341 (N_38341,N_23672,N_28081);
nand U38342 (N_38342,N_27582,N_28238);
and U38343 (N_38343,N_29200,N_23667);
nor U38344 (N_38344,N_29150,N_26205);
and U38345 (N_38345,N_24496,N_27339);
xor U38346 (N_38346,N_27322,N_28370);
nor U38347 (N_38347,N_29598,N_28307);
or U38348 (N_38348,N_21076,N_26144);
nor U38349 (N_38349,N_21757,N_28359);
or U38350 (N_38350,N_26390,N_29434);
and U38351 (N_38351,N_26880,N_29538);
nand U38352 (N_38352,N_22928,N_20173);
nand U38353 (N_38353,N_27600,N_22141);
nand U38354 (N_38354,N_26409,N_24784);
nor U38355 (N_38355,N_23464,N_24574);
and U38356 (N_38356,N_25240,N_20198);
and U38357 (N_38357,N_26275,N_28363);
nor U38358 (N_38358,N_25988,N_21061);
or U38359 (N_38359,N_23543,N_26638);
nand U38360 (N_38360,N_24380,N_21360);
and U38361 (N_38361,N_28050,N_28198);
and U38362 (N_38362,N_23921,N_28442);
nand U38363 (N_38363,N_21937,N_21225);
or U38364 (N_38364,N_28258,N_23255);
nor U38365 (N_38365,N_23413,N_22710);
nand U38366 (N_38366,N_21265,N_25484);
nand U38367 (N_38367,N_23400,N_28116);
nand U38368 (N_38368,N_26976,N_28945);
and U38369 (N_38369,N_21009,N_20784);
nand U38370 (N_38370,N_24088,N_27578);
nand U38371 (N_38371,N_23309,N_20095);
nand U38372 (N_38372,N_23285,N_27271);
xnor U38373 (N_38373,N_23636,N_20729);
xor U38374 (N_38374,N_26186,N_22001);
and U38375 (N_38375,N_26654,N_25684);
nor U38376 (N_38376,N_20943,N_23396);
nor U38377 (N_38377,N_27501,N_21954);
nor U38378 (N_38378,N_29310,N_23326);
xor U38379 (N_38379,N_24757,N_29803);
nor U38380 (N_38380,N_29459,N_22649);
or U38381 (N_38381,N_21478,N_27718);
xor U38382 (N_38382,N_22391,N_27918);
xnor U38383 (N_38383,N_25058,N_21916);
xor U38384 (N_38384,N_26155,N_21419);
nand U38385 (N_38385,N_22554,N_22319);
or U38386 (N_38386,N_20554,N_20826);
xor U38387 (N_38387,N_27914,N_27862);
nor U38388 (N_38388,N_23341,N_20460);
xnor U38389 (N_38389,N_23091,N_22228);
nand U38390 (N_38390,N_20405,N_28478);
and U38391 (N_38391,N_21539,N_27708);
and U38392 (N_38392,N_20411,N_27330);
nand U38393 (N_38393,N_24973,N_22973);
nor U38394 (N_38394,N_28456,N_24391);
nand U38395 (N_38395,N_26380,N_25952);
or U38396 (N_38396,N_28903,N_24107);
and U38397 (N_38397,N_24766,N_25325);
and U38398 (N_38398,N_26289,N_20050);
nor U38399 (N_38399,N_28928,N_25584);
or U38400 (N_38400,N_23851,N_24286);
nor U38401 (N_38401,N_26001,N_29951);
nor U38402 (N_38402,N_28391,N_29782);
xor U38403 (N_38403,N_21362,N_22867);
nand U38404 (N_38404,N_20345,N_20007);
nand U38405 (N_38405,N_28743,N_24318);
nor U38406 (N_38406,N_25474,N_23943);
nand U38407 (N_38407,N_22730,N_21789);
xnor U38408 (N_38408,N_23561,N_21077);
nor U38409 (N_38409,N_26470,N_26671);
nand U38410 (N_38410,N_25100,N_27860);
or U38411 (N_38411,N_24875,N_23719);
nor U38412 (N_38412,N_29756,N_27179);
or U38413 (N_38413,N_20082,N_26078);
and U38414 (N_38414,N_24459,N_22821);
or U38415 (N_38415,N_26340,N_21122);
nand U38416 (N_38416,N_20539,N_26146);
nand U38417 (N_38417,N_21393,N_26367);
nor U38418 (N_38418,N_25916,N_24979);
and U38419 (N_38419,N_26353,N_23784);
nor U38420 (N_38420,N_23012,N_21685);
or U38421 (N_38421,N_24174,N_20399);
or U38422 (N_38422,N_22950,N_22117);
and U38423 (N_38423,N_29030,N_23575);
nand U38424 (N_38424,N_25859,N_20473);
nor U38425 (N_38425,N_23597,N_20736);
and U38426 (N_38426,N_24160,N_20739);
and U38427 (N_38427,N_20710,N_28170);
nor U38428 (N_38428,N_20562,N_26489);
nor U38429 (N_38429,N_28217,N_21393);
nor U38430 (N_38430,N_28613,N_29188);
or U38431 (N_38431,N_24148,N_24406);
and U38432 (N_38432,N_22529,N_27255);
nand U38433 (N_38433,N_21843,N_28593);
nor U38434 (N_38434,N_29239,N_25061);
xnor U38435 (N_38435,N_29379,N_29270);
and U38436 (N_38436,N_22170,N_20257);
and U38437 (N_38437,N_24719,N_28629);
nor U38438 (N_38438,N_23314,N_26617);
and U38439 (N_38439,N_27610,N_21592);
nand U38440 (N_38440,N_22676,N_24857);
nor U38441 (N_38441,N_21410,N_20078);
xor U38442 (N_38442,N_24214,N_26740);
or U38443 (N_38443,N_23599,N_23886);
xnor U38444 (N_38444,N_27918,N_28626);
or U38445 (N_38445,N_24320,N_28966);
or U38446 (N_38446,N_21527,N_25355);
or U38447 (N_38447,N_24744,N_20881);
xnor U38448 (N_38448,N_29357,N_23587);
xor U38449 (N_38449,N_22755,N_29157);
xnor U38450 (N_38450,N_28928,N_26673);
and U38451 (N_38451,N_21967,N_22420);
xor U38452 (N_38452,N_27881,N_23539);
and U38453 (N_38453,N_27950,N_29334);
and U38454 (N_38454,N_28937,N_26865);
or U38455 (N_38455,N_25254,N_29248);
or U38456 (N_38456,N_24099,N_20465);
or U38457 (N_38457,N_28179,N_25052);
xnor U38458 (N_38458,N_26529,N_28372);
xor U38459 (N_38459,N_28067,N_24490);
or U38460 (N_38460,N_26442,N_22204);
nor U38461 (N_38461,N_25837,N_28730);
or U38462 (N_38462,N_20675,N_28495);
or U38463 (N_38463,N_24041,N_29621);
nor U38464 (N_38464,N_27280,N_27057);
and U38465 (N_38465,N_28716,N_24967);
and U38466 (N_38466,N_25467,N_29340);
or U38467 (N_38467,N_22997,N_24336);
nor U38468 (N_38468,N_26054,N_22344);
or U38469 (N_38469,N_22456,N_27664);
or U38470 (N_38470,N_21945,N_28090);
nand U38471 (N_38471,N_25184,N_29311);
and U38472 (N_38472,N_29838,N_21429);
xnor U38473 (N_38473,N_26260,N_26232);
nand U38474 (N_38474,N_23857,N_20988);
and U38475 (N_38475,N_25046,N_25220);
nand U38476 (N_38476,N_23224,N_22828);
and U38477 (N_38477,N_24064,N_28281);
nand U38478 (N_38478,N_28648,N_23474);
nor U38479 (N_38479,N_26773,N_27565);
and U38480 (N_38480,N_21472,N_20899);
nand U38481 (N_38481,N_25463,N_27194);
and U38482 (N_38482,N_24844,N_24116);
and U38483 (N_38483,N_27934,N_29863);
and U38484 (N_38484,N_29336,N_29426);
and U38485 (N_38485,N_20808,N_28996);
nor U38486 (N_38486,N_26801,N_25361);
or U38487 (N_38487,N_28441,N_21041);
nor U38488 (N_38488,N_26546,N_25748);
and U38489 (N_38489,N_21422,N_20030);
and U38490 (N_38490,N_28803,N_29584);
nor U38491 (N_38491,N_28763,N_29294);
nor U38492 (N_38492,N_27164,N_28584);
nand U38493 (N_38493,N_23834,N_20402);
nor U38494 (N_38494,N_27856,N_22443);
or U38495 (N_38495,N_29605,N_20199);
or U38496 (N_38496,N_23762,N_25971);
nor U38497 (N_38497,N_22515,N_28097);
and U38498 (N_38498,N_21318,N_21101);
and U38499 (N_38499,N_27869,N_26673);
nand U38500 (N_38500,N_28552,N_27586);
and U38501 (N_38501,N_25252,N_28536);
nor U38502 (N_38502,N_26960,N_26782);
and U38503 (N_38503,N_26579,N_24509);
or U38504 (N_38504,N_21137,N_27524);
nand U38505 (N_38505,N_20531,N_27767);
nor U38506 (N_38506,N_23330,N_20272);
nand U38507 (N_38507,N_28137,N_29621);
nor U38508 (N_38508,N_26415,N_29550);
and U38509 (N_38509,N_22886,N_22039);
nand U38510 (N_38510,N_28947,N_23024);
nand U38511 (N_38511,N_22882,N_23518);
or U38512 (N_38512,N_26952,N_28306);
nand U38513 (N_38513,N_21903,N_24157);
nand U38514 (N_38514,N_29203,N_26255);
xor U38515 (N_38515,N_27202,N_22313);
or U38516 (N_38516,N_24799,N_25323);
or U38517 (N_38517,N_20710,N_21364);
xnor U38518 (N_38518,N_20709,N_21105);
or U38519 (N_38519,N_26470,N_29989);
and U38520 (N_38520,N_20956,N_23760);
nor U38521 (N_38521,N_26543,N_25903);
nor U38522 (N_38522,N_24391,N_20273);
nand U38523 (N_38523,N_25420,N_20130);
nand U38524 (N_38524,N_23519,N_28266);
nand U38525 (N_38525,N_25764,N_23816);
nand U38526 (N_38526,N_27612,N_22350);
or U38527 (N_38527,N_21352,N_24612);
nand U38528 (N_38528,N_20941,N_27517);
nor U38529 (N_38529,N_25311,N_24054);
nand U38530 (N_38530,N_21845,N_26448);
and U38531 (N_38531,N_25536,N_26100);
and U38532 (N_38532,N_27391,N_26964);
nand U38533 (N_38533,N_26162,N_21659);
and U38534 (N_38534,N_28382,N_28064);
nand U38535 (N_38535,N_25112,N_20985);
nor U38536 (N_38536,N_28054,N_22504);
or U38537 (N_38537,N_23457,N_23821);
and U38538 (N_38538,N_27826,N_20584);
nor U38539 (N_38539,N_23890,N_27142);
nand U38540 (N_38540,N_29857,N_21104);
nor U38541 (N_38541,N_23865,N_24420);
or U38542 (N_38542,N_22371,N_20812);
or U38543 (N_38543,N_26141,N_25642);
nor U38544 (N_38544,N_20163,N_26967);
and U38545 (N_38545,N_28853,N_21029);
nand U38546 (N_38546,N_29269,N_20784);
and U38547 (N_38547,N_29724,N_22207);
nor U38548 (N_38548,N_20436,N_23644);
nor U38549 (N_38549,N_26880,N_29892);
nor U38550 (N_38550,N_22172,N_22906);
and U38551 (N_38551,N_28291,N_26444);
and U38552 (N_38552,N_25500,N_24986);
nor U38553 (N_38553,N_22770,N_24586);
nand U38554 (N_38554,N_20713,N_25062);
and U38555 (N_38555,N_20878,N_29978);
nor U38556 (N_38556,N_29994,N_25509);
or U38557 (N_38557,N_27144,N_28650);
and U38558 (N_38558,N_20034,N_28094);
nand U38559 (N_38559,N_21300,N_27669);
or U38560 (N_38560,N_27654,N_27665);
and U38561 (N_38561,N_27989,N_27241);
nor U38562 (N_38562,N_20026,N_28881);
or U38563 (N_38563,N_20820,N_29955);
nand U38564 (N_38564,N_25356,N_26979);
xnor U38565 (N_38565,N_27086,N_22818);
xor U38566 (N_38566,N_29227,N_25113);
nor U38567 (N_38567,N_24487,N_20196);
xnor U38568 (N_38568,N_25006,N_23322);
nand U38569 (N_38569,N_27160,N_22055);
nor U38570 (N_38570,N_21047,N_21254);
and U38571 (N_38571,N_23083,N_24370);
or U38572 (N_38572,N_29002,N_26393);
and U38573 (N_38573,N_27125,N_21272);
nand U38574 (N_38574,N_22870,N_20229);
and U38575 (N_38575,N_28758,N_28901);
nor U38576 (N_38576,N_24281,N_21430);
xnor U38577 (N_38577,N_24584,N_26006);
nor U38578 (N_38578,N_20020,N_28663);
nand U38579 (N_38579,N_21067,N_25970);
and U38580 (N_38580,N_20142,N_27154);
nand U38581 (N_38581,N_22397,N_28811);
nand U38582 (N_38582,N_24396,N_21131);
and U38583 (N_38583,N_22554,N_20665);
and U38584 (N_38584,N_20779,N_23905);
xnor U38585 (N_38585,N_21303,N_20110);
nand U38586 (N_38586,N_25242,N_20203);
xor U38587 (N_38587,N_28160,N_25636);
nor U38588 (N_38588,N_23278,N_29031);
xor U38589 (N_38589,N_21124,N_29924);
nand U38590 (N_38590,N_26046,N_29484);
or U38591 (N_38591,N_21953,N_23891);
nand U38592 (N_38592,N_21910,N_22947);
nand U38593 (N_38593,N_25030,N_27863);
nor U38594 (N_38594,N_21408,N_28568);
nor U38595 (N_38595,N_28278,N_29339);
nor U38596 (N_38596,N_25216,N_23178);
nor U38597 (N_38597,N_24235,N_23417);
nand U38598 (N_38598,N_25204,N_27392);
xnor U38599 (N_38599,N_26253,N_29099);
and U38600 (N_38600,N_26036,N_29959);
and U38601 (N_38601,N_20876,N_24432);
xnor U38602 (N_38602,N_27025,N_22377);
and U38603 (N_38603,N_29793,N_24166);
or U38604 (N_38604,N_22615,N_29782);
nor U38605 (N_38605,N_23762,N_23896);
and U38606 (N_38606,N_20226,N_25875);
or U38607 (N_38607,N_21652,N_25358);
nor U38608 (N_38608,N_29725,N_25191);
and U38609 (N_38609,N_21973,N_20864);
nand U38610 (N_38610,N_28003,N_24114);
xnor U38611 (N_38611,N_29758,N_25566);
nor U38612 (N_38612,N_27471,N_27694);
and U38613 (N_38613,N_21128,N_27633);
nand U38614 (N_38614,N_27661,N_23394);
and U38615 (N_38615,N_28058,N_29149);
or U38616 (N_38616,N_26337,N_27647);
or U38617 (N_38617,N_29088,N_25730);
nand U38618 (N_38618,N_22702,N_27671);
and U38619 (N_38619,N_23430,N_22766);
or U38620 (N_38620,N_20714,N_27416);
and U38621 (N_38621,N_25468,N_22120);
and U38622 (N_38622,N_25155,N_26111);
and U38623 (N_38623,N_20437,N_27630);
nand U38624 (N_38624,N_21321,N_26148);
nor U38625 (N_38625,N_26330,N_23806);
or U38626 (N_38626,N_21873,N_29903);
nand U38627 (N_38627,N_27489,N_21274);
and U38628 (N_38628,N_26922,N_28084);
nor U38629 (N_38629,N_22836,N_21457);
or U38630 (N_38630,N_27558,N_26402);
nand U38631 (N_38631,N_23780,N_24068);
nor U38632 (N_38632,N_25308,N_22980);
nand U38633 (N_38633,N_21908,N_23267);
nor U38634 (N_38634,N_21517,N_23217);
xor U38635 (N_38635,N_29942,N_26914);
xnor U38636 (N_38636,N_29436,N_28017);
nand U38637 (N_38637,N_28377,N_27101);
and U38638 (N_38638,N_20198,N_26218);
nor U38639 (N_38639,N_25207,N_29751);
and U38640 (N_38640,N_23242,N_29697);
nor U38641 (N_38641,N_22229,N_20535);
nand U38642 (N_38642,N_29067,N_21329);
nor U38643 (N_38643,N_27154,N_24082);
and U38644 (N_38644,N_23245,N_29675);
and U38645 (N_38645,N_26413,N_27621);
and U38646 (N_38646,N_29999,N_29740);
or U38647 (N_38647,N_24290,N_21637);
nand U38648 (N_38648,N_22795,N_26909);
xnor U38649 (N_38649,N_25136,N_26565);
or U38650 (N_38650,N_25499,N_24470);
nand U38651 (N_38651,N_25329,N_27864);
or U38652 (N_38652,N_28159,N_26912);
and U38653 (N_38653,N_29685,N_29369);
and U38654 (N_38654,N_21985,N_23986);
nand U38655 (N_38655,N_20742,N_27049);
and U38656 (N_38656,N_21256,N_25377);
nand U38657 (N_38657,N_25147,N_29570);
and U38658 (N_38658,N_27198,N_29126);
and U38659 (N_38659,N_21609,N_29302);
and U38660 (N_38660,N_22811,N_28416);
and U38661 (N_38661,N_25193,N_21708);
nand U38662 (N_38662,N_28737,N_20111);
nand U38663 (N_38663,N_23739,N_28207);
xor U38664 (N_38664,N_20319,N_28205);
and U38665 (N_38665,N_24320,N_29412);
nor U38666 (N_38666,N_21179,N_28214);
nand U38667 (N_38667,N_22659,N_23030);
nand U38668 (N_38668,N_22503,N_28916);
xnor U38669 (N_38669,N_23489,N_28622);
or U38670 (N_38670,N_24550,N_29857);
nand U38671 (N_38671,N_20387,N_20814);
or U38672 (N_38672,N_26360,N_29784);
nand U38673 (N_38673,N_23798,N_20036);
nand U38674 (N_38674,N_29411,N_22177);
xnor U38675 (N_38675,N_24467,N_21846);
and U38676 (N_38676,N_24926,N_26703);
or U38677 (N_38677,N_29684,N_26781);
or U38678 (N_38678,N_21132,N_20537);
or U38679 (N_38679,N_24758,N_22907);
nand U38680 (N_38680,N_21287,N_25399);
or U38681 (N_38681,N_29695,N_20991);
or U38682 (N_38682,N_27240,N_20266);
nand U38683 (N_38683,N_24730,N_24180);
or U38684 (N_38684,N_23946,N_26710);
xor U38685 (N_38685,N_29840,N_27577);
or U38686 (N_38686,N_22993,N_26172);
xnor U38687 (N_38687,N_22189,N_27555);
and U38688 (N_38688,N_27414,N_21076);
nor U38689 (N_38689,N_27868,N_24083);
and U38690 (N_38690,N_22722,N_24997);
and U38691 (N_38691,N_28760,N_21740);
or U38692 (N_38692,N_21361,N_29224);
nand U38693 (N_38693,N_22817,N_20637);
and U38694 (N_38694,N_22416,N_25293);
nor U38695 (N_38695,N_29586,N_20380);
nand U38696 (N_38696,N_29378,N_24649);
or U38697 (N_38697,N_25546,N_25037);
nor U38698 (N_38698,N_27684,N_21612);
nand U38699 (N_38699,N_20077,N_28954);
or U38700 (N_38700,N_26650,N_29043);
and U38701 (N_38701,N_29404,N_21930);
or U38702 (N_38702,N_28018,N_28489);
xnor U38703 (N_38703,N_27341,N_27880);
and U38704 (N_38704,N_27178,N_21817);
and U38705 (N_38705,N_27336,N_23705);
nor U38706 (N_38706,N_23397,N_23092);
nand U38707 (N_38707,N_20597,N_29757);
nor U38708 (N_38708,N_29553,N_24035);
nand U38709 (N_38709,N_23306,N_26414);
or U38710 (N_38710,N_22747,N_26562);
nor U38711 (N_38711,N_20612,N_26945);
xor U38712 (N_38712,N_22347,N_24693);
or U38713 (N_38713,N_27657,N_27236);
and U38714 (N_38714,N_20663,N_29568);
or U38715 (N_38715,N_23431,N_24433);
xor U38716 (N_38716,N_22314,N_28999);
or U38717 (N_38717,N_26615,N_20342);
or U38718 (N_38718,N_20700,N_25788);
or U38719 (N_38719,N_26166,N_24320);
and U38720 (N_38720,N_28642,N_26062);
or U38721 (N_38721,N_22565,N_25099);
and U38722 (N_38722,N_26243,N_20318);
nor U38723 (N_38723,N_20662,N_20132);
and U38724 (N_38724,N_28158,N_22625);
or U38725 (N_38725,N_26198,N_29010);
or U38726 (N_38726,N_28865,N_26950);
xnor U38727 (N_38727,N_28854,N_22215);
and U38728 (N_38728,N_29906,N_21324);
nor U38729 (N_38729,N_23991,N_29613);
nor U38730 (N_38730,N_20077,N_23888);
nand U38731 (N_38731,N_27159,N_29841);
or U38732 (N_38732,N_22582,N_23297);
xnor U38733 (N_38733,N_27185,N_27348);
xnor U38734 (N_38734,N_23003,N_27370);
nor U38735 (N_38735,N_26467,N_29543);
or U38736 (N_38736,N_20468,N_28911);
and U38737 (N_38737,N_23855,N_23686);
nor U38738 (N_38738,N_24568,N_20970);
and U38739 (N_38739,N_20544,N_26048);
nand U38740 (N_38740,N_21310,N_25133);
and U38741 (N_38741,N_27443,N_28604);
nor U38742 (N_38742,N_27941,N_21386);
or U38743 (N_38743,N_28621,N_27399);
or U38744 (N_38744,N_28402,N_23437);
or U38745 (N_38745,N_22792,N_29268);
nand U38746 (N_38746,N_21258,N_28635);
or U38747 (N_38747,N_27131,N_29547);
and U38748 (N_38748,N_23979,N_28907);
nand U38749 (N_38749,N_22685,N_26296);
and U38750 (N_38750,N_22098,N_22902);
and U38751 (N_38751,N_22006,N_20426);
nand U38752 (N_38752,N_25242,N_20642);
or U38753 (N_38753,N_26032,N_28909);
xnor U38754 (N_38754,N_20956,N_26697);
and U38755 (N_38755,N_25954,N_22586);
xnor U38756 (N_38756,N_25137,N_25785);
or U38757 (N_38757,N_25142,N_22686);
or U38758 (N_38758,N_28876,N_29166);
nand U38759 (N_38759,N_27866,N_21395);
and U38760 (N_38760,N_21146,N_20933);
nor U38761 (N_38761,N_29897,N_20002);
nor U38762 (N_38762,N_29907,N_23286);
nor U38763 (N_38763,N_22523,N_23944);
nor U38764 (N_38764,N_25786,N_29109);
nor U38765 (N_38765,N_25582,N_21904);
or U38766 (N_38766,N_20344,N_23958);
nand U38767 (N_38767,N_26526,N_26169);
xnor U38768 (N_38768,N_26377,N_27191);
and U38769 (N_38769,N_21498,N_20735);
or U38770 (N_38770,N_26769,N_25619);
and U38771 (N_38771,N_22424,N_20776);
xnor U38772 (N_38772,N_28547,N_29034);
nand U38773 (N_38773,N_23885,N_21932);
nor U38774 (N_38774,N_26079,N_21132);
and U38775 (N_38775,N_26769,N_25417);
nor U38776 (N_38776,N_29334,N_22573);
nor U38777 (N_38777,N_21240,N_27233);
nor U38778 (N_38778,N_27212,N_24028);
nand U38779 (N_38779,N_27056,N_26806);
or U38780 (N_38780,N_27485,N_27076);
and U38781 (N_38781,N_27946,N_24324);
nand U38782 (N_38782,N_23559,N_21470);
or U38783 (N_38783,N_29092,N_27013);
and U38784 (N_38784,N_20459,N_22623);
and U38785 (N_38785,N_25352,N_27115);
or U38786 (N_38786,N_28307,N_22355);
nand U38787 (N_38787,N_20811,N_27462);
nor U38788 (N_38788,N_29856,N_27009);
and U38789 (N_38789,N_29548,N_29818);
and U38790 (N_38790,N_29954,N_22019);
and U38791 (N_38791,N_20778,N_25489);
xor U38792 (N_38792,N_26765,N_27598);
nand U38793 (N_38793,N_21556,N_20733);
or U38794 (N_38794,N_28409,N_27443);
and U38795 (N_38795,N_21324,N_23000);
or U38796 (N_38796,N_28756,N_20937);
nand U38797 (N_38797,N_27497,N_27243);
xnor U38798 (N_38798,N_24826,N_24296);
or U38799 (N_38799,N_23138,N_23771);
nand U38800 (N_38800,N_22794,N_25813);
and U38801 (N_38801,N_25825,N_28398);
xor U38802 (N_38802,N_24104,N_24296);
xnor U38803 (N_38803,N_20511,N_24975);
and U38804 (N_38804,N_23673,N_21323);
xnor U38805 (N_38805,N_23471,N_28098);
and U38806 (N_38806,N_29641,N_25081);
nor U38807 (N_38807,N_29842,N_23625);
and U38808 (N_38808,N_21799,N_20350);
or U38809 (N_38809,N_20388,N_27099);
and U38810 (N_38810,N_22632,N_23964);
nor U38811 (N_38811,N_23623,N_22471);
or U38812 (N_38812,N_26760,N_20534);
nand U38813 (N_38813,N_25998,N_20569);
nor U38814 (N_38814,N_22336,N_26469);
or U38815 (N_38815,N_21340,N_22356);
and U38816 (N_38816,N_23609,N_22114);
or U38817 (N_38817,N_28029,N_26483);
nor U38818 (N_38818,N_27227,N_22434);
and U38819 (N_38819,N_24665,N_29617);
or U38820 (N_38820,N_26471,N_26558);
nand U38821 (N_38821,N_21790,N_22550);
and U38822 (N_38822,N_23420,N_25922);
nor U38823 (N_38823,N_23969,N_25470);
or U38824 (N_38824,N_23772,N_22147);
nand U38825 (N_38825,N_24399,N_24958);
xnor U38826 (N_38826,N_28286,N_27933);
nand U38827 (N_38827,N_25722,N_27985);
and U38828 (N_38828,N_21904,N_21693);
nor U38829 (N_38829,N_26289,N_25644);
nor U38830 (N_38830,N_23592,N_20384);
or U38831 (N_38831,N_26806,N_27094);
and U38832 (N_38832,N_24081,N_20426);
nand U38833 (N_38833,N_24512,N_28559);
nor U38834 (N_38834,N_26430,N_24784);
nand U38835 (N_38835,N_24766,N_23330);
xor U38836 (N_38836,N_25193,N_20222);
nor U38837 (N_38837,N_24719,N_22859);
and U38838 (N_38838,N_28421,N_24258);
and U38839 (N_38839,N_22062,N_27663);
and U38840 (N_38840,N_27068,N_21105);
xnor U38841 (N_38841,N_24475,N_24997);
nor U38842 (N_38842,N_23139,N_21461);
nor U38843 (N_38843,N_28545,N_20668);
xor U38844 (N_38844,N_20235,N_24287);
xnor U38845 (N_38845,N_25530,N_29013);
nor U38846 (N_38846,N_29857,N_29672);
and U38847 (N_38847,N_24728,N_21993);
nor U38848 (N_38848,N_22362,N_28591);
nand U38849 (N_38849,N_20889,N_25905);
and U38850 (N_38850,N_26010,N_24202);
and U38851 (N_38851,N_23965,N_27289);
nand U38852 (N_38852,N_20968,N_27490);
or U38853 (N_38853,N_23170,N_28377);
and U38854 (N_38854,N_20732,N_20745);
xor U38855 (N_38855,N_29987,N_28313);
nor U38856 (N_38856,N_20468,N_29518);
xor U38857 (N_38857,N_23313,N_27326);
nor U38858 (N_38858,N_22593,N_27911);
or U38859 (N_38859,N_21471,N_25995);
nand U38860 (N_38860,N_24436,N_23660);
and U38861 (N_38861,N_26189,N_25438);
or U38862 (N_38862,N_27617,N_26443);
and U38863 (N_38863,N_28995,N_23091);
nor U38864 (N_38864,N_22894,N_21956);
nor U38865 (N_38865,N_25435,N_28453);
nor U38866 (N_38866,N_26876,N_24377);
nand U38867 (N_38867,N_23952,N_25961);
or U38868 (N_38868,N_26356,N_27804);
or U38869 (N_38869,N_24189,N_22117);
and U38870 (N_38870,N_22764,N_25170);
xor U38871 (N_38871,N_21415,N_21254);
nand U38872 (N_38872,N_25974,N_26557);
nand U38873 (N_38873,N_25189,N_22648);
nor U38874 (N_38874,N_27409,N_29077);
xnor U38875 (N_38875,N_27096,N_23262);
xor U38876 (N_38876,N_24102,N_24842);
or U38877 (N_38877,N_28645,N_22722);
or U38878 (N_38878,N_25622,N_24504);
xor U38879 (N_38879,N_22073,N_26674);
nand U38880 (N_38880,N_21933,N_22696);
nor U38881 (N_38881,N_23918,N_22404);
nand U38882 (N_38882,N_28168,N_21381);
nand U38883 (N_38883,N_24397,N_22188);
or U38884 (N_38884,N_20717,N_26161);
nand U38885 (N_38885,N_20492,N_29319);
and U38886 (N_38886,N_21427,N_29804);
nand U38887 (N_38887,N_26627,N_23713);
nand U38888 (N_38888,N_27314,N_28146);
nor U38889 (N_38889,N_29091,N_28056);
and U38890 (N_38890,N_22863,N_24259);
nand U38891 (N_38891,N_28193,N_27892);
or U38892 (N_38892,N_27242,N_28332);
nand U38893 (N_38893,N_27240,N_27835);
xor U38894 (N_38894,N_21535,N_29316);
and U38895 (N_38895,N_23891,N_29429);
nand U38896 (N_38896,N_23145,N_23201);
nand U38897 (N_38897,N_28937,N_27209);
or U38898 (N_38898,N_20458,N_29911);
nor U38899 (N_38899,N_25413,N_23632);
and U38900 (N_38900,N_29385,N_27588);
nor U38901 (N_38901,N_22456,N_27149);
nand U38902 (N_38902,N_23830,N_28154);
nor U38903 (N_38903,N_26685,N_27003);
or U38904 (N_38904,N_25793,N_23298);
and U38905 (N_38905,N_29685,N_29434);
or U38906 (N_38906,N_23522,N_22543);
nor U38907 (N_38907,N_28839,N_23521);
or U38908 (N_38908,N_29806,N_25723);
nor U38909 (N_38909,N_27467,N_24573);
nand U38910 (N_38910,N_29184,N_21522);
or U38911 (N_38911,N_22299,N_20538);
or U38912 (N_38912,N_21245,N_29571);
or U38913 (N_38913,N_21982,N_20163);
or U38914 (N_38914,N_22938,N_28341);
xnor U38915 (N_38915,N_26399,N_25766);
and U38916 (N_38916,N_23097,N_24512);
nor U38917 (N_38917,N_23116,N_25885);
or U38918 (N_38918,N_23944,N_24191);
nor U38919 (N_38919,N_29408,N_21299);
or U38920 (N_38920,N_20568,N_28666);
nand U38921 (N_38921,N_26079,N_26641);
nand U38922 (N_38922,N_21466,N_20696);
nand U38923 (N_38923,N_25649,N_28456);
nor U38924 (N_38924,N_29726,N_20944);
xnor U38925 (N_38925,N_27659,N_26762);
nand U38926 (N_38926,N_29350,N_24431);
nand U38927 (N_38927,N_28848,N_22947);
or U38928 (N_38928,N_26079,N_28940);
or U38929 (N_38929,N_23848,N_21017);
nand U38930 (N_38930,N_22441,N_28840);
nor U38931 (N_38931,N_26316,N_20665);
nor U38932 (N_38932,N_26503,N_27516);
and U38933 (N_38933,N_28079,N_21646);
nor U38934 (N_38934,N_26910,N_27111);
or U38935 (N_38935,N_20666,N_24818);
nand U38936 (N_38936,N_25060,N_23596);
or U38937 (N_38937,N_28719,N_27251);
or U38938 (N_38938,N_24947,N_20239);
and U38939 (N_38939,N_27801,N_21700);
or U38940 (N_38940,N_24567,N_21139);
nor U38941 (N_38941,N_22466,N_20960);
xor U38942 (N_38942,N_25168,N_29511);
nand U38943 (N_38943,N_28099,N_24040);
and U38944 (N_38944,N_25527,N_24741);
and U38945 (N_38945,N_23418,N_25839);
nor U38946 (N_38946,N_20946,N_29159);
and U38947 (N_38947,N_28012,N_29248);
and U38948 (N_38948,N_23009,N_29514);
nor U38949 (N_38949,N_22134,N_28525);
and U38950 (N_38950,N_25651,N_28641);
and U38951 (N_38951,N_28913,N_22432);
or U38952 (N_38952,N_22781,N_27331);
or U38953 (N_38953,N_24910,N_24456);
nand U38954 (N_38954,N_27854,N_22390);
or U38955 (N_38955,N_24725,N_29862);
xnor U38956 (N_38956,N_28308,N_28910);
and U38957 (N_38957,N_23892,N_26958);
or U38958 (N_38958,N_21175,N_21987);
nor U38959 (N_38959,N_23316,N_24151);
and U38960 (N_38960,N_29037,N_28263);
or U38961 (N_38961,N_24673,N_25309);
or U38962 (N_38962,N_23856,N_22875);
and U38963 (N_38963,N_29633,N_21878);
nand U38964 (N_38964,N_24821,N_24597);
xor U38965 (N_38965,N_27609,N_25524);
and U38966 (N_38966,N_21297,N_29918);
nor U38967 (N_38967,N_29542,N_24641);
nor U38968 (N_38968,N_25511,N_21386);
nor U38969 (N_38969,N_28319,N_29718);
nor U38970 (N_38970,N_20805,N_24178);
xor U38971 (N_38971,N_27119,N_29885);
or U38972 (N_38972,N_24013,N_26578);
nand U38973 (N_38973,N_23588,N_25590);
and U38974 (N_38974,N_20283,N_27806);
or U38975 (N_38975,N_20855,N_20590);
nor U38976 (N_38976,N_26971,N_23873);
xor U38977 (N_38977,N_20561,N_20154);
nor U38978 (N_38978,N_28613,N_22018);
or U38979 (N_38979,N_20459,N_20135);
and U38980 (N_38980,N_23525,N_29088);
and U38981 (N_38981,N_23930,N_25851);
nand U38982 (N_38982,N_28756,N_21297);
nor U38983 (N_38983,N_27481,N_23789);
xor U38984 (N_38984,N_25636,N_22620);
nand U38985 (N_38985,N_21089,N_29679);
xor U38986 (N_38986,N_21856,N_24809);
nor U38987 (N_38987,N_21328,N_27401);
nor U38988 (N_38988,N_25315,N_22859);
nand U38989 (N_38989,N_20575,N_23889);
and U38990 (N_38990,N_20360,N_22011);
nor U38991 (N_38991,N_25437,N_26823);
or U38992 (N_38992,N_21020,N_24065);
nand U38993 (N_38993,N_26375,N_24616);
or U38994 (N_38994,N_24164,N_25771);
and U38995 (N_38995,N_20202,N_22241);
or U38996 (N_38996,N_22477,N_20108);
or U38997 (N_38997,N_21333,N_22092);
nand U38998 (N_38998,N_21950,N_24580);
xor U38999 (N_38999,N_28643,N_24851);
nand U39000 (N_39000,N_26179,N_25615);
or U39001 (N_39001,N_21652,N_25872);
or U39002 (N_39002,N_26108,N_20857);
nand U39003 (N_39003,N_20893,N_23950);
nor U39004 (N_39004,N_23551,N_28199);
and U39005 (N_39005,N_26427,N_21060);
and U39006 (N_39006,N_27756,N_24415);
xnor U39007 (N_39007,N_28311,N_28101);
nor U39008 (N_39008,N_23023,N_20636);
and U39009 (N_39009,N_24314,N_20954);
and U39010 (N_39010,N_22135,N_23923);
nor U39011 (N_39011,N_20935,N_21024);
or U39012 (N_39012,N_25641,N_24084);
and U39013 (N_39013,N_24340,N_26504);
nand U39014 (N_39014,N_27892,N_22909);
nor U39015 (N_39015,N_22223,N_29190);
and U39016 (N_39016,N_25904,N_22678);
nand U39017 (N_39017,N_20516,N_26944);
nand U39018 (N_39018,N_21375,N_21370);
or U39019 (N_39019,N_21204,N_29896);
nand U39020 (N_39020,N_20051,N_28613);
nand U39021 (N_39021,N_23586,N_24125);
nor U39022 (N_39022,N_25517,N_25500);
and U39023 (N_39023,N_20521,N_29734);
nor U39024 (N_39024,N_20453,N_24475);
nor U39025 (N_39025,N_22814,N_25748);
and U39026 (N_39026,N_27820,N_28821);
nor U39027 (N_39027,N_22854,N_21316);
and U39028 (N_39028,N_22113,N_23903);
nand U39029 (N_39029,N_23586,N_22275);
and U39030 (N_39030,N_27808,N_25490);
nor U39031 (N_39031,N_28173,N_23672);
or U39032 (N_39032,N_21586,N_27414);
xnor U39033 (N_39033,N_27372,N_23982);
and U39034 (N_39034,N_25527,N_23564);
and U39035 (N_39035,N_27697,N_23874);
xnor U39036 (N_39036,N_20986,N_25461);
and U39037 (N_39037,N_28505,N_24074);
and U39038 (N_39038,N_26738,N_22008);
nand U39039 (N_39039,N_26897,N_22235);
nand U39040 (N_39040,N_20425,N_20894);
and U39041 (N_39041,N_29956,N_28070);
or U39042 (N_39042,N_25587,N_28358);
or U39043 (N_39043,N_20975,N_26800);
nand U39044 (N_39044,N_28213,N_20336);
and U39045 (N_39045,N_24864,N_20248);
nor U39046 (N_39046,N_28768,N_27954);
or U39047 (N_39047,N_29820,N_27146);
and U39048 (N_39048,N_24435,N_20696);
nand U39049 (N_39049,N_28429,N_27861);
nor U39050 (N_39050,N_22430,N_20357);
and U39051 (N_39051,N_28120,N_27694);
nor U39052 (N_39052,N_23015,N_27824);
or U39053 (N_39053,N_28429,N_29931);
nor U39054 (N_39054,N_22853,N_23511);
nor U39055 (N_39055,N_24821,N_26761);
nor U39056 (N_39056,N_26411,N_22292);
and U39057 (N_39057,N_27051,N_27195);
nand U39058 (N_39058,N_23000,N_25056);
nand U39059 (N_39059,N_23532,N_26811);
xor U39060 (N_39060,N_22196,N_26466);
xor U39061 (N_39061,N_26552,N_22142);
and U39062 (N_39062,N_29530,N_21896);
nor U39063 (N_39063,N_21957,N_22417);
or U39064 (N_39064,N_24098,N_21188);
nor U39065 (N_39065,N_23889,N_26923);
nand U39066 (N_39066,N_22341,N_22564);
nor U39067 (N_39067,N_20387,N_21069);
nor U39068 (N_39068,N_21547,N_25728);
nor U39069 (N_39069,N_29017,N_29215);
and U39070 (N_39070,N_27813,N_20290);
xnor U39071 (N_39071,N_26584,N_21293);
xnor U39072 (N_39072,N_21781,N_27864);
nor U39073 (N_39073,N_21854,N_27626);
or U39074 (N_39074,N_27384,N_25831);
or U39075 (N_39075,N_29558,N_28609);
and U39076 (N_39076,N_25962,N_20405);
nand U39077 (N_39077,N_22591,N_26435);
xor U39078 (N_39078,N_23962,N_23207);
nor U39079 (N_39079,N_22538,N_28602);
nor U39080 (N_39080,N_20596,N_29496);
nand U39081 (N_39081,N_26995,N_27627);
nand U39082 (N_39082,N_21745,N_28040);
xnor U39083 (N_39083,N_20661,N_21755);
nor U39084 (N_39084,N_28995,N_27655);
or U39085 (N_39085,N_26023,N_20892);
nand U39086 (N_39086,N_27155,N_29988);
or U39087 (N_39087,N_24243,N_24840);
or U39088 (N_39088,N_26431,N_27383);
or U39089 (N_39089,N_25144,N_23118);
and U39090 (N_39090,N_25489,N_20480);
nand U39091 (N_39091,N_24038,N_22342);
and U39092 (N_39092,N_25988,N_29391);
nand U39093 (N_39093,N_26048,N_28599);
or U39094 (N_39094,N_28740,N_27499);
or U39095 (N_39095,N_21128,N_22498);
nand U39096 (N_39096,N_20477,N_29622);
or U39097 (N_39097,N_23212,N_23387);
nor U39098 (N_39098,N_24692,N_27308);
xor U39099 (N_39099,N_27566,N_26781);
nand U39100 (N_39100,N_25593,N_29513);
nor U39101 (N_39101,N_25113,N_28753);
or U39102 (N_39102,N_27539,N_22212);
xor U39103 (N_39103,N_20888,N_27477);
nand U39104 (N_39104,N_27452,N_27454);
and U39105 (N_39105,N_25508,N_22858);
nor U39106 (N_39106,N_29536,N_20230);
nor U39107 (N_39107,N_24654,N_22650);
or U39108 (N_39108,N_21034,N_22393);
and U39109 (N_39109,N_23970,N_26084);
or U39110 (N_39110,N_26030,N_27840);
or U39111 (N_39111,N_23359,N_27159);
nand U39112 (N_39112,N_20970,N_29983);
nand U39113 (N_39113,N_20689,N_29918);
or U39114 (N_39114,N_27222,N_26056);
or U39115 (N_39115,N_28564,N_23013);
xor U39116 (N_39116,N_21816,N_28234);
and U39117 (N_39117,N_25965,N_27898);
nor U39118 (N_39118,N_23415,N_23773);
or U39119 (N_39119,N_27872,N_21582);
and U39120 (N_39120,N_25097,N_26959);
and U39121 (N_39121,N_21024,N_27063);
nor U39122 (N_39122,N_21621,N_26752);
and U39123 (N_39123,N_20267,N_20354);
nand U39124 (N_39124,N_28382,N_26261);
xor U39125 (N_39125,N_28876,N_23935);
xnor U39126 (N_39126,N_27789,N_22996);
or U39127 (N_39127,N_26986,N_20112);
or U39128 (N_39128,N_22847,N_29523);
nand U39129 (N_39129,N_21662,N_23275);
xnor U39130 (N_39130,N_25782,N_22044);
nand U39131 (N_39131,N_22531,N_21679);
and U39132 (N_39132,N_23347,N_25220);
nor U39133 (N_39133,N_23942,N_21303);
nor U39134 (N_39134,N_22133,N_22375);
and U39135 (N_39135,N_22414,N_24399);
or U39136 (N_39136,N_29032,N_26175);
nor U39137 (N_39137,N_24743,N_25844);
nand U39138 (N_39138,N_25508,N_28710);
nand U39139 (N_39139,N_28328,N_27949);
nor U39140 (N_39140,N_29782,N_25457);
or U39141 (N_39141,N_23308,N_23394);
nor U39142 (N_39142,N_21310,N_27987);
and U39143 (N_39143,N_22300,N_22502);
nand U39144 (N_39144,N_20356,N_28156);
or U39145 (N_39145,N_26014,N_20644);
or U39146 (N_39146,N_28033,N_21909);
nand U39147 (N_39147,N_20338,N_28307);
and U39148 (N_39148,N_20035,N_22603);
nor U39149 (N_39149,N_24549,N_26789);
nand U39150 (N_39150,N_21718,N_29873);
xnor U39151 (N_39151,N_23252,N_29442);
nor U39152 (N_39152,N_24196,N_28279);
or U39153 (N_39153,N_26100,N_25509);
nor U39154 (N_39154,N_28441,N_27610);
nor U39155 (N_39155,N_25193,N_26836);
nor U39156 (N_39156,N_26575,N_20053);
or U39157 (N_39157,N_22253,N_26287);
xor U39158 (N_39158,N_29884,N_20709);
nor U39159 (N_39159,N_29693,N_25771);
nand U39160 (N_39160,N_28077,N_24693);
xor U39161 (N_39161,N_24226,N_28449);
and U39162 (N_39162,N_21717,N_25511);
nand U39163 (N_39163,N_20874,N_24414);
and U39164 (N_39164,N_29297,N_27595);
nand U39165 (N_39165,N_26946,N_29286);
or U39166 (N_39166,N_21730,N_21209);
or U39167 (N_39167,N_20096,N_29185);
nand U39168 (N_39168,N_28676,N_20736);
nand U39169 (N_39169,N_28984,N_22077);
nand U39170 (N_39170,N_24873,N_20765);
or U39171 (N_39171,N_27031,N_28680);
nor U39172 (N_39172,N_23322,N_24396);
nand U39173 (N_39173,N_24856,N_22522);
or U39174 (N_39174,N_27821,N_29180);
xnor U39175 (N_39175,N_24320,N_28772);
nand U39176 (N_39176,N_29989,N_25680);
or U39177 (N_39177,N_28883,N_27411);
or U39178 (N_39178,N_28541,N_28001);
xnor U39179 (N_39179,N_20431,N_27452);
or U39180 (N_39180,N_21740,N_25440);
nand U39181 (N_39181,N_28402,N_20477);
and U39182 (N_39182,N_28097,N_29002);
nor U39183 (N_39183,N_22195,N_24666);
xnor U39184 (N_39184,N_21733,N_22635);
xor U39185 (N_39185,N_23385,N_21784);
nor U39186 (N_39186,N_23843,N_26898);
xnor U39187 (N_39187,N_26804,N_28236);
and U39188 (N_39188,N_20127,N_21627);
or U39189 (N_39189,N_29005,N_27234);
nand U39190 (N_39190,N_20518,N_24566);
nor U39191 (N_39191,N_26374,N_29437);
nor U39192 (N_39192,N_22244,N_22848);
and U39193 (N_39193,N_22083,N_21432);
nand U39194 (N_39194,N_26096,N_20090);
and U39195 (N_39195,N_25821,N_23714);
and U39196 (N_39196,N_26536,N_20871);
or U39197 (N_39197,N_25158,N_21563);
nand U39198 (N_39198,N_20959,N_21879);
nor U39199 (N_39199,N_26666,N_28283);
nand U39200 (N_39200,N_22525,N_27147);
or U39201 (N_39201,N_25152,N_27661);
nor U39202 (N_39202,N_26685,N_25507);
nand U39203 (N_39203,N_25152,N_23084);
nand U39204 (N_39204,N_28954,N_24291);
nand U39205 (N_39205,N_21100,N_24691);
nand U39206 (N_39206,N_27931,N_28838);
and U39207 (N_39207,N_28938,N_25714);
xor U39208 (N_39208,N_24293,N_22561);
nand U39209 (N_39209,N_24258,N_28539);
nand U39210 (N_39210,N_26237,N_20079);
nor U39211 (N_39211,N_25046,N_28997);
and U39212 (N_39212,N_25009,N_25661);
and U39213 (N_39213,N_22263,N_24092);
nor U39214 (N_39214,N_21488,N_22430);
or U39215 (N_39215,N_29869,N_28880);
or U39216 (N_39216,N_29954,N_21861);
nand U39217 (N_39217,N_27433,N_21081);
nand U39218 (N_39218,N_28690,N_20793);
or U39219 (N_39219,N_20973,N_21263);
xor U39220 (N_39220,N_23319,N_29868);
or U39221 (N_39221,N_27641,N_20421);
xor U39222 (N_39222,N_29928,N_21925);
or U39223 (N_39223,N_26575,N_27697);
nand U39224 (N_39224,N_27106,N_29250);
nand U39225 (N_39225,N_22411,N_21321);
and U39226 (N_39226,N_27415,N_25303);
nand U39227 (N_39227,N_22785,N_26282);
nor U39228 (N_39228,N_29545,N_28271);
xor U39229 (N_39229,N_20831,N_22893);
xor U39230 (N_39230,N_24875,N_28389);
and U39231 (N_39231,N_22768,N_28991);
nand U39232 (N_39232,N_20215,N_20942);
and U39233 (N_39233,N_25416,N_28798);
nand U39234 (N_39234,N_26958,N_27512);
xor U39235 (N_39235,N_20262,N_28007);
or U39236 (N_39236,N_23441,N_24070);
or U39237 (N_39237,N_20247,N_20990);
nor U39238 (N_39238,N_21003,N_21427);
xor U39239 (N_39239,N_23221,N_22672);
nor U39240 (N_39240,N_20922,N_24503);
xnor U39241 (N_39241,N_20671,N_28025);
nor U39242 (N_39242,N_21086,N_28540);
or U39243 (N_39243,N_26103,N_28062);
or U39244 (N_39244,N_28410,N_21778);
or U39245 (N_39245,N_27537,N_21669);
nand U39246 (N_39246,N_27838,N_20025);
and U39247 (N_39247,N_24217,N_20621);
and U39248 (N_39248,N_28337,N_24176);
or U39249 (N_39249,N_21106,N_22121);
nor U39250 (N_39250,N_24266,N_24725);
nor U39251 (N_39251,N_29259,N_28095);
nor U39252 (N_39252,N_27846,N_24975);
nand U39253 (N_39253,N_22020,N_23693);
or U39254 (N_39254,N_20969,N_20716);
or U39255 (N_39255,N_28188,N_25363);
xor U39256 (N_39256,N_20406,N_22553);
and U39257 (N_39257,N_28217,N_20583);
xnor U39258 (N_39258,N_27437,N_28390);
nor U39259 (N_39259,N_29334,N_28856);
nor U39260 (N_39260,N_29947,N_26442);
or U39261 (N_39261,N_22215,N_25654);
and U39262 (N_39262,N_27578,N_21058);
and U39263 (N_39263,N_20770,N_28597);
nor U39264 (N_39264,N_28844,N_28913);
or U39265 (N_39265,N_28810,N_20939);
and U39266 (N_39266,N_21890,N_26393);
xnor U39267 (N_39267,N_25269,N_20016);
nand U39268 (N_39268,N_27758,N_27164);
nand U39269 (N_39269,N_22501,N_29890);
nor U39270 (N_39270,N_28956,N_25405);
and U39271 (N_39271,N_26751,N_29324);
or U39272 (N_39272,N_20005,N_25933);
or U39273 (N_39273,N_20935,N_28738);
or U39274 (N_39274,N_25268,N_22203);
and U39275 (N_39275,N_27027,N_24675);
or U39276 (N_39276,N_28448,N_23174);
nand U39277 (N_39277,N_21451,N_28659);
nor U39278 (N_39278,N_28460,N_20341);
nor U39279 (N_39279,N_28530,N_27713);
nand U39280 (N_39280,N_20391,N_20749);
or U39281 (N_39281,N_26300,N_25320);
nand U39282 (N_39282,N_27933,N_22490);
nor U39283 (N_39283,N_20720,N_27898);
or U39284 (N_39284,N_26906,N_21722);
nand U39285 (N_39285,N_26010,N_27304);
nand U39286 (N_39286,N_20763,N_22735);
or U39287 (N_39287,N_25397,N_23910);
or U39288 (N_39288,N_21101,N_21869);
and U39289 (N_39289,N_29451,N_22195);
nor U39290 (N_39290,N_20484,N_25025);
or U39291 (N_39291,N_20231,N_20504);
nand U39292 (N_39292,N_28977,N_24587);
xnor U39293 (N_39293,N_23053,N_22529);
xnor U39294 (N_39294,N_25259,N_22656);
and U39295 (N_39295,N_20080,N_24327);
or U39296 (N_39296,N_25829,N_23027);
nor U39297 (N_39297,N_28354,N_23946);
and U39298 (N_39298,N_27783,N_23128);
or U39299 (N_39299,N_25029,N_25273);
and U39300 (N_39300,N_29361,N_25390);
and U39301 (N_39301,N_25419,N_20005);
nand U39302 (N_39302,N_26044,N_21069);
nor U39303 (N_39303,N_25036,N_22068);
and U39304 (N_39304,N_29534,N_25416);
xor U39305 (N_39305,N_25010,N_28251);
or U39306 (N_39306,N_28210,N_29653);
or U39307 (N_39307,N_24466,N_28979);
or U39308 (N_39308,N_28463,N_27188);
nand U39309 (N_39309,N_20412,N_24008);
nor U39310 (N_39310,N_27046,N_28841);
or U39311 (N_39311,N_21835,N_23610);
nand U39312 (N_39312,N_29550,N_21599);
xnor U39313 (N_39313,N_24203,N_29841);
or U39314 (N_39314,N_29316,N_20961);
and U39315 (N_39315,N_28904,N_20917);
nand U39316 (N_39316,N_20521,N_24554);
and U39317 (N_39317,N_29545,N_23347);
nor U39318 (N_39318,N_23926,N_28895);
nand U39319 (N_39319,N_22505,N_24519);
xor U39320 (N_39320,N_22480,N_20270);
and U39321 (N_39321,N_22784,N_21284);
and U39322 (N_39322,N_22348,N_28448);
and U39323 (N_39323,N_24614,N_24318);
or U39324 (N_39324,N_20277,N_23460);
nor U39325 (N_39325,N_23710,N_27320);
nor U39326 (N_39326,N_24444,N_28993);
or U39327 (N_39327,N_22583,N_21001);
nand U39328 (N_39328,N_25909,N_28564);
nor U39329 (N_39329,N_23027,N_28102);
xnor U39330 (N_39330,N_23355,N_26861);
and U39331 (N_39331,N_23782,N_22145);
and U39332 (N_39332,N_24227,N_21547);
nor U39333 (N_39333,N_29857,N_29077);
and U39334 (N_39334,N_26080,N_20413);
and U39335 (N_39335,N_24065,N_22172);
nor U39336 (N_39336,N_28978,N_29080);
and U39337 (N_39337,N_27036,N_29449);
nand U39338 (N_39338,N_29531,N_21028);
nand U39339 (N_39339,N_24848,N_27836);
and U39340 (N_39340,N_21411,N_21113);
nand U39341 (N_39341,N_23000,N_29619);
nor U39342 (N_39342,N_27665,N_25211);
nor U39343 (N_39343,N_27865,N_20870);
and U39344 (N_39344,N_25601,N_29176);
nor U39345 (N_39345,N_20397,N_21136);
and U39346 (N_39346,N_25849,N_29346);
and U39347 (N_39347,N_27937,N_27711);
and U39348 (N_39348,N_28653,N_25125);
or U39349 (N_39349,N_20289,N_24201);
or U39350 (N_39350,N_27286,N_27269);
or U39351 (N_39351,N_22631,N_27195);
nand U39352 (N_39352,N_25241,N_25787);
or U39353 (N_39353,N_24740,N_25158);
and U39354 (N_39354,N_28118,N_22082);
nor U39355 (N_39355,N_22639,N_21700);
nor U39356 (N_39356,N_20126,N_23852);
or U39357 (N_39357,N_24506,N_22907);
xnor U39358 (N_39358,N_24883,N_21077);
and U39359 (N_39359,N_25509,N_22168);
or U39360 (N_39360,N_26943,N_25501);
or U39361 (N_39361,N_22194,N_27946);
nand U39362 (N_39362,N_26651,N_22274);
nand U39363 (N_39363,N_23533,N_24459);
nand U39364 (N_39364,N_23710,N_21267);
and U39365 (N_39365,N_22133,N_24675);
and U39366 (N_39366,N_24109,N_29353);
or U39367 (N_39367,N_21620,N_21256);
and U39368 (N_39368,N_22734,N_27135);
xnor U39369 (N_39369,N_26627,N_26862);
or U39370 (N_39370,N_22241,N_20373);
nor U39371 (N_39371,N_20467,N_27219);
nor U39372 (N_39372,N_26390,N_26730);
and U39373 (N_39373,N_21059,N_24143);
and U39374 (N_39374,N_28333,N_27437);
nor U39375 (N_39375,N_29045,N_22295);
and U39376 (N_39376,N_28950,N_22106);
nor U39377 (N_39377,N_20377,N_28711);
and U39378 (N_39378,N_23783,N_20761);
nand U39379 (N_39379,N_23826,N_27746);
nand U39380 (N_39380,N_29221,N_22828);
nand U39381 (N_39381,N_29489,N_29590);
or U39382 (N_39382,N_26417,N_29361);
and U39383 (N_39383,N_24214,N_21777);
nand U39384 (N_39384,N_24928,N_23546);
xnor U39385 (N_39385,N_24493,N_20896);
nand U39386 (N_39386,N_27362,N_28603);
nor U39387 (N_39387,N_25181,N_25165);
nand U39388 (N_39388,N_20930,N_22288);
nor U39389 (N_39389,N_23199,N_23469);
xor U39390 (N_39390,N_26062,N_21959);
nor U39391 (N_39391,N_20817,N_28975);
nand U39392 (N_39392,N_24767,N_24348);
and U39393 (N_39393,N_26555,N_22553);
and U39394 (N_39394,N_20474,N_21137);
and U39395 (N_39395,N_21439,N_26812);
nand U39396 (N_39396,N_23008,N_21603);
nand U39397 (N_39397,N_23689,N_26871);
or U39398 (N_39398,N_21036,N_24341);
nor U39399 (N_39399,N_28478,N_26259);
nor U39400 (N_39400,N_20450,N_27162);
and U39401 (N_39401,N_26899,N_22400);
or U39402 (N_39402,N_22190,N_27546);
nor U39403 (N_39403,N_22452,N_28886);
xnor U39404 (N_39404,N_27336,N_28733);
nor U39405 (N_39405,N_29088,N_28192);
and U39406 (N_39406,N_29055,N_28152);
nand U39407 (N_39407,N_22839,N_28537);
nand U39408 (N_39408,N_27257,N_29126);
nor U39409 (N_39409,N_21613,N_21475);
nand U39410 (N_39410,N_23560,N_29414);
or U39411 (N_39411,N_27581,N_25350);
or U39412 (N_39412,N_25811,N_27657);
and U39413 (N_39413,N_29403,N_23366);
and U39414 (N_39414,N_26803,N_27559);
and U39415 (N_39415,N_29476,N_22055);
nand U39416 (N_39416,N_24666,N_29510);
nand U39417 (N_39417,N_23503,N_24133);
nand U39418 (N_39418,N_23837,N_25780);
nor U39419 (N_39419,N_26507,N_25761);
and U39420 (N_39420,N_24926,N_24803);
or U39421 (N_39421,N_20237,N_25691);
nor U39422 (N_39422,N_26715,N_29063);
nand U39423 (N_39423,N_22663,N_28249);
or U39424 (N_39424,N_22254,N_24101);
xnor U39425 (N_39425,N_28184,N_24414);
or U39426 (N_39426,N_28703,N_26315);
and U39427 (N_39427,N_23554,N_21077);
nor U39428 (N_39428,N_23451,N_22242);
or U39429 (N_39429,N_27363,N_20960);
and U39430 (N_39430,N_26698,N_25012);
nand U39431 (N_39431,N_28074,N_23130);
xnor U39432 (N_39432,N_20467,N_29385);
or U39433 (N_39433,N_26915,N_22916);
or U39434 (N_39434,N_25396,N_25831);
nor U39435 (N_39435,N_21678,N_29354);
or U39436 (N_39436,N_22111,N_20242);
or U39437 (N_39437,N_20640,N_21921);
nand U39438 (N_39438,N_28011,N_24956);
nor U39439 (N_39439,N_22351,N_21042);
nand U39440 (N_39440,N_28661,N_26202);
xnor U39441 (N_39441,N_27490,N_29857);
nand U39442 (N_39442,N_26576,N_23146);
nand U39443 (N_39443,N_21279,N_27169);
nand U39444 (N_39444,N_21646,N_28647);
nor U39445 (N_39445,N_22527,N_28881);
or U39446 (N_39446,N_24527,N_25534);
and U39447 (N_39447,N_28567,N_20768);
nand U39448 (N_39448,N_26555,N_23443);
xnor U39449 (N_39449,N_28467,N_28497);
nor U39450 (N_39450,N_21815,N_22100);
nor U39451 (N_39451,N_26103,N_20701);
nand U39452 (N_39452,N_25956,N_23989);
or U39453 (N_39453,N_29607,N_27405);
or U39454 (N_39454,N_26038,N_20639);
nand U39455 (N_39455,N_26050,N_25862);
or U39456 (N_39456,N_21490,N_23389);
and U39457 (N_39457,N_23854,N_26799);
nor U39458 (N_39458,N_24837,N_28313);
and U39459 (N_39459,N_23083,N_24763);
and U39460 (N_39460,N_27103,N_25405);
xnor U39461 (N_39461,N_28106,N_26882);
and U39462 (N_39462,N_23725,N_24769);
nand U39463 (N_39463,N_29435,N_23833);
and U39464 (N_39464,N_26672,N_27152);
nor U39465 (N_39465,N_26112,N_22641);
nor U39466 (N_39466,N_20975,N_24709);
nand U39467 (N_39467,N_20211,N_23732);
nand U39468 (N_39468,N_26473,N_26678);
nand U39469 (N_39469,N_24770,N_29043);
and U39470 (N_39470,N_26257,N_29295);
and U39471 (N_39471,N_23670,N_22580);
nand U39472 (N_39472,N_22267,N_29984);
nand U39473 (N_39473,N_21324,N_21608);
nor U39474 (N_39474,N_24531,N_26434);
nor U39475 (N_39475,N_27211,N_20447);
nand U39476 (N_39476,N_24339,N_20958);
nand U39477 (N_39477,N_21197,N_25810);
or U39478 (N_39478,N_21468,N_21049);
and U39479 (N_39479,N_28639,N_25690);
nand U39480 (N_39480,N_23804,N_22292);
or U39481 (N_39481,N_20070,N_28232);
and U39482 (N_39482,N_21741,N_24838);
xor U39483 (N_39483,N_23435,N_27437);
and U39484 (N_39484,N_29226,N_23507);
and U39485 (N_39485,N_26911,N_23973);
or U39486 (N_39486,N_21072,N_28275);
or U39487 (N_39487,N_27538,N_28140);
nand U39488 (N_39488,N_29031,N_23277);
nand U39489 (N_39489,N_27957,N_29479);
and U39490 (N_39490,N_22018,N_28487);
nand U39491 (N_39491,N_23144,N_22322);
or U39492 (N_39492,N_23136,N_22223);
nor U39493 (N_39493,N_27165,N_22820);
and U39494 (N_39494,N_21005,N_22864);
nor U39495 (N_39495,N_24026,N_24185);
or U39496 (N_39496,N_25043,N_28571);
nand U39497 (N_39497,N_22894,N_25487);
and U39498 (N_39498,N_24649,N_23386);
nor U39499 (N_39499,N_27014,N_20321);
nand U39500 (N_39500,N_20558,N_29563);
and U39501 (N_39501,N_21924,N_25479);
nor U39502 (N_39502,N_23818,N_29383);
nor U39503 (N_39503,N_27792,N_23997);
nor U39504 (N_39504,N_26911,N_28943);
and U39505 (N_39505,N_22999,N_20843);
or U39506 (N_39506,N_29055,N_23115);
or U39507 (N_39507,N_22696,N_27948);
xor U39508 (N_39508,N_27260,N_28117);
and U39509 (N_39509,N_22741,N_21201);
and U39510 (N_39510,N_24448,N_27156);
nor U39511 (N_39511,N_29692,N_22334);
and U39512 (N_39512,N_25792,N_24937);
nand U39513 (N_39513,N_20616,N_22696);
and U39514 (N_39514,N_20101,N_21192);
nand U39515 (N_39515,N_21934,N_27285);
nor U39516 (N_39516,N_25617,N_29623);
and U39517 (N_39517,N_28960,N_23920);
xnor U39518 (N_39518,N_25667,N_28045);
nand U39519 (N_39519,N_24467,N_24625);
and U39520 (N_39520,N_22193,N_20875);
nand U39521 (N_39521,N_27937,N_24902);
xor U39522 (N_39522,N_25661,N_23896);
and U39523 (N_39523,N_25557,N_22591);
nor U39524 (N_39524,N_24125,N_29247);
and U39525 (N_39525,N_28167,N_23270);
nor U39526 (N_39526,N_27778,N_21343);
or U39527 (N_39527,N_25515,N_23952);
nand U39528 (N_39528,N_24051,N_27804);
and U39529 (N_39529,N_28410,N_22443);
nand U39530 (N_39530,N_23890,N_23337);
nand U39531 (N_39531,N_21841,N_25252);
or U39532 (N_39532,N_23994,N_29746);
nand U39533 (N_39533,N_20135,N_27635);
nor U39534 (N_39534,N_24137,N_23194);
xnor U39535 (N_39535,N_25978,N_25095);
or U39536 (N_39536,N_28234,N_29749);
nand U39537 (N_39537,N_23027,N_22243);
nor U39538 (N_39538,N_29857,N_23800);
nor U39539 (N_39539,N_23153,N_26540);
nor U39540 (N_39540,N_29523,N_29769);
or U39541 (N_39541,N_29562,N_25431);
or U39542 (N_39542,N_28935,N_24117);
nor U39543 (N_39543,N_29021,N_22322);
nor U39544 (N_39544,N_23534,N_20913);
nand U39545 (N_39545,N_28310,N_28077);
nor U39546 (N_39546,N_28394,N_25250);
nor U39547 (N_39547,N_29326,N_24564);
or U39548 (N_39548,N_20366,N_24822);
and U39549 (N_39549,N_29364,N_25817);
nor U39550 (N_39550,N_21397,N_22638);
and U39551 (N_39551,N_27817,N_29911);
nor U39552 (N_39552,N_21933,N_26193);
and U39553 (N_39553,N_23843,N_20127);
nor U39554 (N_39554,N_23998,N_27412);
nand U39555 (N_39555,N_25278,N_28863);
and U39556 (N_39556,N_27204,N_20098);
and U39557 (N_39557,N_20082,N_25963);
nor U39558 (N_39558,N_25167,N_25202);
nand U39559 (N_39559,N_28952,N_29401);
or U39560 (N_39560,N_27982,N_26523);
nor U39561 (N_39561,N_27103,N_23693);
xor U39562 (N_39562,N_25226,N_23607);
nand U39563 (N_39563,N_29078,N_27080);
nand U39564 (N_39564,N_22600,N_22556);
xnor U39565 (N_39565,N_29693,N_29507);
and U39566 (N_39566,N_20497,N_28894);
and U39567 (N_39567,N_24518,N_21291);
nor U39568 (N_39568,N_27344,N_23530);
nand U39569 (N_39569,N_29653,N_23938);
and U39570 (N_39570,N_26471,N_26257);
nand U39571 (N_39571,N_23705,N_28584);
and U39572 (N_39572,N_25807,N_25061);
and U39573 (N_39573,N_23031,N_23421);
and U39574 (N_39574,N_21671,N_21263);
nor U39575 (N_39575,N_27224,N_29990);
or U39576 (N_39576,N_24713,N_25396);
nor U39577 (N_39577,N_25147,N_28284);
nand U39578 (N_39578,N_25236,N_25941);
and U39579 (N_39579,N_23794,N_28427);
nand U39580 (N_39580,N_21852,N_21305);
nor U39581 (N_39581,N_24237,N_25402);
or U39582 (N_39582,N_27225,N_29471);
nor U39583 (N_39583,N_23121,N_22120);
xor U39584 (N_39584,N_21645,N_27279);
or U39585 (N_39585,N_25286,N_23076);
or U39586 (N_39586,N_25062,N_21221);
or U39587 (N_39587,N_25458,N_26033);
nor U39588 (N_39588,N_21966,N_27359);
nand U39589 (N_39589,N_21640,N_21745);
nor U39590 (N_39590,N_24383,N_24775);
nor U39591 (N_39591,N_27103,N_21047);
and U39592 (N_39592,N_26370,N_26295);
xor U39593 (N_39593,N_22821,N_28994);
and U39594 (N_39594,N_23199,N_29504);
or U39595 (N_39595,N_28412,N_22428);
or U39596 (N_39596,N_27243,N_20217);
nor U39597 (N_39597,N_25356,N_28307);
nand U39598 (N_39598,N_28550,N_26875);
nand U39599 (N_39599,N_25734,N_26727);
and U39600 (N_39600,N_22284,N_25535);
xnor U39601 (N_39601,N_20322,N_25587);
or U39602 (N_39602,N_25969,N_25590);
and U39603 (N_39603,N_28965,N_28018);
or U39604 (N_39604,N_27077,N_26264);
nor U39605 (N_39605,N_28751,N_25999);
nand U39606 (N_39606,N_21695,N_20372);
nor U39607 (N_39607,N_25121,N_23960);
xnor U39608 (N_39608,N_24401,N_26050);
and U39609 (N_39609,N_22109,N_25581);
nor U39610 (N_39610,N_22812,N_22958);
and U39611 (N_39611,N_21659,N_23565);
and U39612 (N_39612,N_27787,N_20134);
and U39613 (N_39613,N_23967,N_29540);
or U39614 (N_39614,N_24078,N_20344);
and U39615 (N_39615,N_29023,N_25405);
nor U39616 (N_39616,N_22399,N_20488);
nand U39617 (N_39617,N_27748,N_23135);
and U39618 (N_39618,N_26570,N_26925);
or U39619 (N_39619,N_28800,N_23303);
nor U39620 (N_39620,N_23326,N_28815);
xnor U39621 (N_39621,N_29299,N_20649);
nand U39622 (N_39622,N_28583,N_27034);
or U39623 (N_39623,N_20301,N_23900);
and U39624 (N_39624,N_23060,N_23588);
xor U39625 (N_39625,N_26820,N_20017);
xor U39626 (N_39626,N_21158,N_27613);
nand U39627 (N_39627,N_26994,N_24161);
nand U39628 (N_39628,N_26280,N_22093);
nor U39629 (N_39629,N_25195,N_29658);
nor U39630 (N_39630,N_24280,N_27283);
or U39631 (N_39631,N_29310,N_26624);
and U39632 (N_39632,N_25264,N_21419);
and U39633 (N_39633,N_22752,N_22831);
or U39634 (N_39634,N_21238,N_20287);
xor U39635 (N_39635,N_26911,N_28028);
and U39636 (N_39636,N_22738,N_26551);
nand U39637 (N_39637,N_28632,N_24167);
nor U39638 (N_39638,N_29267,N_20711);
and U39639 (N_39639,N_26400,N_24284);
xor U39640 (N_39640,N_28819,N_20995);
or U39641 (N_39641,N_22995,N_28453);
nor U39642 (N_39642,N_22227,N_22297);
and U39643 (N_39643,N_26839,N_25275);
or U39644 (N_39644,N_20650,N_24196);
nand U39645 (N_39645,N_20923,N_26032);
xor U39646 (N_39646,N_22197,N_25551);
or U39647 (N_39647,N_26599,N_24658);
and U39648 (N_39648,N_20252,N_25453);
and U39649 (N_39649,N_22763,N_21098);
nand U39650 (N_39650,N_23083,N_26629);
xor U39651 (N_39651,N_21042,N_26259);
nand U39652 (N_39652,N_22993,N_29996);
xnor U39653 (N_39653,N_28119,N_24581);
xnor U39654 (N_39654,N_27023,N_28607);
xnor U39655 (N_39655,N_25376,N_27678);
nand U39656 (N_39656,N_20714,N_21705);
and U39657 (N_39657,N_26804,N_28316);
and U39658 (N_39658,N_29220,N_29025);
nor U39659 (N_39659,N_29413,N_29455);
nand U39660 (N_39660,N_24955,N_24263);
xnor U39661 (N_39661,N_26855,N_28573);
nand U39662 (N_39662,N_20213,N_29939);
nor U39663 (N_39663,N_21386,N_27912);
and U39664 (N_39664,N_23622,N_27992);
and U39665 (N_39665,N_27353,N_26126);
nor U39666 (N_39666,N_27725,N_24809);
nand U39667 (N_39667,N_29160,N_21660);
and U39668 (N_39668,N_23834,N_26813);
or U39669 (N_39669,N_24301,N_26465);
nand U39670 (N_39670,N_23630,N_25789);
or U39671 (N_39671,N_26530,N_29074);
nand U39672 (N_39672,N_24993,N_25689);
xnor U39673 (N_39673,N_20308,N_27950);
or U39674 (N_39674,N_23217,N_23468);
or U39675 (N_39675,N_27602,N_20202);
and U39676 (N_39676,N_20436,N_20744);
and U39677 (N_39677,N_23599,N_26136);
and U39678 (N_39678,N_20236,N_21900);
nand U39679 (N_39679,N_29926,N_26421);
and U39680 (N_39680,N_21137,N_23628);
and U39681 (N_39681,N_26113,N_26244);
and U39682 (N_39682,N_22857,N_21967);
nor U39683 (N_39683,N_25036,N_29681);
nand U39684 (N_39684,N_22027,N_20835);
nand U39685 (N_39685,N_24814,N_20309);
or U39686 (N_39686,N_28335,N_21962);
or U39687 (N_39687,N_20748,N_23926);
nor U39688 (N_39688,N_22599,N_29289);
and U39689 (N_39689,N_29627,N_28789);
nor U39690 (N_39690,N_21149,N_28619);
nor U39691 (N_39691,N_29127,N_25784);
and U39692 (N_39692,N_24134,N_21463);
nand U39693 (N_39693,N_23712,N_25782);
or U39694 (N_39694,N_23327,N_24815);
and U39695 (N_39695,N_27275,N_20829);
xor U39696 (N_39696,N_24379,N_20422);
nor U39697 (N_39697,N_22790,N_25253);
nor U39698 (N_39698,N_28705,N_27365);
xor U39699 (N_39699,N_22496,N_24613);
xnor U39700 (N_39700,N_24148,N_27229);
nand U39701 (N_39701,N_27269,N_29880);
xor U39702 (N_39702,N_20453,N_25651);
nand U39703 (N_39703,N_29524,N_25915);
and U39704 (N_39704,N_28508,N_25515);
nor U39705 (N_39705,N_27610,N_25312);
and U39706 (N_39706,N_26945,N_22128);
nand U39707 (N_39707,N_21759,N_20798);
nand U39708 (N_39708,N_25855,N_25517);
and U39709 (N_39709,N_26299,N_28701);
or U39710 (N_39710,N_22120,N_22661);
or U39711 (N_39711,N_25125,N_23215);
or U39712 (N_39712,N_22536,N_23201);
or U39713 (N_39713,N_21415,N_20582);
and U39714 (N_39714,N_25614,N_26339);
xor U39715 (N_39715,N_21199,N_25212);
or U39716 (N_39716,N_23838,N_29137);
or U39717 (N_39717,N_21222,N_29627);
xnor U39718 (N_39718,N_23591,N_21417);
nor U39719 (N_39719,N_27470,N_23887);
nand U39720 (N_39720,N_20051,N_25971);
and U39721 (N_39721,N_21792,N_29964);
nand U39722 (N_39722,N_25021,N_26930);
nand U39723 (N_39723,N_28702,N_22082);
nor U39724 (N_39724,N_27395,N_27282);
xor U39725 (N_39725,N_23047,N_24323);
xor U39726 (N_39726,N_27112,N_20252);
nand U39727 (N_39727,N_20728,N_26349);
or U39728 (N_39728,N_22689,N_29238);
and U39729 (N_39729,N_23880,N_26223);
nand U39730 (N_39730,N_25248,N_27173);
and U39731 (N_39731,N_28286,N_20823);
and U39732 (N_39732,N_25085,N_20999);
and U39733 (N_39733,N_20485,N_22248);
or U39734 (N_39734,N_22587,N_29849);
and U39735 (N_39735,N_23427,N_24294);
nor U39736 (N_39736,N_25728,N_23100);
xnor U39737 (N_39737,N_25114,N_22328);
xor U39738 (N_39738,N_27192,N_21770);
or U39739 (N_39739,N_25667,N_22122);
or U39740 (N_39740,N_23037,N_21227);
and U39741 (N_39741,N_23816,N_22331);
and U39742 (N_39742,N_28784,N_28435);
or U39743 (N_39743,N_21814,N_28010);
nor U39744 (N_39744,N_27099,N_29971);
nand U39745 (N_39745,N_28242,N_20274);
nor U39746 (N_39746,N_21647,N_26576);
nor U39747 (N_39747,N_25386,N_26616);
nor U39748 (N_39748,N_22006,N_25270);
and U39749 (N_39749,N_24281,N_28730);
or U39750 (N_39750,N_27368,N_22353);
xnor U39751 (N_39751,N_22842,N_29499);
xnor U39752 (N_39752,N_21754,N_28592);
nand U39753 (N_39753,N_27409,N_27073);
nand U39754 (N_39754,N_22808,N_23678);
nand U39755 (N_39755,N_23592,N_25133);
or U39756 (N_39756,N_24720,N_29445);
or U39757 (N_39757,N_23900,N_24234);
or U39758 (N_39758,N_24043,N_25844);
nand U39759 (N_39759,N_20294,N_27283);
and U39760 (N_39760,N_28569,N_26906);
nand U39761 (N_39761,N_21378,N_29434);
or U39762 (N_39762,N_21912,N_28483);
nand U39763 (N_39763,N_28260,N_20385);
or U39764 (N_39764,N_24273,N_22631);
nand U39765 (N_39765,N_28074,N_29508);
nand U39766 (N_39766,N_28295,N_24125);
nand U39767 (N_39767,N_22807,N_20863);
and U39768 (N_39768,N_28391,N_24057);
and U39769 (N_39769,N_20865,N_20002);
or U39770 (N_39770,N_22601,N_27013);
nand U39771 (N_39771,N_22945,N_24071);
nand U39772 (N_39772,N_23634,N_26608);
nor U39773 (N_39773,N_21971,N_28632);
or U39774 (N_39774,N_24359,N_28086);
and U39775 (N_39775,N_22640,N_23720);
nor U39776 (N_39776,N_27582,N_25480);
nor U39777 (N_39777,N_23582,N_26165);
or U39778 (N_39778,N_24511,N_28869);
or U39779 (N_39779,N_21920,N_24137);
and U39780 (N_39780,N_27791,N_23656);
xor U39781 (N_39781,N_21791,N_26784);
nand U39782 (N_39782,N_29390,N_23651);
and U39783 (N_39783,N_22196,N_21817);
nand U39784 (N_39784,N_24065,N_24111);
or U39785 (N_39785,N_29856,N_29277);
nand U39786 (N_39786,N_28427,N_22921);
or U39787 (N_39787,N_25557,N_22140);
xor U39788 (N_39788,N_23821,N_22633);
nor U39789 (N_39789,N_24434,N_20817);
or U39790 (N_39790,N_25781,N_20041);
or U39791 (N_39791,N_25491,N_24069);
and U39792 (N_39792,N_28615,N_20937);
nand U39793 (N_39793,N_24631,N_29243);
or U39794 (N_39794,N_28394,N_29746);
nor U39795 (N_39795,N_27143,N_20000);
or U39796 (N_39796,N_26041,N_20295);
nand U39797 (N_39797,N_25476,N_28271);
nand U39798 (N_39798,N_23109,N_24306);
and U39799 (N_39799,N_24270,N_25313);
and U39800 (N_39800,N_29829,N_20635);
or U39801 (N_39801,N_29966,N_22345);
or U39802 (N_39802,N_27386,N_23618);
nand U39803 (N_39803,N_27635,N_29131);
nor U39804 (N_39804,N_26481,N_28769);
nor U39805 (N_39805,N_21980,N_26775);
and U39806 (N_39806,N_22231,N_24217);
or U39807 (N_39807,N_27058,N_23832);
and U39808 (N_39808,N_23207,N_25243);
and U39809 (N_39809,N_21434,N_24798);
and U39810 (N_39810,N_25999,N_20209);
and U39811 (N_39811,N_25474,N_22480);
and U39812 (N_39812,N_28469,N_21067);
nor U39813 (N_39813,N_28366,N_24539);
or U39814 (N_39814,N_29451,N_20054);
and U39815 (N_39815,N_25806,N_21506);
xnor U39816 (N_39816,N_24883,N_24878);
nor U39817 (N_39817,N_22788,N_26212);
nor U39818 (N_39818,N_21864,N_27104);
or U39819 (N_39819,N_22112,N_29751);
or U39820 (N_39820,N_28377,N_26360);
or U39821 (N_39821,N_25191,N_24121);
nor U39822 (N_39822,N_28316,N_24757);
nand U39823 (N_39823,N_20221,N_26319);
nor U39824 (N_39824,N_20377,N_29379);
or U39825 (N_39825,N_29069,N_27236);
nor U39826 (N_39826,N_23192,N_21905);
or U39827 (N_39827,N_21039,N_27952);
or U39828 (N_39828,N_20602,N_21503);
nand U39829 (N_39829,N_24649,N_27559);
nor U39830 (N_39830,N_23701,N_21486);
and U39831 (N_39831,N_23349,N_26986);
or U39832 (N_39832,N_22996,N_22724);
xor U39833 (N_39833,N_23310,N_26437);
nand U39834 (N_39834,N_22043,N_27881);
or U39835 (N_39835,N_27440,N_20500);
xor U39836 (N_39836,N_25745,N_29987);
and U39837 (N_39837,N_27580,N_26174);
and U39838 (N_39838,N_20378,N_23362);
and U39839 (N_39839,N_24283,N_21185);
or U39840 (N_39840,N_27383,N_29842);
or U39841 (N_39841,N_23246,N_28795);
and U39842 (N_39842,N_26886,N_23651);
or U39843 (N_39843,N_29900,N_29157);
and U39844 (N_39844,N_26931,N_23126);
nand U39845 (N_39845,N_24990,N_23810);
and U39846 (N_39846,N_24701,N_20923);
and U39847 (N_39847,N_29451,N_20479);
xor U39848 (N_39848,N_22642,N_29879);
and U39849 (N_39849,N_20976,N_20687);
or U39850 (N_39850,N_22493,N_22343);
nor U39851 (N_39851,N_24692,N_20274);
and U39852 (N_39852,N_25208,N_28626);
xnor U39853 (N_39853,N_20146,N_21115);
or U39854 (N_39854,N_27075,N_22327);
nor U39855 (N_39855,N_27977,N_27103);
and U39856 (N_39856,N_21375,N_29270);
nand U39857 (N_39857,N_21393,N_25876);
or U39858 (N_39858,N_28590,N_26462);
nand U39859 (N_39859,N_25978,N_23254);
xor U39860 (N_39860,N_25480,N_23747);
nand U39861 (N_39861,N_23973,N_28220);
nand U39862 (N_39862,N_22478,N_29910);
nand U39863 (N_39863,N_22997,N_27768);
nor U39864 (N_39864,N_26777,N_22216);
xor U39865 (N_39865,N_23599,N_20069);
or U39866 (N_39866,N_26252,N_29605);
nor U39867 (N_39867,N_28413,N_21621);
nor U39868 (N_39868,N_24436,N_24123);
and U39869 (N_39869,N_26421,N_21471);
nand U39870 (N_39870,N_28281,N_28079);
nand U39871 (N_39871,N_24527,N_28494);
nand U39872 (N_39872,N_21423,N_27138);
or U39873 (N_39873,N_25758,N_23578);
and U39874 (N_39874,N_23185,N_28657);
xnor U39875 (N_39875,N_27020,N_28787);
nor U39876 (N_39876,N_28353,N_21142);
or U39877 (N_39877,N_24796,N_29825);
and U39878 (N_39878,N_24796,N_29835);
nor U39879 (N_39879,N_26616,N_25709);
or U39880 (N_39880,N_24596,N_22082);
and U39881 (N_39881,N_27584,N_27616);
or U39882 (N_39882,N_28348,N_24673);
nor U39883 (N_39883,N_27562,N_28303);
nand U39884 (N_39884,N_22913,N_22624);
or U39885 (N_39885,N_22526,N_28882);
and U39886 (N_39886,N_22031,N_27774);
or U39887 (N_39887,N_29914,N_29525);
nand U39888 (N_39888,N_24313,N_25363);
or U39889 (N_39889,N_26313,N_26079);
nor U39890 (N_39890,N_24785,N_23692);
and U39891 (N_39891,N_26417,N_27144);
and U39892 (N_39892,N_26002,N_27994);
nand U39893 (N_39893,N_28111,N_20871);
xnor U39894 (N_39894,N_29102,N_25742);
or U39895 (N_39895,N_22337,N_24282);
nor U39896 (N_39896,N_24466,N_24395);
and U39897 (N_39897,N_21743,N_27574);
nand U39898 (N_39898,N_27176,N_28061);
nand U39899 (N_39899,N_24927,N_29369);
and U39900 (N_39900,N_20993,N_24339);
nor U39901 (N_39901,N_24535,N_25772);
nor U39902 (N_39902,N_21787,N_24175);
nand U39903 (N_39903,N_22731,N_21026);
nand U39904 (N_39904,N_20583,N_22200);
nand U39905 (N_39905,N_26417,N_26985);
nor U39906 (N_39906,N_22169,N_24070);
nor U39907 (N_39907,N_21923,N_29145);
nor U39908 (N_39908,N_24826,N_29667);
xor U39909 (N_39909,N_21770,N_25634);
xnor U39910 (N_39910,N_25153,N_20564);
and U39911 (N_39911,N_23560,N_20892);
nor U39912 (N_39912,N_20570,N_23460);
and U39913 (N_39913,N_21898,N_21928);
or U39914 (N_39914,N_23984,N_21043);
xnor U39915 (N_39915,N_27060,N_28505);
xor U39916 (N_39916,N_23379,N_26909);
xor U39917 (N_39917,N_24583,N_29699);
nand U39918 (N_39918,N_24774,N_29569);
nor U39919 (N_39919,N_28725,N_25703);
or U39920 (N_39920,N_24572,N_26456);
or U39921 (N_39921,N_25921,N_27685);
xor U39922 (N_39922,N_29972,N_22643);
nand U39923 (N_39923,N_22255,N_28084);
and U39924 (N_39924,N_27393,N_22661);
nor U39925 (N_39925,N_24274,N_24379);
nor U39926 (N_39926,N_28000,N_20802);
xnor U39927 (N_39927,N_22771,N_22676);
nor U39928 (N_39928,N_27721,N_22987);
or U39929 (N_39929,N_23212,N_22116);
and U39930 (N_39930,N_23262,N_21026);
or U39931 (N_39931,N_27602,N_29039);
and U39932 (N_39932,N_22090,N_28021);
or U39933 (N_39933,N_20217,N_28618);
nand U39934 (N_39934,N_29164,N_23864);
or U39935 (N_39935,N_25698,N_26791);
xor U39936 (N_39936,N_26404,N_25986);
or U39937 (N_39937,N_22651,N_28793);
or U39938 (N_39938,N_27514,N_28109);
and U39939 (N_39939,N_27249,N_23684);
xnor U39940 (N_39940,N_25246,N_26988);
nand U39941 (N_39941,N_27868,N_22545);
or U39942 (N_39942,N_22047,N_27118);
and U39943 (N_39943,N_24934,N_21748);
nand U39944 (N_39944,N_28726,N_23154);
nor U39945 (N_39945,N_20170,N_21296);
nand U39946 (N_39946,N_21146,N_21509);
nand U39947 (N_39947,N_22195,N_26598);
nor U39948 (N_39948,N_22468,N_29414);
and U39949 (N_39949,N_23955,N_23882);
nand U39950 (N_39950,N_24652,N_22697);
nor U39951 (N_39951,N_22895,N_26797);
nor U39952 (N_39952,N_20473,N_25280);
or U39953 (N_39953,N_22997,N_22729);
or U39954 (N_39954,N_27955,N_24072);
nor U39955 (N_39955,N_28456,N_29794);
and U39956 (N_39956,N_20606,N_20378);
xor U39957 (N_39957,N_21576,N_24660);
xnor U39958 (N_39958,N_28913,N_24533);
xor U39959 (N_39959,N_22182,N_27258);
nor U39960 (N_39960,N_20385,N_28116);
nand U39961 (N_39961,N_29117,N_24846);
or U39962 (N_39962,N_27706,N_27234);
nor U39963 (N_39963,N_20898,N_22116);
nor U39964 (N_39964,N_28338,N_21098);
or U39965 (N_39965,N_24511,N_29533);
nand U39966 (N_39966,N_21374,N_26922);
nor U39967 (N_39967,N_26958,N_28828);
and U39968 (N_39968,N_22399,N_24338);
nand U39969 (N_39969,N_23698,N_21635);
or U39970 (N_39970,N_25601,N_29656);
nand U39971 (N_39971,N_27905,N_24174);
or U39972 (N_39972,N_22308,N_27338);
nor U39973 (N_39973,N_27994,N_22005);
nand U39974 (N_39974,N_20977,N_26594);
and U39975 (N_39975,N_25705,N_22845);
nor U39976 (N_39976,N_23603,N_25967);
or U39977 (N_39977,N_26192,N_22786);
nand U39978 (N_39978,N_22246,N_28165);
nand U39979 (N_39979,N_20770,N_26881);
nand U39980 (N_39980,N_21681,N_23018);
and U39981 (N_39981,N_22046,N_27862);
nand U39982 (N_39982,N_22125,N_22738);
xnor U39983 (N_39983,N_26007,N_20183);
nand U39984 (N_39984,N_24353,N_28484);
and U39985 (N_39985,N_23494,N_27407);
and U39986 (N_39986,N_21778,N_23441);
and U39987 (N_39987,N_20045,N_21595);
nor U39988 (N_39988,N_22518,N_29717);
nor U39989 (N_39989,N_21139,N_25319);
or U39990 (N_39990,N_22556,N_25768);
nand U39991 (N_39991,N_23179,N_25882);
or U39992 (N_39992,N_22399,N_24026);
and U39993 (N_39993,N_22927,N_23156);
or U39994 (N_39994,N_25839,N_25139);
and U39995 (N_39995,N_20535,N_24759);
and U39996 (N_39996,N_28534,N_20040);
or U39997 (N_39997,N_20465,N_23917);
and U39998 (N_39998,N_24561,N_28864);
or U39999 (N_39999,N_29834,N_24720);
or U40000 (N_40000,N_37236,N_35282);
nor U40001 (N_40001,N_36956,N_36850);
or U40002 (N_40002,N_35841,N_32613);
and U40003 (N_40003,N_36380,N_35740);
xor U40004 (N_40004,N_32575,N_37795);
nor U40005 (N_40005,N_35175,N_33474);
nand U40006 (N_40006,N_33041,N_35207);
or U40007 (N_40007,N_34336,N_35732);
nor U40008 (N_40008,N_39975,N_36487);
and U40009 (N_40009,N_31020,N_35191);
and U40010 (N_40010,N_39938,N_38684);
nand U40011 (N_40011,N_35601,N_30228);
and U40012 (N_40012,N_31828,N_36526);
or U40013 (N_40013,N_31890,N_34128);
and U40014 (N_40014,N_38709,N_31369);
nand U40015 (N_40015,N_31069,N_30368);
and U40016 (N_40016,N_38848,N_32121);
nand U40017 (N_40017,N_35170,N_37925);
nor U40018 (N_40018,N_37093,N_32397);
nor U40019 (N_40019,N_34760,N_36915);
nor U40020 (N_40020,N_36537,N_32873);
nand U40021 (N_40021,N_31200,N_38063);
or U40022 (N_40022,N_34926,N_30338);
or U40023 (N_40023,N_37623,N_33222);
nor U40024 (N_40024,N_36872,N_31303);
xnor U40025 (N_40025,N_35986,N_35677);
or U40026 (N_40026,N_33544,N_33977);
nor U40027 (N_40027,N_38564,N_31634);
and U40028 (N_40028,N_35747,N_34259);
nand U40029 (N_40029,N_31547,N_37940);
nand U40030 (N_40030,N_34087,N_39231);
xnor U40031 (N_40031,N_36221,N_33175);
and U40032 (N_40032,N_37143,N_34764);
nand U40033 (N_40033,N_31745,N_32724);
and U40034 (N_40034,N_33065,N_34110);
nand U40035 (N_40035,N_32094,N_39080);
and U40036 (N_40036,N_36509,N_35178);
nor U40037 (N_40037,N_34670,N_34955);
nand U40038 (N_40038,N_36722,N_36196);
or U40039 (N_40039,N_37352,N_33697);
nand U40040 (N_40040,N_36703,N_30035);
nor U40041 (N_40041,N_37163,N_33213);
xor U40042 (N_40042,N_39304,N_34474);
nand U40043 (N_40043,N_35704,N_39131);
or U40044 (N_40044,N_30537,N_33081);
nand U40045 (N_40045,N_32493,N_38783);
nor U40046 (N_40046,N_33138,N_30987);
and U40047 (N_40047,N_36372,N_30682);
nand U40048 (N_40048,N_35706,N_32100);
nor U40049 (N_40049,N_33567,N_36906);
nor U40050 (N_40050,N_34732,N_30425);
xor U40051 (N_40051,N_32599,N_36449);
xnor U40052 (N_40052,N_30939,N_35298);
and U40053 (N_40053,N_37456,N_35654);
nor U40054 (N_40054,N_38475,N_31009);
and U40055 (N_40055,N_36826,N_39682);
or U40056 (N_40056,N_34473,N_32438);
or U40057 (N_40057,N_32770,N_31687);
and U40058 (N_40058,N_34248,N_39618);
and U40059 (N_40059,N_35711,N_33617);
nand U40060 (N_40060,N_31114,N_30599);
nand U40061 (N_40061,N_34215,N_30762);
or U40062 (N_40062,N_35818,N_38342);
xor U40063 (N_40063,N_35355,N_31161);
or U40064 (N_40064,N_34075,N_32719);
or U40065 (N_40065,N_37274,N_38593);
and U40066 (N_40066,N_37265,N_39768);
nand U40067 (N_40067,N_35213,N_34465);
nor U40068 (N_40068,N_38289,N_36338);
nand U40069 (N_40069,N_31696,N_33683);
and U40070 (N_40070,N_33029,N_31497);
and U40071 (N_40071,N_31544,N_31139);
nand U40072 (N_40072,N_33737,N_31414);
or U40073 (N_40073,N_30417,N_33379);
nand U40074 (N_40074,N_36486,N_35880);
or U40075 (N_40075,N_33185,N_35894);
nand U40076 (N_40076,N_35693,N_35335);
nand U40077 (N_40077,N_31300,N_39773);
or U40078 (N_40078,N_34210,N_38179);
nand U40079 (N_40079,N_31254,N_37576);
and U40080 (N_40080,N_39122,N_37651);
nor U40081 (N_40081,N_36032,N_34530);
nand U40082 (N_40082,N_30723,N_37222);
or U40083 (N_40083,N_38012,N_35583);
nor U40084 (N_40084,N_32998,N_36961);
and U40085 (N_40085,N_38944,N_35428);
nor U40086 (N_40086,N_36737,N_31130);
nand U40087 (N_40087,N_38717,N_30570);
and U40088 (N_40088,N_35200,N_35283);
nand U40089 (N_40089,N_36823,N_34535);
and U40090 (N_40090,N_30517,N_35592);
and U40091 (N_40091,N_38042,N_34296);
nand U40092 (N_40092,N_39255,N_39707);
nand U40093 (N_40093,N_39471,N_31086);
and U40094 (N_40094,N_39303,N_35966);
nand U40095 (N_40095,N_30568,N_39706);
or U40096 (N_40096,N_37323,N_39351);
nor U40097 (N_40097,N_30852,N_35668);
nand U40098 (N_40098,N_38804,N_36400);
nand U40099 (N_40099,N_35679,N_34434);
nand U40100 (N_40100,N_30298,N_30976);
or U40101 (N_40101,N_36269,N_30995);
nor U40102 (N_40102,N_34912,N_36472);
or U40103 (N_40103,N_30093,N_39008);
nor U40104 (N_40104,N_34868,N_32233);
nor U40105 (N_40105,N_34572,N_34830);
nand U40106 (N_40106,N_31673,N_38349);
xor U40107 (N_40107,N_39367,N_37114);
and U40108 (N_40108,N_33673,N_30495);
or U40109 (N_40109,N_31259,N_32628);
nand U40110 (N_40110,N_34217,N_37158);
nand U40111 (N_40111,N_34848,N_31787);
or U40112 (N_40112,N_38852,N_32024);
nand U40113 (N_40113,N_32456,N_35967);
nand U40114 (N_40114,N_39625,N_37695);
or U40115 (N_40115,N_39652,N_39261);
nor U40116 (N_40116,N_38140,N_33387);
nand U40117 (N_40117,N_39480,N_32020);
nand U40118 (N_40118,N_37641,N_32140);
and U40119 (N_40119,N_36650,N_39402);
and U40120 (N_40120,N_32072,N_38947);
and U40121 (N_40121,N_33691,N_33101);
nor U40122 (N_40122,N_30588,N_30316);
or U40123 (N_40123,N_33497,N_33324);
xnor U40124 (N_40124,N_35787,N_30240);
and U40125 (N_40125,N_38101,N_33206);
xor U40126 (N_40126,N_38863,N_37742);
or U40127 (N_40127,N_32970,N_36943);
nand U40128 (N_40128,N_33438,N_30631);
nor U40129 (N_40129,N_32127,N_38741);
or U40130 (N_40130,N_31621,N_33835);
or U40131 (N_40131,N_35936,N_35799);
nor U40132 (N_40132,N_38430,N_39044);
nor U40133 (N_40133,N_30527,N_35314);
or U40134 (N_40134,N_36191,N_33073);
or U40135 (N_40135,N_31038,N_33279);
or U40136 (N_40136,N_36974,N_33895);
nand U40137 (N_40137,N_37038,N_37135);
nor U40138 (N_40138,N_30749,N_32769);
xnor U40139 (N_40139,N_32455,N_35057);
and U40140 (N_40140,N_30810,N_30356);
xnor U40141 (N_40141,N_37823,N_33214);
nand U40142 (N_40142,N_39672,N_37108);
nor U40143 (N_40143,N_38139,N_33625);
or U40144 (N_40144,N_38644,N_30006);
nor U40145 (N_40145,N_36909,N_35297);
nand U40146 (N_40146,N_32312,N_39570);
nor U40147 (N_40147,N_36073,N_33299);
nand U40148 (N_40148,N_33086,N_30235);
and U40149 (N_40149,N_31504,N_39262);
and U40150 (N_40150,N_39776,N_31306);
and U40151 (N_40151,N_34262,N_33883);
nand U40152 (N_40152,N_39528,N_37948);
nand U40153 (N_40153,N_30451,N_33610);
nor U40154 (N_40154,N_34220,N_34792);
nor U40155 (N_40155,N_38460,N_31341);
nor U40156 (N_40156,N_33606,N_32236);
nor U40157 (N_40157,N_32508,N_39515);
nor U40158 (N_40158,N_35135,N_35387);
nor U40159 (N_40159,N_35511,N_37168);
and U40160 (N_40160,N_34849,N_30077);
nand U40161 (N_40161,N_34845,N_31597);
and U40162 (N_40162,N_32075,N_30477);
or U40163 (N_40163,N_32830,N_34659);
nand U40164 (N_40164,N_37762,N_36780);
nand U40165 (N_40165,N_36505,N_30785);
nand U40166 (N_40166,N_32945,N_33083);
nor U40167 (N_40167,N_31106,N_37834);
nor U40168 (N_40168,N_35617,N_35412);
and U40169 (N_40169,N_30410,N_30078);
or U40170 (N_40170,N_37406,N_39420);
nand U40171 (N_40171,N_35481,N_32426);
nand U40172 (N_40172,N_31162,N_37078);
and U40173 (N_40173,N_36188,N_37949);
and U40174 (N_40174,N_37976,N_38299);
xor U40175 (N_40175,N_34829,N_38890);
xnor U40176 (N_40176,N_36018,N_32570);
nand U40177 (N_40177,N_32422,N_39373);
xor U40178 (N_40178,N_33888,N_39711);
or U40179 (N_40179,N_36347,N_35225);
and U40180 (N_40180,N_30372,N_36769);
or U40181 (N_40181,N_35738,N_34023);
or U40182 (N_40182,N_30452,N_39662);
nor U40183 (N_40183,N_30775,N_30536);
nor U40184 (N_40184,N_31994,N_34208);
or U40185 (N_40185,N_39322,N_30564);
and U40186 (N_40186,N_33828,N_36718);
nand U40187 (N_40187,N_36636,N_31233);
and U40188 (N_40188,N_36848,N_37803);
nor U40189 (N_40189,N_39408,N_38596);
and U40190 (N_40190,N_31090,N_30326);
and U40191 (N_40191,N_32500,N_36839);
nor U40192 (N_40192,N_39488,N_39579);
nor U40193 (N_40193,N_37349,N_33447);
xor U40194 (N_40194,N_39530,N_38191);
nor U40195 (N_40195,N_31604,N_30166);
nor U40196 (N_40196,N_33327,N_31593);
or U40197 (N_40197,N_34286,N_37006);
nand U40198 (N_40198,N_37709,N_36896);
nand U40199 (N_40199,N_39175,N_31327);
nand U40200 (N_40200,N_38485,N_35797);
nand U40201 (N_40201,N_36484,N_37400);
or U40202 (N_40202,N_32740,N_37556);
nor U40203 (N_40203,N_32280,N_32165);
nand U40204 (N_40204,N_37788,N_33703);
nor U40205 (N_40205,N_34987,N_32179);
nand U40206 (N_40206,N_32901,N_35792);
and U40207 (N_40207,N_36433,N_35616);
and U40208 (N_40208,N_34475,N_34452);
and U40209 (N_40209,N_39417,N_36558);
xor U40210 (N_40210,N_36840,N_39018);
or U40211 (N_40211,N_30121,N_33698);
or U40212 (N_40212,N_37360,N_39872);
nor U40213 (N_40213,N_32458,N_39151);
and U40214 (N_40214,N_38665,N_34977);
nand U40215 (N_40215,N_37776,N_33509);
nor U40216 (N_40216,N_34950,N_38476);
and U40217 (N_40217,N_30698,N_34935);
or U40218 (N_40218,N_31206,N_36493);
nand U40219 (N_40219,N_37164,N_36480);
or U40220 (N_40220,N_33787,N_35536);
or U40221 (N_40221,N_34275,N_34468);
nor U40222 (N_40222,N_33847,N_37758);
and U40223 (N_40223,N_34225,N_32341);
nand U40224 (N_40224,N_30307,N_37722);
xor U40225 (N_40225,N_34925,N_39891);
and U40226 (N_40226,N_32515,N_30772);
and U40227 (N_40227,N_36868,N_30758);
nand U40228 (N_40228,N_31867,N_30855);
and U40229 (N_40229,N_35606,N_36550);
or U40230 (N_40230,N_38174,N_39961);
and U40231 (N_40231,N_38291,N_38124);
nand U40232 (N_40232,N_32904,N_39495);
nand U40233 (N_40233,N_39412,N_38834);
xnor U40234 (N_40234,N_38689,N_39095);
and U40235 (N_40235,N_38343,N_38339);
nor U40236 (N_40236,N_35430,N_38790);
xnor U40237 (N_40237,N_36330,N_38466);
nor U40238 (N_40238,N_34214,N_35913);
and U40239 (N_40239,N_31496,N_32790);
and U40240 (N_40240,N_30102,N_33619);
nand U40241 (N_40241,N_32888,N_34944);
xnor U40242 (N_40242,N_38880,N_38167);
nor U40243 (N_40243,N_39128,N_31045);
nor U40244 (N_40244,N_39270,N_38180);
nor U40245 (N_40245,N_34951,N_38334);
or U40246 (N_40246,N_38901,N_36949);
and U40247 (N_40247,N_33841,N_31026);
and U40248 (N_40248,N_34313,N_31323);
and U40249 (N_40249,N_33887,N_35538);
and U40250 (N_40250,N_38212,N_34222);
nor U40251 (N_40251,N_38626,N_37771);
or U40252 (N_40252,N_35837,N_39287);
or U40253 (N_40253,N_34138,N_37817);
nor U40254 (N_40254,N_36287,N_34709);
xnor U40255 (N_40255,N_35440,N_32818);
nor U40256 (N_40256,N_35447,N_38631);
or U40257 (N_40257,N_34633,N_34662);
and U40258 (N_40258,N_33609,N_30232);
xor U40259 (N_40259,N_32723,N_31986);
nor U40260 (N_40260,N_36797,N_35094);
nand U40261 (N_40261,N_34634,N_30611);
or U40262 (N_40262,N_30666,N_36232);
nand U40263 (N_40263,N_35071,N_38752);
nand U40264 (N_40264,N_30342,N_31008);
xor U40265 (N_40265,N_36810,N_30142);
nor U40266 (N_40266,N_32738,N_37989);
or U40267 (N_40267,N_39117,N_31070);
nand U40268 (N_40268,N_38781,N_36383);
nor U40269 (N_40269,N_37185,N_38975);
nand U40270 (N_40270,N_34741,N_36436);
xnor U40271 (N_40271,N_35338,N_30300);
and U40272 (N_40272,N_33139,N_35075);
xnor U40273 (N_40273,N_39003,N_35664);
nor U40274 (N_40274,N_32074,N_39167);
nor U40275 (N_40275,N_39669,N_34759);
or U40276 (N_40276,N_32741,N_35410);
or U40277 (N_40277,N_31579,N_30974);
nand U40278 (N_40278,N_38540,N_32835);
and U40279 (N_40279,N_36580,N_34898);
and U40280 (N_40280,N_37698,N_32731);
or U40281 (N_40281,N_32531,N_38133);
or U40282 (N_40282,N_38601,N_31326);
nor U40283 (N_40283,N_33614,N_37020);
nand U40284 (N_40284,N_38568,N_30835);
and U40285 (N_40285,N_36995,N_37263);
or U40286 (N_40286,N_38799,N_36385);
nand U40287 (N_40287,N_38578,N_38616);
or U40288 (N_40288,N_38356,N_33225);
or U40289 (N_40289,N_30849,N_39383);
xor U40290 (N_40290,N_31433,N_39400);
nand U40291 (N_40291,N_33056,N_35288);
or U40292 (N_40292,N_38019,N_38603);
or U40293 (N_40293,N_32812,N_38265);
or U40294 (N_40294,N_33098,N_30213);
nand U40295 (N_40295,N_36375,N_34098);
nand U40296 (N_40296,N_39085,N_30946);
nand U40297 (N_40297,N_38207,N_36093);
nor U40298 (N_40298,N_33232,N_37101);
or U40299 (N_40299,N_34022,N_38780);
or U40300 (N_40300,N_36306,N_30803);
nor U40301 (N_40301,N_35871,N_34334);
and U40302 (N_40302,N_30158,N_30373);
and U40303 (N_40303,N_35516,N_32160);
nor U40304 (N_40304,N_33901,N_36623);
nor U40305 (N_40305,N_39778,N_34233);
xnor U40306 (N_40306,N_31820,N_39917);
nor U40307 (N_40307,N_33329,N_36842);
and U40308 (N_40308,N_32924,N_35708);
nand U40309 (N_40309,N_35366,N_38567);
and U40310 (N_40310,N_39120,N_35650);
and U40311 (N_40311,N_39157,N_39016);
or U40312 (N_40312,N_38261,N_33253);
and U40313 (N_40313,N_37286,N_31140);
nor U40314 (N_40314,N_32197,N_34714);
and U40315 (N_40315,N_39968,N_35442);
nor U40316 (N_40316,N_39384,N_32480);
nor U40317 (N_40317,N_37598,N_38979);
and U40318 (N_40318,N_36539,N_35652);
xnor U40319 (N_40319,N_34481,N_30780);
nor U40320 (N_40320,N_36134,N_31280);
or U40321 (N_40321,N_33858,N_35567);
nand U40322 (N_40322,N_32026,N_37516);
and U40323 (N_40323,N_39661,N_35354);
and U40324 (N_40324,N_31817,N_34006);
or U40325 (N_40325,N_30934,N_37042);
and U40326 (N_40326,N_33983,N_30001);
or U40327 (N_40327,N_32796,N_32528);
and U40328 (N_40328,N_34299,N_34869);
or U40329 (N_40329,N_31612,N_31115);
nor U40330 (N_40330,N_32655,N_36286);
or U40331 (N_40331,N_39845,N_37171);
nand U40332 (N_40332,N_37443,N_39822);
and U40333 (N_40333,N_30560,N_35780);
nor U40334 (N_40334,N_32429,N_32462);
or U40335 (N_40335,N_34685,N_36272);
and U40336 (N_40336,N_32113,N_37885);
nand U40337 (N_40337,N_38130,N_30198);
nand U40338 (N_40338,N_36939,N_36897);
and U40339 (N_40339,N_30439,N_36418);
xor U40340 (N_40340,N_32168,N_36210);
and U40341 (N_40341,N_35319,N_37980);
nor U40342 (N_40342,N_31541,N_32469);
nand U40343 (N_40343,N_37990,N_36328);
nand U40344 (N_40344,N_37692,N_36146);
xor U40345 (N_40345,N_32712,N_38597);
xnor U40346 (N_40346,N_35104,N_35038);
nor U40347 (N_40347,N_37658,N_38363);
or U40348 (N_40348,N_39189,N_30246);
nor U40349 (N_40349,N_31979,N_38041);
nand U40350 (N_40350,N_30685,N_32722);
and U40351 (N_40351,N_39281,N_37860);
nor U40352 (N_40352,N_34020,N_31600);
and U40353 (N_40353,N_33357,N_34167);
nand U40354 (N_40354,N_34733,N_35590);
nand U40355 (N_40355,N_31811,N_32296);
nand U40356 (N_40356,N_38170,N_36235);
nor U40357 (N_40357,N_32365,N_38972);
nand U40358 (N_40358,N_38514,N_33174);
xnor U40359 (N_40359,N_37145,N_38321);
and U40360 (N_40360,N_39761,N_31197);
nand U40361 (N_40361,N_30182,N_36976);
nor U40362 (N_40362,N_35717,N_30947);
and U40363 (N_40363,N_33117,N_35879);
or U40364 (N_40364,N_30687,N_34990);
nand U40365 (N_40365,N_37687,N_30290);
and U40366 (N_40366,N_38016,N_36782);
nor U40367 (N_40367,N_38000,N_38410);
and U40368 (N_40368,N_33770,N_37371);
or U40369 (N_40369,N_38670,N_30136);
nor U40370 (N_40370,N_33863,N_30787);
nand U40371 (N_40371,N_32083,N_34047);
or U40372 (N_40372,N_37469,N_39110);
nor U40373 (N_40373,N_32645,N_34079);
or U40374 (N_40374,N_34024,N_36829);
or U40375 (N_40375,N_33778,N_34147);
nand U40376 (N_40376,N_38882,N_36415);
and U40377 (N_40377,N_34711,N_38753);
xor U40378 (N_40378,N_32217,N_35689);
or U40379 (N_40379,N_39007,N_34350);
and U40380 (N_40380,N_37011,N_36601);
or U40381 (N_40381,N_32816,N_35777);
xor U40382 (N_40382,N_38573,N_38402);
xnor U40383 (N_40383,N_36327,N_39240);
nand U40384 (N_40384,N_32636,N_37956);
xor U40385 (N_40385,N_31435,N_35032);
nor U40386 (N_40386,N_36204,N_32057);
and U40387 (N_40387,N_33388,N_34647);
nor U40388 (N_40388,N_37150,N_37770);
and U40389 (N_40389,N_35852,N_34423);
nand U40390 (N_40390,N_34569,N_37166);
or U40391 (N_40391,N_39945,N_36452);
nand U40392 (N_40392,N_39903,N_30930);
nor U40393 (N_40393,N_33072,N_30129);
and U40394 (N_40394,N_36276,N_30030);
nor U40395 (N_40395,N_35810,N_38995);
or U40396 (N_40396,N_35984,N_32239);
nand U40397 (N_40397,N_35778,N_38653);
nor U40398 (N_40398,N_35855,N_34487);
and U40399 (N_40399,N_37541,N_35063);
nand U40400 (N_40400,N_30911,N_37495);
or U40401 (N_40401,N_35863,N_38094);
nor U40402 (N_40402,N_31610,N_38991);
nor U40403 (N_40403,N_33311,N_35489);
nor U40404 (N_40404,N_35285,N_30002);
and U40405 (N_40405,N_32288,N_35749);
nor U40406 (N_40406,N_30229,N_38087);
nor U40407 (N_40407,N_38982,N_34835);
nor U40408 (N_40408,N_38237,N_36295);
nor U40409 (N_40409,N_33195,N_35620);
nand U40410 (N_40410,N_37506,N_31919);
or U40411 (N_40411,N_30905,N_32189);
or U40412 (N_40412,N_33281,N_31157);
and U40413 (N_40413,N_39655,N_37574);
nor U40414 (N_40414,N_39636,N_39376);
and U40415 (N_40415,N_37766,N_32170);
or U40416 (N_40416,N_35081,N_34072);
nand U40417 (N_40417,N_34844,N_31938);
nand U40418 (N_40418,N_36361,N_35490);
or U40419 (N_40419,N_34886,N_38361);
nor U40420 (N_40420,N_32073,N_32485);
nor U40421 (N_40421,N_35643,N_37376);
or U40422 (N_40422,N_35407,N_39509);
and U40423 (N_40423,N_33019,N_31472);
or U40424 (N_40424,N_37220,N_38622);
nand U40425 (N_40425,N_32664,N_30815);
xnor U40426 (N_40426,N_38222,N_35382);
nor U40427 (N_40427,N_33500,N_35111);
xor U40428 (N_40428,N_33116,N_39227);
nand U40429 (N_40429,N_35321,N_34608);
nand U40430 (N_40430,N_34445,N_30014);
and U40431 (N_40431,N_31351,N_38519);
and U40432 (N_40432,N_37309,N_37606);
and U40433 (N_40433,N_38148,N_37893);
or U40434 (N_40434,N_38484,N_36118);
xnor U40435 (N_40435,N_39319,N_31975);
or U40436 (N_40436,N_34261,N_37806);
nor U40437 (N_40437,N_37172,N_36252);
or U40438 (N_40438,N_33728,N_38894);
nor U40439 (N_40439,N_34228,N_38206);
xor U40440 (N_40440,N_34005,N_32376);
nor U40441 (N_40441,N_33197,N_34192);
nor U40442 (N_40442,N_31924,N_36761);
or U40443 (N_40443,N_38941,N_37311);
or U40444 (N_40444,N_38045,N_36430);
and U40445 (N_40445,N_31767,N_38200);
or U40446 (N_40446,N_37153,N_37672);
and U40447 (N_40447,N_38006,N_34199);
or U40448 (N_40448,N_30876,N_35845);
and U40449 (N_40449,N_34238,N_36612);
or U40450 (N_40450,N_34442,N_39168);
nor U40451 (N_40451,N_39183,N_35350);
and U40452 (N_40452,N_38057,N_39105);
nand U40453 (N_40453,N_38909,N_34639);
nor U40454 (N_40454,N_30399,N_35134);
nor U40455 (N_40455,N_35537,N_38677);
nand U40456 (N_40456,N_35663,N_36546);
nor U40457 (N_40457,N_35155,N_30069);
or U40458 (N_40458,N_35052,N_37290);
nor U40459 (N_40459,N_33973,N_31603);
and U40460 (N_40460,N_33182,N_31887);
nor U40461 (N_40461,N_32021,N_37748);
and U40462 (N_40462,N_36683,N_38026);
and U40463 (N_40463,N_35912,N_33012);
and U40464 (N_40464,N_31196,N_32976);
or U40465 (N_40465,N_39559,N_34385);
and U40466 (N_40466,N_37878,N_31170);
or U40467 (N_40467,N_36173,N_34618);
nor U40468 (N_40468,N_32941,N_34042);
or U40469 (N_40469,N_30859,N_31315);
and U40470 (N_40470,N_35049,N_33031);
nor U40471 (N_40471,N_39726,N_37522);
or U40472 (N_40472,N_39401,N_35388);
nand U40473 (N_40473,N_33573,N_37109);
or U40474 (N_40474,N_39139,N_34283);
or U40475 (N_40475,N_31360,N_36483);
and U40476 (N_40476,N_35621,N_32046);
and U40477 (N_40477,N_31517,N_35524);
and U40478 (N_40478,N_30325,N_38623);
or U40479 (N_40479,N_38964,N_34352);
nor U40480 (N_40480,N_37951,N_38542);
nor U40481 (N_40481,N_38756,N_34636);
nand U40482 (N_40482,N_37739,N_33771);
xnor U40483 (N_40483,N_38215,N_34899);
and U40484 (N_40484,N_35262,N_31599);
or U40485 (N_40485,N_34027,N_31551);
nand U40486 (N_40486,N_38950,N_32001);
nor U40487 (N_40487,N_39666,N_32869);
or U40488 (N_40488,N_37553,N_37995);
nand U40489 (N_40489,N_37609,N_33296);
and U40490 (N_40490,N_36866,N_35463);
or U40491 (N_40491,N_37741,N_33371);
and U40492 (N_40492,N_38032,N_38525);
nor U40493 (N_40493,N_38168,N_33107);
nand U40494 (N_40494,N_34170,N_30916);
nand U40495 (N_40495,N_39499,N_33439);
nand U40496 (N_40496,N_34809,N_30395);
nor U40497 (N_40497,N_32056,N_31740);
and U40498 (N_40498,N_37126,N_32633);
xnor U40499 (N_40499,N_30185,N_35421);
and U40500 (N_40500,N_37375,N_37082);
or U40501 (N_40501,N_37468,N_35775);
nor U40502 (N_40502,N_33008,N_35926);
or U40503 (N_40503,N_33020,N_35823);
nor U40504 (N_40504,N_39634,N_32631);
nor U40505 (N_40505,N_31641,N_32213);
nor U40506 (N_40506,N_39215,N_34235);
and U40507 (N_40507,N_30319,N_34692);
nor U40508 (N_40508,N_30155,N_31838);
nand U40509 (N_40509,N_30701,N_34629);
and U40510 (N_40510,N_38020,N_34542);
and U40511 (N_40511,N_37440,N_30684);
or U40512 (N_40512,N_32049,N_31452);
or U40513 (N_40513,N_36492,N_39126);
xnor U40514 (N_40514,N_36417,N_35073);
nor U40515 (N_40515,N_31309,N_31274);
nor U40516 (N_40516,N_35767,N_30041);
nand U40517 (N_40517,N_33218,N_30841);
and U40518 (N_40518,N_34846,N_36565);
nor U40519 (N_40519,N_33654,N_32918);
nor U40520 (N_40520,N_36567,N_35988);
and U40521 (N_40521,N_31003,N_33341);
and U40522 (N_40522,N_34122,N_30408);
nand U40523 (N_40523,N_31363,N_38407);
and U40524 (N_40524,N_31813,N_36889);
and U40525 (N_40525,N_39997,N_39766);
xor U40526 (N_40526,N_38210,N_39182);
xnor U40527 (N_40527,N_37750,N_30125);
nand U40528 (N_40528,N_36454,N_34405);
or U40529 (N_40529,N_30037,N_39193);
nand U40530 (N_40530,N_37560,N_33459);
and U40531 (N_40531,N_35802,N_30189);
and U40532 (N_40532,N_34218,N_31589);
and U40533 (N_40533,N_33608,N_32683);
nand U40534 (N_40534,N_38826,N_33308);
nor U40535 (N_40535,N_37586,N_39109);
nand U40536 (N_40536,N_37568,N_33644);
nand U40537 (N_40537,N_36388,N_38092);
or U40538 (N_40538,N_31875,N_39578);
or U40539 (N_40539,N_35267,N_36471);
or U40540 (N_40540,N_31771,N_37384);
and U40541 (N_40541,N_32761,N_34881);
nor U40542 (N_40542,N_36525,N_36675);
nor U40543 (N_40543,N_32679,N_34430);
nand U40544 (N_40544,N_30791,N_39112);
nand U40545 (N_40545,N_37826,N_32882);
or U40546 (N_40546,N_35556,N_39244);
nor U40547 (N_40547,N_31729,N_34799);
nand U40548 (N_40548,N_32567,N_34796);
and U40549 (N_40549,N_32329,N_34028);
xnor U40550 (N_40550,N_39298,N_37822);
nor U40551 (N_40551,N_32410,N_30391);
nand U40552 (N_40552,N_31792,N_30466);
xor U40553 (N_40553,N_39724,N_34901);
and U40554 (N_40554,N_36460,N_38939);
or U40555 (N_40555,N_31120,N_35518);
or U40556 (N_40556,N_31866,N_35450);
nor U40557 (N_40557,N_39583,N_36562);
and U40558 (N_40558,N_31132,N_38198);
or U40559 (N_40559,N_35403,N_36136);
and U40560 (N_40560,N_34135,N_37905);
or U40561 (N_40561,N_35836,N_34637);
nand U40562 (N_40562,N_38673,N_35289);
nand U40563 (N_40563,N_39330,N_36987);
nor U40564 (N_40564,N_34085,N_34665);
xnor U40565 (N_40565,N_37582,N_38879);
nor U40566 (N_40566,N_31156,N_33089);
or U40567 (N_40567,N_35422,N_37851);
nor U40568 (N_40568,N_37599,N_34781);
nand U40569 (N_40569,N_38251,N_36644);
and U40570 (N_40570,N_39437,N_37394);
nor U40571 (N_40571,N_38844,N_34745);
nand U40572 (N_40572,N_33226,N_31333);
or U40573 (N_40573,N_34858,N_34998);
nand U40574 (N_40574,N_37012,N_31704);
nor U40575 (N_40575,N_39341,N_32832);
and U40576 (N_40576,N_33779,N_38867);
or U40577 (N_40577,N_33290,N_37483);
and U40578 (N_40578,N_34504,N_32568);
xor U40579 (N_40579,N_30692,N_38223);
and U40580 (N_40580,N_35576,N_31669);
xor U40581 (N_40581,N_34978,N_30725);
xor U40582 (N_40582,N_34577,N_37328);
or U40583 (N_40583,N_31299,N_37954);
or U40584 (N_40584,N_37796,N_38518);
or U40585 (N_40585,N_32615,N_38987);
or U40586 (N_40586,N_35482,N_30747);
or U40587 (N_40587,N_32292,N_37419);
and U40588 (N_40588,N_38372,N_30209);
xnor U40589 (N_40589,N_39793,N_39991);
or U40590 (N_40590,N_32010,N_31923);
and U40591 (N_40591,N_37993,N_37174);
nor U40592 (N_40592,N_30641,N_34402);
nor U40593 (N_40593,N_31824,N_34291);
nand U40594 (N_40594,N_39900,N_32293);
nor U40595 (N_40595,N_39969,N_36003);
and U40596 (N_40596,N_32259,N_30603);
nand U40597 (N_40597,N_30503,N_39971);
nand U40598 (N_40598,N_37154,N_38526);
nand U40599 (N_40599,N_34249,N_30024);
nor U40600 (N_40600,N_38549,N_35586);
or U40601 (N_40601,N_37294,N_35181);
nand U40602 (N_40602,N_31710,N_32836);
nand U40603 (N_40603,N_32821,N_32746);
xor U40604 (N_40604,N_31570,N_34219);
and U40605 (N_40605,N_30994,N_31913);
or U40606 (N_40606,N_31762,N_31925);
nand U40607 (N_40607,N_39756,N_35015);
or U40608 (N_40608,N_35688,N_31554);
xnor U40609 (N_40609,N_39347,N_38495);
nor U40610 (N_40610,N_38143,N_34580);
and U40611 (N_40611,N_32587,N_34196);
nor U40612 (N_40612,N_39587,N_34121);
xor U40613 (N_40613,N_33351,N_31616);
nor U40614 (N_40614,N_33501,N_32389);
nand U40615 (N_40615,N_31963,N_30349);
and U40616 (N_40616,N_38302,N_35028);
or U40617 (N_40617,N_35084,N_33894);
nand U40618 (N_40618,N_35476,N_31455);
nor U40619 (N_40619,N_35983,N_38832);
or U40620 (N_40620,N_32185,N_39463);
xor U40621 (N_40621,N_30516,N_33759);
and U40622 (N_40622,N_30445,N_35235);
nand U40623 (N_40623,N_30441,N_30913);
nor U40624 (N_40624,N_37493,N_32547);
and U40625 (N_40625,N_38398,N_38287);
nor U40626 (N_40626,N_33221,N_36635);
and U40627 (N_40627,N_32616,N_32735);
or U40628 (N_40628,N_38570,N_35096);
xor U40629 (N_40629,N_30548,N_32212);
or U40630 (N_40630,N_32133,N_37324);
or U40631 (N_40631,N_32340,N_37915);
or U40632 (N_40632,N_30428,N_39026);
nand U40633 (N_40633,N_37067,N_37700);
or U40634 (N_40634,N_36331,N_32979);
or U40635 (N_40635,N_31889,N_38282);
and U40636 (N_40636,N_36779,N_35887);
xor U40637 (N_40637,N_37475,N_38517);
or U40638 (N_40638,N_33215,N_39645);
or U40639 (N_40639,N_32947,N_37656);
xor U40640 (N_40640,N_39028,N_32822);
or U40641 (N_40641,N_33519,N_33300);
nor U40642 (N_40642,N_33367,N_39763);
or U40643 (N_40643,N_30369,N_37110);
xor U40644 (N_40644,N_30296,N_31588);
nor U40645 (N_40645,N_38018,N_30676);
nand U40646 (N_40646,N_36336,N_38522);
and U40647 (N_40647,N_30370,N_34476);
xnor U40648 (N_40648,N_32574,N_32305);
or U40649 (N_40649,N_36553,N_30717);
xnor U40650 (N_40650,N_38001,N_30521);
or U40651 (N_40651,N_39113,N_39979);
nand U40652 (N_40652,N_30048,N_33530);
and U40653 (N_40653,N_36548,N_37799);
nor U40654 (N_40654,N_39892,N_38005);
or U40655 (N_40655,N_35310,N_31031);
and U40656 (N_40656,N_37694,N_35827);
nand U40657 (N_40657,N_35199,N_36112);
nor U40658 (N_40658,N_35826,N_32114);
or U40659 (N_40659,N_36994,N_34280);
nand U40660 (N_40660,N_30086,N_34983);
or U40661 (N_40661,N_37686,N_30571);
nor U40662 (N_40662,N_37207,N_37173);
nand U40663 (N_40663,N_37214,N_32792);
nand U40664 (N_40664,N_31947,N_39155);
and U40665 (N_40665,N_30771,N_39038);
xor U40666 (N_40666,N_38487,N_31827);
xor U40667 (N_40667,N_34454,N_36594);
and U40668 (N_40668,N_39108,N_31176);
nor U40669 (N_40669,N_39651,N_31124);
nor U40670 (N_40670,N_33074,N_33796);
nor U40671 (N_40671,N_35667,N_30846);
or U40672 (N_40672,N_37876,N_35789);
or U40673 (N_40673,N_31318,N_38878);
nor U40674 (N_40674,N_39404,N_34963);
or U40675 (N_40675,N_30637,N_31747);
and U40676 (N_40676,N_36519,N_31126);
and U40677 (N_40677,N_38897,N_35798);
nor U40678 (N_40678,N_37409,N_32476);
or U40679 (N_40679,N_34660,N_39544);
and U40680 (N_40680,N_35098,N_30267);
nand U40681 (N_40681,N_34279,N_33724);
and U40682 (N_40682,N_32309,N_32207);
xnor U40683 (N_40683,N_32255,N_39714);
xnor U40684 (N_40684,N_35851,N_39251);
and U40685 (N_40685,N_30046,N_33928);
and U40686 (N_40686,N_34864,N_33584);
nor U40687 (N_40687,N_35746,N_36808);
nand U40688 (N_40688,N_36764,N_37580);
nand U40689 (N_40689,N_38536,N_38954);
nor U40690 (N_40690,N_35578,N_30073);
and U40691 (N_40691,N_37095,N_34537);
and U40692 (N_40692,N_33910,N_35919);
or U40693 (N_40693,N_37992,N_39637);
nand U40694 (N_40694,N_36870,N_32398);
or U40695 (N_40695,N_33940,N_30578);
or U40696 (N_40696,N_38553,N_34783);
or U40697 (N_40697,N_30378,N_30806);
and U40698 (N_40698,N_31285,N_37872);
nand U40699 (N_40699,N_30252,N_38700);
xnor U40700 (N_40700,N_31010,N_34947);
and U40701 (N_40701,N_36044,N_31595);
or U40702 (N_40702,N_30279,N_38942);
xor U40703 (N_40703,N_39069,N_34377);
nand U40704 (N_40704,N_37867,N_32270);
or U40705 (N_40705,N_34523,N_36749);
nor U40706 (N_40706,N_39475,N_34272);
and U40707 (N_40707,N_35202,N_32150);
nand U40708 (N_40708,N_38938,N_33682);
or U40709 (N_40709,N_35909,N_33665);
and U40710 (N_40710,N_30344,N_37216);
and U40711 (N_40711,N_35040,N_34174);
nor U40712 (N_40712,N_33518,N_36245);
or U40713 (N_40713,N_33365,N_34374);
or U40714 (N_40714,N_30436,N_33077);
nand U40715 (N_40715,N_35985,N_30218);
and U40716 (N_40716,N_37671,N_30591);
nand U40717 (N_40717,N_32815,N_30161);
nor U40718 (N_40718,N_32464,N_32944);
nand U40719 (N_40719,N_35238,N_30665);
nor U40720 (N_40720,N_35359,N_38256);
and U40721 (N_40721,N_30461,N_39759);
or U40722 (N_40722,N_31933,N_35993);
or U40723 (N_40723,N_34437,N_33559);
or U40724 (N_40724,N_36529,N_38529);
nor U40725 (N_40725,N_30149,N_33243);
nand U40726 (N_40726,N_38068,N_39628);
xor U40727 (N_40727,N_31705,N_37703);
nor U40728 (N_40728,N_36129,N_39149);
nand U40729 (N_40729,N_32527,N_35552);
and U40730 (N_40730,N_35066,N_36856);
and U40731 (N_40731,N_38530,N_38327);
nand U40732 (N_40732,N_31064,N_30673);
nand U40733 (N_40733,N_33716,N_30856);
or U40734 (N_40734,N_30552,N_34620);
and U40735 (N_40735,N_33942,N_30486);
nand U40736 (N_40736,N_33624,N_39916);
nor U40737 (N_40737,N_33684,N_37736);
nor U40738 (N_40738,N_39957,N_33911);
xnor U40739 (N_40739,N_37055,N_30147);
and U40740 (N_40740,N_36816,N_36348);
or U40741 (N_40741,N_33694,N_31618);
or U40742 (N_40742,N_33205,N_30419);
nand U40743 (N_40743,N_34123,N_35411);
nor U40744 (N_40744,N_38385,N_38608);
and U40745 (N_40745,N_39550,N_35056);
nor U40746 (N_40746,N_34002,N_33768);
or U40747 (N_40747,N_39248,N_37010);
or U40748 (N_40748,N_34242,N_35441);
or U40749 (N_40749,N_32184,N_32997);
nand U40750 (N_40750,N_30478,N_36945);
nand U40751 (N_40751,N_39398,N_36481);
xor U40752 (N_40752,N_31062,N_35483);
xor U40753 (N_40753,N_33816,N_36007);
or U40754 (N_40754,N_33183,N_36849);
and U40755 (N_40755,N_37338,N_36692);
and U40756 (N_40756,N_30789,N_37935);
and U40757 (N_40757,N_31466,N_31895);
nand U40758 (N_40758,N_31322,N_33173);
nor U40759 (N_40759,N_34708,N_34415);
nand U40760 (N_40760,N_36831,N_38108);
or U40761 (N_40761,N_39805,N_39670);
xnor U40762 (N_40762,N_33890,N_39184);
xnor U40763 (N_40763,N_39772,N_36741);
xnor U40764 (N_40764,N_34852,N_35916);
nand U40765 (N_40765,N_35649,N_36236);
or U40766 (N_40766,N_39799,N_30119);
nor U40767 (N_40767,N_38468,N_32385);
xnor U40768 (N_40768,N_32597,N_30660);
and U40769 (N_40769,N_32867,N_33000);
nor U40770 (N_40770,N_33266,N_32444);
nand U40771 (N_40771,N_35465,N_30656);
nor U40772 (N_40772,N_36952,N_30204);
and U40773 (N_40773,N_38002,N_30250);
nand U40774 (N_40774,N_36285,N_31166);
or U40775 (N_40775,N_31643,N_37778);
and U40776 (N_40776,N_37761,N_37079);
and U40777 (N_40777,N_36901,N_30525);
nor U40778 (N_40778,N_38946,N_35255);
or U40779 (N_40779,N_32923,N_31511);
or U40780 (N_40780,N_30031,N_39438);
nor U40781 (N_40781,N_37022,N_35661);
nand U40782 (N_40782,N_37412,N_33316);
nand U40783 (N_40783,N_31635,N_35502);
and U40784 (N_40784,N_38453,N_33668);
and U40785 (N_40785,N_35128,N_35543);
nand U40786 (N_40786,N_35327,N_31955);
or U40787 (N_40787,N_34748,N_38561);
xor U40788 (N_40788,N_39739,N_33260);
or U40789 (N_40789,N_37190,N_37317);
or U40790 (N_40790,N_34627,N_34851);
nand U40791 (N_40791,N_34270,N_35718);
nand U40792 (N_40792,N_37856,N_33079);
or U40793 (N_40793,N_37125,N_34539);
nor U40794 (N_40794,N_36165,N_32685);
or U40795 (N_40795,N_39527,N_31217);
nor U40796 (N_40796,N_37451,N_31651);
nor U40797 (N_40797,N_33892,N_37999);
nand U40798 (N_40798,N_32630,N_37186);
nand U40799 (N_40799,N_31036,N_39521);
and U40800 (N_40800,N_35393,N_31483);
and U40801 (N_40801,N_36397,N_39729);
nand U40802 (N_40802,N_30242,N_38959);
nand U40803 (N_40803,N_33631,N_38661);
xor U40804 (N_40804,N_39567,N_31264);
nand U40805 (N_40805,N_34820,N_31498);
or U40806 (N_40806,N_31984,N_35788);
or U40807 (N_40807,N_33228,N_30907);
and U40808 (N_40808,N_39907,N_34965);
and U40809 (N_40809,N_34180,N_30297);
nor U40810 (N_40810,N_30322,N_30668);
and U40811 (N_40811,N_33685,N_38786);
nand U40812 (N_40812,N_31138,N_39941);
nor U40813 (N_40813,N_37877,N_34801);
xor U40814 (N_40814,N_33837,N_35115);
nor U40815 (N_40815,N_37402,N_39522);
xnor U40816 (N_40816,N_33820,N_35672);
and U40817 (N_40817,N_32954,N_36267);
and U40818 (N_40818,N_33669,N_36753);
or U40819 (N_40819,N_33210,N_35608);
xor U40820 (N_40820,N_37432,N_34347);
and U40821 (N_40821,N_35318,N_37508);
nor U40822 (N_40822,N_36750,N_36140);
nand U40823 (N_40823,N_31869,N_33719);
xor U40824 (N_40824,N_33345,N_31035);
nand U40825 (N_40825,N_30311,N_35290);
or U40826 (N_40826,N_33307,N_33417);
nor U40827 (N_40827,N_36721,N_33626);
nor U40828 (N_40828,N_31505,N_33854);
nor U40829 (N_40829,N_34315,N_30675);
or U40830 (N_40830,N_37000,N_31381);
and U40831 (N_40831,N_35815,N_39023);
xor U40832 (N_40832,N_30358,N_32788);
nand U40833 (N_40833,N_39545,N_39101);
nand U40834 (N_40834,N_39922,N_33601);
and U40835 (N_40835,N_39223,N_30447);
xor U40836 (N_40836,N_31694,N_33135);
nor U40837 (N_40837,N_30921,N_34607);
and U40838 (N_40838,N_32417,N_30545);
and U40839 (N_40839,N_36809,N_39352);
and U40840 (N_40840,N_35816,N_39627);
and U40841 (N_40841,N_36230,N_38990);
nand U40842 (N_40842,N_35974,N_31577);
nand U40843 (N_40843,N_38545,N_39336);
nor U40844 (N_40844,N_32117,N_38575);
nor U40845 (N_40845,N_31212,N_39868);
xnor U40846 (N_40846,N_34290,N_39792);
or U40847 (N_40847,N_39679,N_33389);
nand U40848 (N_40848,N_39689,N_32834);
xnor U40849 (N_40849,N_37536,N_39349);
nor U40850 (N_40850,N_36942,N_36740);
nor U40851 (N_40851,N_33246,N_33564);
nor U40852 (N_40852,N_39111,N_33775);
and U40853 (N_40853,N_35197,N_37049);
and U40854 (N_40854,N_33204,N_33715);
and U40855 (N_40855,N_34326,N_33914);
nor U40856 (N_40856,N_33731,N_38313);
nor U40857 (N_40857,N_33491,N_33493);
or U40858 (N_40858,N_30105,N_33957);
xnor U40859 (N_40859,N_36793,N_33358);
or U40860 (N_40860,N_34224,N_38054);
and U40861 (N_40861,N_33359,N_38808);
or U40862 (N_40862,N_38792,N_31556);
and U40863 (N_40863,N_30972,N_34525);
and U40864 (N_40864,N_38845,N_36476);
and U40865 (N_40865,N_37144,N_32135);
and U40866 (N_40866,N_31784,N_33385);
xnor U40867 (N_40867,N_38663,N_30433);
nand U40868 (N_40868,N_30429,N_32859);
and U40869 (N_40869,N_36803,N_35105);
and U40870 (N_40870,N_39205,N_36796);
nor U40871 (N_40871,N_33686,N_37625);
and U40872 (N_40872,N_32267,N_38591);
nor U40873 (N_40873,N_32391,N_35522);
nand U40874 (N_40874,N_30053,N_31037);
or U40875 (N_40875,N_31178,N_31648);
and U40876 (N_40876,N_33106,N_37615);
nor U40877 (N_40877,N_39973,N_31378);
nor U40878 (N_40878,N_35392,N_33526);
nand U40879 (N_40879,N_37316,N_39406);
xor U40880 (N_40880,N_31681,N_31391);
nor U40881 (N_40881,N_31897,N_31525);
or U40882 (N_40882,N_39492,N_31137);
and U40883 (N_40883,N_36545,N_33967);
or U40884 (N_40884,N_36193,N_30757);
nor U40885 (N_40885,N_34125,N_36591);
nor U40886 (N_40886,N_32079,N_31834);
nand U40887 (N_40887,N_31080,N_33015);
nand U40888 (N_40888,N_38697,N_33781);
or U40889 (N_40889,N_31343,N_39258);
nor U40890 (N_40890,N_39935,N_38512);
or U40891 (N_40891,N_39127,N_33623);
or U40892 (N_40892,N_35183,N_30151);
xor U40893 (N_40893,N_38862,N_36800);
or U40894 (N_40894,N_37753,N_36672);
or U40895 (N_40895,N_37688,N_33353);
nand U40896 (N_40896,N_37199,N_33750);
xor U40897 (N_40897,N_34134,N_35943);
nor U40898 (N_40898,N_38117,N_39229);
nor U40899 (N_40899,N_36302,N_34381);
and U40900 (N_40900,N_31348,N_33740);
nor U40901 (N_40901,N_36504,N_34916);
xor U40902 (N_40902,N_32627,N_35322);
and U40903 (N_40903,N_32736,N_31702);
nor U40904 (N_40904,N_35896,N_30230);
or U40905 (N_40905,N_37934,N_39259);
nand U40906 (N_40906,N_39914,N_36374);
and U40907 (N_40907,N_39195,N_33052);
xor U40908 (N_40908,N_33479,N_32690);
nand U40909 (N_40909,N_36765,N_32534);
nor U40910 (N_40910,N_38425,N_38721);
and U40911 (N_40911,N_37268,N_38691);
xnor U40912 (N_40912,N_32709,N_35675);
xor U40913 (N_40913,N_31836,N_30492);
and U40914 (N_40914,N_31190,N_31282);
or U40915 (N_40915,N_36643,N_38109);
or U40916 (N_40916,N_38813,N_33938);
nand U40917 (N_40917,N_39425,N_32463);
and U40918 (N_40918,N_30793,N_30719);
nor U40919 (N_40919,N_35185,N_32565);
nor U40920 (N_40920,N_32250,N_34062);
nand U40921 (N_40921,N_38935,N_30481);
xnor U40922 (N_40922,N_38877,N_34911);
nor U40923 (N_40923,N_34099,N_32658);
nand U40924 (N_40924,N_39548,N_38093);
nor U40925 (N_40925,N_34365,N_39764);
nor U40926 (N_40926,N_33441,N_33418);
or U40927 (N_40927,N_39103,N_35700);
and U40928 (N_40928,N_33984,N_38771);
nor U40929 (N_40929,N_39715,N_33360);
or U40930 (N_40930,N_30958,N_38443);
xnor U40931 (N_40931,N_34959,N_35521);
or U40932 (N_40932,N_31566,N_37757);
or U40933 (N_40933,N_35540,N_38724);
or U40934 (N_40934,N_35177,N_36895);
and U40935 (N_40935,N_32577,N_32624);
nor U40936 (N_40936,N_37139,N_36424);
nand U40937 (N_40937,N_34755,N_37396);
nor U40938 (N_40938,N_38088,N_35969);
nor U40939 (N_40939,N_37002,N_39674);
nor U40940 (N_40940,N_36159,N_31726);
and U40941 (N_40941,N_39862,N_34439);
or U40942 (N_40942,N_36137,N_39034);
or U40943 (N_40943,N_32330,N_31775);
nand U40944 (N_40944,N_36917,N_32275);
and U40945 (N_40945,N_32584,N_33393);
nand U40946 (N_40946,N_39701,N_39639);
nor U40947 (N_40947,N_39214,N_38535);
nor U40948 (N_40948,N_36629,N_39517);
nand U40949 (N_40949,N_35092,N_33002);
nor U40950 (N_40950,N_39465,N_31012);
xnor U40951 (N_40951,N_32907,N_33108);
nor U40952 (N_40952,N_36569,N_34870);
and U40953 (N_40953,N_39180,N_36024);
nand U40954 (N_40954,N_37932,N_30318);
nand U40955 (N_40955,N_38546,N_34524);
or U40956 (N_40956,N_33658,N_39284);
xor U40957 (N_40957,N_32920,N_37607);
and U40958 (N_40958,N_33998,N_33548);
nor U40959 (N_40959,N_36141,N_32308);
nor U40960 (N_40960,N_31159,N_39596);
or U40961 (N_40961,N_33961,N_34116);
and U40962 (N_40962,N_36568,N_32852);
nor U40963 (N_40963,N_36742,N_38969);
nor U40964 (N_40964,N_39302,N_36107);
xnor U40965 (N_40965,N_34927,N_30261);
or U40966 (N_40966,N_30329,N_38660);
and U40967 (N_40967,N_35735,N_35804);
nand U40968 (N_40968,N_39613,N_39057);
nand U40969 (N_40969,N_31390,N_34360);
and U40970 (N_40970,N_38949,N_35464);
or U40971 (N_40971,N_38474,N_34139);
and U40972 (N_40972,N_35370,N_35041);
nand U40973 (N_40973,N_30981,N_35241);
and U40974 (N_40974,N_33131,N_34496);
xor U40975 (N_40975,N_35331,N_35425);
nand U40976 (N_40976,N_35881,N_38898);
nand U40977 (N_40977,N_35890,N_34469);
nand U40978 (N_40978,N_34891,N_36592);
or U40979 (N_40979,N_34563,N_35158);
nand U40980 (N_40980,N_33209,N_35334);
nor U40981 (N_40981,N_39541,N_35190);
nand U40982 (N_40982,N_33368,N_33535);
nor U40983 (N_40983,N_33945,N_31331);
or U40984 (N_40984,N_32550,N_32879);
nor U40985 (N_40985,N_30488,N_39982);
nor U40986 (N_40986,N_37333,N_33472);
nor U40987 (N_40987,N_39978,N_34478);
and U40988 (N_40988,N_33872,N_31578);
nand U40989 (N_40989,N_34827,N_39056);
nand U40990 (N_40990,N_34310,N_38528);
and U40991 (N_40991,N_35404,N_36355);
nand U40992 (N_40992,N_35587,N_38779);
and U40993 (N_40993,N_30172,N_32732);
nor U40994 (N_40994,N_31549,N_30967);
and U40995 (N_40995,N_30100,N_31721);
and U40996 (N_40996,N_30364,N_32080);
nand U40997 (N_40997,N_33495,N_37660);
nand U40998 (N_40998,N_35286,N_37194);
nor U40999 (N_40999,N_35323,N_34046);
xnor U41000 (N_41000,N_31273,N_35860);
or U41001 (N_41001,N_30998,N_31714);
nor U41002 (N_41002,N_39266,N_31266);
or U41003 (N_41003,N_37653,N_35402);
nand U41004 (N_41004,N_32223,N_39090);
and U41005 (N_41005,N_31067,N_32344);
xor U41006 (N_41006,N_32546,N_37228);
xnor U41007 (N_41007,N_35519,N_34281);
and U41008 (N_41008,N_33154,N_36729);
or U41009 (N_41009,N_36781,N_35803);
and U41010 (N_41010,N_31594,N_39556);
nor U41011 (N_41011,N_33375,N_34923);
nand U41012 (N_41012,N_35107,N_33233);
or U41013 (N_41013,N_34335,N_31005);
xnor U41014 (N_41014,N_34181,N_35865);
or U41015 (N_41015,N_38202,N_33255);
and U41016 (N_41016,N_35642,N_37916);
nor U41017 (N_41017,N_34688,N_31248);
nand U41018 (N_41018,N_34207,N_33332);
and U41019 (N_41019,N_30544,N_36723);
and U41020 (N_41020,N_30434,N_31099);
nand U41021 (N_41021,N_35249,N_38152);
nand U41022 (N_41022,N_35222,N_37489);
nand U41023 (N_41023,N_39767,N_34706);
nand U41024 (N_41024,N_39114,N_30371);
and U41025 (N_41025,N_35722,N_30304);
xnor U41026 (N_41026,N_38427,N_37620);
xor U41027 (N_41027,N_39606,N_35510);
nor U41028 (N_41028,N_39650,N_36448);
nor U41029 (N_41029,N_34663,N_33364);
and U41030 (N_41030,N_37359,N_30638);
or U41031 (N_41031,N_35095,N_39904);
nand U41032 (N_41032,N_35653,N_31546);
or U41033 (N_41033,N_35651,N_31388);
or U41034 (N_41034,N_32781,N_39732);
or U41035 (N_41035,N_37600,N_33651);
xnor U41036 (N_41036,N_35666,N_39164);
and U41037 (N_41037,N_31893,N_38915);
and U41038 (N_41038,N_37884,N_36732);
and U41039 (N_41039,N_33922,N_39738);
nor U41040 (N_41040,N_32734,N_39472);
nor U41041 (N_41041,N_36882,N_30026);
or U41042 (N_41042,N_39075,N_37128);
or U41043 (N_41043,N_39462,N_34455);
nor U41044 (N_41044,N_33772,N_38118);
xnor U41045 (N_41045,N_38315,N_38793);
and U41046 (N_41046,N_35454,N_37296);
nand U41047 (N_41047,N_33730,N_32728);
or U41048 (N_41048,N_34419,N_33845);
or U41049 (N_41049,N_37678,N_38672);
and U41050 (N_41050,N_30302,N_34893);
xnor U41051 (N_41051,N_32348,N_31559);
and U41052 (N_41052,N_35584,N_37044);
nand U41053 (N_41053,N_37028,N_37471);
or U41054 (N_41054,N_30943,N_34750);
and U41055 (N_41055,N_39024,N_33349);
and U41056 (N_41056,N_39861,N_31837);
and U41057 (N_41057,N_31523,N_37341);
nand U41058 (N_41058,N_32112,N_32889);
and U41059 (N_41059,N_33408,N_31185);
and U41060 (N_41060,N_37337,N_33525);
nand U41061 (N_41061,N_35150,N_36503);
or U41062 (N_41062,N_34203,N_31175);
and U41063 (N_41063,N_34435,N_38056);
nand U41064 (N_41064,N_34159,N_30396);
nor U41065 (N_41065,N_36090,N_30903);
nand U41066 (N_41066,N_34994,N_30624);
nor U41067 (N_41067,N_31995,N_37369);
nand U41068 (N_41068,N_39641,N_39762);
and U41069 (N_41069,N_33026,N_39500);
or U41070 (N_41070,N_31800,N_39591);
nand U41071 (N_41071,N_35641,N_31950);
nor U41072 (N_41072,N_34212,N_30426);
or U41073 (N_41073,N_33476,N_31873);
nand U41074 (N_41074,N_30008,N_36602);
and U41075 (N_41075,N_39047,N_34814);
nor U41076 (N_41076,N_37952,N_38205);
or U41077 (N_41077,N_34292,N_30581);
nor U41078 (N_41078,N_30760,N_34343);
nor U41079 (N_41079,N_33613,N_39631);
nor U41080 (N_41080,N_36299,N_30543);
or U41081 (N_41081,N_33536,N_33988);
nor U41082 (N_41082,N_34247,N_36514);
nor U41083 (N_41083,N_37474,N_38937);
or U41084 (N_41084,N_33935,N_36666);
and U41085 (N_41085,N_35648,N_36801);
nor U41086 (N_41086,N_33038,N_33704);
or U41087 (N_41087,N_30193,N_33241);
nor U41088 (N_41088,N_30761,N_39267);
nand U41089 (N_41089,N_31851,N_32129);
nor U41090 (N_41090,N_38441,N_30529);
or U41091 (N_41091,N_33980,N_34393);
and U41092 (N_41092,N_32743,N_37913);
or U41093 (N_41093,N_36508,N_35757);
nor U41094 (N_41094,N_33546,N_30704);
nand U41095 (N_41095,N_38304,N_32704);
or U41096 (N_41096,N_35252,N_37706);
nand U41097 (N_41097,N_30561,N_38652);
nand U41098 (N_41098,N_34137,N_32061);
nand U41099 (N_41099,N_30714,N_39511);
or U41100 (N_41100,N_36724,N_30055);
and U41101 (N_41101,N_35949,N_36518);
or U41102 (N_41102,N_32862,N_38086);
and U41103 (N_41103,N_39863,N_35925);
nand U41104 (N_41104,N_30617,N_39622);
nor U41105 (N_41105,N_32881,N_38404);
and U41106 (N_41106,N_30575,N_34854);
or U41107 (N_41107,N_32772,N_39399);
nor U41108 (N_41108,N_36585,N_39557);
nand U41109 (N_41109,N_30817,N_32622);
nand U41110 (N_41110,N_38579,N_36228);
and U41111 (N_41111,N_39199,N_36845);
nor U41112 (N_41112,N_34237,N_31620);
nor U41113 (N_41113,N_39503,N_36930);
nand U41114 (N_41114,N_31173,N_39035);
nor U41115 (N_41115,N_34300,N_32967);
nand U41116 (N_41116,N_35908,N_33153);
nand U41117 (N_41117,N_36414,N_32540);
nand U41118 (N_41118,N_36805,N_34513);
nor U41119 (N_41119,N_33865,N_34284);
nor U41120 (N_41120,N_32081,N_37165);
nand U41121 (N_41121,N_33095,N_30234);
nand U41122 (N_41122,N_37391,N_37715);
nor U41123 (N_41123,N_31143,N_39846);
or U41124 (N_41124,N_37828,N_32951);
or U41125 (N_41125,N_36593,N_33496);
xnor U41126 (N_41126,N_34396,N_36207);
nand U41127 (N_41127,N_36271,N_31116);
nand U41128 (N_41128,N_31891,N_32037);
and U41129 (N_41129,N_37212,N_35245);
nand U41130 (N_41130,N_37246,N_39575);
or U41131 (N_41131,N_34486,N_34029);
xor U41132 (N_41132,N_38264,N_33804);
nand U41133 (N_41133,N_34341,N_39160);
nand U41134 (N_41134,N_35499,N_38809);
nand U41135 (N_41135,N_30021,N_30720);
nand U41136 (N_41136,N_35180,N_35963);
or U41137 (N_41137,N_31688,N_39357);
nand U41138 (N_41138,N_31302,N_36821);
nor U41139 (N_41139,N_31395,N_38981);
or U41140 (N_41140,N_39933,N_37896);
nor U41141 (N_41141,N_37405,N_38115);
or U41142 (N_41142,N_35284,N_35491);
or U41143 (N_41143,N_37385,N_32496);
and U41144 (N_41144,N_31095,N_35124);
xor U41145 (N_41145,N_37081,N_38236);
nor U41146 (N_41146,N_33337,N_31644);
xnor U41147 (N_41147,N_37160,N_39483);
nand U41148 (N_41148,N_39552,N_32315);
nand U41149 (N_41149,N_36176,N_31431);
nand U41150 (N_41150,N_35214,N_31357);
nand U41151 (N_41151,N_33416,N_30126);
nor U41152 (N_41152,N_39145,N_30255);
nor U41153 (N_41153,N_39317,N_36903);
nand U41154 (N_41154,N_37122,N_31485);
nor U41155 (N_41155,N_34596,N_32227);
nand U41156 (N_41156,N_37629,N_38538);
nor U41157 (N_41157,N_38424,N_39827);
nand U41158 (N_41158,N_39320,N_37830);
and U41159 (N_41159,N_30239,N_35210);
nor U41160 (N_41160,N_38810,N_38423);
and U41161 (N_41161,N_32052,N_37512);
nand U41162 (N_41162,N_31966,N_39321);
nand U41163 (N_41163,N_38323,N_38899);
nor U41164 (N_41164,N_39006,N_39062);
xor U41165 (N_41165,N_36609,N_33764);
nand U41166 (N_41166,N_39345,N_33711);
or U41167 (N_41167,N_37025,N_30965);
or U41168 (N_41168,N_32232,N_32745);
or U41169 (N_41169,N_31290,N_34088);
or U41170 (N_41170,N_38725,N_33414);
nand U41171 (N_41171,N_34017,N_35340);
or U41172 (N_41172,N_31103,N_39011);
nor U41173 (N_41173,N_39308,N_33298);
nor U41174 (N_41174,N_35486,N_32441);
and U41175 (N_41175,N_31249,N_38357);
nor U41176 (N_41176,N_34597,N_31531);
or U41177 (N_41177,N_36531,N_39135);
nand U41178 (N_41178,N_36067,N_33860);
nor U41179 (N_41179,N_36163,N_34001);
and U41180 (N_41180,N_36005,N_31810);
or U41181 (N_41181,N_31516,N_34615);
or U41182 (N_41182,N_37521,N_35487);
xor U41183 (N_41183,N_31075,N_33599);
nor U41184 (N_41184,N_37457,N_33190);
nand U41185 (N_41185,N_38009,N_35627);
or U41186 (N_41186,N_32221,N_30401);
and U41187 (N_41187,N_39377,N_31540);
nand U41188 (N_41188,N_39476,N_37982);
nand U41189 (N_41189,N_33674,N_36535);
and U41190 (N_41190,N_34392,N_35088);
nand U41191 (N_41191,N_34975,N_39553);
nor U41192 (N_41192,N_38513,N_38442);
and U41193 (N_41193,N_31396,N_38352);
nand U41194 (N_41194,N_31349,N_39633);
nand U41195 (N_41195,N_32747,N_38884);
and U41196 (N_41196,N_31653,N_38842);
nand U41197 (N_41197,N_39173,N_36194);
and U41198 (N_41198,N_33236,N_39324);
and U41199 (N_41199,N_39358,N_32420);
and U41200 (N_41200,N_31025,N_31487);
nor U41201 (N_41201,N_36822,N_38983);
and U41202 (N_41202,N_33460,N_37225);
and U41203 (N_41203,N_38030,N_33690);
and U41204 (N_41204,N_33053,N_38841);
and U41205 (N_41205,N_34307,N_38112);
nor U41206 (N_41206,N_34658,N_39609);
nor U41207 (N_41207,N_34550,N_36157);
nor U41208 (N_41208,N_33230,N_34932);
or U41209 (N_41209,N_32672,N_37855);
nor U41210 (N_41210,N_34391,N_31361);
xnor U41211 (N_41211,N_37517,N_30794);
and U41212 (N_41212,N_36105,N_32218);
nand U41213 (N_41213,N_36990,N_37840);
xnor U41214 (N_41214,N_32883,N_30739);
nand U41215 (N_41215,N_34092,N_32430);
and U41216 (N_41216,N_39855,N_30079);
and U41217 (N_41217,N_39307,N_37836);
nor U41218 (N_41218,N_36406,N_36979);
nor U41219 (N_41219,N_37792,N_38314);
and U41220 (N_41220,N_30272,N_34677);
and U41221 (N_41221,N_32372,N_32659);
and U41222 (N_41222,N_38013,N_30738);
or U41223 (N_41223,N_32201,N_38925);
or U41224 (N_41224,N_35932,N_38632);
or U41225 (N_41225,N_39867,N_33265);
nand U41226 (N_41226,N_34130,N_31535);
and U41227 (N_41227,N_38705,N_36128);
or U41228 (N_41228,N_31330,N_33248);
or U41229 (N_41229,N_37242,N_35024);
and U41230 (N_41230,N_34880,N_36168);
and U41231 (N_41231,N_32027,N_34333);
nor U41232 (N_41232,N_39447,N_31432);
nor U41233 (N_41233,N_32483,N_32145);
or U41234 (N_41234,N_34740,N_36303);
nor U41235 (N_41235,N_30076,N_30484);
and U41236 (N_41236,N_30458,N_35039);
nand U41237 (N_41237,N_35902,N_35367);
and U41238 (N_41238,N_34718,N_38737);
nand U41239 (N_41239,N_39211,N_32620);
and U41240 (N_41240,N_32380,N_31084);
or U41241 (N_41241,N_35379,N_36293);
nand U41242 (N_41242,N_37551,N_39880);
or U41243 (N_41243,N_36620,N_31845);
nand U41244 (N_41244,N_37751,N_36887);
xnor U41245 (N_41245,N_32327,N_30672);
nor U41246 (N_41246,N_33767,N_33705);
or U41247 (N_41247,N_31631,N_38395);
nor U41248 (N_41248,N_30456,N_32648);
and U41249 (N_41249,N_36613,N_37486);
nand U41250 (N_41250,N_39623,N_38931);
and U41251 (N_41251,N_38571,N_31586);
nor U41252 (N_41252,N_36783,N_33593);
nand U41253 (N_41253,N_34010,N_31015);
nor U41254 (N_41254,N_32006,N_34093);
nand U41255 (N_41255,N_30015,N_37428);
nor U41256 (N_41256,N_33051,N_37492);
nor U41257 (N_41257,N_38027,N_30830);
nor U41258 (N_41258,N_31503,N_31730);
nor U41259 (N_41259,N_36219,N_36937);
xnor U41260 (N_41260,N_36369,N_34786);
nand U41261 (N_41261,N_33628,N_33586);
nand U41262 (N_41262,N_35196,N_39176);
nor U41263 (N_41263,N_34837,N_37446);
and U41264 (N_41264,N_38135,N_35849);
and U41265 (N_41265,N_31430,N_31293);
and U41266 (N_41266,N_30533,N_39942);
and U41267 (N_41267,N_32187,N_35555);
and U41268 (N_41268,N_38515,N_36673);
and U41269 (N_41269,N_39212,N_30384);
nand U41270 (N_41270,N_36108,N_31614);
and U41271 (N_41271,N_31470,N_34680);
nand U41272 (N_41272,N_32887,N_32324);
nand U41273 (N_41273,N_34431,N_33862);
and U41274 (N_41274,N_39691,N_32600);
nor U41275 (N_41275,N_35613,N_34842);
nand U41276 (N_41276,N_31943,N_34149);
xnor U41277 (N_41277,N_34053,N_30948);
xnor U41278 (N_41278,N_32044,N_34133);
nand U41279 (N_41279,N_30206,N_37933);
nor U41280 (N_41280,N_39683,N_34384);
nand U41281 (N_41281,N_34571,N_34359);
and U41282 (N_41282,N_37874,N_34368);
and U41283 (N_41283,N_35118,N_33811);
nand U41284 (N_41284,N_37947,N_34158);
nand U41285 (N_41285,N_39339,N_39328);
nor U41286 (N_41286,N_34096,N_31420);
or U41287 (N_41287,N_39980,N_38712);
or U41288 (N_41288,N_35676,N_39099);
nor U41289 (N_41289,N_39048,N_38766);
and U41290 (N_41290,N_32188,N_38621);
and U41291 (N_41291,N_37115,N_31642);
nand U41292 (N_41292,N_31047,N_33653);
nor U41293 (N_41293,N_35940,N_39159);
and U41294 (N_41294,N_37683,N_38250);
nand U41295 (N_41295,N_30236,N_35573);
and U41296 (N_41296,N_31613,N_34257);
and U41297 (N_41297,N_36616,N_33788);
nand U41298 (N_41298,N_30315,N_34604);
or U41299 (N_41299,N_32634,N_39427);
nand U41300 (N_41300,N_37937,N_33363);
and U41301 (N_41301,N_37211,N_39141);
nand U41302 (N_41302,N_36166,N_38125);
nand U41303 (N_41303,N_39037,N_31358);
nor U41304 (N_41304,N_35991,N_36178);
and U41305 (N_41305,N_30966,N_37810);
and U41306 (N_41306,N_33549,N_36551);
xnor U41307 (N_41307,N_33882,N_36407);
nand U41308 (N_41308,N_36206,N_33995);
nor U41309 (N_41309,N_33091,N_32623);
or U41310 (N_41310,N_33790,N_30175);
nor U41311 (N_41311,N_31972,N_36345);
and U41312 (N_41312,N_31846,N_32778);
xnor U41313 (N_41313,N_37051,N_33415);
nor U41314 (N_41314,N_31362,N_38996);
xor U41315 (N_41315,N_30607,N_39561);
and U41316 (N_41316,N_31659,N_36794);
nor U41317 (N_41317,N_38980,N_39161);
and U41318 (N_41318,N_37899,N_33164);
xor U41319 (N_41319,N_39659,N_39533);
and U41320 (N_41320,N_38226,N_33156);
nor U41321 (N_41321,N_30502,N_30341);
or U41322 (N_41322,N_34581,N_39271);
nand U41323 (N_41323,N_39614,N_31463);
and U41324 (N_41324,N_33471,N_36662);
nand U41325 (N_41325,N_35341,N_33558);
or U41326 (N_41326,N_32668,N_32539);
or U41327 (N_41327,N_37793,N_37131);
or U41328 (N_41328,N_37198,N_38912);
xor U41329 (N_41329,N_37563,N_38267);
nand U41330 (N_41330,N_36455,N_37041);
xor U41331 (N_41331,N_30848,N_34721);
nand U41332 (N_41332,N_36494,N_39647);
or U41333 (N_41333,N_38448,N_31192);
nand U41334 (N_41334,N_31016,N_37782);
and U41335 (N_41335,N_38533,N_30653);
nor U41336 (N_41336,N_36814,N_38612);
and U41337 (N_41337,N_38288,N_35031);
xor U41338 (N_41338,N_31449,N_33397);
xnor U41339 (N_41339,N_34988,N_35554);
nand U41340 (N_41340,N_39888,N_32585);
nor U41341 (N_41341,N_38367,N_34386);
nor U41342 (N_41342,N_31774,N_34997);
and U41343 (N_41343,N_30375,N_39116);
nand U41344 (N_41344,N_32912,N_34232);
or U41345 (N_41345,N_34734,N_34609);
or U41346 (N_41346,N_34778,N_36450);
xor U41347 (N_41347,N_38816,N_35083);
and U41348 (N_41348,N_37668,N_37289);
nand U41349 (N_41349,N_38787,N_39913);
or U41350 (N_41350,N_39467,N_32523);
nand U41351 (N_41351,N_30559,N_34073);
xor U41352 (N_41352,N_34086,N_37335);
and U41353 (N_41353,N_32693,N_37674);
nand U41354 (N_41354,N_34108,N_38586);
nor U41355 (N_41355,N_31434,N_30901);
xnor U41356 (N_41356,N_33339,N_34025);
nor U41357 (N_41357,N_33211,N_37267);
nor U41358 (N_41358,N_33499,N_34467);
nand U41359 (N_41359,N_38461,N_32196);
nand U41360 (N_41360,N_37424,N_30936);
nand U41361 (N_41361,N_31180,N_39387);
and U41362 (N_41362,N_33792,N_32338);
and U41363 (N_41363,N_33489,N_35050);
or U41364 (N_41364,N_36815,N_35044);
nor U41365 (N_41365,N_35959,N_38051);
xnor U41366 (N_41366,N_37192,N_38977);
nand U41367 (N_41367,N_30421,N_30584);
or U41368 (N_41368,N_32394,N_31230);
or U41369 (N_41369,N_35469,N_33338);
nor U41370 (N_41370,N_30620,N_37559);
nand U41371 (N_41371,N_39265,N_34614);
nor U41372 (N_41372,N_35317,N_35361);
nand U41373 (N_41373,N_38110,N_36312);
nor U41374 (N_41374,N_37538,N_30470);
xnor U41375 (N_41375,N_32994,N_38156);
or U41376 (N_41376,N_36762,N_36246);
or U41377 (N_41377,N_37712,N_39878);
or U41378 (N_41378,N_31782,N_39022);
and U41379 (N_41379,N_33903,N_31281);
nand U41380 (N_41380,N_35103,N_37815);
nand U41381 (N_41381,N_34369,N_38968);
nor U41382 (N_41382,N_35903,N_37791);
nand U41383 (N_41383,N_37098,N_37571);
nor U41384 (N_41384,N_30650,N_39272);
and U41385 (N_41385,N_38902,N_33688);
or U41386 (N_41386,N_32178,N_33795);
nand U41387 (N_41387,N_33666,N_33513);
nand U41388 (N_41388,N_37306,N_32198);
nand U41389 (N_41389,N_37962,N_34648);
nor U41390 (N_41390,N_38521,N_31611);
and U41391 (N_41391,N_35569,N_36216);
nor U41392 (N_41392,N_35203,N_35473);
xnor U41393 (N_41393,N_32225,N_34690);
nor U41394 (N_41394,N_38716,N_31040);
or U41395 (N_41395,N_31286,N_38774);
nor U41396 (N_41396,N_38470,N_39428);
or U41397 (N_41397,N_37179,N_34693);
nor U41398 (N_41398,N_35061,N_31530);
and U41399 (N_41399,N_39657,N_37350);
or U41400 (N_41400,N_37218,N_39937);
or U41401 (N_41401,N_38157,N_30802);
and U41402 (N_41402,N_36921,N_30064);
or U41403 (N_41403,N_36456,N_32829);
nor U41404 (N_41404,N_36106,N_33147);
nand U41405 (N_41405,N_38921,N_35003);
and U41406 (N_41406,N_33076,N_33836);
xor U41407 (N_41407,N_34106,N_32369);
or U41408 (N_41408,N_38023,N_30027);
nor U41409 (N_41409,N_37882,N_32339);
and U41410 (N_41410,N_36300,N_37994);
and U41411 (N_41411,N_34917,N_37581);
and U41412 (N_41412,N_37182,N_37654);
nor U41413 (N_41413,N_38306,N_37614);
xnor U41414 (N_41414,N_37675,N_30980);
and U41415 (N_41415,N_32347,N_35157);
and U41416 (N_41416,N_31928,N_30171);
nand U41417 (N_41417,N_32383,N_34113);
nand U41418 (N_41418,N_39060,N_30915);
and U41419 (N_41419,N_35120,N_31843);
nor U41420 (N_41420,N_36934,N_35060);
nand U41421 (N_41421,N_36019,N_31795);
nor U41422 (N_41422,N_32489,N_39374);
nand U41423 (N_41423,N_37613,N_39356);
nor U41424 (N_41424,N_37585,N_38329);
nor U41425 (N_41425,N_38114,N_32461);
nand U41426 (N_41426,N_34922,N_36289);
nand U41427 (N_41427,N_31839,N_38351);
nor U41428 (N_41428,N_32978,N_35831);
nor U41429 (N_41429,N_32518,N_37304);
xor U41430 (N_41430,N_31868,N_35146);
or U41431 (N_41431,N_37906,N_32559);
or U41432 (N_41432,N_31743,N_34691);
and U41433 (N_41433,N_37988,N_36491);
nor U41434 (N_41434,N_31048,N_31148);
nand U41435 (N_41435,N_31808,N_34502);
nand U41436 (N_41436,N_35242,N_34993);
and U41437 (N_41437,N_30734,N_33974);
nor U41438 (N_41438,N_30084,N_32191);
or U41439 (N_41439,N_31759,N_35097);
or U41440 (N_41440,N_38184,N_37047);
xor U41441 (N_41441,N_34757,N_36599);
or U41442 (N_41442,N_39397,N_34074);
xnor U41443 (N_41443,N_38617,N_36607);
and U41444 (N_41444,N_38701,N_30025);
or U41445 (N_41445,N_32086,N_38669);
and U41446 (N_41446,N_37983,N_30634);
nor U41447 (N_41447,N_35935,N_38523);
or U41448 (N_41448,N_30139,N_32721);
and U41449 (N_41449,N_39490,N_35550);
xor U41450 (N_41450,N_33463,N_34505);
nor U41451 (N_41451,N_35527,N_32614);
nand U41452 (N_41452,N_37520,N_31584);
nand U41453 (N_41453,N_37603,N_34850);
nor U41454 (N_41454,N_30170,N_30782);
nand U41455 (N_41455,N_32671,N_30202);
nand U41456 (N_41456,N_31482,N_39758);
or U41457 (N_41457,N_32478,N_32460);
and U41458 (N_41458,N_36802,N_33906);
nand U41459 (N_41459,N_31936,N_31738);
and U41460 (N_41460,N_34018,N_32857);
or U41461 (N_41461,N_35720,N_39033);
nor U41462 (N_41462,N_36733,N_32423);
and U41463 (N_41463,N_36143,N_34966);
and U41464 (N_41464,N_34754,N_35629);
or U41465 (N_41465,N_38747,N_34873);
or U41466 (N_41466,N_31225,N_33092);
and U41467 (N_41467,N_39088,N_38986);
nand U41468 (N_41468,N_33852,N_33166);
and U41469 (N_41469,N_30534,N_35426);
nand U41470 (N_41470,N_33602,N_37622);
nand U41471 (N_41471,N_34895,N_33710);
xnor U41472 (N_41472,N_34337,N_31304);
xnor U41473 (N_41473,N_33278,N_34105);
and U41474 (N_41474,N_34198,N_38169);
or U41475 (N_41475,N_31245,N_30689);
and U41476 (N_41476,N_34882,N_37843);
and U41477 (N_41477,N_32638,N_35258);
nor U41478 (N_41478,N_37711,N_33282);
nor U41479 (N_41479,N_39966,N_39179);
and U41480 (N_41480,N_37509,N_37974);
and U41481 (N_41481,N_31468,N_35752);
nor U41482 (N_41482,N_35589,N_36638);
nor U41483 (N_41483,N_33370,N_36559);
and U41484 (N_41484,N_39158,N_30208);
and U41485 (N_41485,N_35755,N_31032);
xnor U41486 (N_41486,N_35035,N_35065);
and U41487 (N_41487,N_38873,N_34776);
nor U41488 (N_41488,N_39813,N_38454);
nand U41489 (N_41489,N_37943,N_31922);
xnor U41490 (N_41490,N_30680,N_34161);
nand U41491 (N_41491,N_33596,N_39288);
or U41492 (N_41492,N_35292,N_30821);
nor U41493 (N_41493,N_30192,N_31564);
and U41494 (N_41494,N_39949,N_34644);
nor U41495 (N_41495,N_32090,N_31344);
or U41496 (N_41496,N_31779,N_31988);
and U41497 (N_41497,N_36121,N_39273);
nand U41498 (N_41498,N_34906,N_39413);
xnor U41499 (N_41499,N_32703,N_35614);
or U41500 (N_41500,N_37329,N_34109);
xnor U41501 (N_41501,N_33469,N_33990);
or U41502 (N_41502,N_32023,N_35055);
or U41503 (N_41503,N_34678,N_37502);
nand U41504 (N_41504,N_34642,N_37485);
nand U41505 (N_41505,N_36305,N_34160);
or U41506 (N_41506,N_36475,N_30519);
or U41507 (N_41507,N_36423,N_33109);
nor U41508 (N_41508,N_31770,N_31865);
and U41509 (N_41509,N_31091,N_33725);
nor U41510 (N_41510,N_37890,N_35306);
or U41511 (N_41511,N_35917,N_31332);
xnor U41512 (N_41512,N_39754,N_30424);
nand U41513 (N_41513,N_39144,N_33427);
xnor U41514 (N_41514,N_36349,N_35023);
nand U41515 (N_41515,N_34069,N_38924);
or U41516 (N_41516,N_34527,N_31716);
and U41517 (N_41517,N_39642,N_32491);
nand U41518 (N_41518,N_35036,N_39222);
and U41519 (N_41519,N_33827,N_33049);
or U41520 (N_41520,N_37213,N_34758);
nor U41521 (N_41521,N_32681,N_33068);
and U41522 (N_41522,N_33178,N_31937);
xor U41523 (N_41523,N_39301,N_32850);
and U41524 (N_41524,N_38682,N_36499);
or U41525 (N_41525,N_38940,N_38974);
and U41526 (N_41526,N_31683,N_38011);
and U41527 (N_41527,N_38599,N_35455);
nand U41528 (N_41528,N_39944,N_33070);
nand U41529 (N_41529,N_32425,N_33646);
or U41530 (N_41530,N_32285,N_37140);
and U41531 (N_41531,N_35858,N_31457);
and U41532 (N_41532,N_33579,N_38745);
or U41533 (N_41533,N_39603,N_31723);
and U41534 (N_41534,N_38609,N_31831);
xnor U41535 (N_41535,N_30968,N_30807);
and U41536 (N_41536,N_30212,N_35087);
nor U41537 (N_41537,N_36674,N_37779);
or U41538 (N_41538,N_33452,N_30733);
nor U41539 (N_41539,N_38007,N_31521);
and U41540 (N_41540,N_31355,N_33761);
or U41541 (N_41541,N_34071,N_30099);
xor U41542 (N_41542,N_37477,N_37919);
xnor U41543 (N_41543,N_33605,N_39664);
or U41544 (N_41544,N_34241,N_30716);
nor U41545 (N_41545,N_34763,N_39174);
and U41546 (N_41546,N_36205,N_37116);
nor U41547 (N_41547,N_35965,N_39747);
nand U41548 (N_41548,N_37224,N_33407);
and U41549 (N_41549,N_39479,N_35944);
nor U41550 (N_41550,N_35861,N_36016);
nor U41551 (N_41551,N_32860,N_34411);
and U41552 (N_41552,N_32641,N_36175);
nor U41553 (N_41553,N_33955,N_31065);
nand U41554 (N_41554,N_30403,N_39203);
nor U41555 (N_41555,N_31650,N_37704);
or U41556 (N_41556,N_30605,N_39750);
and U41557 (N_41557,N_38220,N_31386);
nor U41558 (N_41558,N_39192,N_32700);
or U41559 (N_41559,N_30305,N_32276);
xnor U41560 (N_41560,N_39201,N_38097);
and U41561 (N_41561,N_31253,N_32096);
and U41562 (N_41562,N_38204,N_35828);
nand U41563 (N_41563,N_37417,N_32782);
or U41564 (N_41564,N_34394,N_32768);
and U41565 (N_41565,N_35391,N_33203);
or U41566 (N_41566,N_39573,N_33678);
or U41567 (N_41567,N_37073,N_37798);
or U41568 (N_41568,N_31352,N_32605);
nor U41569 (N_41569,N_37390,N_35685);
nand U41570 (N_41570,N_33369,N_34492);
nor U41571 (N_41571,N_37308,N_32268);
or U41572 (N_41572,N_38292,N_33194);
and U41573 (N_41573,N_37052,N_37319);
or U41574 (N_41574,N_31859,N_35588);
nand U41575 (N_41575,N_39788,N_39299);
or U41576 (N_41576,N_35085,N_38341);
nand U41577 (N_41577,N_34643,N_36597);
xnor U41578 (N_41578,N_33846,N_33317);
nand U41579 (N_41579,N_33188,N_35300);
and U41580 (N_41580,N_37821,N_35279);
xor U41581 (N_41581,N_39286,N_37170);
or U41582 (N_41582,N_34011,N_37252);
nand U41583 (N_41583,N_34884,N_32646);
nand U41584 (N_41584,N_38929,N_30402);
nor U41585 (N_41585,N_35737,N_32222);
nor U41586 (N_41586,N_32833,N_39418);
nand U41587 (N_41587,N_36817,N_35136);
or U41588 (N_41588,N_38266,N_31007);
and U41589 (N_41589,N_31405,N_30247);
nor U41590 (N_41590,N_34338,N_33287);
and U41591 (N_41591,N_31232,N_31319);
or U41592 (N_41592,N_39489,N_38613);
nand U41593 (N_41593,N_36910,N_31440);
nand U41594 (N_41594,N_30115,N_34507);
or U41595 (N_41595,N_37967,N_32713);
nand U41596 (N_41596,N_30829,N_39050);
nand U41597 (N_41597,N_39905,N_33510);
nor U41598 (N_41598,N_33350,N_39960);
nand U41599 (N_41599,N_36745,N_36015);
nand U41600 (N_41600,N_33537,N_39771);
and U41601 (N_41601,N_35893,N_39077);
or U41602 (N_41602,N_35781,N_38881);
or U41603 (N_41603,N_30869,N_30163);
nor U41604 (N_41604,N_39459,N_34980);
nor U41605 (N_41605,N_39981,N_31625);
nand U41606 (N_41606,N_32846,N_32817);
nor U41607 (N_41607,N_38126,N_31910);
nand U41608 (N_41608,N_30110,N_33511);
or U41609 (N_41609,N_32800,N_35398);
xor U41610 (N_41610,N_36966,N_38784);
and U41611 (N_41611,N_38142,N_38104);
and U41612 (N_41612,N_39842,N_31506);
nand U41613 (N_41613,N_31720,N_39599);
nor U41614 (N_41614,N_30220,N_38116);
nor U41615 (N_41615,N_34440,N_38049);
and U41616 (N_41616,N_36576,N_31058);
nand U41617 (N_41617,N_36795,N_32843);
nor U41618 (N_41618,N_37984,N_32684);
nand U41619 (N_41619,N_31401,N_36198);
nand U41620 (N_41620,N_33294,N_38541);
and U41621 (N_41621,N_37859,N_38768);
and U41622 (N_41622,N_38388,N_39576);
nand U41623 (N_41623,N_30270,N_36642);
nor U41624 (N_41624,N_33732,N_34429);
or U41625 (N_41625,N_32451,N_32729);
and U41626 (N_41626,N_39970,N_35453);
and U41627 (N_41627,N_37591,N_30526);
or U41628 (N_41628,N_35829,N_30040);
or U41629 (N_41629,N_33736,N_30827);
or U41630 (N_41630,N_31149,N_37262);
and U41631 (N_41631,N_38147,N_32840);
nand U41632 (N_41632,N_34059,N_36637);
nand U41633 (N_41633,N_32935,N_31288);
nand U41634 (N_41634,N_30043,N_36026);
nor U41635 (N_41635,N_31136,N_31275);
nor U41636 (N_41636,N_33919,N_38070);
nand U41637 (N_41637,N_37287,N_34013);
and U41638 (N_41638,N_32823,N_30707);
or U41639 (N_41639,N_39946,N_32804);
nor U41640 (N_41640,N_38071,N_36825);
or U41641 (N_41641,N_36951,N_36329);
nand U41642 (N_41642,N_39196,N_35027);
nor U41643 (N_41643,N_31657,N_38172);
xnor U41644 (N_41644,N_36828,N_38711);
or U41645 (N_41645,N_34095,N_38103);
nand U41646 (N_41646,N_37535,N_34097);
or U41647 (N_41647,N_34021,N_32674);
nor U41648 (N_41648,N_35921,N_30351);
xor U41649 (N_41649,N_33758,N_30249);
and U41650 (N_41650,N_32900,N_38081);
nand U41651 (N_41651,N_38788,N_37863);
nor U41652 (N_41652,N_38544,N_31321);
xor U41653 (N_41653,N_34163,N_39452);
nand U41654 (N_41654,N_33598,N_38562);
xor U41655 (N_41655,N_37716,N_31051);
nor U41656 (N_41656,N_30196,N_39431);
or U41657 (N_41657,N_37273,N_31951);
and U41658 (N_41658,N_35243,N_34862);
nand U41659 (N_41659,N_33216,N_39170);
nand U41660 (N_41660,N_37523,N_38309);
nand U41661 (N_41661,N_33953,N_34480);
nor U41662 (N_41662,N_39828,N_38377);
and U41663 (N_41663,N_32126,N_30409);
nand U41664 (N_41664,N_36209,N_30258);
xor U41665 (N_41665,N_36875,N_39501);
and U41666 (N_41666,N_36179,N_30999);
nor U41667 (N_41667,N_39407,N_38234);
nand U41668 (N_41668,N_31202,N_33062);
or U41669 (N_41669,N_34303,N_34171);
and U41670 (N_41670,N_38895,N_33119);
nand U41671 (N_41671,N_36766,N_31798);
xnor U41672 (N_41672,N_34704,N_36975);
and U41673 (N_41673,N_38710,N_32582);
nand U41674 (N_41674,N_32779,N_32241);
nor U41675 (N_41675,N_33529,N_34450);
and U41676 (N_41676,N_34592,N_35179);
xnor U41677 (N_41677,N_38775,N_34410);
or U41678 (N_41678,N_36704,N_36892);
or U41679 (N_41679,N_35004,N_33696);
or U41680 (N_41680,N_34531,N_34768);
nor U41681 (N_41681,N_30895,N_30550);
and U41682 (N_41682,N_35726,N_39851);
xnor U41683 (N_41683,N_32544,N_39331);
nor U41684 (N_41684,N_31980,N_38886);
and U41685 (N_41685,N_36654,N_37825);
or U41686 (N_41686,N_38550,N_33105);
and U41687 (N_41687,N_39988,N_31373);
nand U41688 (N_41688,N_32431,N_37030);
and U41689 (N_41689,N_36389,N_39019);
and U41690 (N_41690,N_36557,N_38218);
and U41691 (N_41691,N_39667,N_32937);
or U41692 (N_41692,N_37865,N_38763);
xnor U41693 (N_41693,N_38153,N_38034);
nor U41694 (N_41694,N_37515,N_34900);
or U41695 (N_41695,N_39566,N_33376);
or U41696 (N_41696,N_30123,N_36229);
nor U41697 (N_41697,N_33577,N_30397);
and U41698 (N_41698,N_33096,N_30556);
and U41699 (N_41699,N_36911,N_39053);
nand U41700 (N_41700,N_39717,N_35875);
nand U41701 (N_41701,N_33323,N_30259);
nand U41702 (N_41702,N_39746,N_39293);
nand U41703 (N_41703,N_32774,N_32797);
nor U41704 (N_41704,N_39474,N_35076);
or U41705 (N_41705,N_39440,N_33965);
or U41706 (N_41706,N_35968,N_30642);
or U41707 (N_41707,N_32229,N_33042);
or U41708 (N_41708,N_34477,N_37389);
and U41709 (N_41709,N_38160,N_38296);
nor U41710 (N_41710,N_32839,N_39950);
xor U41711 (N_41711,N_35682,N_38740);
or U41712 (N_41712,N_37626,N_32884);
or U41713 (N_41713,N_34545,N_38373);
or U41714 (N_41714,N_39362,N_34082);
nand U41715 (N_41715,N_38232,N_34459);
or U41716 (N_41716,N_35907,N_36890);
nand U41717 (N_41717,N_39643,N_36669);
and U41718 (N_41718,N_31092,N_39249);
nand U41719 (N_41719,N_33477,N_36227);
nor U41720 (N_41720,N_30062,N_38119);
or U41721 (N_41721,N_39782,N_38508);
nand U41722 (N_41722,N_32752,N_32402);
and U41723 (N_41723,N_31708,N_31949);
and U41724 (N_41724,N_33442,N_30501);
and U41725 (N_41725,N_30013,N_32837);
or U41726 (N_41726,N_36877,N_39213);
and U41727 (N_41727,N_32625,N_33645);
nand U41728 (N_41728,N_37733,N_37305);
or U41729 (N_41729,N_34370,N_37313);
or U41730 (N_41730,N_32253,N_31572);
nand U41731 (N_41731,N_30362,N_34190);
and U41732 (N_41732,N_39436,N_30786);
and U41733 (N_41733,N_37942,N_32092);
nand U41734 (N_41734,N_32123,N_37970);
nor U41735 (N_41735,N_39741,N_36095);
and U41736 (N_41736,N_35645,N_35444);
and U41737 (N_41737,N_31246,N_37746);
or U41738 (N_41738,N_31666,N_37215);
xor U41739 (N_41739,N_37259,N_39233);
nand U41740 (N_41740,N_30651,N_32357);
xor U41741 (N_41741,N_34701,N_34035);
or U41742 (N_41742,N_36429,N_33600);
nand U41743 (N_41743,N_31101,N_37914);
nor U41744 (N_41744,N_37422,N_36231);
xnor U41745 (N_41745,N_34561,N_32271);
and U41746 (N_41746,N_30195,N_34956);
or U41747 (N_41747,N_37745,N_37838);
nor U41748 (N_41748,N_35811,N_39165);
and U41749 (N_41749,N_34567,N_34686);
or U41750 (N_41750,N_34243,N_31117);
nand U41751 (N_41751,N_31737,N_37167);
nand U41752 (N_41752,N_32849,N_36555);
nor U41753 (N_41753,N_32824,N_36366);
nand U41754 (N_41754,N_35347,N_35686);
xnor U41755 (N_41755,N_39243,N_32794);
xnor U41756 (N_41756,N_32987,N_39630);
and U41757 (N_41757,N_32696,N_39621);
or U41758 (N_41758,N_38037,N_36686);
nand U41759 (N_41759,N_39409,N_33797);
nand U41760 (N_41760,N_38657,N_37121);
and U41761 (N_41761,N_35915,N_34902);
or U41762 (N_41762,N_39125,N_31734);
nand U41763 (N_41763,N_32062,N_34064);
nor U41764 (N_41764,N_32373,N_31024);
and U41765 (N_41765,N_33946,N_38757);
or U41766 (N_41766,N_34265,N_35233);
nor U41767 (N_41767,N_30796,N_38196);
or U41768 (N_41768,N_37611,N_39217);
xor U41769 (N_41769,N_35423,N_32158);
nor U41770 (N_41770,N_30889,N_36960);
or U41771 (N_41771,N_38746,N_30173);
and U41772 (N_41772,N_30875,N_32553);
and U41773 (N_41773,N_37540,N_37787);
and U41774 (N_41774,N_32432,N_31772);
nor U41775 (N_41775,N_35435,N_33989);
nand U41776 (N_41776,N_37854,N_32643);
nor U41777 (N_41777,N_34640,N_33494);
nor U41778 (N_41778,N_31421,N_34457);
nand U41779 (N_41779,N_34000,N_35294);
and U41780 (N_41780,N_36109,N_39602);
nor U41781 (N_41781,N_34669,N_37437);
or U41782 (N_41782,N_36925,N_36482);
nand U41783 (N_41783,N_39928,N_36982);
nand U41784 (N_41784,N_33805,N_35934);
or U41785 (N_41785,N_38457,N_34631);
nor U41786 (N_41786,N_37007,N_33196);
or U41787 (N_41787,N_39276,N_30067);
nand U41788 (N_41788,N_37518,N_31522);
and U41789 (N_41789,N_33005,N_33934);
nor U41790 (N_41790,N_32831,N_34145);
nor U41791 (N_41791,N_32876,N_31709);
or U41792 (N_41792,N_30608,N_36080);
nand U41793 (N_41793,N_38195,N_37463);
nor U41794 (N_41794,N_34736,N_30833);
nand U41795 (N_41795,N_37250,N_34330);
and U41796 (N_41796,N_33856,N_37504);
and U41797 (N_41797,N_33689,N_33258);
nor U41798 (N_41798,N_33979,N_30622);
or U41799 (N_41799,N_31697,N_30871);
xnor U41800 (N_41800,N_35834,N_37013);
nor U41801 (N_41801,N_39818,N_38885);
nor U41802 (N_41802,N_32297,N_32939);
nor U41803 (N_41803,N_39429,N_35709);
xor U41804 (N_41804,N_32107,N_30944);
nor U41805 (N_41805,N_32964,N_30215);
and U41806 (N_41806,N_30645,N_38492);
nor U41807 (N_41807,N_33794,N_39366);
xor U41808 (N_41808,N_32195,N_32155);
and U41809 (N_41809,N_30277,N_32676);
nor U41810 (N_41810,N_32571,N_36155);
nor U41811 (N_41811,N_39889,N_35878);
or U41812 (N_41812,N_39312,N_38162);
and U41813 (N_41813,N_31453,N_36528);
nand U41814 (N_41814,N_32224,N_30359);
and U41815 (N_41815,N_36967,N_39461);
nor U41816 (N_41816,N_34673,N_31155);
or U41817 (N_41817,N_31964,N_37596);
and U41818 (N_41818,N_39554,N_37930);
nand U41819 (N_41819,N_37846,N_33399);
nand U41820 (N_41820,N_36708,N_38039);
nor U41821 (N_41821,N_36006,N_32554);
nand U41822 (N_41822,N_35655,N_31179);
nor U41823 (N_41823,N_38455,N_30593);
nor U41824 (N_41824,N_33780,N_31901);
nor U41825 (N_41825,N_39721,N_36053);
or U41826 (N_41826,N_36734,N_32302);
nor U41827 (N_41827,N_34375,N_37801);
and U41828 (N_41828,N_35646,N_39585);
nand U41829 (N_41829,N_30632,N_35665);
and U41830 (N_41830,N_34287,N_30962);
and U41831 (N_41831,N_31711,N_35976);
nand U41832 (N_41832,N_37648,N_39534);
xor U41833 (N_41833,N_38958,N_31769);
xnor U41834 (N_41834,N_39811,N_33378);
or U41835 (N_41835,N_37459,N_30224);
nor U41836 (N_41836,N_38328,N_33555);
xor U41837 (N_41837,N_33333,N_39013);
and U41838 (N_41838,N_34016,N_33809);
xnor U41839 (N_41839,N_37088,N_36813);
or U41840 (N_41840,N_38268,N_30132);
nand U41841 (N_41841,N_32413,N_32007);
nor U41842 (N_41842,N_34124,N_33011);
nand U41843 (N_41843,N_37221,N_34540);
or U41844 (N_41844,N_33309,N_36959);
nor U41845 (N_41845,N_36852,N_31471);
nand U41846 (N_41846,N_30843,N_34500);
nor U41847 (N_41847,N_31822,N_33050);
nor U41848 (N_41848,N_38637,N_37566);
nand U41849 (N_41849,N_36657,N_37019);
nor U41850 (N_41850,N_30779,N_36744);
nand U41851 (N_41851,N_39344,N_31829);
or U41852 (N_41852,N_37297,N_34558);
nand U41853 (N_41853,N_39671,N_37635);
or U41854 (N_41854,N_33150,N_34715);
nor U41855 (N_41855,N_30453,N_34191);
nor U41856 (N_41856,N_31113,N_34447);
xor U41857 (N_41857,N_34044,N_37388);
xor U41858 (N_41858,N_38370,N_33331);
or U41859 (N_41859,N_38131,N_36212);
and U41860 (N_41860,N_33102,N_38136);
and U41861 (N_41861,N_36773,N_39615);
nand U41862 (N_41862,N_33884,N_35274);
nor U41863 (N_41863,N_33130,N_35471);
and U41864 (N_41864,N_31061,N_32172);
xnor U41865 (N_41865,N_30914,N_36760);
nand U41866 (N_41866,N_34172,N_33113);
or U41867 (N_41867,N_32583,N_38033);
and U41868 (N_41868,N_30961,N_33033);
nor U41869 (N_41869,N_37235,N_38277);
and U41870 (N_41870,N_32186,N_30083);
and U41871 (N_41871,N_38183,N_38751);
and U41872 (N_41872,N_35074,N_34353);
or U41873 (N_41873,N_33561,N_36410);
nand U41874 (N_41874,N_34358,N_32925);
nor U41875 (N_41875,N_39876,N_38271);
nor U41876 (N_41876,N_33944,N_38189);
xor U41877 (N_41877,N_37526,N_34995);
and U41878 (N_41878,N_38764,N_31328);
and U41879 (N_41879,N_30293,N_39860);
nor U41880 (N_41880,N_35785,N_39665);
and U41881 (N_41881,N_32440,N_30130);
nand U41882 (N_41882,N_39927,N_35431);
or U41883 (N_41883,N_35885,N_31921);
nor U41884 (N_41884,N_37009,N_31222);
or U41885 (N_41885,N_30094,N_35194);
and U41886 (N_41886,N_35951,N_33763);
nor U41887 (N_41887,N_36851,N_34984);
nand U41888 (N_41888,N_38145,N_38674);
nor U41889 (N_41889,N_36710,N_33127);
nand U41890 (N_41890,N_37248,N_31987);
or U41891 (N_41891,N_34295,N_31174);
and U41892 (N_41892,N_37035,N_30124);
nor U41893 (N_41893,N_34973,N_35758);
nor U41894 (N_41894,N_38483,N_39653);
or U41895 (N_41895,N_31088,N_39466);
or U41896 (N_41896,N_32361,N_32200);
nand U41897 (N_41897,N_30991,N_34712);
xnor U41898 (N_41898,N_31231,N_32454);
and U41899 (N_41899,N_32749,N_32626);
nor U41900 (N_41900,N_35864,N_36180);
nand U41901 (N_41901,N_35591,N_34595);
nor U41902 (N_41902,N_39084,N_38252);
nand U41903 (N_41903,N_37205,N_34015);
nand U41904 (N_41904,N_31807,N_37111);
nand U41905 (N_41905,N_35600,N_37958);
nor U41906 (N_41906,N_32045,N_36608);
nor U41907 (N_41907,N_34938,N_32310);
nor U41908 (N_41908,N_33063,N_37040);
or U41909 (N_41909,N_39685,N_35636);
nand U41910 (N_41910,N_33949,N_30866);
and U41911 (N_41911,N_30011,N_33802);
nor U41912 (N_41912,N_32095,N_33936);
and U41913 (N_41913,N_36069,N_31154);
and U41914 (N_41914,N_31068,N_31277);
and U41915 (N_41915,N_33930,N_30834);
and U41916 (N_41916,N_33128,N_39589);
or U41917 (N_41917,N_38107,N_32205);
or U41918 (N_41918,N_33542,N_30009);
nand U41919 (N_41919,N_31833,N_39986);
nor U41920 (N_41920,N_37106,N_30986);
and U41921 (N_41921,N_31465,N_39419);
nor U41922 (N_41922,N_33234,N_31023);
nand U41923 (N_41923,N_35872,N_39078);
nand U41924 (N_41924,N_35110,N_36104);
or U41925 (N_41925,N_31412,N_34204);
or U41926 (N_41926,N_38344,N_33994);
nor U41927 (N_41927,N_39325,N_32359);
xnor U41928 (N_41928,N_30681,N_38178);
nor U41929 (N_41929,N_31622,N_36884);
and U41930 (N_41930,N_33480,N_37539);
and U41931 (N_41931,N_35754,N_39638);
and U41932 (N_41932,N_33283,N_33037);
or U41933 (N_41933,N_32501,N_34034);
nand U41934 (N_41934,N_30097,N_35337);
nand U41935 (N_41935,N_35395,N_37713);
nor U41936 (N_41936,N_33562,N_31074);
nand U41937 (N_41937,N_36131,N_32303);
nand U41938 (N_41938,N_39742,N_32428);
nand U41939 (N_41939,N_30248,N_37997);
nand U41940 (N_41940,N_39334,N_37848);
or U41941 (N_41941,N_39752,N_36789);
and U41942 (N_41942,N_37345,N_33240);
or U41943 (N_41943,N_39241,N_30636);
nand U41944 (N_41944,N_35764,N_37755);
nand U41945 (N_41945,N_31337,N_32050);
nand U41946 (N_41946,N_34107,N_37639);
nor U41947 (N_41947,N_32673,N_39733);
nor U41948 (N_41948,N_35503,N_31443);
and U41949 (N_41949,N_39391,N_39644);
or U41950 (N_41950,N_37255,N_37058);
and U41951 (N_41951,N_37513,N_35610);
or U41952 (N_41952,N_38061,N_38467);
nor U41953 (N_41953,N_36326,N_39102);
xor U41954 (N_41954,N_39744,N_37327);
nand U41955 (N_41955,N_30928,N_37780);
or U41956 (N_41956,N_39629,N_38581);
or U41957 (N_41957,N_32322,N_31379);
or U41958 (N_41958,N_34996,N_31926);
nor U41959 (N_41959,N_34289,N_34779);
or U41960 (N_41960,N_36998,N_30388);
or U41961 (N_41961,N_34649,N_30736);
nor U41962 (N_41962,N_39708,N_35164);
nor U41963 (N_41963,N_33627,N_33305);
nor U41964 (N_41964,N_38506,N_30822);
xor U41965 (N_41965,N_30404,N_36138);
nand U41966 (N_41966,N_31500,N_32950);
nor U41967 (N_41967,N_36502,N_32647);
and U41968 (N_41968,N_32120,N_39730);
and U41969 (N_41969,N_30683,N_38600);
nand U41970 (N_41970,N_30671,N_34856);
and U41971 (N_41971,N_38058,N_31046);
nand U41972 (N_41972,N_35458,N_32362);
nor U41973 (N_41973,N_30551,N_35508);
nand U41974 (N_41974,N_37627,N_38563);
nand U41975 (N_41975,N_35268,N_33465);
xor U41976 (N_41976,N_39202,N_30221);
and U41977 (N_41977,N_30652,N_38989);
xor U41978 (N_41978,N_36818,N_37275);
nor U41979 (N_41979,N_35007,N_37410);
and U41980 (N_41980,N_31777,N_35501);
and U41981 (N_41981,N_32548,N_33929);
nand U41982 (N_41982,N_31182,N_32005);
nor U41983 (N_41983,N_39416,N_31072);
nor U41984 (N_41984,N_32952,N_39494);
xnor U41985 (N_41985,N_38649,N_34771);
and U41986 (N_41986,N_38164,N_36162);
nor U41987 (N_41987,N_31195,N_34942);
nor U41988 (N_41988,N_31186,N_36883);
or U41989 (N_41989,N_36466,N_38422);
nor U41990 (N_41990,N_39893,N_37738);
nor U41991 (N_41991,N_39441,N_32705);
or U41992 (N_41992,N_33176,N_37904);
nand U41993 (N_41993,N_32666,N_35259);
and U41994 (N_41994,N_35141,N_34635);
or U41995 (N_41995,N_34879,N_30630);
and U41996 (N_41996,N_38614,N_38641);
xor U41997 (N_41997,N_34675,N_36238);
and U41998 (N_41998,N_39898,N_38865);
nand U41999 (N_41999,N_32965,N_32342);
or U42000 (N_42000,N_36893,N_31727);
or U42001 (N_42001,N_37034,N_33267);
nor U42002 (N_42002,N_39881,N_34173);
nor U42003 (N_42003,N_37680,N_34009);
nand U42004 (N_42004,N_32388,N_38583);
or U42005 (N_42005,N_32479,N_32060);
and U42006 (N_42006,N_35121,N_30813);
or U42007 (N_42007,N_33663,N_34553);
or U42008 (N_42008,N_30691,N_35911);
xnor U42009 (N_42009,N_30345,N_36046);
or U42010 (N_42010,N_34585,N_39410);
or U42011 (N_42011,N_32927,N_32877);
xnor U42012 (N_42012,N_34632,N_32510);
and U42013 (N_42013,N_35673,N_33456);
nand U42014 (N_42014,N_33701,N_32955);
or U42015 (N_42015,N_31484,N_35477);
xor U42016 (N_42016,N_37652,N_34967);
nor U42017 (N_42017,N_37326,N_33121);
nor U42018 (N_42018,N_35016,N_34012);
nor U42019 (N_42019,N_37004,N_36091);
and U42020 (N_42020,N_34462,N_36244);
or U42021 (N_42021,N_38298,N_39370);
nor U42022 (N_42022,N_36122,N_35373);
nor U42023 (N_42023,N_34883,N_30309);
nor U42024 (N_42024,N_31520,N_38707);
xor U42025 (N_42025,N_31552,N_31722);
or U42026 (N_42026,N_39696,N_33193);
and U42027 (N_42027,N_38754,N_34749);
nor U42028 (N_42028,N_34555,N_39571);
or U42029 (N_42029,N_30072,N_39871);
nor U42030 (N_42030,N_39411,N_30820);
nand U42031 (N_42031,N_35415,N_36711);
nor U42032 (N_42032,N_30826,N_36358);
or U42033 (N_42033,N_32190,N_30162);
or U42034 (N_42034,N_36151,N_31668);
nor U42035 (N_42035,N_34470,N_36807);
or U42036 (N_42036,N_37681,N_30237);
nand U42037 (N_42037,N_38211,N_39323);
and U42038 (N_42038,N_39844,N_32411);
nor U42039 (N_42039,N_39734,N_37033);
nor U42040 (N_42040,N_36993,N_32669);
xnor U42041 (N_42041,N_36262,N_31119);
or U42042 (N_42042,N_33880,N_38576);
nor U42043 (N_42043,N_39245,N_36876);
or U42044 (N_42044,N_38046,N_31243);
nand U42045 (N_42045,N_39392,N_31900);
and U42046 (N_42046,N_39426,N_33909);
xor U42047 (N_42047,N_37929,N_33030);
or U42048 (N_42048,N_31059,N_32371);
and U42049 (N_42049,N_35365,N_31550);
and U42050 (N_42050,N_34981,N_39464);
xnor U42051 (N_42051,N_36973,N_31085);
xor U42052 (N_42052,N_34668,N_32497);
xor U42053 (N_42053,N_39314,N_36902);
nand U42054 (N_42054,N_33201,N_33383);
nand U42055 (N_42055,N_37100,N_37374);
nand U42056 (N_42056,N_30894,N_34782);
and U42057 (N_42057,N_37318,N_30880);
and U42058 (N_42058,N_31977,N_34169);
nand U42059 (N_42059,N_32320,N_34517);
and U42060 (N_42060,N_32880,N_39359);
xor U42061 (N_42061,N_33551,N_39040);
or U42062 (N_42062,N_36950,N_38120);
nand U42063 (N_42063,N_34032,N_35557);
nand U42064 (N_42064,N_37418,N_36087);
or U42065 (N_42065,N_31904,N_39188);
nand U42066 (N_42066,N_39263,N_31909);
nor U42067 (N_42067,N_39815,N_31301);
or U42068 (N_42068,N_32878,N_36681);
and U42069 (N_42069,N_32892,N_37827);
nor U42070 (N_42070,N_37768,N_32070);
xnor U42071 (N_42071,N_33142,N_37924);
nor U42072 (N_42072,N_37802,N_38067);
nor U42073 (N_42073,N_39663,N_39071);
nor U42074 (N_42074,N_39568,N_34302);
or U42075 (N_42075,N_36297,N_32131);
or U42076 (N_42076,N_34785,N_37811);
nor U42077 (N_42077,N_33855,N_32972);
nor U42078 (N_42078,N_32706,N_38920);
nor U42079 (N_42079,N_32427,N_30923);
nor U42080 (N_42080,N_38489,N_32689);
and U42081 (N_42081,N_34532,N_31832);
nor U42082 (N_42082,N_36301,N_30081);
nand U42083 (N_42083,N_36323,N_31247);
nand U42084 (N_42084,N_38392,N_33754);
and U42085 (N_42085,N_36343,N_36192);
or U42086 (N_42086,N_31027,N_33702);
nor U42087 (N_42087,N_38680,N_34695);
nand U42088 (N_42088,N_34612,N_33160);
or U42089 (N_42089,N_37879,N_32798);
or U42090 (N_42090,N_36070,N_38656);
or U42091 (N_42091,N_30669,N_36929);
xor U42092 (N_42092,N_30850,N_33013);
and U42093 (N_42093,N_34216,N_32109);
xor U42094 (N_42094,N_37303,N_39005);
nand U42095 (N_42095,N_33611,N_34790);
or U42096 (N_42096,N_38854,N_38208);
or U42097 (N_42097,N_30116,N_39640);
and U42098 (N_42098,N_32899,N_38509);
nand U42099 (N_42099,N_36392,N_36147);
or U42100 (N_42100,N_31189,N_37430);
and U42101 (N_42101,N_33172,N_30888);
or U42102 (N_42102,N_35939,N_33189);
or U42103 (N_42103,N_30233,N_33247);
and U42104 (N_42104,N_38358,N_32256);
nor U42105 (N_42105,N_38498,N_31512);
or U42106 (N_42106,N_33348,N_32751);
or U42107 (N_42107,N_37767,N_37575);
or U42108 (N_42108,N_35368,N_37861);
nand U42109 (N_42109,N_35558,N_30376);
nor U42110 (N_42110,N_35449,N_31488);
nor U42111 (N_42111,N_33776,N_39723);
or U42112 (N_42112,N_38025,N_38128);
nor U42113 (N_42113,N_39695,N_35329);
or U42114 (N_42114,N_33760,N_39225);
or U42115 (N_42115,N_35495,N_32750);
or U42116 (N_42116,N_35753,N_31446);
and U42117 (N_42117,N_36324,N_35390);
or U42118 (N_42118,N_34828,N_38123);
nor U42119 (N_42119,N_36972,N_31492);
xnor U42120 (N_42120,N_32393,N_37602);
nand U42121 (N_42121,N_37659,N_30449);
xnor U42122 (N_42122,N_33765,N_37964);
nor U42123 (N_42123,N_36001,N_30485);
nor U42124 (N_42124,N_36408,N_39853);
nand U42125 (N_42125,N_37189,N_30993);
or U42126 (N_42126,N_34616,N_36713);
xor U42127 (N_42127,N_33187,N_37546);
nand U42128 (N_42128,N_34774,N_36420);
and U42129 (N_42129,N_31104,N_32384);
nor U42130 (N_42130,N_36064,N_33650);
and U42131 (N_42131,N_32424,N_34578);
nand U42132 (N_42132,N_30348,N_37484);
xor U42133 (N_42133,N_30801,N_39962);
xnor U42134 (N_42134,N_31028,N_37875);
xnor U42135 (N_42135,N_32717,N_33184);
or U42136 (N_42136,N_30854,N_31680);
nor U42137 (N_42137,N_32258,N_38843);
nand U42138 (N_42138,N_36944,N_33552);
nor U42139 (N_42139,N_36441,N_38004);
and U42140 (N_42140,N_32098,N_32353);
or U42141 (N_42141,N_34414,N_38274);
and U42142 (N_42142,N_39004,N_30491);
or U42143 (N_42143,N_33642,N_37912);
nor U42144 (N_42144,N_34888,N_36378);
nor U42145 (N_42145,N_38095,N_31802);
nor U42146 (N_42146,N_32730,N_33676);
nand U42147 (N_42147,N_38472,N_33090);
nand U42148 (N_42148,N_38231,N_37549);
or U42149 (N_42149,N_38574,N_31356);
nand U42150 (N_42150,N_34787,N_38595);
nor U42151 (N_42151,N_35923,N_31847);
nor U42152 (N_42152,N_32071,N_38858);
nand U42153 (N_42153,N_30858,N_35100);
or U42154 (N_42154,N_33110,N_38675);
nand U42155 (N_42155,N_37754,N_37610);
nand U42156 (N_42156,N_39800,N_36682);
nor U42157 (N_42157,N_36578,N_35695);
and U42158 (N_42158,N_33445,N_33793);
and U42159 (N_42159,N_36547,N_36377);
and U42160 (N_42160,N_32513,N_38249);
or U42161 (N_42161,N_34267,N_36133);
nand U42162 (N_42162,N_32294,N_32228);
nand U42163 (N_42163,N_32784,N_30706);
or U42164 (N_42164,N_30583,N_35432);
xor U42165 (N_42165,N_38807,N_39580);
and U42166 (N_42166,N_36356,N_39834);
nor U42167 (N_42167,N_39789,N_30759);
or U42168 (N_42168,N_31467,N_36161);
or U42169 (N_42169,N_38555,N_38582);
or U42170 (N_42170,N_36062,N_33753);
nand U42171 (N_42171,N_31216,N_38241);
and U42172 (N_42172,N_33826,N_31518);
and U42173 (N_42173,N_30952,N_35291);
or U42174 (N_42174,N_33220,N_32036);
nand U42175 (N_42175,N_32564,N_34449);
and U42176 (N_42176,N_33612,N_36627);
and U42177 (N_42177,N_39228,N_38955);
xnor U42178 (N_42178,N_36632,N_32509);
or U42179 (N_42179,N_36150,N_38411);
nand U42180 (N_42180,N_38300,N_33492);
nor U42181 (N_42181,N_32991,N_32017);
and U42182 (N_42182,N_39700,N_37136);
nand U42183 (N_42183,N_32439,N_37505);
and U42184 (N_42184,N_34897,N_36282);
and U42185 (N_42185,N_34970,N_33007);
nand U42186 (N_42186,N_35380,N_36241);
and U42187 (N_42187,N_36488,N_34100);
nor U42188 (N_42188,N_32307,N_31940);
nor U42189 (N_42189,N_33999,N_39646);
nand U42190 (N_42190,N_39045,N_30989);
nor U42191 (N_42191,N_30355,N_36413);
nor U42192 (N_42192,N_39939,N_35854);
nor U42193 (N_42193,N_30354,N_32199);
and U42194 (N_42194,N_37029,N_38911);
or U42195 (N_42195,N_36619,N_33152);
and U42196 (N_42196,N_35605,N_35772);
or U42197 (N_42197,N_35149,N_30393);
or U42198 (N_42198,N_31796,N_31617);
and U42199 (N_42199,N_39453,N_36038);
nand U42200 (N_42200,N_31640,N_30431);
or U42201 (N_42201,N_38762,N_30268);
nand U42202 (N_42202,N_39727,N_38859);
nor U42203 (N_42203,N_36844,N_36940);
or U42204 (N_42204,N_39305,N_35955);
or U42205 (N_42205,N_33553,N_32720);
xor U42206 (N_42206,N_31766,N_37130);
nand U42207 (N_42207,N_37054,N_38021);
nor U42208 (N_42208,N_38319,N_30350);
or U42209 (N_42209,N_34810,N_35795);
nor U42210 (N_42210,N_35796,N_30805);
or U42211 (N_42211,N_31678,N_32536);
nand U42212 (N_42212,N_33288,N_34559);
or U42213 (N_42213,N_33067,N_30090);
and U42214 (N_42214,N_36014,N_34111);
nand U42215 (N_42215,N_35014,N_38406);
and U42216 (N_42216,N_30420,N_39219);
and U42217 (N_42217,N_34797,N_30904);
and U42218 (N_42218,N_36604,N_33769);
xor U42219 (N_42219,N_30392,N_30262);
or U42220 (N_42220,N_39395,N_36658);
nand U42221 (N_42221,N_34271,N_39252);
or U42222 (N_42222,N_38059,N_30415);
nand U42223 (N_42223,N_30120,N_30271);
nor U42224 (N_42224,N_33118,N_30718);
and U42225 (N_42225,N_37673,N_35954);
nand U42226 (N_42226,N_33747,N_33635);
nand U42227 (N_42227,N_37282,N_35025);
or U42228 (N_42228,N_34285,N_37682);
or U42229 (N_42229,N_33941,N_33655);
or U42230 (N_42230,N_33306,N_39187);
nand U42231 (N_42231,N_35883,N_31674);
and U42232 (N_42232,N_33377,N_38552);
and U42233 (N_42233,N_37544,N_30092);
nand U42234 (N_42234,N_32054,N_30784);
or U42235 (N_42235,N_36743,N_35079);
nand U42236 (N_42236,N_31534,N_30992);
and U42237 (N_42237,N_30471,N_34974);
nor U42238 (N_42238,N_36373,N_39065);
and U42239 (N_42239,N_38654,N_36859);
xnor U42240 (N_42240,N_33563,N_32093);
xor U42241 (N_42241,N_33259,N_37377);
nand U42242 (N_42242,N_39115,N_36145);
or U42243 (N_42243,N_30333,N_30792);
nor U42244 (N_42244,N_33958,N_32692);
and U42245 (N_42245,N_39718,N_38322);
xor U42246 (N_42246,N_32759,N_33004);
nor U42247 (N_42247,N_31371,N_31861);
and U42248 (N_42248,N_34722,N_37871);
nor U42249 (N_42249,N_34940,N_37134);
or U42250 (N_42250,N_38029,N_37857);
and U42251 (N_42251,N_32283,N_32193);
or U42252 (N_42252,N_37129,N_35144);
and U42253 (N_42253,N_31076,N_35707);
nor U42254 (N_42254,N_37314,N_32532);
or U42255 (N_42255,N_37649,N_39755);
nor U42256 (N_42256,N_32985,N_35034);
and U42257 (N_42257,N_31536,N_37979);
nand U42258 (N_42258,N_35051,N_33687);
and U42259 (N_42259,N_32576,N_36754);
and U42260 (N_42260,N_31628,N_34197);
nand U42261 (N_42261,N_37264,N_35326);
nand U42262 (N_42262,N_34731,N_39029);
or U42263 (N_42263,N_37973,N_38722);
nand U42264 (N_42264,N_39859,N_34141);
and U42265 (N_42265,N_30346,N_36587);
or U42266 (N_42266,N_35358,N_30690);
nor U42267 (N_42267,N_34154,N_34461);
nor U42268 (N_42268,N_39854,N_32132);
nand U42269 (N_42269,N_34671,N_32252);
or U42270 (N_42270,N_33023,N_31886);
and U42271 (N_42271,N_33782,N_34184);
xor U42272 (N_42272,N_31172,N_30038);
or U42273 (N_42273,N_36083,N_35874);
nand U42274 (N_42274,N_32760,N_33881);
xnor U42275 (N_42275,N_36072,N_31814);
nand U42276 (N_42276,N_37895,N_31508);
nand U42277 (N_42277,N_35330,N_35734);
xnor U42278 (N_42278,N_34681,N_38078);
or U42279 (N_42279,N_36256,N_37898);
and U42280 (N_42280,N_38642,N_31538);
and U42281 (N_42281,N_32780,N_33403);
and U42282 (N_42282,N_34841,N_35363);
nand U42283 (N_42283,N_38749,N_35033);
nand U42284 (N_42284,N_33100,N_36663);
nand U42285 (N_42285,N_31163,N_39216);
nor U42286 (N_42286,N_31387,N_30988);
nand U42287 (N_42287,N_35219,N_34070);
or U42288 (N_42288,N_39516,N_37005);
and U42289 (N_42289,N_34007,N_32993);
nand U42290 (N_42290,N_37926,N_35299);
nor U42291 (N_42291,N_39529,N_31267);
and U42292 (N_42292,N_32008,N_32115);
or U42293 (N_42293,N_38099,N_36881);
or U42294 (N_42294,N_38366,N_38375);
and U42295 (N_42295,N_37403,N_39508);
and U42296 (N_42296,N_37090,N_37975);
or U42297 (N_42297,N_39185,N_39092);
xor U42298 (N_42298,N_33773,N_32529);
nand U42299 (N_42299,N_39740,N_32592);
nand U42300 (N_42300,N_33652,N_39247);
nand U42301 (N_42301,N_35312,N_36281);
or U42302 (N_42302,N_35698,N_32607);
or U42303 (N_42303,N_34905,N_32930);
nand U42304 (N_42304,N_30891,N_32025);
and U42305 (N_42305,N_34084,N_39607);
or U42306 (N_42306,N_34466,N_35743);
and U42307 (N_42307,N_37978,N_34143);
and U42308 (N_42308,N_38316,N_31660);
nand U42309 (N_42309,N_32913,N_34518);
and U42310 (N_42310,N_34726,N_37276);
nor U42311 (N_42311,N_31260,N_30131);
nand U42312 (N_42312,N_32621,N_33604);
and U42313 (N_42313,N_30823,N_35058);
xor U42314 (N_42314,N_33356,N_35611);
or U42315 (N_42315,N_30971,N_30699);
xnor U42316 (N_42316,N_30773,N_36659);
nand U42317 (N_42317,N_32828,N_38284);
nor U42318 (N_42318,N_35189,N_38364);
xor U42319 (N_42319,N_36316,N_37731);
and U42320 (N_42320,N_36920,N_35517);
or U42321 (N_42321,N_39531,N_31367);
nor U42322 (N_42322,N_37637,N_33597);
or U42323 (N_42323,N_34150,N_39751);
nand U42324 (N_42324,N_37881,N_33046);
nand U42325 (N_42325,N_34036,N_36641);
nor U42326 (N_42326,N_35143,N_31221);
and U42327 (N_42327,N_37923,N_38933);
or U42328 (N_42328,N_31257,N_37340);
nand U42329 (N_42329,N_35445,N_34408);
xor U42330 (N_42330,N_32269,N_33406);
nor U42331 (N_42331,N_35862,N_33161);
and U42332 (N_42332,N_36820,N_36440);
nor U42333 (N_42333,N_31996,N_38695);
nand U42334 (N_42334,N_36294,N_35727);
and U42335 (N_42335,N_32459,N_32111);
xnor U42336 (N_42336,N_37747,N_33168);
xor U42337 (N_42337,N_35563,N_37725);
or U42338 (N_42338,N_36273,N_38922);
nand U42339 (N_42339,N_35640,N_30970);
nor U42340 (N_42340,N_32487,N_33786);
and U42341 (N_42341,N_39460,N_33714);
and U42342 (N_42342,N_38393,N_34800);
and U42343 (N_42343,N_31840,N_35351);
and U42344 (N_42344,N_36066,N_33670);
and U42345 (N_42345,N_33227,N_30075);
xor U42346 (N_42346,N_35671,N_36364);
nor U42347 (N_42347,N_31335,N_38496);
and U42348 (N_42348,N_37705,N_30926);
nor U42349 (N_42349,N_37138,N_36865);
and U42350 (N_42350,N_37383,N_31741);
and U42351 (N_42351,N_32482,N_38150);
nor U42352 (N_42352,N_32181,N_39569);
nand U42353 (N_42353,N_38651,N_32336);
and U42354 (N_42354,N_37886,N_39601);
or U42355 (N_42355,N_39435,N_32226);
nand U42356 (N_42356,N_35174,N_32240);
nand U42357 (N_42357,N_35937,N_30113);
nand U42358 (N_42358,N_39147,N_38887);
xor U42359 (N_42359,N_35188,N_30778);
and U42360 (N_42360,N_39230,N_32437);
nand U42361 (N_42361,N_37972,N_33947);
or U42362 (N_42362,N_30023,N_31384);
nor U42363 (N_42363,N_34444,N_39990);
nor U42364 (N_42364,N_36648,N_30938);
and U42365 (N_42365,N_36649,N_34226);
and U42366 (N_42366,N_34808,N_34872);
and U42367 (N_42367,N_36899,N_35958);
nor U42368 (N_42368,N_39592,N_32956);
nand U42369 (N_42369,N_33312,N_30051);
or U42370 (N_42370,N_37279,N_36846);
or U42371 (N_42371,N_31425,N_39803);
or U42372 (N_42372,N_33217,N_39824);
or U42373 (N_42373,N_39309,N_37137);
or U42374 (N_42374,N_32556,N_35400);
nand U42375 (N_42375,N_34276,N_35624);
or U42376 (N_42376,N_38967,N_35710);
or U42377 (N_42377,N_37547,N_39186);
nor U42378 (N_42378,N_36560,N_39239);
and U42379 (N_42379,N_30505,N_39525);
and U42380 (N_42380,N_37597,N_35725);
and U42381 (N_42381,N_36561,N_34551);
or U42382 (N_42382,N_30190,N_35615);
nor U42383 (N_42383,N_36684,N_34142);
or U42384 (N_42384,N_30808,N_31998);
nand U42385 (N_42385,N_35904,N_35716);
xor U42386 (N_42386,N_31718,N_35568);
and U42387 (N_42387,N_33137,N_36120);
nand U42388 (N_42388,N_32910,N_37234);
nor U42389 (N_42389,N_32758,N_33097);
nor U42390 (N_42390,N_35690,N_37151);
or U42391 (N_42391,N_34728,N_33044);
nand U42392 (N_42392,N_34638,N_38554);
nor U42393 (N_42393,N_31607,N_34954);
nand U42394 (N_42394,N_36028,N_37500);
nor U42395 (N_42395,N_39010,N_33303);
and U42396 (N_42396,N_35765,N_30918);
nor U42397 (N_42397,N_31671,N_34511);
nand U42398 (N_42398,N_31857,N_35548);
and U42399 (N_42399,N_32138,N_31905);
xnor U42400 (N_42400,N_31812,N_34703);
nand U42401 (N_42401,N_38829,N_38978);
nand U42402 (N_42402,N_37773,N_35205);
nor U42403 (N_42403,N_35230,N_38440);
nand U42404 (N_42404,N_37634,N_33806);
nor U42405 (N_42405,N_34274,N_33677);
xnor U42406 (N_42406,N_30973,N_37740);
and U42407 (N_42407,N_38566,N_32040);
and U42408 (N_42408,N_31408,N_38729);
or U42409 (N_42409,N_36339,N_37132);
and U42410 (N_42410,N_30482,N_35472);
nand U42411 (N_42411,N_32018,N_36855);
and U42412 (N_42412,N_30276,N_34118);
and U42413 (N_42413,N_38421,N_34031);
nor U42414 (N_42414,N_36516,N_32210);
nand U42415 (N_42415,N_38008,N_39190);
and U42416 (N_42416,N_36130,N_35542);
and U42417 (N_42417,N_36050,N_34037);
or U42418 (N_42418,N_30211,N_33207);
and U42419 (N_42419,N_36465,N_38620);
and U42420 (N_42420,N_39992,N_35278);
and U42421 (N_42421,N_31237,N_34598);
or U42422 (N_42422,N_35153,N_35162);
nor U42423 (N_42423,N_36081,N_30984);
nand U42424 (N_42424,N_36788,N_31778);
or U42425 (N_42425,N_38053,N_30864);
xnor U42426 (N_42426,N_34813,N_30708);
nand U42427 (N_42427,N_34651,N_35211);
nand U42428 (N_42428,N_38805,N_39911);
nand U42429 (N_42429,N_36645,N_34317);
nor U42430 (N_42430,N_39061,N_33745);
nand U42431 (N_42431,N_36928,N_31437);
xnor U42432 (N_42432,N_38861,N_34928);
nand U42433 (N_42433,N_33409,N_36076);
and U42434 (N_42434,N_38889,N_36152);
nor U42435 (N_42435,N_33238,N_36274);
or U42436 (N_42436,N_35773,N_33723);
or U42437 (N_42437,N_30184,N_30328);
and U42438 (N_42438,N_36864,N_30648);
and U42439 (N_42439,N_38326,N_34503);
xnor U42440 (N_42440,N_31532,N_36248);
nand U42441 (N_42441,N_34255,N_34519);
xor U42442 (N_42442,N_32919,N_34329);
or U42443 (N_42443,N_36311,N_32317);
and U42444 (N_42444,N_35623,N_37197);
nand U42445 (N_42445,N_33252,N_30902);
nor U42446 (N_42446,N_38840,N_39221);
nor U42447 (N_42447,N_39797,N_35982);
nand U42448 (N_42448,N_30783,N_36926);
or U42449 (N_42449,N_33589,N_38338);
or U42450 (N_42450,N_35394,N_31125);
or U42451 (N_42451,N_38828,N_30639);
nand U42452 (N_42452,N_33574,N_36125);
nor U42453 (N_42453,N_36304,N_32350);
nand U42454 (N_42454,N_37092,N_39953);
nor U42455 (N_42455,N_37592,N_38085);
and U42456 (N_42456,N_30957,N_34793);
nand U42457 (N_42457,N_37395,N_35042);
nand U42458 (N_42458,N_36257,N_32035);
nor U42459 (N_42459,N_32091,N_38869);
nand U42460 (N_42460,N_31078,N_33291);
nor U42461 (N_42461,N_37545,N_37824);
or U42462 (N_42462,N_36932,N_31368);
and U42463 (N_42463,N_37584,N_33996);
nand U42464 (N_42464,N_34921,N_30713);
nor U42465 (N_42465,N_39635,N_33618);
or U42466 (N_42466,N_38416,N_32902);
and U42467 (N_42467,N_35303,N_37251);
xnor U42468 (N_42468,N_37321,N_39055);
nand U42469 (N_42469,N_38658,N_37981);
nand U42470 (N_42470,N_35022,N_30450);
nor U42471 (N_42471,N_33503,N_32494);
and U42472 (N_42472,N_38426,N_33219);
and U42473 (N_42473,N_32698,N_33043);
nand U42474 (N_42474,N_31261,N_35116);
nand U42475 (N_42475,N_33896,N_33840);
nand U42476 (N_42476,N_38558,N_32164);
nand U42477 (N_42477,N_30274,N_36841);
nand U42478 (N_42478,N_36532,N_37986);
and U42479 (N_42479,N_39506,N_37661);
and U42480 (N_42480,N_37414,N_33392);
or U42481 (N_42481,N_34762,N_35506);
nor U42482 (N_42482,N_36511,N_32961);
and U42483 (N_42483,N_38330,N_31262);
or U42484 (N_42484,N_32555,N_31473);
nor U42485 (N_42485,N_31917,N_38408);
or U42486 (N_42486,N_32465,N_31916);
and U42487 (N_42487,N_35759,N_31806);
or U42488 (N_42488,N_35941,N_39148);
xor U42489 (N_42489,N_31664,N_38040);
or U42490 (N_42490,N_30284,N_35346);
or U42491 (N_42491,N_39919,N_33789);
xor U42492 (N_42492,N_33864,N_30574);
nand U42493 (N_42493,N_31055,N_31135);
xnor U42494 (N_42494,N_31100,N_36913);
xnor U42495 (N_42495,N_31818,N_34866);
and U42496 (N_42496,N_39998,N_31105);
nand U42497 (N_42497,N_36479,N_35514);
or U42498 (N_42498,N_35377,N_32916);
or U42499 (N_42499,N_32157,N_33693);
nand U42500 (N_42500,N_31785,N_33867);
nand U42501 (N_42501,N_35137,N_30347);
nand U42502 (N_42502,N_38504,N_30655);
or U42503 (N_42503,N_38216,N_35807);
xor U42504 (N_42504,N_31153,N_32498);
or U42505 (N_42505,N_39605,N_38345);
or U42506 (N_42506,N_37595,N_37183);
xnor U42507 (N_42507,N_32490,N_31375);
and U42508 (N_42508,N_35429,N_35545);
or U42509 (N_42509,N_38488,N_36043);
nand U42510 (N_42510,N_30592,N_37902);
nand U42511 (N_42511,N_30824,N_39246);
nand U42512 (N_42512,N_38380,N_37123);
and U42513 (N_42513,N_34494,N_32450);
nor U42514 (N_42514,N_30109,N_35349);
or U42515 (N_42515,N_32922,N_36777);
nor U42516 (N_42516,N_30878,N_38151);
xor U42517 (N_42517,N_36862,N_34982);
and U42518 (N_42518,N_39774,N_31374);
xor U42519 (N_42519,N_31526,N_38585);
and U42520 (N_42520,N_30925,N_30308);
or U42521 (N_42521,N_38559,N_33783);
nor U42522 (N_42522,N_36980,N_32580);
and U42523 (N_42523,N_33943,N_34356);
and U42524 (N_42524,N_38998,N_30029);
nand U42525 (N_42525,N_39952,N_31039);
and U42526 (N_42526,N_39745,N_35089);
or U42527 (N_42527,N_38111,N_39132);
nand U42528 (N_42528,N_33006,N_30881);
nor U42529 (N_42529,N_30314,N_32619);
nor U42530 (N_42530,N_30468,N_36728);
xor U42531 (N_42531,N_33517,N_31860);
nor U42532 (N_42532,N_37514,N_36698);
nand U42533 (N_42533,N_33293,N_35546);
or U42534 (N_42534,N_31623,N_32488);
xor U42535 (N_42535,N_37552,N_32806);
and U42536 (N_42536,N_37270,N_37721);
nand U42537 (N_42537,N_36171,N_30686);
nor U42538 (N_42538,N_39481,N_39829);
or U42539 (N_42539,N_35419,N_33229);
and U42540 (N_42540,N_37936,N_36469);
and U42541 (N_42541,N_30870,N_32105);
or U42542 (N_42542,N_38643,N_39491);
nor U42543 (N_42543,N_39220,N_35794);
and U42544 (N_42544,N_39430,N_30104);
or U42545 (N_42545,N_32505,N_31974);
xor U42546 (N_42546,N_30743,N_38914);
or U42547 (N_42547,N_35325,N_35133);
xor U42548 (N_42548,N_36039,N_35980);
nor U42549 (N_42549,N_31788,N_37479);
and U42550 (N_42550,N_30256,N_35547);
nand U42551 (N_42551,N_30263,N_39079);
nand U42552 (N_42552,N_34520,N_35784);
nand U42553 (N_42553,N_37643,N_37689);
nor U42554 (N_42554,N_35562,N_31757);
or U42555 (N_42555,N_30882,N_39257);
and U42556 (N_42556,N_31903,N_36916);
or U42557 (N_42557,N_34451,N_36500);
nand U42558 (N_42558,N_33681,N_32516);
and U42559 (N_42559,N_30612,N_31050);
nor U42560 (N_42560,N_37524,N_39368);
xnor U42561 (N_42561,N_38822,N_36498);
and U42562 (N_42562,N_38606,N_34554);
and U42563 (N_42563,N_39572,N_36914);
and U42564 (N_42564,N_35165,N_39562);
or U42565 (N_42565,N_30164,N_31164);
and U42566 (N_42566,N_30168,N_38806);
nand U42567 (N_42567,N_30059,N_37331);
nor U42568 (N_42568,N_38254,N_38791);
nor U42569 (N_42569,N_38158,N_38934);
and U42570 (N_42570,N_32377,N_33997);
or U42571 (N_42571,N_37759,N_31749);
nor U42572 (N_42572,N_34230,N_37844);
nor U42573 (N_42573,N_31841,N_32446);
nor U42574 (N_42574,N_36751,N_34269);
nand U42575 (N_42575,N_32118,N_37256);
nand U42576 (N_42576,N_36886,N_39676);
or U42577 (N_42577,N_35360,N_37436);
nor U42578 (N_42578,N_39923,N_34112);
nor U42579 (N_42579,N_32390,N_34589);
xor U42580 (N_42580,N_31311,N_37208);
nor U42581 (N_42581,N_37814,N_31340);
xnor U42582 (N_42582,N_38219,N_39346);
nor U42583 (N_42583,N_39064,N_33286);
nand U42584 (N_42584,N_35000,N_35198);
or U42585 (N_42585,N_33885,N_30435);
and U42586 (N_42586,N_37142,N_31920);
and U42587 (N_42587,N_39686,N_33429);
nor U42588 (N_42588,N_30060,N_32316);
or U42589 (N_42589,N_36357,N_37105);
nor U42590 (N_42590,N_36626,N_33060);
nand U42591 (N_42591,N_35080,N_39181);
nand U42592 (N_42592,N_34080,N_38556);
and U42593 (N_42593,N_30383,N_30585);
nand U42594 (N_42594,N_34992,N_38451);
nor U42595 (N_42595,N_31717,N_30186);
nand U42596 (N_42596,N_38645,N_33830);
or U42597 (N_42597,N_32756,N_34245);
and U42598 (N_42598,N_31686,N_35307);
xnor U42599 (N_42599,N_38833,N_38369);
or U42600 (N_42600,N_38687,N_36220);
nand U42601 (N_42601,N_39885,N_33261);
nor U42602 (N_42602,N_38499,N_31314);
and U42603 (N_42603,N_38778,N_35680);
nand U42604 (N_42604,N_36296,N_32254);
and U42605 (N_42605,N_36473,N_31542);
or U42606 (N_42606,N_37808,N_36874);
nand U42607 (N_42607,N_31187,N_38825);
nor U42608 (N_42608,N_38602,N_38379);
nand U42609 (N_42609,N_39760,N_38233);
nand U42610 (N_42610,N_30809,N_35006);
or U42611 (N_42611,N_32861,N_37233);
and U42612 (N_42612,N_35659,N_31220);
nand U42613 (N_42613,N_33875,N_30253);
or U42614 (N_42614,N_36412,N_31241);
or U42615 (N_42615,N_36832,N_36185);
and U42616 (N_42616,N_32167,N_36584);
and U42617 (N_42617,N_31151,N_39253);
xor U42618 (N_42618,N_37099,N_30654);
and U42619 (N_42619,N_31207,N_36399);
xnor U42620 (N_42620,N_36115,N_37690);
nand U42621 (N_42621,N_34033,N_37809);
or U42622 (N_42622,N_31279,N_38290);
nor U42623 (N_42623,N_33394,N_30214);
or U42624 (N_42624,N_30832,N_35660);
or U42625 (N_42625,N_37894,N_35973);
nand U42626 (N_42626,N_38685,N_37364);
nand U42627 (N_42627,N_30933,N_31956);
and U42628 (N_42628,N_39268,N_34723);
and U42629 (N_42629,N_31191,N_31864);
or U42630 (N_42630,N_33017,N_37036);
and U42631 (N_42631,N_38412,N_38731);
nor U42632 (N_42632,N_35763,N_38365);
or U42633 (N_42633,N_39046,N_30004);
nor U42634 (N_42634,N_34903,N_34657);
nand U42635 (N_42635,N_31213,N_36445);
and U42636 (N_42636,N_31476,N_36991);
and U42637 (N_42637,N_37464,N_37657);
xor U42638 (N_42638,N_32066,N_33036);
and U42639 (N_42639,N_36097,N_32495);
xnor U42640 (N_42640,N_36164,N_36068);
xor U42641 (N_42641,N_39977,N_37669);
or U42642 (N_42642,N_34166,N_35159);
nand U42643 (N_42643,N_36717,N_31932);
nand U42644 (N_42644,N_30146,N_35678);
nand U42645 (N_42645,N_38050,N_31754);
and U42646 (N_42646,N_35910,N_35835);
nor U42647 (N_42647,N_37231,N_35647);
nand U42648 (N_42648,N_32470,N_38855);
and U42649 (N_42649,N_35978,N_35996);
or U42650 (N_42650,N_39054,N_37621);
nand U42651 (N_42651,N_35905,N_37381);
and U42652 (N_42652,N_38491,N_30640);
nand U42653 (N_42653,N_38382,N_32891);
nand U42654 (N_42654,N_39327,N_37373);
nor U42655 (N_42655,N_39389,N_35975);
and U42656 (N_42656,N_35068,N_37045);
or U42657 (N_42657,N_33819,N_33275);
or U42658 (N_42658,N_30906,N_35142);
nor U42659 (N_42659,N_31707,N_33622);
and U42660 (N_42660,N_38750,N_32078);
and U42661 (N_42661,N_32526,N_35930);
nor U42662 (N_42662,N_35151,N_36566);
and U42663 (N_42663,N_34847,N_32333);
or U42664 (N_42664,N_31880,N_31555);
xnor U42665 (N_42665,N_36124,N_33643);
nand U42666 (N_42666,N_33473,N_36431);
nor U42667 (N_42667,N_36572,N_31030);
and U42668 (N_42668,N_37987,N_32675);
or U42669 (N_42669,N_31160,N_35324);
and U42670 (N_42670,N_36931,N_38851);
or U42671 (N_42671,N_36025,N_34564);
or U42672 (N_42672,N_33094,N_30414);
nor U42673 (N_42673,N_35674,N_38547);
or U42674 (N_42674,N_35892,N_31537);
or U42675 (N_42675,N_34699,N_38719);
nand U42676 (N_42676,N_30862,N_37343);
or U42677 (N_42677,N_37608,N_33720);
and U42678 (N_42678,N_33478,N_32561);
nor U42679 (N_42679,N_34076,N_38376);
or U42680 (N_42680,N_31878,N_35639);
nand U42681 (N_42681,N_31240,N_36088);
and U42682 (N_42682,N_31619,N_31855);
or U42683 (N_42683,N_39632,N_32572);
xnor U42684 (N_42684,N_30440,N_30799);
nor U42685 (N_42685,N_32906,N_31961);
or U42686 (N_42686,N_34565,N_34250);
and U42687 (N_42687,N_35168,N_30554);
or U42688 (N_42688,N_35820,N_39394);
and U42689 (N_42689,N_34590,N_32435);
nand U42690 (N_42690,N_38917,N_35622);
nand U42691 (N_42691,N_36427,N_36158);
nor U42692 (N_42692,N_36880,N_34055);
xnor U42693 (N_42693,N_35374,N_30154);
and U42694 (N_42694,N_35138,N_38283);
or U42695 (N_42695,N_33325,N_36401);
and U42696 (N_42696,N_36647,N_37141);
and U42697 (N_42697,N_30201,N_39514);
xnor U42698 (N_42698,N_35790,N_35130);
nand U42699 (N_42699,N_38630,N_38480);
or U42700 (N_42700,N_34426,N_36308);
xnor U42701 (N_42701,N_35019,N_34867);
nand U42702 (N_42702,N_37169,N_38769);
nor U42703 (N_42703,N_39143,N_33641);
nor U42704 (N_42704,N_39502,N_31558);
nand U42705 (N_42705,N_30633,N_39083);
or U42706 (N_42706,N_37177,N_30106);
and U42707 (N_42707,N_36135,N_36478);
or U42708 (N_42708,N_32502,N_36099);
and U42709 (N_42709,N_33431,N_36772);
and U42710 (N_42710,N_39296,N_31914);
nand U42711 (N_42711,N_36183,N_37061);
nand U42712 (N_42712,N_39497,N_32557);
nand U42713 (N_42713,N_35582,N_33346);
nor U42714 (N_42714,N_31852,N_39974);
nand U42715 (N_42715,N_37617,N_33785);
or U42716 (N_42716,N_30619,N_30562);
or U42717 (N_42717,N_30446,N_35840);
or U42718 (N_42718,N_31763,N_37527);
nor U42719 (N_42719,N_35154,N_37089);
nand U42720 (N_42720,N_35946,N_34985);
nor U42721 (N_42721,N_32053,N_34251);
nand U42722 (N_42722,N_38279,N_36785);
or U42723 (N_42723,N_35017,N_33554);
nand U42724 (N_42724,N_34528,N_35064);
xor U42725 (N_42725,N_37618,N_31278);
and U42726 (N_42726,N_31265,N_30598);
nor U42727 (N_42727,N_30898,N_39539);
nand U42728 (N_42728,N_32783,N_38065);
or U42729 (N_42729,N_36439,N_35533);
nor U42730 (N_42730,N_34089,N_35397);
or U42731 (N_42731,N_39873,N_35551);
and U42732 (N_42732,N_38872,N_35037);
and U42733 (N_42733,N_34654,N_33330);
or U42734 (N_42734,N_33202,N_33524);
or U42735 (N_42735,N_37839,N_31108);
nor U42736 (N_42736,N_30464,N_30128);
nor U42737 (N_42737,N_31742,N_39850);
and U42738 (N_42738,N_31123,N_36574);
xor U42739 (N_42739,N_37968,N_39586);
or U42740 (N_42740,N_36678,N_38634);
nand U42741 (N_42741,N_35741,N_33120);
nand U42742 (N_42742,N_32219,N_37743);
and U42743 (N_42743,N_37858,N_34914);
nor U42744 (N_42744,N_36962,N_36368);
and U42745 (N_42745,N_35761,N_37064);
nor U42746 (N_42746,N_32940,N_30659);
nand U42747 (N_42747,N_31098,N_34229);
nor U42748 (N_42748,N_36051,N_34720);
nor U42749 (N_42749,N_31350,N_36422);
nand U42750 (N_42750,N_32245,N_38849);
nor U42751 (N_42751,N_34650,N_36501);
xor U42752 (N_42752,N_34312,N_38635);
nor U42753 (N_42753,N_32265,N_31224);
nand U42754 (N_42754,N_32820,N_33893);
and U42755 (N_42755,N_33523,N_35609);
xor U42756 (N_42756,N_35424,N_36391);
and U42757 (N_42757,N_39138,N_33908);
xnor U42758 (N_42758,N_34907,N_39959);
nand U42759 (N_42759,N_36517,N_37569);
or U42760 (N_42760,N_38794,N_33254);
nor U42761 (N_42761,N_38951,N_32161);
and U42762 (N_42762,N_31912,N_39340);
nand U42763 (N_42763,N_39091,N_38714);
xor U42764 (N_42764,N_32169,N_38994);
and U42765 (N_42765,N_31725,N_34509);
or U42766 (N_42766,N_36938,N_31263);
and U42767 (N_42767,N_35870,N_36907);
nor U42768 (N_42768,N_36653,N_30012);
or U42769 (N_42769,N_33924,N_34588);
nor U42770 (N_42770,N_36333,N_30335);
xor U42771 (N_42771,N_37605,N_36341);
nand U42772 (N_42772,N_34282,N_34887);
xor U42773 (N_42773,N_38870,N_30273);
or U42774 (N_42774,N_38761,N_36679);
and U42775 (N_42775,N_34126,N_33718);
and U42776 (N_42776,N_31228,N_31000);
or U42777 (N_42777,N_38437,N_33708);
or U42778 (N_42778,N_30281,N_37048);
nand U42779 (N_42779,N_39484,N_36577);
and U42780 (N_42780,N_38350,N_30203);
nor U42781 (N_42781,N_36398,N_36791);
xor U42782 (N_42782,N_34472,N_39166);
or U42783 (N_42783,N_30922,N_35308);
or U42784 (N_42784,N_39886,N_31112);
and U42785 (N_42785,N_38098,N_33322);
or U42786 (N_42786,N_38713,N_38188);
or U42787 (N_42787,N_39877,N_32247);
or U42788 (N_42788,N_38076,N_35119);
nand U42789 (N_42789,N_30837,N_30282);
or U42790 (N_42790,N_38520,N_33570);
and U42791 (N_42791,N_32314,N_31582);
nand U42792 (N_42792,N_38952,N_34924);
and U42793 (N_42793,N_36738,N_36061);
and U42794 (N_42794,N_36867,N_34791);
and U42795 (N_42795,N_31513,N_39802);
and U42796 (N_42796,N_37572,N_37537);
xor U42797 (N_42797,N_31199,N_30587);
nand U42798 (N_42798,N_30557,N_30275);
nand U42799 (N_42799,N_33366,N_32364);
and U42800 (N_42800,N_39250,N_38155);
and U42801 (N_42801,N_35296,N_38141);
xnor U42802 (N_42802,N_36763,N_32642);
and U42803 (N_42803,N_32667,N_35090);
or U42804 (N_42804,N_38347,N_35683);
nor U42805 (N_42805,N_38624,N_34372);
and U42806 (N_42806,N_39278,N_38175);
nand U42807 (N_42807,N_33151,N_35254);
xnor U42808 (N_42808,N_39510,N_39902);
or U42809 (N_42809,N_39705,N_38932);
and U42810 (N_42810,N_35045,N_32942);
nor U42811 (N_42811,N_39948,N_33565);
xor U42812 (N_42812,N_33208,N_37473);
nor U42813 (N_42813,N_38224,N_37086);
xor U42814 (N_42814,N_31871,N_31235);
nor U42815 (N_42815,N_35192,N_32872);
and U42816 (N_42816,N_34794,N_30741);
xor U42817 (N_42817,N_33145,N_34378);
or U42818 (N_42818,N_39388,N_33620);
nor U42819 (N_42819,N_35532,N_36335);
or U42820 (N_42820,N_36834,N_34453);
and U42821 (N_42821,N_37147,N_35401);
nor U42822 (N_42822,N_31764,N_39693);
and U42823 (N_42823,N_35687,N_30816);
nor U42824 (N_42824,N_31219,N_38735);
nor U42825 (N_42825,N_37069,N_31563);
nand U42826 (N_42826,N_39238,N_36605);
nand U42827 (N_42827,N_31307,N_35813);
nor U42828 (N_42828,N_32436,N_38629);
and U42829 (N_42829,N_39237,N_30960);
or U42830 (N_42830,N_38242,N_34857);
or U42831 (N_42831,N_33058,N_31324);
nand U42832 (N_42832,N_36606,N_30781);
and U42833 (N_42833,N_33756,N_38311);
xor U42834 (N_42834,N_35869,N_39171);
nor U42835 (N_42835,N_32472,N_31034);
and U42836 (N_42836,N_31685,N_30950);
or U42837 (N_42837,N_39929,N_30752);
and U42838 (N_42838,N_33318,N_39318);
nand U42839 (N_42839,N_33277,N_35800);
xor U42840 (N_42840,N_32058,N_31647);
nand U42841 (N_42841,N_34949,N_39396);
and U42842 (N_42842,N_39207,N_36610);
nand U42843 (N_42843,N_34619,N_37181);
or U42844 (N_42844,N_36860,N_30594);
nand U42845 (N_42845,N_38075,N_35596);
nor U42846 (N_42846,N_30577,N_36319);
nor U42847 (N_42847,N_36830,N_37021);
nor U42848 (N_42848,N_33541,N_33422);
or U42849 (N_42849,N_36983,N_33572);
xor U42850 (N_42850,N_31002,N_32610);
and U42851 (N_42851,N_36706,N_36291);
and U42852 (N_42852,N_33927,N_38077);
xnor U42853 (N_42853,N_38285,N_36588);
and U42854 (N_42854,N_30411,N_36079);
and U42855 (N_42855,N_37670,N_39260);
and U42856 (N_42856,N_35564,N_31957);
nor U42857 (N_42857,N_32594,N_33336);
xor U42858 (N_42858,N_35814,N_34380);
nor U42859 (N_42859,N_34826,N_35579);
nand U42860 (N_42860,N_38121,N_34735);
and U42861 (N_42861,N_32608,N_39381);
or U42862 (N_42862,N_37805,N_31849);
or U42863 (N_42863,N_36618,N_32558);
nand U42864 (N_42864,N_34273,N_34268);
or U42865 (N_42865,N_36058,N_33821);
and U42866 (N_42866,N_35713,N_34941);
nand U42867 (N_42867,N_31474,N_30842);
nand U42868 (N_42868,N_39456,N_31242);
nor U42869 (N_42869,N_32591,N_33700);
nand U42870 (N_42870,N_37562,N_37497);
nand U42871 (N_42871,N_34770,N_31733);
nor U42872 (N_42872,N_36792,N_36462);
or U42873 (N_42873,N_37404,N_35928);
nand U42874 (N_42874,N_31158,N_32870);
nor U42875 (N_42875,N_39725,N_31215);
nand U42876 (N_42876,N_38678,N_33582);
or U42877 (N_42877,N_33025,N_34441);
or U42878 (N_42878,N_32176,N_36470);
xor U42879 (N_42879,N_31941,N_33482);
and U42880 (N_42880,N_30187,N_36670);
nor U42881 (N_42881,N_31823,N_32051);
nor U42882 (N_42882,N_31258,N_35705);
and U42883 (N_42883,N_39847,N_37720);
nand U42884 (N_42884,N_34278,N_30886);
xnor U42885 (N_42885,N_39849,N_30590);
or U42886 (N_42886,N_32699,N_30465);
or U42887 (N_42887,N_35730,N_31439);
nor U42888 (N_42888,N_34894,N_35990);
nand U42889 (N_42889,N_34591,N_37152);
or U42890 (N_42890,N_34885,N_34060);
or U42891 (N_42891,N_34351,N_30087);
nor U42892 (N_42892,N_31712,N_37685);
xnor U42893 (N_42893,N_37732,N_35868);
nand U42894 (N_42894,N_32306,N_38132);
nand U42895 (N_42895,N_34667,N_38459);
xor U42896 (N_42896,N_38400,N_34546);
nor U42897 (N_42897,N_36322,N_37085);
and U42898 (N_42898,N_33487,N_37193);
and U42899 (N_42899,N_35362,N_33505);
and U42900 (N_42900,N_34557,N_38022);
or U42901 (N_42901,N_30663,N_31018);
or U42902 (N_42902,N_39577,N_33932);
nand U42903 (N_42903,N_38598,N_32076);
and U42904 (N_42904,N_33024,N_33992);
nor U42905 (N_42905,N_35156,N_36387);
nor U42906 (N_42906,N_36879,N_37579);
nand U42907 (N_42907,N_34357,N_31475);
or U42908 (N_42908,N_30467,N_39235);
nor U42909 (N_42909,N_35953,N_38149);
nor U42910 (N_42910,N_31481,N_36507);
nor U42911 (N_42911,N_30353,N_37229);
xor U42912 (N_42912,N_31204,N_32278);
nand U42913 (N_42913,N_35961,N_34318);
or U42914 (N_42914,N_39887,N_34838);
and U42915 (N_42915,N_33521,N_34617);
nand U42916 (N_42916,N_38244,N_30200);
nand U42917 (N_42917,N_31458,N_30600);
xor U42918 (N_42918,N_30530,N_30389);
and U42919 (N_42919,N_33245,N_37202);
or U42920 (N_42920,N_37783,N_33421);
and U42921 (N_42921,N_39924,N_31400);
and U42922 (N_42922,N_31654,N_32137);
and U42923 (N_42923,N_34277,N_33347);
nand U42924 (N_42924,N_37103,N_33824);
xnor U42925 (N_42925,N_38918,N_32016);
or U42926 (N_42926,N_39512,N_38625);
nand U42927 (N_42927,N_36748,N_32043);
and U42928 (N_42928,N_36251,N_30156);
nor U42929 (N_42929,N_34729,N_32988);
nand U42930 (N_42930,N_31208,N_35434);
nand U42931 (N_42931,N_31223,N_32602);
xor U42932 (N_42932,N_37679,N_36092);
nor U42933 (N_42933,N_35505,N_35694);
nand U42934 (N_42934,N_37708,N_30674);
xnor U42935 (N_42935,N_37087,N_35779);
or U42936 (N_42936,N_38667,N_34264);
and U42937 (N_42937,N_33424,N_31354);
or U42938 (N_42938,N_33373,N_31679);
nand U42939 (N_42939,N_39852,N_38681);
nand U42940 (N_42940,N_39677,N_30874);
and U42941 (N_42941,N_33486,N_34968);
and U42942 (N_42942,N_30836,N_35703);
nand U42943 (N_42943,N_37883,N_33774);
nor U42944 (N_42944,N_38462,N_30444);
nand U42945 (N_42945,N_36552,N_38384);
or U42946 (N_42946,N_37781,N_33021);
nor U42947 (N_42947,N_31329,N_31528);
or U42948 (N_42948,N_38171,N_39218);
or U42949 (N_42949,N_30144,N_36351);
or U42950 (N_42950,N_37842,N_37023);
nand U42951 (N_42951,N_33112,N_33734);
and U42952 (N_42952,N_39918,N_37050);
and U42953 (N_42953,N_30873,N_38246);
nand U42954 (N_42954,N_37847,N_37667);
or U42955 (N_42955,N_36586,N_33993);
and U42956 (N_42956,N_36812,N_35669);
and U42957 (N_42957,N_30000,N_39588);
nor U42958 (N_42958,N_38227,N_33925);
or U42959 (N_42959,N_34610,N_37920);
xnor U42960 (N_42960,N_37195,N_30050);
nor U42961 (N_42961,N_32981,N_33913);
and U42962 (N_42962,N_37961,N_37819);
nand U42963 (N_42963,N_34933,N_36370);
or U42964 (N_42964,N_30924,N_37342);
nor U42965 (N_42965,N_30955,N_35574);
or U42966 (N_42966,N_30443,N_35163);
xnor U42967 (N_42967,N_36918,N_31690);
nor U42968 (N_42968,N_34165,N_35670);
nand U42969 (N_42969,N_36367,N_30722);
or U42970 (N_42970,N_32345,N_31392);
nand U42971 (N_42971,N_31370,N_32237);
or U42972 (N_42972,N_39372,N_30609);
and U42973 (N_42973,N_39595,N_37730);
nand U42974 (N_42974,N_32541,N_37001);
and U42975 (N_42975,N_39866,N_32863);
nand U42976 (N_42976,N_30140,N_37072);
or U42977 (N_42977,N_33453,N_37157);
and U42978 (N_42978,N_35280,N_34625);
nand U42979 (N_42979,N_37900,N_38230);
nor U42980 (N_42980,N_32175,N_35597);
nand U42981 (N_42981,N_34724,N_36954);
and U42982 (N_42982,N_33810,N_39899);
and U42983 (N_42983,N_35239,N_38259);
or U42984 (N_42984,N_39204,N_30330);
and U42985 (N_42985,N_31297,N_30103);
or U42986 (N_42986,N_35523,N_39017);
nand U42987 (N_42987,N_30732,N_37891);
nor U42988 (N_42988,N_33831,N_33344);
nand U42989 (N_42989,N_34498,N_35059);
nand U42990 (N_42990,N_31418,N_30703);
or U42991 (N_42991,N_37496,N_32629);
xnor U42992 (N_42992,N_39049,N_32097);
nand U42993 (N_42993,N_36997,N_33583);
or U42994 (N_42994,N_39306,N_37060);
and U42995 (N_42995,N_39804,N_34806);
nor U42996 (N_42996,N_33361,N_39967);
nor U42997 (N_42997,N_30357,N_38263);
nand U42998 (N_42998,N_35801,N_36634);
nor U42999 (N_42999,N_37315,N_33443);
nand U43000 (N_43000,N_30489,N_37380);
nand U43001 (N_43001,N_33709,N_39897);
or U43002 (N_43002,N_39424,N_31469);
nor U43003 (N_43003,N_34061,N_38458);
nor U43004 (N_43004,N_32318,N_32360);
nand U43005 (N_43005,N_36527,N_39656);
nor U43006 (N_43006,N_37845,N_30977);
and U43007 (N_43007,N_35500,N_32928);
nor U43008 (N_43008,N_33522,N_38490);
nor U43009 (N_43009,N_32202,N_35369);
or U43010 (N_43010,N_31494,N_32069);
nand U43011 (N_43011,N_34176,N_34575);
nand U43012 (N_43012,N_31944,N_37662);
and U43013 (N_43013,N_30508,N_31236);
nor U43014 (N_43014,N_37271,N_30071);
and U43015 (N_43015,N_36239,N_30610);
and U43016 (N_43016,N_39200,N_38403);
nor U43017 (N_43017,N_33069,N_35776);
nor U43018 (N_43018,N_30510,N_39096);
nor U43019 (N_43019,N_39496,N_39104);
or U43020 (N_43020,N_35957,N_39681);
and U43021 (N_43021,N_39042,N_39943);
and U43022 (N_43022,N_30867,N_31198);
and U43023 (N_43023,N_30199,N_30143);
and U43024 (N_43024,N_34536,N_34839);
and U43025 (N_43025,N_31665,N_36102);
xor U43026 (N_43026,N_35581,N_30303);
or U43027 (N_43027,N_37699,N_31141);
nor U43028 (N_43028,N_37299,N_30740);
or U43029 (N_43029,N_38199,N_33515);
and U43030 (N_43030,N_37425,N_36544);
nor U43031 (N_43031,N_31444,N_39784);
nor U43032 (N_43032,N_33297,N_37439);
nor U43033 (N_43033,N_37245,N_38708);
or U43034 (N_43034,N_36250,N_39449);
or U43035 (N_43035,N_36646,N_30540);
nand U43036 (N_43036,N_33738,N_37786);
and U43037 (N_43037,N_37917,N_31781);
and U43038 (N_43038,N_36266,N_36332);
nor U43039 (N_43039,N_37977,N_31761);
and U43040 (N_43040,N_37465,N_35109);
or U43041 (N_43041,N_33706,N_30751);
nor U43042 (N_43042,N_32246,N_33458);
nor U43043 (N_43043,N_31971,N_31973);
nand U43044 (N_43044,N_37590,N_32356);
or U43045 (N_43045,N_32665,N_31041);
nand U43046 (N_43046,N_32102,N_37346);
nand U43047 (N_43047,N_33538,N_32326);
nand U43048 (N_43048,N_30927,N_30056);
or U43049 (N_43049,N_33425,N_37644);
and U43050 (N_43050,N_32162,N_30058);
nor U43051 (N_43051,N_33475,N_32282);
and U43052 (N_43052,N_38387,N_38905);
nand U43053 (N_43053,N_31006,N_33470);
and U43054 (N_43054,N_31562,N_34151);
nand U43055 (N_43055,N_31133,N_32400);
nand U43056 (N_43056,N_34397,N_31416);
nor U43057 (N_43057,N_37280,N_34751);
or U43058 (N_43058,N_35234,N_33273);
and U43059 (N_43059,N_30487,N_35888);
nor U43060 (N_43060,N_34422,N_37774);
nand U43061 (N_43061,N_34822,N_30265);
xor U43062 (N_43062,N_37561,N_33502);
and U43063 (N_43063,N_36362,N_37442);
xor U43064 (N_43064,N_34861,N_31990);
nor U43065 (N_43065,N_32295,N_30604);
nand U43066 (N_43066,N_33134,N_33272);
xor U43067 (N_43067,N_34157,N_39555);
nor U43068 (N_43068,N_30042,N_34464);
xnor U43069 (N_43069,N_31393,N_33832);
nor U43070 (N_43070,N_34816,N_36187);
nand U43071 (N_43071,N_35922,N_39697);
xor U43072 (N_43072,N_33751,N_33869);
or U43073 (N_43073,N_33987,N_37869);
and U43074 (N_43074,N_36676,N_32776);
or U43075 (N_43075,N_33485,N_35715);
and U43076 (N_43076,N_31339,N_33508);
nand U43077 (N_43077,N_34202,N_38736);
and U43078 (N_43078,N_39355,N_33124);
nor U43079 (N_43079,N_36004,N_31609);
nor U43080 (N_43080,N_39458,N_37017);
nor U43081 (N_43081,N_30597,N_33975);
nand U43082 (N_43082,N_33398,N_37831);
nor U43083 (N_43083,N_36600,N_36757);
and U43084 (N_43084,N_35145,N_39965);
and U43085 (N_43085,N_34804,N_36771);
or U43086 (N_43086,N_33326,N_37955);
nand U43087 (N_43087,N_39455,N_38047);
or U43088 (N_43088,N_36888,N_38821);
and U43089 (N_43089,N_32765,N_30283);
nor U43090 (N_43090,N_39810,N_33528);
nor U43091 (N_43091,N_31289,N_39836);
or U43092 (N_43092,N_38190,N_32827);
xnor U43093 (N_43093,N_33560,N_31082);
nand U43094 (N_43094,N_31029,N_32995);
xnor U43095 (N_43095,N_36265,N_30814);
or U43096 (N_43096,N_30618,N_39130);
and U43097 (N_43097,N_30459,N_38945);
or U43098 (N_43098,N_30819,N_31803);
or U43099 (N_43099,N_37480,N_38743);
nor U43100 (N_43100,N_37184,N_35212);
or U43101 (N_43101,N_36298,N_38797);
nor U43102 (N_43102,N_35770,N_38668);
or U43103 (N_43103,N_32552,N_31877);
and U43104 (N_43104,N_34824,N_33539);
xnor U43105 (N_43105,N_31188,N_32545);
nor U43106 (N_43106,N_37301,N_31639);
nor U43107 (N_43107,N_36799,N_37491);
xor U43108 (N_43108,N_35328,N_39316);
nor U43109 (N_43109,N_34398,N_31989);
xnor U43110 (N_43110,N_30818,N_31982);
and U43111 (N_43111,N_35436,N_39119);
or U43112 (N_43112,N_36564,N_33981);
xor U43113 (N_43113,N_38993,N_30520);
nor U43114 (N_43114,N_30167,N_32542);
and U43115 (N_43115,N_35625,N_36520);
or U43116 (N_43116,N_33812,N_32851);
or U43117 (N_43117,N_34773,N_31276);
nor U43118 (N_43118,N_33616,N_30539);
nor U43119 (N_43119,N_36474,N_36824);
nand U43120 (N_43120,N_39423,N_37370);
or U43121 (N_43121,N_33985,N_37091);
and U43122 (N_43122,N_39405,N_30065);
or U43123 (N_43123,N_38572,N_39390);
nor U43124 (N_43124,N_36100,N_34266);
and U43125 (N_43125,N_36595,N_39994);
nand U43126 (N_43126,N_32273,N_31445);
or U43127 (N_43127,N_39375,N_31441);
or U43128 (N_43128,N_38036,N_34231);
and U43129 (N_43129,N_38936,N_35728);
or U43130 (N_43130,N_31227,N_37769);
nor U43131 (N_43131,N_34795,N_34164);
xnor U43132 (N_43132,N_39812,N_32065);
nand U43133 (N_43133,N_36702,N_32032);
xnor U43134 (N_43134,N_37332,N_30205);
or U43135 (N_43135,N_37237,N_30082);
or U43136 (N_43136,N_38997,N_35343);
or U43137 (N_43137,N_36114,N_34301);
nand U43138 (N_43138,N_36247,N_30595);
and U43139 (N_43139,N_33413,N_32063);
nor U43140 (N_43140,N_32449,N_35947);
nor U43141 (N_43141,N_39290,N_33411);
and U43142 (N_43142,N_38592,N_30811);
nand U43143 (N_43143,N_39254,N_33250);
nor U43144 (N_43144,N_38331,N_38703);
nor U43145 (N_43145,N_35468,N_32514);
nor U43146 (N_43146,N_38209,N_30724);
nand U43147 (N_43147,N_35766,N_36919);
and U43148 (N_43148,N_37966,N_31575);
and U43149 (N_43149,N_32009,N_32848);
nand U43150 (N_43150,N_35293,N_33784);
nand U43151 (N_43151,N_37804,N_34877);
and U43152 (N_43152,N_35399,N_35147);
and U43153 (N_43153,N_38699,N_33849);
nor U43154 (N_43154,N_30777,N_30509);
nor U43155 (N_43155,N_31801,N_35333);
and U43156 (N_43156,N_31689,N_37908);
nand U43157 (N_43157,N_38449,N_35635);
nor U43158 (N_43158,N_37829,N_34178);
and U43159 (N_43159,N_39208,N_31630);
or U43160 (N_43160,N_38276,N_35793);
nand U43161 (N_43161,N_35106,N_33898);
nand U43162 (N_43162,N_35531,N_35575);
xnor U43163 (N_43163,N_39121,N_32030);
and U43164 (N_43164,N_31691,N_35072);
or U43165 (N_43165,N_32209,N_33657);
or U43166 (N_43166,N_36521,N_38396);
nand U43167 (N_43167,N_36464,N_36169);
nor U43168 (N_43168,N_37261,N_39403);
nor U43169 (N_43169,N_32171,N_36224);
nor U43170 (N_43170,N_35364,N_30662);
nor U43171 (N_43171,N_33726,N_38217);
and U43172 (N_43172,N_35316,N_34606);
nor U43173 (N_43173,N_31298,N_39735);
and U43174 (N_43174,N_38856,N_30705);
nand U43175 (N_43175,N_31169,N_38096);
xor U43176 (N_43176,N_38336,N_37355);
or U43177 (N_43177,N_34320,N_36963);
or U43178 (N_43178,N_34738,N_32272);
nand U43179 (N_43179,N_37790,N_31413);
and U43180 (N_43180,N_37120,N_37631);
and U43181 (N_43181,N_31881,N_38960);
nor U43182 (N_43182,N_31256,N_34964);
xnor U43183 (N_43183,N_31879,N_31442);
nor U43184 (N_43184,N_34339,N_33301);
nor U43185 (N_43185,N_37003,N_33851);
or U43186 (N_43186,N_35684,N_35632);
nor U43187 (N_43187,N_38738,N_35140);
or U43188 (N_43188,N_34463,N_30108);
nand U43189 (N_43189,N_32838,N_33103);
nor U43190 (N_43190,N_32447,N_30222);
and U43191 (N_43191,N_37281,N_35171);
xor U43192 (N_43192,N_37724,N_32290);
nor U43193 (N_43193,N_32519,N_31353);
nand U43194 (N_43194,N_33733,N_35093);
nor U43195 (N_43195,N_30278,N_37322);
nand U43196 (N_43196,N_39703,N_32854);
and U43197 (N_43197,N_36320,N_34727);
xnor U43198 (N_43198,N_30678,N_31835);
or U43199 (N_43199,N_36714,N_37062);
or U43200 (N_43200,N_30374,N_33959);
nand U43201 (N_43201,N_39608,N_39363);
or U43202 (N_43202,N_32277,N_30997);
nand U43203 (N_43203,N_38812,N_32249);
and U43204 (N_43204,N_30982,N_36908);
or U43205 (N_43205,N_30191,N_35805);
and U43206 (N_43206,N_37269,N_38831);
nor U43207 (N_43207,N_35656,N_39931);
or U43208 (N_43208,N_30179,N_36290);
nand U43209 (N_43209,N_31756,N_32596);
nand U43210 (N_43210,N_32593,N_30475);
nor U43211 (N_43211,N_38381,N_35167);
and U43212 (N_43212,N_37117,N_39002);
nand U43213 (N_43213,N_37260,N_34443);
xor U43214 (N_43214,N_31402,N_32180);
nand U43215 (N_43215,N_36758,N_38083);
nand U43216 (N_43216,N_35987,N_37950);
nand U43217 (N_43217,N_30697,N_32134);
nand U43218 (N_43218,N_35571,N_33276);
xor U43219 (N_43219,N_38324,N_31495);
or U43220 (N_43220,N_36996,N_37971);
nand U43221 (N_43221,N_37490,N_34904);
xor U43222 (N_43222,N_36086,N_34348);
and U43223 (N_43223,N_34501,N_38090);
and U43224 (N_43224,N_33639,N_38320);
nand U43225 (N_43225,N_34582,N_30323);
xor U43226 (N_43226,N_34403,N_33059);
nor U43227 (N_43227,N_39660,N_31959);
nand U43228 (N_43228,N_38548,N_33419);
or U43229 (N_43229,N_39066,N_35114);
nor U43230 (N_43230,N_31094,N_32651);
and U43231 (N_43231,N_38662,N_30280);
nand U43232 (N_43232,N_31693,N_33640);
xnor U43233 (N_43233,N_39958,N_31226);
and U43234 (N_43234,N_38362,N_32047);
and U43235 (N_43235,N_38414,N_36055);
and U43236 (N_43236,N_35631,N_31876);
or U43237 (N_43237,N_34039,N_34939);
nor U43238 (N_43238,N_31786,N_32825);
and U43239 (N_43239,N_38798,N_30893);
nor U43240 (N_43240,N_30472,N_33434);
and U43241 (N_43241,N_32103,N_39972);
or U43242 (N_43242,N_34929,N_31592);
nand U43243 (N_43243,N_35842,N_30755);
or U43244 (N_43244,N_36459,N_39152);
nand U43245 (N_43245,N_32733,N_30061);
or U43246 (N_43246,N_34514,N_33633);
nor U43247 (N_43247,N_39549,N_33807);
nor U43248 (N_43248,N_36697,N_31129);
xnor U43249 (N_43249,N_34664,N_38337);
nand U43250 (N_43250,N_31981,N_33263);
nor U43251 (N_43251,N_38838,N_30197);
or U43252 (N_43252,N_39360,N_35195);
or U43253 (N_43253,N_37356,N_38903);
nand U43254 (N_43254,N_31464,N_36040);
or U43255 (N_43255,N_39343,N_31699);
nor U43256 (N_43256,N_35492,N_36784);
nor U43257 (N_43257,N_36259,N_35244);
nand U43258 (N_43258,N_39537,N_34040);
or U43259 (N_43259,N_32691,N_33395);
or U43260 (N_43260,N_34878,N_35054);
nor U43261 (N_43261,N_36200,N_35009);
nand U43262 (N_43262,N_31296,N_33978);
nor U43263 (N_43263,N_39434,N_34156);
xnor U43264 (N_43264,N_32739,N_37344);
nor U43265 (N_43265,N_30390,N_36948);
nor U43266 (N_43266,N_30900,N_39020);
nor U43267 (N_43267,N_32787,N_37423);
nand U43268 (N_43268,N_36434,N_38908);
nor U43269 (N_43269,N_37744,N_39070);
xnor U43270 (N_43270,N_30054,N_31410);
and U43271 (N_43271,N_36988,N_39513);
and U43272 (N_43272,N_37113,N_38551);
nand U43273 (N_43273,N_32300,N_31461);
or U43274 (N_43274,N_33729,N_38640);
and U43275 (N_43275,N_37941,N_38930);
or U43276 (N_43276,N_38243,N_37387);
and U43277 (N_43277,N_39597,N_34566);
or U43278 (N_43278,N_37849,N_39076);
and U43279 (N_43279,N_35043,N_37985);
and U43280 (N_43280,N_38835,N_33304);
nand U43281 (N_43281,N_37066,N_30558);
and U43282 (N_43282,N_35846,N_31218);
nand U43283 (N_43283,N_38182,N_31509);
nand U43284 (N_43284,N_34991,N_38144);
nand U43285 (N_43285,N_38240,N_38785);
or U43286 (N_43286,N_36047,N_32286);
nand U43287 (N_43287,N_39378,N_38173);
or U43288 (N_43288,N_33507,N_39123);
nor U43289 (N_43289,N_35161,N_30753);
and U43290 (N_43290,N_37450,N_34753);
or U43291 (N_43291,N_38010,N_30553);
nor U43292 (N_43292,N_38177,N_34702);
nor U43293 (N_43293,N_38628,N_30694);
nor U43294 (N_43294,N_32215,N_32612);
nand U43295 (N_43295,N_37922,N_38297);
nand U43296 (N_43296,N_35721,N_38516);
nor U43297 (N_43297,N_36543,N_34412);
nand U43298 (N_43298,N_36985,N_37097);
and U43299 (N_43299,N_34364,N_32766);
nor U43300 (N_43300,N_38888,N_38505);
nor U43301 (N_43301,N_32352,N_35304);
nor U43302 (N_43302,N_30111,N_31044);
or U43303 (N_43303,N_31316,N_35383);
or U43304 (N_43304,N_34332,N_37928);
and U43305 (N_43305,N_32767,N_36787);
xnor U43306 (N_43306,N_31205,N_31239);
nand U43307 (N_43307,N_32116,N_37083);
and U43308 (N_43308,N_35877,N_36042);
nand U43309 (N_43309,N_33516,N_36898);
and U43310 (N_43310,N_31110,N_38106);
and U43311 (N_43311,N_34661,N_34340);
nand U43312 (N_43312,N_37841,N_34628);
or U43313 (N_43313,N_33444,N_32999);
and U43314 (N_43314,N_39469,N_30299);
nor U43315 (N_43315,N_38543,N_32953);
nand U43316 (N_43316,N_36117,N_33621);
or U43317 (N_43317,N_31667,N_35448);
nor U43318 (N_43318,N_34362,N_30260);
and U43319 (N_43319,N_38100,N_35113);
nor U43320 (N_43320,N_32387,N_33755);
and U43321 (N_43321,N_35997,N_36614);
and U43322 (N_43322,N_35414,N_33035);
xnor U43323 (N_43323,N_30216,N_38773);
nand U43324 (N_43324,N_31652,N_35739);
and U43325 (N_43325,N_32777,N_32220);
nor U43326 (N_43326,N_37642,N_33125);
nor U43327 (N_43327,N_35832,N_38301);
and U43328 (N_43328,N_34515,N_38127);
nor U43329 (N_43329,N_30266,N_32525);
or U43330 (N_43330,N_36029,N_33581);
nor U43331 (N_43331,N_37578,N_35512);
nand U43332 (N_43332,N_38928,N_31724);
or U43333 (N_43333,N_32601,N_35493);
nor U43334 (N_43334,N_32810,N_31967);
nor U43335 (N_43335,N_37577,N_39486);
nand U43336 (N_43336,N_36344,N_34522);
nor U43337 (N_43337,N_32346,N_34777);
or U43338 (N_43338,N_33162,N_31675);
and U43339 (N_43339,N_32795,N_39332);
nor U43340 (N_43340,N_33877,N_37775);
nor U43341 (N_43341,N_31760,N_30711);
nor U43342 (N_43342,N_38028,N_34697);
nor U43343 (N_43343,N_30670,N_37203);
nor U43344 (N_43344,N_31968,N_31052);
nand U43345 (N_43345,N_34543,N_30514);
and U43346 (N_43346,N_32108,N_31748);
nor U43347 (N_43347,N_30507,N_35981);
or U43348 (N_43348,N_38815,N_32637);
nor U43349 (N_43349,N_37498,N_33504);
xor U43350 (N_43350,N_31701,N_34117);
xor U43351 (N_43351,N_39520,N_39289);
and U43352 (N_43352,N_36570,N_31978);
or U43353 (N_43353,N_33592,N_37026);
nand U43354 (N_43354,N_33027,N_32639);
nand U43355 (N_43355,N_38401,N_33001);
or U43356 (N_43356,N_30942,N_39995);
or U43357 (N_43357,N_32130,N_33104);
nor U43358 (N_43358,N_36946,N_34547);
nand U43359 (N_43359,N_31649,N_35479);
nor U43360 (N_43360,N_38772,N_34920);
nor U43361 (N_43361,N_38638,N_37530);
or U43362 (N_43362,N_38565,N_34739);
nand U43363 (N_43363,N_39612,N_36360);
nand U43364 (N_43364,N_30861,N_31312);
and U43365 (N_43365,N_35344,N_30386);
and U43366 (N_43366,N_32598,N_34948);
nand U43367 (N_43367,N_38718,N_38122);
nand U43368 (N_43368,N_39906,N_36379);
and U43369 (N_43369,N_30165,N_39984);
or U43370 (N_43370,N_38374,N_37800);
and U43371 (N_43371,N_32992,N_37873);
xnor U43372 (N_43372,N_36843,N_36457);
xor U43373 (N_43373,N_34354,N_33320);
or U43374 (N_43374,N_34742,N_39688);
and U43375 (N_43375,N_33040,N_31661);
and U43376 (N_43376,N_34401,N_35791);
nor U43377 (N_43377,N_36715,N_31636);
or U43378 (N_43378,N_32503,N_37701);
nor U43379 (N_43379,N_35418,N_32395);
and U43380 (N_43380,N_36432,N_36217);
or U43381 (N_43381,N_39680,N_32408);
nand U43382 (N_43382,N_39821,N_32260);
nor U43383 (N_43383,N_31719,N_32022);
nand U43384 (N_43384,N_34576,N_38235);
and U43385 (N_43385,N_34957,N_32475);
xnor U43386 (N_43386,N_37726,N_37897);
or U43387 (N_43387,N_32973,N_31462);
or U43388 (N_43388,N_31448,N_35427);
nand U43389 (N_43389,N_36428,N_30940);
or U43390 (N_43390,N_34624,N_32392);
and U43391 (N_43391,N_32946,N_30321);
or U43392 (N_43392,N_31902,N_39454);
or U43393 (N_43393,N_37532,N_34244);
and U43394 (N_43394,N_37887,N_36775);
and U43395 (N_43395,N_37162,N_35386);
and U43396 (N_43396,N_37664,N_35565);
nand U43397 (N_43397,N_38537,N_35992);
nand U43398 (N_43398,N_33235,N_38988);
and U43399 (N_43399,N_34819,N_38706);
and U43400 (N_43400,N_35914,N_31489);
nor U43401 (N_43401,N_31060,N_34065);
nor U43402 (N_43402,N_35719,N_33115);
nand U43403 (N_43403,N_31308,N_30141);
and U43404 (N_43404,N_32214,N_35971);
nand U43405 (N_43405,N_39275,N_32996);
nor U43406 (N_43406,N_34930,N_30767);
nor U43407 (N_43407,N_36321,N_38293);
nand U43408 (N_43408,N_39684,N_30020);
nor U43409 (N_43409,N_34240,N_33191);
xnor U43410 (N_43410,N_32533,N_35237);
or U43411 (N_43411,N_34843,N_32003);
nand U43412 (N_43412,N_36000,N_36468);
nand U43413 (N_43413,N_39698,N_30565);
or U43414 (N_43414,N_36425,N_32484);
xor U43415 (N_43415,N_30490,N_37187);
nand U43416 (N_43416,N_34853,N_37180);
and U43417 (N_43417,N_37816,N_31627);
or U43418 (N_43418,N_34483,N_33951);
xnor U43419 (N_43419,N_33722,N_38904);
nor U43420 (N_43420,N_31983,N_33815);
nor U43421 (N_43421,N_32434,N_31698);
nor U43422 (N_43422,N_31181,N_37583);
nor U43423 (N_43423,N_34058,N_39796);
and U43424 (N_43424,N_38348,N_39731);
and U43425 (N_43425,N_33950,N_32986);
nor U43426 (N_43426,N_33192,N_34129);
nor U43427 (N_43427,N_37835,N_31753);
nor U43428 (N_43428,N_37812,N_33321);
nand U43429 (N_43429,N_36534,N_31399);
xnor U43430 (N_43430,N_30320,N_34019);
or U43431 (N_43431,N_35513,N_32144);
nor U43432 (N_43432,N_32753,N_32507);
and U43433 (N_43433,N_33355,N_31404);
or U43434 (N_43434,N_38390,N_38418);
nor U43435 (N_43435,N_33315,N_37903);
and U43436 (N_43436,N_39032,N_33129);
nor U43437 (N_43437,N_36214,N_32139);
nand U43438 (N_43438,N_33833,N_33972);
nor U43439 (N_43439,N_36905,N_37124);
and U43440 (N_43440,N_35117,N_37616);
xor U43441 (N_43441,N_33340,N_34602);
nor U43442 (N_43442,N_34896,N_39015);
or U43443 (N_43443,N_39551,N_30538);
or U43444 (N_43444,N_35756,N_36540);
and U43445 (N_43445,N_35129,N_37071);
and U43446 (N_43446,N_31918,N_38820);
xor U43447 (N_43447,N_36416,N_39779);
xnor U43448 (N_43448,N_34316,N_31001);
or U43449 (N_43449,N_39769,N_36225);
or U43450 (N_43450,N_37445,N_34425);
nand U43451 (N_43451,N_34594,N_37429);
and U43452 (N_43452,N_33587,N_37909);
xor U43453 (N_43453,N_34698,N_33889);
and U43454 (N_43454,N_32084,N_35257);
and U43455 (N_43455,N_36579,N_39574);
nand U43456 (N_43456,N_30677,N_37435);
and U43457 (N_43457,N_38079,N_34236);
nor U43458 (N_43458,N_35534,N_38228);
and U43459 (N_43459,N_35681,N_36126);
or U43460 (N_43460,N_39795,N_36755);
nor U43461 (N_43461,N_37633,N_32716);
nand U43462 (N_43462,N_33099,N_30005);
or U43463 (N_43463,N_33514,N_34687);
nand U43464 (N_43464,N_33915,N_34388);
nand U43465 (N_43465,N_38876,N_37963);
and U43466 (N_43466,N_33803,N_39422);
nand U43467 (N_43467,N_32903,N_39154);
xor U43468 (N_43468,N_37407,N_30127);
and U43469 (N_43469,N_30589,N_39616);
nor U43470 (N_43470,N_31991,N_34725);
or U43471 (N_43471,N_32809,N_37696);
nand U43472 (N_43472,N_32680,N_30730);
nand U43473 (N_43473,N_32299,N_33632);
nor U43474 (N_43474,N_34460,N_39226);
nand U43475 (N_43475,N_35736,N_30910);
and U43476 (N_43476,N_36376,N_32143);
nor U43477 (N_43477,N_32012,N_37156);
or U43478 (N_43478,N_34818,N_30522);
nor U43479 (N_43479,N_39097,N_35644);
nand U43480 (N_43480,N_30788,N_35999);
nor U43481 (N_43481,N_36234,N_35898);
and U43482 (N_43482,N_39870,N_32701);
or U43483 (N_43483,N_31580,N_32579);
nand U43484 (N_43484,N_33054,N_32163);
and U43485 (N_43485,N_37735,N_34676);
and U43486 (N_43486,N_32933,N_30839);
or U43487 (N_43487,N_35439,N_34775);
nand U43488 (N_43488,N_32563,N_30528);
nand U43489 (N_43489,N_35047,N_34382);
and U43490 (N_43490,N_31460,N_32742);
or U43491 (N_43491,N_37938,N_35005);
and U43492 (N_43492,N_38777,N_34652);
nand U43493 (N_43493,N_35559,N_34573);
nor U43494 (N_43494,N_38584,N_32799);
nor U43495 (N_43495,N_33969,N_35236);
nor U43496 (N_43496,N_39912,N_37449);
or U43497 (N_43497,N_38482,N_30863);
or U43498 (N_43498,N_30479,N_37507);
nor U43499 (N_43499,N_31049,N_39137);
nor U43500 (N_43500,N_36707,N_31407);
or U43501 (N_43501,N_38693,N_33712);
nand U43502 (N_43502,N_38758,N_37244);
nand U43503 (N_43503,N_34323,N_33844);
nand U43504 (N_43504,N_38748,N_38069);
and U43505 (N_43505,N_37254,N_33435);
nand U43506 (N_43506,N_39619,N_34253);
or U43507 (N_43507,N_33962,N_35226);
nor U43508 (N_43508,N_37357,N_30569);
and U43509 (N_43509,N_35696,N_33817);
and U43510 (N_43510,N_35507,N_33615);
xnor U43511 (N_43511,N_33014,N_30764);
xnor U43512 (N_43512,N_37272,N_37024);
and U43513 (N_43513,N_39052,N_36384);
nor U43514 (N_43514,N_33034,N_30460);
nand U43515 (N_43515,N_38333,N_32085);
xor U43516 (N_43516,N_39709,N_39823);
or U43517 (N_43517,N_37837,N_33520);
nand U43518 (N_43518,N_33401,N_31892);
and U43519 (N_43519,N_31486,N_37557);
or U43520 (N_43520,N_30223,N_33874);
nand U43521 (N_43521,N_33212,N_38837);
or U43522 (N_43522,N_36035,N_35356);
and U43523 (N_43523,N_34186,N_37444);
and U43524 (N_43524,N_33169,N_37650);
or U43525 (N_43525,N_31706,N_31385);
and U43526 (N_43526,N_32242,N_32477);
and U43527 (N_43527,N_32136,N_32281);
and U43528 (N_43528,N_33853,N_37284);
or U43529 (N_43529,N_34309,N_32656);
nor U43530 (N_43530,N_34298,N_38823);
and U43531 (N_43531,N_39584,N_34424);
nor U43532 (N_43532,N_32755,N_35918);
nor U43533 (N_43533,N_34004,N_39654);
nand U43534 (N_43534,N_38447,N_35018);
xor U43535 (N_43535,N_38803,N_35927);
nand U43536 (N_43536,N_32206,N_31063);
nand U43537 (N_43537,N_33352,N_33578);
nand U43538 (N_43538,N_31765,N_33280);
nor U43539 (N_43539,N_35488,N_37529);
or U43540 (N_43540,N_36340,N_34710);
or U43541 (N_43541,N_34400,N_30032);
nand U43542 (N_43542,N_36590,N_34656);
or U43543 (N_43543,N_32156,N_30937);
and U43544 (N_43544,N_39523,N_39954);
xor U43545 (N_43545,N_31602,N_39864);
or U43546 (N_43546,N_31380,N_39858);
and U43547 (N_43547,N_39955,N_33952);
and U43548 (N_43548,N_31545,N_30696);
nor U43549 (N_43549,N_34717,N_31397);
or U43550 (N_43550,N_30181,N_36819);
or U43551 (N_43551,N_31477,N_31152);
and U43552 (N_43552,N_36226,N_32099);
xor U43553 (N_43553,N_39036,N_34831);
nor U43554 (N_43554,N_38432,N_39786);
nor U43555 (N_43555,N_38479,N_36195);
nor U43556 (N_43556,N_34052,N_38796);
or U43557 (N_43557,N_36350,N_31209);
and U43558 (N_43558,N_32064,N_30658);
nand U43559 (N_43559,N_30763,N_35008);
nand U43560 (N_43560,N_34404,N_37031);
and U43561 (N_43561,N_33141,N_35906);
nor U43562 (N_43562,N_36947,N_39285);
and U43563 (N_43563,N_36524,N_39675);
nand U43564 (N_43564,N_36013,N_35443);
nand U43565 (N_43565,N_31896,N_37310);
or U43566 (N_43566,N_32959,N_37397);
nand U43567 (N_43567,N_32039,N_39604);
xnor U43568 (N_43568,N_32014,N_31422);
and U43569 (N_43569,N_32407,N_38420);
and U43570 (N_43570,N_36363,N_37910);
xnor U43571 (N_43571,N_38052,N_32266);
nor U43572 (N_43572,N_37604,N_39146);
or U43573 (N_43573,N_32368,N_36279);
nand U43574 (N_43574,N_34976,N_38014);
xnor U43575 (N_43575,N_33886,N_38963);
or U43576 (N_43576,N_36767,N_36186);
and U43577 (N_43577,N_34931,N_32466);
nand U43578 (N_43578,N_32146,N_33242);
xnor U43579 (N_43579,N_32581,N_31403);
nand U43580 (N_43580,N_33462,N_38113);
and U43581 (N_43581,N_38868,N_36030);
nor U43582 (N_43582,N_39089,N_30935);
xor U43583 (N_43583,N_31168,N_30532);
and U43584 (N_43584,N_31271,N_35046);
nor U43585 (N_43585,N_35485,N_32975);
and U43586 (N_43586,N_30499,N_32640);
nand U43587 (N_43587,N_36237,N_36085);
and U43588 (N_43588,N_38759,N_36022);
nand U43589 (N_43589,N_39477,N_33223);
xnor U43590 (N_43590,N_34784,N_30812);
nand U43591 (N_43591,N_35750,N_33766);
and U43592 (N_43592,N_30646,N_32029);
or U43593 (N_43593,N_30695,N_36404);
nand U43594 (N_43594,N_30735,N_36075);
nor U43595 (N_43595,N_34136,N_34131);
nand U43596 (N_43596,N_31478,N_30766);
nor U43597 (N_43597,N_30367,N_36181);
or U43598 (N_43598,N_36010,N_36933);
and U43599 (N_43599,N_31804,N_34432);
and U43600 (N_43600,N_31663,N_38811);
or U43601 (N_43601,N_31376,N_35768);
nor U43602 (N_43602,N_32492,N_33550);
nand U43603 (N_43603,N_33661,N_39896);
and U43604 (N_43604,N_38354,N_34102);
nand U43605 (N_43605,N_38892,N_31945);
or U43606 (N_43606,N_37056,N_30343);
and U43607 (N_43607,N_32418,N_36253);
nor U43608 (N_43608,N_33569,N_31252);
and U43609 (N_43609,N_32909,N_30996);
and U43610 (N_43610,N_33163,N_35460);
and U43611 (N_43611,N_36664,N_39274);
and U43612 (N_43612,N_31287,N_33672);
and U43613 (N_43613,N_39073,N_32885);
xor U43614 (N_43614,N_39582,N_35026);
nand U43615 (N_43615,N_37238,N_39694);
nor U43616 (N_43616,N_31906,N_38494);
nand U43617 (N_43617,N_32468,N_35628);
nand U43618 (N_43618,N_32354,N_35184);
nor U43619 (N_43619,N_31456,N_34613);
nor U43620 (N_43620,N_32984,N_35723);
and U43621 (N_43621,N_32538,N_31269);
and U43622 (N_43622,N_31423,N_31883);
and U43623 (N_43623,N_37723,N_34495);
or U43624 (N_43624,N_32504,N_35240);
nand U43625 (N_43625,N_34484,N_31145);
and U43626 (N_43626,N_33032,N_31997);
or U43627 (N_43627,N_36575,N_35897);
nand U43628 (N_43628,N_33362,N_36981);
nor U43629 (N_43629,N_32311,N_35924);
nor U43630 (N_43630,N_36031,N_33897);
nand U43631 (N_43631,N_37367,N_36421);
nor U43632 (N_43632,N_33912,N_30549);
or U43633 (N_43633,N_30339,N_31071);
nand U43634 (N_43634,N_30795,N_34067);
or U43635 (N_43635,N_30667,N_31102);
or U43636 (N_43636,N_33664,N_32764);
or U43637 (N_43637,N_33834,N_31251);
nor U43638 (N_43638,N_30865,N_39051);
xor U43639 (N_43639,N_39234,N_33314);
nor U43640 (N_43640,N_34766,N_39737);
nand U43641 (N_43641,N_31960,N_37907);
and U43642 (N_43642,N_36280,N_32896);
and U43643 (N_43643,N_30292,N_37200);
nand U43644 (N_43644,N_34104,N_30406);
nand U43645 (N_43645,N_33966,N_38194);
and U43646 (N_43646,N_30931,N_33744);
nor U43647 (N_43647,N_36603,N_38891);
and U43648 (N_43648,N_31081,N_33839);
or U43649 (N_43649,N_37209,N_38192);
and U43650 (N_43650,N_30580,N_38471);
and U43651 (N_43651,N_35594,N_32963);
or U43652 (N_43652,N_32124,N_33269);
nor U43653 (N_43653,N_32650,N_38248);
or U43654 (N_43654,N_39690,N_33437);
xor U43655 (N_43655,N_39936,N_38024);
nand U43656 (N_43656,N_37285,N_33575);
xor U43657 (N_43657,N_33464,N_32238);
nor U43658 (N_43658,N_38692,N_31799);
and U43659 (N_43659,N_31598,N_31346);
and U43660 (N_43660,N_34185,N_35261);
nor U43661 (N_43661,N_32367,N_32718);
or U43662 (N_43662,N_33412,N_37094);
nand U43663 (N_43663,N_31638,N_30210);
nor U43664 (N_43664,N_38346,N_31436);
nor U43665 (N_43665,N_37519,N_38688);
and U43666 (N_43666,N_30301,N_33540);
nor U43667 (N_43667,N_32351,N_30890);
nand U43668 (N_43668,N_38355,N_32028);
and U43669 (N_43669,N_35139,N_37737);
or U43670 (N_43670,N_39879,N_36541);
nor U43671 (N_43671,N_34056,N_35176);
nand U43672 (N_43672,N_30851,N_30036);
or U43673 (N_43673,N_35247,N_30398);
or U43674 (N_43674,N_37312,N_38038);
nand U43675 (N_43675,N_34263,N_36023);
or U43676 (N_43676,N_34510,N_33224);
nor U43677 (N_43677,N_31794,N_34115);
and U43678 (N_43678,N_31447,N_36730);
or U43679 (N_43679,N_39059,N_34048);
and U43680 (N_43680,N_37293,N_33671);
nor U43681 (N_43681,N_30576,N_36021);
or U43682 (N_43682,N_38973,N_30366);
and U43683 (N_43683,N_38875,N_30917);
or U43684 (N_43684,N_37554,N_31672);
nand U43685 (N_43685,N_35273,N_36497);
xnor U43686 (N_43686,N_30573,N_31931);
and U43687 (N_43687,N_33239,N_39947);
and U43688 (N_43688,N_38943,N_34803);
and U43689 (N_43689,N_33126,N_33970);
and U43690 (N_43690,N_37888,N_38611);
nor U43691 (N_43691,N_37295,N_37749);
and U43692 (N_43692,N_33132,N_33512);
nor U43693 (N_43693,N_38694,N_34646);
or U43694 (N_43694,N_35320,N_31684);
or U43695 (N_43695,N_36263,N_35416);
nor U43696 (N_43696,N_33904,N_37074);
or U43697 (N_43697,N_33739,N_31543);
nor U43698 (N_43698,N_39498,N_35662);
xnor U43699 (N_43699,N_39843,N_31411);
nor U43700 (N_43700,N_32654,N_30790);
xnor U43701 (N_43701,N_34889,N_36442);
nor U43702 (N_43702,N_34327,N_37624);
xnor U43703 (N_43703,N_37080,N_37230);
nor U43704 (N_43704,N_36720,N_34909);
nand U43705 (N_43705,N_32971,N_31850);
or U43706 (N_43706,N_34297,N_32917);
or U43707 (N_43707,N_38394,N_31364);
nor U43708 (N_43708,N_36571,N_30602);
xnor U43709 (N_43709,N_32015,N_34193);
or U43710 (N_43710,N_31692,N_33630);
or U43711 (N_43711,N_36891,N_31193);
nand U43712 (N_43712,N_31587,N_31929);
nand U43713 (N_43713,N_38154,N_32725);
nand U43714 (N_43714,N_34875,N_32355);
or U43715 (N_43715,N_35498,N_32974);
or U43716 (N_43716,N_36292,N_35461);
xnor U43717 (N_43717,N_31406,N_36223);
and U43718 (N_43718,N_32262,N_37764);
or U43719 (N_43719,N_31507,N_39300);
nand U43720 (N_43720,N_34603,N_34910);
and U43721 (N_43721,N_32682,N_36098);
nor U43722 (N_43722,N_35535,N_30469);
or U43723 (N_43723,N_33649,N_31848);
and U43724 (N_43724,N_39169,N_35001);
or U43725 (N_43725,N_35572,N_34962);
xor U43726 (N_43726,N_37283,N_36142);
nand U43727 (N_43727,N_30627,N_34485);
nand U43728 (N_43728,N_32033,N_31097);
nor U43729 (N_43729,N_37729,N_37478);
xnor U43730 (N_43730,N_33061,N_35270);
or U43731 (N_43731,N_38776,N_34325);
nand U43732 (N_43732,N_35187,N_35315);
nor U43733 (N_43733,N_30052,N_32328);
nor U43734 (N_43734,N_32874,N_39450);
nand U43735 (N_43735,N_38847,N_36111);
nand U43736 (N_43736,N_39791,N_31821);
nand U43737 (N_43737,N_37852,N_31171);
nor U43738 (N_43738,N_36660,N_33848);
xnor U43739 (N_43739,N_37188,N_37718);
and U43740 (N_43740,N_34003,N_34825);
and U43741 (N_43741,N_34119,N_35626);
nand U43742 (N_43742,N_32159,N_32762);
or U43743 (N_43743,N_37567,N_34574);
or U43744 (N_43744,N_38853,N_33842);
and U43745 (N_43745,N_32894,N_39869);
and U43746 (N_43746,N_32578,N_32826);
and U43747 (N_43747,N_37232,N_34063);
and U43748 (N_43748,N_30122,N_31211);
or U43749 (N_43749,N_32977,N_38818);
or U43750 (N_43750,N_34953,N_38539);
nor U43751 (N_43751,N_36873,N_34322);
nand U43752 (N_43752,N_32962,N_38102);
xor U43753 (N_43753,N_33466,N_30180);
nor U43754 (N_43754,N_32617,N_31533);
nor U43755 (N_43755,N_35352,N_31183);
and U43756 (N_43756,N_34132,N_35475);
nand U43757 (N_43757,N_36652,N_30498);
and U43758 (N_43758,N_33433,N_33432);
or U43759 (N_43759,N_36258,N_34623);
nand U43760 (N_43760,N_30153,N_33871);
nor U43761 (N_43761,N_35929,N_32914);
nor U43762 (N_43762,N_37353,N_33532);
nor U43763 (N_43763,N_38280,N_39393);
or U43764 (N_43764,N_31524,N_31131);
nand U43765 (N_43765,N_39041,N_32726);
nor U43766 (N_43766,N_36716,N_36655);
and U43767 (N_43767,N_39439,N_33629);
and U43768 (N_43768,N_30289,N_32793);
xor U43769 (N_43769,N_38619,N_32819);
nor U43770 (N_43770,N_36386,N_30101);
and U43771 (N_43771,N_33873,N_32174);
and U43772 (N_43772,N_39025,N_37944);
nand U43773 (N_43773,N_36426,N_31561);
and U43774 (N_43774,N_33455,N_34747);
or U43775 (N_43775,N_39985,N_39457);
and U43776 (N_43776,N_34491,N_36334);
or U43777 (N_43777,N_32034,N_34114);
or U43778 (N_43778,N_38604,N_30068);
nor U43779 (N_43779,N_37348,N_39909);
nand U43780 (N_43780,N_31773,N_30049);
xnor U43781 (N_43781,N_31911,N_35125);
nand U43782 (N_43782,N_30254,N_35376);
nor U43783 (N_43783,N_32378,N_33662);
nor U43784 (N_43784,N_30010,N_31429);
nand U43785 (N_43785,N_38317,N_38245);
nor U43786 (N_43786,N_38846,N_38594);
or U43787 (N_43787,N_39444,N_33721);
nand U43788 (N_43788,N_35478,N_36218);
nand U43789 (N_43789,N_32611,N_30959);
or U43790 (N_43790,N_36197,N_31780);
or U43791 (N_43791,N_37880,N_33271);
nand U43792 (N_43792,N_34014,N_31606);
nand U43793 (N_43793,N_38415,N_33177);
and U43794 (N_43794,N_39832,N_31954);
nand U43795 (N_43795,N_36622,N_33171);
nand U43796 (N_43796,N_31450,N_35462);
nand U43797 (N_43797,N_32004,N_30613);
nand U43798 (N_43798,N_32802,N_39719);
and U43799 (N_43799,N_36989,N_38325);
or U43800 (N_43800,N_39365,N_36154);
and U43801 (N_43801,N_30978,N_34626);
nand U43802 (N_43802,N_33251,N_34767);
and U43803 (N_43803,N_39142,N_36786);
nand U43804 (N_43804,N_34311,N_32670);
or U43805 (N_43805,N_36685,N_36640);
and U43806 (N_43806,N_35451,N_37075);
nand U43807 (N_43807,N_38965,N_37292);
or U43808 (N_43808,N_39380,N_37510);
and U43809 (N_43809,N_33488,N_32499);
and U43810 (N_43810,N_30137,N_31632);
and U43811 (N_43811,N_39337,N_34252);
nor U43812 (N_43812,N_32059,N_37697);
xnor U43813 (N_43813,N_32858,N_37027);
and U43814 (N_43814,N_37249,N_32443);
nor U43815 (N_43815,N_30715,N_39094);
nor U43816 (N_43816,N_30765,N_32618);
nand U43817 (N_43817,N_38666,N_38857);
or U43818 (N_43818,N_34508,N_33857);
and U43819 (N_43819,N_37226,N_31320);
nor U43820 (N_43820,N_30555,N_34512);
nor U43821 (N_43821,N_30324,N_37862);
or U43822 (N_43822,N_30176,N_32382);
or U43823 (N_43823,N_37772,N_31755);
xnor U43824 (N_43824,N_38532,N_31942);
or U43825 (N_43825,N_36199,N_39658);
xor U43826 (N_43826,N_38962,N_39687);
and U43827 (N_43827,N_30956,N_37601);
nor U43828 (N_43828,N_31645,N_30754);
or U43829 (N_43829,N_38465,N_38966);
xor U43830 (N_43830,N_32204,N_32486);
and U43831 (N_43831,N_37448,N_34324);
or U43832 (N_43832,N_37965,N_31768);
nor U43833 (N_43833,N_35336,N_37565);
and U43834 (N_43834,N_32230,N_32343);
or U43835 (N_43835,N_36510,N_34653);
nor U43836 (N_43836,N_30647,N_37494);
and U43837 (N_43837,N_35515,N_38186);
nor U43838 (N_43838,N_37959,N_32471);
and U43839 (N_43839,N_37636,N_33093);
and U43840 (N_43840,N_39710,N_36523);
nor U43841 (N_43841,N_32379,N_35812);
nand U43842 (N_43842,N_37361,N_32695);
and U43843 (N_43843,N_32926,N_35786);
and U43844 (N_43844,N_39001,N_34367);
nand U43845 (N_43845,N_36756,N_34256);
nor U43846 (N_43846,N_39433,N_35529);
xor U43847 (N_43847,N_31479,N_34694);
nor U43848 (N_43848,N_36353,N_34433);
nor U43849 (N_43849,N_32067,N_36275);
and U43850 (N_43850,N_33149,N_35602);
or U43851 (N_43851,N_39536,N_31882);
or U43852 (N_43852,N_35899,N_36549);
or U43853 (N_43853,N_39875,N_34593);
or U43854 (N_43854,N_35504,N_36222);
nand U43855 (N_43855,N_32687,N_32845);
xor U43856 (N_43856,N_38105,N_31295);
or U43857 (N_43857,N_35843,N_31728);
nor U43858 (N_43858,N_30007,N_39926);
and U43859 (N_43859,N_31677,N_30679);
or U43860 (N_43860,N_33798,N_36060);
nor U43861 (N_43861,N_38450,N_38789);
nor U43862 (N_43862,N_32211,N_37892);
nand U43863 (N_43863,N_36057,N_30457);
nor U43864 (N_43864,N_38720,N_32520);
or U43865 (N_43865,N_33264,N_30567);
or U43866 (N_43866,N_30177,N_38531);
or U43867 (N_43867,N_39326,N_31713);
xnor U43868 (N_43868,N_30334,N_31089);
nor U43869 (N_43869,N_34807,N_38253);
or U43870 (N_43870,N_30288,N_35053);
and U43871 (N_43871,N_35637,N_35633);
or U43872 (N_43872,N_31976,N_35544);
nor U43873 (N_43873,N_35598,N_36747);
and U43874 (N_43874,N_38627,N_30798);
nor U43875 (N_43875,N_34234,N_36624);
nor U43876 (N_43876,N_30400,N_32960);
nor U43877 (N_43877,N_36695,N_33902);
or U43878 (N_43878,N_32841,N_30512);
nand U43879 (N_43879,N_32748,N_37057);
or U43880 (N_43880,N_35972,N_38134);
or U43881 (N_43881,N_31907,N_30241);
nor U43882 (N_43882,N_31419,N_33818);
or U43883 (N_43883,N_31057,N_32284);
and U43884 (N_43884,N_32248,N_38383);
nand U43885 (N_43885,N_35375,N_31109);
and U43886 (N_43886,N_30541,N_36582);
or U43887 (N_43887,N_36243,N_38163);
xnor U43888 (N_43888,N_39743,N_39581);
and U43889 (N_43889,N_33825,N_30853);
and U43890 (N_43890,N_35186,N_38161);
nand U43891 (N_43891,N_34409,N_36667);
and U43892 (N_43892,N_37693,N_37918);
and U43893 (N_43893,N_33808,N_34730);
and U43894 (N_43894,N_30480,N_32763);
nor U43895 (N_43895,N_39712,N_39831);
nor U43896 (N_43896,N_32231,N_39264);
nor U43897 (N_43897,N_34871,N_30883);
nor U43898 (N_43898,N_33976,N_35497);
nand U43899 (N_43899,N_32104,N_34834);
and U43900 (N_43900,N_35948,N_30621);
nor U43901 (N_43901,N_34482,N_39692);
nand U43902 (N_43902,N_36573,N_33692);
nand U43903 (N_43903,N_36074,N_30463);
nand U43904 (N_43904,N_34583,N_39835);
nand U43905 (N_43905,N_37487,N_35002);
or U43906 (N_43906,N_30629,N_31515);
and U43907 (N_43907,N_34534,N_32442);
or U43908 (N_43908,N_35962,N_32414);
and U43909 (N_43909,N_32864,N_31915);
and U43910 (N_43910,N_39976,N_37415);
nand U43911 (N_43911,N_33968,N_38431);
nor U43912 (N_43912,N_32068,N_39783);
xor U43913 (N_43913,N_33960,N_38817);
and U43914 (N_43914,N_37646,N_35277);
xor U43915 (N_43915,N_32807,N_39194);
or U43916 (N_43916,N_30285,N_34913);
and U43917 (N_43917,N_35082,N_34972);
nand U43918 (N_43918,N_34552,N_35577);
nor U43919 (N_43919,N_30405,N_39932);
or U43920 (N_43920,N_30941,N_33843);
or U43921 (N_43921,N_31952,N_35193);
xor U43922 (N_43922,N_37684,N_39781);
nand U43923 (N_43923,N_37533,N_34260);
or U43924 (N_43924,N_39364,N_32710);
or U43925 (N_43925,N_31338,N_30896);
and U43926 (N_43926,N_35173,N_32474);
nor U43927 (N_43927,N_35246,N_39560);
nand U43928 (N_43928,N_31732,N_38618);
nor U43929 (N_43929,N_33179,N_38615);
nand U43930 (N_43930,N_31927,N_36052);
nor U43931 (N_43931,N_34908,N_34051);
nor U43932 (N_43932,N_36615,N_33667);
and U43933 (N_43933,N_35960,N_39720);
xor U43934 (N_43934,N_35406,N_37112);
or U43935 (N_43935,N_31383,N_32588);
xor U43936 (N_43936,N_37719,N_34155);
xnor U43937 (N_43937,N_38446,N_34418);
nand U43938 (N_43938,N_34544,N_33879);
nand U43939 (N_43939,N_31739,N_34304);
or U43940 (N_43940,N_36172,N_35938);
nor U43941 (N_43941,N_30985,N_35525);
or U43942 (N_43942,N_33813,N_36489);
and U43943 (N_43943,N_33410,N_37043);
and U43944 (N_43944,N_39280,N_33982);
nand U43945 (N_43945,N_38671,N_33143);
nand U43946 (N_43946,N_35339,N_37476);
nor U43947 (N_43947,N_34239,N_37665);
and U43948 (N_43948,N_37046,N_36912);
nor U43949 (N_43949,N_31825,N_35217);
nor U43950 (N_43950,N_36149,N_38587);
nand U43951 (N_43951,N_38782,N_35762);
nand U43952 (N_43952,N_32653,N_35160);
or U43953 (N_43953,N_37785,N_35457);
nand U43954 (N_43954,N_34420,N_38273);
and U43955 (N_43955,N_35630,N_33186);
nand U43956 (N_43956,N_30089,N_31601);
nand U43957 (N_43957,N_33274,N_37441);
nand U43958 (N_43958,N_30416,N_38800);
nor U43959 (N_43959,N_38502,N_35769);
nor U43960 (N_43960,N_31576,N_30003);
or U43961 (N_43961,N_36153,N_31842);
or U43962 (N_43962,N_33868,N_34943);
xor U43963 (N_43963,N_39209,N_32289);
or U43964 (N_43964,N_36617,N_33450);
nand U43965 (N_43965,N_35580,N_33918);
and U43966 (N_43966,N_32649,N_36836);
and U43967 (N_43967,N_32421,N_35287);
and U43968 (N_43968,N_38557,N_32711);
xnor U43969 (N_43969,N_32560,N_31359);
nor U43970 (N_43970,N_36009,N_33467);
xor U43971 (N_43971,N_35994,N_32785);
nor U43972 (N_43972,N_33866,N_32890);
or U43973 (N_43973,N_34780,N_36242);
nor U43974 (N_43974,N_37542,N_39277);
nand U43975 (N_43975,N_34361,N_38159);
and U43976 (N_43976,N_34293,N_38260);
nor U43977 (N_43977,N_37589,N_33822);
nand U43978 (N_43978,N_34934,N_38080);
and U43979 (N_43979,N_30909,N_37931);
and U43980 (N_43980,N_30975,N_35822);
and U43981 (N_43981,N_33634,N_39558);
or U43982 (N_43982,N_30327,N_32562);
nand U43983 (N_43983,N_34211,N_30847);
and U43984 (N_43984,N_32274,N_39063);
and U43985 (N_43985,N_36701,N_31557);
and U43986 (N_43986,N_30964,N_31815);
nand U43987 (N_43987,N_31394,N_38066);
nor U43988 (N_43988,N_31908,N_32055);
nand U43989 (N_43989,N_34705,N_31776);
xnor U43990 (N_43990,N_39563,N_32969);
xnor U43991 (N_43991,N_32938,N_33133);
and U43992 (N_43992,N_37155,N_36736);
nor U43993 (N_43993,N_30257,N_31415);
nor U43994 (N_43994,N_38082,N_35560);
nor U43995 (N_43995,N_31819,N_34421);
nand U43996 (N_43996,N_37889,N_35264);
xnor U43997 (N_43997,N_30774,N_32141);
nor U43998 (N_43998,N_34183,N_30145);
and U43999 (N_43999,N_39964,N_30710);
and U44000 (N_44000,N_38839,N_32370);
or U44001 (N_44001,N_33568,N_35309);
nor U44002 (N_44002,N_38043,N_33386);
nand U44003 (N_44003,N_34177,N_36438);
nor U44004 (N_44004,N_32148,N_31560);
nand U44005 (N_44005,N_34918,N_36694);
nor U44006 (N_44006,N_39894,N_36054);
and U44007 (N_44007,N_36110,N_39819);
nand U44008 (N_44008,N_31377,N_35227);
or U44009 (N_44009,N_36261,N_33920);
and U44010 (N_44010,N_31493,N_36396);
or U44011 (N_44011,N_30135,N_39785);
or U44012 (N_44012,N_34406,N_34144);
nor U44013 (N_44013,N_32657,N_36633);
xor U44014 (N_44014,N_36941,N_33543);
or U44015 (N_44015,N_33405,N_38999);
nand U44016 (N_44016,N_30566,N_37253);
xnor U44017 (N_44017,N_34417,N_35206);
and U44018 (N_44018,N_31793,N_34195);
or U44019 (N_44019,N_36359,N_30727);
and U44020 (N_44020,N_37358,N_38916);
nand U44021 (N_44021,N_39780,N_34489);
and U44022 (N_44022,N_36144,N_39385);
and U44023 (N_44023,N_30887,N_39901);
and U44024 (N_44024,N_34979,N_39478);
or U44025 (N_44025,N_32921,N_36776);
nor U44026 (N_44026,N_31121,N_30742);
or U44027 (N_44027,N_36283,N_33167);
nand U44028 (N_44028,N_35494,N_30643);
or U44029 (N_44029,N_30579,N_32908);
nand U44030 (N_44030,N_31294,N_31930);
nor U44031 (N_44031,N_39841,N_38445);
or U44032 (N_44032,N_39067,N_39177);
and U44033 (N_44033,N_30310,N_38510);
nand U44034 (N_44034,N_33200,N_32775);
and U44035 (N_44035,N_33262,N_32013);
nand U44036 (N_44036,N_39031,N_31862);
or U44037 (N_44037,N_34413,N_36598);
and U44038 (N_44038,N_32125,N_33468);
nand U44039 (N_44039,N_38910,N_35825);
or U44040 (N_44040,N_36665,N_34863);
nand U44041 (N_44041,N_35848,N_35520);
nor U44042 (N_44042,N_31310,N_34586);
nor U44043 (N_44043,N_34428,N_33123);
or U44044 (N_44044,N_34223,N_35221);
nor U44045 (N_44045,N_35970,N_37501);
nand U44046 (N_44046,N_38527,N_34865);
or U44047 (N_44047,N_31858,N_34682);
nor U44048 (N_44048,N_39519,N_36390);
and U44049 (N_44049,N_35265,N_39021);
and U44050 (N_44050,N_36313,N_31992);
nor U44051 (N_44051,N_33080,N_30047);
nor U44052 (N_44052,N_38906,N_32943);
nand U44053 (N_44053,N_34605,N_38335);
and U44054 (N_44054,N_39648,N_38073);
or U44055 (N_44055,N_32737,N_32948);
or U44056 (N_44056,N_34101,N_35809);
nand U44057 (N_44057,N_36986,N_32349);
nand U44058 (N_44058,N_36712,N_35371);
or U44059 (N_44059,N_39350,N_34521);
nor U44060 (N_44060,N_39068,N_36002);
nand U44061 (N_44061,N_39279,N_33199);
nor U44062 (N_44062,N_37366,N_31480);
nor U44063 (N_44063,N_33391,N_37065);
nand U44064 (N_44064,N_30194,N_36148);
and U44065 (N_44065,N_38493,N_38830);
nor U44066 (N_44066,N_39598,N_38795);
nand U44067 (N_44067,N_32632,N_34986);
xnor U44068 (N_44068,N_38507,N_33956);
or U44069 (N_44069,N_34120,N_30340);
nor U44070 (N_44070,N_36969,N_39311);
nand U44071 (N_44071,N_33396,N_30750);
nor U44072 (N_44072,N_37807,N_33748);
or U44073 (N_44073,N_36726,N_34008);
and U44074 (N_44074,N_33374,N_37119);
and U44075 (N_44075,N_32128,N_31305);
and U44076 (N_44076,N_38648,N_31752);
nor U44077 (N_44077,N_32173,N_39794);
or U44078 (N_44078,N_33146,N_35619);
and U44079 (N_44079,N_39856,N_36693);
or U44080 (N_44080,N_36689,N_33971);
nand U44081 (N_44081,N_39386,N_30382);
and U44082 (N_44082,N_37991,N_30601);
nand U44083 (N_44083,N_39728,N_38308);
nor U44084 (N_44084,N_35724,N_38074);
nand U44085 (N_44085,N_38281,N_32077);
xor U44086 (N_44086,N_34789,N_30118);
and U44087 (N_44087,N_33302,N_30287);
xnor U44088 (N_44088,N_35783,N_35127);
or U44089 (N_44089,N_33801,N_37632);
xnor U44090 (N_44090,N_30582,N_31165);
or U44091 (N_44091,N_36170,N_31999);
or U44092 (N_44092,N_36725,N_30134);
and U44093 (N_44093,N_34855,N_31292);
nand U44094 (N_44094,N_37921,N_30969);
nor U44095 (N_44095,N_31735,N_36208);
and U44096 (N_44096,N_30547,N_30731);
and U44097 (N_44097,N_36631,N_37818);
or U44098 (N_44098,N_31203,N_39801);
and U44099 (N_44099,N_38340,N_36522);
and U44100 (N_44100,N_38589,N_37434);
nand U44101 (N_44101,N_35771,N_38896);
xnor U44102 (N_44102,N_33342,N_38970);
nor U44103 (N_44103,N_37548,N_32771);
or U44104 (N_44104,N_34026,N_39027);
and U44105 (N_44105,N_37015,N_30352);
nor U44106 (N_44106,N_39775,N_31946);
nand U44107 (N_44107,N_34533,N_33461);
xnor U44108 (N_44108,N_38146,N_34162);
nand U44109 (N_44109,N_36806,N_37503);
nand U44110 (N_44110,N_38238,N_35612);
and U44111 (N_44111,N_38444,N_30804);
and U44112 (N_44112,N_35253,N_34587);
and U44113 (N_44113,N_33861,N_31365);
or U44114 (N_44114,N_37488,N_34389);
and U44115 (N_44115,N_35010,N_37998);
and U44116 (N_44116,N_34390,N_39269);
nor U44117 (N_44117,N_35817,N_35342);
or U44118 (N_44118,N_39996,N_35067);
nand U44119 (N_44119,N_35470,N_32521);
and U44120 (N_44120,N_37734,N_36160);
or U44121 (N_44121,N_36853,N_31144);
nand U44122 (N_44122,N_36201,N_33917);
xnor U44123 (N_44123,N_34696,N_36337);
nand U44124 (N_44124,N_36240,N_39713);
or U44125 (N_44125,N_30095,N_30644);
or U44126 (N_44126,N_34761,N_30286);
and U44127 (N_44127,N_32853,N_34200);
and U44128 (N_44128,N_32697,N_34383);
nand U44129 (N_44129,N_39482,N_36671);
nand U44130 (N_44130,N_33585,N_37393);
nor U44131 (N_44131,N_34168,N_36924);
nand U44132 (N_44132,N_35069,N_36045);
nor U44133 (N_44133,N_39825,N_34707);
or U44134 (N_44134,N_35607,N_34919);
or U44135 (N_44135,N_37037,N_35808);
nand U44136 (N_44136,N_33390,N_35348);
xor U44137 (N_44137,N_38221,N_34258);
or U44138 (N_44138,N_33045,N_34209);
nor U44139 (N_44139,N_37107,N_36971);
or U44140 (N_44140,N_30518,N_34288);
xnor U44141 (N_44141,N_32535,N_36461);
xnor U44142 (N_44142,N_35824,N_34254);
nand U44143 (N_44143,N_35933,N_38275);
or U44144 (N_44144,N_39890,N_35964);
nor U44145 (N_44145,N_38295,N_32530);
xnor U44146 (N_44146,N_34331,N_37240);
and U44147 (N_44147,N_36885,N_39848);
nor U44148 (N_44148,N_33284,N_34376);
nand U44149 (N_44149,N_31150,N_31809);
xnor U44150 (N_44150,N_35220,N_39371);
and U44151 (N_44151,N_36437,N_35012);
nand U44152 (N_44152,N_31127,N_34529);
xor U44153 (N_44153,N_32847,N_38732);
xor U44154 (N_44154,N_37870,N_33576);
nor U44155 (N_44155,N_35433,N_33777);
and U44156 (N_44156,N_36411,N_36651);
nor U44157 (N_44157,N_36485,N_38976);
nand U44158 (N_44158,N_33679,N_36854);
nand U44159 (N_44159,N_36255,N_32019);
and U44160 (N_44160,N_39451,N_34041);
nand U44161 (N_44161,N_38953,N_37833);
nand U44162 (N_44162,N_36318,N_38214);
and U44163 (N_44163,N_34446,N_33746);
nand U44164 (N_44164,N_30207,N_30474);
and U44165 (N_44165,N_34314,N_37868);
nand U44166 (N_44166,N_31317,N_35539);
nor U44167 (N_44167,N_33954,N_36264);
or U44168 (N_44168,N_32678,N_36365);
or U44169 (N_44169,N_39133,N_36530);
and U44170 (N_44170,N_34958,N_37148);
and U44171 (N_44171,N_32358,N_38650);
nor U44172 (N_44172,N_39809,N_39136);
nor U44173 (N_44173,N_33876,N_37320);
or U44174 (N_44174,N_36904,N_34672);
and U44175 (N_44175,N_33085,N_33270);
nand U44176 (N_44176,N_32932,N_35459);
or U44177 (N_44177,N_38883,N_35381);
nor U44178 (N_44178,N_35733,N_32110);
and U44179 (N_44179,N_36968,N_31283);
nor U44180 (N_44180,N_36639,N_34103);
nor U44181 (N_44181,N_32811,N_34068);
and U44182 (N_44182,N_37794,N_38948);
or U44183 (N_44183,N_30336,N_35839);
and U44184 (N_44184,N_39129,N_34611);
nor U44185 (N_44185,N_39765,N_37014);
or U44186 (N_44186,N_30455,N_34342);
nand U44187 (N_44187,N_33566,N_38371);
nand U44188 (N_44188,N_36827,N_36477);
nor U44189 (N_44189,N_30623,N_33457);
or U44190 (N_44190,N_39895,N_35231);
nand U44191 (N_44191,N_38770,N_35553);
nor U44192 (N_44192,N_33527,N_36554);
nand U44193 (N_44193,N_33931,N_33986);
nand U44194 (N_44194,N_32511,N_34366);
and U44195 (N_44195,N_37677,N_37461);
and U44196 (N_44196,N_33165,N_39840);
nor U44197 (N_44197,N_37570,N_33948);
nor U44198 (N_44198,N_33964,N_31250);
nand U44199 (N_44199,N_38435,N_31939);
nor U44200 (N_44200,N_34305,N_38434);
nand U44201 (N_44201,N_31872,N_34148);
nor U44202 (N_44202,N_31789,N_39354);
nand U44203 (N_44203,N_38062,N_38500);
nor U44204 (N_44204,N_30768,N_39678);
nor U44205 (N_44205,N_32805,N_34221);
and U44206 (N_44206,N_35744,N_38225);
nand U44207 (N_44207,N_31011,N_33937);
nand U44208 (N_44208,N_39163,N_30332);
nor U44209 (N_44209,N_35229,N_31700);
nand U44210 (N_44210,N_39626,N_30879);
and U44211 (N_44211,N_33636,N_37587);
xnor U44212 (N_44212,N_36254,N_35658);
or U44213 (N_44213,N_36538,N_37691);
or U44214 (N_44214,N_35604,N_37176);
and U44215 (N_44215,N_38229,N_39807);
xor U44216 (N_44216,N_35821,N_30045);
nand U44217 (N_44217,N_33916,N_33285);
and U44218 (N_44218,N_30770,N_30096);
xnor U44219 (N_44219,N_33891,N_35409);
and U44220 (N_44220,N_36556,N_35850);
or U44221 (N_44221,N_39624,N_32363);
or U44222 (N_44222,N_33158,N_34427);
nand U44223 (N_44223,N_32011,N_37257);
nand U44224 (N_44224,N_33656,N_38655);
xor U44225 (N_44225,N_31569,N_33878);
or U44226 (N_44226,N_31695,N_39198);
nor U44227 (N_44227,N_33310,N_33498);
or U44228 (N_44228,N_30493,N_30188);
and U44229 (N_44229,N_36857,N_39134);
nor U44230 (N_44230,N_36691,N_38360);
and U44231 (N_44231,N_35420,N_30515);
nor U44232 (N_44232,N_34043,N_34752);
or U44233 (N_44233,N_30430,N_38850);
or U44234 (N_44234,N_30379,N_33591);
nor U44235 (N_44235,N_32243,N_36127);
nand U44236 (N_44236,N_37008,N_34549);
nand U44237 (N_44237,N_30657,N_31856);
and U44238 (N_44238,N_36381,N_39790);
nand U44239 (N_44239,N_31167,N_39446);
or U44240 (N_44240,N_35099,N_33244);
nand U44241 (N_44241,N_32604,N_31043);
nor U44242 (N_44242,N_34213,N_37063);
xor U44243 (N_44243,N_36668,N_38907);
and U44244 (N_44244,N_37452,N_33047);
or U44245 (N_44245,N_37960,N_37564);
and U44246 (N_44246,N_35474,N_37866);
nor U44247 (N_44247,N_32087,N_34506);
and U44248 (N_44248,N_39421,N_30387);
or U44249 (N_44249,N_36700,N_34833);
and U44250 (N_44250,N_33660,N_39617);
or U44251 (N_44251,N_35509,N_35692);
xor U44252 (N_44252,N_38193,N_39295);
or U44253 (N_44253,N_32661,N_30919);
or U44254 (N_44254,N_38405,N_37528);
xor U44255 (N_44255,N_30427,N_31791);
nor U44256 (N_44256,N_33256,N_36746);
and U44257 (N_44257,N_30028,N_35467);
nand U44258 (N_44258,N_36059,N_32122);
nor U44259 (N_44259,N_30513,N_39820);
and U44260 (N_44260,N_38704,N_39757);
nor U44261 (N_44261,N_37363,N_33647);
nand U44262 (N_44262,N_34744,N_35857);
and U44263 (N_44263,N_32803,N_36116);
and U44264 (N_44264,N_32686,N_33699);
xor U44265 (N_44265,N_38577,N_30951);
or U44266 (N_44266,N_30702,N_39493);
nand U44267 (N_44267,N_35263,N_31888);
or U44268 (N_44268,N_32589,N_34630);
nor U44269 (N_44269,N_34471,N_38463);
xor U44270 (N_44270,N_35048,N_31958);
nand U44271 (N_44271,N_31255,N_35873);
nor U44272 (N_44272,N_30473,N_36625);
xnor U44273 (N_44273,N_37032,N_31017);
or U44274 (N_44274,N_30872,N_31053);
nand U44275 (N_44275,N_36078,N_33923);
xor U44276 (N_44276,N_34057,N_39857);
nand U44277 (N_44277,N_38698,N_37161);
or U44278 (N_44278,N_37850,N_36838);
or U44279 (N_44279,N_36927,N_35408);
or U44280 (N_44280,N_37573,N_32786);
and U44281 (N_44281,N_32000,N_33114);
xnor U44282 (N_44282,N_38439,N_33449);
nand U44283 (N_44283,N_31334,N_32898);
nand U44284 (N_44284,N_30912,N_36790);
and U44285 (N_44285,N_35021,N_34945);
nor U44286 (N_44286,N_37277,N_31201);
xor U44287 (N_44287,N_33003,N_31014);
nor U44288 (N_44288,N_30892,N_30360);
nor U44289 (N_44289,N_38255,N_37351);
xor U44290 (N_44290,N_33533,N_30098);
and U44291 (N_44291,N_39000,N_37543);
or U44292 (N_44292,N_31022,N_35745);
and U44293 (N_44293,N_32261,N_39058);
and U44294 (N_44294,N_39297,N_34363);
nor U44295 (N_44295,N_32147,N_36453);
and U44296 (N_44296,N_39993,N_35742);
nor U44297 (N_44297,N_31077,N_38726);
nand U44298 (N_44298,N_33545,N_39540);
or U44299 (N_44299,N_34538,N_34146);
nor U44300 (N_44300,N_34999,N_30523);
or U44301 (N_44301,N_32989,N_35702);
nand U44302 (N_44302,N_30828,N_36965);
and U44303 (N_44303,N_32652,N_30885);
nand U44304 (N_44304,N_32234,N_32813);
and U44305 (N_44305,N_32298,N_35126);
and U44306 (N_44306,N_36774,N_39673);
nor U44307 (N_44307,N_30066,N_37482);
and U44308 (N_44308,N_35078,N_37372);
nand U44309 (N_44309,N_39348,N_38723);
and U44310 (N_44310,N_33157,N_37247);
nor U44311 (N_44311,N_35528,N_35853);
and U44312 (N_44312,N_34349,N_30243);
or U44313 (N_44313,N_38742,N_37334);
or U44314 (N_44314,N_36096,N_38956);
or U44315 (N_44315,N_35895,N_39565);
nor U44316 (N_44316,N_39593,N_35691);
or U44317 (N_44317,N_37104,N_35956);
and U44318 (N_44318,N_37227,N_32789);
xnor U44319 (N_44319,N_35859,N_30070);
and U44320 (N_44320,N_38176,N_32644);
nor U44321 (N_44321,N_31935,N_35833);
or U44322 (N_44322,N_34345,N_36871);
nand U44323 (N_44323,N_35224,N_37777);
and U44324 (N_44324,N_38031,N_34772);
or U44325 (N_44325,N_31934,N_36563);
and U44326 (N_44326,N_33531,N_35311);
or U44327 (N_44327,N_35712,N_30112);
nand U44328 (N_44328,N_39838,N_31590);
and U44329 (N_44329,N_36869,N_36103);
nand U44330 (N_44330,N_32551,N_38664);
and U44331 (N_44331,N_32566,N_31985);
nor U44332 (N_44332,N_33707,N_31744);
nor U44333 (N_44333,N_39722,N_31134);
and U44334 (N_44334,N_36089,N_32871);
or U44335 (N_44335,N_34811,N_37760);
and U44336 (N_44336,N_31884,N_35977);
and U44337 (N_44337,N_37996,N_38913);
xnor U44338 (N_44338,N_34346,N_32708);
xnor U44339 (N_44339,N_36759,N_30929);
or U44340 (N_44340,N_36113,N_34308);
nor U44341 (N_44341,N_31863,N_31596);
nor U44342 (N_44342,N_30034,N_38185);
or U44343 (N_44343,N_38900,N_30063);
or U44344 (N_44344,N_35275,N_34737);
nor U44345 (N_44345,N_35272,N_34946);
or U44346 (N_44346,N_31345,N_31816);
and U44347 (N_44347,N_38203,N_30313);
nand U44348 (N_44348,N_37096,N_32331);
nand U44349 (N_44349,N_38607,N_32452);
and U44350 (N_44350,N_39485,N_38213);
nand U44351 (N_44351,N_33319,N_33588);
xnor U44352 (N_44352,N_37204,N_36463);
or U44353 (N_44353,N_34719,N_30746);
nand U44354 (N_44354,N_32396,N_39883);
nand U44355 (N_44355,N_38048,N_32142);
nand U44356 (N_44356,N_35332,N_30091);
nand U44357 (N_44357,N_34355,N_32154);
or U44358 (N_44358,N_32042,N_38386);
nor U44359 (N_44359,N_33814,N_34622);
and U44360 (N_44360,N_31783,N_37525);
nand U44361 (N_44361,N_39098,N_31459);
and U44362 (N_44362,N_31313,N_39153);
nand U44363 (N_44363,N_35385,N_32856);
xor U44364 (N_44364,N_32082,N_36027);
nor U44365 (N_44365,N_33594,N_30437);
and U44366 (N_44366,N_37728,N_36719);
nor U44367 (N_44367,N_36033,N_30044);
nand U44368 (N_44368,N_38286,N_38690);
nor U44369 (N_44369,N_31056,N_39736);
nand U44370 (N_44370,N_37756,N_33426);
xnor U44371 (N_44371,N_37447,N_39546);
or U44372 (N_44372,N_36182,N_33899);
nor U44373 (N_44373,N_36202,N_34952);
xor U44374 (N_44374,N_38686,N_30476);
nor U44375 (N_44375,N_30423,N_36278);
xnor U44376 (N_44376,N_39817,N_38438);
and U44377 (N_44377,N_32522,N_33140);
xnor U44378 (N_44378,N_33800,N_37411);
or U44379 (N_44379,N_32549,N_32694);
and U44380 (N_44380,N_37454,N_33022);
xor U44381 (N_44381,N_37300,N_37325);
nor U44382 (N_44382,N_33180,N_34570);
nand U44383 (N_44383,N_35714,N_30844);
or U44384 (N_44384,N_36628,N_36382);
or U44385 (N_44385,N_35480,N_34054);
or U44386 (N_44386,N_37765,N_33181);
and U44387 (N_44387,N_37378,N_34448);
and U44388 (N_44388,N_33436,N_31042);
nor U44389 (N_44389,N_38676,N_32337);
nor U44390 (N_44390,N_39649,N_39611);
nor U44391 (N_44391,N_37210,N_33850);
nor U44392 (N_44392,N_38332,N_30868);
and U44393 (N_44393,N_38511,N_38647);
or U44394 (N_44394,N_30017,N_32149);
nor U44395 (N_44395,N_36451,N_34526);
xor U44396 (N_44396,N_30712,N_30954);
nand U44397 (N_44397,N_36189,N_39702);
or U44398 (N_44398,N_30385,N_38926);
or U44399 (N_44399,N_37953,N_36008);
and U44400 (N_44400,N_31111,N_36656);
or U44401 (N_44401,N_32677,N_35456);
nand U44402 (N_44402,N_31118,N_30838);
nand U44403 (N_44403,N_37813,N_38258);
nand U44404 (N_44404,N_38824,N_39329);
or U44405 (N_44405,N_38137,N_30726);
and U44406 (N_44406,N_30563,N_36309);
or U44407 (N_44407,N_31347,N_32773);
nor U44408 (N_44408,N_31398,N_31854);
and U44409 (N_44409,N_32905,N_35228);
nor U44410 (N_44410,N_34497,N_30160);
nor U44411 (N_44411,N_39940,N_37427);
nor U44412 (N_44412,N_34836,N_38478);
nand U44413 (N_44413,N_35302,N_32151);
and U44414 (N_44414,N_36405,N_30462);
and U44415 (N_44415,N_30178,N_37458);
nor U44416 (N_44416,N_36342,N_39156);
or U44417 (N_44417,N_33071,N_31519);
and U44418 (N_44418,N_37588,N_36861);
nor U44419 (N_44419,N_32895,N_33590);
nand U44420 (N_44420,N_38269,N_30983);
nor U44421 (N_44421,N_38138,N_34077);
and U44422 (N_44422,N_34488,N_39039);
nand U44423 (N_44423,N_33078,N_38469);
nand U44424 (N_44424,N_38397,N_37438);
or U44425 (N_44425,N_37717,N_37927);
or U44426 (N_44426,N_34621,N_38428);
nor U44427 (N_44427,N_37789,N_36977);
nand U44428 (N_44428,N_30756,N_30057);
nand U44429 (N_44429,N_34294,N_39989);
or U44430 (N_44430,N_34493,N_30074);
and U44431 (N_44431,N_32381,N_35248);
nor U44432 (N_44432,N_31953,N_30418);
nor U44433 (N_44433,N_31970,N_39564);
and U44434 (N_44434,N_37853,N_33039);
and U44435 (N_44435,N_35900,N_30264);
or U44436 (N_44436,N_39830,N_37945);
nor U44437 (N_44437,N_39777,N_37201);
and U44438 (N_44438,N_33547,N_34989);
nor U44439 (N_44439,N_35920,N_31885);
xnor U44440 (N_44440,N_39874,N_35945);
nor U44441 (N_44441,N_34769,N_35091);
and U44442 (N_44442,N_33155,N_33381);
or U44443 (N_44443,N_34860,N_34490);
or U44444 (N_44444,N_35599,N_37392);
or U44445 (N_44445,N_31054,N_33384);
xor U44446 (N_44446,N_33446,N_34045);
or U44447 (N_44447,N_36847,N_32335);
nand U44448 (N_44448,N_37466,N_39808);
or U44449 (N_44449,N_37118,N_31122);
nand U44450 (N_44450,N_37178,N_33506);
nor U44451 (N_44451,N_33009,N_39770);
nand U44452 (N_44452,N_33420,N_36611);
xor U44453 (N_44453,N_36992,N_37076);
and U44454 (N_44454,N_33556,N_31682);
nor U44455 (N_44455,N_31229,N_33870);
nor U44456 (N_44456,N_31894,N_37550);
nand U44457 (N_44457,N_39753,N_39081);
nor U44458 (N_44458,N_36490,N_32966);
xor U44459 (N_44459,N_30337,N_33838);
nand U44460 (N_44460,N_37666,N_32153);
nor U44461 (N_44461,N_33343,N_36596);
nor U44462 (N_44462,N_36249,N_31670);
and U44463 (N_44463,N_33404,N_32754);
nor U44464 (N_44464,N_35131,N_39313);
nor U44465 (N_44465,N_31750,N_35585);
xor U44466 (N_44466,N_31529,N_38501);
xor U44467 (N_44467,N_39014,N_39787);
nand U44468 (N_44468,N_31021,N_30664);
and U44469 (N_44469,N_35396,N_30080);
or U44470 (N_44470,N_36798,N_36011);
or U44471 (N_44471,N_35699,N_38378);
nand U44472 (N_44472,N_31539,N_36393);
or U44473 (N_44473,N_32301,N_38262);
and U44474 (N_44474,N_36041,N_34874);
or U44475 (N_44475,N_31948,N_36589);
or U44476 (N_44476,N_33727,N_34666);
nand U44477 (N_44477,N_30269,N_32590);
or U44478 (N_44478,N_39921,N_36536);
and U44479 (N_44479,N_36444,N_35889);
nand U44480 (N_44480,N_35378,N_32453);
or U44481 (N_44481,N_36435,N_32801);
nor U44482 (N_44482,N_34645,N_34600);
nor U44483 (N_44483,N_39072,N_38819);
nor U44484 (N_44484,N_30317,N_31874);
or U44485 (N_44485,N_31128,N_32119);
nor U44486 (N_44486,N_32216,N_34516);
and U44487 (N_44487,N_38765,N_33295);
nand U44488 (N_44488,N_30897,N_30442);
nand U44489 (N_44489,N_34416,N_39547);
or U44490 (N_44490,N_32403,N_33380);
nor U44491 (N_44491,N_33481,N_39505);
nand U44492 (N_44492,N_30963,N_36680);
and U44493 (N_44493,N_33648,N_36071);
nand U44494 (N_44494,N_33382,N_38318);
or U44495 (N_44495,N_30217,N_33159);
or U44496 (N_44496,N_31797,N_39087);
and U44497 (N_44497,N_30174,N_30016);
nor U44498 (N_44498,N_36768,N_36533);
or U44499 (N_44499,N_37797,N_39012);
nor U44500 (N_44500,N_34038,N_33198);
nand U44501 (N_44501,N_36268,N_34969);
nor U44502 (N_44502,N_39415,N_35152);
and U44503 (N_44503,N_33580,N_38433);
nand U44504 (N_44504,N_31629,N_35030);
or U44505 (N_44505,N_33440,N_39379);
xnor U44506 (N_44506,N_32088,N_39925);
and U44507 (N_44507,N_37191,N_31633);
and U44508 (N_44508,N_37278,N_31703);
nor U44509 (N_44509,N_33136,N_31490);
and U44510 (N_44510,N_32325,N_30159);
xor U44511 (N_44511,N_37946,N_38715);
xor U44512 (N_44512,N_31548,N_36077);
xor U44513 (N_44513,N_39518,N_32405);
xnor U44514 (N_44514,N_35122,N_36621);
nand U44515 (N_44515,N_31454,N_31214);
xor U44516 (N_44516,N_37939,N_36661);
or U44517 (N_44517,N_36512,N_34560);
nand U44518 (N_44518,N_32714,N_35701);
nor U44519 (N_44519,N_30877,N_32980);
and U44520 (N_44520,N_33249,N_31527);
nand U44521 (N_44521,N_37241,N_37159);
nand U44522 (N_44522,N_35389,N_31087);
and U44523 (N_44523,N_31107,N_33268);
nand U44524 (N_44524,N_35634,N_31147);
or U44525 (N_44525,N_39999,N_31646);
or U44526 (N_44526,N_36513,N_35148);
and U44527 (N_44527,N_35353,N_37399);
or U44528 (N_44528,N_30033,N_35998);
nor U44529 (N_44529,N_35169,N_33448);
and U44530 (N_44530,N_35250,N_32366);
and U44531 (N_44531,N_32457,N_32983);
or U44532 (N_44532,N_35102,N_37039);
or U44533 (N_44533,N_37426,N_35256);
nor U44534 (N_44534,N_36900,N_30748);
or U44535 (N_44535,N_31844,N_32958);
and U44536 (N_44536,N_36063,N_38739);
and U44537 (N_44537,N_31502,N_33451);
or U44538 (N_44538,N_31655,N_33289);
and U44539 (N_44539,N_34716,N_34373);
nor U44540 (N_44540,N_37702,N_34227);
nand U44541 (N_44541,N_36835,N_39369);
and U44542 (N_44542,N_35295,N_30361);
xor U44543 (N_44543,N_33743,N_35593);
nand U44544 (N_44544,N_30294,N_34815);
xor U44545 (N_44545,N_36739,N_39191);
xnor U44546 (N_44546,N_37619,N_30331);
or U44547 (N_44547,N_37676,N_34821);
and U44548 (N_44548,N_33237,N_33791);
and U44549 (N_44549,N_36084,N_30138);
and U44550 (N_44550,N_34683,N_39315);
nand U44551 (N_44551,N_37455,N_32406);
xnor U44552 (N_44552,N_33595,N_36955);
nor U44553 (N_44553,N_34306,N_35216);
and U44554 (N_44554,N_35123,N_34030);
or U44555 (N_44555,N_39150,N_37146);
or U44556 (N_44556,N_32404,N_31083);
and U44557 (N_44557,N_31790,N_31177);
nand U44558 (N_44558,N_32543,N_38417);
nand U44559 (N_44559,N_33400,N_30413);
or U44560 (N_44560,N_34344,N_37068);
or U44561 (N_44561,N_34090,N_38534);
nor U44562 (N_44562,N_32936,N_30831);
nor U44563 (N_44563,N_37266,N_38310);
nor U44564 (N_44564,N_32808,N_33064);
nand U44565 (N_44565,N_39837,N_37481);
or U44566 (N_44566,N_39668,N_39448);
nand U44567 (N_44567,N_30700,N_32663);
nand U44568 (N_44568,N_35204,N_39748);
and U44569 (N_44569,N_39030,N_35561);
nor U44570 (N_44570,N_31066,N_30117);
or U44571 (N_44571,N_37243,N_30744);
nor U44572 (N_44572,N_35313,N_34083);
nand U44573 (N_44573,N_39140,N_36409);
nor U44574 (N_44574,N_36804,N_36447);
nor U44575 (N_44575,N_38270,N_34743);
nand U44576 (N_44576,N_32595,N_33148);
xor U44577 (N_44577,N_39468,N_37832);
or U44578 (N_44578,N_34152,N_37339);
or U44579 (N_44579,N_33741,N_30157);
or U44580 (N_44580,N_30745,N_36443);
nor U44581 (N_44581,N_34050,N_37663);
or U44582 (N_44582,N_30231,N_38312);
and U44583 (N_44583,N_38473,N_36811);
xor U44584 (N_44584,N_36307,N_38197);
nand U44585 (N_44585,N_32957,N_39930);
nor U44586 (N_44586,N_38391,N_30596);
nor U44587 (N_44587,N_35281,N_38129);
xor U44588 (N_44588,N_35101,N_37864);
nor U44589 (N_44589,N_32257,N_33659);
or U44590 (N_44590,N_37175,N_32183);
or U44591 (N_44591,N_30884,N_36034);
nand U44592 (N_44592,N_36953,N_30380);
xor U44593 (N_44593,N_32512,N_30797);
and U44594 (N_44594,N_32934,N_36770);
nand U44595 (N_44595,N_35438,N_32002);
nor U44596 (N_44596,N_36184,N_36630);
or U44597 (N_44597,N_39335,N_36174);
or U44598 (N_44598,N_37288,N_36310);
nand U44599 (N_44599,N_31325,N_33752);
nor U44600 (N_44600,N_33402,N_37362);
xor U44601 (N_44601,N_37330,N_33335);
and U44602 (N_44602,N_30840,N_30226);
nor U44603 (N_44603,N_39353,N_39704);
nand U44604 (N_44604,N_31637,N_31272);
and U44605 (N_44605,N_36048,N_39162);
xnor U44606 (N_44606,N_30295,N_34179);
nor U44607 (N_44607,N_34499,N_33762);
nor U44608 (N_44608,N_30245,N_35541);
or U44609 (N_44609,N_30407,N_32715);
nor U44610 (N_44610,N_38064,N_39934);
nor U44611 (N_44611,N_34541,N_37593);
nor U44612 (N_44612,N_30504,N_37714);
and U44613 (N_44613,N_38874,N_36677);
xnor U44614 (N_44614,N_38639,N_35271);
or U44615 (N_44615,N_38486,N_38305);
nor U44616 (N_44616,N_36837,N_31073);
nand U44617 (N_44617,N_31805,N_31019);
or U44618 (N_44618,N_38923,N_32609);
nand U44619 (N_44619,N_31585,N_38503);
nand U44620 (N_44620,N_38278,N_30422);
xor U44621 (N_44621,N_39242,N_38727);
and U44622 (N_44622,N_37219,N_32375);
and U44623 (N_44623,N_32192,N_35266);
and U44624 (N_44624,N_36542,N_38984);
and U44625 (N_44625,N_39009,N_31715);
nand U44626 (N_44626,N_33082,N_39118);
and U44627 (N_44627,N_38866,N_33454);
or U44628 (N_44628,N_36156,N_37630);
and U44629 (N_44629,N_33066,N_38089);
xnor U44630 (N_44630,N_35901,N_34175);
and U44631 (N_44631,N_30496,N_30085);
nand U44632 (N_44632,N_35884,N_35942);
or U44633 (N_44633,N_31656,N_31615);
or U44634 (N_44634,N_36049,N_35269);
nor U44635 (N_44635,N_37638,N_37594);
nor U44636 (N_44636,N_33757,N_30546);
xnor U44637 (N_44637,N_39210,N_37084);
or U44638 (N_44638,N_34655,N_38247);
and U44639 (N_44639,N_39526,N_33055);
nor U44640 (N_44640,N_32844,N_37408);
or U44641 (N_44641,N_33991,N_39610);
nor U44642 (N_44642,N_32182,N_38524);
and U44643 (N_44643,N_36203,N_33905);
or U44644 (N_44644,N_30800,N_38017);
and U44645 (N_44645,N_37070,N_32606);
nand U44646 (N_44646,N_35405,N_39074);
and U44647 (N_44647,N_32727,N_36065);
nor U44648 (N_44648,N_35657,N_31142);
and U44649 (N_44649,N_35979,N_39224);
nand U44650 (N_44650,N_31284,N_35466);
and U44651 (N_44651,N_36123,N_32791);
nand U44652 (N_44652,N_38814,N_37059);
nor U44653 (N_44653,N_36752,N_32332);
nor U44654 (N_44654,N_34679,N_31096);
xnor U44655 (N_44655,N_35952,N_35995);
xor U44656 (N_44656,N_39798,N_38755);
and U44657 (N_44657,N_31093,N_37149);
and U44658 (N_44658,N_32968,N_33742);
and U44659 (N_44659,N_38165,N_35251);
and U44660 (N_44660,N_36132,N_33859);
nand U44661 (N_44661,N_39538,N_34049);
nand U44662 (N_44662,N_35856,N_39816);
nor U44663 (N_44663,N_31658,N_36581);
and U44664 (N_44664,N_32031,N_38633);
nor U44665 (N_44665,N_32445,N_36395);
nor U44666 (N_44666,N_36496,N_33926);
or U44667 (N_44667,N_33354,N_34788);
nor U44668 (N_44668,N_30661,N_37239);
nand U44669 (N_44669,N_35223,N_36687);
nand U44670 (N_44670,N_34399,N_34684);
nor U44671 (N_44671,N_38560,N_37307);
nand U44672 (N_44672,N_33907,N_38927);
or U44673 (N_44673,N_31736,N_30860);
and U44674 (N_44674,N_32166,N_37531);
nand U44675 (N_44675,N_32524,N_34321);
nand U44676 (N_44676,N_36858,N_33084);
nor U44677 (N_44677,N_31751,N_39236);
xnor U44678 (N_44678,N_30729,N_39414);
nor U44679 (N_44679,N_33430,N_37302);
nand U44680 (N_44680,N_30535,N_30908);
or U44681 (N_44681,N_39543,N_38303);
or U44682 (N_44682,N_38353,N_38733);
nor U44683 (N_44683,N_30572,N_32386);
nand U44684 (N_44684,N_32401,N_36863);
or U44685 (N_44685,N_36284,N_31079);
nor U44686 (N_44686,N_32929,N_36833);
nor U44687 (N_44687,N_39542,N_37453);
nand U44688 (N_44688,N_39106,N_39338);
or U44689 (N_44689,N_39983,N_35603);
or U44690 (N_44690,N_32897,N_32635);
and U44691 (N_44691,N_36446,N_38683);
nand U44692 (N_44692,N_34961,N_34936);
xnor U44693 (N_44693,N_32194,N_31426);
or U44694 (N_44694,N_34937,N_30244);
nor U44695 (N_44695,N_35062,N_35950);
nand U44696 (N_44696,N_32517,N_35437);
nand U44697 (N_44697,N_35208,N_32291);
nand U44698 (N_44698,N_33111,N_33534);
xor U44699 (N_44699,N_35729,N_39443);
xor U44700 (N_44700,N_35086,N_34438);
and U44701 (N_44701,N_38419,N_36352);
and U44702 (N_44702,N_32374,N_36999);
nand U44703 (N_44703,N_33921,N_37462);
and U44704 (N_44704,N_37365,N_35215);
and U44705 (N_44705,N_37420,N_33484);
nand U44706 (N_44706,N_32990,N_38702);
and U44707 (N_44707,N_32041,N_37612);
nand U44708 (N_44708,N_37433,N_34798);
and U44709 (N_44709,N_35549,N_31184);
nor U44710 (N_44710,N_39197,N_38760);
or U44711 (N_44711,N_33423,N_39535);
and U44712 (N_44712,N_39342,N_34890);
or U44713 (N_44713,N_38015,N_36731);
nand U44714 (N_44714,N_39473,N_30312);
xnor U44715 (N_44715,N_31424,N_38464);
nand U44716 (N_44716,N_30524,N_30114);
and U44717 (N_44717,N_38827,N_35751);
nand U44718 (N_44718,N_30857,N_39442);
and U44719 (N_44719,N_35276,N_31676);
nand U44720 (N_44720,N_35166,N_34201);
nor U44721 (N_44721,N_35638,N_34700);
nand U44722 (N_44722,N_39600,N_33075);
and U44723 (N_44723,N_37558,N_35260);
nand U44724 (N_44724,N_30251,N_37727);
and U44725 (N_44725,N_36325,N_35774);
nor U44726 (N_44726,N_36167,N_33372);
nor U44727 (N_44727,N_39282,N_38744);
nor U44728 (N_44728,N_32868,N_38893);
nor U44729 (N_44729,N_36260,N_34584);
nor U44730 (N_44730,N_36458,N_32235);
nor U44731 (N_44731,N_30454,N_30776);
nand U44732 (N_44732,N_30614,N_36957);
nand U44733 (N_44733,N_39283,N_33144);
or U44734 (N_44734,N_32931,N_34153);
nor U44735 (N_44735,N_35182,N_30721);
or U44736 (N_44736,N_33603,N_39291);
nand U44737 (N_44737,N_30953,N_34188);
and U44738 (N_44738,N_37382,N_31870);
nand U44739 (N_44739,N_32893,N_33571);
nand U44740 (N_44740,N_34458,N_38659);
nor U44741 (N_44741,N_37957,N_34765);
or U44742 (N_44742,N_32586,N_39833);
and U44743 (N_44743,N_35819,N_35595);
xor U44744 (N_44744,N_31210,N_30709);
nand U44745 (N_44745,N_38413,N_32263);
nor U44746 (N_44746,N_37470,N_39920);
nor U44747 (N_44747,N_30635,N_30394);
and U44748 (N_44748,N_35218,N_32537);
nor U44749 (N_44749,N_34579,N_39908);
xor U44750 (N_44750,N_36288,N_36371);
and U44751 (N_44751,N_37421,N_35570);
nor U44752 (N_44752,N_35452,N_33170);
nor U44753 (N_44753,N_32304,N_34094);
xor U44754 (N_44754,N_32949,N_37655);
nor U44755 (N_44755,N_37298,N_32855);
nand U44756 (N_44756,N_37016,N_33680);
or U44757 (N_44757,N_35301,N_34812);
nor U44758 (N_44758,N_34206,N_30825);
or U44759 (N_44759,N_35782,N_34599);
nand U44760 (N_44760,N_38307,N_38730);
or U44761 (N_44761,N_32203,N_34078);
nand U44762 (N_44762,N_31491,N_30845);
nand U44763 (N_44763,N_33088,N_39814);
and U44764 (N_44764,N_37053,N_37784);
or U44765 (N_44765,N_33490,N_36017);
or U44766 (N_44766,N_35866,N_31342);
nand U44767 (N_44767,N_38044,N_39093);
nand U44768 (N_44768,N_35417,N_33257);
nand U44769 (N_44769,N_35345,N_34328);
nand U44770 (N_44770,N_35305,N_35876);
and U44771 (N_44771,N_39963,N_34817);
nand U44772 (N_44772,N_38801,N_37217);
nor U44773 (N_44773,N_36696,N_31583);
nand U44774 (N_44774,N_35618,N_30628);
or U44775 (N_44775,N_36970,N_34479);
xor U44776 (N_44776,N_33963,N_30088);
or U44777 (N_44777,N_32744,N_38429);
nor U44778 (N_44778,N_31389,N_30363);
nor U44779 (N_44779,N_34091,N_31428);
nand U44780 (N_44780,N_31567,N_35013);
nor U44781 (N_44781,N_37223,N_39382);
or U44782 (N_44782,N_31013,N_34568);
nand U44783 (N_44783,N_31746,N_38734);
nand U44784 (N_44784,N_32506,N_33028);
xor U44785 (N_44785,N_32448,N_34756);
nand U44786 (N_44786,N_34713,N_33823);
and U44787 (N_44787,N_34319,N_31238);
nand U44788 (N_44788,N_31244,N_30306);
and U44789 (N_44789,N_39524,N_36709);
nor U44790 (N_44790,N_34971,N_36727);
nand U44791 (N_44791,N_36346,N_38497);
and U44792 (N_44792,N_33557,N_38971);
and U44793 (N_44793,N_39590,N_38084);
or U44794 (N_44794,N_36211,N_36036);
or U44795 (N_44795,N_35496,N_31731);
nor U44796 (N_44796,N_36213,N_39107);
or U44797 (N_44797,N_36082,N_30225);
nand U44798 (N_44798,N_33018,N_37534);
and U44799 (N_44799,N_37472,N_31899);
or U44800 (N_44800,N_36403,N_36978);
xor U44801 (N_44801,N_35070,N_38239);
or U44802 (N_44802,N_30737,N_37628);
and U44803 (N_44803,N_37640,N_32106);
and U44804 (N_44804,N_34436,N_34960);
nand U44805 (N_44805,N_31270,N_30506);
nand U44806 (N_44806,N_30511,N_36984);
nor U44807 (N_44807,N_32662,N_31965);
nand U44808 (N_44808,N_32416,N_30979);
or U44809 (N_44809,N_30381,N_31336);
and U44810 (N_44810,N_30150,N_36688);
nand U44811 (N_44811,N_38257,N_32334);
nand U44812 (N_44812,N_32573,N_30148);
nand U44813 (N_44813,N_34205,N_30625);
nor U44814 (N_44814,N_30615,N_30019);
or U44815 (N_44815,N_35867,N_37413);
or U44816 (N_44816,N_35413,N_37196);
nand U44817 (N_44817,N_38864,N_37911);
or U44818 (N_44818,N_37206,N_36037);
and U44819 (N_44819,N_36467,N_31581);
or U44820 (N_44820,N_31451,N_39256);
nand U44821 (N_44821,N_32419,N_39915);
or U44822 (N_44822,N_30018,N_35844);
nor U44823 (N_44823,N_33607,N_30626);
and U44824 (N_44824,N_32757,N_31626);
nor U44825 (N_44825,N_38181,N_39620);
or U44826 (N_44826,N_38580,N_37710);
and U44827 (N_44827,N_33638,N_36705);
or U44828 (N_44828,N_33328,N_31427);
and U44829 (N_44829,N_35201,N_36515);
or U44830 (N_44830,N_30899,N_39206);
nor U44831 (N_44831,N_34601,N_34674);
nor U44832 (N_44832,N_39806,N_31574);
and U44833 (N_44833,N_34066,N_31993);
nor U44834 (N_44834,N_34081,N_38860);
or U44835 (N_44835,N_39172,N_37398);
or U44836 (N_44836,N_39043,N_33122);
and U44837 (N_44837,N_39507,N_38456);
nand U44838 (N_44838,N_39082,N_37379);
or U44839 (N_44839,N_38590,N_35526);
and U44840 (N_44840,N_36119,N_35172);
and U44841 (N_44841,N_32875,N_35446);
or U44842 (N_44842,N_35847,N_39504);
and U44843 (N_44843,N_32101,N_33048);
and U44844 (N_44844,N_30945,N_32177);
nand U44845 (N_44845,N_32319,N_32264);
and U44846 (N_44846,N_33016,N_36878);
or U44847 (N_44847,N_35891,N_31898);
and U44848 (N_44848,N_36394,N_39432);
and U44849 (N_44849,N_38569,N_32038);
or U44850 (N_44850,N_36894,N_32089);
nor U44851 (N_44851,N_31438,N_30990);
nand U44852 (N_44852,N_34562,N_30238);
nand U44853 (N_44853,N_38201,N_36101);
nand U44854 (N_44854,N_30531,N_33829);
or U44855 (N_44855,N_32323,N_32702);
nor U44856 (N_44856,N_31033,N_36317);
nor U44857 (N_44857,N_32842,N_34802);
nor U44858 (N_44858,N_34127,N_35806);
or U44859 (N_44859,N_32473,N_39445);
xnor U44860 (N_44860,N_37018,N_39839);
and U44861 (N_44861,N_34395,N_35989);
or U44862 (N_44862,N_32251,N_38359);
or U44863 (N_44863,N_39292,N_34746);
or U44864 (N_44864,N_31366,N_37354);
and U44865 (N_44865,N_35384,N_31382);
and U44866 (N_44866,N_31510,N_31624);
and U44867 (N_44867,N_36923,N_39594);
and U44868 (N_44868,N_34456,N_39716);
or U44869 (N_44869,N_38072,N_31499);
or U44870 (N_44870,N_30133,N_31662);
or U44871 (N_44871,N_32321,N_36012);
and U44872 (N_44872,N_37752,N_31853);
nand U44873 (N_44873,N_38409,N_31514);
or U44874 (N_44874,N_34189,N_30920);
xor U44875 (N_44875,N_32814,N_39294);
nand U44876 (N_44876,N_33087,N_35882);
xor U44877 (N_44877,N_34379,N_37460);
nand U44878 (N_44878,N_35838,N_32660);
or U44879 (N_44879,N_37368,N_32409);
or U44880 (N_44880,N_34805,N_34387);
and U44881 (N_44881,N_38679,N_34823);
xnor U44882 (N_44882,N_30483,N_39865);
nor U44883 (N_44883,N_30542,N_38588);
nand U44884 (N_44884,N_36778,N_36735);
nand U44885 (N_44885,N_39100,N_38696);
nor U44886 (N_44886,N_30586,N_30107);
and U44887 (N_44887,N_32399,N_35232);
and U44888 (N_44888,N_36277,N_30497);
nand U44889 (N_44889,N_37431,N_32481);
and U44890 (N_44890,N_32433,N_34194);
and U44891 (N_44891,N_37707,N_30448);
and U44892 (N_44892,N_32208,N_36215);
nand U44893 (N_44893,N_35530,N_31591);
xor U44894 (N_44894,N_33231,N_31573);
and U44895 (N_44895,N_38060,N_31571);
nor U44896 (N_44896,N_36233,N_30688);
nand U44897 (N_44897,N_39333,N_36506);
and U44898 (N_44898,N_30291,N_36177);
nand U44899 (N_44899,N_38452,N_39699);
nor U44900 (N_44900,N_33428,N_39882);
nor U44901 (N_44901,N_37291,N_38294);
and U44902 (N_44902,N_31146,N_30500);
nor U44903 (N_44903,N_31553,N_33749);
and U44904 (N_44904,N_33713,N_33292);
nand U44905 (N_44905,N_39086,N_39487);
and U44906 (N_44906,N_38187,N_37401);
nor U44907 (N_44907,N_31004,N_30494);
and U44908 (N_44908,N_33717,N_36354);
nand U44909 (N_44909,N_31194,N_34915);
and U44910 (N_44910,N_31501,N_30769);
and U44911 (N_44911,N_37969,N_30039);
nor U44912 (N_44912,N_39232,N_38957);
xnor U44913 (N_44913,N_33313,N_32412);
and U44914 (N_44914,N_35372,N_30152);
nand U44915 (N_44915,N_36190,N_32152);
and U44916 (N_44916,N_31969,N_34832);
nand U44917 (N_44917,N_36922,N_39178);
nor U44918 (N_44918,N_38272,N_39987);
nor U44919 (N_44919,N_31234,N_33010);
nor U44920 (N_44920,N_34641,N_33900);
nor U44921 (N_44921,N_35357,N_30432);
nand U44922 (N_44922,N_37467,N_37763);
and U44923 (N_44923,N_35132,N_38836);
nor U44924 (N_44924,N_36020,N_37347);
or U44925 (N_44925,N_30022,N_36964);
and U44926 (N_44926,N_39124,N_38477);
nand U44927 (N_44927,N_34689,N_34876);
and U44928 (N_44928,N_36139,N_38919);
nand U44929 (N_44929,N_31758,N_31962);
and U44930 (N_44930,N_30438,N_32244);
or U44931 (N_44931,N_34407,N_39956);
or U44932 (N_44932,N_35830,N_32467);
xor U44933 (N_44933,N_35484,N_33483);
and U44934 (N_44934,N_30169,N_35077);
nand U44935 (N_44935,N_38399,N_39361);
and U44936 (N_44936,N_39951,N_37511);
and U44937 (N_44937,N_34187,N_34140);
xor U44938 (N_44938,N_32911,N_32048);
or U44939 (N_44939,N_34548,N_30949);
xor U44940 (N_44940,N_37416,N_36690);
nor U44941 (N_44941,N_37386,N_30606);
and U44942 (N_44942,N_38802,N_35931);
and U44943 (N_44943,N_30377,N_37102);
or U44944 (N_44944,N_39749,N_38961);
or U44945 (N_44945,N_36583,N_38436);
nor U44946 (N_44946,N_33675,N_32313);
and U44947 (N_44947,N_35209,N_34182);
or U44948 (N_44948,N_38767,N_31568);
and U44949 (N_44949,N_31830,N_30616);
xnor U44950 (N_44950,N_37647,N_36270);
or U44951 (N_44951,N_30365,N_38003);
nand U44952 (N_44952,N_33334,N_34859);
or U44953 (N_44953,N_35697,N_33735);
nor U44954 (N_44954,N_31291,N_35112);
nor U44955 (N_44955,N_38992,N_37077);
or U44956 (N_44956,N_31372,N_30932);
nor U44957 (N_44957,N_38610,N_31565);
or U44958 (N_44958,N_37820,N_34371);
nand U44959 (N_44959,N_34892,N_33695);
or U44960 (N_44960,N_35566,N_34246);
nor U44961 (N_44961,N_31268,N_33939);
nor U44962 (N_44962,N_32707,N_31826);
and U44963 (N_44963,N_36935,N_35760);
xnor U44964 (N_44964,N_36314,N_38368);
xor U44965 (N_44965,N_36094,N_32982);
nor U44966 (N_44966,N_35886,N_31605);
nor U44967 (N_44967,N_38035,N_39470);
nor U44968 (N_44968,N_35029,N_38055);
and U44969 (N_44969,N_32603,N_38481);
xnor U44970 (N_44970,N_38646,N_31417);
nor U44971 (N_44971,N_32886,N_30412);
or U44972 (N_44972,N_33057,N_32865);
and U44973 (N_44973,N_39910,N_31608);
nand U44974 (N_44974,N_38985,N_33799);
nand U44975 (N_44975,N_37127,N_39532);
nand U44976 (N_44976,N_30227,N_36056);
or U44977 (N_44977,N_32866,N_30728);
nor U44978 (N_44978,N_31409,N_32688);
nor U44979 (N_44979,N_36958,N_36936);
and U44980 (N_44980,N_34556,N_37645);
nand U44981 (N_44981,N_32279,N_37336);
nor U44982 (N_44982,N_30219,N_32915);
nand U44983 (N_44983,N_35748,N_32287);
xnor U44984 (N_44984,N_38605,N_35020);
or U44985 (N_44985,N_35011,N_38166);
and U44986 (N_44986,N_38389,N_38728);
or U44987 (N_44987,N_37258,N_33933);
nand U44988 (N_44988,N_30649,N_35731);
nand U44989 (N_44989,N_38636,N_32415);
and U44990 (N_44990,N_36315,N_36419);
and U44991 (N_44991,N_38091,N_30183);
or U44992 (N_44992,N_36495,N_37555);
and U44993 (N_44993,N_30693,N_36699);
nor U44994 (N_44994,N_39884,N_35108);
or U44995 (N_44995,N_37499,N_34840);
nor U44996 (N_44996,N_37133,N_32569);
or U44997 (N_44997,N_36402,N_39826);
xor U44998 (N_44998,N_37901,N_33637);
and U44999 (N_44999,N_39310,N_38871);
nor U45000 (N_45000,N_39346,N_35043);
xor U45001 (N_45001,N_30460,N_30261);
or U45002 (N_45002,N_30687,N_32448);
and U45003 (N_45003,N_39549,N_35531);
and U45004 (N_45004,N_33525,N_37886);
or U45005 (N_45005,N_35027,N_39027);
and U45006 (N_45006,N_31130,N_39046);
xor U45007 (N_45007,N_31483,N_32945);
and U45008 (N_45008,N_33316,N_37248);
or U45009 (N_45009,N_38714,N_35594);
xor U45010 (N_45010,N_39058,N_34352);
nand U45011 (N_45011,N_33381,N_34785);
xnor U45012 (N_45012,N_37993,N_38704);
and U45013 (N_45013,N_33568,N_33219);
xor U45014 (N_45014,N_30329,N_39393);
or U45015 (N_45015,N_33335,N_31056);
nor U45016 (N_45016,N_33058,N_39650);
nand U45017 (N_45017,N_32867,N_39681);
xnor U45018 (N_45018,N_32481,N_37756);
nand U45019 (N_45019,N_39146,N_34699);
and U45020 (N_45020,N_32529,N_30902);
nand U45021 (N_45021,N_31075,N_31190);
nand U45022 (N_45022,N_36348,N_37480);
or U45023 (N_45023,N_33977,N_35574);
xnor U45024 (N_45024,N_39542,N_39727);
or U45025 (N_45025,N_31044,N_34032);
nand U45026 (N_45026,N_35805,N_35157);
or U45027 (N_45027,N_33445,N_36334);
nand U45028 (N_45028,N_30269,N_31525);
nand U45029 (N_45029,N_37894,N_34951);
nand U45030 (N_45030,N_36010,N_33693);
or U45031 (N_45031,N_39521,N_39632);
and U45032 (N_45032,N_36612,N_31877);
xnor U45033 (N_45033,N_32941,N_30418);
or U45034 (N_45034,N_38344,N_33884);
nor U45035 (N_45035,N_39740,N_36036);
nor U45036 (N_45036,N_39609,N_33985);
nor U45037 (N_45037,N_32522,N_33096);
xnor U45038 (N_45038,N_38782,N_37978);
nor U45039 (N_45039,N_32126,N_39437);
or U45040 (N_45040,N_39388,N_38217);
xnor U45041 (N_45041,N_37415,N_35059);
nor U45042 (N_45042,N_32999,N_37444);
nor U45043 (N_45043,N_32455,N_37938);
and U45044 (N_45044,N_32098,N_31097);
and U45045 (N_45045,N_37153,N_31076);
nor U45046 (N_45046,N_37702,N_39886);
nand U45047 (N_45047,N_34073,N_31968);
nand U45048 (N_45048,N_33004,N_39526);
nand U45049 (N_45049,N_31559,N_31415);
and U45050 (N_45050,N_39198,N_37790);
nand U45051 (N_45051,N_38860,N_36484);
nand U45052 (N_45052,N_35793,N_37674);
nand U45053 (N_45053,N_39516,N_30648);
nand U45054 (N_45054,N_39294,N_32592);
xor U45055 (N_45055,N_38336,N_35247);
and U45056 (N_45056,N_39259,N_31904);
or U45057 (N_45057,N_36437,N_38528);
or U45058 (N_45058,N_38087,N_35939);
nand U45059 (N_45059,N_39249,N_33121);
nand U45060 (N_45060,N_32690,N_32939);
xor U45061 (N_45061,N_39955,N_35622);
and U45062 (N_45062,N_37232,N_38228);
and U45063 (N_45063,N_37914,N_36288);
nor U45064 (N_45064,N_35575,N_38465);
or U45065 (N_45065,N_35905,N_36373);
nor U45066 (N_45066,N_35890,N_37055);
nor U45067 (N_45067,N_30430,N_36332);
and U45068 (N_45068,N_36615,N_31363);
nand U45069 (N_45069,N_32640,N_31504);
nand U45070 (N_45070,N_31582,N_31474);
nor U45071 (N_45071,N_32940,N_34247);
nor U45072 (N_45072,N_33441,N_38207);
and U45073 (N_45073,N_34240,N_39998);
and U45074 (N_45074,N_37301,N_33616);
or U45075 (N_45075,N_37794,N_39797);
and U45076 (N_45076,N_30622,N_33144);
and U45077 (N_45077,N_37825,N_32048);
and U45078 (N_45078,N_33827,N_36844);
or U45079 (N_45079,N_33383,N_34938);
or U45080 (N_45080,N_38130,N_38177);
and U45081 (N_45081,N_31889,N_37229);
or U45082 (N_45082,N_34736,N_30572);
and U45083 (N_45083,N_38909,N_37287);
and U45084 (N_45084,N_35393,N_35695);
and U45085 (N_45085,N_39029,N_35351);
and U45086 (N_45086,N_33992,N_39460);
or U45087 (N_45087,N_38997,N_36283);
and U45088 (N_45088,N_30681,N_30223);
nand U45089 (N_45089,N_38940,N_31033);
nor U45090 (N_45090,N_35733,N_32973);
or U45091 (N_45091,N_38059,N_36549);
nand U45092 (N_45092,N_34117,N_32111);
nand U45093 (N_45093,N_35235,N_33373);
or U45094 (N_45094,N_35635,N_36384);
or U45095 (N_45095,N_37919,N_33978);
or U45096 (N_45096,N_33104,N_35552);
nor U45097 (N_45097,N_30464,N_32256);
nand U45098 (N_45098,N_33032,N_32516);
nand U45099 (N_45099,N_36170,N_38001);
and U45100 (N_45100,N_38400,N_32671);
and U45101 (N_45101,N_30723,N_31933);
nand U45102 (N_45102,N_35090,N_34947);
nand U45103 (N_45103,N_33708,N_38651);
xnor U45104 (N_45104,N_39591,N_33102);
and U45105 (N_45105,N_31160,N_37486);
nor U45106 (N_45106,N_37680,N_31542);
xor U45107 (N_45107,N_34033,N_34414);
nor U45108 (N_45108,N_32234,N_32473);
or U45109 (N_45109,N_36610,N_37932);
nand U45110 (N_45110,N_33467,N_32735);
and U45111 (N_45111,N_38684,N_39268);
nor U45112 (N_45112,N_31764,N_38531);
or U45113 (N_45113,N_38347,N_36176);
and U45114 (N_45114,N_33225,N_33389);
nand U45115 (N_45115,N_35748,N_30732);
nor U45116 (N_45116,N_34905,N_37137);
or U45117 (N_45117,N_38774,N_36100);
nor U45118 (N_45118,N_38381,N_33081);
nor U45119 (N_45119,N_37046,N_36644);
nand U45120 (N_45120,N_33898,N_33395);
xnor U45121 (N_45121,N_35349,N_35499);
nand U45122 (N_45122,N_32898,N_38784);
and U45123 (N_45123,N_33748,N_35249);
and U45124 (N_45124,N_38613,N_31535);
or U45125 (N_45125,N_35681,N_31028);
nand U45126 (N_45126,N_34569,N_33990);
and U45127 (N_45127,N_39287,N_38479);
nand U45128 (N_45128,N_37374,N_35660);
and U45129 (N_45129,N_36264,N_39957);
xnor U45130 (N_45130,N_30853,N_36067);
nor U45131 (N_45131,N_36253,N_35482);
and U45132 (N_45132,N_38349,N_39464);
nor U45133 (N_45133,N_37542,N_31341);
nand U45134 (N_45134,N_34742,N_31435);
and U45135 (N_45135,N_34663,N_32175);
and U45136 (N_45136,N_33659,N_38414);
nor U45137 (N_45137,N_38373,N_34281);
nand U45138 (N_45138,N_34204,N_37687);
and U45139 (N_45139,N_37893,N_35759);
or U45140 (N_45140,N_38402,N_31469);
nor U45141 (N_45141,N_36463,N_36066);
nand U45142 (N_45142,N_33134,N_32968);
and U45143 (N_45143,N_36584,N_30184);
or U45144 (N_45144,N_32754,N_30188);
and U45145 (N_45145,N_39789,N_34282);
and U45146 (N_45146,N_37383,N_37761);
and U45147 (N_45147,N_36597,N_39113);
and U45148 (N_45148,N_30218,N_34188);
nand U45149 (N_45149,N_38221,N_31577);
or U45150 (N_45150,N_36768,N_39282);
nand U45151 (N_45151,N_37462,N_38969);
nor U45152 (N_45152,N_33796,N_34061);
and U45153 (N_45153,N_39685,N_33793);
or U45154 (N_45154,N_39494,N_32908);
and U45155 (N_45155,N_35033,N_37554);
nand U45156 (N_45156,N_33498,N_38875);
nand U45157 (N_45157,N_37465,N_38173);
nor U45158 (N_45158,N_30238,N_36791);
or U45159 (N_45159,N_33554,N_32652);
nor U45160 (N_45160,N_35193,N_39683);
or U45161 (N_45161,N_31155,N_38858);
nor U45162 (N_45162,N_38287,N_32100);
nand U45163 (N_45163,N_39628,N_39513);
nand U45164 (N_45164,N_37236,N_37233);
and U45165 (N_45165,N_34111,N_36203);
nand U45166 (N_45166,N_35576,N_36823);
or U45167 (N_45167,N_31594,N_36394);
xor U45168 (N_45168,N_34444,N_33730);
nand U45169 (N_45169,N_35194,N_38367);
nor U45170 (N_45170,N_34378,N_35166);
or U45171 (N_45171,N_36780,N_33590);
xnor U45172 (N_45172,N_31347,N_32868);
and U45173 (N_45173,N_35186,N_36251);
xnor U45174 (N_45174,N_33558,N_36681);
or U45175 (N_45175,N_36210,N_32754);
nand U45176 (N_45176,N_31218,N_32481);
and U45177 (N_45177,N_36437,N_34601);
or U45178 (N_45178,N_37414,N_35385);
nand U45179 (N_45179,N_30009,N_37633);
nor U45180 (N_45180,N_31139,N_30345);
and U45181 (N_45181,N_34968,N_35463);
and U45182 (N_45182,N_33133,N_33397);
or U45183 (N_45183,N_34200,N_31093);
nor U45184 (N_45184,N_35621,N_35867);
nand U45185 (N_45185,N_37022,N_34606);
nor U45186 (N_45186,N_31563,N_32343);
nor U45187 (N_45187,N_32321,N_30475);
nand U45188 (N_45188,N_39735,N_36652);
and U45189 (N_45189,N_35458,N_36434);
xor U45190 (N_45190,N_37474,N_30252);
or U45191 (N_45191,N_33013,N_37985);
and U45192 (N_45192,N_37678,N_30949);
nor U45193 (N_45193,N_30379,N_39416);
nor U45194 (N_45194,N_32063,N_31168);
and U45195 (N_45195,N_35458,N_31209);
or U45196 (N_45196,N_31499,N_32884);
and U45197 (N_45197,N_35162,N_34206);
and U45198 (N_45198,N_39935,N_30350);
or U45199 (N_45199,N_36487,N_30586);
nand U45200 (N_45200,N_35106,N_30574);
nor U45201 (N_45201,N_38264,N_32328);
xor U45202 (N_45202,N_31069,N_36877);
xnor U45203 (N_45203,N_39155,N_30677);
and U45204 (N_45204,N_33656,N_32566);
nor U45205 (N_45205,N_34505,N_35186);
nor U45206 (N_45206,N_35186,N_30307);
nand U45207 (N_45207,N_31756,N_36338);
nor U45208 (N_45208,N_36311,N_31188);
and U45209 (N_45209,N_36612,N_32478);
and U45210 (N_45210,N_37180,N_30631);
nand U45211 (N_45211,N_38454,N_38321);
or U45212 (N_45212,N_39711,N_35267);
nor U45213 (N_45213,N_36752,N_35973);
nand U45214 (N_45214,N_34131,N_33731);
nand U45215 (N_45215,N_36727,N_34363);
or U45216 (N_45216,N_33577,N_30660);
nor U45217 (N_45217,N_35236,N_32245);
and U45218 (N_45218,N_38606,N_37826);
nor U45219 (N_45219,N_34841,N_33809);
nand U45220 (N_45220,N_31484,N_33221);
nor U45221 (N_45221,N_35684,N_35143);
nand U45222 (N_45222,N_38095,N_35039);
nand U45223 (N_45223,N_37421,N_33854);
and U45224 (N_45224,N_30927,N_36069);
nor U45225 (N_45225,N_35301,N_32574);
or U45226 (N_45226,N_39032,N_35609);
and U45227 (N_45227,N_33416,N_39743);
and U45228 (N_45228,N_38466,N_34560);
and U45229 (N_45229,N_39897,N_35090);
nor U45230 (N_45230,N_37667,N_38682);
nor U45231 (N_45231,N_32659,N_38623);
nand U45232 (N_45232,N_34475,N_38551);
nand U45233 (N_45233,N_38088,N_36350);
or U45234 (N_45234,N_33412,N_30599);
or U45235 (N_45235,N_38099,N_37784);
nand U45236 (N_45236,N_36009,N_34458);
or U45237 (N_45237,N_33980,N_32997);
xor U45238 (N_45238,N_30845,N_35689);
nand U45239 (N_45239,N_31385,N_32247);
or U45240 (N_45240,N_36216,N_34787);
nor U45241 (N_45241,N_38835,N_37309);
or U45242 (N_45242,N_32592,N_30467);
or U45243 (N_45243,N_33869,N_39716);
nand U45244 (N_45244,N_35323,N_37392);
nor U45245 (N_45245,N_37975,N_39946);
and U45246 (N_45246,N_34115,N_33061);
or U45247 (N_45247,N_33501,N_32715);
nor U45248 (N_45248,N_34438,N_33857);
or U45249 (N_45249,N_37979,N_38706);
and U45250 (N_45250,N_33900,N_32668);
nand U45251 (N_45251,N_33545,N_31763);
nand U45252 (N_45252,N_32895,N_34896);
xor U45253 (N_45253,N_39057,N_33549);
xnor U45254 (N_45254,N_36108,N_37405);
and U45255 (N_45255,N_37778,N_33512);
nand U45256 (N_45256,N_31141,N_37876);
and U45257 (N_45257,N_32868,N_37411);
or U45258 (N_45258,N_35333,N_31587);
xor U45259 (N_45259,N_37628,N_39514);
nand U45260 (N_45260,N_38521,N_33065);
or U45261 (N_45261,N_31255,N_31228);
and U45262 (N_45262,N_34965,N_34030);
or U45263 (N_45263,N_35540,N_32413);
nand U45264 (N_45264,N_38875,N_34418);
and U45265 (N_45265,N_37401,N_35628);
nand U45266 (N_45266,N_39577,N_32974);
nand U45267 (N_45267,N_35513,N_33174);
nor U45268 (N_45268,N_35172,N_36558);
nand U45269 (N_45269,N_35414,N_36560);
or U45270 (N_45270,N_36260,N_38804);
and U45271 (N_45271,N_34448,N_39692);
nand U45272 (N_45272,N_35190,N_30639);
nor U45273 (N_45273,N_37172,N_38150);
or U45274 (N_45274,N_36454,N_34548);
nand U45275 (N_45275,N_30883,N_37123);
nor U45276 (N_45276,N_32065,N_32426);
and U45277 (N_45277,N_30392,N_34072);
nor U45278 (N_45278,N_31641,N_31073);
nor U45279 (N_45279,N_38633,N_38775);
xnor U45280 (N_45280,N_35923,N_38077);
nand U45281 (N_45281,N_39509,N_35846);
or U45282 (N_45282,N_39890,N_34813);
nand U45283 (N_45283,N_37462,N_32462);
or U45284 (N_45284,N_36921,N_37550);
or U45285 (N_45285,N_35941,N_39302);
and U45286 (N_45286,N_38875,N_32179);
nor U45287 (N_45287,N_39544,N_33562);
nand U45288 (N_45288,N_34774,N_38387);
nor U45289 (N_45289,N_30252,N_39987);
or U45290 (N_45290,N_38564,N_37674);
and U45291 (N_45291,N_33688,N_36050);
nand U45292 (N_45292,N_30787,N_34663);
and U45293 (N_45293,N_38372,N_30397);
or U45294 (N_45294,N_36764,N_37494);
or U45295 (N_45295,N_39540,N_39767);
or U45296 (N_45296,N_37077,N_37052);
or U45297 (N_45297,N_34065,N_34726);
nor U45298 (N_45298,N_33624,N_33017);
nand U45299 (N_45299,N_36275,N_33750);
xor U45300 (N_45300,N_31640,N_34783);
and U45301 (N_45301,N_38650,N_39129);
nand U45302 (N_45302,N_31592,N_35832);
and U45303 (N_45303,N_37377,N_31090);
and U45304 (N_45304,N_32661,N_33099);
nor U45305 (N_45305,N_36110,N_35358);
or U45306 (N_45306,N_32411,N_34815);
or U45307 (N_45307,N_36910,N_39769);
and U45308 (N_45308,N_32263,N_36573);
or U45309 (N_45309,N_33191,N_38416);
nand U45310 (N_45310,N_30052,N_37972);
nor U45311 (N_45311,N_35468,N_31418);
and U45312 (N_45312,N_32619,N_33183);
or U45313 (N_45313,N_35373,N_33987);
nand U45314 (N_45314,N_35150,N_36848);
or U45315 (N_45315,N_37839,N_39534);
nand U45316 (N_45316,N_34448,N_30116);
and U45317 (N_45317,N_30859,N_39433);
nand U45318 (N_45318,N_35830,N_32401);
nand U45319 (N_45319,N_34250,N_30835);
nand U45320 (N_45320,N_35805,N_39778);
or U45321 (N_45321,N_30303,N_33131);
and U45322 (N_45322,N_37056,N_37276);
or U45323 (N_45323,N_39254,N_32576);
and U45324 (N_45324,N_36034,N_36199);
xnor U45325 (N_45325,N_32243,N_37554);
nand U45326 (N_45326,N_32638,N_34099);
and U45327 (N_45327,N_32719,N_34088);
and U45328 (N_45328,N_38100,N_33016);
xor U45329 (N_45329,N_37050,N_35957);
nor U45330 (N_45330,N_31092,N_35621);
nand U45331 (N_45331,N_34618,N_36136);
xnor U45332 (N_45332,N_37749,N_36507);
or U45333 (N_45333,N_30325,N_34565);
and U45334 (N_45334,N_31565,N_36109);
nor U45335 (N_45335,N_31874,N_34032);
nand U45336 (N_45336,N_37581,N_31436);
or U45337 (N_45337,N_32866,N_30944);
nand U45338 (N_45338,N_39957,N_32034);
nand U45339 (N_45339,N_37162,N_30444);
nand U45340 (N_45340,N_39248,N_33845);
and U45341 (N_45341,N_31015,N_38547);
and U45342 (N_45342,N_35967,N_36540);
and U45343 (N_45343,N_32644,N_34205);
or U45344 (N_45344,N_38089,N_39666);
nand U45345 (N_45345,N_39102,N_38269);
xor U45346 (N_45346,N_36915,N_37345);
and U45347 (N_45347,N_35098,N_35418);
and U45348 (N_45348,N_34718,N_37859);
xnor U45349 (N_45349,N_34295,N_38561);
nand U45350 (N_45350,N_33607,N_30760);
nor U45351 (N_45351,N_33977,N_32959);
or U45352 (N_45352,N_39655,N_38089);
or U45353 (N_45353,N_36743,N_37524);
or U45354 (N_45354,N_35655,N_33402);
nand U45355 (N_45355,N_36192,N_32303);
or U45356 (N_45356,N_31819,N_37099);
nand U45357 (N_45357,N_35889,N_31144);
nand U45358 (N_45358,N_38806,N_39537);
and U45359 (N_45359,N_32126,N_31296);
nor U45360 (N_45360,N_36811,N_35234);
or U45361 (N_45361,N_35466,N_31312);
or U45362 (N_45362,N_35554,N_33877);
and U45363 (N_45363,N_37667,N_35888);
xor U45364 (N_45364,N_32022,N_36811);
nand U45365 (N_45365,N_35731,N_39356);
nand U45366 (N_45366,N_30910,N_30592);
nand U45367 (N_45367,N_30468,N_39728);
nor U45368 (N_45368,N_35544,N_35758);
nor U45369 (N_45369,N_32777,N_33843);
and U45370 (N_45370,N_39422,N_37354);
xnor U45371 (N_45371,N_38398,N_32512);
nor U45372 (N_45372,N_30789,N_30106);
or U45373 (N_45373,N_31118,N_37431);
or U45374 (N_45374,N_38714,N_39724);
nand U45375 (N_45375,N_31370,N_39469);
or U45376 (N_45376,N_31796,N_38970);
and U45377 (N_45377,N_38956,N_31331);
or U45378 (N_45378,N_38925,N_32003);
xor U45379 (N_45379,N_39018,N_38553);
nand U45380 (N_45380,N_31431,N_36782);
xor U45381 (N_45381,N_37004,N_33876);
nand U45382 (N_45382,N_38014,N_34780);
nor U45383 (N_45383,N_35438,N_32484);
and U45384 (N_45384,N_32947,N_37944);
nand U45385 (N_45385,N_34579,N_34047);
nand U45386 (N_45386,N_36164,N_36025);
or U45387 (N_45387,N_39190,N_38436);
or U45388 (N_45388,N_32558,N_31497);
nand U45389 (N_45389,N_37623,N_30596);
nor U45390 (N_45390,N_34602,N_34016);
nand U45391 (N_45391,N_39319,N_34667);
or U45392 (N_45392,N_35246,N_36891);
xnor U45393 (N_45393,N_32801,N_36211);
nor U45394 (N_45394,N_39736,N_33513);
nor U45395 (N_45395,N_31307,N_33976);
nor U45396 (N_45396,N_33751,N_31176);
and U45397 (N_45397,N_34370,N_30220);
nand U45398 (N_45398,N_33604,N_34443);
and U45399 (N_45399,N_38026,N_34476);
nor U45400 (N_45400,N_39079,N_37140);
and U45401 (N_45401,N_33755,N_33460);
or U45402 (N_45402,N_30097,N_39676);
nor U45403 (N_45403,N_36352,N_36928);
xnor U45404 (N_45404,N_38984,N_36601);
or U45405 (N_45405,N_30657,N_31131);
nand U45406 (N_45406,N_38778,N_38391);
and U45407 (N_45407,N_36873,N_33570);
nor U45408 (N_45408,N_34745,N_37577);
nor U45409 (N_45409,N_33301,N_36071);
and U45410 (N_45410,N_33631,N_31890);
and U45411 (N_45411,N_39876,N_35702);
or U45412 (N_45412,N_37109,N_34507);
and U45413 (N_45413,N_39308,N_37711);
or U45414 (N_45414,N_35213,N_39415);
and U45415 (N_45415,N_32037,N_34435);
or U45416 (N_45416,N_35670,N_34949);
nand U45417 (N_45417,N_38733,N_33233);
or U45418 (N_45418,N_36547,N_35513);
and U45419 (N_45419,N_38311,N_30952);
and U45420 (N_45420,N_35069,N_32310);
nand U45421 (N_45421,N_36785,N_38853);
and U45422 (N_45422,N_38628,N_38348);
and U45423 (N_45423,N_34247,N_35152);
nand U45424 (N_45424,N_37322,N_39125);
and U45425 (N_45425,N_37384,N_35359);
or U45426 (N_45426,N_31215,N_30434);
nand U45427 (N_45427,N_33708,N_39464);
and U45428 (N_45428,N_33731,N_38210);
xnor U45429 (N_45429,N_30227,N_39798);
and U45430 (N_45430,N_39914,N_38629);
nand U45431 (N_45431,N_30668,N_30126);
and U45432 (N_45432,N_36501,N_38888);
nand U45433 (N_45433,N_35260,N_38406);
xnor U45434 (N_45434,N_34199,N_36600);
or U45435 (N_45435,N_39817,N_37376);
nand U45436 (N_45436,N_38887,N_35190);
nand U45437 (N_45437,N_33463,N_39068);
xnor U45438 (N_45438,N_30484,N_32791);
nor U45439 (N_45439,N_35492,N_37704);
and U45440 (N_45440,N_32990,N_36179);
or U45441 (N_45441,N_39314,N_35680);
or U45442 (N_45442,N_34420,N_34177);
nand U45443 (N_45443,N_37223,N_39448);
nand U45444 (N_45444,N_33582,N_37193);
nor U45445 (N_45445,N_34470,N_31045);
nor U45446 (N_45446,N_30874,N_34616);
and U45447 (N_45447,N_36787,N_33631);
and U45448 (N_45448,N_37222,N_34163);
nand U45449 (N_45449,N_35385,N_33374);
xor U45450 (N_45450,N_35463,N_37295);
or U45451 (N_45451,N_35474,N_35493);
nand U45452 (N_45452,N_32382,N_38455);
nand U45453 (N_45453,N_34486,N_36212);
nand U45454 (N_45454,N_37209,N_30789);
nand U45455 (N_45455,N_38681,N_34834);
nand U45456 (N_45456,N_33832,N_34999);
or U45457 (N_45457,N_30471,N_33116);
nand U45458 (N_45458,N_33018,N_36238);
nor U45459 (N_45459,N_37797,N_36452);
nor U45460 (N_45460,N_39624,N_38471);
xor U45461 (N_45461,N_36748,N_37613);
and U45462 (N_45462,N_39216,N_31182);
or U45463 (N_45463,N_31854,N_35867);
nand U45464 (N_45464,N_36702,N_37085);
and U45465 (N_45465,N_38612,N_38091);
xnor U45466 (N_45466,N_34314,N_30522);
nand U45467 (N_45467,N_38091,N_35908);
or U45468 (N_45468,N_33815,N_35299);
or U45469 (N_45469,N_34335,N_37226);
nor U45470 (N_45470,N_34222,N_34252);
or U45471 (N_45471,N_35420,N_39741);
or U45472 (N_45472,N_31147,N_31119);
and U45473 (N_45473,N_33899,N_32932);
nor U45474 (N_45474,N_32212,N_35265);
or U45475 (N_45475,N_33989,N_36740);
nand U45476 (N_45476,N_35368,N_35445);
or U45477 (N_45477,N_39933,N_30351);
or U45478 (N_45478,N_34563,N_37324);
nor U45479 (N_45479,N_39015,N_34526);
nand U45480 (N_45480,N_30784,N_38795);
nor U45481 (N_45481,N_39992,N_33524);
or U45482 (N_45482,N_33083,N_30527);
or U45483 (N_45483,N_35200,N_37820);
nand U45484 (N_45484,N_30202,N_31234);
nor U45485 (N_45485,N_30269,N_35262);
and U45486 (N_45486,N_35488,N_32266);
nor U45487 (N_45487,N_39139,N_36702);
nand U45488 (N_45488,N_31574,N_39919);
nor U45489 (N_45489,N_33279,N_32378);
nand U45490 (N_45490,N_35925,N_34955);
xnor U45491 (N_45491,N_37476,N_30019);
nand U45492 (N_45492,N_36896,N_33338);
and U45493 (N_45493,N_39144,N_30389);
nand U45494 (N_45494,N_33226,N_38017);
or U45495 (N_45495,N_38550,N_32131);
nor U45496 (N_45496,N_34812,N_37724);
nor U45497 (N_45497,N_30500,N_31709);
and U45498 (N_45498,N_34929,N_37125);
xor U45499 (N_45499,N_31892,N_31998);
nand U45500 (N_45500,N_39437,N_39830);
and U45501 (N_45501,N_38946,N_30760);
xnor U45502 (N_45502,N_34367,N_38828);
and U45503 (N_45503,N_33156,N_35629);
and U45504 (N_45504,N_33337,N_33878);
and U45505 (N_45505,N_31342,N_31889);
nand U45506 (N_45506,N_32200,N_32797);
and U45507 (N_45507,N_32320,N_32681);
nor U45508 (N_45508,N_36229,N_35183);
nand U45509 (N_45509,N_33121,N_37218);
and U45510 (N_45510,N_39221,N_37730);
and U45511 (N_45511,N_33447,N_39204);
or U45512 (N_45512,N_33376,N_38098);
or U45513 (N_45513,N_33872,N_31786);
nand U45514 (N_45514,N_31230,N_33997);
nor U45515 (N_45515,N_34251,N_39933);
and U45516 (N_45516,N_30657,N_31852);
or U45517 (N_45517,N_37858,N_32144);
or U45518 (N_45518,N_30561,N_38606);
or U45519 (N_45519,N_39078,N_31565);
nor U45520 (N_45520,N_33043,N_30755);
and U45521 (N_45521,N_32570,N_38192);
or U45522 (N_45522,N_36917,N_35428);
and U45523 (N_45523,N_38949,N_35922);
nor U45524 (N_45524,N_32662,N_37330);
or U45525 (N_45525,N_31206,N_36578);
nand U45526 (N_45526,N_31077,N_34237);
nand U45527 (N_45527,N_37615,N_32812);
nor U45528 (N_45528,N_38428,N_35163);
xor U45529 (N_45529,N_37463,N_30566);
nor U45530 (N_45530,N_37880,N_35997);
nor U45531 (N_45531,N_32111,N_31146);
nor U45532 (N_45532,N_37954,N_33965);
nor U45533 (N_45533,N_34101,N_34295);
and U45534 (N_45534,N_34450,N_34321);
or U45535 (N_45535,N_31011,N_35730);
or U45536 (N_45536,N_32600,N_32539);
xnor U45537 (N_45537,N_37612,N_37709);
nand U45538 (N_45538,N_32268,N_39140);
and U45539 (N_45539,N_36961,N_37097);
nand U45540 (N_45540,N_37033,N_35379);
nor U45541 (N_45541,N_33785,N_39741);
nand U45542 (N_45542,N_35430,N_33846);
or U45543 (N_45543,N_34787,N_39374);
nand U45544 (N_45544,N_35179,N_34341);
xnor U45545 (N_45545,N_37274,N_37400);
nand U45546 (N_45546,N_37485,N_35646);
or U45547 (N_45547,N_34903,N_33827);
nor U45548 (N_45548,N_33186,N_32810);
and U45549 (N_45549,N_32746,N_39086);
and U45550 (N_45550,N_37713,N_31815);
nor U45551 (N_45551,N_36969,N_32806);
xor U45552 (N_45552,N_37957,N_36311);
nand U45553 (N_45553,N_37820,N_33219);
nor U45554 (N_45554,N_32835,N_34384);
nand U45555 (N_45555,N_35696,N_39024);
or U45556 (N_45556,N_30241,N_34574);
nor U45557 (N_45557,N_31601,N_36597);
nor U45558 (N_45558,N_39902,N_37490);
nor U45559 (N_45559,N_32956,N_30183);
nor U45560 (N_45560,N_39592,N_33821);
nor U45561 (N_45561,N_31667,N_39876);
nor U45562 (N_45562,N_30609,N_34498);
nor U45563 (N_45563,N_34360,N_36256);
and U45564 (N_45564,N_37661,N_38685);
nor U45565 (N_45565,N_38348,N_39110);
and U45566 (N_45566,N_33407,N_33874);
or U45567 (N_45567,N_32714,N_37261);
or U45568 (N_45568,N_35339,N_34575);
or U45569 (N_45569,N_30910,N_36788);
or U45570 (N_45570,N_30146,N_32725);
nand U45571 (N_45571,N_39133,N_30652);
or U45572 (N_45572,N_31945,N_39477);
xnor U45573 (N_45573,N_36606,N_35209);
nand U45574 (N_45574,N_35952,N_34938);
or U45575 (N_45575,N_33698,N_31489);
and U45576 (N_45576,N_30880,N_31676);
nor U45577 (N_45577,N_37557,N_36183);
xnor U45578 (N_45578,N_30640,N_34231);
and U45579 (N_45579,N_34190,N_35998);
nand U45580 (N_45580,N_38843,N_35419);
nor U45581 (N_45581,N_38284,N_30627);
nor U45582 (N_45582,N_37878,N_39445);
xnor U45583 (N_45583,N_37180,N_36364);
nor U45584 (N_45584,N_33878,N_36300);
or U45585 (N_45585,N_35410,N_32150);
and U45586 (N_45586,N_39424,N_31517);
nand U45587 (N_45587,N_36892,N_30202);
and U45588 (N_45588,N_32208,N_35719);
or U45589 (N_45589,N_33663,N_39935);
or U45590 (N_45590,N_39322,N_30644);
nor U45591 (N_45591,N_38427,N_39514);
and U45592 (N_45592,N_30540,N_35547);
or U45593 (N_45593,N_34392,N_38737);
xnor U45594 (N_45594,N_38000,N_34289);
xnor U45595 (N_45595,N_33865,N_32640);
or U45596 (N_45596,N_36742,N_39319);
or U45597 (N_45597,N_39501,N_36475);
xnor U45598 (N_45598,N_38517,N_37703);
nand U45599 (N_45599,N_31100,N_37582);
nand U45600 (N_45600,N_32049,N_33884);
and U45601 (N_45601,N_30317,N_33635);
or U45602 (N_45602,N_37790,N_38328);
nor U45603 (N_45603,N_33682,N_31165);
or U45604 (N_45604,N_31750,N_37305);
and U45605 (N_45605,N_34119,N_32176);
or U45606 (N_45606,N_39890,N_39775);
xor U45607 (N_45607,N_39238,N_34140);
or U45608 (N_45608,N_35213,N_30113);
and U45609 (N_45609,N_37402,N_37153);
xor U45610 (N_45610,N_36206,N_31717);
nand U45611 (N_45611,N_36160,N_36012);
nand U45612 (N_45612,N_31357,N_34772);
xor U45613 (N_45613,N_37188,N_32716);
and U45614 (N_45614,N_34399,N_37049);
xor U45615 (N_45615,N_35552,N_36556);
nor U45616 (N_45616,N_39044,N_35029);
nor U45617 (N_45617,N_39535,N_36553);
and U45618 (N_45618,N_31007,N_36381);
xor U45619 (N_45619,N_33474,N_37503);
or U45620 (N_45620,N_37540,N_38300);
or U45621 (N_45621,N_39783,N_35613);
nor U45622 (N_45622,N_32072,N_32951);
nor U45623 (N_45623,N_34822,N_37525);
and U45624 (N_45624,N_30969,N_36649);
nand U45625 (N_45625,N_38405,N_38231);
or U45626 (N_45626,N_33102,N_38041);
or U45627 (N_45627,N_32456,N_31863);
or U45628 (N_45628,N_31235,N_33689);
and U45629 (N_45629,N_32854,N_30819);
or U45630 (N_45630,N_39053,N_35925);
and U45631 (N_45631,N_31983,N_35124);
nor U45632 (N_45632,N_33894,N_37576);
and U45633 (N_45633,N_32769,N_33466);
or U45634 (N_45634,N_31830,N_34834);
nor U45635 (N_45635,N_32586,N_32030);
or U45636 (N_45636,N_32091,N_39615);
or U45637 (N_45637,N_31169,N_36929);
nand U45638 (N_45638,N_30979,N_30392);
and U45639 (N_45639,N_39954,N_31848);
xor U45640 (N_45640,N_30073,N_32134);
and U45641 (N_45641,N_35479,N_36142);
and U45642 (N_45642,N_39831,N_35951);
xnor U45643 (N_45643,N_33190,N_37395);
or U45644 (N_45644,N_39281,N_32513);
xnor U45645 (N_45645,N_37319,N_31964);
xor U45646 (N_45646,N_33374,N_34444);
and U45647 (N_45647,N_34520,N_31236);
and U45648 (N_45648,N_33724,N_35953);
or U45649 (N_45649,N_34327,N_31476);
nor U45650 (N_45650,N_30243,N_34021);
and U45651 (N_45651,N_38793,N_33571);
nor U45652 (N_45652,N_35280,N_34928);
or U45653 (N_45653,N_35968,N_33602);
nor U45654 (N_45654,N_35962,N_30674);
nand U45655 (N_45655,N_39620,N_31133);
nor U45656 (N_45656,N_31707,N_39816);
and U45657 (N_45657,N_31225,N_31328);
or U45658 (N_45658,N_37720,N_31785);
and U45659 (N_45659,N_36708,N_38403);
nor U45660 (N_45660,N_36978,N_38553);
or U45661 (N_45661,N_31541,N_37920);
and U45662 (N_45662,N_32432,N_36385);
and U45663 (N_45663,N_37430,N_37534);
nor U45664 (N_45664,N_31887,N_34351);
or U45665 (N_45665,N_39084,N_34369);
or U45666 (N_45666,N_34985,N_37178);
and U45667 (N_45667,N_36006,N_35838);
and U45668 (N_45668,N_30895,N_35342);
and U45669 (N_45669,N_33544,N_34458);
nor U45670 (N_45670,N_30965,N_35482);
nor U45671 (N_45671,N_37100,N_31416);
nor U45672 (N_45672,N_31897,N_32142);
nand U45673 (N_45673,N_38694,N_35540);
nand U45674 (N_45674,N_30196,N_37807);
or U45675 (N_45675,N_36718,N_37403);
nand U45676 (N_45676,N_31725,N_35257);
nor U45677 (N_45677,N_33678,N_38611);
nor U45678 (N_45678,N_33961,N_32339);
nand U45679 (N_45679,N_35437,N_36908);
and U45680 (N_45680,N_32334,N_30227);
xor U45681 (N_45681,N_36565,N_32067);
or U45682 (N_45682,N_39977,N_30694);
nor U45683 (N_45683,N_37557,N_39849);
and U45684 (N_45684,N_34039,N_31875);
nor U45685 (N_45685,N_39158,N_36751);
or U45686 (N_45686,N_37081,N_33435);
nand U45687 (N_45687,N_39325,N_39794);
or U45688 (N_45688,N_33302,N_39105);
and U45689 (N_45689,N_35411,N_33741);
nand U45690 (N_45690,N_31575,N_30588);
and U45691 (N_45691,N_34084,N_39312);
or U45692 (N_45692,N_33618,N_39674);
nand U45693 (N_45693,N_39436,N_33429);
nand U45694 (N_45694,N_34420,N_36887);
nand U45695 (N_45695,N_31850,N_30587);
or U45696 (N_45696,N_35032,N_30783);
xor U45697 (N_45697,N_32233,N_36801);
or U45698 (N_45698,N_34390,N_39809);
nand U45699 (N_45699,N_36229,N_31723);
nor U45700 (N_45700,N_33475,N_39914);
and U45701 (N_45701,N_39411,N_39969);
or U45702 (N_45702,N_31488,N_36504);
and U45703 (N_45703,N_30576,N_30967);
and U45704 (N_45704,N_32764,N_35921);
xnor U45705 (N_45705,N_31118,N_35198);
or U45706 (N_45706,N_36792,N_35477);
and U45707 (N_45707,N_36208,N_33640);
and U45708 (N_45708,N_34370,N_39963);
and U45709 (N_45709,N_39500,N_32952);
xnor U45710 (N_45710,N_35509,N_32610);
nor U45711 (N_45711,N_36778,N_37225);
or U45712 (N_45712,N_30089,N_37609);
and U45713 (N_45713,N_39995,N_35616);
and U45714 (N_45714,N_39888,N_39291);
nor U45715 (N_45715,N_39343,N_38812);
or U45716 (N_45716,N_36364,N_31201);
nand U45717 (N_45717,N_31668,N_32451);
nor U45718 (N_45718,N_38687,N_35808);
xor U45719 (N_45719,N_39800,N_39356);
nand U45720 (N_45720,N_39292,N_32040);
nor U45721 (N_45721,N_39979,N_36492);
nand U45722 (N_45722,N_35214,N_31496);
nor U45723 (N_45723,N_38699,N_37357);
nor U45724 (N_45724,N_30366,N_33895);
nor U45725 (N_45725,N_34952,N_30144);
xor U45726 (N_45726,N_36184,N_31279);
nand U45727 (N_45727,N_33368,N_38121);
nand U45728 (N_45728,N_37463,N_32448);
nand U45729 (N_45729,N_31931,N_33363);
nor U45730 (N_45730,N_33905,N_35302);
nor U45731 (N_45731,N_35005,N_32170);
xnor U45732 (N_45732,N_33085,N_39544);
nand U45733 (N_45733,N_34315,N_32445);
and U45734 (N_45734,N_39171,N_39462);
and U45735 (N_45735,N_38006,N_36270);
or U45736 (N_45736,N_38690,N_38777);
nor U45737 (N_45737,N_30488,N_34470);
xor U45738 (N_45738,N_30383,N_36964);
and U45739 (N_45739,N_39276,N_32616);
and U45740 (N_45740,N_30807,N_30712);
or U45741 (N_45741,N_33663,N_35001);
nand U45742 (N_45742,N_33320,N_33755);
nand U45743 (N_45743,N_36449,N_30581);
or U45744 (N_45744,N_37099,N_31097);
and U45745 (N_45745,N_33639,N_38124);
nor U45746 (N_45746,N_31485,N_33722);
or U45747 (N_45747,N_32631,N_31060);
and U45748 (N_45748,N_37181,N_37862);
and U45749 (N_45749,N_31256,N_34192);
nand U45750 (N_45750,N_30822,N_37945);
or U45751 (N_45751,N_37410,N_36585);
and U45752 (N_45752,N_37209,N_31838);
nor U45753 (N_45753,N_30984,N_39613);
and U45754 (N_45754,N_38066,N_37695);
nor U45755 (N_45755,N_33525,N_35610);
nor U45756 (N_45756,N_35337,N_30814);
xnor U45757 (N_45757,N_36820,N_33110);
or U45758 (N_45758,N_34720,N_32952);
nand U45759 (N_45759,N_34400,N_35701);
nand U45760 (N_45760,N_30372,N_38377);
nor U45761 (N_45761,N_36138,N_30685);
nor U45762 (N_45762,N_39449,N_33978);
nand U45763 (N_45763,N_34202,N_33249);
nand U45764 (N_45764,N_34628,N_39973);
nor U45765 (N_45765,N_31812,N_36813);
or U45766 (N_45766,N_37422,N_38216);
or U45767 (N_45767,N_36124,N_39931);
nor U45768 (N_45768,N_34570,N_34039);
or U45769 (N_45769,N_39471,N_37121);
nor U45770 (N_45770,N_39165,N_39837);
and U45771 (N_45771,N_37166,N_38842);
nor U45772 (N_45772,N_34730,N_38772);
nor U45773 (N_45773,N_31390,N_38285);
and U45774 (N_45774,N_31248,N_30294);
nand U45775 (N_45775,N_39775,N_30985);
or U45776 (N_45776,N_32502,N_38977);
xnor U45777 (N_45777,N_31073,N_34951);
nand U45778 (N_45778,N_30839,N_35390);
nand U45779 (N_45779,N_33912,N_33272);
and U45780 (N_45780,N_31708,N_34678);
or U45781 (N_45781,N_37177,N_38449);
or U45782 (N_45782,N_38317,N_31868);
nor U45783 (N_45783,N_36091,N_37106);
and U45784 (N_45784,N_35461,N_34101);
nand U45785 (N_45785,N_38553,N_32924);
nor U45786 (N_45786,N_38885,N_36177);
nand U45787 (N_45787,N_38343,N_35334);
nor U45788 (N_45788,N_37021,N_36552);
or U45789 (N_45789,N_34781,N_33823);
nor U45790 (N_45790,N_33119,N_31750);
nand U45791 (N_45791,N_35671,N_35860);
or U45792 (N_45792,N_31152,N_33085);
and U45793 (N_45793,N_30390,N_34447);
nand U45794 (N_45794,N_30311,N_30551);
nor U45795 (N_45795,N_37726,N_32496);
nand U45796 (N_45796,N_36068,N_36483);
xnor U45797 (N_45797,N_37315,N_35579);
nor U45798 (N_45798,N_36423,N_30395);
nand U45799 (N_45799,N_39981,N_36584);
nor U45800 (N_45800,N_30335,N_32893);
nand U45801 (N_45801,N_37446,N_35821);
and U45802 (N_45802,N_31551,N_37558);
nor U45803 (N_45803,N_36735,N_39287);
and U45804 (N_45804,N_39837,N_38626);
or U45805 (N_45805,N_34602,N_35499);
xor U45806 (N_45806,N_34725,N_32285);
or U45807 (N_45807,N_37103,N_32975);
nor U45808 (N_45808,N_35720,N_34659);
nor U45809 (N_45809,N_39743,N_37628);
and U45810 (N_45810,N_36263,N_35260);
nor U45811 (N_45811,N_31730,N_32087);
or U45812 (N_45812,N_35013,N_38676);
and U45813 (N_45813,N_35984,N_36700);
nor U45814 (N_45814,N_37570,N_33573);
or U45815 (N_45815,N_31584,N_38698);
xnor U45816 (N_45816,N_34816,N_33125);
and U45817 (N_45817,N_30044,N_34633);
xnor U45818 (N_45818,N_33619,N_38946);
or U45819 (N_45819,N_31293,N_31287);
or U45820 (N_45820,N_31988,N_31311);
nand U45821 (N_45821,N_39127,N_39007);
nor U45822 (N_45822,N_38513,N_38236);
and U45823 (N_45823,N_34298,N_34495);
xnor U45824 (N_45824,N_39702,N_32396);
nor U45825 (N_45825,N_31613,N_34399);
or U45826 (N_45826,N_31607,N_34926);
and U45827 (N_45827,N_31683,N_33153);
xor U45828 (N_45828,N_33836,N_32628);
nor U45829 (N_45829,N_32894,N_39100);
nor U45830 (N_45830,N_37557,N_34548);
and U45831 (N_45831,N_36706,N_37034);
and U45832 (N_45832,N_31626,N_32185);
or U45833 (N_45833,N_37644,N_32047);
and U45834 (N_45834,N_39195,N_34239);
nand U45835 (N_45835,N_32014,N_39844);
nand U45836 (N_45836,N_36417,N_35757);
nor U45837 (N_45837,N_34593,N_36263);
nand U45838 (N_45838,N_32430,N_32089);
nand U45839 (N_45839,N_35363,N_34203);
or U45840 (N_45840,N_39349,N_32145);
and U45841 (N_45841,N_37743,N_37933);
xnor U45842 (N_45842,N_34308,N_39202);
and U45843 (N_45843,N_39667,N_35681);
or U45844 (N_45844,N_34066,N_34475);
nand U45845 (N_45845,N_33897,N_37261);
or U45846 (N_45846,N_34508,N_31935);
nand U45847 (N_45847,N_34944,N_36561);
nand U45848 (N_45848,N_37038,N_31910);
nand U45849 (N_45849,N_33941,N_39898);
and U45850 (N_45850,N_38824,N_32688);
or U45851 (N_45851,N_36557,N_35832);
nor U45852 (N_45852,N_39644,N_30310);
xnor U45853 (N_45853,N_38385,N_35457);
or U45854 (N_45854,N_39275,N_34562);
nand U45855 (N_45855,N_37237,N_33379);
nor U45856 (N_45856,N_31556,N_34034);
xnor U45857 (N_45857,N_33921,N_33050);
nand U45858 (N_45858,N_33862,N_30625);
xnor U45859 (N_45859,N_37412,N_36694);
or U45860 (N_45860,N_32634,N_33417);
or U45861 (N_45861,N_31160,N_34342);
nand U45862 (N_45862,N_37764,N_32786);
and U45863 (N_45863,N_32673,N_38175);
nor U45864 (N_45864,N_34980,N_37494);
nand U45865 (N_45865,N_32575,N_31197);
nand U45866 (N_45866,N_39009,N_31757);
and U45867 (N_45867,N_32729,N_34077);
nand U45868 (N_45868,N_38295,N_30325);
xnor U45869 (N_45869,N_38343,N_31620);
or U45870 (N_45870,N_35215,N_31674);
nand U45871 (N_45871,N_37958,N_30271);
and U45872 (N_45872,N_36763,N_33057);
or U45873 (N_45873,N_35449,N_33463);
and U45874 (N_45874,N_36445,N_33055);
nand U45875 (N_45875,N_36602,N_34837);
or U45876 (N_45876,N_38328,N_34827);
and U45877 (N_45877,N_32610,N_35358);
nand U45878 (N_45878,N_36395,N_39731);
nor U45879 (N_45879,N_33155,N_30086);
nor U45880 (N_45880,N_34939,N_31135);
or U45881 (N_45881,N_33472,N_32983);
or U45882 (N_45882,N_36368,N_32115);
nand U45883 (N_45883,N_33277,N_31151);
nand U45884 (N_45884,N_32451,N_38429);
and U45885 (N_45885,N_33850,N_30260);
nand U45886 (N_45886,N_39157,N_30677);
nor U45887 (N_45887,N_34939,N_34256);
or U45888 (N_45888,N_38559,N_36428);
and U45889 (N_45889,N_34827,N_38271);
or U45890 (N_45890,N_31685,N_30546);
nor U45891 (N_45891,N_31512,N_33766);
or U45892 (N_45892,N_30332,N_39779);
or U45893 (N_45893,N_33175,N_37879);
nor U45894 (N_45894,N_30290,N_33304);
xor U45895 (N_45895,N_37981,N_30803);
nand U45896 (N_45896,N_33827,N_32039);
or U45897 (N_45897,N_35571,N_31603);
xnor U45898 (N_45898,N_31417,N_33527);
nand U45899 (N_45899,N_30108,N_37235);
or U45900 (N_45900,N_33998,N_37176);
nor U45901 (N_45901,N_37471,N_34815);
nor U45902 (N_45902,N_38129,N_38273);
nand U45903 (N_45903,N_36357,N_32449);
nor U45904 (N_45904,N_31422,N_35771);
or U45905 (N_45905,N_35379,N_38917);
and U45906 (N_45906,N_34589,N_38263);
xor U45907 (N_45907,N_30833,N_31408);
nor U45908 (N_45908,N_39953,N_37756);
xor U45909 (N_45909,N_32136,N_32302);
nand U45910 (N_45910,N_35189,N_36862);
or U45911 (N_45911,N_36625,N_34237);
or U45912 (N_45912,N_34434,N_32127);
nor U45913 (N_45913,N_34269,N_35369);
or U45914 (N_45914,N_36944,N_37029);
nand U45915 (N_45915,N_37400,N_34934);
or U45916 (N_45916,N_34417,N_34654);
nand U45917 (N_45917,N_31238,N_35863);
or U45918 (N_45918,N_38644,N_34115);
nor U45919 (N_45919,N_32774,N_30501);
or U45920 (N_45920,N_30228,N_32531);
and U45921 (N_45921,N_33557,N_37132);
or U45922 (N_45922,N_33116,N_35749);
xnor U45923 (N_45923,N_30251,N_31363);
nand U45924 (N_45924,N_35361,N_36580);
or U45925 (N_45925,N_39741,N_36125);
or U45926 (N_45926,N_31791,N_32155);
or U45927 (N_45927,N_38389,N_30746);
nor U45928 (N_45928,N_33637,N_36154);
nand U45929 (N_45929,N_35515,N_36670);
and U45930 (N_45930,N_35056,N_36659);
nor U45931 (N_45931,N_37819,N_32162);
xor U45932 (N_45932,N_34625,N_35812);
or U45933 (N_45933,N_36860,N_37242);
xnor U45934 (N_45934,N_38682,N_36785);
nand U45935 (N_45935,N_30761,N_35231);
or U45936 (N_45936,N_31215,N_31090);
and U45937 (N_45937,N_30130,N_35032);
nand U45938 (N_45938,N_37092,N_39691);
and U45939 (N_45939,N_34855,N_30800);
nand U45940 (N_45940,N_38214,N_35531);
and U45941 (N_45941,N_35072,N_39871);
nor U45942 (N_45942,N_34570,N_34485);
or U45943 (N_45943,N_36417,N_36924);
or U45944 (N_45944,N_30963,N_31335);
or U45945 (N_45945,N_33802,N_39798);
and U45946 (N_45946,N_37667,N_31001);
nor U45947 (N_45947,N_33163,N_30153);
nand U45948 (N_45948,N_38563,N_35450);
nor U45949 (N_45949,N_39570,N_33764);
or U45950 (N_45950,N_37264,N_33738);
or U45951 (N_45951,N_36023,N_34668);
or U45952 (N_45952,N_39745,N_30695);
or U45953 (N_45953,N_33990,N_37487);
or U45954 (N_45954,N_30875,N_35168);
nor U45955 (N_45955,N_35170,N_32425);
nand U45956 (N_45956,N_37869,N_30742);
and U45957 (N_45957,N_30492,N_36751);
nor U45958 (N_45958,N_39164,N_36743);
nand U45959 (N_45959,N_39259,N_30030);
and U45960 (N_45960,N_30826,N_31866);
nor U45961 (N_45961,N_32314,N_35129);
nand U45962 (N_45962,N_34790,N_38586);
nor U45963 (N_45963,N_33924,N_36020);
nand U45964 (N_45964,N_39125,N_33773);
xnor U45965 (N_45965,N_36675,N_31713);
nor U45966 (N_45966,N_38816,N_31522);
and U45967 (N_45967,N_36599,N_36743);
nand U45968 (N_45968,N_36119,N_36094);
xnor U45969 (N_45969,N_36478,N_32605);
xnor U45970 (N_45970,N_31434,N_33386);
nor U45971 (N_45971,N_32653,N_30082);
nand U45972 (N_45972,N_36244,N_36885);
nor U45973 (N_45973,N_34716,N_39349);
or U45974 (N_45974,N_38770,N_32615);
nand U45975 (N_45975,N_34709,N_35004);
nor U45976 (N_45976,N_38654,N_37901);
nand U45977 (N_45977,N_33432,N_31951);
and U45978 (N_45978,N_34136,N_31150);
nor U45979 (N_45979,N_37748,N_34877);
nor U45980 (N_45980,N_30855,N_30884);
nor U45981 (N_45981,N_30398,N_38969);
or U45982 (N_45982,N_38922,N_34782);
or U45983 (N_45983,N_32639,N_37189);
or U45984 (N_45984,N_36113,N_36244);
and U45985 (N_45985,N_36060,N_31262);
and U45986 (N_45986,N_35557,N_39257);
or U45987 (N_45987,N_35777,N_30356);
nor U45988 (N_45988,N_39566,N_35819);
nand U45989 (N_45989,N_31082,N_39729);
xnor U45990 (N_45990,N_39829,N_39267);
xor U45991 (N_45991,N_37729,N_39669);
nor U45992 (N_45992,N_38507,N_32394);
nor U45993 (N_45993,N_32366,N_36332);
and U45994 (N_45994,N_32070,N_31221);
or U45995 (N_45995,N_39330,N_33929);
xor U45996 (N_45996,N_32087,N_34379);
and U45997 (N_45997,N_38068,N_30269);
xor U45998 (N_45998,N_37995,N_39659);
nand U45999 (N_45999,N_33851,N_30457);
and U46000 (N_46000,N_36432,N_35264);
and U46001 (N_46001,N_39517,N_34572);
and U46002 (N_46002,N_36773,N_36817);
nand U46003 (N_46003,N_36748,N_31832);
nand U46004 (N_46004,N_39950,N_36609);
nand U46005 (N_46005,N_33449,N_35331);
nand U46006 (N_46006,N_32805,N_37306);
and U46007 (N_46007,N_31619,N_36162);
nor U46008 (N_46008,N_32949,N_39967);
nor U46009 (N_46009,N_31820,N_34396);
nor U46010 (N_46010,N_34482,N_34549);
or U46011 (N_46011,N_38896,N_36992);
or U46012 (N_46012,N_37371,N_35139);
nand U46013 (N_46013,N_35906,N_36456);
and U46014 (N_46014,N_34838,N_33797);
nor U46015 (N_46015,N_38343,N_34923);
or U46016 (N_46016,N_31550,N_34347);
and U46017 (N_46017,N_39301,N_38522);
or U46018 (N_46018,N_36905,N_30820);
and U46019 (N_46019,N_30608,N_36810);
nor U46020 (N_46020,N_34761,N_32609);
and U46021 (N_46021,N_34202,N_33299);
xor U46022 (N_46022,N_33422,N_37044);
nand U46023 (N_46023,N_30790,N_31666);
or U46024 (N_46024,N_37748,N_34840);
and U46025 (N_46025,N_35929,N_31508);
and U46026 (N_46026,N_39658,N_33281);
nor U46027 (N_46027,N_32011,N_36735);
and U46028 (N_46028,N_36191,N_36754);
or U46029 (N_46029,N_31908,N_37916);
and U46030 (N_46030,N_36431,N_30628);
nand U46031 (N_46031,N_32056,N_39516);
nand U46032 (N_46032,N_30534,N_36217);
and U46033 (N_46033,N_33386,N_36342);
xor U46034 (N_46034,N_32679,N_38785);
nand U46035 (N_46035,N_33423,N_32011);
xor U46036 (N_46036,N_32944,N_30746);
nand U46037 (N_46037,N_34639,N_30454);
and U46038 (N_46038,N_36946,N_36513);
and U46039 (N_46039,N_37294,N_35912);
xnor U46040 (N_46040,N_38861,N_35658);
nor U46041 (N_46041,N_37674,N_30943);
nand U46042 (N_46042,N_37891,N_36000);
xnor U46043 (N_46043,N_30423,N_37891);
xor U46044 (N_46044,N_30620,N_31874);
and U46045 (N_46045,N_38994,N_31459);
and U46046 (N_46046,N_37901,N_31447);
or U46047 (N_46047,N_38345,N_31837);
nand U46048 (N_46048,N_37207,N_37866);
or U46049 (N_46049,N_30634,N_39778);
or U46050 (N_46050,N_32141,N_31387);
xor U46051 (N_46051,N_39699,N_33069);
or U46052 (N_46052,N_37636,N_32256);
nand U46053 (N_46053,N_38047,N_35654);
nor U46054 (N_46054,N_39820,N_33995);
and U46055 (N_46055,N_30270,N_38298);
and U46056 (N_46056,N_30781,N_30941);
xor U46057 (N_46057,N_33857,N_36948);
and U46058 (N_46058,N_32260,N_30126);
or U46059 (N_46059,N_36023,N_35023);
xnor U46060 (N_46060,N_33264,N_35438);
or U46061 (N_46061,N_30907,N_30914);
nor U46062 (N_46062,N_34524,N_36242);
xor U46063 (N_46063,N_39022,N_34760);
and U46064 (N_46064,N_30416,N_35788);
and U46065 (N_46065,N_32883,N_34066);
nand U46066 (N_46066,N_31674,N_37302);
and U46067 (N_46067,N_34181,N_31713);
nor U46068 (N_46068,N_31637,N_30806);
and U46069 (N_46069,N_34503,N_35736);
nor U46070 (N_46070,N_33863,N_39689);
nand U46071 (N_46071,N_37440,N_38340);
nor U46072 (N_46072,N_34313,N_31512);
or U46073 (N_46073,N_38795,N_31267);
or U46074 (N_46074,N_33351,N_35223);
or U46075 (N_46075,N_38821,N_32822);
nor U46076 (N_46076,N_35910,N_35836);
nand U46077 (N_46077,N_38973,N_39641);
nor U46078 (N_46078,N_30558,N_32522);
or U46079 (N_46079,N_36264,N_39081);
nor U46080 (N_46080,N_33739,N_37461);
nand U46081 (N_46081,N_35419,N_33326);
and U46082 (N_46082,N_37323,N_34158);
nand U46083 (N_46083,N_39449,N_31767);
nand U46084 (N_46084,N_32361,N_36400);
nor U46085 (N_46085,N_35736,N_36324);
and U46086 (N_46086,N_35325,N_38266);
xnor U46087 (N_46087,N_39409,N_33199);
nand U46088 (N_46088,N_39974,N_35969);
or U46089 (N_46089,N_36581,N_38656);
xor U46090 (N_46090,N_36350,N_38874);
nand U46091 (N_46091,N_38620,N_38795);
or U46092 (N_46092,N_33609,N_34375);
and U46093 (N_46093,N_33665,N_39867);
nand U46094 (N_46094,N_31774,N_34895);
nand U46095 (N_46095,N_39073,N_37905);
nand U46096 (N_46096,N_31177,N_36794);
nand U46097 (N_46097,N_35980,N_34243);
and U46098 (N_46098,N_36887,N_36490);
nor U46099 (N_46099,N_30331,N_38381);
and U46100 (N_46100,N_36796,N_34921);
or U46101 (N_46101,N_30614,N_32370);
or U46102 (N_46102,N_36940,N_35876);
nand U46103 (N_46103,N_38507,N_31509);
nand U46104 (N_46104,N_34196,N_30770);
xnor U46105 (N_46105,N_37306,N_39405);
xnor U46106 (N_46106,N_35604,N_33077);
nand U46107 (N_46107,N_36781,N_32326);
xor U46108 (N_46108,N_37945,N_31304);
nor U46109 (N_46109,N_34112,N_32411);
or U46110 (N_46110,N_37257,N_32179);
nand U46111 (N_46111,N_33180,N_35816);
nor U46112 (N_46112,N_33839,N_35042);
and U46113 (N_46113,N_37479,N_31283);
and U46114 (N_46114,N_37344,N_30108);
nor U46115 (N_46115,N_35391,N_34590);
nand U46116 (N_46116,N_36178,N_31681);
xor U46117 (N_46117,N_37111,N_31012);
nand U46118 (N_46118,N_38795,N_33211);
xnor U46119 (N_46119,N_31515,N_30617);
nand U46120 (N_46120,N_35671,N_32744);
nand U46121 (N_46121,N_30411,N_39477);
or U46122 (N_46122,N_39489,N_32928);
or U46123 (N_46123,N_33283,N_36436);
nor U46124 (N_46124,N_33649,N_32934);
nor U46125 (N_46125,N_35212,N_34951);
nor U46126 (N_46126,N_32046,N_37668);
nand U46127 (N_46127,N_36612,N_33693);
nand U46128 (N_46128,N_37720,N_31405);
and U46129 (N_46129,N_32299,N_30780);
nand U46130 (N_46130,N_31659,N_37890);
and U46131 (N_46131,N_34107,N_39131);
nor U46132 (N_46132,N_38053,N_38121);
or U46133 (N_46133,N_37775,N_31907);
nand U46134 (N_46134,N_38582,N_35477);
nand U46135 (N_46135,N_31619,N_30122);
xor U46136 (N_46136,N_32784,N_34364);
nor U46137 (N_46137,N_38054,N_38138);
or U46138 (N_46138,N_36221,N_37290);
nand U46139 (N_46139,N_34202,N_33508);
and U46140 (N_46140,N_32199,N_39766);
and U46141 (N_46141,N_31584,N_31290);
nand U46142 (N_46142,N_37047,N_39899);
or U46143 (N_46143,N_31752,N_34076);
nor U46144 (N_46144,N_37019,N_37711);
nor U46145 (N_46145,N_34586,N_30752);
xnor U46146 (N_46146,N_31250,N_37778);
nand U46147 (N_46147,N_38558,N_37423);
and U46148 (N_46148,N_39331,N_38927);
xnor U46149 (N_46149,N_35999,N_37066);
nor U46150 (N_46150,N_38760,N_36112);
or U46151 (N_46151,N_39808,N_31112);
nand U46152 (N_46152,N_30058,N_37376);
xnor U46153 (N_46153,N_36348,N_34464);
nor U46154 (N_46154,N_36516,N_39808);
nor U46155 (N_46155,N_39417,N_39012);
and U46156 (N_46156,N_36413,N_37973);
or U46157 (N_46157,N_34544,N_39604);
xnor U46158 (N_46158,N_39740,N_38714);
nand U46159 (N_46159,N_38680,N_32198);
and U46160 (N_46160,N_36160,N_34247);
and U46161 (N_46161,N_33698,N_33103);
or U46162 (N_46162,N_33632,N_31578);
nand U46163 (N_46163,N_32386,N_36472);
nand U46164 (N_46164,N_38404,N_36512);
or U46165 (N_46165,N_38503,N_39804);
nand U46166 (N_46166,N_32411,N_39580);
nor U46167 (N_46167,N_38706,N_35329);
or U46168 (N_46168,N_35318,N_39545);
nor U46169 (N_46169,N_33901,N_38167);
and U46170 (N_46170,N_36738,N_36399);
xnor U46171 (N_46171,N_30717,N_36663);
xor U46172 (N_46172,N_38994,N_31311);
nor U46173 (N_46173,N_39129,N_31986);
and U46174 (N_46174,N_38825,N_32972);
nand U46175 (N_46175,N_35603,N_36288);
nor U46176 (N_46176,N_30784,N_31515);
nor U46177 (N_46177,N_32806,N_34899);
and U46178 (N_46178,N_35480,N_35287);
and U46179 (N_46179,N_30241,N_37614);
or U46180 (N_46180,N_36375,N_34723);
nor U46181 (N_46181,N_33949,N_37130);
and U46182 (N_46182,N_39743,N_31946);
nor U46183 (N_46183,N_38166,N_35350);
or U46184 (N_46184,N_35734,N_37460);
or U46185 (N_46185,N_37562,N_35034);
nand U46186 (N_46186,N_30206,N_38756);
or U46187 (N_46187,N_36668,N_37785);
nand U46188 (N_46188,N_33104,N_38280);
nand U46189 (N_46189,N_38987,N_37724);
nor U46190 (N_46190,N_34719,N_37918);
nor U46191 (N_46191,N_34907,N_30672);
and U46192 (N_46192,N_32564,N_31735);
xnor U46193 (N_46193,N_38760,N_34059);
and U46194 (N_46194,N_36687,N_31701);
nor U46195 (N_46195,N_30865,N_34431);
or U46196 (N_46196,N_35865,N_35435);
xor U46197 (N_46197,N_32867,N_32977);
nand U46198 (N_46198,N_30344,N_39509);
nand U46199 (N_46199,N_30546,N_36449);
and U46200 (N_46200,N_35418,N_38840);
nand U46201 (N_46201,N_31109,N_36303);
and U46202 (N_46202,N_34578,N_38973);
and U46203 (N_46203,N_35105,N_37572);
and U46204 (N_46204,N_34868,N_34844);
xnor U46205 (N_46205,N_39458,N_39290);
nor U46206 (N_46206,N_33608,N_32460);
nand U46207 (N_46207,N_34713,N_32724);
nor U46208 (N_46208,N_33497,N_33098);
nand U46209 (N_46209,N_36606,N_38944);
or U46210 (N_46210,N_31267,N_37050);
nor U46211 (N_46211,N_31530,N_30624);
or U46212 (N_46212,N_37261,N_35113);
and U46213 (N_46213,N_31606,N_33910);
or U46214 (N_46214,N_34371,N_34880);
nand U46215 (N_46215,N_36687,N_31509);
and U46216 (N_46216,N_32458,N_35904);
nor U46217 (N_46217,N_34134,N_39233);
nor U46218 (N_46218,N_38384,N_32775);
and U46219 (N_46219,N_37967,N_34765);
and U46220 (N_46220,N_31393,N_31220);
nand U46221 (N_46221,N_31953,N_37192);
nand U46222 (N_46222,N_32994,N_33789);
nor U46223 (N_46223,N_37030,N_31441);
or U46224 (N_46224,N_36992,N_36594);
or U46225 (N_46225,N_33397,N_37585);
nor U46226 (N_46226,N_36584,N_30071);
and U46227 (N_46227,N_31765,N_33444);
nor U46228 (N_46228,N_30743,N_33053);
and U46229 (N_46229,N_34160,N_37813);
and U46230 (N_46230,N_38329,N_36192);
or U46231 (N_46231,N_32935,N_35588);
nor U46232 (N_46232,N_32602,N_35569);
xnor U46233 (N_46233,N_38076,N_30906);
nand U46234 (N_46234,N_35271,N_31818);
or U46235 (N_46235,N_30737,N_36652);
and U46236 (N_46236,N_31796,N_31204);
nand U46237 (N_46237,N_30722,N_31836);
xnor U46238 (N_46238,N_37299,N_33773);
and U46239 (N_46239,N_35053,N_33858);
and U46240 (N_46240,N_34862,N_32732);
nor U46241 (N_46241,N_34645,N_34150);
nor U46242 (N_46242,N_36000,N_31026);
nand U46243 (N_46243,N_31148,N_38943);
nand U46244 (N_46244,N_34373,N_38402);
and U46245 (N_46245,N_33165,N_38688);
or U46246 (N_46246,N_32910,N_30181);
or U46247 (N_46247,N_37916,N_35688);
nand U46248 (N_46248,N_35850,N_36743);
nand U46249 (N_46249,N_32675,N_37812);
nor U46250 (N_46250,N_37815,N_30187);
nand U46251 (N_46251,N_37925,N_38157);
nor U46252 (N_46252,N_36955,N_39282);
nor U46253 (N_46253,N_30777,N_31728);
and U46254 (N_46254,N_39865,N_31354);
and U46255 (N_46255,N_39365,N_38017);
or U46256 (N_46256,N_36969,N_38379);
nand U46257 (N_46257,N_38554,N_37392);
or U46258 (N_46258,N_31732,N_31771);
and U46259 (N_46259,N_37804,N_32049);
or U46260 (N_46260,N_37646,N_37162);
nor U46261 (N_46261,N_34417,N_36524);
nor U46262 (N_46262,N_32492,N_38757);
nor U46263 (N_46263,N_33144,N_34274);
and U46264 (N_46264,N_35657,N_38645);
nor U46265 (N_46265,N_34970,N_30897);
xnor U46266 (N_46266,N_30410,N_36800);
or U46267 (N_46267,N_34954,N_37611);
or U46268 (N_46268,N_35921,N_38193);
nor U46269 (N_46269,N_31605,N_39462);
nand U46270 (N_46270,N_34665,N_37756);
or U46271 (N_46271,N_32740,N_31584);
xor U46272 (N_46272,N_32249,N_34462);
nor U46273 (N_46273,N_39748,N_31497);
nor U46274 (N_46274,N_30326,N_31300);
or U46275 (N_46275,N_34371,N_34699);
nand U46276 (N_46276,N_34462,N_34032);
xnor U46277 (N_46277,N_38350,N_30983);
nor U46278 (N_46278,N_39231,N_31713);
nor U46279 (N_46279,N_38336,N_35760);
and U46280 (N_46280,N_39704,N_36451);
and U46281 (N_46281,N_30687,N_33353);
nand U46282 (N_46282,N_34189,N_39665);
and U46283 (N_46283,N_37003,N_36638);
xor U46284 (N_46284,N_37443,N_38136);
and U46285 (N_46285,N_37444,N_34535);
nand U46286 (N_46286,N_36259,N_32570);
nand U46287 (N_46287,N_33555,N_38926);
and U46288 (N_46288,N_32592,N_34942);
nand U46289 (N_46289,N_32984,N_35233);
nand U46290 (N_46290,N_31443,N_32437);
and U46291 (N_46291,N_33575,N_34627);
and U46292 (N_46292,N_32191,N_37621);
and U46293 (N_46293,N_35900,N_37689);
nor U46294 (N_46294,N_36401,N_38271);
nor U46295 (N_46295,N_30890,N_32045);
nor U46296 (N_46296,N_36422,N_38683);
or U46297 (N_46297,N_32848,N_38064);
and U46298 (N_46298,N_36987,N_38281);
nor U46299 (N_46299,N_37688,N_39319);
and U46300 (N_46300,N_35917,N_35925);
nand U46301 (N_46301,N_31353,N_35443);
nand U46302 (N_46302,N_33155,N_39229);
and U46303 (N_46303,N_35447,N_31654);
and U46304 (N_46304,N_37797,N_38282);
nand U46305 (N_46305,N_39302,N_34830);
or U46306 (N_46306,N_37023,N_34622);
xor U46307 (N_46307,N_36518,N_33573);
and U46308 (N_46308,N_35597,N_35409);
nor U46309 (N_46309,N_38813,N_33216);
and U46310 (N_46310,N_34703,N_34482);
nor U46311 (N_46311,N_30995,N_39773);
or U46312 (N_46312,N_30165,N_30799);
nor U46313 (N_46313,N_37721,N_39362);
or U46314 (N_46314,N_34104,N_35104);
nand U46315 (N_46315,N_38326,N_33100);
or U46316 (N_46316,N_34470,N_34752);
nor U46317 (N_46317,N_31682,N_32853);
nand U46318 (N_46318,N_32389,N_34042);
and U46319 (N_46319,N_30377,N_38959);
and U46320 (N_46320,N_37369,N_38625);
nor U46321 (N_46321,N_34884,N_35693);
nand U46322 (N_46322,N_33362,N_32435);
or U46323 (N_46323,N_34923,N_31419);
nand U46324 (N_46324,N_34669,N_31230);
and U46325 (N_46325,N_34056,N_39299);
nor U46326 (N_46326,N_31380,N_31303);
xnor U46327 (N_46327,N_32322,N_34187);
xor U46328 (N_46328,N_37925,N_37626);
and U46329 (N_46329,N_37022,N_39271);
nor U46330 (N_46330,N_30134,N_38556);
nand U46331 (N_46331,N_36459,N_35318);
and U46332 (N_46332,N_30309,N_33713);
or U46333 (N_46333,N_34050,N_38823);
nand U46334 (N_46334,N_39878,N_30016);
and U46335 (N_46335,N_37369,N_31716);
or U46336 (N_46336,N_38381,N_31845);
xnor U46337 (N_46337,N_30220,N_38236);
nor U46338 (N_46338,N_37178,N_38610);
and U46339 (N_46339,N_30786,N_36956);
xnor U46340 (N_46340,N_39539,N_36158);
xnor U46341 (N_46341,N_39990,N_30627);
nor U46342 (N_46342,N_37731,N_39539);
nand U46343 (N_46343,N_34367,N_36352);
and U46344 (N_46344,N_37164,N_39060);
and U46345 (N_46345,N_39874,N_30466);
and U46346 (N_46346,N_37620,N_37339);
or U46347 (N_46347,N_38183,N_39566);
or U46348 (N_46348,N_31003,N_34259);
nor U46349 (N_46349,N_36311,N_33202);
nor U46350 (N_46350,N_31979,N_31609);
xor U46351 (N_46351,N_37787,N_38490);
or U46352 (N_46352,N_31277,N_37090);
nor U46353 (N_46353,N_39527,N_39034);
nand U46354 (N_46354,N_32519,N_36610);
nand U46355 (N_46355,N_35219,N_39370);
and U46356 (N_46356,N_36650,N_31069);
or U46357 (N_46357,N_36048,N_31618);
nand U46358 (N_46358,N_38926,N_34524);
nand U46359 (N_46359,N_31002,N_38672);
or U46360 (N_46360,N_37819,N_38719);
or U46361 (N_46361,N_37025,N_39956);
or U46362 (N_46362,N_35087,N_36532);
and U46363 (N_46363,N_31014,N_31369);
xor U46364 (N_46364,N_31491,N_38248);
and U46365 (N_46365,N_33376,N_32008);
or U46366 (N_46366,N_39893,N_31876);
and U46367 (N_46367,N_30165,N_35633);
and U46368 (N_46368,N_37275,N_32589);
or U46369 (N_46369,N_30228,N_32671);
nand U46370 (N_46370,N_34479,N_37918);
or U46371 (N_46371,N_39388,N_34866);
xnor U46372 (N_46372,N_39207,N_34607);
nand U46373 (N_46373,N_39564,N_36699);
nand U46374 (N_46374,N_34404,N_35847);
nand U46375 (N_46375,N_34167,N_34055);
nand U46376 (N_46376,N_39189,N_38720);
nand U46377 (N_46377,N_36623,N_34038);
and U46378 (N_46378,N_32282,N_39790);
nor U46379 (N_46379,N_36316,N_30294);
and U46380 (N_46380,N_31801,N_35848);
xor U46381 (N_46381,N_30879,N_33404);
and U46382 (N_46382,N_37023,N_38594);
nand U46383 (N_46383,N_37440,N_33982);
nor U46384 (N_46384,N_36127,N_32056);
nor U46385 (N_46385,N_39384,N_36463);
xor U46386 (N_46386,N_30697,N_37810);
xor U46387 (N_46387,N_34407,N_38721);
nor U46388 (N_46388,N_30441,N_35252);
nor U46389 (N_46389,N_35815,N_31681);
and U46390 (N_46390,N_33518,N_32201);
and U46391 (N_46391,N_32091,N_31713);
nor U46392 (N_46392,N_37657,N_35693);
or U46393 (N_46393,N_30626,N_36221);
and U46394 (N_46394,N_39441,N_36205);
or U46395 (N_46395,N_31305,N_37986);
xor U46396 (N_46396,N_34717,N_35830);
nand U46397 (N_46397,N_31194,N_36826);
and U46398 (N_46398,N_39866,N_37349);
nand U46399 (N_46399,N_38512,N_36900);
or U46400 (N_46400,N_34395,N_31736);
nor U46401 (N_46401,N_36463,N_38412);
or U46402 (N_46402,N_31279,N_30214);
nand U46403 (N_46403,N_31953,N_34853);
nand U46404 (N_46404,N_33335,N_35355);
or U46405 (N_46405,N_39295,N_35330);
nor U46406 (N_46406,N_33038,N_30381);
xnor U46407 (N_46407,N_32441,N_34715);
nand U46408 (N_46408,N_30778,N_37633);
and U46409 (N_46409,N_38470,N_36991);
nand U46410 (N_46410,N_36383,N_38400);
nand U46411 (N_46411,N_37396,N_32413);
or U46412 (N_46412,N_34534,N_30659);
nand U46413 (N_46413,N_33664,N_31068);
nor U46414 (N_46414,N_38121,N_34595);
nand U46415 (N_46415,N_37192,N_32138);
nor U46416 (N_46416,N_34366,N_35042);
nand U46417 (N_46417,N_37370,N_30789);
nor U46418 (N_46418,N_39270,N_33409);
nand U46419 (N_46419,N_30655,N_38606);
or U46420 (N_46420,N_39450,N_36682);
nand U46421 (N_46421,N_34475,N_37851);
nand U46422 (N_46422,N_31118,N_32750);
or U46423 (N_46423,N_38801,N_31200);
nor U46424 (N_46424,N_36161,N_37719);
xor U46425 (N_46425,N_36147,N_33518);
or U46426 (N_46426,N_33903,N_32060);
nand U46427 (N_46427,N_39075,N_39630);
or U46428 (N_46428,N_32523,N_34062);
or U46429 (N_46429,N_37078,N_35831);
nand U46430 (N_46430,N_31212,N_36710);
or U46431 (N_46431,N_34555,N_32990);
nor U46432 (N_46432,N_33159,N_36705);
nor U46433 (N_46433,N_38429,N_30549);
xnor U46434 (N_46434,N_33800,N_35657);
nand U46435 (N_46435,N_35043,N_31951);
or U46436 (N_46436,N_32401,N_39693);
or U46437 (N_46437,N_38385,N_32258);
and U46438 (N_46438,N_35691,N_38887);
or U46439 (N_46439,N_36907,N_30958);
and U46440 (N_46440,N_37601,N_31390);
nor U46441 (N_46441,N_39842,N_39936);
nor U46442 (N_46442,N_38919,N_32290);
or U46443 (N_46443,N_38372,N_38037);
or U46444 (N_46444,N_31311,N_31967);
and U46445 (N_46445,N_36319,N_37205);
or U46446 (N_46446,N_31935,N_36287);
and U46447 (N_46447,N_32274,N_39452);
and U46448 (N_46448,N_31022,N_37527);
nor U46449 (N_46449,N_32509,N_39946);
xnor U46450 (N_46450,N_35278,N_39680);
and U46451 (N_46451,N_38506,N_35313);
nor U46452 (N_46452,N_39759,N_34713);
and U46453 (N_46453,N_35749,N_35526);
nand U46454 (N_46454,N_35806,N_32250);
xor U46455 (N_46455,N_37309,N_33482);
or U46456 (N_46456,N_31841,N_30354);
nand U46457 (N_46457,N_30333,N_30519);
or U46458 (N_46458,N_34481,N_38958);
xor U46459 (N_46459,N_37587,N_35123);
nand U46460 (N_46460,N_34428,N_35238);
and U46461 (N_46461,N_35662,N_32197);
and U46462 (N_46462,N_30353,N_38950);
nand U46463 (N_46463,N_34367,N_31529);
or U46464 (N_46464,N_31409,N_34711);
nand U46465 (N_46465,N_35097,N_38494);
nand U46466 (N_46466,N_36040,N_36206);
xnor U46467 (N_46467,N_32690,N_38554);
or U46468 (N_46468,N_32444,N_39396);
and U46469 (N_46469,N_38814,N_35857);
nand U46470 (N_46470,N_36907,N_39542);
nor U46471 (N_46471,N_31236,N_37343);
and U46472 (N_46472,N_30506,N_35223);
nor U46473 (N_46473,N_38715,N_37790);
and U46474 (N_46474,N_33318,N_33253);
nand U46475 (N_46475,N_35419,N_38122);
nand U46476 (N_46476,N_32421,N_35855);
nor U46477 (N_46477,N_31366,N_36376);
or U46478 (N_46478,N_38158,N_30113);
or U46479 (N_46479,N_32455,N_37758);
or U46480 (N_46480,N_35842,N_39277);
nor U46481 (N_46481,N_35617,N_35053);
or U46482 (N_46482,N_34472,N_34461);
xnor U46483 (N_46483,N_34791,N_37457);
nand U46484 (N_46484,N_37199,N_39444);
nor U46485 (N_46485,N_30485,N_39147);
and U46486 (N_46486,N_37886,N_39283);
or U46487 (N_46487,N_39545,N_38375);
nand U46488 (N_46488,N_36875,N_35374);
and U46489 (N_46489,N_34286,N_33410);
nor U46490 (N_46490,N_32577,N_31850);
nand U46491 (N_46491,N_37460,N_35438);
nand U46492 (N_46492,N_30995,N_34959);
nand U46493 (N_46493,N_32475,N_33133);
nand U46494 (N_46494,N_34435,N_37038);
nand U46495 (N_46495,N_38315,N_33233);
and U46496 (N_46496,N_30836,N_35655);
nor U46497 (N_46497,N_31733,N_34493);
or U46498 (N_46498,N_34598,N_30674);
or U46499 (N_46499,N_33289,N_32718);
nor U46500 (N_46500,N_31395,N_33723);
or U46501 (N_46501,N_37073,N_34453);
and U46502 (N_46502,N_36453,N_36319);
nand U46503 (N_46503,N_34098,N_37234);
or U46504 (N_46504,N_34952,N_34692);
and U46505 (N_46505,N_37039,N_36287);
nor U46506 (N_46506,N_37870,N_32134);
and U46507 (N_46507,N_38681,N_37704);
or U46508 (N_46508,N_31078,N_33484);
nor U46509 (N_46509,N_38499,N_38788);
nand U46510 (N_46510,N_31847,N_38539);
nand U46511 (N_46511,N_39218,N_31844);
or U46512 (N_46512,N_38361,N_36961);
nor U46513 (N_46513,N_37998,N_36753);
xnor U46514 (N_46514,N_36856,N_30381);
and U46515 (N_46515,N_33846,N_39113);
nand U46516 (N_46516,N_37284,N_32664);
nand U46517 (N_46517,N_37938,N_32790);
nor U46518 (N_46518,N_37995,N_38590);
and U46519 (N_46519,N_35359,N_36298);
nor U46520 (N_46520,N_34451,N_31529);
nand U46521 (N_46521,N_35834,N_31389);
or U46522 (N_46522,N_36113,N_33691);
nor U46523 (N_46523,N_30495,N_38421);
xnor U46524 (N_46524,N_35212,N_30051);
nand U46525 (N_46525,N_39531,N_33752);
or U46526 (N_46526,N_30005,N_37639);
nor U46527 (N_46527,N_39927,N_32554);
or U46528 (N_46528,N_35413,N_37199);
nand U46529 (N_46529,N_38504,N_37524);
and U46530 (N_46530,N_30637,N_36331);
or U46531 (N_46531,N_32937,N_38034);
nor U46532 (N_46532,N_35109,N_38342);
or U46533 (N_46533,N_34171,N_38896);
and U46534 (N_46534,N_31798,N_38775);
nand U46535 (N_46535,N_36759,N_34695);
or U46536 (N_46536,N_30834,N_31941);
nor U46537 (N_46537,N_34358,N_38721);
or U46538 (N_46538,N_37251,N_32012);
nand U46539 (N_46539,N_33146,N_38981);
nor U46540 (N_46540,N_39611,N_30362);
or U46541 (N_46541,N_36349,N_39465);
nor U46542 (N_46542,N_37660,N_39685);
xnor U46543 (N_46543,N_39541,N_33004);
or U46544 (N_46544,N_36143,N_37985);
or U46545 (N_46545,N_34417,N_37923);
nand U46546 (N_46546,N_36082,N_38249);
nand U46547 (N_46547,N_33387,N_38391);
nand U46548 (N_46548,N_39273,N_35668);
nor U46549 (N_46549,N_31352,N_30987);
or U46550 (N_46550,N_35360,N_30758);
or U46551 (N_46551,N_34404,N_35589);
and U46552 (N_46552,N_31304,N_31339);
or U46553 (N_46553,N_39433,N_32194);
or U46554 (N_46554,N_37797,N_39251);
xnor U46555 (N_46555,N_34279,N_34696);
nand U46556 (N_46556,N_35292,N_34451);
or U46557 (N_46557,N_31153,N_36506);
or U46558 (N_46558,N_37619,N_36388);
nand U46559 (N_46559,N_38842,N_34719);
and U46560 (N_46560,N_39184,N_33331);
nor U46561 (N_46561,N_39096,N_39152);
nand U46562 (N_46562,N_38004,N_34698);
nor U46563 (N_46563,N_31458,N_38418);
xnor U46564 (N_46564,N_35476,N_31468);
nor U46565 (N_46565,N_39664,N_35082);
xnor U46566 (N_46566,N_33906,N_37185);
xor U46567 (N_46567,N_36839,N_38033);
and U46568 (N_46568,N_38228,N_34630);
nor U46569 (N_46569,N_33984,N_39630);
or U46570 (N_46570,N_37797,N_35213);
nand U46571 (N_46571,N_30905,N_36970);
nor U46572 (N_46572,N_33223,N_33365);
and U46573 (N_46573,N_35314,N_38242);
nor U46574 (N_46574,N_31039,N_36454);
or U46575 (N_46575,N_34191,N_32685);
nor U46576 (N_46576,N_37637,N_31305);
or U46577 (N_46577,N_32692,N_30648);
and U46578 (N_46578,N_39667,N_36605);
nand U46579 (N_46579,N_32578,N_37916);
nand U46580 (N_46580,N_39746,N_39533);
nor U46581 (N_46581,N_39642,N_37733);
or U46582 (N_46582,N_39375,N_31688);
or U46583 (N_46583,N_32657,N_34035);
nand U46584 (N_46584,N_32378,N_37697);
or U46585 (N_46585,N_30538,N_35471);
or U46586 (N_46586,N_37648,N_36501);
nand U46587 (N_46587,N_37493,N_32821);
or U46588 (N_46588,N_36833,N_31279);
or U46589 (N_46589,N_30542,N_30760);
nand U46590 (N_46590,N_38217,N_31808);
and U46591 (N_46591,N_33988,N_32883);
and U46592 (N_46592,N_30065,N_37550);
nor U46593 (N_46593,N_33295,N_33656);
and U46594 (N_46594,N_37936,N_36078);
nand U46595 (N_46595,N_32233,N_35771);
xnor U46596 (N_46596,N_32287,N_35636);
or U46597 (N_46597,N_37090,N_36171);
nand U46598 (N_46598,N_39023,N_30396);
and U46599 (N_46599,N_37293,N_31454);
or U46600 (N_46600,N_33674,N_36095);
or U46601 (N_46601,N_34290,N_32122);
and U46602 (N_46602,N_35808,N_38418);
nand U46603 (N_46603,N_38162,N_33051);
nor U46604 (N_46604,N_38189,N_36959);
nand U46605 (N_46605,N_32692,N_37092);
nor U46606 (N_46606,N_30034,N_34786);
or U46607 (N_46607,N_35240,N_35323);
nand U46608 (N_46608,N_38376,N_35964);
or U46609 (N_46609,N_31950,N_36994);
and U46610 (N_46610,N_30651,N_38793);
xnor U46611 (N_46611,N_30434,N_33028);
or U46612 (N_46612,N_39440,N_35811);
nor U46613 (N_46613,N_32546,N_30328);
or U46614 (N_46614,N_38546,N_37509);
nor U46615 (N_46615,N_31287,N_33585);
xnor U46616 (N_46616,N_39745,N_36717);
or U46617 (N_46617,N_39055,N_35349);
nand U46618 (N_46618,N_39400,N_37298);
nor U46619 (N_46619,N_38279,N_35550);
xor U46620 (N_46620,N_34154,N_39175);
and U46621 (N_46621,N_37843,N_36528);
or U46622 (N_46622,N_33939,N_30904);
nand U46623 (N_46623,N_35781,N_32678);
or U46624 (N_46624,N_34197,N_31854);
nor U46625 (N_46625,N_36147,N_39234);
or U46626 (N_46626,N_38885,N_31225);
nand U46627 (N_46627,N_33555,N_38025);
or U46628 (N_46628,N_38146,N_34945);
or U46629 (N_46629,N_37148,N_32509);
nor U46630 (N_46630,N_38888,N_31159);
xor U46631 (N_46631,N_33444,N_32018);
nand U46632 (N_46632,N_31105,N_31806);
nor U46633 (N_46633,N_33105,N_36135);
xnor U46634 (N_46634,N_31245,N_36049);
nor U46635 (N_46635,N_32283,N_32914);
and U46636 (N_46636,N_37223,N_35635);
or U46637 (N_46637,N_39291,N_39410);
and U46638 (N_46638,N_31619,N_34578);
and U46639 (N_46639,N_30877,N_38354);
or U46640 (N_46640,N_32206,N_34006);
and U46641 (N_46641,N_32335,N_30461);
nor U46642 (N_46642,N_39586,N_31488);
nor U46643 (N_46643,N_36380,N_35435);
xnor U46644 (N_46644,N_37291,N_31774);
or U46645 (N_46645,N_36224,N_38198);
nand U46646 (N_46646,N_31045,N_39929);
or U46647 (N_46647,N_32532,N_39524);
nand U46648 (N_46648,N_39597,N_30766);
nand U46649 (N_46649,N_38080,N_36559);
nor U46650 (N_46650,N_36395,N_33681);
nand U46651 (N_46651,N_33523,N_35983);
or U46652 (N_46652,N_31445,N_39526);
nand U46653 (N_46653,N_33725,N_34581);
xnor U46654 (N_46654,N_36368,N_31311);
and U46655 (N_46655,N_32150,N_33664);
or U46656 (N_46656,N_36330,N_31779);
nor U46657 (N_46657,N_39748,N_36109);
and U46658 (N_46658,N_36790,N_35376);
nor U46659 (N_46659,N_36341,N_34867);
nand U46660 (N_46660,N_35262,N_36679);
nand U46661 (N_46661,N_33866,N_35584);
nor U46662 (N_46662,N_33451,N_31087);
or U46663 (N_46663,N_30111,N_38802);
nor U46664 (N_46664,N_33668,N_34259);
nor U46665 (N_46665,N_38923,N_31940);
or U46666 (N_46666,N_31631,N_33252);
nor U46667 (N_46667,N_34489,N_37653);
nor U46668 (N_46668,N_30225,N_31598);
or U46669 (N_46669,N_39229,N_30325);
or U46670 (N_46670,N_36649,N_30897);
nand U46671 (N_46671,N_31843,N_38211);
nand U46672 (N_46672,N_38966,N_35605);
or U46673 (N_46673,N_35451,N_39674);
xnor U46674 (N_46674,N_37176,N_31774);
nor U46675 (N_46675,N_30807,N_32337);
or U46676 (N_46676,N_36778,N_34922);
nand U46677 (N_46677,N_38672,N_32878);
or U46678 (N_46678,N_39779,N_34208);
nand U46679 (N_46679,N_33412,N_34112);
nor U46680 (N_46680,N_34403,N_39187);
nand U46681 (N_46681,N_33269,N_35286);
nor U46682 (N_46682,N_36320,N_36550);
nor U46683 (N_46683,N_39918,N_36076);
nor U46684 (N_46684,N_35279,N_35446);
and U46685 (N_46685,N_34504,N_39646);
nor U46686 (N_46686,N_34620,N_30971);
nor U46687 (N_46687,N_33631,N_38527);
or U46688 (N_46688,N_39190,N_38065);
and U46689 (N_46689,N_35256,N_34399);
nor U46690 (N_46690,N_32838,N_30383);
nor U46691 (N_46691,N_35444,N_33529);
or U46692 (N_46692,N_38258,N_35583);
nand U46693 (N_46693,N_34206,N_36388);
or U46694 (N_46694,N_38547,N_37488);
nor U46695 (N_46695,N_31944,N_30555);
or U46696 (N_46696,N_34008,N_34268);
nand U46697 (N_46697,N_34703,N_33062);
xor U46698 (N_46698,N_36199,N_36233);
nand U46699 (N_46699,N_35575,N_37328);
nand U46700 (N_46700,N_32870,N_37133);
nor U46701 (N_46701,N_32188,N_35105);
and U46702 (N_46702,N_38732,N_39779);
or U46703 (N_46703,N_38424,N_36646);
nor U46704 (N_46704,N_38818,N_32503);
nand U46705 (N_46705,N_37254,N_38654);
nand U46706 (N_46706,N_37808,N_33689);
and U46707 (N_46707,N_33528,N_36596);
and U46708 (N_46708,N_33026,N_39186);
and U46709 (N_46709,N_31584,N_38549);
and U46710 (N_46710,N_35464,N_39783);
nor U46711 (N_46711,N_33988,N_30647);
nand U46712 (N_46712,N_35898,N_33097);
and U46713 (N_46713,N_30668,N_39406);
nand U46714 (N_46714,N_33742,N_33483);
and U46715 (N_46715,N_39129,N_35800);
or U46716 (N_46716,N_39715,N_32957);
nand U46717 (N_46717,N_37614,N_37873);
or U46718 (N_46718,N_32090,N_38078);
and U46719 (N_46719,N_33786,N_39153);
and U46720 (N_46720,N_32462,N_36785);
nand U46721 (N_46721,N_37356,N_32941);
and U46722 (N_46722,N_36462,N_35547);
nand U46723 (N_46723,N_30148,N_39941);
xnor U46724 (N_46724,N_34017,N_37502);
or U46725 (N_46725,N_38945,N_35413);
and U46726 (N_46726,N_30092,N_37406);
or U46727 (N_46727,N_37963,N_39344);
xor U46728 (N_46728,N_36218,N_37021);
and U46729 (N_46729,N_34494,N_35061);
and U46730 (N_46730,N_30477,N_31972);
nand U46731 (N_46731,N_34931,N_39211);
nand U46732 (N_46732,N_39545,N_32163);
or U46733 (N_46733,N_36334,N_31382);
xnor U46734 (N_46734,N_30968,N_31854);
nor U46735 (N_46735,N_35642,N_36588);
or U46736 (N_46736,N_39144,N_32961);
or U46737 (N_46737,N_39327,N_30544);
or U46738 (N_46738,N_35819,N_32211);
or U46739 (N_46739,N_31491,N_30829);
nand U46740 (N_46740,N_36256,N_31731);
xnor U46741 (N_46741,N_37564,N_38113);
xor U46742 (N_46742,N_36592,N_33376);
nand U46743 (N_46743,N_39830,N_32297);
nand U46744 (N_46744,N_33757,N_38757);
or U46745 (N_46745,N_39516,N_39701);
nor U46746 (N_46746,N_30427,N_38716);
and U46747 (N_46747,N_30885,N_35956);
and U46748 (N_46748,N_30597,N_34070);
xnor U46749 (N_46749,N_31060,N_33745);
xnor U46750 (N_46750,N_30372,N_31012);
or U46751 (N_46751,N_39856,N_35636);
and U46752 (N_46752,N_31348,N_38729);
and U46753 (N_46753,N_35938,N_37738);
and U46754 (N_46754,N_36622,N_36769);
or U46755 (N_46755,N_31078,N_34214);
and U46756 (N_46756,N_38819,N_36435);
nor U46757 (N_46757,N_39919,N_36023);
and U46758 (N_46758,N_38455,N_39465);
nor U46759 (N_46759,N_35530,N_30154);
and U46760 (N_46760,N_30220,N_36601);
or U46761 (N_46761,N_39290,N_32481);
and U46762 (N_46762,N_38247,N_36243);
nand U46763 (N_46763,N_37579,N_37933);
and U46764 (N_46764,N_38255,N_30940);
nor U46765 (N_46765,N_36338,N_39483);
xnor U46766 (N_46766,N_33734,N_34289);
nand U46767 (N_46767,N_38690,N_36399);
or U46768 (N_46768,N_33255,N_34328);
and U46769 (N_46769,N_35885,N_33812);
nand U46770 (N_46770,N_34601,N_35179);
nand U46771 (N_46771,N_31410,N_36822);
and U46772 (N_46772,N_39094,N_31474);
or U46773 (N_46773,N_39775,N_37068);
nand U46774 (N_46774,N_30701,N_30559);
nand U46775 (N_46775,N_31661,N_39018);
or U46776 (N_46776,N_35571,N_34928);
nor U46777 (N_46777,N_31282,N_33692);
nand U46778 (N_46778,N_31947,N_38081);
or U46779 (N_46779,N_37578,N_32865);
nand U46780 (N_46780,N_37014,N_37009);
and U46781 (N_46781,N_35517,N_30691);
or U46782 (N_46782,N_31330,N_32384);
nor U46783 (N_46783,N_35312,N_35645);
nand U46784 (N_46784,N_35973,N_39117);
and U46785 (N_46785,N_30906,N_32502);
and U46786 (N_46786,N_35238,N_38649);
nand U46787 (N_46787,N_31565,N_34434);
nand U46788 (N_46788,N_33793,N_32019);
and U46789 (N_46789,N_36612,N_36273);
and U46790 (N_46790,N_32354,N_30763);
and U46791 (N_46791,N_39712,N_32396);
xor U46792 (N_46792,N_36071,N_38102);
nand U46793 (N_46793,N_33511,N_35231);
nor U46794 (N_46794,N_38377,N_37469);
nand U46795 (N_46795,N_36825,N_33618);
or U46796 (N_46796,N_38375,N_33556);
and U46797 (N_46797,N_35461,N_37509);
or U46798 (N_46798,N_31779,N_30227);
nor U46799 (N_46799,N_39909,N_30746);
nor U46800 (N_46800,N_38868,N_37950);
or U46801 (N_46801,N_30610,N_33042);
nand U46802 (N_46802,N_36749,N_36847);
nor U46803 (N_46803,N_39805,N_38236);
or U46804 (N_46804,N_37449,N_39531);
or U46805 (N_46805,N_30845,N_36051);
xnor U46806 (N_46806,N_30701,N_35243);
nand U46807 (N_46807,N_32525,N_37373);
nor U46808 (N_46808,N_34857,N_32181);
and U46809 (N_46809,N_30357,N_39538);
nor U46810 (N_46810,N_35849,N_37137);
or U46811 (N_46811,N_31168,N_36724);
or U46812 (N_46812,N_33474,N_38280);
and U46813 (N_46813,N_33683,N_37275);
nor U46814 (N_46814,N_39092,N_32205);
or U46815 (N_46815,N_35182,N_30905);
nand U46816 (N_46816,N_31311,N_33274);
nor U46817 (N_46817,N_35899,N_35090);
nand U46818 (N_46818,N_34009,N_35904);
nor U46819 (N_46819,N_39484,N_39599);
nor U46820 (N_46820,N_37168,N_35415);
and U46821 (N_46821,N_33831,N_32813);
nor U46822 (N_46822,N_38741,N_36408);
and U46823 (N_46823,N_32108,N_35282);
nor U46824 (N_46824,N_31059,N_31962);
nand U46825 (N_46825,N_37264,N_37538);
or U46826 (N_46826,N_33378,N_39334);
nand U46827 (N_46827,N_36692,N_35182);
nand U46828 (N_46828,N_38510,N_36150);
nor U46829 (N_46829,N_36823,N_30060);
nand U46830 (N_46830,N_37391,N_39660);
and U46831 (N_46831,N_31007,N_30582);
nor U46832 (N_46832,N_30249,N_34934);
or U46833 (N_46833,N_37863,N_33178);
nand U46834 (N_46834,N_38714,N_32109);
or U46835 (N_46835,N_38977,N_32976);
nand U46836 (N_46836,N_31622,N_33837);
or U46837 (N_46837,N_32391,N_37141);
nand U46838 (N_46838,N_37383,N_35895);
nand U46839 (N_46839,N_37243,N_35407);
or U46840 (N_46840,N_32336,N_38126);
nor U46841 (N_46841,N_32129,N_39408);
or U46842 (N_46842,N_32785,N_31323);
xor U46843 (N_46843,N_32738,N_32759);
or U46844 (N_46844,N_39704,N_35323);
nand U46845 (N_46845,N_31218,N_38650);
xor U46846 (N_46846,N_39258,N_38298);
nor U46847 (N_46847,N_38206,N_36413);
nor U46848 (N_46848,N_30600,N_34464);
or U46849 (N_46849,N_39693,N_35707);
and U46850 (N_46850,N_38506,N_30809);
nor U46851 (N_46851,N_35859,N_34114);
and U46852 (N_46852,N_33440,N_36287);
and U46853 (N_46853,N_39369,N_39826);
xor U46854 (N_46854,N_39073,N_36711);
nor U46855 (N_46855,N_38853,N_33128);
nor U46856 (N_46856,N_37526,N_34674);
nor U46857 (N_46857,N_33744,N_35396);
or U46858 (N_46858,N_33726,N_32283);
nor U46859 (N_46859,N_32075,N_39231);
xor U46860 (N_46860,N_35539,N_37296);
or U46861 (N_46861,N_34848,N_38442);
and U46862 (N_46862,N_38490,N_30659);
or U46863 (N_46863,N_31917,N_33258);
nand U46864 (N_46864,N_36544,N_34413);
xnor U46865 (N_46865,N_39913,N_35989);
or U46866 (N_46866,N_35233,N_35275);
and U46867 (N_46867,N_30035,N_39418);
and U46868 (N_46868,N_32536,N_33892);
and U46869 (N_46869,N_37510,N_31315);
and U46870 (N_46870,N_31744,N_37629);
and U46871 (N_46871,N_35381,N_30844);
or U46872 (N_46872,N_30663,N_39302);
nand U46873 (N_46873,N_37042,N_39213);
nor U46874 (N_46874,N_34222,N_35426);
nor U46875 (N_46875,N_35405,N_38834);
or U46876 (N_46876,N_39535,N_39017);
nor U46877 (N_46877,N_33239,N_30841);
and U46878 (N_46878,N_39929,N_37601);
or U46879 (N_46879,N_36426,N_36481);
nand U46880 (N_46880,N_30800,N_32518);
or U46881 (N_46881,N_33665,N_33371);
or U46882 (N_46882,N_35093,N_39174);
nand U46883 (N_46883,N_33219,N_31674);
nor U46884 (N_46884,N_37709,N_35130);
nor U46885 (N_46885,N_37045,N_37916);
nand U46886 (N_46886,N_30700,N_34395);
nand U46887 (N_46887,N_35362,N_39594);
nand U46888 (N_46888,N_34042,N_34008);
nand U46889 (N_46889,N_33166,N_36437);
nand U46890 (N_46890,N_30308,N_35017);
nor U46891 (N_46891,N_35499,N_37396);
nor U46892 (N_46892,N_39459,N_31167);
nor U46893 (N_46893,N_31417,N_37494);
nor U46894 (N_46894,N_30447,N_35443);
and U46895 (N_46895,N_39625,N_35140);
nor U46896 (N_46896,N_33767,N_33431);
nand U46897 (N_46897,N_39314,N_38053);
and U46898 (N_46898,N_35399,N_30984);
nor U46899 (N_46899,N_34089,N_35196);
nand U46900 (N_46900,N_36310,N_32814);
or U46901 (N_46901,N_37341,N_37282);
nand U46902 (N_46902,N_31899,N_37816);
nand U46903 (N_46903,N_31308,N_34347);
nand U46904 (N_46904,N_36318,N_36001);
or U46905 (N_46905,N_31136,N_33059);
or U46906 (N_46906,N_35116,N_31005);
nand U46907 (N_46907,N_30462,N_32588);
nand U46908 (N_46908,N_30000,N_34239);
and U46909 (N_46909,N_39633,N_36188);
and U46910 (N_46910,N_32852,N_34281);
nor U46911 (N_46911,N_31542,N_34009);
xor U46912 (N_46912,N_37907,N_35336);
nor U46913 (N_46913,N_33980,N_35870);
nand U46914 (N_46914,N_38741,N_32703);
and U46915 (N_46915,N_36336,N_32186);
nor U46916 (N_46916,N_37214,N_32127);
xor U46917 (N_46917,N_33079,N_35664);
xnor U46918 (N_46918,N_39893,N_33700);
nor U46919 (N_46919,N_35285,N_36070);
nor U46920 (N_46920,N_39849,N_31493);
nor U46921 (N_46921,N_35144,N_37051);
nor U46922 (N_46922,N_30477,N_32321);
nand U46923 (N_46923,N_31741,N_31398);
and U46924 (N_46924,N_33270,N_32693);
or U46925 (N_46925,N_36404,N_34058);
nor U46926 (N_46926,N_33256,N_36595);
nand U46927 (N_46927,N_33677,N_39020);
and U46928 (N_46928,N_30301,N_30395);
xnor U46929 (N_46929,N_32544,N_30966);
nor U46930 (N_46930,N_35831,N_37463);
xor U46931 (N_46931,N_36012,N_30057);
and U46932 (N_46932,N_31745,N_33858);
and U46933 (N_46933,N_34383,N_32344);
or U46934 (N_46934,N_34940,N_39651);
nor U46935 (N_46935,N_30953,N_31702);
nor U46936 (N_46936,N_35769,N_33788);
and U46937 (N_46937,N_31446,N_33474);
nand U46938 (N_46938,N_30242,N_33990);
nor U46939 (N_46939,N_32472,N_35203);
and U46940 (N_46940,N_39707,N_39461);
nor U46941 (N_46941,N_31435,N_31624);
nor U46942 (N_46942,N_30424,N_39752);
xnor U46943 (N_46943,N_34137,N_33749);
nor U46944 (N_46944,N_34082,N_32407);
nor U46945 (N_46945,N_37572,N_36713);
nand U46946 (N_46946,N_32197,N_32190);
nand U46947 (N_46947,N_37988,N_36739);
and U46948 (N_46948,N_39970,N_32046);
nand U46949 (N_46949,N_34777,N_33271);
nand U46950 (N_46950,N_35927,N_38568);
or U46951 (N_46951,N_35420,N_33374);
nand U46952 (N_46952,N_38431,N_32365);
nand U46953 (N_46953,N_33901,N_34265);
or U46954 (N_46954,N_34016,N_38706);
or U46955 (N_46955,N_31419,N_35560);
xor U46956 (N_46956,N_37623,N_31352);
nor U46957 (N_46957,N_36401,N_36030);
nor U46958 (N_46958,N_37012,N_32430);
nor U46959 (N_46959,N_33142,N_37155);
and U46960 (N_46960,N_35513,N_32325);
and U46961 (N_46961,N_33776,N_30966);
and U46962 (N_46962,N_30122,N_34037);
and U46963 (N_46963,N_33889,N_33090);
or U46964 (N_46964,N_31916,N_32264);
or U46965 (N_46965,N_39839,N_31675);
or U46966 (N_46966,N_39880,N_39967);
xor U46967 (N_46967,N_32154,N_34585);
and U46968 (N_46968,N_37736,N_39092);
nand U46969 (N_46969,N_39723,N_34244);
and U46970 (N_46970,N_31239,N_36691);
nand U46971 (N_46971,N_33578,N_34584);
nor U46972 (N_46972,N_38978,N_34191);
nor U46973 (N_46973,N_37474,N_31690);
or U46974 (N_46974,N_38244,N_34129);
and U46975 (N_46975,N_36432,N_31101);
nor U46976 (N_46976,N_38693,N_32917);
or U46977 (N_46977,N_34037,N_32624);
and U46978 (N_46978,N_39157,N_35487);
nor U46979 (N_46979,N_38456,N_33342);
nor U46980 (N_46980,N_31897,N_30668);
or U46981 (N_46981,N_37157,N_34234);
nand U46982 (N_46982,N_39080,N_33468);
and U46983 (N_46983,N_34038,N_31150);
nor U46984 (N_46984,N_38594,N_35764);
and U46985 (N_46985,N_36535,N_36093);
or U46986 (N_46986,N_39959,N_33108);
nor U46987 (N_46987,N_39688,N_39489);
nor U46988 (N_46988,N_35637,N_33043);
and U46989 (N_46989,N_37671,N_39004);
xnor U46990 (N_46990,N_38068,N_34497);
nand U46991 (N_46991,N_35591,N_34025);
and U46992 (N_46992,N_32516,N_38739);
xor U46993 (N_46993,N_34533,N_30946);
nand U46994 (N_46994,N_32996,N_30435);
nand U46995 (N_46995,N_39770,N_36382);
nand U46996 (N_46996,N_35525,N_38570);
or U46997 (N_46997,N_32887,N_35635);
or U46998 (N_46998,N_36582,N_30673);
and U46999 (N_46999,N_37586,N_33821);
xor U47000 (N_47000,N_33370,N_37088);
nor U47001 (N_47001,N_37499,N_32975);
or U47002 (N_47002,N_35377,N_34579);
nor U47003 (N_47003,N_30389,N_36220);
and U47004 (N_47004,N_32737,N_36102);
nand U47005 (N_47005,N_31487,N_39291);
nand U47006 (N_47006,N_36586,N_31883);
nand U47007 (N_47007,N_39527,N_39142);
and U47008 (N_47008,N_36211,N_31517);
nor U47009 (N_47009,N_33344,N_32888);
nor U47010 (N_47010,N_38046,N_35933);
nor U47011 (N_47011,N_31732,N_36945);
nor U47012 (N_47012,N_39382,N_34031);
xnor U47013 (N_47013,N_39335,N_37250);
nor U47014 (N_47014,N_32713,N_39080);
and U47015 (N_47015,N_31323,N_33784);
or U47016 (N_47016,N_37760,N_35636);
or U47017 (N_47017,N_30358,N_30593);
and U47018 (N_47018,N_36192,N_31279);
nand U47019 (N_47019,N_30893,N_39361);
or U47020 (N_47020,N_39961,N_39525);
nor U47021 (N_47021,N_38621,N_37268);
nand U47022 (N_47022,N_32431,N_36368);
nor U47023 (N_47023,N_30149,N_30667);
or U47024 (N_47024,N_36688,N_36636);
or U47025 (N_47025,N_38740,N_35795);
nand U47026 (N_47026,N_34469,N_38477);
or U47027 (N_47027,N_31260,N_36974);
and U47028 (N_47028,N_33613,N_37477);
nand U47029 (N_47029,N_30313,N_32098);
xnor U47030 (N_47030,N_38697,N_34825);
nand U47031 (N_47031,N_39809,N_38370);
nand U47032 (N_47032,N_30435,N_32754);
xor U47033 (N_47033,N_39574,N_35876);
nand U47034 (N_47034,N_35136,N_31582);
nand U47035 (N_47035,N_38449,N_39370);
or U47036 (N_47036,N_36701,N_34451);
and U47037 (N_47037,N_38961,N_34579);
xor U47038 (N_47038,N_35554,N_37931);
nor U47039 (N_47039,N_32496,N_32481);
and U47040 (N_47040,N_38686,N_36247);
or U47041 (N_47041,N_33194,N_32596);
and U47042 (N_47042,N_36625,N_31138);
and U47043 (N_47043,N_34699,N_34122);
or U47044 (N_47044,N_35813,N_37939);
and U47045 (N_47045,N_31338,N_32010);
or U47046 (N_47046,N_31386,N_32650);
nor U47047 (N_47047,N_39541,N_38187);
and U47048 (N_47048,N_34593,N_31150);
nor U47049 (N_47049,N_37597,N_38832);
and U47050 (N_47050,N_30593,N_35725);
nand U47051 (N_47051,N_31896,N_33699);
and U47052 (N_47052,N_38604,N_34365);
or U47053 (N_47053,N_35459,N_32705);
or U47054 (N_47054,N_37378,N_34475);
nor U47055 (N_47055,N_34155,N_35972);
or U47056 (N_47056,N_30235,N_31364);
and U47057 (N_47057,N_33052,N_32734);
or U47058 (N_47058,N_32851,N_35479);
nor U47059 (N_47059,N_32333,N_32392);
and U47060 (N_47060,N_34879,N_31902);
nand U47061 (N_47061,N_38438,N_31717);
and U47062 (N_47062,N_39043,N_36014);
or U47063 (N_47063,N_38976,N_36253);
or U47064 (N_47064,N_34464,N_31321);
or U47065 (N_47065,N_33335,N_33145);
or U47066 (N_47066,N_37406,N_39525);
xnor U47067 (N_47067,N_35114,N_34071);
xnor U47068 (N_47068,N_33281,N_30965);
nand U47069 (N_47069,N_38823,N_34363);
xnor U47070 (N_47070,N_35048,N_32400);
and U47071 (N_47071,N_37514,N_39536);
or U47072 (N_47072,N_35217,N_36580);
nor U47073 (N_47073,N_39046,N_32088);
nand U47074 (N_47074,N_31124,N_32525);
nor U47075 (N_47075,N_36228,N_32184);
and U47076 (N_47076,N_38511,N_30030);
and U47077 (N_47077,N_31779,N_36362);
nand U47078 (N_47078,N_37813,N_38294);
nor U47079 (N_47079,N_34969,N_33637);
or U47080 (N_47080,N_35772,N_34198);
nor U47081 (N_47081,N_36773,N_37360);
nor U47082 (N_47082,N_30076,N_35683);
nor U47083 (N_47083,N_31948,N_35056);
nor U47084 (N_47084,N_38016,N_30277);
and U47085 (N_47085,N_39630,N_31908);
nand U47086 (N_47086,N_31743,N_32872);
and U47087 (N_47087,N_37205,N_38416);
nor U47088 (N_47088,N_32988,N_31574);
nor U47089 (N_47089,N_39414,N_37104);
nor U47090 (N_47090,N_38562,N_37295);
or U47091 (N_47091,N_38920,N_30487);
and U47092 (N_47092,N_39500,N_35457);
xnor U47093 (N_47093,N_36064,N_37855);
nor U47094 (N_47094,N_32564,N_35952);
nand U47095 (N_47095,N_35553,N_37913);
and U47096 (N_47096,N_36457,N_31274);
and U47097 (N_47097,N_33164,N_34656);
and U47098 (N_47098,N_33668,N_38840);
nor U47099 (N_47099,N_35014,N_39796);
and U47100 (N_47100,N_38304,N_32179);
and U47101 (N_47101,N_39872,N_31167);
nor U47102 (N_47102,N_37828,N_30238);
and U47103 (N_47103,N_38096,N_33951);
and U47104 (N_47104,N_35923,N_32592);
nor U47105 (N_47105,N_32304,N_35827);
xnor U47106 (N_47106,N_38254,N_36108);
nand U47107 (N_47107,N_30477,N_39125);
or U47108 (N_47108,N_32441,N_37687);
nor U47109 (N_47109,N_39943,N_30208);
nand U47110 (N_47110,N_35567,N_36950);
nor U47111 (N_47111,N_37870,N_34970);
nand U47112 (N_47112,N_38314,N_30100);
xor U47113 (N_47113,N_39589,N_30829);
nand U47114 (N_47114,N_33122,N_31434);
xor U47115 (N_47115,N_35872,N_30275);
nand U47116 (N_47116,N_38790,N_38504);
nand U47117 (N_47117,N_31181,N_36797);
nand U47118 (N_47118,N_33666,N_35712);
nor U47119 (N_47119,N_34451,N_35372);
nor U47120 (N_47120,N_34945,N_39058);
or U47121 (N_47121,N_36839,N_33222);
nand U47122 (N_47122,N_38218,N_36573);
nand U47123 (N_47123,N_37505,N_38501);
nand U47124 (N_47124,N_33646,N_30550);
and U47125 (N_47125,N_39656,N_31059);
nand U47126 (N_47126,N_37859,N_35467);
and U47127 (N_47127,N_33684,N_30186);
and U47128 (N_47128,N_38184,N_33302);
and U47129 (N_47129,N_30612,N_30242);
or U47130 (N_47130,N_39228,N_34034);
xnor U47131 (N_47131,N_37451,N_32774);
and U47132 (N_47132,N_39414,N_39117);
and U47133 (N_47133,N_30766,N_39308);
nor U47134 (N_47134,N_39369,N_31965);
nand U47135 (N_47135,N_30781,N_35129);
or U47136 (N_47136,N_31125,N_33641);
nor U47137 (N_47137,N_39703,N_30965);
nor U47138 (N_47138,N_36418,N_39852);
nand U47139 (N_47139,N_31636,N_36290);
or U47140 (N_47140,N_33368,N_37271);
or U47141 (N_47141,N_38666,N_32210);
nor U47142 (N_47142,N_36595,N_34622);
nor U47143 (N_47143,N_33039,N_31612);
or U47144 (N_47144,N_30388,N_32838);
nor U47145 (N_47145,N_31809,N_35711);
nand U47146 (N_47146,N_38793,N_34788);
or U47147 (N_47147,N_33738,N_38616);
nor U47148 (N_47148,N_31141,N_30511);
nor U47149 (N_47149,N_31795,N_34685);
and U47150 (N_47150,N_33106,N_33658);
nor U47151 (N_47151,N_32567,N_33959);
and U47152 (N_47152,N_30228,N_32934);
nand U47153 (N_47153,N_31229,N_32048);
or U47154 (N_47154,N_37192,N_31029);
and U47155 (N_47155,N_34782,N_30048);
nor U47156 (N_47156,N_30857,N_39642);
or U47157 (N_47157,N_30401,N_31855);
and U47158 (N_47158,N_38268,N_36736);
xor U47159 (N_47159,N_37841,N_36080);
nand U47160 (N_47160,N_32540,N_36807);
nor U47161 (N_47161,N_30204,N_36711);
nand U47162 (N_47162,N_39659,N_37759);
nor U47163 (N_47163,N_39020,N_39881);
nor U47164 (N_47164,N_35468,N_34631);
or U47165 (N_47165,N_39408,N_38572);
nand U47166 (N_47166,N_33620,N_37145);
nand U47167 (N_47167,N_34280,N_31947);
or U47168 (N_47168,N_38364,N_38134);
nor U47169 (N_47169,N_33044,N_31595);
xnor U47170 (N_47170,N_39850,N_37405);
nor U47171 (N_47171,N_31839,N_38182);
and U47172 (N_47172,N_31344,N_32413);
nor U47173 (N_47173,N_35009,N_32995);
nor U47174 (N_47174,N_39332,N_35000);
nand U47175 (N_47175,N_30405,N_31623);
or U47176 (N_47176,N_35464,N_32959);
or U47177 (N_47177,N_30430,N_33075);
or U47178 (N_47178,N_31081,N_32104);
and U47179 (N_47179,N_37818,N_32075);
nand U47180 (N_47180,N_37500,N_37021);
nor U47181 (N_47181,N_34972,N_37354);
nor U47182 (N_47182,N_36289,N_39478);
nor U47183 (N_47183,N_31229,N_36304);
or U47184 (N_47184,N_32557,N_35118);
and U47185 (N_47185,N_37326,N_32265);
nor U47186 (N_47186,N_34329,N_37280);
nand U47187 (N_47187,N_30210,N_35418);
nand U47188 (N_47188,N_37117,N_38786);
or U47189 (N_47189,N_32617,N_33100);
nor U47190 (N_47190,N_38601,N_33901);
nand U47191 (N_47191,N_35732,N_31563);
nand U47192 (N_47192,N_37842,N_38770);
and U47193 (N_47193,N_35265,N_38234);
nor U47194 (N_47194,N_32950,N_34660);
or U47195 (N_47195,N_36644,N_37955);
and U47196 (N_47196,N_39915,N_32543);
nand U47197 (N_47197,N_37778,N_31382);
nand U47198 (N_47198,N_31204,N_31683);
xnor U47199 (N_47199,N_35880,N_34624);
xor U47200 (N_47200,N_37445,N_34260);
nand U47201 (N_47201,N_34493,N_36293);
nand U47202 (N_47202,N_30493,N_39009);
nor U47203 (N_47203,N_30197,N_34608);
nor U47204 (N_47204,N_34166,N_37500);
nand U47205 (N_47205,N_34200,N_35033);
nor U47206 (N_47206,N_33690,N_35970);
nand U47207 (N_47207,N_33618,N_30681);
nor U47208 (N_47208,N_37221,N_35068);
or U47209 (N_47209,N_37018,N_37183);
nor U47210 (N_47210,N_37302,N_38276);
nor U47211 (N_47211,N_39210,N_38503);
nor U47212 (N_47212,N_37722,N_33273);
nand U47213 (N_47213,N_38519,N_38809);
nand U47214 (N_47214,N_32347,N_36498);
and U47215 (N_47215,N_37642,N_34414);
nor U47216 (N_47216,N_33202,N_32349);
nand U47217 (N_47217,N_39396,N_35380);
nor U47218 (N_47218,N_31965,N_31505);
nor U47219 (N_47219,N_37154,N_36840);
or U47220 (N_47220,N_32459,N_33532);
or U47221 (N_47221,N_34572,N_35867);
or U47222 (N_47222,N_35708,N_32193);
nor U47223 (N_47223,N_30128,N_37670);
nand U47224 (N_47224,N_32716,N_32035);
and U47225 (N_47225,N_39522,N_31672);
and U47226 (N_47226,N_32431,N_39019);
nand U47227 (N_47227,N_36324,N_36448);
nor U47228 (N_47228,N_31683,N_38741);
and U47229 (N_47229,N_34828,N_35027);
and U47230 (N_47230,N_30417,N_36203);
and U47231 (N_47231,N_37223,N_32538);
or U47232 (N_47232,N_36988,N_38952);
and U47233 (N_47233,N_33734,N_39099);
and U47234 (N_47234,N_34607,N_30993);
and U47235 (N_47235,N_36179,N_39401);
or U47236 (N_47236,N_36503,N_31340);
nand U47237 (N_47237,N_33056,N_36285);
nor U47238 (N_47238,N_34918,N_31469);
or U47239 (N_47239,N_36129,N_36132);
and U47240 (N_47240,N_39978,N_32292);
or U47241 (N_47241,N_35772,N_33336);
xnor U47242 (N_47242,N_36563,N_38032);
or U47243 (N_47243,N_36522,N_35247);
or U47244 (N_47244,N_30832,N_39716);
nand U47245 (N_47245,N_39795,N_33520);
or U47246 (N_47246,N_37230,N_35318);
nand U47247 (N_47247,N_39474,N_30655);
and U47248 (N_47248,N_38903,N_30378);
xnor U47249 (N_47249,N_35885,N_39092);
nand U47250 (N_47250,N_31203,N_30211);
or U47251 (N_47251,N_38098,N_31607);
nand U47252 (N_47252,N_30962,N_34169);
or U47253 (N_47253,N_38373,N_39282);
or U47254 (N_47254,N_35085,N_34702);
and U47255 (N_47255,N_38514,N_32917);
xnor U47256 (N_47256,N_38032,N_34642);
nor U47257 (N_47257,N_34236,N_34151);
and U47258 (N_47258,N_33315,N_32126);
or U47259 (N_47259,N_31905,N_31906);
or U47260 (N_47260,N_30606,N_33182);
and U47261 (N_47261,N_32089,N_31575);
nor U47262 (N_47262,N_37973,N_39425);
or U47263 (N_47263,N_38892,N_32270);
and U47264 (N_47264,N_37336,N_39080);
or U47265 (N_47265,N_31567,N_34444);
nand U47266 (N_47266,N_33046,N_38589);
or U47267 (N_47267,N_30116,N_30891);
nor U47268 (N_47268,N_35291,N_32163);
nor U47269 (N_47269,N_31463,N_36091);
nand U47270 (N_47270,N_30625,N_38305);
nor U47271 (N_47271,N_35338,N_31974);
and U47272 (N_47272,N_30314,N_35649);
nor U47273 (N_47273,N_30972,N_31609);
or U47274 (N_47274,N_33980,N_33564);
and U47275 (N_47275,N_39884,N_31586);
nor U47276 (N_47276,N_37532,N_36661);
and U47277 (N_47277,N_34408,N_35214);
xor U47278 (N_47278,N_33218,N_30531);
xnor U47279 (N_47279,N_32358,N_30703);
and U47280 (N_47280,N_37482,N_35112);
or U47281 (N_47281,N_31524,N_31741);
nor U47282 (N_47282,N_37918,N_36996);
nor U47283 (N_47283,N_37767,N_33941);
or U47284 (N_47284,N_37020,N_31292);
xnor U47285 (N_47285,N_34105,N_38612);
nor U47286 (N_47286,N_36033,N_38754);
xnor U47287 (N_47287,N_33948,N_35195);
nand U47288 (N_47288,N_36699,N_39465);
and U47289 (N_47289,N_30163,N_32564);
or U47290 (N_47290,N_31022,N_36942);
and U47291 (N_47291,N_35627,N_32894);
nor U47292 (N_47292,N_38572,N_32711);
xnor U47293 (N_47293,N_32291,N_36178);
nand U47294 (N_47294,N_35106,N_39906);
nor U47295 (N_47295,N_30051,N_39325);
or U47296 (N_47296,N_35011,N_39008);
nor U47297 (N_47297,N_38651,N_32662);
or U47298 (N_47298,N_35793,N_34973);
xnor U47299 (N_47299,N_35592,N_39192);
nand U47300 (N_47300,N_33008,N_34691);
and U47301 (N_47301,N_35311,N_31326);
xor U47302 (N_47302,N_32527,N_39265);
nor U47303 (N_47303,N_39882,N_30453);
or U47304 (N_47304,N_36529,N_36780);
or U47305 (N_47305,N_32160,N_37384);
nand U47306 (N_47306,N_36629,N_38536);
or U47307 (N_47307,N_38635,N_39191);
nand U47308 (N_47308,N_39526,N_33301);
and U47309 (N_47309,N_32087,N_36808);
nor U47310 (N_47310,N_31631,N_38807);
or U47311 (N_47311,N_38255,N_32507);
nor U47312 (N_47312,N_33176,N_34588);
and U47313 (N_47313,N_38824,N_39895);
or U47314 (N_47314,N_37950,N_35559);
nor U47315 (N_47315,N_39137,N_30878);
nand U47316 (N_47316,N_36359,N_34257);
nor U47317 (N_47317,N_31087,N_31590);
or U47318 (N_47318,N_38372,N_34556);
nor U47319 (N_47319,N_31605,N_37697);
nand U47320 (N_47320,N_35058,N_33489);
and U47321 (N_47321,N_35628,N_30439);
xnor U47322 (N_47322,N_30864,N_33483);
nor U47323 (N_47323,N_36379,N_36217);
nor U47324 (N_47324,N_33945,N_30403);
nor U47325 (N_47325,N_34171,N_31613);
nor U47326 (N_47326,N_33846,N_31611);
and U47327 (N_47327,N_33152,N_39424);
or U47328 (N_47328,N_39554,N_30564);
nand U47329 (N_47329,N_39866,N_33290);
xor U47330 (N_47330,N_34528,N_38809);
xor U47331 (N_47331,N_31552,N_38228);
and U47332 (N_47332,N_36207,N_33815);
or U47333 (N_47333,N_35122,N_31860);
nand U47334 (N_47334,N_36427,N_38785);
and U47335 (N_47335,N_30248,N_39772);
nand U47336 (N_47336,N_35541,N_38257);
xnor U47337 (N_47337,N_32723,N_37321);
and U47338 (N_47338,N_39441,N_33811);
nand U47339 (N_47339,N_38070,N_39448);
or U47340 (N_47340,N_37359,N_37091);
nand U47341 (N_47341,N_35250,N_36165);
or U47342 (N_47342,N_36219,N_31547);
and U47343 (N_47343,N_31292,N_33513);
nor U47344 (N_47344,N_30226,N_39110);
and U47345 (N_47345,N_35022,N_39669);
nor U47346 (N_47346,N_31300,N_33733);
or U47347 (N_47347,N_30307,N_35156);
nor U47348 (N_47348,N_32017,N_35898);
or U47349 (N_47349,N_37993,N_32065);
or U47350 (N_47350,N_34384,N_30740);
xnor U47351 (N_47351,N_33720,N_37615);
or U47352 (N_47352,N_30224,N_31842);
nor U47353 (N_47353,N_34295,N_38782);
xnor U47354 (N_47354,N_39517,N_33251);
or U47355 (N_47355,N_36546,N_35149);
or U47356 (N_47356,N_30873,N_38180);
nor U47357 (N_47357,N_32531,N_38718);
nand U47358 (N_47358,N_30752,N_37676);
nor U47359 (N_47359,N_36778,N_39133);
nor U47360 (N_47360,N_36897,N_32788);
and U47361 (N_47361,N_34824,N_39015);
xor U47362 (N_47362,N_34662,N_30588);
or U47363 (N_47363,N_34549,N_33677);
nor U47364 (N_47364,N_37586,N_38051);
nand U47365 (N_47365,N_30046,N_32924);
or U47366 (N_47366,N_36030,N_31873);
nor U47367 (N_47367,N_35105,N_39724);
nor U47368 (N_47368,N_39984,N_34314);
nand U47369 (N_47369,N_31496,N_39739);
xnor U47370 (N_47370,N_37886,N_39816);
xor U47371 (N_47371,N_34571,N_35222);
nand U47372 (N_47372,N_32472,N_31741);
or U47373 (N_47373,N_33915,N_32336);
and U47374 (N_47374,N_31031,N_36191);
nand U47375 (N_47375,N_30760,N_33188);
nor U47376 (N_47376,N_30372,N_33229);
nand U47377 (N_47377,N_36246,N_32828);
nand U47378 (N_47378,N_36075,N_30163);
nand U47379 (N_47379,N_34041,N_31082);
and U47380 (N_47380,N_34307,N_35049);
nand U47381 (N_47381,N_30036,N_37558);
and U47382 (N_47382,N_37467,N_39781);
or U47383 (N_47383,N_31577,N_31899);
nand U47384 (N_47384,N_36663,N_32168);
nor U47385 (N_47385,N_36469,N_30243);
and U47386 (N_47386,N_39191,N_30272);
nor U47387 (N_47387,N_35376,N_38889);
and U47388 (N_47388,N_36318,N_35744);
nand U47389 (N_47389,N_31005,N_39524);
and U47390 (N_47390,N_37601,N_31810);
nor U47391 (N_47391,N_30769,N_32809);
and U47392 (N_47392,N_32552,N_30173);
nand U47393 (N_47393,N_31562,N_37683);
and U47394 (N_47394,N_30677,N_39996);
and U47395 (N_47395,N_33869,N_31914);
and U47396 (N_47396,N_37773,N_39430);
or U47397 (N_47397,N_38215,N_35610);
and U47398 (N_47398,N_34480,N_32109);
nor U47399 (N_47399,N_37159,N_38090);
nand U47400 (N_47400,N_37219,N_34242);
nor U47401 (N_47401,N_35084,N_36271);
nor U47402 (N_47402,N_33159,N_36043);
nand U47403 (N_47403,N_32469,N_33655);
or U47404 (N_47404,N_37034,N_31340);
nor U47405 (N_47405,N_31879,N_31693);
nor U47406 (N_47406,N_36250,N_31340);
nor U47407 (N_47407,N_38472,N_30315);
and U47408 (N_47408,N_36926,N_32246);
nor U47409 (N_47409,N_35141,N_33854);
and U47410 (N_47410,N_32283,N_32849);
nand U47411 (N_47411,N_30952,N_31130);
and U47412 (N_47412,N_37955,N_38994);
nor U47413 (N_47413,N_36243,N_34254);
nor U47414 (N_47414,N_37902,N_32099);
or U47415 (N_47415,N_35021,N_38347);
nor U47416 (N_47416,N_39653,N_36765);
xor U47417 (N_47417,N_38410,N_33957);
nand U47418 (N_47418,N_39527,N_36015);
nor U47419 (N_47419,N_31470,N_38004);
nor U47420 (N_47420,N_32921,N_37289);
and U47421 (N_47421,N_38425,N_36241);
nor U47422 (N_47422,N_38202,N_35051);
and U47423 (N_47423,N_36984,N_36897);
and U47424 (N_47424,N_32895,N_32455);
and U47425 (N_47425,N_34184,N_32581);
or U47426 (N_47426,N_38725,N_36930);
nor U47427 (N_47427,N_34177,N_33709);
nand U47428 (N_47428,N_30881,N_36217);
xor U47429 (N_47429,N_38960,N_33288);
xor U47430 (N_47430,N_32741,N_37565);
nor U47431 (N_47431,N_37672,N_31038);
nand U47432 (N_47432,N_37683,N_31714);
and U47433 (N_47433,N_36072,N_33157);
or U47434 (N_47434,N_32136,N_37790);
nand U47435 (N_47435,N_36463,N_33379);
and U47436 (N_47436,N_35095,N_32197);
and U47437 (N_47437,N_30446,N_37255);
nand U47438 (N_47438,N_30919,N_39200);
and U47439 (N_47439,N_38111,N_34766);
xnor U47440 (N_47440,N_36506,N_39858);
nor U47441 (N_47441,N_37830,N_31514);
nand U47442 (N_47442,N_33541,N_35701);
nand U47443 (N_47443,N_35749,N_36297);
or U47444 (N_47444,N_36642,N_35440);
xor U47445 (N_47445,N_37621,N_30974);
nor U47446 (N_47446,N_32128,N_36762);
nor U47447 (N_47447,N_39923,N_35996);
nor U47448 (N_47448,N_39911,N_35618);
nand U47449 (N_47449,N_36666,N_37650);
xnor U47450 (N_47450,N_37487,N_35678);
and U47451 (N_47451,N_36635,N_38144);
nand U47452 (N_47452,N_34536,N_32622);
and U47453 (N_47453,N_39715,N_39416);
nand U47454 (N_47454,N_37668,N_37632);
xor U47455 (N_47455,N_36646,N_32588);
nor U47456 (N_47456,N_39801,N_34213);
nand U47457 (N_47457,N_33480,N_37267);
nor U47458 (N_47458,N_30302,N_31064);
nor U47459 (N_47459,N_30634,N_39665);
or U47460 (N_47460,N_37987,N_36890);
nor U47461 (N_47461,N_34011,N_30344);
nand U47462 (N_47462,N_30076,N_36036);
xnor U47463 (N_47463,N_37992,N_32592);
nand U47464 (N_47464,N_34402,N_30085);
nor U47465 (N_47465,N_30122,N_34749);
nor U47466 (N_47466,N_31403,N_33250);
or U47467 (N_47467,N_39337,N_35762);
and U47468 (N_47468,N_30320,N_38201);
or U47469 (N_47469,N_35664,N_34068);
xnor U47470 (N_47470,N_30973,N_38725);
or U47471 (N_47471,N_37505,N_32120);
nor U47472 (N_47472,N_39127,N_39956);
and U47473 (N_47473,N_36678,N_33479);
nand U47474 (N_47474,N_31810,N_35612);
and U47475 (N_47475,N_33115,N_31245);
nand U47476 (N_47476,N_39339,N_32628);
nand U47477 (N_47477,N_35499,N_32064);
and U47478 (N_47478,N_35853,N_39586);
or U47479 (N_47479,N_37780,N_32557);
nand U47480 (N_47480,N_34435,N_33231);
nand U47481 (N_47481,N_36179,N_31967);
or U47482 (N_47482,N_33043,N_30289);
nand U47483 (N_47483,N_38244,N_33194);
nor U47484 (N_47484,N_37420,N_37540);
and U47485 (N_47485,N_31681,N_35210);
and U47486 (N_47486,N_33310,N_34713);
nor U47487 (N_47487,N_30638,N_38110);
xor U47488 (N_47488,N_31104,N_38506);
and U47489 (N_47489,N_30921,N_34728);
nor U47490 (N_47490,N_34698,N_30372);
or U47491 (N_47491,N_36515,N_34210);
nand U47492 (N_47492,N_35527,N_31165);
and U47493 (N_47493,N_37188,N_39547);
nor U47494 (N_47494,N_39442,N_31873);
and U47495 (N_47495,N_36992,N_38133);
and U47496 (N_47496,N_31942,N_39921);
nand U47497 (N_47497,N_39308,N_31744);
or U47498 (N_47498,N_36241,N_38802);
nand U47499 (N_47499,N_32872,N_38897);
and U47500 (N_47500,N_35893,N_34269);
nor U47501 (N_47501,N_32245,N_33557);
or U47502 (N_47502,N_32275,N_34076);
nor U47503 (N_47503,N_31708,N_37502);
nand U47504 (N_47504,N_32266,N_37738);
nand U47505 (N_47505,N_33947,N_38283);
nor U47506 (N_47506,N_39992,N_39958);
nor U47507 (N_47507,N_35348,N_35142);
nor U47508 (N_47508,N_32787,N_32933);
nor U47509 (N_47509,N_30612,N_38627);
nor U47510 (N_47510,N_31789,N_37891);
and U47511 (N_47511,N_32408,N_30777);
or U47512 (N_47512,N_38660,N_36246);
nand U47513 (N_47513,N_31739,N_39896);
or U47514 (N_47514,N_36847,N_36892);
nand U47515 (N_47515,N_39361,N_35222);
nand U47516 (N_47516,N_30747,N_31855);
nor U47517 (N_47517,N_38100,N_35637);
nor U47518 (N_47518,N_37808,N_33016);
or U47519 (N_47519,N_33316,N_30115);
xor U47520 (N_47520,N_30967,N_36865);
or U47521 (N_47521,N_35778,N_36894);
or U47522 (N_47522,N_39607,N_35414);
nor U47523 (N_47523,N_32099,N_36299);
and U47524 (N_47524,N_39153,N_31563);
or U47525 (N_47525,N_35357,N_33307);
or U47526 (N_47526,N_39782,N_32124);
nand U47527 (N_47527,N_32082,N_33568);
nand U47528 (N_47528,N_31353,N_35696);
and U47529 (N_47529,N_33115,N_30693);
nand U47530 (N_47530,N_33412,N_30067);
nand U47531 (N_47531,N_33387,N_30180);
nor U47532 (N_47532,N_38864,N_32441);
or U47533 (N_47533,N_38783,N_35256);
nor U47534 (N_47534,N_32524,N_39393);
and U47535 (N_47535,N_36414,N_33270);
and U47536 (N_47536,N_30951,N_36483);
and U47537 (N_47537,N_34636,N_37419);
and U47538 (N_47538,N_32617,N_38732);
nand U47539 (N_47539,N_39949,N_34229);
and U47540 (N_47540,N_34739,N_38344);
or U47541 (N_47541,N_37889,N_35929);
nor U47542 (N_47542,N_34042,N_37045);
and U47543 (N_47543,N_34861,N_32097);
nand U47544 (N_47544,N_31796,N_36397);
or U47545 (N_47545,N_32315,N_34640);
nand U47546 (N_47546,N_34008,N_38075);
nand U47547 (N_47547,N_36886,N_39774);
xnor U47548 (N_47548,N_35684,N_30770);
and U47549 (N_47549,N_32547,N_38252);
nand U47550 (N_47550,N_35199,N_39913);
nand U47551 (N_47551,N_31840,N_30949);
or U47552 (N_47552,N_30137,N_31623);
and U47553 (N_47553,N_30794,N_36849);
nor U47554 (N_47554,N_33940,N_32039);
or U47555 (N_47555,N_31929,N_32392);
nor U47556 (N_47556,N_33268,N_35984);
nor U47557 (N_47557,N_32181,N_39184);
and U47558 (N_47558,N_35460,N_36515);
nor U47559 (N_47559,N_34749,N_36554);
or U47560 (N_47560,N_30851,N_33811);
and U47561 (N_47561,N_39346,N_35966);
or U47562 (N_47562,N_36023,N_31139);
and U47563 (N_47563,N_36150,N_36990);
nor U47564 (N_47564,N_39128,N_32831);
xnor U47565 (N_47565,N_32541,N_30614);
nor U47566 (N_47566,N_33386,N_39734);
nor U47567 (N_47567,N_31343,N_38944);
nand U47568 (N_47568,N_34603,N_36911);
and U47569 (N_47569,N_37380,N_30764);
nand U47570 (N_47570,N_31855,N_34328);
nor U47571 (N_47571,N_32366,N_31719);
nor U47572 (N_47572,N_33507,N_35601);
or U47573 (N_47573,N_35019,N_34663);
nor U47574 (N_47574,N_34366,N_33031);
or U47575 (N_47575,N_36507,N_34030);
nand U47576 (N_47576,N_38597,N_36651);
xor U47577 (N_47577,N_34158,N_31700);
or U47578 (N_47578,N_38142,N_34034);
nand U47579 (N_47579,N_39509,N_31060);
xnor U47580 (N_47580,N_39206,N_39793);
and U47581 (N_47581,N_36634,N_32317);
xor U47582 (N_47582,N_37518,N_39236);
and U47583 (N_47583,N_30506,N_31066);
or U47584 (N_47584,N_31970,N_30739);
and U47585 (N_47585,N_38702,N_38390);
nand U47586 (N_47586,N_36828,N_35042);
or U47587 (N_47587,N_39255,N_32760);
and U47588 (N_47588,N_37133,N_39808);
or U47589 (N_47589,N_33772,N_32734);
and U47590 (N_47590,N_31586,N_34242);
and U47591 (N_47591,N_37083,N_37013);
or U47592 (N_47592,N_38785,N_36905);
nand U47593 (N_47593,N_39499,N_32788);
or U47594 (N_47594,N_32493,N_37791);
and U47595 (N_47595,N_36270,N_35178);
nor U47596 (N_47596,N_34155,N_39845);
and U47597 (N_47597,N_32397,N_34314);
xnor U47598 (N_47598,N_31302,N_36032);
or U47599 (N_47599,N_36904,N_36434);
or U47600 (N_47600,N_38671,N_38949);
and U47601 (N_47601,N_35412,N_37354);
or U47602 (N_47602,N_35994,N_33822);
nand U47603 (N_47603,N_31897,N_35872);
nor U47604 (N_47604,N_35991,N_36641);
or U47605 (N_47605,N_34530,N_36666);
xnor U47606 (N_47606,N_36042,N_35775);
nor U47607 (N_47607,N_31045,N_37737);
nand U47608 (N_47608,N_31656,N_37903);
nand U47609 (N_47609,N_39709,N_33629);
nand U47610 (N_47610,N_32004,N_32302);
nand U47611 (N_47611,N_31809,N_35342);
nand U47612 (N_47612,N_30270,N_31173);
nand U47613 (N_47613,N_31551,N_35705);
or U47614 (N_47614,N_35029,N_37960);
or U47615 (N_47615,N_32643,N_38592);
nand U47616 (N_47616,N_39283,N_34031);
or U47617 (N_47617,N_34650,N_37854);
nand U47618 (N_47618,N_39733,N_31703);
nand U47619 (N_47619,N_30270,N_35904);
and U47620 (N_47620,N_32874,N_37037);
or U47621 (N_47621,N_33527,N_31381);
nor U47622 (N_47622,N_36277,N_34972);
nand U47623 (N_47623,N_38720,N_32213);
and U47624 (N_47624,N_32100,N_38301);
nor U47625 (N_47625,N_32920,N_32444);
nor U47626 (N_47626,N_38687,N_35161);
nand U47627 (N_47627,N_36519,N_35758);
xnor U47628 (N_47628,N_34303,N_37030);
and U47629 (N_47629,N_38218,N_30979);
xnor U47630 (N_47630,N_32739,N_37993);
nand U47631 (N_47631,N_34587,N_35354);
and U47632 (N_47632,N_37775,N_30205);
nand U47633 (N_47633,N_38881,N_30493);
and U47634 (N_47634,N_33440,N_35457);
nor U47635 (N_47635,N_32957,N_38578);
nand U47636 (N_47636,N_32484,N_36245);
xor U47637 (N_47637,N_32107,N_33477);
nand U47638 (N_47638,N_31193,N_35760);
nor U47639 (N_47639,N_32843,N_30477);
xor U47640 (N_47640,N_33268,N_31675);
nand U47641 (N_47641,N_39955,N_32237);
or U47642 (N_47642,N_39891,N_36220);
nor U47643 (N_47643,N_30431,N_34061);
nor U47644 (N_47644,N_35984,N_31479);
nand U47645 (N_47645,N_39599,N_37243);
or U47646 (N_47646,N_35845,N_30513);
nor U47647 (N_47647,N_33719,N_37063);
or U47648 (N_47648,N_30323,N_34545);
nor U47649 (N_47649,N_35970,N_38963);
or U47650 (N_47650,N_33719,N_33868);
xor U47651 (N_47651,N_33453,N_36228);
or U47652 (N_47652,N_30680,N_38814);
or U47653 (N_47653,N_30130,N_33145);
nand U47654 (N_47654,N_35434,N_30948);
nor U47655 (N_47655,N_34930,N_34201);
xor U47656 (N_47656,N_32139,N_37958);
nor U47657 (N_47657,N_39606,N_34685);
and U47658 (N_47658,N_34774,N_35262);
or U47659 (N_47659,N_34929,N_37400);
xnor U47660 (N_47660,N_34726,N_32410);
and U47661 (N_47661,N_33735,N_34801);
xnor U47662 (N_47662,N_36574,N_37466);
nor U47663 (N_47663,N_39965,N_37020);
and U47664 (N_47664,N_39919,N_34526);
nand U47665 (N_47665,N_39226,N_36523);
or U47666 (N_47666,N_32757,N_38073);
nand U47667 (N_47667,N_39187,N_34348);
nand U47668 (N_47668,N_36613,N_39503);
and U47669 (N_47669,N_33560,N_30373);
or U47670 (N_47670,N_36396,N_38747);
and U47671 (N_47671,N_32020,N_39057);
and U47672 (N_47672,N_30049,N_36187);
nor U47673 (N_47673,N_32020,N_32833);
or U47674 (N_47674,N_30204,N_36264);
and U47675 (N_47675,N_30589,N_39890);
or U47676 (N_47676,N_39214,N_36581);
or U47677 (N_47677,N_38117,N_34073);
and U47678 (N_47678,N_39318,N_31672);
and U47679 (N_47679,N_32762,N_33460);
and U47680 (N_47680,N_30896,N_32353);
nand U47681 (N_47681,N_32825,N_35071);
nor U47682 (N_47682,N_31429,N_32530);
nand U47683 (N_47683,N_35513,N_39518);
and U47684 (N_47684,N_39541,N_34766);
nand U47685 (N_47685,N_38800,N_33796);
or U47686 (N_47686,N_35047,N_30514);
nor U47687 (N_47687,N_38587,N_38401);
nand U47688 (N_47688,N_39241,N_33683);
nand U47689 (N_47689,N_35089,N_32230);
nor U47690 (N_47690,N_37162,N_36501);
or U47691 (N_47691,N_38151,N_35010);
or U47692 (N_47692,N_35908,N_34562);
nand U47693 (N_47693,N_36472,N_31748);
nor U47694 (N_47694,N_31567,N_39451);
nand U47695 (N_47695,N_30199,N_39989);
and U47696 (N_47696,N_31597,N_39413);
or U47697 (N_47697,N_34688,N_36802);
or U47698 (N_47698,N_30493,N_39825);
or U47699 (N_47699,N_34008,N_34155);
nor U47700 (N_47700,N_34748,N_30037);
and U47701 (N_47701,N_39397,N_39795);
xnor U47702 (N_47702,N_37949,N_31168);
and U47703 (N_47703,N_31228,N_34030);
nand U47704 (N_47704,N_30341,N_35284);
nor U47705 (N_47705,N_37195,N_38569);
nor U47706 (N_47706,N_30222,N_34810);
and U47707 (N_47707,N_32508,N_33150);
and U47708 (N_47708,N_33118,N_37463);
and U47709 (N_47709,N_35944,N_32425);
or U47710 (N_47710,N_34479,N_39781);
and U47711 (N_47711,N_35757,N_34974);
xor U47712 (N_47712,N_33831,N_35345);
nand U47713 (N_47713,N_35172,N_30732);
and U47714 (N_47714,N_35051,N_39148);
nor U47715 (N_47715,N_39835,N_39587);
or U47716 (N_47716,N_35205,N_39488);
xnor U47717 (N_47717,N_34538,N_37840);
or U47718 (N_47718,N_36422,N_33280);
or U47719 (N_47719,N_39431,N_39376);
and U47720 (N_47720,N_38355,N_34160);
and U47721 (N_47721,N_30719,N_31576);
and U47722 (N_47722,N_35975,N_33210);
xor U47723 (N_47723,N_34761,N_33363);
xnor U47724 (N_47724,N_36485,N_33257);
and U47725 (N_47725,N_38366,N_30324);
and U47726 (N_47726,N_32500,N_39584);
nor U47727 (N_47727,N_36571,N_38614);
and U47728 (N_47728,N_35506,N_32086);
nor U47729 (N_47729,N_34056,N_35457);
nand U47730 (N_47730,N_39758,N_38964);
or U47731 (N_47731,N_32815,N_33270);
and U47732 (N_47732,N_39225,N_31275);
nand U47733 (N_47733,N_39881,N_39615);
nor U47734 (N_47734,N_37657,N_36570);
and U47735 (N_47735,N_36923,N_33923);
nand U47736 (N_47736,N_31151,N_34949);
and U47737 (N_47737,N_33382,N_36770);
and U47738 (N_47738,N_37717,N_34673);
or U47739 (N_47739,N_38887,N_30286);
and U47740 (N_47740,N_32081,N_37040);
or U47741 (N_47741,N_31313,N_38285);
and U47742 (N_47742,N_37995,N_38166);
and U47743 (N_47743,N_34705,N_35127);
nand U47744 (N_47744,N_35226,N_39037);
or U47745 (N_47745,N_34018,N_39436);
and U47746 (N_47746,N_39517,N_30871);
nand U47747 (N_47747,N_30126,N_33690);
or U47748 (N_47748,N_32786,N_36974);
nand U47749 (N_47749,N_30611,N_31082);
or U47750 (N_47750,N_34473,N_37393);
nand U47751 (N_47751,N_30826,N_30382);
nand U47752 (N_47752,N_33380,N_37612);
or U47753 (N_47753,N_37147,N_31432);
and U47754 (N_47754,N_39118,N_36347);
and U47755 (N_47755,N_34054,N_38565);
and U47756 (N_47756,N_38833,N_35759);
and U47757 (N_47757,N_34742,N_38176);
xor U47758 (N_47758,N_30078,N_30925);
xnor U47759 (N_47759,N_37200,N_34264);
nand U47760 (N_47760,N_33508,N_36542);
nor U47761 (N_47761,N_33541,N_33166);
nand U47762 (N_47762,N_33678,N_33968);
xnor U47763 (N_47763,N_38851,N_36381);
and U47764 (N_47764,N_36742,N_30831);
or U47765 (N_47765,N_35267,N_32667);
nor U47766 (N_47766,N_35947,N_38864);
and U47767 (N_47767,N_34911,N_37141);
or U47768 (N_47768,N_39054,N_33656);
and U47769 (N_47769,N_34784,N_34706);
nor U47770 (N_47770,N_38684,N_31869);
nor U47771 (N_47771,N_33141,N_35614);
xor U47772 (N_47772,N_32425,N_38275);
xnor U47773 (N_47773,N_30443,N_39000);
and U47774 (N_47774,N_35094,N_37616);
nand U47775 (N_47775,N_32261,N_38026);
nor U47776 (N_47776,N_32703,N_33427);
or U47777 (N_47777,N_31935,N_36450);
nand U47778 (N_47778,N_30648,N_33487);
and U47779 (N_47779,N_33620,N_30318);
or U47780 (N_47780,N_31649,N_31804);
nor U47781 (N_47781,N_38466,N_33708);
nand U47782 (N_47782,N_36024,N_37172);
nor U47783 (N_47783,N_39215,N_36211);
or U47784 (N_47784,N_37867,N_36601);
nand U47785 (N_47785,N_36470,N_38320);
and U47786 (N_47786,N_33633,N_31331);
and U47787 (N_47787,N_30386,N_32230);
nand U47788 (N_47788,N_38005,N_37794);
or U47789 (N_47789,N_34244,N_36812);
or U47790 (N_47790,N_38349,N_32645);
nand U47791 (N_47791,N_38507,N_35516);
xor U47792 (N_47792,N_31266,N_36961);
nor U47793 (N_47793,N_36917,N_30591);
nand U47794 (N_47794,N_38152,N_35433);
nand U47795 (N_47795,N_36467,N_35622);
nand U47796 (N_47796,N_35861,N_37981);
nand U47797 (N_47797,N_32535,N_30132);
xor U47798 (N_47798,N_34034,N_31083);
nand U47799 (N_47799,N_30459,N_34628);
nor U47800 (N_47800,N_39126,N_39998);
nor U47801 (N_47801,N_39311,N_31272);
or U47802 (N_47802,N_30789,N_30878);
or U47803 (N_47803,N_37863,N_30017);
and U47804 (N_47804,N_37369,N_31795);
nand U47805 (N_47805,N_37881,N_31927);
or U47806 (N_47806,N_33629,N_38030);
nand U47807 (N_47807,N_30818,N_37455);
nand U47808 (N_47808,N_38063,N_37702);
nand U47809 (N_47809,N_36287,N_39573);
xor U47810 (N_47810,N_34543,N_31306);
nor U47811 (N_47811,N_31401,N_30999);
or U47812 (N_47812,N_32905,N_31403);
xor U47813 (N_47813,N_32449,N_39207);
or U47814 (N_47814,N_34828,N_36407);
xor U47815 (N_47815,N_30644,N_33922);
xnor U47816 (N_47816,N_37422,N_37379);
nand U47817 (N_47817,N_36982,N_30912);
or U47818 (N_47818,N_38865,N_33238);
xnor U47819 (N_47819,N_36358,N_37575);
nand U47820 (N_47820,N_32266,N_34859);
xnor U47821 (N_47821,N_36974,N_32379);
nor U47822 (N_47822,N_30979,N_31768);
nor U47823 (N_47823,N_37376,N_34635);
and U47824 (N_47824,N_34835,N_39007);
or U47825 (N_47825,N_39107,N_31255);
nand U47826 (N_47826,N_37345,N_39718);
and U47827 (N_47827,N_37250,N_36405);
and U47828 (N_47828,N_33349,N_31861);
or U47829 (N_47829,N_35637,N_32288);
nor U47830 (N_47830,N_33877,N_32284);
xor U47831 (N_47831,N_35860,N_33115);
and U47832 (N_47832,N_32007,N_31246);
or U47833 (N_47833,N_33608,N_35529);
or U47834 (N_47834,N_39037,N_33910);
or U47835 (N_47835,N_37441,N_30883);
or U47836 (N_47836,N_31727,N_33939);
nor U47837 (N_47837,N_38101,N_32911);
nor U47838 (N_47838,N_31428,N_34191);
or U47839 (N_47839,N_35249,N_38753);
and U47840 (N_47840,N_30537,N_37225);
or U47841 (N_47841,N_31459,N_35641);
and U47842 (N_47842,N_32449,N_30301);
nor U47843 (N_47843,N_36093,N_35807);
or U47844 (N_47844,N_38799,N_33037);
or U47845 (N_47845,N_34531,N_30514);
or U47846 (N_47846,N_39893,N_34491);
or U47847 (N_47847,N_38896,N_32505);
and U47848 (N_47848,N_36852,N_38960);
and U47849 (N_47849,N_31610,N_38656);
and U47850 (N_47850,N_39090,N_37007);
nor U47851 (N_47851,N_32078,N_37573);
nor U47852 (N_47852,N_35832,N_33967);
or U47853 (N_47853,N_32456,N_33798);
or U47854 (N_47854,N_31476,N_30509);
or U47855 (N_47855,N_35350,N_37027);
or U47856 (N_47856,N_33594,N_36050);
or U47857 (N_47857,N_32833,N_33183);
and U47858 (N_47858,N_34298,N_35498);
or U47859 (N_47859,N_34532,N_31073);
nand U47860 (N_47860,N_37478,N_33422);
nand U47861 (N_47861,N_35107,N_31423);
nand U47862 (N_47862,N_39313,N_38403);
or U47863 (N_47863,N_34251,N_35600);
xnor U47864 (N_47864,N_39339,N_39939);
or U47865 (N_47865,N_35443,N_32217);
nor U47866 (N_47866,N_31776,N_35635);
and U47867 (N_47867,N_32950,N_34894);
and U47868 (N_47868,N_39320,N_39973);
xnor U47869 (N_47869,N_39700,N_38165);
nand U47870 (N_47870,N_35269,N_32594);
and U47871 (N_47871,N_36781,N_30458);
and U47872 (N_47872,N_37494,N_33909);
and U47873 (N_47873,N_34254,N_30911);
nor U47874 (N_47874,N_31936,N_38984);
xor U47875 (N_47875,N_32761,N_36151);
nand U47876 (N_47876,N_35586,N_30784);
or U47877 (N_47877,N_37674,N_35554);
nor U47878 (N_47878,N_33905,N_39843);
and U47879 (N_47879,N_32663,N_38973);
nor U47880 (N_47880,N_32868,N_35077);
nor U47881 (N_47881,N_30834,N_32237);
and U47882 (N_47882,N_38212,N_37970);
and U47883 (N_47883,N_35114,N_35083);
nor U47884 (N_47884,N_33384,N_39444);
or U47885 (N_47885,N_38787,N_30706);
nor U47886 (N_47886,N_32503,N_37600);
or U47887 (N_47887,N_36356,N_37406);
and U47888 (N_47888,N_35727,N_35162);
nand U47889 (N_47889,N_30864,N_34218);
or U47890 (N_47890,N_35465,N_32409);
nand U47891 (N_47891,N_31007,N_36706);
nor U47892 (N_47892,N_37415,N_35221);
or U47893 (N_47893,N_35399,N_34321);
and U47894 (N_47894,N_32611,N_35830);
nand U47895 (N_47895,N_38527,N_30874);
nor U47896 (N_47896,N_39327,N_33167);
nand U47897 (N_47897,N_36607,N_33790);
xor U47898 (N_47898,N_34206,N_38148);
nand U47899 (N_47899,N_35834,N_36028);
nor U47900 (N_47900,N_39919,N_36510);
nand U47901 (N_47901,N_36003,N_30372);
xor U47902 (N_47902,N_32142,N_34315);
nand U47903 (N_47903,N_39660,N_32745);
and U47904 (N_47904,N_31029,N_36896);
nor U47905 (N_47905,N_37067,N_36163);
xnor U47906 (N_47906,N_38033,N_30618);
nor U47907 (N_47907,N_34791,N_34339);
nand U47908 (N_47908,N_38393,N_38248);
xnor U47909 (N_47909,N_33653,N_34204);
and U47910 (N_47910,N_37499,N_30111);
nor U47911 (N_47911,N_34248,N_33390);
xnor U47912 (N_47912,N_35853,N_37019);
nor U47913 (N_47913,N_39212,N_39868);
or U47914 (N_47914,N_31355,N_38610);
nand U47915 (N_47915,N_37818,N_35450);
or U47916 (N_47916,N_36431,N_36780);
nor U47917 (N_47917,N_31863,N_34840);
nand U47918 (N_47918,N_33760,N_30668);
and U47919 (N_47919,N_38101,N_39570);
nor U47920 (N_47920,N_32411,N_38208);
nor U47921 (N_47921,N_34212,N_31866);
and U47922 (N_47922,N_39713,N_30826);
nand U47923 (N_47923,N_38162,N_34880);
nand U47924 (N_47924,N_37806,N_38537);
nand U47925 (N_47925,N_37981,N_37459);
xnor U47926 (N_47926,N_37244,N_32651);
or U47927 (N_47927,N_31736,N_32877);
or U47928 (N_47928,N_30469,N_38084);
and U47929 (N_47929,N_37158,N_32329);
and U47930 (N_47930,N_30346,N_30599);
and U47931 (N_47931,N_34027,N_30587);
and U47932 (N_47932,N_31506,N_33552);
nand U47933 (N_47933,N_30625,N_35946);
nor U47934 (N_47934,N_39353,N_31639);
or U47935 (N_47935,N_39329,N_37075);
or U47936 (N_47936,N_38457,N_31146);
and U47937 (N_47937,N_31366,N_32708);
and U47938 (N_47938,N_33269,N_34203);
nand U47939 (N_47939,N_38370,N_30196);
and U47940 (N_47940,N_31181,N_34395);
xnor U47941 (N_47941,N_37226,N_38643);
nor U47942 (N_47942,N_30018,N_30564);
nand U47943 (N_47943,N_37850,N_31581);
or U47944 (N_47944,N_31867,N_34447);
and U47945 (N_47945,N_37500,N_33475);
nor U47946 (N_47946,N_34775,N_38574);
nand U47947 (N_47947,N_34830,N_35393);
nor U47948 (N_47948,N_39028,N_36121);
nand U47949 (N_47949,N_33634,N_30486);
nor U47950 (N_47950,N_32724,N_33342);
or U47951 (N_47951,N_39500,N_31076);
and U47952 (N_47952,N_30645,N_32311);
nand U47953 (N_47953,N_38744,N_35456);
or U47954 (N_47954,N_33035,N_38870);
nand U47955 (N_47955,N_33593,N_37173);
xnor U47956 (N_47956,N_39216,N_36996);
nor U47957 (N_47957,N_30824,N_32026);
and U47958 (N_47958,N_30381,N_39543);
and U47959 (N_47959,N_34533,N_36577);
or U47960 (N_47960,N_33613,N_30142);
or U47961 (N_47961,N_37685,N_34787);
nor U47962 (N_47962,N_30296,N_36629);
and U47963 (N_47963,N_33429,N_35661);
or U47964 (N_47964,N_38821,N_30847);
nand U47965 (N_47965,N_30617,N_38389);
nor U47966 (N_47966,N_30186,N_39624);
or U47967 (N_47967,N_34837,N_32374);
and U47968 (N_47968,N_36966,N_39819);
and U47969 (N_47969,N_39249,N_33126);
and U47970 (N_47970,N_31453,N_33572);
xor U47971 (N_47971,N_31299,N_34807);
xor U47972 (N_47972,N_34280,N_39695);
nand U47973 (N_47973,N_35287,N_30312);
nor U47974 (N_47974,N_33790,N_32936);
and U47975 (N_47975,N_39831,N_34700);
and U47976 (N_47976,N_38560,N_30710);
and U47977 (N_47977,N_34012,N_38099);
or U47978 (N_47978,N_33287,N_35237);
or U47979 (N_47979,N_34605,N_37757);
nand U47980 (N_47980,N_36341,N_38009);
nor U47981 (N_47981,N_35592,N_30286);
xnor U47982 (N_47982,N_36738,N_36268);
and U47983 (N_47983,N_35027,N_32775);
and U47984 (N_47984,N_39912,N_38502);
nand U47985 (N_47985,N_38601,N_37249);
nand U47986 (N_47986,N_39591,N_31012);
and U47987 (N_47987,N_30889,N_35418);
or U47988 (N_47988,N_31873,N_33047);
xnor U47989 (N_47989,N_33648,N_39262);
or U47990 (N_47990,N_38989,N_35096);
and U47991 (N_47991,N_31863,N_35581);
or U47992 (N_47992,N_36279,N_31487);
xnor U47993 (N_47993,N_37442,N_30556);
and U47994 (N_47994,N_32349,N_30287);
nand U47995 (N_47995,N_38770,N_33095);
and U47996 (N_47996,N_36402,N_38351);
and U47997 (N_47997,N_39957,N_39833);
or U47998 (N_47998,N_33898,N_38619);
and U47999 (N_47999,N_34362,N_36731);
nor U48000 (N_48000,N_30633,N_33329);
nand U48001 (N_48001,N_36706,N_35470);
xnor U48002 (N_48002,N_32543,N_35424);
or U48003 (N_48003,N_38816,N_32202);
or U48004 (N_48004,N_36701,N_31485);
or U48005 (N_48005,N_30712,N_33148);
xnor U48006 (N_48006,N_35431,N_39182);
or U48007 (N_48007,N_36139,N_36697);
nor U48008 (N_48008,N_32378,N_31005);
or U48009 (N_48009,N_34778,N_36783);
and U48010 (N_48010,N_39296,N_34856);
and U48011 (N_48011,N_33116,N_36671);
or U48012 (N_48012,N_32462,N_31524);
nand U48013 (N_48013,N_31074,N_35680);
and U48014 (N_48014,N_31296,N_32729);
and U48015 (N_48015,N_35320,N_30862);
nand U48016 (N_48016,N_38498,N_31172);
nor U48017 (N_48017,N_36349,N_33208);
xnor U48018 (N_48018,N_36749,N_37809);
nand U48019 (N_48019,N_36738,N_33081);
or U48020 (N_48020,N_33216,N_35347);
nor U48021 (N_48021,N_36556,N_38002);
xnor U48022 (N_48022,N_34937,N_35828);
nor U48023 (N_48023,N_36098,N_35633);
and U48024 (N_48024,N_30537,N_37035);
nand U48025 (N_48025,N_39163,N_36957);
or U48026 (N_48026,N_33288,N_30407);
nand U48027 (N_48027,N_37805,N_33954);
xor U48028 (N_48028,N_34315,N_32309);
and U48029 (N_48029,N_37728,N_32127);
nor U48030 (N_48030,N_37681,N_34897);
nand U48031 (N_48031,N_36299,N_35142);
xnor U48032 (N_48032,N_39784,N_32170);
and U48033 (N_48033,N_37805,N_38967);
and U48034 (N_48034,N_30108,N_31650);
or U48035 (N_48035,N_32355,N_32918);
nand U48036 (N_48036,N_37120,N_39844);
or U48037 (N_48037,N_37163,N_30285);
nand U48038 (N_48038,N_31018,N_36074);
nor U48039 (N_48039,N_30899,N_32215);
or U48040 (N_48040,N_35097,N_32182);
and U48041 (N_48041,N_33758,N_33208);
nor U48042 (N_48042,N_36521,N_31067);
and U48043 (N_48043,N_32280,N_32998);
nor U48044 (N_48044,N_35527,N_38990);
and U48045 (N_48045,N_34542,N_39652);
and U48046 (N_48046,N_34753,N_38492);
or U48047 (N_48047,N_35921,N_32381);
nor U48048 (N_48048,N_33376,N_37021);
and U48049 (N_48049,N_35345,N_35948);
xor U48050 (N_48050,N_31198,N_34072);
xor U48051 (N_48051,N_39221,N_37211);
nand U48052 (N_48052,N_34303,N_37523);
and U48053 (N_48053,N_36147,N_36644);
nand U48054 (N_48054,N_32273,N_34701);
nor U48055 (N_48055,N_34686,N_37034);
and U48056 (N_48056,N_31134,N_38443);
and U48057 (N_48057,N_35532,N_38196);
or U48058 (N_48058,N_37309,N_32459);
and U48059 (N_48059,N_30975,N_35071);
xnor U48060 (N_48060,N_34960,N_34402);
and U48061 (N_48061,N_31644,N_33356);
or U48062 (N_48062,N_39050,N_35601);
nand U48063 (N_48063,N_39375,N_37306);
nor U48064 (N_48064,N_34829,N_35176);
and U48065 (N_48065,N_30060,N_37503);
xor U48066 (N_48066,N_35680,N_38556);
nand U48067 (N_48067,N_32420,N_30988);
or U48068 (N_48068,N_30449,N_36086);
nand U48069 (N_48069,N_32085,N_32736);
and U48070 (N_48070,N_30688,N_36364);
and U48071 (N_48071,N_30793,N_33769);
or U48072 (N_48072,N_33144,N_32710);
nor U48073 (N_48073,N_30727,N_38055);
or U48074 (N_48074,N_36617,N_32215);
or U48075 (N_48075,N_39616,N_33490);
nor U48076 (N_48076,N_35137,N_34192);
nand U48077 (N_48077,N_35399,N_32729);
nand U48078 (N_48078,N_33095,N_30891);
nor U48079 (N_48079,N_39671,N_39292);
nand U48080 (N_48080,N_33790,N_34326);
or U48081 (N_48081,N_39649,N_38038);
nand U48082 (N_48082,N_39409,N_34297);
and U48083 (N_48083,N_39561,N_39492);
and U48084 (N_48084,N_36413,N_34390);
and U48085 (N_48085,N_39125,N_34473);
or U48086 (N_48086,N_38950,N_33303);
nor U48087 (N_48087,N_34839,N_33666);
or U48088 (N_48088,N_33313,N_34887);
nor U48089 (N_48089,N_35494,N_35809);
nor U48090 (N_48090,N_35047,N_32950);
and U48091 (N_48091,N_38400,N_32325);
and U48092 (N_48092,N_31032,N_34784);
and U48093 (N_48093,N_35003,N_39175);
nand U48094 (N_48094,N_34826,N_31063);
nor U48095 (N_48095,N_30888,N_39302);
nor U48096 (N_48096,N_35181,N_38685);
xor U48097 (N_48097,N_30934,N_37190);
nor U48098 (N_48098,N_30298,N_38733);
and U48099 (N_48099,N_32747,N_30619);
nor U48100 (N_48100,N_39312,N_37934);
nand U48101 (N_48101,N_33493,N_37516);
nand U48102 (N_48102,N_37974,N_34751);
nand U48103 (N_48103,N_38833,N_39365);
nor U48104 (N_48104,N_32879,N_39942);
nand U48105 (N_48105,N_38101,N_32063);
nand U48106 (N_48106,N_37713,N_31770);
and U48107 (N_48107,N_39357,N_31730);
nor U48108 (N_48108,N_33653,N_37211);
xor U48109 (N_48109,N_39814,N_36070);
and U48110 (N_48110,N_30550,N_38821);
nor U48111 (N_48111,N_35300,N_37324);
and U48112 (N_48112,N_35796,N_37047);
nor U48113 (N_48113,N_31268,N_33255);
nand U48114 (N_48114,N_38313,N_35349);
nor U48115 (N_48115,N_30300,N_38518);
xor U48116 (N_48116,N_34207,N_37203);
and U48117 (N_48117,N_37749,N_37099);
nor U48118 (N_48118,N_33796,N_38894);
xnor U48119 (N_48119,N_34969,N_31079);
nand U48120 (N_48120,N_31963,N_37211);
and U48121 (N_48121,N_32698,N_33320);
and U48122 (N_48122,N_36094,N_32054);
and U48123 (N_48123,N_33634,N_39349);
nand U48124 (N_48124,N_38417,N_39734);
nand U48125 (N_48125,N_35055,N_32338);
and U48126 (N_48126,N_34553,N_38741);
or U48127 (N_48127,N_32621,N_39002);
nand U48128 (N_48128,N_39117,N_39399);
or U48129 (N_48129,N_36588,N_37186);
nand U48130 (N_48130,N_37399,N_32180);
or U48131 (N_48131,N_36944,N_38041);
nand U48132 (N_48132,N_39030,N_31004);
nor U48133 (N_48133,N_31000,N_33746);
or U48134 (N_48134,N_30442,N_32520);
nor U48135 (N_48135,N_36882,N_33925);
nand U48136 (N_48136,N_38154,N_30023);
nor U48137 (N_48137,N_38700,N_38505);
xor U48138 (N_48138,N_30782,N_30342);
or U48139 (N_48139,N_30457,N_38224);
or U48140 (N_48140,N_34876,N_39797);
or U48141 (N_48141,N_30866,N_32747);
or U48142 (N_48142,N_37847,N_35376);
nand U48143 (N_48143,N_34982,N_33593);
and U48144 (N_48144,N_35799,N_37958);
nand U48145 (N_48145,N_38272,N_30891);
nor U48146 (N_48146,N_31919,N_31243);
nand U48147 (N_48147,N_31329,N_37233);
nand U48148 (N_48148,N_38970,N_31282);
and U48149 (N_48149,N_39945,N_35549);
nand U48150 (N_48150,N_31811,N_31586);
nand U48151 (N_48151,N_37987,N_30293);
nor U48152 (N_48152,N_32274,N_31589);
or U48153 (N_48153,N_34140,N_35738);
nand U48154 (N_48154,N_37532,N_34011);
nand U48155 (N_48155,N_35640,N_39829);
nor U48156 (N_48156,N_34067,N_31598);
xor U48157 (N_48157,N_35125,N_33045);
and U48158 (N_48158,N_39865,N_35459);
or U48159 (N_48159,N_38249,N_36775);
and U48160 (N_48160,N_33050,N_30035);
nand U48161 (N_48161,N_35984,N_35176);
nand U48162 (N_48162,N_33579,N_39849);
xor U48163 (N_48163,N_38048,N_34819);
nor U48164 (N_48164,N_31522,N_34009);
and U48165 (N_48165,N_33443,N_34653);
or U48166 (N_48166,N_34647,N_38243);
and U48167 (N_48167,N_34431,N_39294);
and U48168 (N_48168,N_31727,N_38383);
nand U48169 (N_48169,N_38308,N_30879);
or U48170 (N_48170,N_30997,N_33650);
nand U48171 (N_48171,N_39991,N_30855);
nand U48172 (N_48172,N_32943,N_31407);
or U48173 (N_48173,N_33931,N_30047);
and U48174 (N_48174,N_35813,N_35654);
or U48175 (N_48175,N_32158,N_30841);
nor U48176 (N_48176,N_34978,N_39634);
and U48177 (N_48177,N_37903,N_39000);
and U48178 (N_48178,N_36209,N_31591);
or U48179 (N_48179,N_39144,N_30432);
or U48180 (N_48180,N_33676,N_33275);
and U48181 (N_48181,N_37054,N_38333);
and U48182 (N_48182,N_30934,N_33585);
nor U48183 (N_48183,N_33195,N_37863);
nand U48184 (N_48184,N_39475,N_37794);
and U48185 (N_48185,N_34732,N_30668);
nor U48186 (N_48186,N_38231,N_33590);
or U48187 (N_48187,N_35325,N_35024);
or U48188 (N_48188,N_31645,N_39670);
or U48189 (N_48189,N_30603,N_33609);
and U48190 (N_48190,N_37048,N_32913);
nor U48191 (N_48191,N_38364,N_37018);
and U48192 (N_48192,N_34277,N_35034);
and U48193 (N_48193,N_31053,N_30729);
and U48194 (N_48194,N_33566,N_35631);
nor U48195 (N_48195,N_37504,N_36150);
and U48196 (N_48196,N_37338,N_35228);
xor U48197 (N_48197,N_30122,N_37021);
nor U48198 (N_48198,N_31972,N_34965);
and U48199 (N_48199,N_35338,N_38154);
xor U48200 (N_48200,N_35949,N_31763);
nor U48201 (N_48201,N_30436,N_33322);
and U48202 (N_48202,N_33093,N_31069);
nor U48203 (N_48203,N_39817,N_32957);
or U48204 (N_48204,N_34397,N_34053);
and U48205 (N_48205,N_39502,N_36554);
nand U48206 (N_48206,N_31770,N_37533);
nand U48207 (N_48207,N_37736,N_35346);
xnor U48208 (N_48208,N_34701,N_37016);
or U48209 (N_48209,N_31294,N_30954);
xnor U48210 (N_48210,N_33213,N_36824);
xnor U48211 (N_48211,N_35820,N_37670);
nor U48212 (N_48212,N_34466,N_31729);
and U48213 (N_48213,N_30965,N_31382);
nand U48214 (N_48214,N_37443,N_39125);
and U48215 (N_48215,N_36815,N_36991);
and U48216 (N_48216,N_32129,N_31449);
nand U48217 (N_48217,N_30906,N_39179);
nor U48218 (N_48218,N_34636,N_34212);
xnor U48219 (N_48219,N_35039,N_31153);
nand U48220 (N_48220,N_34721,N_38050);
nand U48221 (N_48221,N_37372,N_32612);
or U48222 (N_48222,N_33814,N_33894);
and U48223 (N_48223,N_30692,N_35290);
nor U48224 (N_48224,N_34314,N_32110);
xnor U48225 (N_48225,N_37184,N_36851);
nor U48226 (N_48226,N_30493,N_31332);
nor U48227 (N_48227,N_32786,N_30089);
nor U48228 (N_48228,N_32555,N_33164);
nor U48229 (N_48229,N_31872,N_35800);
nand U48230 (N_48230,N_33227,N_37642);
nand U48231 (N_48231,N_37261,N_33009);
nand U48232 (N_48232,N_33202,N_32447);
xnor U48233 (N_48233,N_33701,N_34431);
nand U48234 (N_48234,N_39222,N_37034);
and U48235 (N_48235,N_37858,N_32103);
nand U48236 (N_48236,N_34422,N_31351);
and U48237 (N_48237,N_30323,N_30880);
nor U48238 (N_48238,N_31323,N_36259);
or U48239 (N_48239,N_34043,N_30066);
nand U48240 (N_48240,N_35751,N_37677);
nand U48241 (N_48241,N_35142,N_38735);
or U48242 (N_48242,N_33777,N_36122);
and U48243 (N_48243,N_35598,N_30432);
nor U48244 (N_48244,N_37048,N_33229);
nand U48245 (N_48245,N_35786,N_32691);
and U48246 (N_48246,N_30062,N_33979);
and U48247 (N_48247,N_39896,N_33857);
or U48248 (N_48248,N_38705,N_37554);
nand U48249 (N_48249,N_38676,N_35807);
or U48250 (N_48250,N_38374,N_38084);
and U48251 (N_48251,N_33519,N_31520);
nor U48252 (N_48252,N_35532,N_31946);
nor U48253 (N_48253,N_31929,N_33371);
and U48254 (N_48254,N_30999,N_33735);
nor U48255 (N_48255,N_38839,N_34262);
nor U48256 (N_48256,N_37938,N_36898);
or U48257 (N_48257,N_33759,N_37314);
or U48258 (N_48258,N_38451,N_31631);
and U48259 (N_48259,N_39046,N_32207);
and U48260 (N_48260,N_36334,N_31466);
or U48261 (N_48261,N_32374,N_36766);
nand U48262 (N_48262,N_30944,N_32748);
or U48263 (N_48263,N_30018,N_31344);
nand U48264 (N_48264,N_35800,N_35428);
and U48265 (N_48265,N_31122,N_33227);
nor U48266 (N_48266,N_36625,N_38543);
or U48267 (N_48267,N_39494,N_37003);
or U48268 (N_48268,N_37924,N_30186);
nand U48269 (N_48269,N_38698,N_32816);
nand U48270 (N_48270,N_38805,N_34479);
or U48271 (N_48271,N_36857,N_34055);
or U48272 (N_48272,N_33249,N_32886);
nor U48273 (N_48273,N_37941,N_30090);
and U48274 (N_48274,N_30921,N_32475);
or U48275 (N_48275,N_36416,N_33032);
nor U48276 (N_48276,N_37819,N_38071);
nand U48277 (N_48277,N_31361,N_34082);
nor U48278 (N_48278,N_31765,N_39158);
or U48279 (N_48279,N_35150,N_31558);
or U48280 (N_48280,N_34917,N_38331);
nand U48281 (N_48281,N_31377,N_31419);
nor U48282 (N_48282,N_36183,N_31411);
nand U48283 (N_48283,N_31331,N_38640);
nand U48284 (N_48284,N_34687,N_36468);
nand U48285 (N_48285,N_39187,N_33807);
nand U48286 (N_48286,N_34508,N_35151);
nor U48287 (N_48287,N_30933,N_30572);
or U48288 (N_48288,N_30681,N_30107);
and U48289 (N_48289,N_37652,N_38383);
or U48290 (N_48290,N_35865,N_39234);
and U48291 (N_48291,N_30670,N_35048);
nor U48292 (N_48292,N_34391,N_32530);
or U48293 (N_48293,N_38969,N_37998);
and U48294 (N_48294,N_36643,N_39181);
or U48295 (N_48295,N_35150,N_31739);
and U48296 (N_48296,N_32514,N_39948);
xor U48297 (N_48297,N_31370,N_36770);
nand U48298 (N_48298,N_39223,N_32335);
or U48299 (N_48299,N_37543,N_36901);
and U48300 (N_48300,N_35052,N_37245);
or U48301 (N_48301,N_34465,N_37984);
nand U48302 (N_48302,N_31328,N_33425);
or U48303 (N_48303,N_33628,N_39395);
xnor U48304 (N_48304,N_37074,N_31671);
or U48305 (N_48305,N_32459,N_39739);
nor U48306 (N_48306,N_37177,N_37448);
nor U48307 (N_48307,N_30540,N_38292);
nand U48308 (N_48308,N_36176,N_33828);
or U48309 (N_48309,N_35764,N_35528);
nor U48310 (N_48310,N_39279,N_37262);
or U48311 (N_48311,N_35170,N_31978);
and U48312 (N_48312,N_31939,N_32759);
and U48313 (N_48313,N_36136,N_30355);
and U48314 (N_48314,N_36464,N_31599);
nor U48315 (N_48315,N_31916,N_37384);
nor U48316 (N_48316,N_35894,N_37740);
or U48317 (N_48317,N_34590,N_39786);
xor U48318 (N_48318,N_36759,N_33553);
nand U48319 (N_48319,N_39967,N_38792);
nand U48320 (N_48320,N_39170,N_36004);
or U48321 (N_48321,N_34423,N_31563);
and U48322 (N_48322,N_34776,N_33398);
nor U48323 (N_48323,N_32361,N_39403);
nor U48324 (N_48324,N_39210,N_33291);
and U48325 (N_48325,N_35076,N_35884);
and U48326 (N_48326,N_37247,N_32075);
nand U48327 (N_48327,N_34734,N_37686);
or U48328 (N_48328,N_35316,N_30567);
or U48329 (N_48329,N_30746,N_31331);
and U48330 (N_48330,N_36090,N_33434);
xnor U48331 (N_48331,N_37721,N_36748);
and U48332 (N_48332,N_34070,N_39697);
nand U48333 (N_48333,N_35471,N_34569);
or U48334 (N_48334,N_38794,N_37022);
or U48335 (N_48335,N_32800,N_34599);
nor U48336 (N_48336,N_34973,N_33342);
or U48337 (N_48337,N_38290,N_30786);
nor U48338 (N_48338,N_34174,N_35661);
nand U48339 (N_48339,N_35446,N_34437);
and U48340 (N_48340,N_31735,N_32000);
nand U48341 (N_48341,N_35760,N_32952);
nor U48342 (N_48342,N_32504,N_37918);
and U48343 (N_48343,N_30110,N_36604);
nand U48344 (N_48344,N_34260,N_30450);
or U48345 (N_48345,N_37558,N_35140);
nor U48346 (N_48346,N_35615,N_38532);
nand U48347 (N_48347,N_37397,N_38411);
nand U48348 (N_48348,N_38659,N_31358);
nor U48349 (N_48349,N_31182,N_30751);
and U48350 (N_48350,N_39491,N_39402);
or U48351 (N_48351,N_31211,N_35349);
or U48352 (N_48352,N_31229,N_30576);
and U48353 (N_48353,N_36177,N_32445);
nand U48354 (N_48354,N_39601,N_32714);
or U48355 (N_48355,N_38876,N_31808);
or U48356 (N_48356,N_31376,N_33394);
xor U48357 (N_48357,N_37959,N_30249);
and U48358 (N_48358,N_33466,N_30656);
or U48359 (N_48359,N_31342,N_34873);
or U48360 (N_48360,N_37260,N_30970);
and U48361 (N_48361,N_35427,N_34162);
nand U48362 (N_48362,N_36975,N_36065);
or U48363 (N_48363,N_32867,N_30144);
and U48364 (N_48364,N_36028,N_34286);
nor U48365 (N_48365,N_33377,N_35910);
or U48366 (N_48366,N_36082,N_37185);
nand U48367 (N_48367,N_36923,N_35669);
or U48368 (N_48368,N_39885,N_32140);
or U48369 (N_48369,N_38100,N_30881);
nor U48370 (N_48370,N_32810,N_36153);
and U48371 (N_48371,N_34294,N_36851);
or U48372 (N_48372,N_34177,N_37492);
or U48373 (N_48373,N_32250,N_35013);
nor U48374 (N_48374,N_30225,N_33146);
and U48375 (N_48375,N_37161,N_35713);
and U48376 (N_48376,N_34302,N_30677);
and U48377 (N_48377,N_37155,N_39494);
xnor U48378 (N_48378,N_37875,N_35232);
and U48379 (N_48379,N_38341,N_39116);
xnor U48380 (N_48380,N_32148,N_31703);
xor U48381 (N_48381,N_30176,N_35482);
xor U48382 (N_48382,N_39210,N_35146);
nor U48383 (N_48383,N_33106,N_38559);
nand U48384 (N_48384,N_38615,N_34121);
and U48385 (N_48385,N_37424,N_38145);
and U48386 (N_48386,N_39237,N_33824);
nor U48387 (N_48387,N_33593,N_39753);
or U48388 (N_48388,N_36730,N_33208);
nand U48389 (N_48389,N_33488,N_33565);
nand U48390 (N_48390,N_38664,N_37593);
xor U48391 (N_48391,N_34557,N_39773);
and U48392 (N_48392,N_36081,N_39275);
nor U48393 (N_48393,N_35235,N_38365);
nand U48394 (N_48394,N_33116,N_32724);
and U48395 (N_48395,N_32179,N_33872);
and U48396 (N_48396,N_35617,N_35703);
nand U48397 (N_48397,N_36657,N_34764);
and U48398 (N_48398,N_35382,N_37000);
and U48399 (N_48399,N_39012,N_38428);
nand U48400 (N_48400,N_36538,N_34891);
or U48401 (N_48401,N_39549,N_39662);
nand U48402 (N_48402,N_34426,N_32091);
and U48403 (N_48403,N_31877,N_38749);
or U48404 (N_48404,N_31795,N_30152);
nor U48405 (N_48405,N_32555,N_31433);
or U48406 (N_48406,N_39609,N_30387);
or U48407 (N_48407,N_31308,N_32785);
nand U48408 (N_48408,N_31617,N_39027);
xor U48409 (N_48409,N_37454,N_33638);
and U48410 (N_48410,N_35304,N_30382);
xor U48411 (N_48411,N_39673,N_33923);
nor U48412 (N_48412,N_33974,N_32228);
or U48413 (N_48413,N_39421,N_33215);
nor U48414 (N_48414,N_36623,N_32703);
nand U48415 (N_48415,N_35734,N_34135);
and U48416 (N_48416,N_33877,N_36739);
and U48417 (N_48417,N_36996,N_33143);
or U48418 (N_48418,N_37478,N_39829);
or U48419 (N_48419,N_36788,N_34042);
xor U48420 (N_48420,N_33809,N_37423);
nand U48421 (N_48421,N_39837,N_32396);
nor U48422 (N_48422,N_36621,N_38437);
and U48423 (N_48423,N_34949,N_37610);
or U48424 (N_48424,N_30679,N_31580);
xor U48425 (N_48425,N_36774,N_38734);
or U48426 (N_48426,N_35025,N_35231);
nor U48427 (N_48427,N_30364,N_38243);
xnor U48428 (N_48428,N_32427,N_38429);
or U48429 (N_48429,N_38927,N_37517);
nand U48430 (N_48430,N_35627,N_35676);
nor U48431 (N_48431,N_38973,N_30170);
or U48432 (N_48432,N_35046,N_31347);
and U48433 (N_48433,N_33357,N_36674);
nand U48434 (N_48434,N_39277,N_32568);
nand U48435 (N_48435,N_39929,N_36601);
nor U48436 (N_48436,N_36947,N_33985);
nor U48437 (N_48437,N_37464,N_32604);
or U48438 (N_48438,N_30180,N_31531);
nand U48439 (N_48439,N_30798,N_39818);
nor U48440 (N_48440,N_38391,N_34780);
nor U48441 (N_48441,N_34792,N_32989);
and U48442 (N_48442,N_31190,N_31324);
nor U48443 (N_48443,N_30402,N_32773);
or U48444 (N_48444,N_33447,N_39543);
or U48445 (N_48445,N_35400,N_32729);
and U48446 (N_48446,N_36391,N_39120);
and U48447 (N_48447,N_34543,N_31958);
and U48448 (N_48448,N_36184,N_37535);
or U48449 (N_48449,N_39998,N_33986);
nor U48450 (N_48450,N_30270,N_32881);
nor U48451 (N_48451,N_35269,N_30691);
nand U48452 (N_48452,N_30046,N_34934);
nand U48453 (N_48453,N_32107,N_32953);
or U48454 (N_48454,N_38269,N_35360);
xnor U48455 (N_48455,N_38465,N_34926);
nand U48456 (N_48456,N_35625,N_35381);
nand U48457 (N_48457,N_34140,N_32716);
nor U48458 (N_48458,N_37964,N_35931);
or U48459 (N_48459,N_33258,N_39651);
and U48460 (N_48460,N_31057,N_31850);
or U48461 (N_48461,N_31743,N_32513);
and U48462 (N_48462,N_37093,N_32193);
nor U48463 (N_48463,N_39657,N_31850);
and U48464 (N_48464,N_35593,N_32436);
and U48465 (N_48465,N_38127,N_32817);
or U48466 (N_48466,N_32382,N_39451);
nand U48467 (N_48467,N_39060,N_32514);
nand U48468 (N_48468,N_30747,N_35159);
nor U48469 (N_48469,N_32457,N_34953);
nand U48470 (N_48470,N_38114,N_33280);
and U48471 (N_48471,N_37823,N_31886);
nor U48472 (N_48472,N_34521,N_31836);
xor U48473 (N_48473,N_36965,N_39682);
nand U48474 (N_48474,N_31730,N_35158);
nand U48475 (N_48475,N_38983,N_39740);
nor U48476 (N_48476,N_38743,N_34398);
nand U48477 (N_48477,N_33237,N_31642);
nor U48478 (N_48478,N_30375,N_36873);
xor U48479 (N_48479,N_38582,N_34885);
or U48480 (N_48480,N_35489,N_39028);
and U48481 (N_48481,N_37928,N_39260);
and U48482 (N_48482,N_39085,N_31866);
xor U48483 (N_48483,N_36298,N_31849);
nor U48484 (N_48484,N_32307,N_35637);
and U48485 (N_48485,N_36597,N_35220);
nor U48486 (N_48486,N_33534,N_38297);
nand U48487 (N_48487,N_39883,N_30397);
nand U48488 (N_48488,N_33468,N_36573);
nand U48489 (N_48489,N_33303,N_32181);
nor U48490 (N_48490,N_39198,N_39796);
nand U48491 (N_48491,N_30258,N_31791);
nand U48492 (N_48492,N_33358,N_34505);
xnor U48493 (N_48493,N_35274,N_30753);
nand U48494 (N_48494,N_35419,N_37080);
nand U48495 (N_48495,N_39101,N_38484);
nor U48496 (N_48496,N_36158,N_32680);
nor U48497 (N_48497,N_39123,N_32184);
nor U48498 (N_48498,N_31690,N_38357);
nand U48499 (N_48499,N_32835,N_30562);
or U48500 (N_48500,N_35183,N_36595);
and U48501 (N_48501,N_37915,N_36285);
or U48502 (N_48502,N_30905,N_32524);
nand U48503 (N_48503,N_31867,N_31634);
nand U48504 (N_48504,N_39492,N_34624);
or U48505 (N_48505,N_31896,N_30663);
nand U48506 (N_48506,N_37760,N_38990);
or U48507 (N_48507,N_35673,N_31989);
nand U48508 (N_48508,N_35774,N_37505);
and U48509 (N_48509,N_31317,N_39973);
or U48510 (N_48510,N_30533,N_30292);
or U48511 (N_48511,N_34450,N_34985);
xor U48512 (N_48512,N_34232,N_31231);
and U48513 (N_48513,N_39655,N_36261);
and U48514 (N_48514,N_32080,N_38425);
xnor U48515 (N_48515,N_38381,N_37080);
xor U48516 (N_48516,N_30252,N_33747);
or U48517 (N_48517,N_30912,N_36696);
and U48518 (N_48518,N_31252,N_33562);
or U48519 (N_48519,N_37529,N_38201);
or U48520 (N_48520,N_31485,N_35106);
nor U48521 (N_48521,N_35644,N_38740);
nand U48522 (N_48522,N_36596,N_31628);
nor U48523 (N_48523,N_30868,N_30902);
nand U48524 (N_48524,N_39276,N_39189);
nor U48525 (N_48525,N_36141,N_33863);
nand U48526 (N_48526,N_30641,N_33442);
nor U48527 (N_48527,N_34070,N_36161);
nand U48528 (N_48528,N_31230,N_30331);
nor U48529 (N_48529,N_37890,N_32417);
or U48530 (N_48530,N_37253,N_35307);
nor U48531 (N_48531,N_36124,N_31719);
and U48532 (N_48532,N_38555,N_36353);
nand U48533 (N_48533,N_33476,N_31045);
nand U48534 (N_48534,N_35029,N_39793);
and U48535 (N_48535,N_33364,N_30634);
and U48536 (N_48536,N_31465,N_39392);
nor U48537 (N_48537,N_36780,N_38922);
or U48538 (N_48538,N_33076,N_33117);
nor U48539 (N_48539,N_33977,N_31726);
nand U48540 (N_48540,N_36106,N_33134);
and U48541 (N_48541,N_32371,N_30310);
or U48542 (N_48542,N_38955,N_30450);
nor U48543 (N_48543,N_37757,N_38072);
nor U48544 (N_48544,N_35714,N_36222);
nor U48545 (N_48545,N_32161,N_31101);
or U48546 (N_48546,N_30390,N_35616);
and U48547 (N_48547,N_34315,N_35395);
nor U48548 (N_48548,N_37640,N_35739);
and U48549 (N_48549,N_34607,N_34691);
nand U48550 (N_48550,N_34672,N_37513);
and U48551 (N_48551,N_31228,N_30048);
nand U48552 (N_48552,N_37485,N_39603);
nor U48553 (N_48553,N_34468,N_33326);
or U48554 (N_48554,N_36812,N_31458);
nor U48555 (N_48555,N_33885,N_33502);
or U48556 (N_48556,N_37589,N_31345);
nor U48557 (N_48557,N_32908,N_36004);
nand U48558 (N_48558,N_36021,N_31824);
or U48559 (N_48559,N_30677,N_34165);
or U48560 (N_48560,N_34450,N_32780);
nor U48561 (N_48561,N_37309,N_33729);
nand U48562 (N_48562,N_31314,N_34629);
xor U48563 (N_48563,N_35969,N_38203);
nand U48564 (N_48564,N_39075,N_38614);
or U48565 (N_48565,N_31709,N_33442);
or U48566 (N_48566,N_33493,N_33781);
or U48567 (N_48567,N_37218,N_31846);
or U48568 (N_48568,N_32776,N_38076);
nand U48569 (N_48569,N_33790,N_39390);
nand U48570 (N_48570,N_37651,N_38115);
nor U48571 (N_48571,N_37527,N_37686);
and U48572 (N_48572,N_35874,N_35125);
nand U48573 (N_48573,N_35521,N_30802);
xor U48574 (N_48574,N_30244,N_38943);
nand U48575 (N_48575,N_38480,N_34728);
and U48576 (N_48576,N_36007,N_39050);
nand U48577 (N_48577,N_30346,N_36356);
or U48578 (N_48578,N_33105,N_31555);
xor U48579 (N_48579,N_39677,N_32554);
and U48580 (N_48580,N_35607,N_36011);
nand U48581 (N_48581,N_35322,N_36617);
and U48582 (N_48582,N_35336,N_35631);
and U48583 (N_48583,N_35051,N_34625);
and U48584 (N_48584,N_32132,N_34682);
and U48585 (N_48585,N_34228,N_39695);
nor U48586 (N_48586,N_38523,N_34691);
and U48587 (N_48587,N_32968,N_37193);
nand U48588 (N_48588,N_36170,N_30249);
nand U48589 (N_48589,N_39031,N_32693);
nor U48590 (N_48590,N_32729,N_34532);
or U48591 (N_48591,N_39114,N_31989);
nor U48592 (N_48592,N_32065,N_33453);
nand U48593 (N_48593,N_32342,N_30149);
and U48594 (N_48594,N_38371,N_33422);
nor U48595 (N_48595,N_37524,N_38889);
nand U48596 (N_48596,N_37371,N_32250);
nand U48597 (N_48597,N_33653,N_33720);
or U48598 (N_48598,N_32844,N_33992);
or U48599 (N_48599,N_36362,N_34701);
nand U48600 (N_48600,N_30153,N_35696);
or U48601 (N_48601,N_32156,N_37689);
or U48602 (N_48602,N_38598,N_34976);
xor U48603 (N_48603,N_37822,N_39022);
nor U48604 (N_48604,N_30639,N_38705);
xor U48605 (N_48605,N_33999,N_32017);
and U48606 (N_48606,N_36161,N_37763);
nand U48607 (N_48607,N_34985,N_31969);
nor U48608 (N_48608,N_32133,N_38644);
and U48609 (N_48609,N_30175,N_35448);
and U48610 (N_48610,N_39079,N_34862);
or U48611 (N_48611,N_39631,N_33298);
or U48612 (N_48612,N_33273,N_32811);
nand U48613 (N_48613,N_31912,N_39759);
or U48614 (N_48614,N_38015,N_34560);
and U48615 (N_48615,N_31735,N_34897);
nand U48616 (N_48616,N_38958,N_37901);
and U48617 (N_48617,N_30858,N_31410);
or U48618 (N_48618,N_31278,N_36649);
nand U48619 (N_48619,N_37009,N_30994);
and U48620 (N_48620,N_32199,N_38794);
nand U48621 (N_48621,N_36340,N_33879);
nand U48622 (N_48622,N_33560,N_36351);
or U48623 (N_48623,N_38162,N_38749);
and U48624 (N_48624,N_32665,N_34001);
nand U48625 (N_48625,N_33701,N_31506);
or U48626 (N_48626,N_31886,N_38137);
nor U48627 (N_48627,N_37807,N_36677);
and U48628 (N_48628,N_35138,N_30714);
and U48629 (N_48629,N_33153,N_31919);
nand U48630 (N_48630,N_38273,N_31369);
xnor U48631 (N_48631,N_34793,N_30686);
nor U48632 (N_48632,N_37868,N_35791);
nor U48633 (N_48633,N_31767,N_38158);
or U48634 (N_48634,N_32301,N_38648);
and U48635 (N_48635,N_32769,N_37651);
nand U48636 (N_48636,N_34895,N_30426);
nor U48637 (N_48637,N_32767,N_37843);
or U48638 (N_48638,N_37626,N_30488);
and U48639 (N_48639,N_34493,N_38504);
xnor U48640 (N_48640,N_36769,N_38539);
nor U48641 (N_48641,N_30076,N_33012);
nand U48642 (N_48642,N_32410,N_33911);
or U48643 (N_48643,N_37978,N_34608);
and U48644 (N_48644,N_30099,N_36657);
or U48645 (N_48645,N_34779,N_33749);
xnor U48646 (N_48646,N_39617,N_33477);
and U48647 (N_48647,N_33244,N_32300);
nand U48648 (N_48648,N_37958,N_34159);
and U48649 (N_48649,N_31765,N_30363);
nand U48650 (N_48650,N_32758,N_39374);
nand U48651 (N_48651,N_31887,N_34202);
nand U48652 (N_48652,N_33003,N_31132);
nor U48653 (N_48653,N_31416,N_33553);
and U48654 (N_48654,N_35692,N_37042);
nand U48655 (N_48655,N_30463,N_39525);
and U48656 (N_48656,N_32398,N_31728);
and U48657 (N_48657,N_30390,N_30492);
or U48658 (N_48658,N_31628,N_31693);
or U48659 (N_48659,N_33607,N_38759);
and U48660 (N_48660,N_33743,N_30002);
or U48661 (N_48661,N_37244,N_37380);
nand U48662 (N_48662,N_33005,N_35872);
or U48663 (N_48663,N_37110,N_37920);
or U48664 (N_48664,N_35760,N_37478);
nor U48665 (N_48665,N_33599,N_39443);
nand U48666 (N_48666,N_39131,N_32600);
and U48667 (N_48667,N_34128,N_38194);
or U48668 (N_48668,N_36174,N_32281);
and U48669 (N_48669,N_35175,N_32148);
nor U48670 (N_48670,N_31376,N_39904);
or U48671 (N_48671,N_38008,N_33424);
nand U48672 (N_48672,N_30492,N_32409);
xor U48673 (N_48673,N_33017,N_36563);
nand U48674 (N_48674,N_32539,N_30492);
and U48675 (N_48675,N_30264,N_31909);
and U48676 (N_48676,N_31527,N_33623);
xnor U48677 (N_48677,N_39105,N_38971);
and U48678 (N_48678,N_32846,N_38490);
xor U48679 (N_48679,N_33649,N_33422);
or U48680 (N_48680,N_30882,N_35097);
nor U48681 (N_48681,N_34346,N_31464);
nand U48682 (N_48682,N_33254,N_30677);
nor U48683 (N_48683,N_36259,N_30927);
nor U48684 (N_48684,N_33345,N_37263);
nor U48685 (N_48685,N_34078,N_35387);
nor U48686 (N_48686,N_31204,N_31894);
xor U48687 (N_48687,N_38420,N_33667);
and U48688 (N_48688,N_39071,N_36394);
or U48689 (N_48689,N_38235,N_34233);
or U48690 (N_48690,N_36781,N_33580);
and U48691 (N_48691,N_32794,N_39155);
nor U48692 (N_48692,N_37342,N_32510);
nand U48693 (N_48693,N_32073,N_37955);
nand U48694 (N_48694,N_38502,N_31876);
nor U48695 (N_48695,N_33271,N_33921);
nor U48696 (N_48696,N_38272,N_30889);
nand U48697 (N_48697,N_33429,N_38508);
xnor U48698 (N_48698,N_35140,N_31477);
nor U48699 (N_48699,N_30684,N_39246);
nand U48700 (N_48700,N_38875,N_35640);
nor U48701 (N_48701,N_36018,N_34081);
and U48702 (N_48702,N_39600,N_39460);
or U48703 (N_48703,N_32566,N_38409);
nand U48704 (N_48704,N_32265,N_35185);
nor U48705 (N_48705,N_37339,N_31395);
and U48706 (N_48706,N_36708,N_35434);
or U48707 (N_48707,N_38776,N_33840);
nor U48708 (N_48708,N_31530,N_30427);
and U48709 (N_48709,N_33546,N_34604);
and U48710 (N_48710,N_33918,N_39514);
or U48711 (N_48711,N_39000,N_37881);
or U48712 (N_48712,N_39032,N_33081);
and U48713 (N_48713,N_39178,N_38795);
or U48714 (N_48714,N_36866,N_35348);
and U48715 (N_48715,N_39686,N_30731);
xor U48716 (N_48716,N_37711,N_34955);
nor U48717 (N_48717,N_35767,N_34037);
and U48718 (N_48718,N_35495,N_36478);
and U48719 (N_48719,N_32388,N_39665);
nor U48720 (N_48720,N_39640,N_34743);
nor U48721 (N_48721,N_32679,N_36146);
xor U48722 (N_48722,N_38396,N_30295);
or U48723 (N_48723,N_33088,N_38069);
nor U48724 (N_48724,N_33797,N_38492);
or U48725 (N_48725,N_33163,N_36660);
nor U48726 (N_48726,N_32237,N_31322);
or U48727 (N_48727,N_30254,N_37830);
or U48728 (N_48728,N_33377,N_34895);
and U48729 (N_48729,N_39059,N_38001);
or U48730 (N_48730,N_32836,N_37116);
nor U48731 (N_48731,N_39613,N_38064);
xnor U48732 (N_48732,N_34407,N_36146);
or U48733 (N_48733,N_31859,N_35954);
nand U48734 (N_48734,N_34631,N_36637);
and U48735 (N_48735,N_32991,N_34023);
xor U48736 (N_48736,N_38547,N_38944);
xor U48737 (N_48737,N_31780,N_36996);
xnor U48738 (N_48738,N_36798,N_38173);
and U48739 (N_48739,N_35705,N_36457);
or U48740 (N_48740,N_36491,N_39959);
and U48741 (N_48741,N_35433,N_36504);
nor U48742 (N_48742,N_32454,N_35753);
or U48743 (N_48743,N_38600,N_39424);
nand U48744 (N_48744,N_38208,N_38102);
or U48745 (N_48745,N_31228,N_36793);
xor U48746 (N_48746,N_38099,N_33257);
nand U48747 (N_48747,N_31284,N_36769);
nor U48748 (N_48748,N_32048,N_37953);
and U48749 (N_48749,N_36490,N_39457);
nand U48750 (N_48750,N_30534,N_34176);
and U48751 (N_48751,N_36533,N_30981);
xor U48752 (N_48752,N_36068,N_33363);
nor U48753 (N_48753,N_35028,N_31828);
nor U48754 (N_48754,N_31165,N_39589);
nand U48755 (N_48755,N_35403,N_39551);
or U48756 (N_48756,N_33939,N_37127);
nor U48757 (N_48757,N_34518,N_30973);
or U48758 (N_48758,N_39113,N_32021);
and U48759 (N_48759,N_39007,N_30434);
and U48760 (N_48760,N_32560,N_32520);
nor U48761 (N_48761,N_31993,N_37023);
nor U48762 (N_48762,N_39461,N_32330);
and U48763 (N_48763,N_35135,N_31610);
and U48764 (N_48764,N_36019,N_30009);
nand U48765 (N_48765,N_37328,N_32739);
nand U48766 (N_48766,N_38850,N_37752);
xnor U48767 (N_48767,N_33922,N_36563);
nor U48768 (N_48768,N_32392,N_32975);
nor U48769 (N_48769,N_33720,N_30067);
and U48770 (N_48770,N_39661,N_39494);
or U48771 (N_48771,N_32157,N_32685);
nand U48772 (N_48772,N_31259,N_39855);
nand U48773 (N_48773,N_33836,N_34495);
nand U48774 (N_48774,N_33290,N_31704);
xor U48775 (N_48775,N_37381,N_37808);
and U48776 (N_48776,N_36491,N_36190);
nand U48777 (N_48777,N_30120,N_31047);
nand U48778 (N_48778,N_31683,N_33604);
or U48779 (N_48779,N_39293,N_35192);
nor U48780 (N_48780,N_31542,N_38762);
or U48781 (N_48781,N_36582,N_38076);
nand U48782 (N_48782,N_31893,N_31874);
and U48783 (N_48783,N_33980,N_34605);
or U48784 (N_48784,N_35938,N_33991);
and U48785 (N_48785,N_30654,N_34830);
or U48786 (N_48786,N_37216,N_38582);
nand U48787 (N_48787,N_36984,N_31111);
and U48788 (N_48788,N_37113,N_31463);
or U48789 (N_48789,N_38898,N_38140);
nor U48790 (N_48790,N_32016,N_30645);
xor U48791 (N_48791,N_38721,N_39966);
xnor U48792 (N_48792,N_33916,N_39321);
nand U48793 (N_48793,N_31761,N_37169);
and U48794 (N_48794,N_36295,N_37007);
nand U48795 (N_48795,N_38246,N_35398);
and U48796 (N_48796,N_36163,N_39394);
and U48797 (N_48797,N_33587,N_34254);
or U48798 (N_48798,N_37164,N_39594);
nor U48799 (N_48799,N_37419,N_31780);
nor U48800 (N_48800,N_36530,N_30108);
nand U48801 (N_48801,N_30727,N_30875);
nor U48802 (N_48802,N_32739,N_35943);
or U48803 (N_48803,N_31235,N_33277);
and U48804 (N_48804,N_38889,N_36620);
nor U48805 (N_48805,N_38819,N_35427);
and U48806 (N_48806,N_37770,N_30257);
or U48807 (N_48807,N_39234,N_32215);
nor U48808 (N_48808,N_34883,N_39857);
nor U48809 (N_48809,N_38427,N_37759);
nand U48810 (N_48810,N_38494,N_30560);
or U48811 (N_48811,N_30853,N_38943);
nor U48812 (N_48812,N_34532,N_35349);
or U48813 (N_48813,N_35207,N_37125);
xor U48814 (N_48814,N_34384,N_39229);
nand U48815 (N_48815,N_33672,N_39731);
and U48816 (N_48816,N_30516,N_38381);
or U48817 (N_48817,N_38482,N_34682);
nand U48818 (N_48818,N_32176,N_39741);
xnor U48819 (N_48819,N_34982,N_33837);
nor U48820 (N_48820,N_32717,N_36922);
nor U48821 (N_48821,N_32552,N_32693);
and U48822 (N_48822,N_34505,N_33326);
nand U48823 (N_48823,N_38242,N_38060);
or U48824 (N_48824,N_34633,N_31936);
nand U48825 (N_48825,N_33727,N_39688);
or U48826 (N_48826,N_37565,N_39091);
and U48827 (N_48827,N_31732,N_35735);
nand U48828 (N_48828,N_39454,N_32105);
or U48829 (N_48829,N_36822,N_31275);
and U48830 (N_48830,N_39984,N_37912);
xor U48831 (N_48831,N_34869,N_37917);
nand U48832 (N_48832,N_34544,N_32033);
and U48833 (N_48833,N_39519,N_33140);
nor U48834 (N_48834,N_38777,N_38389);
and U48835 (N_48835,N_30489,N_35028);
or U48836 (N_48836,N_37911,N_36105);
xor U48837 (N_48837,N_38664,N_33359);
and U48838 (N_48838,N_37592,N_37452);
xor U48839 (N_48839,N_32065,N_31478);
xor U48840 (N_48840,N_34085,N_34982);
nand U48841 (N_48841,N_30840,N_39214);
nor U48842 (N_48842,N_38092,N_38839);
or U48843 (N_48843,N_30926,N_35303);
and U48844 (N_48844,N_35094,N_38731);
or U48845 (N_48845,N_37955,N_36419);
nand U48846 (N_48846,N_34512,N_30013);
nand U48847 (N_48847,N_36780,N_38830);
xor U48848 (N_48848,N_32564,N_33021);
xnor U48849 (N_48849,N_39639,N_39050);
nor U48850 (N_48850,N_39929,N_32805);
nand U48851 (N_48851,N_33600,N_30389);
nand U48852 (N_48852,N_39137,N_32013);
nand U48853 (N_48853,N_35945,N_37440);
xnor U48854 (N_48854,N_38388,N_39939);
and U48855 (N_48855,N_32468,N_32626);
or U48856 (N_48856,N_33775,N_30691);
xor U48857 (N_48857,N_33489,N_34361);
nand U48858 (N_48858,N_33083,N_38190);
xnor U48859 (N_48859,N_37197,N_38938);
nand U48860 (N_48860,N_30372,N_38216);
or U48861 (N_48861,N_36055,N_33172);
or U48862 (N_48862,N_36240,N_33383);
nor U48863 (N_48863,N_35835,N_34746);
or U48864 (N_48864,N_37009,N_30121);
and U48865 (N_48865,N_38174,N_37673);
nor U48866 (N_48866,N_31464,N_32964);
nor U48867 (N_48867,N_34109,N_34071);
nor U48868 (N_48868,N_36694,N_37130);
and U48869 (N_48869,N_35115,N_37817);
or U48870 (N_48870,N_36107,N_34948);
or U48871 (N_48871,N_39647,N_32849);
and U48872 (N_48872,N_37853,N_37893);
xnor U48873 (N_48873,N_31679,N_36997);
nor U48874 (N_48874,N_36891,N_36822);
nand U48875 (N_48875,N_34585,N_39650);
and U48876 (N_48876,N_34172,N_31240);
and U48877 (N_48877,N_33487,N_30658);
and U48878 (N_48878,N_31165,N_31470);
xnor U48879 (N_48879,N_36591,N_34314);
xnor U48880 (N_48880,N_31425,N_35624);
or U48881 (N_48881,N_39528,N_38763);
or U48882 (N_48882,N_39986,N_38987);
and U48883 (N_48883,N_37300,N_37674);
or U48884 (N_48884,N_35357,N_37487);
nand U48885 (N_48885,N_35457,N_31570);
nor U48886 (N_48886,N_36862,N_33101);
or U48887 (N_48887,N_38708,N_32339);
xor U48888 (N_48888,N_31199,N_32155);
or U48889 (N_48889,N_39963,N_33080);
nand U48890 (N_48890,N_38118,N_37143);
nand U48891 (N_48891,N_30850,N_37804);
nor U48892 (N_48892,N_35153,N_31779);
nor U48893 (N_48893,N_35293,N_34407);
or U48894 (N_48894,N_35293,N_38385);
xor U48895 (N_48895,N_37890,N_38219);
nor U48896 (N_48896,N_33221,N_34828);
and U48897 (N_48897,N_30372,N_36182);
or U48898 (N_48898,N_33288,N_39462);
nor U48899 (N_48899,N_36811,N_32166);
and U48900 (N_48900,N_30161,N_35567);
and U48901 (N_48901,N_33663,N_38888);
nor U48902 (N_48902,N_39014,N_30301);
nor U48903 (N_48903,N_38588,N_33065);
nor U48904 (N_48904,N_35181,N_31956);
nor U48905 (N_48905,N_32708,N_33340);
nor U48906 (N_48906,N_33570,N_32078);
nor U48907 (N_48907,N_39040,N_32091);
and U48908 (N_48908,N_31243,N_37806);
and U48909 (N_48909,N_39791,N_30758);
xor U48910 (N_48910,N_32253,N_35532);
or U48911 (N_48911,N_34127,N_38609);
and U48912 (N_48912,N_30523,N_39226);
nor U48913 (N_48913,N_31317,N_37429);
nand U48914 (N_48914,N_35222,N_38706);
or U48915 (N_48915,N_30830,N_33371);
nand U48916 (N_48916,N_37135,N_34520);
or U48917 (N_48917,N_38283,N_36935);
nor U48918 (N_48918,N_30944,N_32786);
or U48919 (N_48919,N_30790,N_33674);
nand U48920 (N_48920,N_39888,N_32740);
nor U48921 (N_48921,N_35222,N_32459);
or U48922 (N_48922,N_35304,N_30419);
nor U48923 (N_48923,N_38781,N_38506);
nand U48924 (N_48924,N_39529,N_34628);
xor U48925 (N_48925,N_39443,N_34480);
and U48926 (N_48926,N_39662,N_30683);
or U48927 (N_48927,N_31954,N_33788);
and U48928 (N_48928,N_34939,N_36649);
nor U48929 (N_48929,N_32007,N_35922);
and U48930 (N_48930,N_37231,N_38872);
xor U48931 (N_48931,N_36286,N_36067);
nand U48932 (N_48932,N_30588,N_31709);
nor U48933 (N_48933,N_32613,N_30312);
nand U48934 (N_48934,N_32223,N_36331);
nand U48935 (N_48935,N_38189,N_37364);
nand U48936 (N_48936,N_31641,N_38855);
nor U48937 (N_48937,N_34897,N_36512);
nor U48938 (N_48938,N_32840,N_37615);
xor U48939 (N_48939,N_31961,N_35800);
or U48940 (N_48940,N_34460,N_33874);
xor U48941 (N_48941,N_32933,N_36081);
xnor U48942 (N_48942,N_30950,N_30066);
xnor U48943 (N_48943,N_37764,N_37802);
nor U48944 (N_48944,N_31777,N_32278);
and U48945 (N_48945,N_38695,N_35051);
or U48946 (N_48946,N_35478,N_33641);
nand U48947 (N_48947,N_38710,N_32792);
nand U48948 (N_48948,N_37110,N_31457);
nor U48949 (N_48949,N_30257,N_37662);
nand U48950 (N_48950,N_39487,N_35607);
nor U48951 (N_48951,N_30442,N_31429);
or U48952 (N_48952,N_39210,N_33489);
or U48953 (N_48953,N_32667,N_35005);
and U48954 (N_48954,N_32754,N_33984);
nand U48955 (N_48955,N_37763,N_33320);
nand U48956 (N_48956,N_32568,N_31790);
nor U48957 (N_48957,N_39066,N_37614);
nand U48958 (N_48958,N_37760,N_39885);
or U48959 (N_48959,N_31669,N_34560);
and U48960 (N_48960,N_38508,N_38252);
nor U48961 (N_48961,N_39223,N_30251);
xnor U48962 (N_48962,N_37094,N_32071);
nor U48963 (N_48963,N_30347,N_30344);
nor U48964 (N_48964,N_36717,N_34676);
and U48965 (N_48965,N_37862,N_33741);
or U48966 (N_48966,N_39460,N_31676);
nor U48967 (N_48967,N_35013,N_30752);
or U48968 (N_48968,N_38083,N_38210);
xor U48969 (N_48969,N_32735,N_34571);
nand U48970 (N_48970,N_39168,N_37085);
or U48971 (N_48971,N_30100,N_35669);
and U48972 (N_48972,N_31680,N_34021);
nor U48973 (N_48973,N_33550,N_33370);
nor U48974 (N_48974,N_33716,N_32203);
and U48975 (N_48975,N_37293,N_32855);
nand U48976 (N_48976,N_39679,N_38323);
nand U48977 (N_48977,N_37198,N_32927);
or U48978 (N_48978,N_34806,N_31407);
and U48979 (N_48979,N_38060,N_33696);
or U48980 (N_48980,N_30476,N_32246);
nor U48981 (N_48981,N_31724,N_32923);
nand U48982 (N_48982,N_33493,N_37911);
xor U48983 (N_48983,N_32691,N_38946);
and U48984 (N_48984,N_31639,N_36297);
nor U48985 (N_48985,N_36285,N_37126);
nand U48986 (N_48986,N_33308,N_31342);
nor U48987 (N_48987,N_31431,N_30997);
nand U48988 (N_48988,N_34941,N_30984);
or U48989 (N_48989,N_30070,N_36052);
nand U48990 (N_48990,N_38798,N_32863);
nand U48991 (N_48991,N_31323,N_38841);
and U48992 (N_48992,N_32461,N_34809);
and U48993 (N_48993,N_30517,N_37536);
and U48994 (N_48994,N_30812,N_35292);
and U48995 (N_48995,N_33207,N_37562);
or U48996 (N_48996,N_39113,N_33238);
or U48997 (N_48997,N_33807,N_31061);
or U48998 (N_48998,N_32568,N_35024);
nand U48999 (N_48999,N_32878,N_33992);
nand U49000 (N_49000,N_38593,N_35999);
or U49001 (N_49001,N_31491,N_36084);
nor U49002 (N_49002,N_36679,N_36508);
and U49003 (N_49003,N_35376,N_38764);
and U49004 (N_49004,N_37786,N_34855);
nand U49005 (N_49005,N_35565,N_31004);
and U49006 (N_49006,N_38361,N_33442);
xor U49007 (N_49007,N_36204,N_30359);
and U49008 (N_49008,N_33233,N_39173);
and U49009 (N_49009,N_32971,N_38397);
xnor U49010 (N_49010,N_30267,N_34453);
xnor U49011 (N_49011,N_35734,N_33721);
nor U49012 (N_49012,N_35911,N_30528);
nor U49013 (N_49013,N_33232,N_37365);
nor U49014 (N_49014,N_37599,N_30439);
nand U49015 (N_49015,N_32721,N_39869);
xor U49016 (N_49016,N_33152,N_31006);
and U49017 (N_49017,N_31128,N_38855);
or U49018 (N_49018,N_33097,N_37333);
or U49019 (N_49019,N_39073,N_39650);
and U49020 (N_49020,N_39772,N_30203);
nand U49021 (N_49021,N_33354,N_33363);
nand U49022 (N_49022,N_39222,N_39759);
or U49023 (N_49023,N_38957,N_36859);
or U49024 (N_49024,N_36156,N_30905);
xor U49025 (N_49025,N_31228,N_33169);
and U49026 (N_49026,N_38337,N_33118);
or U49027 (N_49027,N_38552,N_38106);
nor U49028 (N_49028,N_33018,N_35222);
nand U49029 (N_49029,N_30197,N_35742);
nor U49030 (N_49030,N_32826,N_34219);
nand U49031 (N_49031,N_31462,N_39482);
and U49032 (N_49032,N_31196,N_35916);
xor U49033 (N_49033,N_38160,N_36652);
nand U49034 (N_49034,N_38583,N_36105);
nor U49035 (N_49035,N_33360,N_36080);
nand U49036 (N_49036,N_30368,N_36412);
or U49037 (N_49037,N_32129,N_30870);
and U49038 (N_49038,N_35288,N_37473);
or U49039 (N_49039,N_39681,N_30372);
and U49040 (N_49040,N_35565,N_38412);
or U49041 (N_49041,N_36503,N_30259);
xor U49042 (N_49042,N_34914,N_30410);
nor U49043 (N_49043,N_32746,N_33780);
and U49044 (N_49044,N_35045,N_36563);
and U49045 (N_49045,N_35146,N_39205);
nand U49046 (N_49046,N_32536,N_37425);
or U49047 (N_49047,N_36741,N_38222);
nand U49048 (N_49048,N_39148,N_39372);
or U49049 (N_49049,N_37336,N_38061);
or U49050 (N_49050,N_36482,N_30119);
nor U49051 (N_49051,N_39261,N_30061);
or U49052 (N_49052,N_31595,N_30862);
xnor U49053 (N_49053,N_38973,N_35119);
or U49054 (N_49054,N_30119,N_37680);
and U49055 (N_49055,N_34367,N_34193);
and U49056 (N_49056,N_30605,N_34076);
xnor U49057 (N_49057,N_39944,N_31158);
or U49058 (N_49058,N_34091,N_37724);
nand U49059 (N_49059,N_30349,N_32167);
xnor U49060 (N_49060,N_33518,N_34880);
xor U49061 (N_49061,N_35190,N_30414);
nor U49062 (N_49062,N_35802,N_31271);
nand U49063 (N_49063,N_39611,N_36469);
and U49064 (N_49064,N_30223,N_37170);
nand U49065 (N_49065,N_30900,N_34147);
or U49066 (N_49066,N_31366,N_31368);
nand U49067 (N_49067,N_31897,N_38416);
and U49068 (N_49068,N_34102,N_31512);
xor U49069 (N_49069,N_33141,N_36093);
nor U49070 (N_49070,N_39682,N_37762);
and U49071 (N_49071,N_35985,N_32017);
and U49072 (N_49072,N_36001,N_37315);
nand U49073 (N_49073,N_30500,N_32332);
nand U49074 (N_49074,N_36439,N_34104);
nand U49075 (N_49075,N_39511,N_39505);
and U49076 (N_49076,N_39809,N_30244);
nor U49077 (N_49077,N_38032,N_31754);
nor U49078 (N_49078,N_39726,N_31280);
nor U49079 (N_49079,N_33704,N_35614);
xor U49080 (N_49080,N_36980,N_36541);
and U49081 (N_49081,N_30654,N_34175);
or U49082 (N_49082,N_34793,N_39155);
nand U49083 (N_49083,N_34213,N_31713);
or U49084 (N_49084,N_31296,N_34328);
and U49085 (N_49085,N_30489,N_36065);
nand U49086 (N_49086,N_31044,N_30200);
and U49087 (N_49087,N_31169,N_35645);
and U49088 (N_49088,N_35101,N_38141);
nor U49089 (N_49089,N_31653,N_31216);
and U49090 (N_49090,N_30908,N_31347);
xor U49091 (N_49091,N_32972,N_36644);
and U49092 (N_49092,N_37689,N_33827);
and U49093 (N_49093,N_36699,N_37773);
nor U49094 (N_49094,N_39255,N_35423);
and U49095 (N_49095,N_34047,N_30109);
nor U49096 (N_49096,N_31200,N_35781);
or U49097 (N_49097,N_39967,N_30449);
nor U49098 (N_49098,N_31725,N_37437);
nor U49099 (N_49099,N_30542,N_31653);
xor U49100 (N_49100,N_32583,N_36167);
and U49101 (N_49101,N_30839,N_38148);
nor U49102 (N_49102,N_39149,N_33085);
nand U49103 (N_49103,N_30268,N_35502);
nor U49104 (N_49104,N_36142,N_30619);
xor U49105 (N_49105,N_30326,N_38150);
and U49106 (N_49106,N_32702,N_35065);
nand U49107 (N_49107,N_34262,N_31944);
nor U49108 (N_49108,N_34252,N_37998);
nor U49109 (N_49109,N_34207,N_33894);
nand U49110 (N_49110,N_32915,N_31111);
or U49111 (N_49111,N_31383,N_32001);
nand U49112 (N_49112,N_36530,N_38946);
nand U49113 (N_49113,N_31026,N_36098);
and U49114 (N_49114,N_34968,N_39954);
nand U49115 (N_49115,N_30371,N_34923);
and U49116 (N_49116,N_34324,N_36989);
xor U49117 (N_49117,N_38664,N_36913);
nand U49118 (N_49118,N_34631,N_35872);
and U49119 (N_49119,N_35967,N_38152);
and U49120 (N_49120,N_33071,N_32642);
and U49121 (N_49121,N_32874,N_39468);
or U49122 (N_49122,N_35821,N_37544);
nand U49123 (N_49123,N_30793,N_36819);
or U49124 (N_49124,N_39612,N_36518);
nand U49125 (N_49125,N_31151,N_30434);
or U49126 (N_49126,N_39487,N_32992);
or U49127 (N_49127,N_36609,N_33814);
nor U49128 (N_49128,N_39558,N_36940);
nor U49129 (N_49129,N_39755,N_30308);
and U49130 (N_49130,N_35811,N_35854);
nand U49131 (N_49131,N_32918,N_33009);
and U49132 (N_49132,N_35116,N_33416);
nand U49133 (N_49133,N_38244,N_38680);
or U49134 (N_49134,N_32364,N_33201);
nor U49135 (N_49135,N_35963,N_37034);
and U49136 (N_49136,N_32611,N_35384);
or U49137 (N_49137,N_31293,N_36858);
and U49138 (N_49138,N_30207,N_32970);
and U49139 (N_49139,N_31697,N_38648);
and U49140 (N_49140,N_32878,N_38541);
nand U49141 (N_49141,N_36198,N_36509);
and U49142 (N_49142,N_37007,N_36216);
nand U49143 (N_49143,N_31814,N_34530);
nor U49144 (N_49144,N_36219,N_31876);
nand U49145 (N_49145,N_32135,N_30222);
nand U49146 (N_49146,N_34676,N_35181);
and U49147 (N_49147,N_33896,N_33573);
nand U49148 (N_49148,N_38186,N_39775);
and U49149 (N_49149,N_30800,N_37362);
and U49150 (N_49150,N_35760,N_38506);
and U49151 (N_49151,N_32586,N_39097);
or U49152 (N_49152,N_36782,N_35416);
nand U49153 (N_49153,N_30404,N_33974);
xnor U49154 (N_49154,N_35255,N_33703);
nand U49155 (N_49155,N_36269,N_35126);
and U49156 (N_49156,N_32635,N_33412);
nor U49157 (N_49157,N_30405,N_30996);
and U49158 (N_49158,N_32916,N_38019);
nor U49159 (N_49159,N_37918,N_32885);
nor U49160 (N_49160,N_37958,N_35615);
nor U49161 (N_49161,N_31230,N_36802);
nand U49162 (N_49162,N_32350,N_37445);
nand U49163 (N_49163,N_32106,N_31514);
and U49164 (N_49164,N_34516,N_31076);
or U49165 (N_49165,N_34386,N_34059);
nand U49166 (N_49166,N_36481,N_34586);
nor U49167 (N_49167,N_32440,N_37936);
nand U49168 (N_49168,N_35279,N_31308);
and U49169 (N_49169,N_38327,N_32373);
nand U49170 (N_49170,N_32411,N_37208);
nor U49171 (N_49171,N_31402,N_33602);
nand U49172 (N_49172,N_37791,N_39430);
xnor U49173 (N_49173,N_31866,N_34960);
nand U49174 (N_49174,N_31050,N_31179);
and U49175 (N_49175,N_31464,N_30170);
nand U49176 (N_49176,N_33213,N_32690);
or U49177 (N_49177,N_33638,N_31708);
nand U49178 (N_49178,N_37919,N_32212);
nand U49179 (N_49179,N_39541,N_33139);
nand U49180 (N_49180,N_33072,N_34438);
and U49181 (N_49181,N_34894,N_35014);
or U49182 (N_49182,N_35266,N_33823);
nor U49183 (N_49183,N_38996,N_36582);
and U49184 (N_49184,N_38594,N_32684);
and U49185 (N_49185,N_38555,N_32072);
or U49186 (N_49186,N_39164,N_34913);
nor U49187 (N_49187,N_31789,N_39212);
nor U49188 (N_49188,N_36762,N_33606);
and U49189 (N_49189,N_31380,N_30786);
nand U49190 (N_49190,N_36758,N_39242);
or U49191 (N_49191,N_39334,N_38056);
or U49192 (N_49192,N_35016,N_36439);
nor U49193 (N_49193,N_36740,N_33365);
and U49194 (N_49194,N_34501,N_33013);
nor U49195 (N_49195,N_32341,N_31523);
nand U49196 (N_49196,N_30215,N_37617);
or U49197 (N_49197,N_34314,N_39178);
or U49198 (N_49198,N_30637,N_36486);
or U49199 (N_49199,N_33971,N_31554);
xnor U49200 (N_49200,N_33134,N_34723);
nand U49201 (N_49201,N_36513,N_37432);
nor U49202 (N_49202,N_36962,N_31869);
and U49203 (N_49203,N_37792,N_39574);
and U49204 (N_49204,N_32136,N_38464);
nand U49205 (N_49205,N_37522,N_38115);
nor U49206 (N_49206,N_38623,N_32802);
or U49207 (N_49207,N_35307,N_32401);
nor U49208 (N_49208,N_31980,N_34167);
and U49209 (N_49209,N_31960,N_39526);
xor U49210 (N_49210,N_31882,N_34474);
or U49211 (N_49211,N_35626,N_33954);
and U49212 (N_49212,N_32660,N_39331);
and U49213 (N_49213,N_36321,N_35126);
or U49214 (N_49214,N_30678,N_32040);
or U49215 (N_49215,N_36676,N_33317);
nand U49216 (N_49216,N_32167,N_34843);
nor U49217 (N_49217,N_34635,N_30869);
and U49218 (N_49218,N_34574,N_30373);
or U49219 (N_49219,N_39637,N_36263);
and U49220 (N_49220,N_39128,N_31122);
xnor U49221 (N_49221,N_31223,N_35755);
or U49222 (N_49222,N_37453,N_38081);
or U49223 (N_49223,N_38949,N_34087);
nand U49224 (N_49224,N_30290,N_33142);
and U49225 (N_49225,N_37632,N_36916);
nand U49226 (N_49226,N_37135,N_34937);
nand U49227 (N_49227,N_36584,N_39186);
nor U49228 (N_49228,N_38707,N_33707);
nand U49229 (N_49229,N_35373,N_37366);
nor U49230 (N_49230,N_33210,N_39067);
nand U49231 (N_49231,N_38352,N_31485);
or U49232 (N_49232,N_30755,N_31706);
nor U49233 (N_49233,N_30641,N_34948);
nor U49234 (N_49234,N_36010,N_31832);
and U49235 (N_49235,N_38465,N_34718);
and U49236 (N_49236,N_38777,N_35311);
nor U49237 (N_49237,N_34592,N_35119);
and U49238 (N_49238,N_34058,N_38722);
nand U49239 (N_49239,N_33869,N_31607);
nand U49240 (N_49240,N_32892,N_31666);
nand U49241 (N_49241,N_37983,N_31982);
and U49242 (N_49242,N_34388,N_37782);
nand U49243 (N_49243,N_32179,N_39502);
or U49244 (N_49244,N_34213,N_32871);
xnor U49245 (N_49245,N_31898,N_35142);
and U49246 (N_49246,N_39643,N_32657);
or U49247 (N_49247,N_38894,N_31571);
or U49248 (N_49248,N_30264,N_36931);
and U49249 (N_49249,N_34110,N_33426);
and U49250 (N_49250,N_34044,N_39939);
nand U49251 (N_49251,N_32292,N_39038);
and U49252 (N_49252,N_35075,N_34395);
and U49253 (N_49253,N_35973,N_38222);
and U49254 (N_49254,N_32727,N_36509);
or U49255 (N_49255,N_38916,N_38782);
or U49256 (N_49256,N_31136,N_33582);
nor U49257 (N_49257,N_37267,N_37648);
xor U49258 (N_49258,N_34901,N_33281);
or U49259 (N_49259,N_35676,N_38879);
and U49260 (N_49260,N_30367,N_35615);
nand U49261 (N_49261,N_34601,N_36300);
nor U49262 (N_49262,N_30981,N_30952);
nand U49263 (N_49263,N_33725,N_39610);
nor U49264 (N_49264,N_35566,N_32892);
nor U49265 (N_49265,N_31183,N_33015);
xor U49266 (N_49266,N_32549,N_35659);
and U49267 (N_49267,N_36924,N_34359);
and U49268 (N_49268,N_35274,N_38754);
xor U49269 (N_49269,N_34408,N_38654);
nor U49270 (N_49270,N_35143,N_34837);
xor U49271 (N_49271,N_39585,N_31977);
nand U49272 (N_49272,N_36396,N_36157);
nor U49273 (N_49273,N_36750,N_37522);
or U49274 (N_49274,N_30472,N_38258);
nor U49275 (N_49275,N_34135,N_31781);
or U49276 (N_49276,N_39270,N_34159);
nor U49277 (N_49277,N_37101,N_37096);
and U49278 (N_49278,N_32143,N_37416);
xor U49279 (N_49279,N_31965,N_36364);
or U49280 (N_49280,N_30192,N_32613);
or U49281 (N_49281,N_31181,N_39780);
or U49282 (N_49282,N_37620,N_32806);
xor U49283 (N_49283,N_31660,N_33732);
and U49284 (N_49284,N_39518,N_39552);
xor U49285 (N_49285,N_36867,N_32833);
nand U49286 (N_49286,N_38221,N_30767);
and U49287 (N_49287,N_36299,N_32249);
nor U49288 (N_49288,N_30536,N_39364);
xor U49289 (N_49289,N_32014,N_35696);
nand U49290 (N_49290,N_30702,N_33959);
and U49291 (N_49291,N_31620,N_39719);
and U49292 (N_49292,N_30695,N_37005);
and U49293 (N_49293,N_37081,N_30028);
and U49294 (N_49294,N_39274,N_32369);
nor U49295 (N_49295,N_35593,N_34894);
nor U49296 (N_49296,N_34832,N_38990);
nand U49297 (N_49297,N_32993,N_35052);
or U49298 (N_49298,N_30190,N_36574);
and U49299 (N_49299,N_38766,N_36268);
nand U49300 (N_49300,N_30932,N_37645);
nand U49301 (N_49301,N_34309,N_30149);
and U49302 (N_49302,N_36899,N_33215);
or U49303 (N_49303,N_32678,N_32259);
nor U49304 (N_49304,N_31545,N_38774);
xnor U49305 (N_49305,N_34650,N_31294);
and U49306 (N_49306,N_36700,N_32822);
and U49307 (N_49307,N_35438,N_30746);
and U49308 (N_49308,N_32185,N_36116);
nand U49309 (N_49309,N_39900,N_36560);
or U49310 (N_49310,N_30693,N_37550);
nor U49311 (N_49311,N_33245,N_39580);
nor U49312 (N_49312,N_39108,N_37202);
nor U49313 (N_49313,N_35487,N_32731);
nand U49314 (N_49314,N_32124,N_33321);
nor U49315 (N_49315,N_35802,N_38256);
and U49316 (N_49316,N_36178,N_32194);
nand U49317 (N_49317,N_32719,N_33369);
and U49318 (N_49318,N_32544,N_38997);
nor U49319 (N_49319,N_30897,N_34717);
xnor U49320 (N_49320,N_33041,N_30741);
and U49321 (N_49321,N_35005,N_35938);
nand U49322 (N_49322,N_36600,N_35856);
nor U49323 (N_49323,N_34877,N_36340);
xnor U49324 (N_49324,N_33922,N_32298);
or U49325 (N_49325,N_31566,N_36882);
xor U49326 (N_49326,N_36104,N_35533);
or U49327 (N_49327,N_39275,N_35352);
nand U49328 (N_49328,N_35736,N_37020);
nand U49329 (N_49329,N_37010,N_33526);
nand U49330 (N_49330,N_31168,N_37551);
and U49331 (N_49331,N_39170,N_39807);
nor U49332 (N_49332,N_39136,N_38560);
nor U49333 (N_49333,N_39307,N_38644);
or U49334 (N_49334,N_36551,N_39820);
nor U49335 (N_49335,N_31125,N_35066);
xor U49336 (N_49336,N_39692,N_31632);
or U49337 (N_49337,N_36482,N_34011);
nor U49338 (N_49338,N_33827,N_30861);
or U49339 (N_49339,N_31770,N_33996);
or U49340 (N_49340,N_34786,N_32200);
nor U49341 (N_49341,N_35795,N_31996);
nor U49342 (N_49342,N_31111,N_32188);
and U49343 (N_49343,N_35246,N_38460);
nor U49344 (N_49344,N_33938,N_37098);
xor U49345 (N_49345,N_39878,N_30759);
and U49346 (N_49346,N_36197,N_30998);
or U49347 (N_49347,N_39821,N_35893);
or U49348 (N_49348,N_36064,N_37167);
xnor U49349 (N_49349,N_33605,N_34951);
nand U49350 (N_49350,N_35294,N_31310);
nor U49351 (N_49351,N_38262,N_30965);
nand U49352 (N_49352,N_33778,N_31623);
or U49353 (N_49353,N_36696,N_38238);
nor U49354 (N_49354,N_33914,N_39440);
or U49355 (N_49355,N_37718,N_36066);
xor U49356 (N_49356,N_37574,N_39547);
and U49357 (N_49357,N_38086,N_39127);
or U49358 (N_49358,N_38953,N_36284);
nand U49359 (N_49359,N_36781,N_32414);
and U49360 (N_49360,N_34403,N_37661);
or U49361 (N_49361,N_38583,N_35503);
and U49362 (N_49362,N_30094,N_39016);
nand U49363 (N_49363,N_30610,N_36497);
xor U49364 (N_49364,N_31071,N_32133);
or U49365 (N_49365,N_38955,N_32455);
nor U49366 (N_49366,N_31853,N_31049);
nor U49367 (N_49367,N_35846,N_37207);
nor U49368 (N_49368,N_31943,N_36133);
and U49369 (N_49369,N_35829,N_36187);
nand U49370 (N_49370,N_34096,N_30551);
or U49371 (N_49371,N_30717,N_34358);
and U49372 (N_49372,N_33453,N_36365);
and U49373 (N_49373,N_34059,N_34912);
and U49374 (N_49374,N_32071,N_35327);
nand U49375 (N_49375,N_35587,N_30599);
and U49376 (N_49376,N_33844,N_39985);
and U49377 (N_49377,N_39667,N_34714);
and U49378 (N_49378,N_32253,N_37210);
nand U49379 (N_49379,N_35028,N_31400);
nand U49380 (N_49380,N_38649,N_35055);
xor U49381 (N_49381,N_34074,N_31623);
or U49382 (N_49382,N_37699,N_34538);
and U49383 (N_49383,N_39615,N_37830);
xor U49384 (N_49384,N_38202,N_39020);
or U49385 (N_49385,N_37206,N_32406);
nor U49386 (N_49386,N_37041,N_30121);
and U49387 (N_49387,N_35235,N_30938);
and U49388 (N_49388,N_35525,N_32378);
or U49389 (N_49389,N_35120,N_32312);
and U49390 (N_49390,N_37108,N_36640);
nand U49391 (N_49391,N_31174,N_34349);
or U49392 (N_49392,N_30677,N_39089);
nand U49393 (N_49393,N_39995,N_39282);
xnor U49394 (N_49394,N_30605,N_38836);
nor U49395 (N_49395,N_34453,N_31058);
and U49396 (N_49396,N_33799,N_36837);
nand U49397 (N_49397,N_39441,N_34324);
nand U49398 (N_49398,N_39818,N_33247);
or U49399 (N_49399,N_34648,N_35922);
and U49400 (N_49400,N_32191,N_39932);
nand U49401 (N_49401,N_33364,N_38828);
nand U49402 (N_49402,N_31617,N_31912);
nor U49403 (N_49403,N_30512,N_33271);
and U49404 (N_49404,N_31450,N_31110);
nor U49405 (N_49405,N_32342,N_38811);
xor U49406 (N_49406,N_36587,N_32688);
and U49407 (N_49407,N_38978,N_38378);
nand U49408 (N_49408,N_34574,N_38293);
nor U49409 (N_49409,N_37817,N_33987);
and U49410 (N_49410,N_39777,N_39212);
nor U49411 (N_49411,N_32414,N_35530);
nor U49412 (N_49412,N_37163,N_36274);
or U49413 (N_49413,N_31972,N_31176);
or U49414 (N_49414,N_32636,N_30614);
xnor U49415 (N_49415,N_33905,N_36645);
nand U49416 (N_49416,N_31364,N_36235);
xor U49417 (N_49417,N_37100,N_39185);
and U49418 (N_49418,N_37961,N_39904);
nand U49419 (N_49419,N_30085,N_36786);
and U49420 (N_49420,N_39318,N_32325);
xnor U49421 (N_49421,N_36619,N_33842);
and U49422 (N_49422,N_30083,N_33028);
and U49423 (N_49423,N_30474,N_33599);
nand U49424 (N_49424,N_38570,N_36523);
nor U49425 (N_49425,N_32415,N_37568);
nand U49426 (N_49426,N_31543,N_37859);
xnor U49427 (N_49427,N_33869,N_36884);
nor U49428 (N_49428,N_38357,N_32159);
nor U49429 (N_49429,N_38699,N_33090);
or U49430 (N_49430,N_31587,N_35538);
and U49431 (N_49431,N_38618,N_36634);
and U49432 (N_49432,N_30514,N_30052);
nor U49433 (N_49433,N_30733,N_33810);
and U49434 (N_49434,N_33178,N_34739);
nand U49435 (N_49435,N_38966,N_39638);
and U49436 (N_49436,N_31235,N_32319);
or U49437 (N_49437,N_38067,N_30562);
nand U49438 (N_49438,N_30490,N_33772);
nor U49439 (N_49439,N_37808,N_31639);
or U49440 (N_49440,N_33300,N_34321);
nor U49441 (N_49441,N_30907,N_38274);
nor U49442 (N_49442,N_33802,N_35848);
and U49443 (N_49443,N_31617,N_31613);
nor U49444 (N_49444,N_33251,N_36774);
xor U49445 (N_49445,N_39526,N_35782);
and U49446 (N_49446,N_33993,N_36262);
xnor U49447 (N_49447,N_38017,N_39008);
nor U49448 (N_49448,N_34616,N_35700);
or U49449 (N_49449,N_33475,N_36640);
nor U49450 (N_49450,N_33416,N_38385);
xor U49451 (N_49451,N_35416,N_36315);
nand U49452 (N_49452,N_38031,N_33228);
nor U49453 (N_49453,N_30769,N_33582);
and U49454 (N_49454,N_31669,N_31452);
or U49455 (N_49455,N_37825,N_33655);
nand U49456 (N_49456,N_37077,N_34813);
and U49457 (N_49457,N_35763,N_39104);
or U49458 (N_49458,N_31902,N_32419);
nor U49459 (N_49459,N_38595,N_37078);
nand U49460 (N_49460,N_35605,N_34089);
or U49461 (N_49461,N_31526,N_32953);
nand U49462 (N_49462,N_32426,N_35682);
xnor U49463 (N_49463,N_38464,N_39441);
nor U49464 (N_49464,N_31728,N_38587);
nor U49465 (N_49465,N_31435,N_37176);
nor U49466 (N_49466,N_31939,N_33965);
nor U49467 (N_49467,N_36224,N_33393);
nor U49468 (N_49468,N_31294,N_36985);
nor U49469 (N_49469,N_31561,N_35395);
nor U49470 (N_49470,N_32721,N_37824);
nor U49471 (N_49471,N_34428,N_38731);
nor U49472 (N_49472,N_39979,N_36319);
and U49473 (N_49473,N_34852,N_30995);
nor U49474 (N_49474,N_37714,N_34558);
nor U49475 (N_49475,N_39438,N_35096);
nor U49476 (N_49476,N_37664,N_32419);
or U49477 (N_49477,N_36048,N_38579);
nand U49478 (N_49478,N_37602,N_31469);
and U49479 (N_49479,N_37809,N_37937);
and U49480 (N_49480,N_34051,N_31425);
nand U49481 (N_49481,N_39221,N_38365);
nand U49482 (N_49482,N_38703,N_34882);
nor U49483 (N_49483,N_36704,N_36290);
or U49484 (N_49484,N_36234,N_38578);
or U49485 (N_49485,N_32931,N_37302);
or U49486 (N_49486,N_32461,N_36172);
or U49487 (N_49487,N_36725,N_35614);
xor U49488 (N_49488,N_39351,N_36796);
xnor U49489 (N_49489,N_37767,N_34487);
and U49490 (N_49490,N_33262,N_36066);
nand U49491 (N_49491,N_36329,N_34739);
nand U49492 (N_49492,N_38900,N_30914);
nor U49493 (N_49493,N_35606,N_36537);
or U49494 (N_49494,N_38196,N_35925);
xnor U49495 (N_49495,N_36581,N_30407);
nand U49496 (N_49496,N_31892,N_33360);
and U49497 (N_49497,N_37655,N_33440);
nor U49498 (N_49498,N_35343,N_31133);
xnor U49499 (N_49499,N_30716,N_39260);
nand U49500 (N_49500,N_32227,N_37364);
and U49501 (N_49501,N_33462,N_32019);
nand U49502 (N_49502,N_36008,N_32986);
nand U49503 (N_49503,N_30598,N_34564);
or U49504 (N_49504,N_35906,N_36173);
nand U49505 (N_49505,N_30127,N_38714);
nand U49506 (N_49506,N_38287,N_35187);
or U49507 (N_49507,N_35584,N_33142);
nor U49508 (N_49508,N_32166,N_32147);
and U49509 (N_49509,N_37910,N_36096);
nand U49510 (N_49510,N_32923,N_34221);
and U49511 (N_49511,N_39142,N_33878);
and U49512 (N_49512,N_30145,N_34043);
nor U49513 (N_49513,N_32180,N_31532);
nor U49514 (N_49514,N_31914,N_35830);
and U49515 (N_49515,N_33861,N_33070);
nor U49516 (N_49516,N_37885,N_36576);
or U49517 (N_49517,N_30750,N_38414);
or U49518 (N_49518,N_37802,N_37909);
xnor U49519 (N_49519,N_30743,N_36426);
xnor U49520 (N_49520,N_33618,N_35035);
and U49521 (N_49521,N_30516,N_33005);
and U49522 (N_49522,N_36289,N_35878);
nor U49523 (N_49523,N_37874,N_36366);
nor U49524 (N_49524,N_37811,N_38284);
nand U49525 (N_49525,N_38843,N_37410);
or U49526 (N_49526,N_39171,N_32307);
nor U49527 (N_49527,N_32444,N_37686);
or U49528 (N_49528,N_35927,N_30349);
nor U49529 (N_49529,N_31388,N_30591);
or U49530 (N_49530,N_32714,N_34102);
and U49531 (N_49531,N_37613,N_33473);
and U49532 (N_49532,N_30292,N_38148);
or U49533 (N_49533,N_31057,N_37478);
or U49534 (N_49534,N_32976,N_31055);
nand U49535 (N_49535,N_36845,N_39940);
or U49536 (N_49536,N_38458,N_34180);
nand U49537 (N_49537,N_32351,N_35298);
or U49538 (N_49538,N_36747,N_30489);
nor U49539 (N_49539,N_35219,N_35341);
or U49540 (N_49540,N_38180,N_35921);
and U49541 (N_49541,N_36018,N_31986);
nand U49542 (N_49542,N_30385,N_35752);
xor U49543 (N_49543,N_39883,N_33029);
or U49544 (N_49544,N_33690,N_37513);
or U49545 (N_49545,N_32542,N_37886);
nor U49546 (N_49546,N_38606,N_30786);
nand U49547 (N_49547,N_38407,N_32372);
nor U49548 (N_49548,N_39183,N_30451);
nor U49549 (N_49549,N_38571,N_34019);
or U49550 (N_49550,N_32570,N_39454);
and U49551 (N_49551,N_34721,N_35685);
nand U49552 (N_49552,N_33715,N_31553);
or U49553 (N_49553,N_32330,N_30061);
nor U49554 (N_49554,N_35510,N_30830);
and U49555 (N_49555,N_30215,N_31208);
and U49556 (N_49556,N_34921,N_37825);
or U49557 (N_49557,N_34555,N_35240);
nor U49558 (N_49558,N_35282,N_39297);
nand U49559 (N_49559,N_34051,N_30165);
nor U49560 (N_49560,N_31042,N_31192);
nand U49561 (N_49561,N_34412,N_36199);
nor U49562 (N_49562,N_37578,N_30174);
nor U49563 (N_49563,N_31694,N_32397);
nor U49564 (N_49564,N_38068,N_34772);
nand U49565 (N_49565,N_37591,N_36260);
nand U49566 (N_49566,N_38674,N_31125);
and U49567 (N_49567,N_33904,N_34070);
or U49568 (N_49568,N_35045,N_31017);
xnor U49569 (N_49569,N_33135,N_34742);
xnor U49570 (N_49570,N_37179,N_33927);
or U49571 (N_49571,N_37471,N_37709);
or U49572 (N_49572,N_30734,N_32401);
or U49573 (N_49573,N_36514,N_30822);
nand U49574 (N_49574,N_34810,N_36690);
nand U49575 (N_49575,N_36911,N_32680);
or U49576 (N_49576,N_39554,N_38354);
nand U49577 (N_49577,N_31493,N_37933);
and U49578 (N_49578,N_35985,N_32804);
nand U49579 (N_49579,N_34816,N_35275);
xor U49580 (N_49580,N_37792,N_30440);
xor U49581 (N_49581,N_30930,N_32617);
nand U49582 (N_49582,N_35708,N_30457);
xnor U49583 (N_49583,N_39622,N_39150);
and U49584 (N_49584,N_31758,N_35539);
and U49585 (N_49585,N_36804,N_31180);
xor U49586 (N_49586,N_33670,N_33653);
or U49587 (N_49587,N_36960,N_31329);
nand U49588 (N_49588,N_34187,N_31129);
nand U49589 (N_49589,N_39851,N_33161);
and U49590 (N_49590,N_38344,N_35238);
xor U49591 (N_49591,N_34555,N_34256);
or U49592 (N_49592,N_39938,N_37216);
nor U49593 (N_49593,N_30544,N_30512);
or U49594 (N_49594,N_32454,N_31360);
and U49595 (N_49595,N_31062,N_32572);
or U49596 (N_49596,N_38431,N_36389);
nor U49597 (N_49597,N_30525,N_36029);
nand U49598 (N_49598,N_31535,N_36107);
nor U49599 (N_49599,N_34198,N_33581);
and U49600 (N_49600,N_35497,N_37646);
and U49601 (N_49601,N_35074,N_37019);
xor U49602 (N_49602,N_30148,N_35000);
xor U49603 (N_49603,N_33772,N_39841);
or U49604 (N_49604,N_39737,N_34210);
nor U49605 (N_49605,N_30975,N_31929);
nor U49606 (N_49606,N_33692,N_39258);
nor U49607 (N_49607,N_39237,N_33174);
or U49608 (N_49608,N_34286,N_35250);
and U49609 (N_49609,N_30307,N_39161);
xor U49610 (N_49610,N_35601,N_34905);
nand U49611 (N_49611,N_30236,N_34535);
and U49612 (N_49612,N_34008,N_33036);
nor U49613 (N_49613,N_34184,N_30747);
nand U49614 (N_49614,N_35657,N_31651);
nor U49615 (N_49615,N_34808,N_33861);
or U49616 (N_49616,N_35542,N_32872);
nor U49617 (N_49617,N_33666,N_33785);
or U49618 (N_49618,N_33182,N_30729);
nor U49619 (N_49619,N_33815,N_30769);
nand U49620 (N_49620,N_37056,N_35838);
nor U49621 (N_49621,N_35594,N_31561);
nor U49622 (N_49622,N_31429,N_30095);
and U49623 (N_49623,N_38426,N_38245);
nand U49624 (N_49624,N_37427,N_31823);
and U49625 (N_49625,N_37484,N_31447);
nor U49626 (N_49626,N_37269,N_37760);
and U49627 (N_49627,N_37360,N_38848);
nand U49628 (N_49628,N_33721,N_34912);
nor U49629 (N_49629,N_39315,N_36488);
or U49630 (N_49630,N_39719,N_32111);
nor U49631 (N_49631,N_32146,N_36612);
or U49632 (N_49632,N_32982,N_34653);
or U49633 (N_49633,N_33862,N_30188);
or U49634 (N_49634,N_35187,N_38439);
or U49635 (N_49635,N_33092,N_35764);
nor U49636 (N_49636,N_38277,N_37542);
nor U49637 (N_49637,N_39833,N_31870);
nor U49638 (N_49638,N_34151,N_34382);
or U49639 (N_49639,N_35792,N_32659);
nand U49640 (N_49640,N_30504,N_32312);
or U49641 (N_49641,N_30370,N_39573);
nor U49642 (N_49642,N_33150,N_32969);
nor U49643 (N_49643,N_32864,N_31514);
and U49644 (N_49644,N_34912,N_32811);
xor U49645 (N_49645,N_35111,N_38399);
nor U49646 (N_49646,N_36500,N_34419);
and U49647 (N_49647,N_38089,N_30905);
nand U49648 (N_49648,N_33355,N_32621);
or U49649 (N_49649,N_35282,N_31295);
and U49650 (N_49650,N_39977,N_35333);
or U49651 (N_49651,N_31657,N_37513);
or U49652 (N_49652,N_32549,N_34069);
nor U49653 (N_49653,N_38372,N_32056);
nor U49654 (N_49654,N_32730,N_32421);
xor U49655 (N_49655,N_33435,N_36678);
or U49656 (N_49656,N_38082,N_34076);
nor U49657 (N_49657,N_36477,N_32943);
nor U49658 (N_49658,N_35668,N_34763);
and U49659 (N_49659,N_38698,N_39935);
nor U49660 (N_49660,N_36684,N_37218);
nor U49661 (N_49661,N_31621,N_32458);
or U49662 (N_49662,N_32531,N_30261);
or U49663 (N_49663,N_30050,N_33909);
nor U49664 (N_49664,N_36551,N_38034);
or U49665 (N_49665,N_36886,N_36059);
xnor U49666 (N_49666,N_36798,N_39422);
xor U49667 (N_49667,N_31365,N_32175);
nor U49668 (N_49668,N_37266,N_37493);
or U49669 (N_49669,N_36497,N_33986);
or U49670 (N_49670,N_35494,N_31136);
nor U49671 (N_49671,N_39709,N_38543);
nand U49672 (N_49672,N_31463,N_31439);
or U49673 (N_49673,N_32472,N_37195);
xnor U49674 (N_49674,N_37643,N_32497);
and U49675 (N_49675,N_36264,N_39759);
or U49676 (N_49676,N_30604,N_38787);
nand U49677 (N_49677,N_36387,N_34905);
or U49678 (N_49678,N_38473,N_34006);
and U49679 (N_49679,N_34811,N_30811);
nand U49680 (N_49680,N_38460,N_34627);
xnor U49681 (N_49681,N_36081,N_37049);
nor U49682 (N_49682,N_36567,N_32184);
or U49683 (N_49683,N_33710,N_32966);
nor U49684 (N_49684,N_38401,N_32234);
nand U49685 (N_49685,N_34100,N_34308);
xor U49686 (N_49686,N_32846,N_33642);
or U49687 (N_49687,N_36278,N_39479);
or U49688 (N_49688,N_35739,N_35933);
and U49689 (N_49689,N_32923,N_36146);
nor U49690 (N_49690,N_32592,N_36563);
and U49691 (N_49691,N_39108,N_33126);
nand U49692 (N_49692,N_32017,N_33797);
and U49693 (N_49693,N_34617,N_33134);
or U49694 (N_49694,N_37052,N_31082);
or U49695 (N_49695,N_33877,N_33123);
or U49696 (N_49696,N_32114,N_31411);
nand U49697 (N_49697,N_35055,N_37458);
nor U49698 (N_49698,N_39562,N_39097);
xor U49699 (N_49699,N_35275,N_38420);
nand U49700 (N_49700,N_32612,N_32379);
xor U49701 (N_49701,N_33054,N_35292);
nor U49702 (N_49702,N_36722,N_34375);
and U49703 (N_49703,N_32921,N_33230);
nor U49704 (N_49704,N_38345,N_38754);
nand U49705 (N_49705,N_34051,N_37207);
and U49706 (N_49706,N_37856,N_33194);
and U49707 (N_49707,N_32621,N_35785);
nand U49708 (N_49708,N_39692,N_39651);
and U49709 (N_49709,N_34118,N_35334);
nand U49710 (N_49710,N_34605,N_38692);
or U49711 (N_49711,N_36260,N_38053);
or U49712 (N_49712,N_31711,N_30158);
and U49713 (N_49713,N_37799,N_31379);
nand U49714 (N_49714,N_31153,N_39624);
and U49715 (N_49715,N_33987,N_35710);
and U49716 (N_49716,N_33508,N_36210);
xnor U49717 (N_49717,N_38610,N_38637);
and U49718 (N_49718,N_36607,N_37597);
nand U49719 (N_49719,N_34639,N_38877);
nand U49720 (N_49720,N_35854,N_38035);
or U49721 (N_49721,N_30261,N_35931);
nand U49722 (N_49722,N_39692,N_33611);
nor U49723 (N_49723,N_33840,N_36853);
nand U49724 (N_49724,N_35387,N_31412);
nor U49725 (N_49725,N_37822,N_31651);
nor U49726 (N_49726,N_35618,N_32741);
or U49727 (N_49727,N_32194,N_36881);
and U49728 (N_49728,N_35637,N_37213);
and U49729 (N_49729,N_32774,N_38659);
or U49730 (N_49730,N_37046,N_38660);
nor U49731 (N_49731,N_39597,N_35880);
nor U49732 (N_49732,N_38168,N_31941);
xor U49733 (N_49733,N_39168,N_37172);
or U49734 (N_49734,N_35066,N_30438);
or U49735 (N_49735,N_31937,N_39113);
nor U49736 (N_49736,N_34439,N_38898);
or U49737 (N_49737,N_30825,N_35215);
and U49738 (N_49738,N_35567,N_39890);
nand U49739 (N_49739,N_31492,N_33989);
nand U49740 (N_49740,N_37199,N_34815);
nand U49741 (N_49741,N_39586,N_34973);
or U49742 (N_49742,N_35266,N_38563);
nor U49743 (N_49743,N_33079,N_36675);
nor U49744 (N_49744,N_34282,N_33648);
xnor U49745 (N_49745,N_30918,N_39055);
xor U49746 (N_49746,N_30643,N_39486);
xor U49747 (N_49747,N_35137,N_31125);
or U49748 (N_49748,N_35540,N_31104);
and U49749 (N_49749,N_33132,N_36008);
and U49750 (N_49750,N_38523,N_33433);
nand U49751 (N_49751,N_38395,N_35732);
and U49752 (N_49752,N_31885,N_34548);
and U49753 (N_49753,N_35051,N_30315);
xnor U49754 (N_49754,N_31867,N_38172);
and U49755 (N_49755,N_38475,N_36127);
or U49756 (N_49756,N_30370,N_31535);
nand U49757 (N_49757,N_37385,N_36732);
nand U49758 (N_49758,N_32854,N_35503);
nand U49759 (N_49759,N_33383,N_37228);
or U49760 (N_49760,N_34906,N_32124);
xor U49761 (N_49761,N_32601,N_36859);
nor U49762 (N_49762,N_34850,N_38264);
nand U49763 (N_49763,N_36769,N_35780);
and U49764 (N_49764,N_38362,N_34283);
and U49765 (N_49765,N_37814,N_32669);
and U49766 (N_49766,N_39329,N_30681);
nor U49767 (N_49767,N_34904,N_36593);
nand U49768 (N_49768,N_30046,N_35479);
and U49769 (N_49769,N_35932,N_35254);
and U49770 (N_49770,N_35498,N_38797);
nor U49771 (N_49771,N_33343,N_30662);
nor U49772 (N_49772,N_33520,N_37110);
or U49773 (N_49773,N_32686,N_31034);
and U49774 (N_49774,N_30483,N_35361);
and U49775 (N_49775,N_31753,N_35214);
nand U49776 (N_49776,N_30628,N_39061);
and U49777 (N_49777,N_32798,N_35899);
nor U49778 (N_49778,N_39764,N_35026);
and U49779 (N_49779,N_39418,N_33775);
nor U49780 (N_49780,N_36500,N_37826);
nand U49781 (N_49781,N_36725,N_39176);
and U49782 (N_49782,N_32647,N_34590);
nand U49783 (N_49783,N_39144,N_34939);
xor U49784 (N_49784,N_30082,N_37815);
nand U49785 (N_49785,N_35016,N_31459);
nand U49786 (N_49786,N_31334,N_37120);
nor U49787 (N_49787,N_39653,N_36648);
nor U49788 (N_49788,N_37430,N_38875);
nor U49789 (N_49789,N_34368,N_35995);
nor U49790 (N_49790,N_31703,N_39168);
and U49791 (N_49791,N_35349,N_37043);
and U49792 (N_49792,N_39493,N_32145);
or U49793 (N_49793,N_34909,N_30671);
nor U49794 (N_49794,N_34411,N_36356);
nor U49795 (N_49795,N_37730,N_33816);
and U49796 (N_49796,N_34167,N_31485);
and U49797 (N_49797,N_39565,N_33757);
nor U49798 (N_49798,N_30497,N_38501);
nand U49799 (N_49799,N_39486,N_34196);
or U49800 (N_49800,N_35533,N_33333);
xor U49801 (N_49801,N_33392,N_32110);
nor U49802 (N_49802,N_35298,N_31361);
and U49803 (N_49803,N_36367,N_30718);
nand U49804 (N_49804,N_33683,N_31535);
and U49805 (N_49805,N_34563,N_34335);
or U49806 (N_49806,N_37693,N_35540);
and U49807 (N_49807,N_31158,N_34244);
nor U49808 (N_49808,N_30048,N_35971);
xnor U49809 (N_49809,N_34512,N_34863);
nor U49810 (N_49810,N_36166,N_37603);
nand U49811 (N_49811,N_30411,N_34898);
or U49812 (N_49812,N_39329,N_33489);
and U49813 (N_49813,N_38102,N_38892);
nor U49814 (N_49814,N_38083,N_39966);
xor U49815 (N_49815,N_39626,N_37808);
or U49816 (N_49816,N_31840,N_34032);
xor U49817 (N_49817,N_35063,N_34576);
xnor U49818 (N_49818,N_31197,N_39174);
and U49819 (N_49819,N_35883,N_38577);
nor U49820 (N_49820,N_30883,N_32451);
or U49821 (N_49821,N_34331,N_30408);
nand U49822 (N_49822,N_37889,N_33182);
and U49823 (N_49823,N_37817,N_38229);
xor U49824 (N_49824,N_32751,N_32495);
nand U49825 (N_49825,N_31175,N_35025);
and U49826 (N_49826,N_37793,N_32024);
and U49827 (N_49827,N_32146,N_30041);
xnor U49828 (N_49828,N_36546,N_39692);
nor U49829 (N_49829,N_30257,N_32191);
nand U49830 (N_49830,N_38859,N_34475);
nand U49831 (N_49831,N_38875,N_30593);
and U49832 (N_49832,N_35237,N_37563);
nor U49833 (N_49833,N_33733,N_31683);
nor U49834 (N_49834,N_34459,N_31902);
xor U49835 (N_49835,N_35540,N_34598);
nor U49836 (N_49836,N_38596,N_31776);
or U49837 (N_49837,N_34574,N_34109);
and U49838 (N_49838,N_36951,N_36649);
and U49839 (N_49839,N_39985,N_33059);
nand U49840 (N_49840,N_30345,N_32825);
or U49841 (N_49841,N_33070,N_34733);
nor U49842 (N_49842,N_36106,N_34655);
and U49843 (N_49843,N_36464,N_35786);
or U49844 (N_49844,N_32825,N_37674);
and U49845 (N_49845,N_36607,N_31666);
nand U49846 (N_49846,N_39898,N_37388);
or U49847 (N_49847,N_37954,N_39098);
or U49848 (N_49848,N_37291,N_35264);
or U49849 (N_49849,N_34342,N_38468);
xor U49850 (N_49850,N_34745,N_37393);
and U49851 (N_49851,N_31383,N_34083);
nand U49852 (N_49852,N_39846,N_36622);
or U49853 (N_49853,N_34558,N_36405);
xor U49854 (N_49854,N_32753,N_35091);
xnor U49855 (N_49855,N_38256,N_38039);
xor U49856 (N_49856,N_35340,N_33351);
and U49857 (N_49857,N_35824,N_33959);
nor U49858 (N_49858,N_39032,N_37753);
and U49859 (N_49859,N_30887,N_35603);
and U49860 (N_49860,N_39233,N_31242);
and U49861 (N_49861,N_30493,N_33266);
xor U49862 (N_49862,N_36116,N_35102);
nor U49863 (N_49863,N_39458,N_39188);
and U49864 (N_49864,N_34702,N_35460);
nand U49865 (N_49865,N_30646,N_33632);
nand U49866 (N_49866,N_32573,N_35115);
xor U49867 (N_49867,N_36977,N_32734);
nand U49868 (N_49868,N_38807,N_39393);
nand U49869 (N_49869,N_37012,N_33281);
or U49870 (N_49870,N_33110,N_32871);
or U49871 (N_49871,N_36777,N_36121);
or U49872 (N_49872,N_31198,N_34877);
nor U49873 (N_49873,N_37858,N_38626);
nor U49874 (N_49874,N_32705,N_37144);
or U49875 (N_49875,N_35681,N_35100);
nor U49876 (N_49876,N_33108,N_34863);
or U49877 (N_49877,N_37662,N_35037);
or U49878 (N_49878,N_33173,N_30389);
and U49879 (N_49879,N_32944,N_38050);
nor U49880 (N_49880,N_32089,N_39463);
xnor U49881 (N_49881,N_39216,N_33748);
and U49882 (N_49882,N_33569,N_33428);
nand U49883 (N_49883,N_38854,N_36852);
nand U49884 (N_49884,N_32163,N_31416);
and U49885 (N_49885,N_35832,N_36839);
nor U49886 (N_49886,N_33721,N_34515);
and U49887 (N_49887,N_36015,N_34085);
nor U49888 (N_49888,N_32533,N_39285);
or U49889 (N_49889,N_35008,N_35543);
nand U49890 (N_49890,N_34432,N_37871);
or U49891 (N_49891,N_30133,N_34724);
and U49892 (N_49892,N_33369,N_35698);
or U49893 (N_49893,N_30890,N_30719);
and U49894 (N_49894,N_32799,N_33730);
nand U49895 (N_49895,N_32850,N_34277);
nor U49896 (N_49896,N_36911,N_33610);
or U49897 (N_49897,N_37778,N_31138);
nor U49898 (N_49898,N_30599,N_33447);
nand U49899 (N_49899,N_37363,N_38673);
and U49900 (N_49900,N_30807,N_31401);
or U49901 (N_49901,N_38296,N_36580);
and U49902 (N_49902,N_33072,N_39025);
nor U49903 (N_49903,N_30776,N_34918);
nor U49904 (N_49904,N_36245,N_35940);
or U49905 (N_49905,N_30197,N_38540);
nor U49906 (N_49906,N_36187,N_37878);
xor U49907 (N_49907,N_34701,N_31795);
or U49908 (N_49908,N_37878,N_30001);
or U49909 (N_49909,N_30314,N_36938);
and U49910 (N_49910,N_33679,N_31993);
nor U49911 (N_49911,N_30501,N_34660);
nor U49912 (N_49912,N_31547,N_39966);
nor U49913 (N_49913,N_30605,N_31186);
xor U49914 (N_49914,N_32212,N_37982);
nand U49915 (N_49915,N_33052,N_35978);
or U49916 (N_49916,N_36034,N_39225);
or U49917 (N_49917,N_30927,N_36622);
nand U49918 (N_49918,N_36446,N_39817);
and U49919 (N_49919,N_31619,N_38069);
and U49920 (N_49920,N_34876,N_34379);
and U49921 (N_49921,N_34735,N_32809);
xor U49922 (N_49922,N_35057,N_31855);
or U49923 (N_49923,N_30359,N_31060);
nand U49924 (N_49924,N_39890,N_30516);
or U49925 (N_49925,N_30213,N_39645);
or U49926 (N_49926,N_37572,N_38490);
xnor U49927 (N_49927,N_32208,N_35832);
and U49928 (N_49928,N_33047,N_31528);
nor U49929 (N_49929,N_36893,N_32219);
or U49930 (N_49930,N_30141,N_37105);
nor U49931 (N_49931,N_36471,N_39734);
nor U49932 (N_49932,N_39284,N_39272);
nand U49933 (N_49933,N_36986,N_34965);
nor U49934 (N_49934,N_34526,N_35371);
and U49935 (N_49935,N_38278,N_30942);
and U49936 (N_49936,N_34309,N_36266);
and U49937 (N_49937,N_31414,N_37807);
and U49938 (N_49938,N_32346,N_33973);
xor U49939 (N_49939,N_38915,N_37997);
nand U49940 (N_49940,N_38485,N_37545);
nor U49941 (N_49941,N_31373,N_34106);
xnor U49942 (N_49942,N_36281,N_33232);
nor U49943 (N_49943,N_34093,N_36925);
and U49944 (N_49944,N_39276,N_33999);
xor U49945 (N_49945,N_36282,N_36346);
nand U49946 (N_49946,N_34719,N_38123);
xnor U49947 (N_49947,N_33543,N_39507);
xnor U49948 (N_49948,N_35258,N_36454);
xor U49949 (N_49949,N_35685,N_30508);
or U49950 (N_49950,N_31922,N_36758);
and U49951 (N_49951,N_35763,N_39407);
or U49952 (N_49952,N_36415,N_33230);
nand U49953 (N_49953,N_39967,N_38578);
and U49954 (N_49954,N_34014,N_30339);
and U49955 (N_49955,N_38549,N_38476);
and U49956 (N_49956,N_38253,N_34775);
nand U49957 (N_49957,N_39745,N_38032);
and U49958 (N_49958,N_38088,N_38207);
nor U49959 (N_49959,N_33506,N_39128);
and U49960 (N_49960,N_33153,N_38220);
nor U49961 (N_49961,N_38854,N_33301);
or U49962 (N_49962,N_35791,N_31275);
and U49963 (N_49963,N_34579,N_35551);
and U49964 (N_49964,N_30796,N_35084);
and U49965 (N_49965,N_35383,N_38478);
and U49966 (N_49966,N_32820,N_34229);
nor U49967 (N_49967,N_31859,N_32243);
and U49968 (N_49968,N_37692,N_31075);
nor U49969 (N_49969,N_37934,N_36204);
and U49970 (N_49970,N_39687,N_36278);
or U49971 (N_49971,N_32391,N_36840);
nand U49972 (N_49972,N_33220,N_31485);
or U49973 (N_49973,N_33732,N_31812);
or U49974 (N_49974,N_38771,N_30711);
and U49975 (N_49975,N_35517,N_38072);
or U49976 (N_49976,N_38799,N_30747);
and U49977 (N_49977,N_32770,N_39606);
or U49978 (N_49978,N_32220,N_39294);
nand U49979 (N_49979,N_34525,N_36298);
or U49980 (N_49980,N_33125,N_30720);
nand U49981 (N_49981,N_38352,N_32014);
and U49982 (N_49982,N_35925,N_39992);
nor U49983 (N_49983,N_37337,N_35489);
xnor U49984 (N_49984,N_32274,N_32476);
xnor U49985 (N_49985,N_34534,N_38172);
and U49986 (N_49986,N_35197,N_32540);
nor U49987 (N_49987,N_39621,N_37225);
or U49988 (N_49988,N_39594,N_31078);
and U49989 (N_49989,N_34988,N_39335);
or U49990 (N_49990,N_32798,N_30485);
nand U49991 (N_49991,N_31749,N_37108);
nand U49992 (N_49992,N_37901,N_39015);
and U49993 (N_49993,N_38387,N_36999);
xor U49994 (N_49994,N_30111,N_38936);
xnor U49995 (N_49995,N_35934,N_31999);
and U49996 (N_49996,N_39707,N_31681);
or U49997 (N_49997,N_39523,N_32824);
and U49998 (N_49998,N_32361,N_33320);
nand U49999 (N_49999,N_33603,N_39225);
and UO_0 (O_0,N_42696,N_42664);
nand UO_1 (O_1,N_48589,N_49741);
xor UO_2 (O_2,N_45480,N_41688);
or UO_3 (O_3,N_40989,N_47510);
nor UO_4 (O_4,N_43771,N_45621);
or UO_5 (O_5,N_44887,N_43032);
and UO_6 (O_6,N_49114,N_44431);
or UO_7 (O_7,N_47908,N_41483);
or UO_8 (O_8,N_41351,N_41172);
nor UO_9 (O_9,N_45036,N_47631);
and UO_10 (O_10,N_49762,N_49421);
nand UO_11 (O_11,N_43426,N_41042);
and UO_12 (O_12,N_46556,N_40771);
or UO_13 (O_13,N_45128,N_43370);
nor UO_14 (O_14,N_42119,N_47824);
or UO_15 (O_15,N_42151,N_43683);
nand UO_16 (O_16,N_44151,N_47242);
and UO_17 (O_17,N_40744,N_41786);
and UO_18 (O_18,N_40904,N_43815);
or UO_19 (O_19,N_43203,N_45364);
and UO_20 (O_20,N_42300,N_45537);
nand UO_21 (O_21,N_46446,N_46583);
or UO_22 (O_22,N_48414,N_42335);
xor UO_23 (O_23,N_41685,N_46823);
or UO_24 (O_24,N_42910,N_48082);
and UO_25 (O_25,N_45176,N_43424);
nand UO_26 (O_26,N_43462,N_40219);
nor UO_27 (O_27,N_46425,N_46919);
nor UO_28 (O_28,N_49335,N_43357);
nor UO_29 (O_29,N_40275,N_41503);
nand UO_30 (O_30,N_47929,N_46064);
nor UO_31 (O_31,N_46688,N_45986);
nor UO_32 (O_32,N_40630,N_45589);
and UO_33 (O_33,N_49424,N_46994);
nand UO_34 (O_34,N_41652,N_42692);
xnor UO_35 (O_35,N_49394,N_49919);
nor UO_36 (O_36,N_41429,N_49026);
and UO_37 (O_37,N_43379,N_42852);
nor UO_38 (O_38,N_43856,N_43708);
or UO_39 (O_39,N_43481,N_45242);
xnor UO_40 (O_40,N_43187,N_43245);
nand UO_41 (O_41,N_45733,N_46992);
and UO_42 (O_42,N_45546,N_43513);
or UO_43 (O_43,N_43799,N_47200);
nor UO_44 (O_44,N_46609,N_48013);
and UO_45 (O_45,N_47494,N_48982);
or UO_46 (O_46,N_46793,N_46828);
nor UO_47 (O_47,N_41080,N_44763);
and UO_48 (O_48,N_47093,N_42257);
or UO_49 (O_49,N_46124,N_42178);
or UO_50 (O_50,N_44133,N_45812);
or UO_51 (O_51,N_42958,N_48996);
or UO_52 (O_52,N_45517,N_48363);
xor UO_53 (O_53,N_48678,N_45063);
and UO_54 (O_54,N_40268,N_43041);
and UO_55 (O_55,N_41173,N_45641);
nand UO_56 (O_56,N_47312,N_43564);
or UO_57 (O_57,N_42713,N_45634);
or UO_58 (O_58,N_42954,N_43959);
and UO_59 (O_59,N_46502,N_47323);
nand UO_60 (O_60,N_49453,N_43729);
nand UO_61 (O_61,N_41621,N_44807);
xor UO_62 (O_62,N_43570,N_48057);
nand UO_63 (O_63,N_46822,N_42641);
xnor UO_64 (O_64,N_41096,N_45366);
xnor UO_65 (O_65,N_45246,N_40036);
nand UO_66 (O_66,N_42551,N_49481);
and UO_67 (O_67,N_43456,N_42019);
nand UO_68 (O_68,N_42404,N_47559);
and UO_69 (O_69,N_47883,N_48604);
and UO_70 (O_70,N_43810,N_46861);
xor UO_71 (O_71,N_41408,N_45963);
and UO_72 (O_72,N_40843,N_43943);
and UO_73 (O_73,N_48388,N_40419);
nor UO_74 (O_74,N_44155,N_48289);
nand UO_75 (O_75,N_43969,N_45191);
nand UO_76 (O_76,N_45208,N_41713);
and UO_77 (O_77,N_44302,N_49122);
or UO_78 (O_78,N_47153,N_41884);
and UO_79 (O_79,N_48266,N_45576);
xnor UO_80 (O_80,N_43169,N_43993);
xor UO_81 (O_81,N_41896,N_49707);
nand UO_82 (O_82,N_45972,N_44741);
and UO_83 (O_83,N_44262,N_47893);
or UO_84 (O_84,N_40503,N_40525);
nand UO_85 (O_85,N_41935,N_45585);
and UO_86 (O_86,N_42920,N_44776);
nor UO_87 (O_87,N_42053,N_46803);
nand UO_88 (O_88,N_40171,N_47493);
or UO_89 (O_89,N_48440,N_40163);
nor UO_90 (O_90,N_47944,N_40612);
nand UO_91 (O_91,N_41211,N_45170);
or UO_92 (O_92,N_40686,N_43742);
nor UO_93 (O_93,N_46755,N_49474);
or UO_94 (O_94,N_42307,N_46888);
nor UO_95 (O_95,N_47948,N_41524);
or UO_96 (O_96,N_41677,N_43700);
or UO_97 (O_97,N_48207,N_40211);
nor UO_98 (O_98,N_40511,N_49177);
and UO_99 (O_99,N_46060,N_43093);
or UO_100 (O_100,N_46790,N_48722);
and UO_101 (O_101,N_44386,N_45133);
nand UO_102 (O_102,N_41229,N_49570);
or UO_103 (O_103,N_46869,N_45074);
nand UO_104 (O_104,N_45401,N_40308);
and UO_105 (O_105,N_44743,N_49382);
nand UO_106 (O_106,N_43420,N_44245);
nand UO_107 (O_107,N_40790,N_40181);
nor UO_108 (O_108,N_43869,N_44137);
and UO_109 (O_109,N_45427,N_42767);
and UO_110 (O_110,N_45215,N_43410);
xor UO_111 (O_111,N_42754,N_42979);
nor UO_112 (O_112,N_44110,N_49594);
and UO_113 (O_113,N_47939,N_46907);
xor UO_114 (O_114,N_41395,N_42511);
nand UO_115 (O_115,N_43928,N_43224);
and UO_116 (O_116,N_43642,N_44844);
nand UO_117 (O_117,N_40690,N_44559);
nor UO_118 (O_118,N_40773,N_44703);
nor UO_119 (O_119,N_49609,N_41320);
nor UO_120 (O_120,N_47937,N_43659);
or UO_121 (O_121,N_43834,N_44552);
nand UO_122 (O_122,N_49371,N_43673);
nor UO_123 (O_123,N_42984,N_45791);
and UO_124 (O_124,N_48368,N_40089);
nand UO_125 (O_125,N_48071,N_49281);
or UO_126 (O_126,N_43950,N_42678);
or UO_127 (O_127,N_48592,N_46340);
nor UO_128 (O_128,N_48839,N_48342);
nand UO_129 (O_129,N_46927,N_46883);
nor UO_130 (O_130,N_42850,N_45345);
nor UO_131 (O_131,N_44358,N_46945);
nand UO_132 (O_132,N_43393,N_44173);
nand UO_133 (O_133,N_45387,N_41510);
or UO_134 (O_134,N_46240,N_40902);
xor UO_135 (O_135,N_46905,N_42513);
or UO_136 (O_136,N_48404,N_41291);
nor UO_137 (O_137,N_46619,N_43303);
or UO_138 (O_138,N_48499,N_47408);
nand UO_139 (O_139,N_44746,N_47066);
nand UO_140 (O_140,N_40215,N_42201);
and UO_141 (O_141,N_40860,N_45057);
and UO_142 (O_142,N_43244,N_47571);
and UO_143 (O_143,N_48016,N_41855);
or UO_144 (O_144,N_43806,N_40868);
and UO_145 (O_145,N_47081,N_42423);
and UO_146 (O_146,N_41934,N_46133);
or UO_147 (O_147,N_42563,N_42647);
nand UO_148 (O_148,N_49681,N_48731);
nor UO_149 (O_149,N_49030,N_45195);
or UO_150 (O_150,N_43355,N_40376);
or UO_151 (O_151,N_41137,N_48462);
nand UO_152 (O_152,N_44616,N_49184);
nand UO_153 (O_153,N_41060,N_40195);
and UO_154 (O_154,N_47725,N_42565);
and UO_155 (O_155,N_43568,N_47434);
nor UO_156 (O_156,N_45219,N_45165);
nand UO_157 (O_157,N_42816,N_47722);
nand UO_158 (O_158,N_42415,N_41146);
or UO_159 (O_159,N_46379,N_45013);
xnor UO_160 (O_160,N_49361,N_48554);
and UO_161 (O_161,N_48895,N_49337);
nor UO_162 (O_162,N_47421,N_45188);
or UO_163 (O_163,N_45040,N_42576);
and UO_164 (O_164,N_42614,N_44018);
or UO_165 (O_165,N_43575,N_46887);
nor UO_166 (O_166,N_47507,N_48714);
or UO_167 (O_167,N_45107,N_48339);
xor UO_168 (O_168,N_43211,N_46552);
nand UO_169 (O_169,N_43276,N_41602);
nor UO_170 (O_170,N_47912,N_48491);
nand UO_171 (O_171,N_46788,N_43933);
nor UO_172 (O_172,N_46511,N_46929);
and UO_173 (O_173,N_46058,N_41201);
nand UO_174 (O_174,N_43754,N_44352);
or UO_175 (O_175,N_41259,N_47680);
nor UO_176 (O_176,N_41402,N_41116);
and UO_177 (O_177,N_46461,N_44187);
xor UO_178 (O_178,N_40292,N_47634);
nor UO_179 (O_179,N_49610,N_43764);
nand UO_180 (O_180,N_41389,N_49555);
nor UO_181 (O_181,N_45676,N_41922);
and UO_182 (O_182,N_41352,N_49370);
or UO_183 (O_183,N_42126,N_49931);
or UO_184 (O_184,N_47989,N_43098);
or UO_185 (O_185,N_43396,N_42129);
nor UO_186 (O_186,N_42539,N_47451);
nor UO_187 (O_187,N_42328,N_49841);
nor UO_188 (O_188,N_42853,N_49706);
nand UO_189 (O_189,N_40415,N_47640);
nand UO_190 (O_190,N_45530,N_45079);
or UO_191 (O_191,N_48978,N_43318);
or UO_192 (O_192,N_43202,N_49790);
xor UO_193 (O_193,N_45931,N_49347);
or UO_194 (O_194,N_40269,N_46951);
xnor UO_195 (O_195,N_48838,N_44577);
or UO_196 (O_196,N_41633,N_48919);
nand UO_197 (O_197,N_49280,N_47616);
nor UO_198 (O_198,N_46965,N_40019);
nand UO_199 (O_199,N_47519,N_49265);
and UO_200 (O_200,N_41777,N_47746);
nor UO_201 (O_201,N_40286,N_43835);
nand UO_202 (O_202,N_44486,N_46308);
nor UO_203 (O_203,N_44476,N_49772);
and UO_204 (O_204,N_43209,N_49994);
and UO_205 (O_205,N_44996,N_49461);
or UO_206 (O_206,N_49220,N_43688);
and UO_207 (O_207,N_42690,N_47349);
nor UO_208 (O_208,N_47768,N_41244);
and UO_209 (O_209,N_47872,N_41655);
xor UO_210 (O_210,N_42054,N_47765);
and UO_211 (O_211,N_47992,N_48928);
nor UO_212 (O_212,N_42488,N_45131);
nor UO_213 (O_213,N_44667,N_46862);
and UO_214 (O_214,N_40578,N_49082);
nor UO_215 (O_215,N_44898,N_42985);
nand UO_216 (O_216,N_42961,N_48235);
xnor UO_217 (O_217,N_43766,N_48726);
nand UO_218 (O_218,N_49812,N_44414);
nor UO_219 (O_219,N_44533,N_45702);
xor UO_220 (O_220,N_44069,N_46632);
and UO_221 (O_221,N_45948,N_46193);
nand UO_222 (O_222,N_46186,N_42859);
xnor UO_223 (O_223,N_45588,N_46660);
or UO_224 (O_224,N_41029,N_45636);
or UO_225 (O_225,N_47363,N_47582);
nand UO_226 (O_226,N_49605,N_43183);
and UO_227 (O_227,N_44906,N_45056);
nand UO_228 (O_228,N_47648,N_47804);
and UO_229 (O_229,N_41459,N_44409);
or UO_230 (O_230,N_49884,N_47467);
nand UO_231 (O_231,N_40177,N_43509);
nand UO_232 (O_232,N_43632,N_48497);
or UO_233 (O_233,N_41221,N_40194);
and UO_234 (O_234,N_49846,N_42062);
and UO_235 (O_235,N_41810,N_40403);
and UO_236 (O_236,N_49304,N_44064);
and UO_237 (O_237,N_48723,N_42096);
nand UO_238 (O_238,N_45988,N_47412);
nand UO_239 (O_239,N_41959,N_42680);
and UO_240 (O_240,N_48992,N_44450);
xor UO_241 (O_241,N_48463,N_42067);
nand UO_242 (O_242,N_47838,N_44960);
nor UO_243 (O_243,N_49447,N_45201);
and UO_244 (O_244,N_49124,N_44466);
and UO_245 (O_245,N_43618,N_44865);
nand UO_246 (O_246,N_47596,N_47877);
nor UO_247 (O_247,N_41644,N_40465);
xnor UO_248 (O_248,N_47202,N_40558);
or UO_249 (O_249,N_43987,N_46387);
and UO_250 (O_250,N_42135,N_44167);
nand UO_251 (O_251,N_45760,N_48543);
or UO_252 (O_252,N_41719,N_46617);
nand UO_253 (O_253,N_40009,N_47377);
or UO_254 (O_254,N_44516,N_43066);
xor UO_255 (O_255,N_42015,N_45510);
or UO_256 (O_256,N_49500,N_40916);
xor UO_257 (O_257,N_46260,N_40872);
nor UO_258 (O_258,N_40619,N_49291);
and UO_259 (O_259,N_47713,N_40967);
nor UO_260 (O_260,N_40853,N_45374);
and UO_261 (O_261,N_45727,N_43499);
nor UO_262 (O_262,N_48576,N_45493);
xor UO_263 (O_263,N_44881,N_42124);
xor UO_264 (O_264,N_46066,N_49312);
nand UO_265 (O_265,N_45077,N_40021);
and UO_266 (O_266,N_47546,N_43177);
nand UO_267 (O_267,N_48479,N_48527);
or UO_268 (O_268,N_40646,N_47524);
xor UO_269 (O_269,N_42219,N_48674);
nor UO_270 (O_270,N_43983,N_44598);
nand UO_271 (O_271,N_49121,N_44231);
or UO_272 (O_272,N_41393,N_42851);
xnor UO_273 (O_273,N_42068,N_49622);
xnor UO_274 (O_274,N_46262,N_49223);
nor UO_275 (O_275,N_47907,N_43817);
nand UO_276 (O_276,N_43455,N_40841);
or UO_277 (O_277,N_48127,N_49657);
nor UO_278 (O_278,N_45938,N_49091);
xnor UO_279 (O_279,N_41383,N_44537);
nand UO_280 (O_280,N_40486,N_49008);
and UO_281 (O_281,N_42489,N_45968);
nor UO_282 (O_282,N_46247,N_42166);
nor UO_283 (O_283,N_45894,N_42439);
and UO_284 (O_284,N_45998,N_40150);
nor UO_285 (O_285,N_45446,N_46695);
nor UO_286 (O_286,N_47403,N_44794);
or UO_287 (O_287,N_46519,N_40608);
nand UO_288 (O_288,N_41192,N_46194);
and UO_289 (O_289,N_41347,N_43332);
nor UO_290 (O_290,N_47688,N_45973);
nor UO_291 (O_291,N_49794,N_41338);
nand UO_292 (O_292,N_46955,N_41197);
or UO_293 (O_293,N_40104,N_47455);
nor UO_294 (O_294,N_46986,N_41369);
or UO_295 (O_295,N_45649,N_42360);
nor UO_296 (O_296,N_40603,N_40451);
nand UO_297 (O_297,N_46482,N_41846);
and UO_298 (O_298,N_48693,N_47051);
or UO_299 (O_299,N_44118,N_46809);
nand UO_300 (O_300,N_49173,N_47933);
nand UO_301 (O_301,N_47378,N_41945);
and UO_302 (O_302,N_44401,N_49298);
nor UO_303 (O_303,N_47864,N_45763);
or UO_304 (O_304,N_41168,N_43954);
nand UO_305 (O_305,N_46713,N_42526);
or UO_306 (O_306,N_42693,N_40447);
nand UO_307 (O_307,N_41461,N_49066);
or UO_308 (O_308,N_48624,N_42034);
nand UO_309 (O_309,N_42375,N_41977);
or UO_310 (O_310,N_40271,N_47290);
and UO_311 (O_311,N_40530,N_45308);
or UO_312 (O_312,N_47799,N_46720);
or UO_313 (O_313,N_45276,N_42081);
and UO_314 (O_314,N_48953,N_47182);
or UO_315 (O_315,N_41741,N_47031);
nor UO_316 (O_316,N_46816,N_49996);
nand UO_317 (O_317,N_48819,N_45738);
xnor UO_318 (O_318,N_45061,N_47737);
nor UO_319 (O_319,N_48900,N_45307);
xor UO_320 (O_320,N_45524,N_43978);
and UO_321 (O_321,N_41920,N_47719);
and UO_322 (O_322,N_40866,N_44526);
or UO_323 (O_323,N_41511,N_42742);
nand UO_324 (O_324,N_47744,N_45434);
nand UO_325 (O_325,N_42617,N_45837);
nand UO_326 (O_326,N_47052,N_43866);
and UO_327 (O_327,N_40559,N_40848);
or UO_328 (O_328,N_45320,N_40482);
nand UO_329 (O_329,N_42532,N_43117);
or UO_330 (O_330,N_40059,N_46787);
or UO_331 (O_331,N_48089,N_41410);
nand UO_332 (O_332,N_43468,N_40032);
nor UO_333 (O_333,N_47979,N_46101);
or UO_334 (O_334,N_49467,N_41753);
nand UO_335 (O_335,N_46358,N_44631);
or UO_336 (O_336,N_48586,N_49917);
and UO_337 (O_337,N_46961,N_49271);
or UO_338 (O_338,N_47329,N_45193);
or UO_339 (O_339,N_41264,N_42517);
or UO_340 (O_340,N_44388,N_43005);
or UO_341 (O_341,N_48201,N_44560);
and UO_342 (O_342,N_45504,N_41944);
and UO_343 (O_343,N_45032,N_49317);
and UO_344 (O_344,N_49226,N_42058);
or UO_345 (O_345,N_42223,N_44030);
nand UO_346 (O_346,N_42554,N_45810);
xnor UO_347 (O_347,N_43094,N_40284);
and UO_348 (O_348,N_49663,N_44875);
nor UO_349 (O_349,N_44980,N_40556);
nor UO_350 (O_350,N_45102,N_44742);
or UO_351 (O_351,N_46223,N_45205);
nand UO_352 (O_352,N_47576,N_42987);
xnor UO_353 (O_353,N_41588,N_45863);
nor UO_354 (O_354,N_45121,N_40554);
nand UO_355 (O_355,N_41195,N_46669);
nor UO_356 (O_356,N_45799,N_46032);
xnor UO_357 (O_357,N_42741,N_46968);
xnor UO_358 (O_358,N_41720,N_40944);
or UO_359 (O_359,N_43034,N_42558);
nand UO_360 (O_360,N_42909,N_41658);
or UO_361 (O_361,N_46819,N_48835);
and UO_362 (O_362,N_41206,N_40543);
nor UO_363 (O_363,N_47629,N_48573);
nand UO_364 (O_364,N_43444,N_45376);
nor UO_365 (O_365,N_45732,N_48062);
nand UO_366 (O_366,N_45509,N_46155);
nor UO_367 (O_367,N_41456,N_42412);
nor UO_368 (O_368,N_45868,N_40481);
or UO_369 (O_369,N_47819,N_42580);
nand UO_370 (O_370,N_40116,N_40987);
and UO_371 (O_371,N_46352,N_45111);
xor UO_372 (O_372,N_44511,N_42587);
or UO_373 (O_373,N_44719,N_44979);
and UO_374 (O_374,N_47873,N_44689);
nand UO_375 (O_375,N_48975,N_47554);
and UO_376 (O_376,N_46002,N_44085);
nand UO_377 (O_377,N_49580,N_47776);
xor UO_378 (O_378,N_42679,N_43715);
xnor UO_379 (O_379,N_40851,N_44208);
or UO_380 (O_380,N_40243,N_44654);
or UO_381 (O_381,N_49269,N_49214);
or UO_382 (O_382,N_48262,N_46139);
nor UO_383 (O_383,N_41025,N_43971);
nor UO_384 (O_384,N_44171,N_49138);
or UO_385 (O_385,N_40126,N_44109);
nor UO_386 (O_386,N_47856,N_44858);
or UO_387 (O_387,N_42654,N_42147);
or UO_388 (O_388,N_49478,N_48804);
or UO_389 (O_389,N_46756,N_44249);
nor UO_390 (O_390,N_46896,N_45018);
nand UO_391 (O_391,N_44866,N_46325);
or UO_392 (O_392,N_42305,N_45156);
or UO_393 (O_393,N_45667,N_40257);
nand UO_394 (O_394,N_46228,N_45066);
or UO_395 (O_395,N_49528,N_40653);
and UO_396 (O_396,N_48889,N_46694);
nor UO_397 (O_397,N_48378,N_44802);
or UO_398 (O_398,N_44297,N_49459);
nand UO_399 (O_399,N_46612,N_42369);
or UO_400 (O_400,N_48595,N_41055);
and UO_401 (O_401,N_43501,N_42640);
xnor UO_402 (O_402,N_40178,N_42026);
nor UO_403 (O_403,N_49839,N_47414);
and UO_404 (O_404,N_46204,N_41910);
nor UO_405 (O_405,N_45829,N_48174);
nor UO_406 (O_406,N_44705,N_42612);
and UO_407 (O_407,N_48293,N_41041);
and UO_408 (O_408,N_46981,N_40348);
and UO_409 (O_409,N_43188,N_43192);
or UO_410 (O_410,N_46424,N_40367);
xnor UO_411 (O_411,N_44904,N_44091);
or UO_412 (O_412,N_41379,N_43168);
nor UO_413 (O_413,N_49715,N_41784);
and UO_414 (O_414,N_44550,N_45142);
or UO_415 (O_415,N_46882,N_45839);
nand UO_416 (O_416,N_47201,N_47046);
and UO_417 (O_417,N_48261,N_40945);
nor UO_418 (O_418,N_43327,N_49092);
or UO_419 (O_419,N_49272,N_43920);
xnor UO_420 (O_420,N_47544,N_47362);
nor UO_421 (O_421,N_41585,N_43573);
nor UO_422 (O_422,N_41913,N_48651);
nand UO_423 (O_423,N_42064,N_45984);
or UO_424 (O_424,N_46966,N_45802);
nand UO_425 (O_425,N_45691,N_48259);
and UO_426 (O_426,N_46123,N_45355);
and UO_427 (O_427,N_44747,N_46798);
nor UO_428 (O_428,N_48137,N_48517);
nand UO_429 (O_429,N_49458,N_45101);
nor UO_430 (O_430,N_41220,N_45160);
nand UO_431 (O_431,N_44581,N_40909);
and UO_432 (O_432,N_41522,N_43490);
nand UO_433 (O_433,N_46333,N_41234);
or UO_434 (O_434,N_42794,N_42508);
nand UO_435 (O_435,N_42383,N_47564);
nor UO_436 (O_436,N_42572,N_42547);
xor UO_437 (O_437,N_49439,N_42073);
nor UO_438 (O_438,N_41049,N_48665);
or UO_439 (O_439,N_48119,N_41199);
and UO_440 (O_440,N_48433,N_40940);
or UO_441 (O_441,N_47529,N_43486);
nand UO_442 (O_442,N_40002,N_40737);
and UO_443 (O_443,N_40557,N_41594);
xnor UO_444 (O_444,N_43527,N_40088);
xor UO_445 (O_445,N_45072,N_40207);
and UO_446 (O_446,N_45245,N_43171);
xor UO_447 (O_447,N_43480,N_40218);
nor UO_448 (O_448,N_46303,N_41500);
nor UO_449 (O_449,N_40547,N_48865);
or UO_450 (O_450,N_48407,N_40533);
and UO_451 (O_451,N_48175,N_43397);
nand UO_452 (O_452,N_46661,N_44277);
or UO_453 (O_453,N_44435,N_47891);
xor UO_454 (O_454,N_46726,N_47498);
nor UO_455 (O_455,N_49718,N_42483);
xnor UO_456 (O_456,N_49838,N_45261);
or UO_457 (O_457,N_46160,N_47174);
xor UO_458 (O_458,N_44661,N_47197);
nor UO_459 (O_459,N_45474,N_48795);
and UO_460 (O_460,N_42107,N_46513);
nand UO_461 (O_461,N_43328,N_43916);
and UO_462 (O_462,N_47946,N_47283);
and UO_463 (O_463,N_49113,N_46535);
and UO_464 (O_464,N_47982,N_42487);
nand UO_465 (O_465,N_42763,N_40970);
and UO_466 (O_466,N_48286,N_46736);
or UO_467 (O_467,N_46776,N_48771);
xor UO_468 (O_468,N_48641,N_43930);
and UO_469 (O_469,N_47021,N_46766);
or UO_470 (O_470,N_41344,N_47383);
nand UO_471 (O_471,N_43794,N_42280);
or UO_472 (O_472,N_47224,N_44129);
and UO_473 (O_473,N_40346,N_45349);
nand UO_474 (O_474,N_42299,N_43340);
or UO_475 (O_475,N_44329,N_43922);
and UO_476 (O_476,N_40832,N_49851);
nor UO_477 (O_477,N_47905,N_42993);
or UO_478 (O_478,N_47649,N_43976);
and UO_479 (O_479,N_42638,N_47468);
xnor UO_480 (O_480,N_45847,N_40487);
nor UO_481 (O_481,N_42501,N_43326);
nor UO_482 (O_482,N_40228,N_41120);
or UO_483 (O_483,N_45244,N_42527);
or UO_484 (O_484,N_46690,N_45442);
or UO_485 (O_485,N_45042,N_41779);
nor UO_486 (O_486,N_42673,N_43061);
nor UO_487 (O_487,N_48039,N_46527);
nand UO_488 (O_488,N_42233,N_47117);
nor UO_489 (O_489,N_44744,N_44872);
xnor UO_490 (O_490,N_45670,N_46309);
and UO_491 (O_491,N_42992,N_40253);
or UO_492 (O_492,N_44941,N_46851);
nand UO_493 (O_493,N_49844,N_42943);
nand UO_494 (O_494,N_40295,N_42140);
nor UO_495 (O_495,N_48002,N_45598);
nand UO_496 (O_496,N_43807,N_45919);
xnor UO_497 (O_497,N_43653,N_46836);
and UO_498 (O_498,N_43440,N_45786);
nand UO_499 (O_499,N_48875,N_47198);
and UO_500 (O_500,N_46348,N_40393);
nor UO_501 (O_501,N_47180,N_47286);
nand UO_502 (O_502,N_47015,N_42196);
nor UO_503 (O_503,N_40734,N_48371);
nand UO_504 (O_504,N_42967,N_42376);
xor UO_505 (O_505,N_45443,N_43448);
and UO_506 (O_506,N_40439,N_46267);
nor UO_507 (O_507,N_41082,N_47586);
nand UO_508 (O_508,N_45009,N_44061);
or UO_509 (O_509,N_42373,N_45248);
nor UO_510 (O_510,N_46875,N_47391);
and UO_511 (O_511,N_43975,N_48790);
nor UO_512 (O_512,N_48751,N_45048);
nor UO_513 (O_513,N_46047,N_42361);
nand UO_514 (O_514,N_48947,N_46254);
nand UO_515 (O_515,N_45390,N_47995);
nand UO_516 (O_516,N_47213,N_41823);
or UO_517 (O_517,N_49129,N_47422);
and UO_518 (O_518,N_46902,N_42272);
xnor UO_519 (O_519,N_49722,N_44126);
or UO_520 (O_520,N_44902,N_47590);
nand UO_521 (O_521,N_45452,N_48252);
and UO_522 (O_522,N_41826,N_41482);
xnor UO_523 (O_523,N_44619,N_47622);
nand UO_524 (O_524,N_46298,N_41703);
nor UO_525 (O_525,N_46516,N_41019);
xor UO_526 (O_526,N_47328,N_47078);
nor UO_527 (O_527,N_43837,N_49843);
nand UO_528 (O_528,N_40910,N_46627);
and UO_529 (O_529,N_48749,N_46443);
nor UO_530 (O_530,N_40762,N_49418);
nor UO_531 (O_531,N_43464,N_46538);
or UO_532 (O_532,N_46956,N_47038);
and UO_533 (O_533,N_45392,N_47825);
or UO_534 (O_534,N_48896,N_48610);
nor UO_535 (O_535,N_47769,N_43752);
or UO_536 (O_536,N_46971,N_44079);
nand UO_537 (O_537,N_46366,N_48796);
nand UO_538 (O_538,N_47897,N_45301);
and UO_539 (O_539,N_46699,N_41852);
or UO_540 (O_540,N_49456,N_43445);
nor UO_541 (O_541,N_45323,N_49203);
nand UO_542 (O_542,N_43184,N_47300);
and UO_543 (O_543,N_43017,N_41629);
nand UO_544 (O_544,N_42001,N_43053);
nor UO_545 (O_545,N_44555,N_42089);
xor UO_546 (O_546,N_43110,N_43058);
xor UO_547 (O_547,N_40520,N_40984);
or UO_548 (O_548,N_43057,N_46412);
nor UO_549 (O_549,N_48232,N_44615);
or UO_550 (O_550,N_43980,N_40983);
or UO_551 (O_551,N_46655,N_40622);
xnor UO_552 (O_552,N_48027,N_45391);
or UO_553 (O_553,N_46585,N_44340);
xor UO_554 (O_554,N_44180,N_44097);
or UO_555 (O_555,N_48961,N_40952);
or UO_556 (O_556,N_49218,N_48979);
nand UO_557 (O_557,N_49991,N_43567);
and UO_558 (O_558,N_44602,N_42188);
or UO_559 (O_559,N_46417,N_41831);
xnor UO_560 (O_560,N_41519,N_47230);
and UO_561 (O_561,N_40606,N_41785);
nor UO_562 (O_562,N_45080,N_44043);
or UO_563 (O_563,N_47090,N_47957);
nand UO_564 (O_564,N_42567,N_43804);
or UO_565 (O_565,N_45327,N_40813);
nand UO_566 (O_566,N_40615,N_40338);
and UO_567 (O_567,N_47235,N_41654);
and UO_568 (O_568,N_40416,N_46892);
xor UO_569 (O_569,N_42768,N_44638);
nand UO_570 (O_570,N_43656,N_49219);
nor UO_571 (O_571,N_47029,N_42437);
and UO_572 (O_572,N_47840,N_41479);
and UO_573 (O_573,N_46963,N_48650);
nor UO_574 (O_574,N_47604,N_44544);
and UO_575 (O_575,N_45884,N_45828);
or UO_576 (O_576,N_48337,N_42861);
nor UO_577 (O_577,N_42521,N_47001);
or UO_578 (O_578,N_41820,N_41994);
and UO_579 (O_579,N_41054,N_49549);
nand UO_580 (O_580,N_48011,N_44737);
nand UO_581 (O_581,N_47866,N_42799);
nand UO_582 (O_582,N_48776,N_44334);
xnor UO_583 (O_583,N_46528,N_46141);
or UO_584 (O_584,N_44846,N_42154);
or UO_585 (O_585,N_49699,N_40185);
or UO_586 (O_586,N_42738,N_43082);
nor UO_587 (O_587,N_48489,N_47826);
and UO_588 (O_588,N_40997,N_40660);
xor UO_589 (O_589,N_47319,N_40740);
or UO_590 (O_590,N_45478,N_45492);
and UO_591 (O_591,N_40052,N_42101);
or UO_592 (O_592,N_45186,N_43115);
nand UO_593 (O_593,N_44330,N_45264);
and UO_594 (O_594,N_47010,N_43477);
and UO_595 (O_595,N_42368,N_42273);
and UO_596 (O_596,N_44896,N_46932);
nor UO_597 (O_597,N_42266,N_48090);
and UO_598 (O_598,N_49209,N_45380);
and UO_599 (O_599,N_40745,N_49085);
xor UO_600 (O_600,N_46643,N_41084);
nand UO_601 (O_601,N_44928,N_43600);
or UO_602 (O_602,N_47666,N_44493);
and UO_603 (O_603,N_48719,N_48128);
or UO_604 (O_604,N_47110,N_46570);
or UO_605 (O_605,N_46171,N_43054);
or UO_606 (O_606,N_47237,N_47704);
and UO_607 (O_607,N_45526,N_48311);
or UO_608 (O_608,N_48296,N_48083);
xnor UO_609 (O_609,N_47176,N_49989);
nor UO_610 (O_610,N_40887,N_42541);
or UO_611 (O_611,N_49727,N_45124);
or UO_612 (O_612,N_43295,N_40564);
or UO_613 (O_613,N_45615,N_46030);
and UO_614 (O_614,N_42787,N_42821);
xor UO_615 (O_615,N_46979,N_44140);
nand UO_616 (O_616,N_47857,N_48335);
or UO_617 (O_617,N_42938,N_48298);
nor UO_618 (O_618,N_49744,N_45268);
or UO_619 (O_619,N_41795,N_41691);
nor UO_620 (O_620,N_42079,N_47234);
nand UO_621 (O_621,N_49958,N_47248);
nand UO_622 (O_622,N_42914,N_40550);
nor UO_623 (O_623,N_41215,N_43830);
nor UO_624 (O_624,N_40260,N_41067);
and UO_625 (O_625,N_48954,N_40682);
and UO_626 (O_626,N_45352,N_45249);
nor UO_627 (O_627,N_47361,N_43893);
and UO_628 (O_628,N_43157,N_40787);
nor UO_629 (O_629,N_47293,N_47070);
nor UO_630 (O_630,N_46054,N_44525);
and UO_631 (O_631,N_44817,N_42382);
nand UO_632 (O_632,N_44662,N_41458);
nor UO_633 (O_633,N_48471,N_49971);
and UO_634 (O_634,N_46406,N_44448);
nand UO_635 (O_635,N_47164,N_41191);
nor UO_636 (O_636,N_45618,N_47126);
or UO_637 (O_637,N_48374,N_45561);
nor UO_638 (O_638,N_46452,N_48073);
and UO_639 (O_639,N_47012,N_46747);
and UO_640 (O_640,N_40937,N_46203);
or UO_641 (O_641,N_40494,N_45337);
or UO_642 (O_642,N_40109,N_47695);
and UO_643 (O_643,N_49014,N_46953);
and UO_644 (O_644,N_42259,N_45022);
nand UO_645 (O_645,N_48441,N_45295);
nand UO_646 (O_646,N_47311,N_43281);
or UO_647 (O_647,N_48753,N_44868);
xor UO_648 (O_648,N_46997,N_43228);
nand UO_649 (O_649,N_41657,N_41941);
and UO_650 (O_650,N_42894,N_46293);
nand UO_651 (O_651,N_43145,N_45539);
nand UO_652 (O_652,N_43887,N_46495);
and UO_653 (O_653,N_49542,N_40863);
and UO_654 (O_654,N_45385,N_44853);
nor UO_655 (O_655,N_44961,N_45765);
nor UO_656 (O_656,N_45275,N_41506);
and UO_657 (O_657,N_48942,N_45104);
and UO_658 (O_658,N_41819,N_48167);
xnor UO_659 (O_659,N_47822,N_43626);
or UO_660 (O_660,N_42467,N_44540);
nand UO_661 (O_661,N_44294,N_49126);
or UO_662 (O_662,N_49833,N_47896);
and UO_663 (O_663,N_44236,N_40441);
and UO_664 (O_664,N_41551,N_41508);
and UO_665 (O_665,N_41155,N_41707);
or UO_666 (O_666,N_41792,N_47387);
nor UO_667 (O_667,N_40858,N_43662);
nor UO_668 (O_668,N_48410,N_47192);
nand UO_669 (O_669,N_49147,N_49168);
nor UO_670 (O_670,N_45226,N_42120);
nand UO_671 (O_671,N_45484,N_49773);
nor UO_672 (O_672,N_47643,N_46301);
and UO_673 (O_673,N_42245,N_40118);
xnor UO_674 (O_674,N_43210,N_41187);
or UO_675 (O_675,N_44433,N_47085);
or UO_676 (O_676,N_42379,N_49353);
or UO_677 (O_677,N_46978,N_47123);
nor UO_678 (O_678,N_41494,N_42836);
and UO_679 (O_679,N_44570,N_46457);
nor UO_680 (O_680,N_45627,N_42637);
or UO_681 (O_681,N_49901,N_48068);
and UO_682 (O_682,N_49259,N_45051);
and UO_683 (O_683,N_46881,N_42505);
and UO_684 (O_684,N_47265,N_45921);
or UO_685 (O_685,N_40251,N_45039);
xor UO_686 (O_686,N_49227,N_43453);
nand UO_687 (O_687,N_49638,N_41706);
and UO_688 (O_688,N_41608,N_47053);
and UO_689 (O_689,N_49734,N_47351);
nor UO_690 (O_690,N_40536,N_40781);
or UO_691 (O_691,N_43515,N_44732);
nand UO_692 (O_692,N_42080,N_42330);
nor UO_693 (O_693,N_42074,N_44890);
nand UO_694 (O_694,N_46630,N_44179);
or UO_695 (O_695,N_40475,N_42121);
or UO_696 (O_696,N_46624,N_46752);
nor UO_697 (O_697,N_45979,N_45204);
nor UO_698 (O_698,N_44027,N_47282);
or UO_699 (O_699,N_43011,N_40350);
xor UO_700 (O_700,N_46488,N_44717);
and UO_701 (O_701,N_43696,N_40471);
nor UO_702 (O_702,N_45648,N_45334);
or UO_703 (O_703,N_41357,N_48461);
nor UO_704 (O_704,N_47222,N_44190);
nand UO_705 (O_705,N_47813,N_49872);
or UO_706 (O_706,N_49038,N_46939);
or UO_707 (O_707,N_48692,N_41561);
xor UO_708 (O_708,N_47006,N_47189);
nor UO_709 (O_709,N_48826,N_49405);
nor UO_710 (O_710,N_43215,N_45293);
nand UO_711 (O_711,N_43489,N_44244);
nand UO_712 (O_712,N_43261,N_45558);
or UO_713 (O_713,N_41873,N_45356);
and UO_714 (O_714,N_40061,N_41812);
and UO_715 (O_715,N_44288,N_44016);
xnor UO_716 (O_716,N_48629,N_46245);
nor UO_717 (O_717,N_45095,N_42193);
nand UO_718 (O_718,N_42445,N_49899);
and UO_719 (O_719,N_45218,N_44477);
nor UO_720 (O_720,N_40143,N_46185);
and UO_721 (O_721,N_47517,N_41609);
nand UO_722 (O_722,N_46941,N_47095);
or UO_723 (O_723,N_47430,N_42009);
or UO_724 (O_724,N_48748,N_48026);
nand UO_725 (O_725,N_48281,N_40064);
and UO_726 (O_726,N_44347,N_46868);
and UO_727 (O_727,N_48578,N_46925);
or UO_728 (O_728,N_48233,N_43580);
or UO_729 (O_729,N_41876,N_47796);
and UO_730 (O_730,N_43849,N_42028);
or UO_731 (O_731,N_44077,N_43667);
or UO_732 (O_732,N_43763,N_44757);
nand UO_733 (O_733,N_41743,N_49410);
or UO_734 (O_734,N_47865,N_44740);
or UO_735 (O_735,N_44071,N_46041);
or UO_736 (O_736,N_40324,N_44812);
and UO_737 (O_737,N_45874,N_49890);
and UO_738 (O_738,N_47909,N_47303);
nor UO_739 (O_739,N_48255,N_49392);
nand UO_740 (O_740,N_44217,N_41076);
nor UO_741 (O_741,N_45947,N_42449);
or UO_742 (O_742,N_44736,N_45818);
or UO_743 (O_743,N_42407,N_48052);
nand UO_744 (O_744,N_44437,N_47431);
and UO_745 (O_745,N_48894,N_43851);
nand UO_746 (O_746,N_43150,N_42017);
and UO_747 (O_747,N_45306,N_49742);
and UO_748 (O_748,N_49378,N_46739);
nor UO_749 (O_749,N_44471,N_44020);
nand UO_750 (O_750,N_42337,N_48998);
or UO_751 (O_751,N_42128,N_45935);
xor UO_752 (O_752,N_47523,N_42189);
nand UO_753 (O_753,N_42030,N_40086);
nand UO_754 (O_754,N_42341,N_46322);
xnor UO_755 (O_755,N_41005,N_41647);
nand UO_756 (O_756,N_42977,N_48870);
nand UO_757 (O_757,N_48890,N_47731);
nand UO_758 (O_758,N_43159,N_47928);
nand UO_759 (O_759,N_48080,N_45950);
or UO_760 (O_760,N_48423,N_40574);
xor UO_761 (O_761,N_47400,N_49853);
or UO_762 (O_762,N_46543,N_43216);
nand UO_763 (O_763,N_40809,N_45339);
or UO_764 (O_764,N_45612,N_42846);
nor UO_765 (O_765,N_48643,N_45571);
and UO_766 (O_766,N_47560,N_45168);
or UO_767 (O_767,N_40026,N_40688);
nand UO_768 (O_768,N_43739,N_46717);
nand UO_769 (O_769,N_42157,N_47060);
and UO_770 (O_770,N_46813,N_47512);
nor UO_771 (O_771,N_43088,N_40972);
nand UO_772 (O_772,N_42970,N_40753);
nand UO_773 (O_773,N_47665,N_47787);
nor UO_774 (O_774,N_46754,N_47869);
or UO_775 (O_775,N_46866,N_45663);
or UO_776 (O_776,N_45741,N_45021);
or UO_777 (O_777,N_42806,N_41679);
nand UO_778 (O_778,N_43825,N_47459);
nor UO_779 (O_779,N_45548,N_47423);
or UO_780 (O_780,N_47918,N_44546);
or UO_781 (O_781,N_40396,N_42148);
nand UO_782 (O_782,N_44176,N_44063);
or UO_783 (O_783,N_49629,N_40862);
and UO_784 (O_784,N_49904,N_47138);
and UO_785 (O_785,N_40410,N_44172);
or UO_786 (O_786,N_40828,N_49096);
xnor UO_787 (O_787,N_46104,N_46211);
nand UO_788 (O_788,N_40167,N_46581);
nor UO_789 (O_789,N_48035,N_48196);
nand UO_790 (O_790,N_48076,N_44995);
nor UO_791 (O_791,N_46323,N_43740);
nand UO_792 (O_792,N_41627,N_44031);
and UO_793 (O_793,N_44321,N_44869);
nor UO_794 (O_794,N_40823,N_41354);
and UO_795 (O_795,N_43728,N_45453);
nor UO_796 (O_796,N_42999,N_49376);
or UO_797 (O_797,N_40896,N_48647);
and UO_798 (O_798,N_41047,N_49240);
or UO_799 (O_799,N_41591,N_44975);
nand UO_800 (O_800,N_40950,N_47655);
xnor UO_801 (O_801,N_49028,N_47450);
nand UO_802 (O_802,N_40034,N_45901);
and UO_803 (O_803,N_44078,N_45983);
or UO_804 (O_804,N_43335,N_48190);
or UO_805 (O_805,N_48421,N_43770);
nand UO_806 (O_806,N_40373,N_44735);
or UO_807 (O_807,N_48077,N_49055);
or UO_808 (O_808,N_49065,N_47132);
xnor UO_809 (O_809,N_46814,N_42729);
nor UO_810 (O_810,N_48189,N_49040);
or UO_811 (O_811,N_44965,N_41899);
nor UO_812 (O_812,N_49831,N_43719);
or UO_813 (O_813,N_40186,N_43929);
nor UO_814 (O_814,N_40650,N_45626);
or UO_815 (O_815,N_47089,N_41587);
nor UO_816 (O_816,N_49005,N_42962);
nand UO_817 (O_817,N_48861,N_48381);
nor UO_818 (O_818,N_40593,N_43660);
nand UO_819 (O_819,N_46216,N_45235);
or UO_820 (O_820,N_49749,N_42197);
xnor UO_821 (O_821,N_42808,N_42456);
nor UO_822 (O_822,N_49352,N_49330);
nand UO_823 (O_823,N_48871,N_42747);
and UO_824 (O_824,N_43608,N_42983);
or UO_825 (O_825,N_42210,N_42765);
or UO_826 (O_826,N_40518,N_42869);
and UO_827 (O_827,N_40996,N_42651);
or UO_828 (O_828,N_42759,N_49182);
or UO_829 (O_829,N_44573,N_47255);
and UO_830 (O_830,N_40774,N_48392);
nor UO_831 (O_831,N_41902,N_44752);
nor UO_832 (O_832,N_40361,N_46163);
nor UO_833 (O_833,N_41075,N_48626);
or UO_834 (O_834,N_45384,N_45592);
nand UO_835 (O_835,N_47924,N_40919);
xor UO_836 (O_836,N_41023,N_45959);
nand UO_837 (O_837,N_44710,N_44963);
xnor UO_838 (O_838,N_48824,N_45325);
nand UO_839 (O_839,N_47063,N_49604);
xor UO_840 (O_840,N_48256,N_44942);
nand UO_841 (O_841,N_43709,N_42020);
and UO_842 (O_842,N_41537,N_43757);
or UO_843 (O_843,N_41923,N_40674);
xor UO_844 (O_844,N_41401,N_47756);
nand UO_845 (O_845,N_47273,N_42399);
nand UO_846 (O_846,N_48858,N_42907);
or UO_847 (O_847,N_43732,N_42136);
nor UO_848 (O_848,N_41095,N_49581);
nand UO_849 (O_849,N_41993,N_49704);
nand UO_850 (O_850,N_41782,N_41062);
and UO_851 (O_851,N_46750,N_41930);
and UO_852 (O_852,N_47364,N_41426);
and UO_853 (O_853,N_49425,N_48652);
or UO_854 (O_854,N_47860,N_48422);
nor UO_855 (O_855,N_43675,N_46658);
nand UO_856 (O_856,N_41690,N_47981);
or UO_857 (O_857,N_43222,N_41619);
or UO_858 (O_858,N_46378,N_41130);
xor UO_859 (O_859,N_46514,N_44644);
nand UO_860 (O_860,N_47045,N_42349);
or UO_861 (O_861,N_40081,N_41287);
and UO_862 (O_862,N_42573,N_41767);
nand UO_863 (O_863,N_48536,N_46602);
or UO_864 (O_864,N_41372,N_40231);
nor UO_865 (O_865,N_48166,N_42625);
and UO_866 (O_866,N_45329,N_46733);
nor UO_867 (O_867,N_46614,N_46879);
nand UO_868 (O_868,N_40128,N_47062);
and UO_869 (O_869,N_43531,N_47802);
and UO_870 (O_870,N_43970,N_46948);
nand UO_871 (O_871,N_45368,N_44021);
and UO_872 (O_872,N_47170,N_42238);
or UO_873 (O_873,N_42618,N_46043);
nand UO_874 (O_874,N_44225,N_48520);
and UO_875 (O_875,N_46933,N_47205);
or UO_876 (O_876,N_45619,N_42012);
and UO_877 (O_877,N_46050,N_41111);
or UO_878 (O_878,N_41735,N_49504);
xnor UO_879 (O_879,N_49922,N_48676);
or UO_880 (O_880,N_49664,N_41415);
or UO_881 (O_881,N_41053,N_48882);
xor UO_882 (O_882,N_49123,N_48677);
and UO_883 (O_883,N_48012,N_42717);
nor UO_884 (O_884,N_46522,N_47464);
nor UO_885 (O_885,N_42355,N_41108);
nand UO_886 (O_886,N_42591,N_49977);
nor UO_887 (O_887,N_44931,N_43986);
or UO_888 (O_888,N_44421,N_40663);
xnor UO_889 (O_889,N_45081,N_44407);
nor UO_890 (O_890,N_43428,N_49671);
and UO_891 (O_891,N_47218,N_41700);
or UO_892 (O_892,N_44913,N_46354);
nand UO_893 (O_893,N_41781,N_46423);
or UO_894 (O_894,N_42108,N_42228);
and UO_895 (O_895,N_43597,N_48032);
and UO_896 (O_896,N_44089,N_45253);
or UO_897 (O_897,N_41214,N_42339);
xor UO_898 (O_898,N_42477,N_43331);
nand UO_899 (O_899,N_45298,N_45668);
nor UO_900 (O_900,N_47854,N_48144);
or UO_901 (O_901,N_45928,N_42442);
xor UO_902 (O_902,N_42766,N_41433);
and UO_903 (O_903,N_45678,N_46157);
or UO_904 (O_904,N_46074,N_46279);
nand UO_905 (O_905,N_47993,N_46382);
or UO_906 (O_906,N_40247,N_41274);
nor UO_907 (O_907,N_48521,N_40750);
nor UO_908 (O_908,N_44455,N_42814);
or UO_909 (O_909,N_46052,N_40926);
nand UO_910 (O_910,N_41742,N_45572);
nand UO_911 (O_911,N_40200,N_45211);
nor UO_912 (O_912,N_48814,N_40467);
nor UO_913 (O_913,N_43664,N_45853);
and UO_914 (O_914,N_49913,N_48341);
or UO_915 (O_915,N_49941,N_47134);
nor UO_916 (O_916,N_42706,N_48817);
and UO_917 (O_917,N_44429,N_41170);
nor UO_918 (O_918,N_47579,N_47878);
or UO_919 (O_919,N_47591,N_47914);
and UO_920 (O_920,N_47416,N_44910);
nor UO_921 (O_921,N_45015,N_46817);
or UO_922 (O_922,N_48560,N_46873);
nand UO_923 (O_923,N_44131,N_48915);
nor UO_924 (O_924,N_40842,N_45502);
and UO_925 (O_925,N_47445,N_44988);
and UO_926 (O_926,N_45239,N_47667);
nor UO_927 (O_927,N_41530,N_41417);
nor UO_928 (O_928,N_40894,N_49946);
nor UO_929 (O_929,N_46786,N_40385);
or UO_930 (O_930,N_43957,N_46751);
nand UO_931 (O_931,N_44218,N_44630);
nor UO_932 (O_932,N_44527,N_42235);
and UO_933 (O_933,N_47920,N_40613);
xnor UO_934 (O_934,N_41306,N_43361);
or UO_935 (O_935,N_43681,N_43948);
nor UO_936 (O_936,N_40192,N_42211);
nand UO_937 (O_937,N_41915,N_45362);
or UO_938 (O_938,N_41514,N_49443);
or UO_939 (O_939,N_44125,N_41988);
nor UO_940 (O_940,N_47435,N_42877);
and UO_941 (O_941,N_47721,N_44697);
and UO_942 (O_942,N_49069,N_43864);
nor UO_943 (O_943,N_45562,N_40964);
or UO_944 (O_944,N_45012,N_45400);
nor UO_945 (O_945,N_48377,N_45735);
and UO_946 (O_946,N_47702,N_49907);
nor UO_947 (O_947,N_44884,N_49480);
or UO_948 (O_948,N_47146,N_44099);
nand UO_949 (O_949,N_41620,N_49484);
nand UO_950 (O_950,N_46577,N_46476);
nor UO_951 (O_951,N_44645,N_45693);
nor UO_952 (O_952,N_45920,N_40458);
nor UO_953 (O_953,N_49985,N_47221);
nor UO_954 (O_954,N_41467,N_49262);
nand UO_955 (O_955,N_45888,N_42905);
or UO_956 (O_956,N_48314,N_43153);
nand UO_957 (O_957,N_49109,N_41255);
and UO_958 (O_958,N_42455,N_45098);
and UO_959 (O_959,N_42988,N_43079);
nand UO_960 (O_960,N_49589,N_45154);
and UO_961 (O_961,N_45472,N_43095);
nor UO_962 (O_962,N_44936,N_47102);
nor UO_963 (O_963,N_40223,N_45908);
nand UO_964 (O_964,N_48437,N_41373);
or UO_965 (O_965,N_42297,N_42919);
nor UO_966 (O_966,N_42046,N_49705);
nand UO_967 (O_967,N_48114,N_43347);
nand UO_968 (O_968,N_47740,N_41603);
nor UO_969 (O_969,N_40029,N_41015);
or UO_970 (O_970,N_44349,N_44480);
and UO_971 (O_971,N_46824,N_49541);
nor UO_972 (O_972,N_44864,N_43591);
and UO_973 (O_973,N_48195,N_44469);
nor UO_974 (O_974,N_48593,N_48219);
nand UO_975 (O_975,N_44826,N_46549);
or UO_976 (O_976,N_40301,N_40981);
nor UO_977 (O_977,N_48005,N_42699);
nor UO_978 (O_978,N_41683,N_40095);
and UO_979 (O_979,N_42843,N_41457);
nor UO_980 (O_980,N_42720,N_48303);
or UO_981 (O_981,N_44849,N_42665);
nand UO_982 (O_982,N_48897,N_40133);
xnor UO_983 (O_983,N_41895,N_40699);
nand UO_984 (O_984,N_41477,N_46789);
nand UO_985 (O_985,N_44301,N_40048);
nand UO_986 (O_986,N_46367,N_47142);
nor UO_987 (O_987,N_41216,N_42888);
nand UO_988 (O_988,N_40226,N_42248);
nor UO_989 (O_989,N_46377,N_49559);
or UO_990 (O_990,N_47048,N_45411);
nor UO_991 (O_991,N_45647,N_40876);
nand UO_992 (O_992,N_40401,N_48964);
or UO_993 (O_993,N_41466,N_47030);
nor UO_994 (O_994,N_42377,N_46448);
and UO_995 (O_995,N_43279,N_42860);
or UO_996 (O_996,N_41453,N_48169);
or UO_997 (O_997,N_40905,N_45962);
xor UO_998 (O_998,N_44191,N_43346);
and UO_999 (O_999,N_45789,N_41878);
and UO_1000 (O_1000,N_45547,N_43774);
nor UO_1001 (O_1001,N_41493,N_48660);
and UO_1002 (O_1002,N_48888,N_42342);
xnor UO_1003 (O_1003,N_43321,N_48778);
or UO_1004 (O_1004,N_45644,N_40169);
or UO_1005 (O_1005,N_49660,N_43582);
nor UO_1006 (O_1006,N_41260,N_40664);
nand UO_1007 (O_1007,N_46013,N_48939);
nor UO_1008 (O_1008,N_42214,N_41841);
nor UO_1009 (O_1009,N_43935,N_48874);
or UO_1010 (O_1010,N_45234,N_46487);
nor UO_1011 (O_1011,N_44727,N_40889);
or UO_1012 (O_1012,N_42024,N_40474);
nand UO_1013 (O_1013,N_45426,N_43306);
xor UO_1014 (O_1014,N_42187,N_46973);
nand UO_1015 (O_1015,N_41697,N_46936);
or UO_1016 (O_1016,N_48878,N_43915);
nor UO_1017 (O_1017,N_40974,N_44575);
or UO_1018 (O_1018,N_40013,N_48282);
nand UO_1019 (O_1019,N_40320,N_41687);
nor UO_1020 (O_1020,N_46116,N_46550);
and UO_1021 (O_1021,N_46533,N_45977);
nand UO_1022 (O_1022,N_47888,N_45565);
and UO_1023 (O_1023,N_43824,N_49191);
nor UO_1024 (O_1024,N_42695,N_47759);
or UO_1025 (O_1025,N_40122,N_41481);
or UO_1026 (O_1026,N_40060,N_44760);
and UO_1027 (O_1027,N_47505,N_47971);
and UO_1028 (O_1028,N_45737,N_43996);
and UO_1029 (O_1029,N_48716,N_47317);
and UO_1030 (O_1030,N_41593,N_48843);
and UO_1031 (O_1031,N_40668,N_42854);
and UO_1032 (O_1032,N_42609,N_43272);
nand UO_1033 (O_1033,N_40085,N_41300);
and UO_1034 (O_1034,N_44625,N_45139);
or UO_1035 (O_1035,N_49070,N_43840);
nand UO_1036 (O_1036,N_44214,N_46682);
and UO_1037 (O_1037,N_40199,N_44847);
and UO_1038 (O_1038,N_44453,N_47959);
nor UO_1039 (O_1039,N_42354,N_42725);
xnor UO_1040 (O_1040,N_44611,N_45194);
nand UO_1041 (O_1041,N_44009,N_45360);
and UO_1042 (O_1042,N_49128,N_48515);
nand UO_1043 (O_1043,N_42599,N_46988);
nor UO_1044 (O_1044,N_45196,N_47209);
and UO_1045 (O_1045,N_45055,N_45444);
and UO_1046 (O_1046,N_40112,N_48464);
nor UO_1047 (O_1047,N_47471,N_40265);
nand UO_1048 (O_1048,N_48791,N_41147);
nor UO_1049 (O_1049,N_40532,N_40020);
xnor UO_1050 (O_1050,N_41801,N_42265);
xnor UO_1051 (O_1051,N_48666,N_43612);
nor UO_1052 (O_1052,N_48054,N_42406);
nand UO_1053 (O_1053,N_47309,N_40056);
nor UO_1054 (O_1054,N_49457,N_44926);
xor UO_1055 (O_1055,N_44394,N_41643);
nor UO_1056 (O_1056,N_49379,N_41787);
or UO_1057 (O_1057,N_42438,N_43488);
or UO_1058 (O_1058,N_42764,N_41850);
or UO_1059 (O_1059,N_41961,N_45867);
and UO_1060 (O_1060,N_42875,N_40281);
and UO_1061 (O_1061,N_45207,N_44999);
nor UO_1062 (O_1062,N_46106,N_41505);
nand UO_1063 (O_1063,N_47545,N_41434);
nor UO_1064 (O_1064,N_41018,N_46840);
and UO_1065 (O_1065,N_46328,N_43703);
or UO_1066 (O_1066,N_40931,N_49569);
or UO_1067 (O_1067,N_43146,N_48191);
nand UO_1068 (O_1068,N_46604,N_42133);
and UO_1069 (O_1069,N_40957,N_45817);
nand UO_1070 (O_1070,N_41079,N_41193);
nor UO_1071 (O_1071,N_49951,N_41268);
and UO_1072 (O_1072,N_48136,N_42276);
nor UO_1073 (O_1073,N_42839,N_47515);
nand UO_1074 (O_1074,N_48822,N_42366);
nand UO_1075 (O_1075,N_49287,N_48450);
and UO_1076 (O_1076,N_46783,N_45896);
or UO_1077 (O_1077,N_40703,N_40545);
nor UO_1078 (O_1078,N_42522,N_42236);
nand UO_1079 (O_1079,N_45028,N_48434);
nor UO_1080 (O_1080,N_42003,N_41110);
or UO_1081 (O_1081,N_41044,N_44378);
xnor UO_1082 (O_1082,N_40852,N_41889);
or UO_1083 (O_1083,N_42380,N_45610);
nor UO_1084 (O_1084,N_44258,N_49039);
nand UO_1085 (O_1085,N_41370,N_47476);
and UO_1086 (O_1086,N_45333,N_46130);
nor UO_1087 (O_1087,N_46770,N_42862);
and UO_1088 (O_1088,N_45026,N_49302);
nand UO_1089 (O_1089,N_48006,N_42705);
nor UO_1090 (O_1090,N_46906,N_45940);
xor UO_1091 (O_1091,N_44952,N_41931);
nand UO_1092 (O_1092,N_47785,N_42388);
and UO_1093 (O_1093,N_42728,N_41118);
and UO_1094 (O_1094,N_42163,N_44905);
or UO_1095 (O_1095,N_41435,N_47953);
xnor UO_1096 (O_1096,N_47711,N_44361);
or UO_1097 (O_1097,N_49969,N_43572);
or UO_1098 (O_1098,N_40799,N_46547);
xor UO_1099 (O_1099,N_45907,N_43936);
nand UO_1100 (O_1100,N_47204,N_42320);
or UO_1101 (O_1101,N_49975,N_49333);
or UO_1102 (O_1102,N_43301,N_46484);
and UO_1103 (O_1103,N_47233,N_43846);
xor UO_1104 (O_1104,N_40582,N_46026);
or UO_1105 (O_1105,N_41887,N_46069);
nor UO_1106 (O_1106,N_49534,N_43630);
nand UO_1107 (O_1107,N_47250,N_46189);
and UO_1108 (O_1108,N_44595,N_49650);
nand UO_1109 (O_1109,N_44034,N_46231);
or UO_1110 (O_1110,N_48940,N_42575);
nand UO_1111 (O_1111,N_43025,N_47771);
and UO_1112 (O_1112,N_40834,N_46773);
nor UO_1113 (O_1113,N_40424,N_47760);
or UO_1114 (O_1114,N_43174,N_43596);
and UO_1115 (O_1115,N_43260,N_43151);
xnor UO_1116 (O_1116,N_43543,N_48856);
or UO_1117 (O_1117,N_41058,N_44406);
nand UO_1118 (O_1118,N_46149,N_48644);
nor UO_1119 (O_1119,N_45956,N_40182);
and UO_1120 (O_1120,N_41570,N_42200);
or UO_1121 (O_1121,N_48494,N_45177);
or UO_1122 (O_1122,N_45137,N_46456);
nor UO_1123 (O_1123,N_41366,N_44770);
nor UO_1124 (O_1124,N_47931,N_49020);
and UO_1125 (O_1125,N_44372,N_42677);
nand UO_1126 (O_1126,N_49822,N_46019);
nor UO_1127 (O_1127,N_41744,N_45774);
nor UO_1128 (O_1128,N_43538,N_42100);
and UO_1129 (O_1129,N_43561,N_46251);
xor UO_1130 (O_1130,N_45725,N_40671);
or UO_1131 (O_1131,N_42347,N_47227);
nor UO_1132 (O_1132,N_48924,N_40001);
nor UO_1133 (O_1133,N_41166,N_42966);
xnor UO_1134 (O_1134,N_45752,N_45855);
nor UO_1135 (O_1135,N_46078,N_47797);
and UO_1136 (O_1136,N_45184,N_40428);
nand UO_1137 (O_1137,N_41364,N_45519);
nand UO_1138 (O_1138,N_49537,N_49661);
nand UO_1139 (O_1139,N_47527,N_45155);
or UO_1140 (O_1140,N_45312,N_45281);
nand UO_1141 (O_1141,N_42639,N_41388);
or UO_1142 (O_1142,N_46270,N_47846);
xor UO_1143 (O_1143,N_41185,N_47469);
nor UO_1144 (O_1144,N_46435,N_42704);
nand UO_1145 (O_1145,N_49207,N_44810);
nor UO_1146 (O_1146,N_45981,N_41837);
or UO_1147 (O_1147,N_48063,N_48157);
or UO_1148 (O_1148,N_41521,N_44175);
nor UO_1149 (O_1149,N_44405,N_46055);
and UO_1150 (O_1150,N_45936,N_41992);
nand UO_1151 (O_1151,N_49015,N_43892);
nor UO_1152 (O_1152,N_42669,N_40144);
nor UO_1153 (O_1153,N_40795,N_45159);
nor UO_1154 (O_1154,N_42653,N_43233);
nor UO_1155 (O_1155,N_42416,N_48004);
or UO_1156 (O_1156,N_45041,N_45259);
nand UO_1157 (O_1157,N_42569,N_47585);
and UO_1158 (O_1158,N_45632,N_43045);
or UO_1159 (O_1159,N_41262,N_49700);
nand UO_1160 (O_1160,N_42545,N_49998);
xnor UO_1161 (O_1161,N_45890,N_43334);
or UO_1162 (O_1162,N_45263,N_41938);
nand UO_1163 (O_1163,N_40148,N_49870);
or UO_1164 (O_1164,N_48699,N_41772);
and UO_1165 (O_1165,N_41783,N_41418);
and UO_1166 (O_1166,N_42312,N_43194);
nor UO_1167 (O_1167,N_41038,N_41269);
nor UO_1168 (O_1168,N_43549,N_44044);
xnor UO_1169 (O_1169,N_46964,N_43694);
and UO_1170 (O_1170,N_43666,N_41768);
nor UO_1171 (O_1171,N_42138,N_43938);
or UO_1172 (O_1172,N_48704,N_48829);
or UO_1173 (O_1173,N_48182,N_44283);
or UO_1174 (O_1174,N_48164,N_42542);
and UO_1175 (O_1175,N_46621,N_44424);
nor UO_1176 (O_1176,N_46889,N_47168);
and UO_1177 (O_1177,N_47727,N_40220);
nor UO_1178 (O_1178,N_42615,N_45841);
nor UO_1179 (O_1179,N_44215,N_48669);
nor UO_1180 (O_1180,N_44666,N_42585);
xnor UO_1181 (O_1181,N_45531,N_47998);
nand UO_1182 (O_1182,N_45872,N_47271);
nand UO_1183 (O_1183,N_43250,N_40273);
xor UO_1184 (O_1184,N_47342,N_40731);
nor UO_1185 (O_1185,N_44798,N_43826);
nand UO_1186 (O_1186,N_44226,N_41569);
or UO_1187 (O_1187,N_40254,N_47701);
nor UO_1188 (O_1188,N_45359,N_41851);
nand UO_1189 (O_1189,N_45379,N_49252);
or UO_1190 (O_1190,N_49151,N_40715);
or UO_1191 (O_1191,N_40277,N_44092);
and UO_1192 (O_1192,N_48096,N_40567);
nor UO_1193 (O_1193,N_45553,N_41888);
xor UO_1194 (O_1194,N_43234,N_49862);
nor UO_1195 (O_1195,N_42727,N_43676);
or UO_1196 (O_1196,N_48040,N_49397);
nor UO_1197 (O_1197,N_44387,N_47034);
or UO_1198 (O_1198,N_44449,N_49525);
nand UO_1199 (O_1199,N_44761,N_41546);
and UO_1200 (O_1200,N_46005,N_41445);
nand UO_1201 (O_1201,N_45525,N_46995);
or UO_1202 (O_1202,N_44383,N_45047);
and UO_1203 (O_1203,N_44422,N_44261);
xnor UO_1204 (O_1204,N_40625,N_40669);
nand UO_1205 (O_1205,N_46506,N_49245);
nor UO_1206 (O_1206,N_40540,N_41919);
xnor UO_1207 (O_1207,N_44927,N_47118);
nor UO_1208 (O_1208,N_42288,N_40569);
and UO_1209 (O_1209,N_44184,N_45749);
or UO_1210 (O_1210,N_41333,N_40097);
or UO_1211 (O_1211,N_47306,N_40892);
nand UO_1212 (O_1212,N_48078,N_40713);
and UO_1213 (O_1213,N_45250,N_41660);
nand UO_1214 (O_1214,N_44545,N_48885);
nand UO_1215 (O_1215,N_44313,N_41802);
nor UO_1216 (O_1216,N_47987,N_44293);
nor UO_1217 (O_1217,N_44571,N_44076);
and UO_1218 (O_1218,N_42935,N_43152);
or UO_1219 (O_1219,N_47101,N_41443);
nor UO_1220 (O_1220,N_46771,N_47565);
nand UO_1221 (O_1221,N_41816,N_45736);
nand UO_1222 (O_1222,N_43416,N_48873);
nor UO_1223 (O_1223,N_49585,N_46855);
and UO_1224 (O_1224,N_43307,N_42324);
and UO_1225 (O_1225,N_41709,N_45336);
and UO_1226 (O_1226,N_47594,N_49691);
and UO_1227 (O_1227,N_40847,N_45620);
xor UO_1228 (O_1228,N_41972,N_42566);
nor UO_1229 (O_1229,N_44291,N_44366);
nor UO_1230 (O_1230,N_47668,N_44112);
and UO_1231 (O_1231,N_41698,N_47849);
nor UO_1232 (O_1232,N_49908,N_48507);
nor UO_1233 (O_1233,N_45179,N_48808);
nand UO_1234 (O_1234,N_44782,N_41914);
nand UO_1235 (O_1235,N_41814,N_40689);
xor UO_1236 (O_1236,N_48395,N_49685);
or UO_1237 (O_1237,N_49548,N_47406);
nand UO_1238 (O_1238,N_49948,N_48728);
xnor UO_1239 (O_1239,N_45462,N_44720);
nor UO_1240 (O_1240,N_40624,N_48912);
or UO_1241 (O_1241,N_47904,N_47911);
or UO_1242 (O_1242,N_41692,N_42986);
nand UO_1243 (O_1243,N_49210,N_40632);
nand UO_1244 (O_1244,N_48484,N_48761);
xor UO_1245 (O_1245,N_49550,N_41769);
nor UO_1246 (O_1246,N_42384,N_47105);
and UO_1247 (O_1247,N_48708,N_45568);
or UO_1248 (O_1248,N_44488,N_42094);
nor UO_1249 (O_1249,N_49412,N_40635);
nor UO_1250 (O_1250,N_42606,N_41689);
nor UO_1251 (O_1251,N_48633,N_47506);
and UO_1252 (O_1252,N_40811,N_42540);
xor UO_1253 (O_1253,N_41675,N_48980);
nand UO_1254 (O_1254,N_43386,N_45227);
and UO_1255 (O_1255,N_47212,N_44566);
or UO_1256 (O_1256,N_43769,N_49285);
or UO_1257 (O_1257,N_47223,N_47940);
nor UO_1258 (O_1258,N_42689,N_49961);
nand UO_1259 (O_1259,N_46253,N_40357);
nand UO_1260 (O_1260,N_46083,N_47122);
xor UO_1261 (O_1261,N_40855,N_41386);
or UO_1262 (O_1262,N_40033,N_40053);
or UO_1263 (O_1263,N_41027,N_43023);
nand UO_1264 (O_1264,N_44565,N_45999);
or UO_1265 (O_1265,N_46541,N_47899);
or UO_1266 (O_1266,N_40881,N_45824);
xor UO_1267 (O_1267,N_43949,N_41854);
or UO_1268 (O_1268,N_45370,N_43297);
or UO_1269 (O_1269,N_49614,N_43821);
nand UO_1270 (O_1270,N_44100,N_44499);
nand UO_1271 (O_1271,N_45456,N_49101);
nand UO_1272 (O_1272,N_46926,N_42885);
or UO_1273 (O_1273,N_42942,N_41721);
or UO_1274 (O_1274,N_43376,N_40900);
or UO_1275 (O_1275,N_48621,N_44704);
nor UO_1276 (O_1276,N_40204,N_44840);
and UO_1277 (O_1277,N_41391,N_43305);
or UO_1278 (O_1278,N_41975,N_45150);
or UO_1279 (O_1279,N_42820,N_40783);
and UO_1280 (O_1280,N_40297,N_46481);
nor UO_1281 (O_1281,N_46212,N_49413);
nand UO_1282 (O_1282,N_47834,N_45941);
or UO_1283 (O_1283,N_47938,N_43981);
xor UO_1284 (O_1284,N_42149,N_42267);
or UO_1285 (O_1285,N_43429,N_45490);
and UO_1286 (O_1286,N_42903,N_43052);
nor UO_1287 (O_1287,N_49840,N_47767);
nor UO_1288 (O_1288,N_44319,N_41298);
xor UO_1289 (O_1289,N_46913,N_42191);
or UO_1290 (O_1290,N_41632,N_42113);
or UO_1291 (O_1291,N_48891,N_40528);
nor UO_1292 (O_1292,N_41249,N_41153);
or UO_1293 (O_1293,N_44170,N_43291);
or UO_1294 (O_1294,N_49199,N_44095);
or UO_1295 (O_1295,N_45637,N_45232);
nor UO_1296 (O_1296,N_48943,N_47650);
nand UO_1297 (O_1297,N_42876,N_46318);
or UO_1298 (O_1298,N_45851,N_40037);
nor UO_1299 (O_1299,N_42646,N_43767);
or UO_1300 (O_1300,N_48382,N_42895);
nor UO_1301 (O_1301,N_46579,N_45115);
and UO_1302 (O_1302,N_45344,N_41882);
xnor UO_1303 (O_1303,N_46530,N_49367);
and UO_1304 (O_1304,N_49830,N_44088);
nand UO_1305 (O_1305,N_49196,N_46847);
xnor UO_1306 (O_1306,N_40717,N_46289);
nand UO_1307 (O_1307,N_47297,N_42134);
or UO_1308 (O_1308,N_40918,N_47736);
and UO_1309 (O_1309,N_43924,N_44506);
nor UO_1310 (O_1310,N_46686,N_49309);
or UO_1311 (O_1311,N_44818,N_44473);
or UO_1312 (O_1312,N_48879,N_43965);
xor UO_1313 (O_1313,N_49800,N_41825);
and UO_1314 (O_1314,N_40979,N_40588);
nand UO_1315 (O_1315,N_47016,N_42497);
nand UO_1316 (O_1316,N_44276,N_42746);
and UO_1317 (O_1317,N_49402,N_48725);
or UO_1318 (O_1318,N_41254,N_42872);
and UO_1319 (O_1319,N_48709,N_42864);
nor UO_1320 (O_1320,N_46274,N_42234);
nor UO_1321 (O_1321,N_47207,N_41488);
or UO_1322 (O_1322,N_45551,N_43449);
nand UO_1323 (O_1323,N_49434,N_49683);
nand UO_1324 (O_1324,N_42586,N_48620);
and UO_1325 (O_1325,N_44939,N_45586);
nor UO_1326 (O_1326,N_42911,N_46347);
or UO_1327 (O_1327,N_41414,N_45054);
nor UO_1328 (O_1328,N_49776,N_40857);
xor UO_1329 (O_1329,N_40433,N_44836);
or UO_1330 (O_1330,N_47735,N_48226);
or UO_1331 (O_1331,N_42448,N_49086);
nor UO_1332 (O_1332,N_46775,N_41455);
and UO_1333 (O_1333,N_49475,N_48037);
or UO_1334 (O_1334,N_41732,N_49815);
nand UO_1335 (O_1335,N_43875,N_49938);
or UO_1336 (O_1336,N_47381,N_46562);
and UO_1337 (O_1337,N_47491,N_43362);
and UO_1338 (O_1338,N_49090,N_44520);
nand UO_1339 (O_1339,N_47610,N_42109);
or UO_1340 (O_1340,N_40743,N_40131);
nor UO_1341 (O_1341,N_49266,N_41104);
nand UO_1342 (O_1342,N_45091,N_44312);
nand UO_1343 (O_1343,N_48325,N_49865);
nor UO_1344 (O_1344,N_45783,N_43921);
nand UO_1345 (O_1345,N_49509,N_43175);
and UO_1346 (O_1346,N_48683,N_45405);
nor UO_1347 (O_1347,N_49868,N_40358);
and UO_1348 (O_1348,N_49883,N_40736);
xor UO_1349 (O_1349,N_49381,N_44597);
and UO_1350 (O_1350,N_41276,N_40164);
nor UO_1351 (O_1351,N_45300,N_46257);
and UO_1352 (O_1352,N_43895,N_45117);
or UO_1353 (O_1353,N_43024,N_42115);
nand UO_1354 (O_1354,N_44316,N_44124);
nand UO_1355 (O_1355,N_40638,N_40208);
nand UO_1356 (O_1356,N_48929,N_45834);
or UO_1357 (O_1357,N_48048,N_48941);
or UO_1358 (O_1358,N_43348,N_48230);
and UO_1359 (O_1359,N_49746,N_40038);
nand UO_1360 (O_1360,N_47963,N_43253);
nor UO_1361 (O_1361,N_48323,N_45236);
nand UO_1362 (O_1362,N_49095,N_49306);
nor UO_1363 (O_1363,N_43748,N_41091);
nand UO_1364 (O_1364,N_45285,N_45684);
nor UO_1365 (O_1365,N_48574,N_44911);
nor UO_1366 (O_1366,N_41980,N_49983);
and UO_1367 (O_1367,N_47626,N_46126);
nor UO_1368 (O_1368,N_47975,N_42411);
nand UO_1369 (O_1369,N_44371,N_42229);
nor UO_1370 (O_1370,N_41484,N_42293);
and UO_1371 (O_1371,N_48553,N_49384);
nor UO_1372 (O_1372,N_43350,N_40043);
and UO_1373 (O_1373,N_45937,N_47627);
nand UO_1374 (O_1374,N_49910,N_49820);
and UO_1375 (O_1375,N_49881,N_49360);
nor UO_1376 (O_1376,N_47805,N_43050);
or UO_1377 (O_1377,N_40698,N_49952);
nand UO_1378 (O_1378,N_46764,N_40659);
nor UO_1379 (O_1379,N_41773,N_46294);
or UO_1380 (O_1380,N_41890,N_44578);
nand UO_1381 (O_1381,N_41083,N_40800);
or UO_1382 (O_1382,N_42630,N_43384);
or UO_1383 (O_1383,N_48546,N_45485);
and UO_1384 (O_1384,N_40074,N_43925);
xnor UO_1385 (O_1385,N_47427,N_40856);
nor UO_1386 (O_1386,N_45172,N_42400);
or UO_1387 (O_1387,N_48935,N_40258);
nand UO_1388 (O_1388,N_43689,N_47339);
xor UO_1389 (O_1389,N_44503,N_46937);
and UO_1390 (O_1390,N_41392,N_46410);
nor UO_1391 (O_1391,N_48163,N_43725);
nor UO_1392 (O_1392,N_43552,N_41515);
nand UO_1393 (O_1393,N_46780,N_48470);
xnor UO_1394 (O_1394,N_40874,N_40568);
and UO_1395 (O_1395,N_48500,N_43019);
nand UO_1396 (O_1396,N_41469,N_46122);
nor UO_1397 (O_1397,N_40551,N_40279);
and UO_1398 (O_1398,N_48333,N_40864);
xnor UO_1399 (O_1399,N_44464,N_43967);
xnor UO_1400 (O_1400,N_48218,N_49519);
nor UO_1401 (O_1401,N_45438,N_49787);
or UO_1402 (O_1402,N_43128,N_47707);
nor UO_1403 (O_1403,N_45030,N_42059);
nand UO_1404 (O_1404,N_48123,N_40242);
and UO_1405 (O_1405,N_45772,N_42740);
nor UO_1406 (O_1406,N_43818,N_47354);
xnor UO_1407 (O_1407,N_46025,N_48880);
or UO_1408 (O_1408,N_43958,N_46172);
nor UO_1409 (O_1409,N_40976,N_42577);
or UO_1410 (O_1410,N_43792,N_44938);
xnor UO_1411 (O_1411,N_46062,N_45415);
nand UO_1412 (O_1412,N_48584,N_43063);
nand UO_1413 (O_1413,N_44143,N_47386);
xnor UO_1414 (O_1414,N_48836,N_45464);
or UO_1415 (O_1415,N_40580,N_41646);
or UO_1416 (O_1416,N_46337,N_45407);
nand UO_1417 (O_1417,N_49225,N_44094);
or UO_1418 (O_1418,N_44718,N_43092);
nand UO_1419 (O_1419,N_49949,N_44523);
or UO_1420 (O_1420,N_48702,N_44062);
nor UO_1421 (O_1421,N_48766,N_43067);
xor UO_1422 (O_1422,N_48271,N_45719);
nor UO_1423 (O_1423,N_41425,N_47892);
xor UO_1424 (O_1424,N_45292,N_49687);
and UO_1425 (O_1425,N_49684,N_47082);
nand UO_1426 (O_1426,N_41936,N_49942);
nor UO_1427 (O_1427,N_41871,N_44800);
or UO_1428 (O_1428,N_40246,N_48664);
and UO_1429 (O_1429,N_49263,N_43891);
nand UO_1430 (O_1430,N_44317,N_46777);
and UO_1431 (O_1431,N_47786,N_48350);
or UO_1432 (O_1432,N_44871,N_42205);
nand UO_1433 (O_1433,N_47530,N_42132);
nand UO_1434 (O_1434,N_45744,N_43508);
nor UO_1435 (O_1435,N_44144,N_41791);
nor UO_1436 (O_1436,N_49318,N_48265);
nand UO_1437 (O_1437,N_41673,N_42997);
and UO_1438 (O_1438,N_42429,N_49582);
or UO_1439 (O_1439,N_41476,N_45062);
nor UO_1440 (O_1440,N_49804,N_42424);
nand UO_1441 (O_1441,N_48840,N_47380);
or UO_1442 (O_1442,N_40572,N_41636);
xnor UO_1443 (O_1443,N_48744,N_48280);
xor UO_1444 (O_1444,N_40640,N_46108);
or UO_1445 (O_1445,N_49292,N_49445);
and UO_1446 (O_1446,N_41335,N_41007);
nor UO_1447 (O_1447,N_43167,N_49201);
or UO_1448 (O_1448,N_49400,N_43182);
xor UO_1449 (O_1449,N_44640,N_40661);
nor UO_1450 (O_1450,N_46278,N_43338);
nand UO_1451 (O_1451,N_41990,N_43443);
nor UO_1452 (O_1452,N_40241,N_48898);
and UO_1453 (O_1453,N_40390,N_40453);
nor UO_1454 (O_1454,N_49583,N_40431);
and UO_1455 (O_1455,N_45152,N_41420);
or UO_1456 (O_1456,N_41965,N_47935);
nand UO_1457 (O_1457,N_48415,N_41803);
nor UO_1458 (O_1458,N_43018,N_44997);
and UO_1459 (O_1459,N_40051,N_40948);
nand UO_1460 (O_1460,N_49237,N_45049);
nand UO_1461 (O_1461,N_46560,N_48238);
and UO_1462 (O_1462,N_48257,N_44655);
or UO_1463 (O_1463,N_45457,N_41545);
and UO_1464 (O_1464,N_44985,N_46708);
and UO_1465 (O_1465,N_41289,N_41520);
nor UO_1466 (O_1466,N_49027,N_47502);
and UO_1467 (O_1467,N_45784,N_48737);
nand UO_1468 (O_1468,N_49836,N_40884);
and UO_1469 (O_1469,N_44223,N_44600);
or UO_1470 (O_1470,N_47466,N_48249);
and UO_1471 (O_1471,N_46147,N_41844);
nor UO_1472 (O_1472,N_40662,N_42881);
nand UO_1473 (O_1473,N_48094,N_43905);
or UO_1474 (O_1474,N_47183,N_43939);
nand UO_1475 (O_1475,N_49579,N_44793);
nand UO_1476 (O_1476,N_40602,N_42608);
and UO_1477 (O_1477,N_42428,N_44612);
or UO_1478 (O_1478,N_49970,N_49756);
or UO_1479 (O_1479,N_48023,N_44627);
and UO_1480 (O_1480,N_45423,N_49779);
and UO_1481 (O_1481,N_48030,N_44903);
and UO_1482 (O_1482,N_44146,N_45650);
and UO_1483 (O_1483,N_43655,N_46846);
nor UO_1484 (O_1484,N_41979,N_44673);
xnor UO_1485 (O_1485,N_42648,N_43469);
or UO_1486 (O_1486,N_42146,N_43988);
and UO_1487 (O_1487,N_44093,N_43620);
and UO_1488 (O_1488,N_49083,N_41722);
and UO_1489 (O_1489,N_49321,N_48029);
nor UO_1490 (O_1490,N_48950,N_42481);
nor UO_1491 (O_1491,N_45905,N_42295);
and UO_1492 (O_1492,N_46138,N_40105);
and UO_1493 (O_1493,N_46712,N_45704);
nand UO_1494 (O_1494,N_49502,N_43047);
nor UO_1495 (O_1495,N_46845,N_43956);
or UO_1496 (O_1496,N_47097,N_40507);
or UO_1497 (O_1497,N_46399,N_48542);
nand UO_1498 (O_1498,N_44233,N_42292);
and UO_1499 (O_1499,N_40498,N_46950);
or UO_1500 (O_1500,N_42792,N_42417);
or UO_1501 (O_1501,N_45059,N_44695);
xor UO_1502 (O_1502,N_40801,N_46225);
and UO_1503 (O_1503,N_41833,N_42365);
or UO_1504 (O_1504,N_43684,N_43896);
and UO_1505 (O_1505,N_46403,N_42232);
xor UO_1506 (O_1506,N_45701,N_42518);
or UO_1507 (O_1507,N_40667,N_42774);
xor UO_1508 (O_1508,N_46072,N_43472);
and UO_1509 (O_1509,N_44790,N_41813);
or UO_1510 (O_1510,N_42574,N_43422);
nand UO_1511 (O_1511,N_45153,N_41046);
xnor UO_1512 (O_1512,N_47821,N_45479);
or UO_1513 (O_1513,N_47710,N_47056);
or UO_1514 (O_1514,N_42250,N_43784);
or UO_1515 (O_1515,N_49736,N_47836);
nor UO_1516 (O_1516,N_46503,N_44583);
and UO_1517 (O_1517,N_49757,N_45840);
nor UO_1518 (O_1518,N_48539,N_43749);
and UO_1519 (O_1519,N_43711,N_40041);
xnor UO_1520 (O_1520,N_47974,N_40079);
nand UO_1521 (O_1521,N_41013,N_48425);
or UO_1522 (O_1522,N_49932,N_46000);
nand UO_1523 (O_1523,N_43258,N_44348);
nor UO_1524 (O_1524,N_46722,N_49231);
and UO_1525 (O_1525,N_41378,N_49940);
or UO_1526 (O_1526,N_42345,N_48360);
or UO_1527 (O_1527,N_43475,N_41754);
nor UO_1528 (O_1528,N_40655,N_45795);
nand UO_1529 (O_1529,N_49531,N_44438);
nor UO_1530 (O_1530,N_48171,N_46011);
nor UO_1531 (O_1531,N_43755,N_46009);
and UO_1532 (O_1532,N_44353,N_45523);
nor UO_1533 (O_1533,N_47440,N_46703);
and UO_1534 (O_1534,N_41885,N_43619);
or UO_1535 (O_1535,N_49544,N_40383);
or UO_1536 (O_1536,N_43087,N_44163);
or UO_1537 (O_1537,N_49607,N_46107);
nor UO_1538 (O_1538,N_43156,N_40115);
nor UO_1539 (O_1539,N_41648,N_47480);
nor UO_1540 (O_1540,N_46302,N_48351);
nor UO_1541 (O_1541,N_40008,N_47708);
and UO_1542 (O_1542,N_49813,N_47550);
nand UO_1543 (O_1543,N_44775,N_41471);
or UO_1544 (O_1544,N_46633,N_42557);
nor UO_1545 (O_1545,N_45550,N_44491);
nand UO_1546 (O_1546,N_45822,N_47613);
or UO_1547 (O_1547,N_47645,N_48513);
or UO_1548 (O_1548,N_43521,N_48067);
nor UO_1549 (O_1549,N_45274,N_41628);
or UO_1550 (O_1550,N_45751,N_40444);
nor UO_1551 (O_1551,N_49279,N_41929);
xnor UO_1552 (O_1552,N_44012,N_46497);
nand UO_1553 (O_1553,N_41869,N_48482);
or UO_1554 (O_1554,N_44678,N_45758);
nand UO_1555 (O_1555,N_42865,N_49782);
nand UO_1556 (O_1556,N_49655,N_40816);
xor UO_1557 (O_1557,N_49108,N_41305);
nand UO_1558 (O_1558,N_43880,N_40833);
nor UO_1559 (O_1559,N_40319,N_49396);
nand UO_1560 (O_1560,N_49462,N_48069);
nor UO_1561 (O_1561,N_49567,N_48366);
nor UO_1562 (O_1562,N_42180,N_44888);
or UO_1563 (O_1563,N_43487,N_47167);
nor UO_1564 (O_1564,N_48579,N_47086);
or UO_1565 (O_1565,N_44336,N_43616);
and UO_1566 (O_1566,N_47065,N_42441);
and UO_1567 (O_1567,N_42568,N_49556);
nand UO_1568 (O_1568,N_49654,N_48662);
and UO_1569 (O_1569,N_41807,N_40248);
and UO_1570 (O_1570,N_44428,N_45536);
nor UO_1571 (O_1571,N_47800,N_45584);
nand UO_1572 (O_1572,N_47770,N_48053);
nand UO_1573 (O_1573,N_42697,N_45138);
nand UO_1574 (O_1574,N_49523,N_41793);
xnor UO_1575 (O_1575,N_41547,N_43736);
and UO_1576 (O_1576,N_46129,N_40212);
and UO_1577 (O_1577,N_41446,N_46326);
nand UO_1578 (O_1578,N_48937,N_43613);
nand UO_1579 (O_1579,N_43497,N_49597);
nor UO_1580 (O_1580,N_44639,N_43130);
and UO_1581 (O_1581,N_44585,N_41862);
or UO_1582 (O_1582,N_49963,N_42385);
xor UO_1583 (O_1583,N_40705,N_48700);
or UO_1584 (O_1584,N_45087,N_41696);
nand UO_1585 (O_1585,N_47206,N_44513);
or UO_1586 (O_1586,N_42866,N_44257);
nor UO_1587 (O_1587,N_44984,N_42170);
or UO_1588 (O_1588,N_48884,N_49723);
and UO_1589 (O_1589,N_49176,N_41614);
or UO_1590 (O_1590,N_48854,N_49966);
nor UO_1591 (O_1591,N_47231,N_47738);
and UO_1592 (O_1592,N_47343,N_40718);
and UO_1593 (O_1593,N_43434,N_48845);
nor UO_1594 (O_1594,N_40513,N_43400);
nand UO_1595 (O_1595,N_44758,N_41571);
or UO_1596 (O_1596,N_48225,N_40149);
nand UO_1597 (O_1597,N_46620,N_40552);
nand UO_1598 (O_1598,N_46675,N_41442);
or UO_1599 (O_1599,N_44153,N_43858);
and UO_1600 (O_1600,N_43706,N_41310);
nand UO_1601 (O_1601,N_43285,N_46159);
xor UO_1602 (O_1602,N_44166,N_46300);
and UO_1603 (O_1603,N_41423,N_43990);
nor UO_1604 (O_1604,N_47074,N_49527);
nand UO_1605 (O_1605,N_45532,N_46304);
and UO_1606 (O_1606,N_46759,N_40125);
and UO_1607 (O_1607,N_44698,N_41452);
xor UO_1608 (O_1608,N_45198,N_41680);
nand UO_1609 (O_1609,N_49643,N_43158);
or UO_1610 (O_1610,N_42671,N_44642);
nand UO_1611 (O_1611,N_49911,N_45419);
nand UO_1612 (O_1612,N_49539,N_46718);
xnor UO_1613 (O_1613,N_44474,N_49730);
nand UO_1614 (O_1614,N_42994,N_40778);
and UO_1615 (O_1615,N_46668,N_48442);
nand UO_1616 (O_1616,N_46707,N_49613);
nand UO_1617 (O_1617,N_42694,N_44901);
or UO_1618 (O_1618,N_43599,N_48042);
and UO_1619 (O_1619,N_46629,N_40135);
nand UO_1620 (O_1620,N_47347,N_41424);
and UO_1621 (O_1621,N_47902,N_40217);
and UO_1622 (O_1622,N_46714,N_44728);
nor UO_1623 (O_1623,N_46812,N_45291);
and UO_1624 (O_1624,N_44156,N_44839);
nand UO_1625 (O_1625,N_42515,N_40332);
nor UO_1626 (O_1626,N_49793,N_45875);
xnor UO_1627 (O_1627,N_40066,N_43734);
xor UO_1628 (O_1628,N_45496,N_40555);
nor UO_1629 (O_1629,N_42921,N_43417);
nor UO_1630 (O_1630,N_40817,N_43827);
nor UO_1631 (O_1631,N_49256,N_46501);
nand UO_1632 (O_1632,N_42256,N_40227);
nor UO_1633 (O_1633,N_42506,N_41230);
nor UO_1634 (O_1634,N_43532,N_43292);
and UO_1635 (O_1635,N_41158,N_47926);
nor UO_1636 (O_1636,N_42613,N_44381);
nand UO_1637 (O_1637,N_42117,N_40103);
or UO_1638 (O_1638,N_49586,N_49984);
xnor UO_1639 (O_1639,N_43793,N_45304);
nand UO_1640 (O_1640,N_49249,N_46057);
or UO_1641 (O_1641,N_40601,N_49438);
and UO_1642 (O_1642,N_46045,N_41641);
nor UO_1643 (O_1643,N_42960,N_48613);
and UO_1644 (O_1644,N_47516,N_47057);
or UO_1645 (O_1645,N_43745,N_41598);
and UO_1646 (O_1646,N_47379,N_44876);
and UO_1647 (O_1647,N_49149,N_42683);
or UO_1648 (O_1648,N_47547,N_49644);
and UO_1649 (O_1649,N_46974,N_41105);
nand UO_1650 (O_1650,N_41874,N_41321);
nand UO_1651 (O_1651,N_44729,N_41916);
or UO_1652 (O_1652,N_48933,N_40561);
or UO_1653 (O_1653,N_45043,N_47178);
or UO_1654 (O_1654,N_40210,N_44392);
nand UO_1655 (O_1655,N_41322,N_45297);
and UO_1656 (O_1656,N_47076,N_45781);
or UO_1657 (O_1657,N_42031,N_49572);
or UO_1658 (O_1658,N_48658,N_40166);
nand UO_1659 (O_1659,N_45149,N_44877);
nand UO_1660 (O_1660,N_49205,N_40607);
nor UO_1661 (O_1661,N_47741,N_47514);
xnor UO_1662 (O_1662,N_44201,N_45422);
and UO_1663 (O_1663,N_46380,N_44829);
and UO_1664 (O_1664,N_41665,N_48457);
nand UO_1665 (O_1665,N_49835,N_40585);
nor UO_1666 (O_1666,N_40516,N_44411);
or UO_1667 (O_1667,N_43423,N_42344);
and UO_1668 (O_1668,N_40165,N_43842);
and UO_1669 (O_1669,N_42139,N_44326);
or UO_1670 (O_1670,N_44379,N_49809);
nor UO_1671 (O_1671,N_41832,N_46586);
or UO_1672 (O_1672,N_47100,N_45477);
or UO_1673 (O_1673,N_49788,N_44460);
nand UO_1674 (O_1674,N_48571,N_42739);
and UO_1675 (O_1675,N_47141,N_48240);
nand UO_1676 (O_1676,N_42294,N_43247);
nor UO_1677 (O_1677,N_46179,N_47019);
xnor UO_1678 (O_1678,N_45416,N_46834);
or UO_1679 (O_1679,N_47040,N_41106);
nand UO_1680 (O_1680,N_49283,N_47357);
and UO_1681 (O_1681,N_43776,N_47748);
or UO_1682 (O_1682,N_49662,N_46061);
and UO_1683 (O_1683,N_41449,N_44267);
or UO_1684 (O_1684,N_42088,N_48384);
or UO_1685 (O_1685,N_41541,N_46479);
xnor UO_1686 (O_1686,N_49774,N_49073);
nand UO_1687 (O_1687,N_46746,N_43796);
or UO_1688 (O_1688,N_44750,N_43026);
xor UO_1689 (O_1689,N_46854,N_43645);
and UO_1690 (O_1690,N_47280,N_42183);
and UO_1691 (O_1691,N_45836,N_49933);
nand UO_1692 (O_1692,N_48837,N_42298);
and UO_1693 (O_1693,N_47069,N_44529);
and UO_1694 (O_1694,N_49380,N_43217);
or UO_1695 (O_1695,N_43707,N_43465);
or UO_1696 (O_1696,N_44056,N_49162);
nand UO_1697 (O_1697,N_45209,N_44164);
or UO_1698 (O_1698,N_46908,N_41630);
and UO_1699 (O_1699,N_43178,N_41563);
or UO_1700 (O_1700,N_43320,N_40333);
and UO_1701 (O_1701,N_42398,N_46276);
nor UO_1702 (O_1702,N_46022,N_40355);
nor UO_1703 (O_1703,N_40680,N_45581);
and UO_1704 (O_1704,N_42504,N_40627);
nor UO_1705 (O_1705,N_46438,N_40399);
xor UO_1706 (O_1706,N_49267,N_48121);
xor UO_1707 (O_1707,N_47113,N_46373);
nand UO_1708 (O_1708,N_49390,N_43271);
and UO_1709 (O_1709,N_42306,N_46117);
xnor UO_1710 (O_1710,N_48901,N_44649);
and UO_1711 (O_1711,N_40724,N_42736);
or UO_1712 (O_1712,N_45756,N_44919);
and UO_1713 (O_1713,N_48065,N_47531);
and UO_1714 (O_1714,N_48188,N_47161);
nand UO_1715 (O_1715,N_44986,N_41336);
and UO_1716 (O_1716,N_49755,N_44543);
and UO_1717 (O_1717,N_43718,N_40484);
or UO_1718 (O_1718,N_40685,N_42008);
and UO_1719 (O_1719,N_46800,N_42440);
and UO_1720 (O_1720,N_41334,N_44141);
or UO_1721 (O_1721,N_44958,N_42581);
or UO_1722 (O_1722,N_42393,N_40235);
and UO_1723 (O_1723,N_49248,N_44426);
and UO_1724 (O_1724,N_41581,N_42462);
nand UO_1725 (O_1725,N_42950,N_45000);
and UO_1726 (O_1726,N_49520,N_45016);
nor UO_1727 (O_1727,N_49592,N_47646);
and UO_1728 (O_1728,N_40641,N_44591);
nand UO_1729 (O_1729,N_48631,N_44389);
or UO_1730 (O_1730,N_48107,N_44841);
or UO_1731 (O_1731,N_42771,N_47832);
or UO_1732 (O_1732,N_44886,N_44452);
nor UO_1733 (O_1733,N_46428,N_46006);
xor UO_1734 (O_1734,N_44889,N_42974);
or UO_1735 (O_1735,N_47669,N_42721);
or UO_1736 (O_1736,N_43583,N_43072);
or UO_1737 (O_1737,N_42603,N_44148);
and UO_1738 (O_1738,N_41342,N_42968);
or UO_1739 (O_1739,N_45989,N_47942);
or UO_1740 (O_1740,N_46266,N_49719);
nand UO_1741 (O_1741,N_44949,N_43551);
and UO_1742 (O_1742,N_46802,N_47429);
nor UO_1743 (O_1743,N_45646,N_40678);
nor UO_1744 (O_1744,N_45324,N_43339);
nor UO_1745 (O_1745,N_47352,N_48883);
nand UO_1746 (O_1746,N_42857,N_44536);
nor UO_1747 (O_1747,N_45708,N_41419);
and UO_1748 (O_1748,N_41892,N_43229);
and UO_1749 (O_1749,N_41937,N_49215);
nor UO_1750 (O_1750,N_43530,N_48074);
nor UO_1751 (O_1751,N_47497,N_44111);
and UO_1752 (O_1752,N_43865,N_47067);
or UO_1753 (O_1753,N_44530,N_46870);
and UO_1754 (O_1754,N_47394,N_48406);
nor UO_1755 (O_1755,N_47382,N_42837);
or UO_1756 (O_1756,N_40162,N_42397);
xor UO_1757 (O_1757,N_40371,N_44007);
or UO_1758 (O_1758,N_45580,N_46729);
or UO_1759 (O_1759,N_44002,N_47061);
or UO_1760 (O_1760,N_48841,N_44001);
nor UO_1761 (O_1761,N_42509,N_48622);
and UO_1762 (O_1762,N_46349,N_49632);
nor UO_1763 (O_1763,N_45180,N_40111);
or UO_1764 (O_1764,N_42991,N_46982);
nand UO_1765 (O_1765,N_42716,N_45653);
nor UO_1766 (O_1766,N_47728,N_47715);
nand UO_1767 (O_1767,N_41328,N_44586);
xor UO_1768 (O_1768,N_47321,N_48646);
nand UO_1769 (O_1769,N_48316,N_41849);
or UO_1770 (O_1770,N_44264,N_46698);
nor UO_1771 (O_1771,N_41375,N_40988);
nor UO_1772 (O_1772,N_40879,N_47044);
nor UO_1773 (O_1773,N_47154,N_41986);
or UO_1774 (O_1774,N_41149,N_47533);
nor UO_1775 (O_1775,N_42844,N_44019);
or UO_1776 (O_1776,N_47239,N_44948);
nor UO_1777 (O_1777,N_43107,N_49628);
nand UO_1778 (O_1778,N_48612,N_42039);
or UO_1779 (O_1779,N_49859,N_40735);
nor UO_1780 (O_1780,N_42972,N_47792);
xor UO_1781 (O_1781,N_40942,N_43269);
nand UO_1782 (O_1782,N_44779,N_49659);
nor UO_1783 (O_1783,N_45552,N_40575);
nand UO_1784 (O_1784,N_48999,N_43144);
xnor UO_1785 (O_1785,N_44239,N_48396);
nand UO_1786 (O_1786,N_42845,N_46258);
nand UO_1787 (O_1787,N_47791,N_40384);
or UO_1788 (O_1788,N_49805,N_45835);
nor UO_1789 (O_1789,N_48590,N_44182);
nand UO_1790 (O_1790,N_41949,N_43518);
and UO_1791 (O_1791,N_48844,N_45858);
nor UO_1792 (O_1792,N_42975,N_42331);
nand UO_1793 (O_1793,N_46465,N_49491);
xor UO_1794 (O_1794,N_41470,N_46111);
or UO_1795 (O_1795,N_49934,N_44900);
or UO_1796 (O_1796,N_47103,N_41991);
or UO_1797 (O_1797,N_40146,N_40693);
nand UO_1798 (O_1798,N_42751,N_47794);
nand UO_1799 (O_1799,N_43315,N_48815);
nor UO_1800 (O_1800,N_49099,N_44622);
nor UO_1801 (O_1801,N_41536,N_44929);
nand UO_1802 (O_1802,N_43116,N_47461);
and UO_1803 (O_1803,N_40761,N_46092);
and UO_1804 (O_1804,N_45113,N_45093);
or UO_1805 (O_1805,N_45845,N_41761);
nand UO_1806 (O_1806,N_47859,N_46016);
and UO_1807 (O_1807,N_47017,N_46312);
xor UO_1808 (O_1808,N_48706,N_42561);
and UO_1809 (O_1809,N_41583,N_45877);
nor UO_1810 (O_1810,N_42681,N_41710);
nor UO_1811 (O_1811,N_42492,N_49444);
nand UO_1812 (O_1812,N_40716,N_47890);
or UO_1813 (O_1813,N_46681,N_44465);
or UO_1814 (O_1814,N_40468,N_40387);
and UO_1815 (O_1815,N_47967,N_44032);
nand UO_1816 (O_1816,N_42066,N_49960);
or UO_1817 (O_1817,N_45657,N_47305);
or UO_1818 (O_1818,N_42833,N_47108);
nor UO_1819 (O_1819,N_46969,N_46085);
nor UO_1820 (O_1820,N_45076,N_49411);
or UO_1821 (O_1821,N_41189,N_44721);
and UO_1822 (O_1822,N_43536,N_41565);
nand UO_1823 (O_1823,N_47615,N_43585);
and UO_1824 (O_1824,N_42422,N_49731);
xnor UO_1825 (O_1825,N_44270,N_49450);
and UO_1826 (O_1826,N_44331,N_43037);
nor UO_1827 (O_1827,N_40489,N_46483);
xnor UO_1828 (O_1828,N_43111,N_49867);
or UO_1829 (O_1829,N_48146,N_48003);
nand UO_1830 (O_1830,N_42004,N_43973);
nand UO_1831 (O_1831,N_46490,N_41799);
or UO_1832 (O_1832,N_42788,N_49875);
or UO_1833 (O_1833,N_47664,N_48951);
and UO_1834 (O_1834,N_48519,N_44738);
nand UO_1835 (O_1835,N_46537,N_43526);
nor UO_1836 (O_1836,N_48305,N_48635);
and UO_1837 (O_1837,N_44508,N_48472);
and UO_1838 (O_1838,N_46651,N_49155);
or UO_1839 (O_1839,N_40541,N_41717);
nor UO_1840 (O_1840,N_45614,N_41759);
nand UO_1841 (O_1841,N_49134,N_47734);
nor UO_1842 (O_1842,N_46405,N_48994);
nand UO_1843 (O_1843,N_47927,N_41359);
and UO_1844 (O_1844,N_41712,N_40303);
nand UO_1845 (O_1845,N_40628,N_46510);
nand UO_1846 (O_1846,N_48911,N_49688);
xor UO_1847 (O_1847,N_44863,N_43697);
xor UO_1848 (O_1848,N_46167,N_49230);
or UO_1849 (O_1849,N_47426,N_46924);
or UO_1850 (O_1850,N_47833,N_41828);
or UO_1851 (O_1851,N_46491,N_41663);
or UO_1852 (O_1852,N_40353,N_49914);
or UO_1853 (O_1853,N_43744,N_48159);
or UO_1854 (O_1854,N_40327,N_49216);
nand UO_1855 (O_1855,N_43577,N_46693);
and UO_1856 (O_1856,N_42243,N_46144);
or UO_1857 (O_1857,N_45543,N_42093);
and UO_1858 (O_1858,N_43883,N_43040);
and UO_1859 (O_1859,N_49968,N_43135);
nor UO_1860 (O_1860,N_44186,N_45448);
or UO_1861 (O_1861,N_40311,N_43823);
nand UO_1862 (O_1862,N_45272,N_47353);
and UO_1863 (O_1863,N_42620,N_48617);
nand UO_1864 (O_1864,N_46039,N_45243);
or UO_1865 (O_1865,N_42924,N_45161);
and UO_1866 (O_1866,N_46753,N_47642);
nand UO_1867 (O_1867,N_43588,N_42032);
nand UO_1868 (O_1868,N_46957,N_43765);
xnor UO_1869 (O_1869,N_48100,N_48455);
and UO_1870 (O_1870,N_42682,N_46532);
and UO_1871 (O_1871,N_40515,N_44342);
nor UO_1872 (O_1872,N_41099,N_47425);
nor UO_1873 (O_1873,N_48408,N_42685);
nand UO_1874 (O_1874,N_41724,N_45135);
or UO_1875 (O_1875,N_47160,N_48739);
nand UO_1876 (O_1876,N_46599,N_42848);
and UO_1877 (O_1877,N_44273,N_40672);
or UO_1878 (O_1878,N_49422,N_40947);
nor UO_1879 (O_1879,N_40589,N_42333);
nand UO_1880 (O_1880,N_41917,N_45927);
or UO_1881 (O_1881,N_44004,N_41396);
and UO_1882 (O_1882,N_42503,N_49721);
nand UO_1883 (O_1883,N_43955,N_44251);
nor UO_1884 (O_1884,N_40798,N_40966);
nor UO_1885 (O_1885,N_43919,N_46242);
and UO_1886 (O_1886,N_44498,N_46210);
nor UO_1887 (O_1887,N_46264,N_40347);
nor UO_1888 (O_1888,N_40738,N_49282);
or UO_1889 (O_1889,N_47417,N_43431);
and UO_1890 (O_1890,N_44861,N_49545);
nand UO_1891 (O_1891,N_40719,N_42486);
or UO_1892 (O_1892,N_49993,N_40302);
or UO_1893 (O_1893,N_42269,N_49886);
and UO_1894 (O_1894,N_48818,N_43200);
or UO_1895 (O_1895,N_41734,N_42687);
nor UO_1896 (O_1896,N_42917,N_44613);
nor UO_1897 (O_1897,N_44556,N_49955);
nor UO_1898 (O_1898,N_45971,N_40928);
xor UO_1899 (O_1899,N_40897,N_47266);
nor UO_1900 (O_1900,N_40140,N_43716);
and UO_1901 (O_1901,N_46398,N_41066);
and UO_1902 (O_1902,N_43977,N_42040);
nor UO_1903 (O_1903,N_49153,N_43566);
nor UO_1904 (O_1904,N_41213,N_46859);
nand UO_1905 (O_1905,N_48764,N_45514);
and UO_1906 (O_1906,N_45608,N_49119);
or UO_1907 (O_1907,N_42818,N_47698);
or UO_1908 (O_1908,N_42048,N_48743);
or UO_1909 (O_1909,N_45451,N_40007);
nand UO_1910 (O_1910,N_46691,N_40898);
xor UO_1911 (O_1911,N_47272,N_46706);
and UO_1912 (O_1912,N_46897,N_44851);
and UO_1913 (O_1913,N_46222,N_46474);
nand UO_1914 (O_1914,N_45705,N_40652);
nor UO_1915 (O_1915,N_44241,N_46909);
nor UO_1916 (O_1916,N_40510,N_47442);
and UO_1917 (O_1917,N_43120,N_45058);
or UO_1918 (O_1918,N_48103,N_42106);
nor UO_1919 (O_1919,N_47150,N_40120);
xnor UO_1920 (O_1920,N_48411,N_48695);
nor UO_1921 (O_1921,N_48987,N_40093);
and UO_1922 (O_1922,N_49499,N_41390);
and UO_1923 (O_1923,N_42498,N_47229);
and UO_1924 (O_1924,N_42143,N_47482);
nor UO_1925 (O_1925,N_43374,N_44593);
xor UO_1926 (O_1926,N_48405,N_45776);
and UO_1927 (O_1927,N_49979,N_41074);
and UO_1928 (O_1928,N_43070,N_49365);
or UO_1929 (O_1929,N_41272,N_45798);
or UO_1930 (O_1930,N_47397,N_48668);
nor UO_1931 (O_1931,N_42436,N_47943);
xor UO_1932 (O_1932,N_46335,N_47842);
and UO_1933 (O_1933,N_40457,N_41403);
or UO_1934 (O_1934,N_42198,N_41204);
and UO_1935 (O_1935,N_40917,N_41422);
or UO_1936 (O_1936,N_43779,N_44374);
nand UO_1937 (O_1937,N_44716,N_46362);
nand UO_1938 (O_1938,N_43592,N_42161);
nand UO_1939 (O_1939,N_42325,N_43227);
nand UO_1940 (O_1940,N_45886,N_41489);
and UO_1941 (O_1941,N_43427,N_45488);
nor UO_1942 (O_1942,N_46422,N_41954);
xor UO_1943 (O_1943,N_46649,N_43242);
and UO_1944 (O_1944,N_46640,N_49241);
nand UO_1945 (O_1945,N_47165,N_43071);
or UO_1946 (O_1946,N_49368,N_42753);
and UO_1947 (O_1947,N_44375,N_46455);
nor UO_1948 (O_1948,N_43311,N_47601);
nor UO_1949 (O_1949,N_47487,N_47092);
nand UO_1950 (O_1950,N_43208,N_41811);
or UO_1951 (O_1951,N_41374,N_46338);
nor UO_1952 (O_1952,N_40463,N_47171);
nor UO_1953 (O_1953,N_44914,N_48049);
nor UO_1954 (O_1954,N_43758,N_48516);
or UO_1955 (O_1955,N_42159,N_40861);
nand UO_1956 (O_1956,N_42386,N_45820);
and UO_1957 (O_1957,N_44954,N_42584);
xnor UO_1958 (O_1958,N_48227,N_45808);
or UO_1959 (O_1959,N_47773,N_41495);
nand UO_1960 (O_1960,N_42056,N_45132);
xor UO_1961 (O_1961,N_41280,N_46343);
nand UO_1962 (O_1962,N_46439,N_40101);
or UO_1963 (O_1963,N_42610,N_41634);
or UO_1964 (O_1964,N_45869,N_44489);
and UO_1965 (O_1965,N_45904,N_45461);
and UO_1966 (O_1966,N_47962,N_49116);
xor UO_1967 (O_1967,N_42082,N_47921);
and UO_1968 (O_1968,N_48445,N_46526);
xnor UO_1969 (O_1969,N_40378,N_48715);
xnor UO_1970 (O_1970,N_45052,N_44668);
and UO_1971 (O_1971,N_49677,N_44053);
or UO_1972 (O_1972,N_47079,N_40933);
nand UO_1973 (O_1973,N_43205,N_45266);
or UO_1974 (O_1974,N_45328,N_46645);
nor UO_1975 (O_1975,N_45361,N_44013);
and UO_1976 (O_1976,N_46922,N_43160);
nor UO_1977 (O_1977,N_43809,N_47861);
or UO_1978 (O_1978,N_45916,N_43687);
and UO_1979 (O_1979,N_47714,N_47446);
xor UO_1980 (O_1980,N_41226,N_44279);
nor UO_1981 (O_1981,N_46090,N_44633);
xor UO_1982 (O_1982,N_46161,N_42536);
nor UO_1983 (O_1983,N_41126,N_42989);
xor UO_1984 (O_1984,N_48092,N_44850);
or UO_1985 (O_1985,N_45569,N_45404);
and UO_1986 (O_1986,N_40727,N_46272);
or UO_1987 (O_1987,N_43290,N_42813);
and UO_1988 (O_1988,N_43899,N_40076);
or UO_1989 (O_1989,N_47841,N_41526);
or UO_1990 (O_1990,N_46102,N_49338);
nor UO_1991 (O_1991,N_44500,N_47258);
or UO_1992 (O_1992,N_44185,N_47116);
or UO_1993 (O_1993,N_47433,N_46762);
xnor UO_1994 (O_1994,N_49314,N_42055);
nor UO_1995 (O_1995,N_45880,N_45037);
nor UO_1996 (O_1996,N_48655,N_45964);
or UO_1997 (O_1997,N_48514,N_46206);
nor UO_1998 (O_1998,N_49152,N_41875);
nor UO_1999 (O_1999,N_42710,N_46880);
or UO_2000 (O_2000,N_49081,N_44663);
and UO_2001 (O_2001,N_48550,N_47671);
nor UO_2002 (O_2002,N_43882,N_44207);
xor UO_2003 (O_2003,N_46832,N_49167);
nand UO_2004 (O_2004,N_45109,N_41437);
or UO_2005 (O_2005,N_42930,N_46099);
nor UO_2006 (O_2006,N_48785,N_40720);
xor UO_2007 (O_2007,N_46395,N_47584);
or UO_2008 (O_2008,N_41377,N_46350);
nor UO_2009 (O_2009,N_40796,N_41757);
nand UO_2010 (O_2010,N_42578,N_43710);
xor UO_2011 (O_2011,N_47055,N_44892);
nor UO_2012 (O_2012,N_44924,N_40985);
nor UO_2013 (O_2013,N_48608,N_45271);
nor UO_2014 (O_2014,N_43640,N_49437);
nand UO_2015 (O_2015,N_42414,N_43238);
nor UO_2016 (O_2016,N_45240,N_45167);
and UO_2017 (O_2017,N_44842,N_40233);
nor UO_2018 (O_2018,N_46740,N_47949);
nand UO_2019 (O_2019,N_42628,N_44959);
xnor UO_2020 (O_2020,N_44054,N_46137);
nor UO_2021 (O_2021,N_47145,N_48215);
or UO_2022 (O_2022,N_42607,N_40922);
xnor UO_2023 (O_2023,N_47325,N_40083);
xor UO_2024 (O_2024,N_42458,N_48021);
xnor UO_2025 (O_2025,N_43436,N_42718);
nand UO_2026 (O_2026,N_48867,N_48449);
or UO_2027 (O_2027,N_47839,N_40626);
nor UO_2028 (O_2028,N_48413,N_46697);
and UO_2029 (O_2029,N_44305,N_49565);
or UO_2030 (O_2030,N_43540,N_40117);
nand UO_2031 (O_2031,N_48125,N_45424);
or UO_2032 (O_2032,N_41450,N_48673);
and UO_2033 (O_2033,N_48705,N_48060);
or UO_2034 (O_2034,N_47274,N_40389);
nor UO_2035 (O_2035,N_48558,N_43119);
nor UO_2036 (O_2036,N_48435,N_40883);
xnor UO_2037 (O_2037,N_43302,N_45946);
nand UO_2038 (O_2038,N_49097,N_49324);
nand UO_2039 (O_2039,N_40407,N_40449);
nand UO_2040 (O_2040,N_42945,N_47186);
and UO_2041 (O_2041,N_48830,N_41454);
nand UO_2042 (O_2042,N_45224,N_48354);
nand UO_2043 (O_2043,N_43467,N_45541);
nor UO_2044 (O_2044,N_41198,N_42263);
nand UO_2045 (O_2045,N_44303,N_43682);
or UO_2046 (O_2046,N_41538,N_44814);
or UO_2047 (O_2047,N_48906,N_42164);
xnor UO_2048 (O_2048,N_40010,N_42217);
nand UO_2049 (O_2049,N_47399,N_46394);
xnor UO_2050 (O_2050,N_47739,N_47685);
or UO_2051 (O_2051,N_43593,N_49446);
nand UO_2052 (O_2052,N_49823,N_49295);
nand UO_2053 (O_2053,N_46381,N_47689);
and UO_2054 (O_2054,N_41398,N_42748);
and UO_2055 (O_2055,N_49854,N_48345);
or UO_2056 (O_2056,N_43960,N_44653);
nand UO_2057 (O_2057,N_46952,N_40495);
or UO_2058 (O_2058,N_48565,N_49503);
nor UO_2059 (O_2059,N_48362,N_45166);
xor UO_2060 (O_2060,N_41848,N_48153);
nor UO_2061 (O_2061,N_47693,N_41745);
or UO_2062 (O_2062,N_46287,N_44132);
nor UO_2063 (O_2063,N_49515,N_45396);
or UO_2064 (O_2064,N_40058,N_42045);
nand UO_2065 (O_2065,N_48970,N_42215);
nor UO_2066 (O_2066,N_47823,N_46734);
and UO_2067 (O_2067,N_44972,N_46431);
xor UO_2068 (O_2068,N_49711,N_49132);
or UO_2069 (O_2069,N_45906,N_40476);
nor UO_2070 (O_2070,N_43847,N_40113);
or UO_2071 (O_2071,N_46890,N_43255);
xor UO_2072 (O_2072,N_41141,N_42104);
nand UO_2073 (O_2073,N_41968,N_46413);
or UO_2074 (O_2074,N_47910,N_42514);
and UO_2075 (O_2075,N_49460,N_47181);
nand UO_2076 (O_2076,N_44436,N_42796);
nand UO_2077 (O_2077,N_49164,N_46237);
nand UO_2078 (O_2078,N_47439,N_45197);
or UO_2079 (O_2079,N_40707,N_44969);
and UO_2080 (O_2080,N_42253,N_49036);
or UO_2081 (O_2081,N_49257,N_49229);
nor UO_2082 (O_2082,N_41109,N_41963);
or UO_2083 (O_2083,N_40312,N_45185);
nand UO_2084 (O_2084,N_43027,N_43554);
or UO_2085 (O_2085,N_47005,N_44564);
and UO_2086 (O_2086,N_47096,N_42644);
nand UO_2087 (O_2087,N_44610,N_48264);
or UO_2088 (O_2088,N_46970,N_46217);
or UO_2089 (O_2089,N_47112,N_47778);
nor UO_2090 (O_2090,N_42479,N_43598);
or UO_2091 (O_2091,N_42251,N_48931);
xor UO_2092 (O_2092,N_45363,N_47798);
nor UO_2093 (O_2093,N_42254,N_45694);
or UO_2094 (O_2094,N_48561,N_44272);
or UO_2095 (O_2095,N_41731,N_45288);
nor UO_2096 (O_2096,N_45712,N_42097);
nor UO_2097 (O_2097,N_45833,N_41140);
or UO_2098 (O_2098,N_45463,N_42005);
nor UO_2099 (O_2099,N_45377,N_49157);
nand UO_2100 (O_2100,N_42461,N_49307);
and UO_2101 (O_2101,N_47508,N_47270);
nand UO_2102 (O_2102,N_48893,N_43042);
and UO_2103 (O_2103,N_49751,N_48921);
and UO_2104 (O_2104,N_46248,N_45486);
and UO_2105 (O_2105,N_45023,N_44073);
nor UO_2106 (O_2106,N_48851,N_45726);
and UO_2107 (O_2107,N_44538,N_45600);
nand UO_2108 (O_2108,N_47807,N_43284);
and UO_2109 (O_2109,N_49244,N_40696);
xnor UO_2110 (O_2110,N_49016,N_42810);
nand UO_2111 (O_2111,N_45883,N_48108);
and UO_2112 (O_2112,N_44442,N_45321);
nand UO_2113 (O_2113,N_47396,N_48597);
and UO_2114 (O_2114,N_46521,N_46900);
nand UO_2115 (O_2115,N_42402,N_45178);
and UO_2116 (O_2116,N_49784,N_49745);
or UO_2117 (O_2117,N_46324,N_47609);
and UO_2118 (O_2118,N_48380,N_47143);
and UO_2119 (O_2119,N_48926,N_40831);
nor UO_2120 (O_2120,N_41217,N_47605);
or UO_2121 (O_2121,N_46259,N_49666);
or UO_2122 (O_2122,N_43907,N_40237);
nand UO_2123 (O_2123,N_49143,N_46059);
nand UO_2124 (O_2124,N_44596,N_40448);
nor UO_2125 (O_2125,N_42083,N_47444);
nor UO_2126 (O_2126,N_41798,N_42070);
nand UO_2127 (O_2127,N_45910,N_45014);
and UO_2128 (O_2128,N_41405,N_48852);
nor UO_2129 (O_2129,N_48860,N_49505);
and UO_2130 (O_2130,N_43358,N_49832);
or UO_2131 (O_2131,N_45669,N_41251);
xnor UO_2132 (O_2132,N_48802,N_43665);
and UO_2133 (O_2133,N_42372,N_42199);
nand UO_2134 (O_2134,N_44286,N_48206);
and UO_2135 (O_2135,N_46531,N_44501);
or UO_2136 (O_2136,N_40959,N_46351);
or UO_2137 (O_2137,N_40779,N_48161);
nor UO_2138 (O_2138,N_48549,N_47526);
or UO_2139 (O_2139,N_48557,N_44376);
nor UO_2140 (O_2140,N_40342,N_40502);
xor UO_2141 (O_2141,N_43677,N_49950);
xnor UO_2142 (O_2142,N_41092,N_49172);
nor UO_2143 (O_2143,N_42915,N_45747);
nor UO_2144 (O_2144,N_43946,N_49233);
xor UO_2145 (O_2145,N_47370,N_45163);
nand UO_2146 (O_2146,N_42773,N_40906);
nor UO_2147 (O_2147,N_43204,N_46369);
or UO_2148 (O_2148,N_46634,N_46190);
nand UO_2149 (O_2149,N_42582,N_46364);
and UO_2150 (O_2150,N_42918,N_44973);
nor UO_2151 (O_2151,N_41343,N_40570);
xor UO_2152 (O_2152,N_45162,N_47699);
nor UO_2153 (O_2153,N_49735,N_42627);
nand UO_2154 (O_2154,N_46411,N_49898);
and UO_2155 (O_2155,N_47022,N_48126);
nand UO_2156 (O_2156,N_49902,N_44160);
nand UO_2157 (O_2157,N_44440,N_44856);
nor UO_2158 (O_2158,N_48149,N_44117);
nor UO_2159 (O_2159,N_48155,N_41567);
and UO_2160 (O_2160,N_43470,N_47880);
nand UO_2161 (O_2161,N_49084,N_48253);
nor UO_2162 (O_2162,N_46938,N_41097);
nor UO_2163 (O_2163,N_40065,N_42173);
and UO_2164 (O_2164,N_43009,N_40317);
or UO_2165 (O_2165,N_44723,N_42760);
xnor UO_2166 (O_2166,N_41385,N_42660);
or UO_2167 (O_2167,N_44005,N_44893);
nor UO_2168 (O_2168,N_43314,N_43342);
and UO_2169 (O_2169,N_44685,N_47289);
and UO_2170 (O_2170,N_46444,N_47895);
or UO_2171 (O_2171,N_44964,N_48275);
xnor UO_2172 (O_2172,N_41222,N_40591);
nand UO_2173 (O_2173,N_48269,N_41599);
or UO_2174 (O_2174,N_46480,N_47717);
xnor UO_2175 (O_2175,N_40565,N_41555);
or UO_2176 (O_2176,N_45521,N_48762);
nor UO_2177 (O_2177,N_46131,N_45689);
nand UO_2178 (O_2178,N_49694,N_45743);
or UO_2179 (O_2179,N_45570,N_42652);
nand UO_2180 (O_2180,N_43048,N_46120);
and UO_2181 (O_2181,N_45024,N_41133);
and UO_2182 (O_2182,N_45690,N_41539);
xor UO_2183 (O_2183,N_49876,N_48292);
nand UO_2184 (O_2184,N_40849,N_40810);
or UO_2185 (O_2185,N_43020,N_41788);
and UO_2186 (O_2186,N_44136,N_40354);
xnor UO_2187 (O_2187,N_46709,N_40402);
or UO_2188 (O_2188,N_42604,N_44082);
nor UO_2189 (O_2189,N_41143,N_42322);
nand UO_2190 (O_2190,N_40187,N_45100);
xnor UO_2191 (O_2191,N_41664,N_43862);
and UO_2192 (O_2192,N_46143,N_40604);
nand UO_2193 (O_2193,N_48033,N_40244);
and UO_2194 (O_2194,N_48041,N_43550);
nor UO_2195 (O_2195,N_40764,N_46820);
nor UO_2196 (O_2196,N_43647,N_45476);
or UO_2197 (O_2197,N_43861,N_42334);
nor UO_2198 (O_2198,N_46678,N_44921);
nand UO_2199 (O_2199,N_40822,N_42825);
nor UO_2200 (O_2200,N_40445,N_45282);
nor UO_2201 (O_2201,N_45216,N_41051);
and UO_2202 (O_2202,N_44815,N_43693);
or UO_2203 (O_2203,N_41202,N_46566);
or UO_2204 (O_2204,N_49224,N_46040);
nor UO_2205 (O_2205,N_49964,N_44774);
nand UO_2206 (O_2206,N_45800,N_48132);
nor UO_2207 (O_2207,N_45876,N_44907);
or UO_2208 (O_2208,N_40280,N_42374);
nand UO_2209 (O_2209,N_46170,N_42904);
or UO_2210 (O_2210,N_48601,N_46663);
and UO_2211 (O_2211,N_48204,N_48657);
xor UO_2212 (O_2212,N_44989,N_45435);
or UO_2213 (O_2213,N_40189,N_43257);
nor UO_2214 (O_2214,N_42277,N_49098);
or UO_2215 (O_2215,N_43517,N_46316);
xor UO_2216 (O_2216,N_48945,N_47947);
and UO_2217 (O_2217,N_46799,N_43797);
xnor UO_2218 (O_2218,N_46077,N_41903);
nor UO_2219 (O_2219,N_46871,N_45930);
and UO_2220 (O_2220,N_47976,N_41285);
or UO_2221 (O_2221,N_47375,N_48385);
nand UO_2222 (O_2222,N_47569,N_42901);
or UO_2223 (O_2223,N_42663,N_48525);
nand UO_2224 (O_2224,N_42507,N_40617);
nand UO_2225 (O_2225,N_41764,N_49879);
nor UO_2226 (O_2226,N_48254,N_40328);
nor UO_2227 (O_2227,N_48684,N_49495);
nor UO_2228 (O_2228,N_40412,N_48139);
and UO_2229 (O_2229,N_40584,N_41163);
nand UO_2230 (O_2230,N_47572,N_42303);
nor UO_2231 (O_2231,N_42934,N_48710);
or UO_2232 (O_2232,N_42733,N_41180);
and UO_2233 (O_2233,N_46008,N_42761);
xor UO_2234 (O_2234,N_40576,N_40634);
and UO_2235 (O_2235,N_45809,N_49388);
nand UO_2236 (O_2236,N_41088,N_48653);
nand UO_2237 (O_2237,N_49897,N_48393);
or UO_2238 (O_2238,N_47345,N_43043);
or UO_2239 (O_2239,N_41231,N_43104);
and UO_2240 (O_2240,N_44161,N_46153);
xnor UO_2241 (O_2241,N_40421,N_46168);
xor UO_2242 (O_2242,N_42749,N_43454);
and UO_2243 (O_2243,N_48359,N_44681);
or UO_2244 (O_2244,N_49080,N_45792);
nand UO_2245 (O_2245,N_40067,N_44425);
nand UO_2246 (O_2246,N_45034,N_41542);
nand UO_2247 (O_2247,N_45433,N_44855);
xnor UO_2248 (O_2248,N_42769,N_42050);
or UO_2249 (O_2249,N_45088,N_48786);
and UO_2250 (O_2250,N_48736,N_44121);
nand UO_2251 (O_2251,N_43702,N_45740);
nor UO_2252 (O_2252,N_43014,N_42370);
nand UO_2253 (O_2253,N_45730,N_48800);
or UO_2254 (O_2254,N_49763,N_46700);
and UO_2255 (O_2255,N_45314,N_48475);
nor UO_2256 (O_2256,N_48112,N_47344);
xnor UO_2257 (O_2257,N_42313,N_49448);
and UO_2258 (O_2258,N_43855,N_46496);
and UO_2259 (O_2259,N_42559,N_48104);
xor UO_2260 (O_2260,N_44976,N_42925);
nor UO_2261 (O_2261,N_46319,N_41409);
nor UO_2262 (O_2262,N_46115,N_43267);
and UO_2263 (O_2263,N_42512,N_45460);
nor UO_2264 (O_2264,N_43329,N_41323);
nand UO_2265 (O_2265,N_44894,N_44310);
xnor UO_2266 (O_2266,N_49473,N_47700);
nor UO_2267 (O_2267,N_48913,N_46551);
or UO_2268 (O_2268,N_43873,N_41473);
or UO_2269 (O_2269,N_42783,N_47287);
and UO_2270 (O_2270,N_46404,N_48522);
or UO_2271 (O_2271,N_46434,N_45865);
or UO_2272 (O_2272,N_49759,N_48572);
xnor UO_2273 (O_2273,N_49401,N_49817);
or UO_2274 (O_2274,N_45123,N_40321);
nand UO_2275 (O_2275,N_40935,N_45985);
or UO_2276 (O_2276,N_40299,N_41809);
or UO_2277 (O_2277,N_48297,N_41948);
and UO_2278 (O_2278,N_49194,N_40334);
nor UO_2279 (O_2279,N_49496,N_41164);
nor UO_2280 (O_2280,N_43246,N_40082);
nand UO_2281 (O_2281,N_49533,N_48010);
or UO_2282 (O_2282,N_40134,N_44955);
nor UO_2283 (O_2283,N_41770,N_40153);
or UO_2284 (O_2284,N_49050,N_48000);
or UO_2285 (O_2285,N_46176,N_40666);
nand UO_2286 (O_2286,N_41924,N_43473);
or UO_2287 (O_2287,N_41616,N_46744);
xnor UO_2288 (O_2288,N_46299,N_42937);
or UO_2289 (O_2289,N_40854,N_42378);
and UO_2290 (O_2290,N_44628,N_45709);
and UO_2291 (O_2291,N_42340,N_45642);
and UO_2292 (O_2292,N_40145,N_43994);
xnor UO_2293 (O_2293,N_44490,N_44920);
or UO_2294 (O_2294,N_48857,N_45431);
or UO_2295 (O_2295,N_47262,N_49315);
nand UO_2296 (O_2296,N_41893,N_43399);
or UO_2297 (O_2297,N_42797,N_44834);
nor UO_2298 (O_2298,N_46288,N_43900);
nand UO_2299 (O_2299,N_49924,N_45371);
xnor UO_2300 (O_2300,N_45286,N_49785);
and UO_2301 (O_2301,N_48329,N_49329);
nor UO_2302 (O_2302,N_46796,N_43560);
and UO_2303 (O_2303,N_47803,N_48239);
or UO_2304 (O_2304,N_41107,N_47745);
or UO_2305 (O_2305,N_44159,N_46539);
and UO_2306 (O_2306,N_45319,N_45958);
nor UO_2307 (O_2307,N_41154,N_49403);
nand UO_2308 (O_2308,N_48864,N_42181);
and UO_2309 (O_2309,N_47449,N_47608);
and UO_2310 (O_2310,N_45583,N_41758);
nand UO_2311 (O_2311,N_44339,N_46285);
or UO_2312 (O_2312,N_44314,N_45628);
nor UO_2313 (O_2313,N_46265,N_49208);
nand UO_2314 (O_2314,N_40132,N_47036);
nand UO_2315 (O_2315,N_49920,N_46282);
and UO_2316 (O_2316,N_48178,N_43857);
nand UO_2317 (O_2317,N_42116,N_49470);
or UO_2318 (O_2318,N_48955,N_43259);
nor UO_2319 (O_2319,N_43413,N_46768);
nand UO_2320 (O_2320,N_46255,N_43492);
nor UO_2321 (O_2321,N_44444,N_46843);
or UO_2322 (O_2322,N_44797,N_45807);
or UO_2323 (O_2323,N_42670,N_46166);
or UO_2324 (O_2324,N_40276,N_48458);
xor UO_2325 (O_2325,N_49294,N_47709);
or UO_2326 (O_2326,N_48343,N_40806);
nor UO_2327 (O_2327,N_46475,N_48045);
nand UO_2328 (O_2328,N_48568,N_42530);
nand UO_2329 (O_2329,N_46701,N_45549);
xnor UO_2330 (O_2330,N_44192,N_43657);
nor UO_2331 (O_2331,N_44454,N_45997);
nand UO_2332 (O_2332,N_41129,N_46575);
nand UO_2333 (O_2333,N_44281,N_44135);
nand UO_2334 (O_2334,N_42352,N_49169);
or UO_2335 (O_2335,N_46605,N_49341);
nand UO_2336 (O_2336,N_42444,N_43196);
nand UO_2337 (O_2337,N_42709,N_47575);
nand UO_2338 (O_2338,N_42830,N_47681);
nor UO_2339 (O_2339,N_49339,N_45108);
and UO_2340 (O_2340,N_49962,N_49004);
nand UO_2341 (O_2341,N_44328,N_46769);
nor UO_2342 (O_2342,N_42936,N_49150);
nor UO_2343 (O_2343,N_45357,N_42430);
nor UO_2344 (O_2344,N_44104,N_41463);
or UO_2345 (O_2345,N_48278,N_46445);
or UO_2346 (O_2346,N_45934,N_41235);
xnor UO_2347 (O_2347,N_44978,N_42500);
nand UO_2348 (O_2348,N_40325,N_40232);
and UO_2349 (O_2349,N_46763,N_44373);
and UO_2350 (O_2350,N_49362,N_42916);
nand UO_2351 (O_2351,N_40427,N_48770);
xnor UO_2352 (O_2352,N_48799,N_40616);
nand UO_2353 (O_2353,N_47196,N_42022);
nand UO_2354 (O_2354,N_42956,N_40365);
nor UO_2355 (O_2355,N_40127,N_44831);
nor UO_2356 (O_2356,N_49079,N_40927);
nand UO_2357 (O_2357,N_47663,N_49486);
or UO_2358 (O_2358,N_44528,N_43638);
xnor UO_2359 (O_2359,N_47917,N_47612);
nor UO_2360 (O_2360,N_43652,N_45873);
or UO_2361 (O_2361,N_40611,N_40337);
or UO_2362 (O_2362,N_45222,N_40290);
nand UO_2363 (O_2363,N_46402,N_43280);
and UO_2364 (O_2364,N_48295,N_43392);
xor UO_2365 (O_2365,N_48184,N_45017);
or UO_2366 (O_2366,N_40702,N_47106);
nand UO_2367 (O_2367,N_49590,N_46214);
nand UO_2368 (O_2368,N_46791,N_48734);
nand UO_2369 (O_2369,N_44183,N_48220);
xor UO_2370 (O_2370,N_44670,N_40840);
and UO_2371 (O_2371,N_47259,N_45893);
or UO_2372 (O_2372,N_40138,N_47509);
nor UO_2373 (O_2373,N_40980,N_41584);
or UO_2374 (O_2374,N_40978,N_43288);
nand UO_2375 (O_2375,N_49717,N_48476);
or UO_2376 (O_2376,N_43312,N_44557);
or UO_2377 (O_2377,N_40759,N_48172);
nand UO_2378 (O_2378,N_49243,N_46031);
nand UO_2379 (O_2379,N_49186,N_45473);
nand UO_2380 (O_2380,N_40142,N_42434);
and UO_2381 (O_2381,N_49293,N_47003);
or UO_2382 (O_2382,N_43743,N_47228);
nand UO_2383 (O_2383,N_42549,N_43775);
or UO_2384 (O_2384,N_45918,N_46150);
and UO_2385 (O_2385,N_44764,N_40958);
and UO_2386 (O_2386,N_49944,N_43241);
and UO_2387 (O_2387,N_43803,N_42611);
nand UO_2388 (O_2388,N_41843,N_49006);
nand UO_2389 (O_2389,N_47930,N_44298);
and UO_2390 (O_2390,N_44269,N_49806);
nor UO_2391 (O_2391,N_45716,N_43966);
or UO_2392 (O_2392,N_46355,N_47986);
nand UO_2393 (O_2393,N_49408,N_40436);
xor UO_2394 (O_2394,N_49146,N_44590);
nand UO_2395 (O_2395,N_41523,N_45814);
nor UO_2396 (O_2396,N_44909,N_49562);
and UO_2397 (O_2397,N_41695,N_41699);
or UO_2398 (O_2398,N_46386,N_41010);
or UO_2399 (O_2399,N_45280,N_44879);
nor UO_2400 (O_2400,N_40768,N_42735);
xnor UO_2401 (O_2401,N_43123,N_49423);
xnor UO_2402 (O_2402,N_44680,N_49013);
nand UO_2403 (O_2403,N_43751,N_49093);
nor UO_2404 (O_2404,N_47551,N_45805);
nand UO_2405 (O_2405,N_42356,N_40954);
or UO_2406 (O_2406,N_41400,N_48962);
xor UO_2407 (O_2407,N_45399,N_41497);
and UO_2408 (O_2408,N_48355,N_41867);
nor UO_2409 (O_2409,N_46959,N_48438);
nor UO_2410 (O_2410,N_40004,N_43495);
or UO_2411 (O_2411,N_48217,N_43623);
or UO_2412 (O_2412,N_48486,N_44482);
nor UO_2413 (O_2413,N_47602,N_45126);
and UO_2414 (O_2414,N_46749,N_40080);
or UO_2415 (O_2415,N_48070,N_40923);
nand UO_2416 (O_2416,N_49011,N_40962);
nor UO_2417 (O_2417,N_45338,N_48623);
nand UO_2418 (O_2418,N_44816,N_46418);
nor UO_2419 (O_2419,N_44351,N_40430);
nor UO_2420 (O_2420,N_49232,N_44049);
or UO_2421 (O_2421,N_40372,N_46096);
nor UO_2422 (O_2422,N_46635,N_41282);
and UO_2423 (O_2423,N_49331,N_40749);
nand UO_2424 (O_2424,N_43727,N_41723);
xor UO_2425 (O_2425,N_48718,N_41774);
xnor UO_2426 (O_2426,N_46652,N_42756);
and UO_2427 (O_2427,N_42457,N_45780);
nor UO_2428 (O_2428,N_41368,N_40379);
xnor UO_2429 (O_2429,N_48179,N_44532);
or UO_2430 (O_2430,N_47292,N_47542);
or UO_2431 (O_2431,N_45454,N_40249);
and UO_2432 (O_2432,N_44362,N_44614);
xor UO_2433 (O_2433,N_43516,N_48585);
xnor UO_2434 (O_2434,N_43699,N_40658);
or UO_2435 (O_2435,N_40600,N_46898);
or UO_2436 (O_2436,N_46113,N_49874);
and UO_2437 (O_2437,N_49485,N_47624);
or UO_2438 (O_2438,N_41771,N_49808);
nand UO_2439 (O_2439,N_46436,N_44127);
xor UO_2440 (O_2440,N_46540,N_47887);
and UO_2441 (O_2441,N_41485,N_44402);
nand UO_2442 (O_2442,N_40488,N_46314);
nor UO_2443 (O_2443,N_41250,N_40886);
nand UO_2444 (O_2444,N_43081,N_43419);
nor UO_2445 (O_2445,N_49350,N_42090);
nand UO_2446 (O_2446,N_49768,N_45785);
or UO_2447 (O_2447,N_40130,N_46613);
and UO_2448 (O_2448,N_46365,N_40797);
or UO_2449 (O_2449,N_47676,N_44042);
and UO_2450 (O_2450,N_43225,N_45302);
nand UO_2451 (O_2451,N_48531,N_45500);
nand UO_2452 (O_2452,N_42260,N_43103);
or UO_2453 (O_2453,N_48367,N_44664);
and UO_2454 (O_2454,N_45773,N_45143);
nor UO_2455 (O_2455,N_45961,N_41040);
nor UO_2456 (O_2456,N_45289,N_40499);
nor UO_2457 (O_2457,N_44200,N_45633);
and UO_2458 (O_2458,N_41012,N_48110);
nand UO_2459 (O_2459,N_46863,N_43829);
nand UO_2460 (O_2460,N_40069,N_48971);
and UO_2461 (O_2461,N_43705,N_49419);
nand UO_2462 (O_2462,N_42063,N_48079);
and UO_2463 (O_2463,N_49133,N_42829);
nor UO_2464 (O_2464,N_40300,N_46145);
and UO_2465 (O_2465,N_45655,N_42871);
and UO_2466 (O_2466,N_48231,N_47599);
nand UO_2467 (O_2467,N_44652,N_41286);
xnor UO_2468 (O_2468,N_40780,N_48473);
nand UO_2469 (O_2469,N_49885,N_49656);
nor UO_2470 (O_2470,N_40456,N_46674);
or UO_2471 (O_2471,N_42819,N_44086);
and UO_2472 (O_2472,N_45468,N_43432);
and UO_2473 (O_2473,N_41790,N_47483);
or UO_2474 (O_2474,N_43375,N_44679);
or UO_2475 (O_2475,N_46946,N_43747);
and UO_2476 (O_2476,N_40158,N_42296);
nor UO_2477 (O_2477,N_47674,N_44103);
nand UO_2478 (O_2478,N_44335,N_42118);
nor UO_2479 (O_2479,N_46631,N_43859);
and UO_2480 (O_2480,N_41159,N_46414);
nor UO_2481 (O_2481,N_46534,N_45294);
nor UO_2482 (O_2482,N_41776,N_45003);
nor UO_2483 (O_2483,N_41063,N_41203);
nand UO_2484 (O_2484,N_42051,N_47470);
or UO_2485 (O_2485,N_42655,N_41582);
nand UO_2486 (O_2486,N_41151,N_49024);
nor UO_2487 (O_2487,N_48452,N_40259);
nor UO_2488 (O_2488,N_45878,N_49154);
or UO_2489 (O_2489,N_48154,N_47965);
or UO_2490 (O_2490,N_42381,N_43055);
nor UO_2491 (O_2491,N_45778,N_40969);
nand UO_2492 (O_2492,N_41412,N_45540);
or UO_2493 (O_2493,N_48914,N_46076);
nor UO_2494 (O_2494,N_41704,N_45214);
or UO_2495 (O_2495,N_42283,N_47124);
nand UO_2496 (O_2496,N_41277,N_45202);
and UO_2497 (O_2497,N_47662,N_47712);
or UO_2498 (O_2498,N_45617,N_43406);
nor UO_2499 (O_2499,N_44694,N_42556);
and UO_2500 (O_2500,N_46046,N_49848);
nand UO_2501 (O_2501,N_46087,N_48344);
or UO_2502 (O_2502,N_44730,N_45347);
nand UO_2503 (O_2503,N_46910,N_43265);
nor UO_2504 (O_2504,N_40359,N_40028);
and UO_2505 (O_2505,N_41071,N_40381);
and UO_2506 (O_2506,N_48214,N_44918);
or UO_2507 (O_2507,N_49053,N_49689);
nand UO_2508 (O_2508,N_47922,N_46275);
nor UO_2509 (O_2509,N_46654,N_45332);
and UO_2510 (O_2510,N_49936,N_42656);
xor UO_2511 (O_2511,N_48923,N_45529);
and UO_2512 (O_2512,N_40730,N_44485);
nor UO_2513 (O_2513,N_45715,N_49855);
and UO_2514 (O_2514,N_42222,N_41830);
and UO_2515 (O_2515,N_42387,N_45351);
or UO_2516 (O_2516,N_42662,N_43524);
xnor UO_2517 (O_2517,N_40620,N_40946);
or UO_2518 (O_2518,N_42207,N_42137);
and UO_2519 (O_2519,N_45796,N_43059);
and UO_2520 (O_2520,N_43918,N_41257);
or UO_2521 (O_2521,N_45683,N_49264);
nor UO_2522 (O_2522,N_47301,N_47496);
or UO_2523 (O_2523,N_44534,N_41349);
xnor UO_2524 (O_2524,N_47660,N_41113);
nand UO_2525 (O_2525,N_43407,N_40386);
nor UO_2526 (O_2526,N_49426,N_44417);
and UO_2527 (O_2527,N_41605,N_46292);
nand UO_2528 (O_2528,N_48625,N_42858);
xor UO_2529 (O_2529,N_47385,N_45560);
xnor UO_2530 (O_2530,N_42227,N_44561);
nand UO_2531 (O_2531,N_49641,N_41529);
or UO_2532 (O_2532,N_40461,N_46672);
xor UO_2533 (O_2533,N_49547,N_45534);
or UO_2534 (O_2534,N_45436,N_44971);
nor UO_2535 (O_2535,N_44859,N_47589);
and UO_2536 (O_2536,N_45624,N_47566);
and UO_2537 (O_2537,N_40491,N_49297);
or UO_2538 (O_2538,N_45071,N_42463);
or UO_2539 (O_2539,N_49516,N_45759);
xnor UO_2540 (O_2540,N_48948,N_44365);
nor UO_2541 (O_2541,N_48505,N_48134);
nand UO_2542 (O_2542,N_48892,N_45508);
nor UO_2543 (O_2543,N_43336,N_40173);
or UO_2544 (O_2544,N_42789,N_49651);
nor UO_2545 (O_2545,N_40050,N_47479);
or UO_2546 (O_2546,N_45734,N_46735);
nor UO_2547 (O_2547,N_42329,N_40352);
nand UO_2548 (O_2548,N_47870,N_46464);
and UO_2549 (O_2549,N_48242,N_49110);
and UO_2550 (O_2550,N_49819,N_46327);
or UO_2551 (O_2551,N_45410,N_43783);
nor UO_2552 (O_2552,N_42286,N_40154);
nand UO_2553 (O_2553,N_44247,N_44138);
nor UO_2554 (O_2554,N_43494,N_49873);
and UO_2555 (O_2555,N_40156,N_45378);
nor UO_2556 (O_2556,N_42832,N_41981);
or UO_2557 (O_2557,N_47961,N_42951);
nor UO_2558 (O_2558,N_40870,N_43897);
xor UO_2559 (O_2559,N_49882,N_42883);
or UO_2560 (O_2560,N_47815,N_42944);
nand UO_2561 (O_2561,N_41662,N_40137);
nor UO_2562 (O_2562,N_41580,N_44142);
nor UO_2563 (O_2563,N_48346,N_40504);
or UO_2564 (O_2564,N_49251,N_45267);
nor UO_2565 (O_2565,N_45505,N_43992);
nor UO_2566 (O_2566,N_40289,N_45475);
and UO_2567 (O_2567,N_40587,N_44046);
and UO_2568 (O_2568,N_42095,N_48792);
xnor UO_2569 (O_2569,N_49163,N_47847);
and UO_2570 (O_2570,N_46529,N_41427);
nand UO_2571 (O_2571,N_43964,N_49560);
nand UO_2572 (O_2572,N_42842,N_47488);
nand UO_2573 (O_2573,N_45605,N_47187);
nand UO_2574 (O_2574,N_46416,N_42931);
nor UO_2575 (O_2575,N_48588,N_40519);
or UO_2576 (O_2576,N_45844,N_43914);
nand UO_2577 (O_2577,N_41177,N_47098);
nand UO_2578 (O_2578,N_41035,N_41148);
or UO_2579 (O_2579,N_48304,N_46650);
nor UO_2580 (O_2580,N_48545,N_48868);
nand UO_2581 (O_2581,N_41367,N_47867);
nor UO_2582 (O_2582,N_46230,N_40546);
nor UO_2583 (O_2583,N_45660,N_44260);
nor UO_2584 (O_2584,N_46371,N_42886);
and UO_2585 (O_2585,N_41337,N_46224);
or UO_2586 (O_2586,N_42203,N_45069);
or UO_2587 (O_2587,N_46891,N_40741);
xor UO_2588 (O_2588,N_46188,N_40789);
and UO_2589 (O_2589,N_45164,N_48607);
or UO_2590 (O_2590,N_48241,N_45742);
or UO_2591 (O_2591,N_48397,N_45953);
xnor UO_2592 (O_2592,N_40859,N_46164);
xor UO_2593 (O_2593,N_42980,N_48712);
nor UO_2594 (O_2594,N_48451,N_48109);
xnor UO_2595 (O_2595,N_42310,N_49732);
or UO_2596 (O_2596,N_46588,N_43322);
nand UO_2597 (O_2597,N_47831,N_42452);
or UO_2598 (O_2598,N_47294,N_45173);
nand UO_2599 (O_2599,N_43753,N_40930);
and UO_2600 (O_2600,N_44299,N_42564);
nand UO_2601 (O_2601,N_44835,N_41145);
or UO_2602 (O_2602,N_47304,N_48162);
nand UO_2603 (O_2603,N_44992,N_42714);
nor UO_2604 (O_2604,N_46363,N_48135);
nor UO_2605 (O_2605,N_41908,N_47462);
xnor UO_2606 (O_2606,N_41891,N_44067);
or UO_2607 (O_2607,N_42835,N_48276);
xor UO_2608 (O_2608,N_44023,N_47956);
nor UO_2609 (O_2609,N_43911,N_48224);
nand UO_2610 (O_2610,N_45421,N_41227);
nand UO_2611 (O_2611,N_40924,N_43670);
nand UO_2612 (O_2612,N_45604,N_44308);
nand UO_2613 (O_2613,N_48250,N_40351);
and UO_2614 (O_2614,N_48386,N_49250);
xor UO_2615 (O_2615,N_48834,N_42702);
or UO_2616 (O_2616,N_40594,N_49551);
or UO_2617 (O_2617,N_42363,N_41705);
nor UO_2618 (O_2618,N_48430,N_46284);
and UO_2619 (O_2619,N_48097,N_47580);
and UO_2620 (O_2620,N_46283,N_46518);
nand UO_2621 (O_2621,N_40077,N_43364);
nand UO_2622 (O_2622,N_42571,N_43333);
nand UO_2623 (O_2623,N_44075,N_44266);
nor UO_2624 (O_2624,N_45766,N_47454);
nor UO_2625 (O_2625,N_41114,N_45105);
and UO_2626 (O_2626,N_48916,N_42922);
nand UO_2627 (O_2627,N_47954,N_43641);
or UO_2628 (O_2628,N_49682,N_42700);
xor UO_2629 (O_2629,N_42887,N_48091);
nand UO_2630 (O_2630,N_44827,N_41475);
and UO_2631 (O_2631,N_45145,N_40368);
nor UO_2632 (O_2632,N_47175,N_48156);
or UO_2633 (O_2633,N_41715,N_41371);
and UO_2634 (O_2634,N_42274,N_41365);
or UO_2635 (O_2635,N_44235,N_41883);
nor UO_2636 (O_2636,N_49042,N_49187);
and UO_2637 (O_2637,N_49574,N_47598);
nand UO_2638 (O_2638,N_41239,N_44709);
and UO_2639 (O_2639,N_42459,N_42014);
or UO_2640 (O_2640,N_46467,N_44895);
nand UO_2641 (O_2641,N_41052,N_42529);
and UO_2642 (O_2642,N_46928,N_41312);
and UO_2643 (O_2643,N_41332,N_49923);
nor UO_2644 (O_2644,N_46696,N_43853);
nand UO_2645 (O_2645,N_48842,N_45754);
and UO_2646 (O_2646,N_47285,N_48960);
or UO_2647 (O_2647,N_45577,N_47567);
and UO_2648 (O_2648,N_49606,N_47749);
nor UO_2649 (O_2649,N_48887,N_42252);
nor UO_2650 (O_2650,N_40239,N_45004);
or UO_2651 (O_2651,N_42218,N_45578);
nor UO_2652 (O_2652,N_46544,N_45067);
or UO_2653 (O_2653,N_42016,N_43741);
or UO_2654 (O_2654,N_41006,N_46091);
nand UO_2655 (O_2655,N_48809,N_46089);
nand UO_2656 (O_2656,N_41399,N_48288);
and UO_2657 (O_2657,N_45671,N_49334);
and UO_2658 (O_2658,N_41223,N_44515);
nor UO_2659 (O_2659,N_45939,N_46947);
nand UO_2660 (O_2660,N_44722,N_43056);
xnor UO_2661 (O_2661,N_44268,N_42239);
xor UO_2662 (O_2662,N_44228,N_41952);
or UO_2663 (O_2663,N_49513,N_44706);
or UO_2664 (O_2664,N_46893,N_40782);
nand UO_2665 (O_2665,N_40877,N_46794);
and UO_2666 (O_2666,N_47555,N_44265);
and UO_2667 (O_2667,N_45090,N_48605);
nand UO_2668 (O_2668,N_47809,N_42098);
or UO_2669 (O_2669,N_48268,N_44637);
or UO_2670 (O_2670,N_46459,N_48976);
or UO_2671 (O_2671,N_43004,N_49529);
nand UO_2672 (O_2672,N_41238,N_49810);
nand UO_2673 (O_2673,N_49658,N_40804);
nor UO_2674 (O_2674,N_48707,N_49786);
and UO_2675 (O_2675,N_46673,N_41725);
xnor UO_2676 (O_2676,N_44993,N_41858);
and UO_2677 (O_2677,N_48575,N_40206);
nor UO_2678 (O_2678,N_44535,N_40114);
nand UO_2679 (O_2679,N_44463,N_45085);
nor UO_2680 (O_2680,N_48938,N_46853);
nor UO_2681 (O_2681,N_48580,N_42482);
nor UO_2682 (O_2682,N_43972,N_40479);
and UO_2683 (O_2683,N_46504,N_44669);
or UO_2684 (O_2684,N_43091,N_44588);
nand UO_2685 (O_2685,N_42391,N_49054);
nand UO_2686 (O_2686,N_41898,N_43411);
or UO_2687 (O_2687,N_41139,N_48085);
nand UO_2688 (O_2688,N_41003,N_44967);
and UO_2689 (O_2689,N_40747,N_41958);
and UO_2690 (O_2690,N_49451,N_43863);
nor UO_2691 (O_2691,N_40141,N_47984);
xor UO_2692 (O_2692,N_48730,N_43813);
and UO_2693 (O_2693,N_49693,N_40679);
nor UO_2694 (O_2694,N_46191,N_45010);
xor UO_2695 (O_2695,N_49145,N_41800);
nor UO_2696 (O_2696,N_47256,N_40003);
nand UO_2697 (O_2697,N_46361,N_44122);
or UO_2698 (O_2698,N_44636,N_45718);
and UO_2699 (O_2699,N_43576,N_47157);
nor UO_2700 (O_2700,N_45903,N_48872);
and UO_2701 (O_2701,N_40345,N_46478);
or UO_2702 (O_2702,N_42593,N_43122);
nand UO_2703 (O_2703,N_47156,N_41527);
and UO_2704 (O_2704,N_42552,N_44250);
or UO_2705 (O_2705,N_49435,N_41739);
nand UO_2706 (O_2706,N_45367,N_41341);
nor UO_2707 (O_2707,N_42595,N_48530);
nor UO_2708 (O_2708,N_49325,N_41974);
nand UO_2709 (O_2709,N_46181,N_42184);
nand UO_2710 (O_2710,N_48599,N_42301);
nand UO_2711 (O_2711,N_47332,N_47068);
and UO_2712 (O_2712,N_45597,N_45680);
or UO_2713 (O_2713,N_42358,N_49222);
or UO_2714 (O_2714,N_44084,N_45651);
nor UO_2715 (O_2715,N_45506,N_47169);
nand UO_2716 (O_2716,N_46336,N_48735);
and UO_2717 (O_2717,N_43430,N_40234);
or UO_2718 (O_2718,N_49180,N_47684);
nor UO_2719 (O_2719,N_46071,N_41472);
or UO_2720 (O_2720,N_41360,N_45471);
nor UO_2721 (O_2721,N_48358,N_44154);
and UO_2722 (O_2722,N_43451,N_40991);
and UO_2723 (O_2723,N_45951,N_49943);
nand UO_2724 (O_2724,N_49860,N_45498);
xor UO_2725 (O_2725,N_42160,N_48713);
nand UO_2726 (O_2726,N_43629,N_47324);
xor UO_2727 (O_2727,N_44799,N_44592);
and UO_2728 (O_2728,N_41350,N_45717);
nor UO_2729 (O_2729,N_48504,N_48118);
or UO_2730 (O_2730,N_45151,N_46877);
nor UO_2731 (O_2731,N_47151,N_47647);
xnor UO_2732 (O_2732,N_43236,N_47525);
and UO_2733 (O_2733,N_48619,N_46943);
and UO_2734 (O_2734,N_42493,N_41953);
and UO_2735 (O_2735,N_47950,N_40170);
xor UO_2736 (O_2736,N_42432,N_43876);
and UO_2737 (O_2737,N_43565,N_49640);
nand UO_2738 (O_2738,N_43888,N_40318);
or UO_2739 (O_2739,N_40459,N_43266);
nand UO_2740 (O_2740,N_46765,N_44461);
or UO_2741 (O_2741,N_45279,N_42757);
nand UO_2742 (O_2742,N_45247,N_43541);
xor UO_2743 (O_2743,N_43323,N_40656);
or UO_2744 (O_2744,N_43069,N_43648);
or UO_2745 (O_2745,N_45980,N_43685);
or UO_2746 (O_2746,N_48548,N_48099);
nor UO_2747 (O_2747,N_44617,N_48956);
and UO_2748 (O_2748,N_48014,N_47845);
and UO_2749 (O_2749,N_48420,N_41626);
and UO_2750 (O_2750,N_49482,N_46664);
nor UO_2751 (O_2751,N_43917,N_40538);
or UO_2752 (O_2752,N_44065,N_45856);
nand UO_2753 (O_2753,N_46118,N_41574);
or UO_2754 (O_2754,N_47651,N_45203);
nand UO_2755 (O_2755,N_44350,N_43124);
nand UO_2756 (O_2756,N_48142,N_43433);
and UO_2757 (O_2757,N_41439,N_41008);
xnor UO_2758 (O_2758,N_46296,N_48949);
nor UO_2759 (O_2759,N_49336,N_40152);
or UO_2760 (O_2760,N_43902,N_47047);
nand UO_2761 (O_2761,N_41345,N_46606);
or UO_2762 (O_2762,N_49903,N_45746);
or UO_2763 (O_2763,N_48187,N_47960);
xnor UO_2764 (O_2764,N_42037,N_45967);
nor UO_2765 (O_2765,N_43997,N_45881);
xnor UO_2766 (O_2766,N_42249,N_43594);
and UO_2767 (O_2767,N_42998,N_46596);
nor UO_2768 (O_2768,N_43579,N_43781);
or UO_2769 (O_2769,N_43064,N_41085);
nor UO_2770 (O_2770,N_41380,N_46517);
nand UO_2771 (O_2771,N_43692,N_48247);
nor UO_2772 (O_2772,N_49680,N_49566);
nor UO_2773 (O_2773,N_49992,N_42047);
or UO_2774 (O_2774,N_42550,N_45664);
or UO_2775 (O_2775,N_49624,N_43643);
nor UO_2776 (O_2776,N_46469,N_40397);
or UO_2777 (O_2777,N_42734,N_43903);
nand UO_2778 (O_2778,N_49059,N_47641);
nor UO_2779 (O_2779,N_41184,N_40155);
xnor UO_2780 (O_2780,N_48402,N_44385);
nor UO_2781 (O_2781,N_46745,N_44025);
nor UO_2782 (O_2782,N_48361,N_48453);
nand UO_2783 (O_2783,N_46346,N_46505);
or UO_2784 (O_2784,N_42231,N_45283);
or UO_2785 (O_2785,N_45414,N_48627);
nand UO_2786 (O_2786,N_46330,N_48518);
nor UO_2787 (O_2787,N_45127,N_44671);
nor UO_2788 (O_2788,N_46221,N_49300);
and UO_2789 (O_2789,N_44315,N_42212);
and UO_2790 (O_2790,N_43506,N_41468);
or UO_2791 (O_2791,N_44237,N_49892);
or UO_2792 (O_2792,N_41407,N_47563);
and UO_2793 (O_2793,N_49105,N_43785);
or UO_2794 (O_2794,N_48780,N_41865);
nor UO_2795 (O_2795,N_48183,N_44574);
nand UO_2796 (O_2796,N_43674,N_45199);
nand UO_2797 (O_2797,N_49258,N_41037);
and UO_2798 (O_2798,N_42490,N_42464);
nor UO_2799 (O_2799,N_49127,N_46563);
nor UO_2800 (O_2800,N_46196,N_49278);
nor UO_2801 (O_2801,N_42302,N_41670);
nor UO_2802 (O_2802,N_47972,N_42666);
and UO_2803 (O_2803,N_40446,N_40236);
or UO_2804 (O_2804,N_46685,N_47107);
nand UO_2805 (O_2805,N_45103,N_47855);
nand UO_2806 (O_2806,N_40006,N_46692);
xor UO_2807 (O_2807,N_43118,N_45859);
nor UO_2808 (O_2808,N_41651,N_48807);
or UO_2809 (O_2809,N_47775,N_43491);
nor UO_2810 (O_2810,N_40455,N_46169);
or UO_2811 (O_2811,N_44119,N_45309);
nor UO_2812 (O_2812,N_46027,N_44567);
xor UO_2813 (O_2813,N_45942,N_47687);
xor UO_2814 (O_2814,N_48424,N_49915);
or UO_2815 (O_2815,N_48733,N_45501);
nor UO_2816 (O_2816,N_41101,N_40645);
nand UO_2817 (O_2817,N_46360,N_43221);
and UO_2818 (O_2818,N_48502,N_47269);
nand UO_2819 (O_2819,N_45770,N_42268);
xnor UO_2820 (O_2820,N_45993,N_41942);
nand UO_2821 (O_2821,N_45313,N_46568);
and UO_2822 (O_2822,N_43294,N_45764);
and UO_2823 (O_2823,N_44912,N_43904);
nand UO_2824 (O_2824,N_49490,N_43590);
xor UO_2825 (O_2825,N_42643,N_48825);
nand UO_2826 (O_2826,N_41579,N_43109);
nand UO_2827 (O_2827,N_46782,N_48562);
nand UO_2828 (O_2828,N_47581,N_47173);
and UO_2829 (O_2829,N_40406,N_42103);
and UO_2830 (O_2830,N_44198,N_47558);
nor UO_2831 (O_2831,N_42605,N_49464);
or UO_2832 (O_2832,N_47968,N_49765);
or UO_2833 (O_2833,N_46112,N_48015);
nor UO_2834 (O_2834,N_46261,N_45909);
nor UO_2835 (O_2835,N_49136,N_49864);
nor UO_2836 (O_2836,N_43507,N_47619);
or UO_2837 (O_2837,N_40934,N_49695);
nand UO_2838 (O_2838,N_42939,N_46638);
or UO_2839 (O_2839,N_40452,N_44443);
xor UO_2840 (O_2840,N_49254,N_41969);
and UO_2841 (O_2841,N_44755,N_42394);
or UO_2842 (O_2842,N_47570,N_40961);
and UO_2843 (O_2843,N_40229,N_48058);
and UO_2844 (O_2844,N_45353,N_44015);
nand UO_2845 (O_2845,N_49737,N_46151);
or UO_2846 (O_2846,N_43884,N_43062);
nand UO_2847 (O_2847,N_49406,N_48294);
and UO_2848 (O_2848,N_43910,N_43528);
xor UO_2849 (O_2849,N_44107,N_47436);
nor UO_2850 (O_2850,N_41886,N_44950);
xor UO_2851 (O_2851,N_46578,N_48481);
xor UO_2852 (O_2852,N_40537,N_45665);
and UO_2853 (O_2853,N_48779,N_42078);
nor UO_2854 (O_2854,N_44036,N_45711);
or UO_2855 (O_2855,N_44885,N_44692);
or UO_2856 (O_2856,N_43373,N_43555);
nand UO_2857 (O_2857,N_48969,N_48566);
nand UO_2858 (O_2858,N_40965,N_46784);
nor UO_2859 (O_2859,N_42636,N_42528);
and UO_2860 (O_2860,N_43354,N_42304);
and UO_2861 (O_2861,N_46595,N_41864);
and UO_2862 (O_2862,N_42291,N_41794);
or UO_2863 (O_2863,N_45499,N_42485);
nor UO_2864 (O_2864,N_43437,N_40408);
xnor UO_2865 (O_2865,N_42750,N_41755);
or UO_2866 (O_2866,N_43438,N_46850);
or UO_2867 (O_2867,N_42035,N_49826);
nor UO_2868 (O_2868,N_48679,N_47251);
and UO_2869 (O_2869,N_42896,N_43772);
nand UO_2870 (O_2870,N_49141,N_46097);
or UO_2871 (O_2871,N_46500,N_45857);
and UO_2872 (O_2872,N_49621,N_49356);
or UO_2873 (O_2873,N_44848,N_44707);
nor UO_2874 (O_2874,N_48850,N_49982);
and UO_2875 (O_2875,N_49935,N_43542);
or UO_2876 (O_2876,N_47128,N_47913);
nor UO_2877 (O_2877,N_44098,N_46105);
and UO_2878 (O_2878,N_44259,N_41868);
nand UO_2879 (O_2879,N_40878,N_40882);
or UO_2880 (O_2880,N_41714,N_43680);
and UO_2881 (O_2881,N_45082,N_49535);
nand UO_2882 (O_2882,N_44801,N_47177);
nand UO_2883 (O_2883,N_42182,N_41441);
and UO_2884 (O_2884,N_46295,N_46849);
or UO_2885 (O_2885,N_42033,N_45192);
xor UO_2886 (O_2886,N_45635,N_41669);
nor UO_2887 (O_2887,N_46238,N_40769);
nand UO_2888 (O_2888,N_42240,N_46680);
nor UO_2889 (O_2889,N_47808,N_47848);
nand UO_2890 (O_2890,N_49103,N_48848);
xor UO_2891 (O_2891,N_47679,N_47522);
nand UO_2892 (O_2892,N_41946,N_48246);
nor UO_2893 (O_2893,N_48511,N_40262);
or UO_2894 (O_2894,N_47133,N_41209);
nor UO_2895 (O_2895,N_44395,N_42940);
and UO_2896 (O_2896,N_45832,N_49242);
nor UO_2897 (O_2897,N_49803,N_48533);
and UO_2898 (O_2898,N_40394,N_48903);
xor UO_2899 (O_2899,N_42634,N_45995);
or UO_2900 (O_2900,N_48877,N_42317);
nor UO_2901 (O_2901,N_43512,N_48495);
xor UO_2902 (O_2902,N_48598,N_42494);
nand UO_2903 (O_2903,N_48582,N_46554);
and UO_2904 (O_2904,N_42314,N_47246);
xnor UO_2905 (O_2905,N_40070,N_48656);
or UO_2906 (O_2906,N_40030,N_40314);
and UO_2907 (O_2907,N_48983,N_44930);
and UO_2908 (O_2908,N_41827,N_46128);
nor UO_2909 (O_2909,N_49391,N_46070);
or UO_2910 (O_2910,N_41577,N_48528);
or UO_2911 (O_2911,N_40099,N_45721);
nor UO_2912 (O_2912,N_40951,N_45230);
nor UO_2913 (O_2913,N_48046,N_49161);
or UO_2914 (O_2914,N_46826,N_41748);
xnor UO_2915 (O_2915,N_41314,N_45978);
nand UO_2916 (O_2916,N_46636,N_41623);
and UO_2917 (O_2917,N_40899,N_46297);
or UO_2918 (O_2918,N_43366,N_48399);
and UO_2919 (O_2919,N_42165,N_47595);
nor UO_2920 (O_2920,N_46569,N_43016);
and UO_2921 (O_2921,N_45944,N_45200);
or UO_2922 (O_2922,N_48587,N_44702);
nor UO_2923 (O_2923,N_42807,N_48365);
nand UO_2924 (O_2924,N_40203,N_40309);
nand UO_2925 (O_2925,N_41947,N_43525);
or UO_2926 (O_2926,N_40469,N_47781);
or UO_2927 (O_2927,N_40423,N_45046);
or UO_2928 (O_2928,N_45447,N_45466);
or UO_2929 (O_2929,N_44934,N_46433);
or UO_2930 (O_2930,N_40939,N_40920);
xnor UO_2931 (O_2931,N_40250,N_45389);
nand UO_2932 (O_2932,N_44158,N_41746);
or UO_2933 (O_2933,N_41728,N_49130);
nor UO_2934 (O_2934,N_47568,N_40492);
and UO_2935 (O_2935,N_49619,N_41733);
or UO_2936 (O_2936,N_48687,N_42777);
nor UO_2937 (O_2937,N_40395,N_46830);
and UO_2938 (O_2938,N_47216,N_43273);
nor UO_2939 (O_2939,N_44199,N_48130);
and UO_2940 (O_2940,N_45083,N_47724);
xnor UO_2941 (O_2941,N_44659,N_41182);
nand UO_2942 (O_2942,N_46383,N_47084);
nor UO_2943 (O_2943,N_47457,N_46372);
or UO_2944 (O_2944,N_48783,N_42826);
or UO_2945 (O_2945,N_46842,N_49796);
nor UO_2946 (O_2946,N_42809,N_40681);
or UO_2947 (O_2947,N_40238,N_44604);
or UO_2948 (O_2948,N_48428,N_44193);
and UO_2949 (O_2949,N_45996,N_41964);
and UO_2950 (O_2950,N_40315,N_45882);
xnor UO_2951 (O_2951,N_49834,N_49488);
nor UO_2952 (O_2952,N_45714,N_41474);
and UO_2953 (O_2953,N_43701,N_45440);
nor UO_2954 (O_2954,N_47879,N_49630);
nor UO_2955 (O_2955,N_44447,N_40544);
and UO_2956 (O_2956,N_41550,N_46810);
nor UO_2957 (O_2957,N_43786,N_41169);
or UO_2958 (O_2958,N_40123,N_42225);
nor UO_2959 (O_2959,N_42110,N_48729);
and UO_2960 (O_2960,N_45403,N_47562);
or UO_2961 (O_2961,N_40914,N_47024);
nand UO_2962 (O_2962,N_42036,N_40599);
or UO_2963 (O_2963,N_44232,N_44998);
or UO_2964 (O_2964,N_42908,N_40035);
and UO_2965 (O_2965,N_40205,N_47691);
and UO_2966 (O_2966,N_44011,N_46646);
nand UO_2967 (O_2967,N_41928,N_42744);
or UO_2968 (O_2968,N_40296,N_45449);
or UO_2969 (O_2969,N_42029,N_48526);
nor UO_2970 (O_2970,N_48474,N_41050);
nand UO_2971 (O_2971,N_48273,N_40274);
or UO_2972 (O_2972,N_47980,N_47925);
nor UO_2973 (O_2973,N_44213,N_49517);
nor UO_2974 (O_2974,N_46241,N_46356);
and UO_2975 (O_2975,N_45119,N_46385);
and UO_2976 (O_2976,N_49051,N_49557);
nand UO_2977 (O_2977,N_40092,N_49633);
or UO_2978 (O_2978,N_46996,N_45860);
nor UO_2979 (O_2979,N_44282,N_45960);
and UO_2980 (O_2980,N_47758,N_49648);
and UO_2981 (O_2981,N_45925,N_49385);
nand UO_2982 (O_2982,N_47335,N_41716);
nor UO_2983 (O_2983,N_44795,N_48902);
nand UO_2984 (O_2984,N_48211,N_40949);
nand UO_2985 (O_2985,N_48263,N_48907);
nor UO_2986 (O_2986,N_40911,N_45220);
or UO_2987 (O_2987,N_46042,N_41224);
and UO_2988 (O_2988,N_46462,N_41030);
and UO_2989 (O_2989,N_40907,N_41613);
or UO_2990 (O_2990,N_47073,N_40992);
nor UO_2991 (O_2991,N_45987,N_49414);
nor UO_2992 (O_2992,N_43951,N_42350);
nor UO_2993 (O_2993,N_44083,N_42420);
and UO_2994 (O_2994,N_44307,N_43544);
and UO_2995 (O_2995,N_43545,N_46345);
and UO_2996 (O_2996,N_42880,N_47214);
nand UO_2997 (O_2997,N_47654,N_48849);
nand UO_2998 (O_2998,N_49811,N_47127);
or UO_2999 (O_2999,N_41749,N_48968);
and UO_3000 (O_3000,N_49845,N_41325);
xor UO_3001 (O_3001,N_41070,N_48691);
nand UO_3002 (O_3002,N_46705,N_48387);
and UO_3003 (O_3003,N_41525,N_45078);
nand UO_3004 (O_3004,N_46667,N_41956);
and UO_3005 (O_3005,N_42242,N_47193);
or UO_3006 (O_3006,N_47659,N_47428);
and UO_3007 (O_3007,N_44589,N_44311);
nand UO_3008 (O_3008,N_47002,N_41653);
and UO_3009 (O_3009,N_45094,N_49031);
nor UO_3010 (O_3010,N_42537,N_49313);
or UO_3011 (O_3011,N_44860,N_45575);
nand UO_3012 (O_3012,N_44360,N_41738);
and UO_3013 (O_3013,N_41208,N_42092);
nand UO_3014 (O_3014,N_49316,N_48401);
xor UO_3015 (O_3015,N_40590,N_44977);
nand UO_3016 (O_3016,N_45594,N_42091);
xor UO_3017 (O_3017,N_41904,N_47083);
and UO_3018 (O_3018,N_44943,N_43646);
nor UO_3019 (O_3019,N_41112,N_47033);
nor UO_3020 (O_3020,N_47635,N_42174);
and UO_3021 (O_3021,N_42144,N_43733);
and UO_3022 (O_3022,N_46864,N_40760);
or UO_3023 (O_3023,N_46202,N_47588);
and UO_3024 (O_3024,N_41982,N_40011);
and UO_3025 (O_3025,N_42177,N_45025);
nand UO_3026 (O_3026,N_48614,N_47894);
and UO_3027 (O_3027,N_49033,N_46485);
nor UO_3028 (O_3028,N_43522,N_44874);
nor UO_3029 (O_3029,N_43148,N_49754);
nor UO_3030 (O_3030,N_47288,N_41436);
nor UO_3031 (O_3031,N_47934,N_47587);
and UO_3032 (O_3032,N_49019,N_49895);
and UO_3033 (O_3033,N_44041,N_43239);
nor UO_3034 (O_3034,N_41397,N_47367);
and UO_3035 (O_3035,N_47088,N_42061);
nor UO_3036 (O_3036,N_41243,N_40548);
nand UO_3037 (O_3037,N_49159,N_41176);
nor UO_3038 (O_3038,N_49431,N_43368);
or UO_3039 (O_3039,N_40473,N_43351);
or UO_3040 (O_3040,N_41901,N_46165);
and UO_3041 (O_3041,N_41912,N_41533);
nor UO_3042 (O_3042,N_43051,N_40684);
and UO_3043 (O_3043,N_42758,N_47371);
nand UO_3044 (O_3044,N_40193,N_49332);
nor UO_3045 (O_3045,N_49455,N_45900);
nand UO_3046 (O_3046,N_42470,N_42812);
or UO_3047 (O_3047,N_47672,N_41136);
nand UO_3048 (O_3048,N_49041,N_48251);
nor UO_3049 (O_3049,N_43274,N_47670);
and UO_3050 (O_3050,N_46904,N_42451);
and UO_3051 (O_3051,N_49299,N_40000);
or UO_3052 (O_3052,N_47360,N_45418);
or UO_3053 (O_3053,N_47263,N_43414);
nor UO_3054 (O_3054,N_42762,N_44504);
nand UO_3055 (O_3055,N_43161,N_46608);
and UO_3056 (O_3056,N_45491,N_47783);
nand UO_3057 (O_3057,N_44787,N_42570);
nand UO_3058 (O_3058,N_40643,N_44957);
nand UO_3059 (O_3059,N_40752,N_47148);
nor UO_3060 (O_3060,N_49976,N_48740);
nand UO_3061 (O_3061,N_44648,N_42601);
and UO_3062 (O_3062,N_41339,N_49301);
nor UO_3063 (O_3063,N_43571,N_42285);
and UO_3064 (O_3064,N_43547,N_45652);
nor UO_3065 (O_3065,N_40336,N_45645);
or UO_3066 (O_3066,N_48717,N_40304);
nand UO_3067 (O_3067,N_41241,N_43819);
and UO_3068 (O_3068,N_47338,N_40119);
or UO_3069 (O_3069,N_40432,N_41622);
nand UO_3070 (O_3070,N_48018,N_49740);
and UO_3071 (O_3071,N_47064,N_48372);
or UO_3072 (O_3072,N_49305,N_44149);
nor UO_3073 (O_3073,N_49637,N_43021);
xnor UO_3074 (O_3074,N_47366,N_41815);
nand UO_3075 (O_3075,N_40637,N_48448);
nand UO_3076 (O_3076,N_49847,N_48319);
nor UO_3077 (O_3077,N_49115,N_46158);
nor UO_3078 (O_3078,N_47441,N_42343);
nor UO_3079 (O_3079,N_49144,N_41465);
nand UO_3080 (O_3080,N_48443,N_45311);
nand UO_3081 (O_3081,N_49511,N_49018);
nand UO_3082 (O_3082,N_41978,N_49524);
nand UO_3083 (O_3083,N_42776,N_42318);
xnor UO_3084 (O_3084,N_40827,N_48469);
and UO_3085 (O_3085,N_43777,N_48977);
nand UO_3086 (O_3086,N_42805,N_44945);
nor UO_3087 (O_3087,N_49789,N_47390);
xor UO_3088 (O_3088,N_48694,N_41590);
nor UO_3089 (O_3089,N_45522,N_48326);
or UO_3090 (O_3090,N_43668,N_46317);
and UO_3091 (O_3091,N_47025,N_43479);
or UO_3092 (O_3092,N_46392,N_47155);
xor UO_3093 (O_3093,N_40102,N_48616);
or UO_3094 (O_3094,N_45106,N_49777);
and UO_3095 (O_3095,N_49465,N_42346);
xor UO_3096 (O_3096,N_44806,N_44803);
nand UO_3097 (O_3097,N_46914,N_44341);
nor UO_3098 (O_3098,N_41501,N_45975);
and UO_3099 (O_3099,N_46884,N_49571);
nand UO_3100 (O_3100,N_49997,N_48370);
xor UO_3101 (O_3101,N_49916,N_49795);
nand UO_3102 (O_3102,N_44690,N_41247);
and UO_3103 (O_3103,N_49373,N_49001);
or UO_3104 (O_3104,N_49852,N_47037);
nor UO_3105 (O_3105,N_48813,N_42867);
nand UO_3106 (O_3106,N_46835,N_42519);
xor UO_3107 (O_3107,N_44786,N_46972);
nor UO_3108 (O_3108,N_42827,N_49003);
nand UO_3109 (O_3109,N_44396,N_41225);
nand UO_3110 (O_3110,N_41045,N_46591);
nor UO_3111 (O_3111,N_40818,N_48151);
nand UO_3112 (O_3112,N_49068,N_41125);
and UO_3113 (O_3113,N_42241,N_40472);
xor UO_3114 (O_3114,N_43828,N_43595);
nor UO_3115 (O_3115,N_41939,N_43380);
or UO_3116 (O_3116,N_43624,N_47350);
and UO_3117 (O_3117,N_44554,N_45816);
nand UO_3118 (O_3118,N_48876,N_47007);
nor UO_3119 (O_3119,N_46080,N_47411);
and UO_3120 (O_3120,N_46119,N_49022);
and UO_3121 (O_3121,N_47276,N_48210);
nor UO_3122 (O_3122,N_43463,N_49780);
nor UO_3123 (O_3123,N_43658,N_47541);
nand UO_3124 (O_3124,N_47477,N_49778);
or UO_3125 (O_3125,N_45850,N_42072);
nand UO_3126 (O_3126,N_49797,N_40363);
nand UO_3127 (O_3127,N_46103,N_47492);
or UO_3128 (O_3128,N_42255,N_44087);
and UO_3129 (O_3129,N_47718,N_48738);
nor UO_3130 (O_3130,N_45595,N_46886);
or UO_3131 (O_3131,N_40746,N_47706);
nor UO_3132 (O_3132,N_44572,N_43176);
and UO_3133 (O_3133,N_43878,N_47463);
nor UO_3134 (O_3134,N_49686,N_43633);
and UO_3135 (O_3135,N_47875,N_46865);
nand UO_3136 (O_3136,N_45803,N_46263);
nor UO_3137 (O_3137,N_41549,N_47901);
and UO_3138 (O_3138,N_40222,N_41989);
xnor UO_3139 (O_3139,N_47013,N_47410);
and UO_3140 (O_3140,N_47004,N_40649);
nor UO_3141 (O_3141,N_49837,N_42543);
and UO_3142 (O_3142,N_41853,N_49818);
or UO_3143 (O_3143,N_41645,N_47232);
and UO_3144 (O_3144,N_44246,N_49239);
nor UO_3145 (O_3145,N_42791,N_42018);
or UO_3146 (O_3146,N_49311,N_41056);
nand UO_3147 (O_3147,N_40994,N_49667);
or UO_3148 (O_3148,N_48628,N_42538);
or UO_3149 (O_3149,N_44106,N_47539);
nand UO_3150 (O_3150,N_46125,N_40072);
or UO_3151 (O_3151,N_45849,N_41693);
nor UO_3152 (O_3152,N_42496,N_46135);
nand UO_3153 (O_3153,N_40500,N_48698);
or UO_3154 (O_3154,N_40147,N_47969);
xnor UO_3155 (O_3155,N_41134,N_48317);
nor UO_3156 (O_3156,N_41293,N_43300);
nor UO_3157 (O_3157,N_49047,N_40266);
or UO_3158 (O_3158,N_40198,N_42123);
or UO_3159 (O_3159,N_49386,N_41121);
nor UO_3160 (O_3160,N_40330,N_41765);
nand UO_3161 (O_3161,N_48301,N_41668);
nor UO_3162 (O_3162,N_47851,N_45912);
xor UO_3163 (O_3163,N_42431,N_43349);
and UO_3164 (O_3164,N_40213,N_47217);
nor UO_3165 (O_3165,N_41996,N_46127);
or UO_3166 (O_3166,N_43947,N_43143);
xnor UO_3167 (O_3167,N_45609,N_49857);
nor UO_3168 (O_3168,N_49616,N_48328);
nor UO_3169 (O_3169,N_45982,N_40172);
or UO_3170 (O_3170,N_48781,N_47853);
and UO_3171 (O_3171,N_41517,N_48681);
and UO_3172 (O_3172,N_45753,N_46132);
nand UO_3173 (O_3173,N_40278,N_40063);
nor UO_3174 (O_3174,N_49956,N_46199);
nand UO_3175 (O_3175,N_45631,N_42555);
and UO_3176 (O_3176,N_41073,N_46731);
and UO_3177 (O_3177,N_40121,N_41256);
or UO_3178 (O_3178,N_49770,N_45350);
and UO_3179 (O_3179,N_41219,N_47884);
or UO_3180 (O_3180,N_40880,N_41586);
or UO_3181 (O_3181,N_44420,N_42195);
xnor UO_3182 (O_3182,N_49025,N_49489);
nand UO_3183 (O_3183,N_45954,N_45827);
and UO_3184 (O_3184,N_48512,N_42793);
xnor UO_3185 (O_3185,N_42419,N_41278);
nand UO_3186 (O_3186,N_45768,N_42927);
nand UO_3187 (O_3187,N_44066,N_41897);
or UO_3188 (O_3188,N_43256,N_40012);
and UO_3189 (O_3189,N_42775,N_47392);
and UO_3190 (O_3190,N_45075,N_41834);
nor UO_3191 (O_3191,N_40725,N_41228);
nand UO_3192 (O_3192,N_49626,N_42737);
and UO_3193 (O_3193,N_49608,N_42520);
nor UO_3194 (O_3194,N_40888,N_48095);
nor UO_3195 (O_3195,N_47203,N_47898);
xnor UO_3196 (O_3196,N_49595,N_48331);
and UO_3197 (O_3197,N_42701,N_41639);
nor UO_3198 (O_3198,N_40592,N_48569);
xnor UO_3199 (O_3199,N_49842,N_44734);
nand UO_3200 (O_3200,N_41165,N_45625);
or UO_3201 (O_3201,N_45914,N_48696);
nor UO_3202 (O_3202,N_40024,N_40529);
nor UO_3203 (O_3203,N_40015,N_46450);
or UO_3204 (O_3204,N_43605,N_48093);
and UO_3205 (O_3205,N_40405,N_40462);
or UO_3206 (O_3206,N_43139,N_43213);
xnor UO_3207 (O_3207,N_46623,N_43077);
and UO_3208 (O_3208,N_49739,N_45713);
nor UO_3209 (O_3209,N_49743,N_41857);
nand UO_3210 (O_3210,N_44854,N_40836);
or UO_3211 (O_3211,N_45284,N_49957);
xnor UO_3212 (O_3212,N_48279,N_40757);
and UO_3213 (O_3213,N_41554,N_46109);
nor UO_3214 (O_3214,N_48581,N_49323);
nand UO_3215 (O_3215,N_49100,N_42657);
nand UO_3216 (O_3216,N_42011,N_48806);
and UO_3217 (O_3217,N_47316,N_48349);
or UO_3218 (O_3218,N_40216,N_46093);
nor UO_3219 (O_3219,N_43478,N_41026);
or UO_3220 (O_3220,N_45991,N_40464);
nand UO_3221 (O_3221,N_43789,N_49246);
xnor UO_3222 (O_3222,N_46489,N_40791);
nor UO_3223 (O_3223,N_42955,N_49618);
nor UO_3224 (O_3224,N_44296,N_49896);
nor UO_3225 (O_3225,N_42460,N_42579);
nand UO_3226 (O_3226,N_43587,N_41829);
and UO_3227 (O_3227,N_46670,N_41560);
or UO_3228 (O_3228,N_49357,N_40573);
xnor UO_3229 (O_3229,N_45952,N_49236);
nand UO_3230 (O_3230,N_44624,N_40340);
or UO_3231 (O_3231,N_48556,N_49905);
or UO_3232 (O_3232,N_40542,N_47844);
or UO_3233 (O_3233,N_47817,N_43012);
or UO_3234 (O_3234,N_49814,N_49698);
xnor UO_3235 (O_3235,N_42172,N_41444);
or UO_3236 (O_3236,N_45340,N_44551);
or UO_3237 (O_3237,N_49577,N_49965);
or UO_3238 (O_3238,N_42589,N_42597);
nor UO_3239 (O_3239,N_49937,N_47059);
or UO_3240 (O_3240,N_48140,N_40636);
or UO_3241 (O_3241,N_45593,N_48173);
and UO_3242 (O_3242,N_42978,N_42947);
or UO_3243 (O_3243,N_47557,N_49929);
and UO_3244 (O_3244,N_45591,N_48038);
nor UO_3245 (O_3245,N_45495,N_48603);
xor UO_3246 (O_3246,N_40201,N_40732);
xnor UO_3247 (O_3247,N_43879,N_46767);
nand UO_3248 (O_3248,N_48008,N_45686);
and UO_3249 (O_3249,N_42626,N_41822);
and UO_3250 (O_3250,N_41596,N_48690);
or UO_3251 (O_3251,N_40057,N_41072);
or UO_3252 (O_3252,N_43871,N_45383);
nand UO_3253 (O_3253,N_49927,N_49928);
nand UO_3254 (O_3254,N_42868,N_42596);
nand UO_3255 (O_3255,N_49289,N_45223);
nand UO_3256 (O_3256,N_45065,N_41152);
nor UO_3257 (O_3257,N_49344,N_44484);
and UO_3258 (O_3258,N_44691,N_41997);
nand UO_3259 (O_3259,N_41451,N_49383);
nor UO_3260 (O_3260,N_48321,N_46564);
or UO_3261 (O_3261,N_48212,N_42405);
or UO_3262 (O_3262,N_40995,N_47393);
and UO_3263 (O_3263,N_40867,N_49268);
and UO_3264 (O_3264,N_44601,N_44105);
or UO_3265 (O_3265,N_41962,N_45762);
xnor UO_3266 (O_3266,N_47729,N_45020);
nand UO_3267 (O_3267,N_41880,N_49829);
nor UO_3268 (O_3268,N_44398,N_40683);
and UO_3269 (O_3269,N_44791,N_44982);
xnor UO_3270 (O_3270,N_46805,N_48203);
nand UO_3271 (O_3271,N_47726,N_45994);
or UO_3272 (O_3272,N_48248,N_44658);
nor UO_3273 (O_3273,N_44502,N_47358);
and UO_3274 (O_3274,N_44688,N_44725);
nor UO_3275 (O_3275,N_46086,N_46730);
or UO_3276 (O_3276,N_48353,N_44418);
or UO_3277 (O_3277,N_42897,N_40160);
and UO_3278 (O_3278,N_42321,N_44152);
nand UO_3279 (O_3279,N_44656,N_45566);
and UO_3280 (O_3280,N_43112,N_47499);
and UO_3281 (O_3281,N_44096,N_43610);
nor UO_3282 (O_3282,N_42801,N_40413);
or UO_3283 (O_3283,N_45110,N_44843);
nand UO_3284 (O_3284,N_46829,N_42454);
or UO_3285 (O_3285,N_43412,N_40501);
nand UO_3286 (O_3286,N_40912,N_46001);
nor UO_3287 (O_3287,N_41016,N_46175);
nand UO_3288 (O_3288,N_41531,N_47152);
nand UO_3289 (O_3289,N_45862,N_44646);
and UO_3290 (O_3290,N_48701,N_48084);
nand UO_3291 (O_3291,N_40526,N_46542);
nand UO_3292 (O_3292,N_42176,N_48777);
or UO_3293 (O_3293,N_43795,N_48544);
and UO_3294 (O_3294,N_43415,N_49118);
and UO_3295 (O_3295,N_48747,N_47252);
and UO_3296 (O_3296,N_45296,N_41340);
nand UO_3297 (O_3297,N_44629,N_46376);
or UO_3298 (O_3298,N_41207,N_47816);
xor UO_3299 (O_3299,N_42899,N_46183);
nand UO_3300 (O_3300,N_48909,N_48920);
nor UO_3301 (O_3301,N_49359,N_49710);
and UO_3302 (O_3302,N_42668,N_41984);
nand UO_3303 (O_3303,N_48336,N_42246);
or UO_3304 (O_3304,N_40756,N_41258);
and UO_3305 (O_3305,N_46967,N_44211);
and UO_3306 (O_3306,N_47996,N_47511);
xnor UO_3307 (O_3307,N_47042,N_41157);
xor UO_3308 (O_3308,N_48645,N_40073);
or UO_3309 (O_3309,N_45682,N_47424);
nand UO_3310 (O_3310,N_40426,N_45992);
nor UO_3311 (O_3311,N_48752,N_49247);
or UO_3312 (O_3312,N_40657,N_46642);
and UO_3313 (O_3313,N_44222,N_40091);
nand UO_3314 (O_3314,N_45811,N_44128);
or UO_3315 (O_3315,N_48394,N_47801);
nor UO_3316 (O_3316,N_44209,N_49575);
xor UO_3317 (O_3317,N_48056,N_49988);
and UO_3318 (O_3318,N_48963,N_47552);
or UO_3319 (O_3319,N_45823,N_49197);
or UO_3320 (O_3320,N_49476,N_44234);
nand UO_3321 (O_3321,N_49909,N_49343);
nand UO_3322 (O_3322,N_41674,N_44397);
nor UO_3323 (O_3323,N_44413,N_42226);
and UO_3324 (O_3324,N_48784,N_42672);
or UO_3325 (O_3325,N_48416,N_47945);
or UO_3326 (O_3326,N_41036,N_42929);
nand UO_3327 (O_3327,N_40343,N_42220);
or UO_3328 (O_3328,N_44134,N_44937);
nand UO_3329 (O_3329,N_43735,N_40723);
xnor UO_3330 (O_3330,N_42281,N_49501);
and UO_3331 (O_3331,N_41413,N_43090);
xor UO_3332 (O_3332,N_44568,N_44547);
nand UO_3333 (O_3333,N_48671,N_48925);
xnor UO_3334 (O_3334,N_43154,N_45213);
and UO_3335 (O_3335,N_47827,N_47789);
nand UO_3336 (O_3336,N_48803,N_40466);
and UO_3337 (O_3337,N_46559,N_46724);
and UO_3338 (O_3338,N_45661,N_41970);
nand UO_3339 (O_3339,N_44935,N_48120);
nor UO_3340 (O_3340,N_42510,N_42453);
nand UO_3341 (O_3341,N_48221,N_42900);
nand UO_3342 (O_3342,N_40820,N_41271);
xnor UO_3343 (O_3343,N_44194,N_42326);
nand UO_3344 (O_3344,N_46857,N_47489);
nand UO_3345 (O_3345,N_49766,N_43142);
or UO_3346 (O_3346,N_47437,N_44495);
nand UO_3347 (O_3347,N_48379,N_42785);
and UO_3348 (O_3348,N_46949,N_40224);
or UO_3349 (O_3349,N_43890,N_49612);
or UO_3350 (O_3350,N_49508,N_47018);
nand UO_3351 (O_3351,N_47243,N_46207);
and UO_3352 (O_3352,N_44300,N_46121);
or UO_3353 (O_3353,N_40288,N_43324);
or UO_3354 (O_3354,N_41534,N_42450);
nor UO_3355 (O_3355,N_43147,N_46018);
nor UO_3356 (O_3356,N_42784,N_49137);
and UO_3357 (O_3357,N_43750,N_46437);
nor UO_3358 (O_3358,N_44400,N_48465);
or UO_3359 (O_3359,N_49354,N_48966);
nand UO_3360 (O_3360,N_46584,N_45096);
or UO_3361 (O_3361,N_45372,N_49973);
and UO_3362 (O_3362,N_48101,N_43553);
nand UO_3363 (O_3363,N_49522,N_46197);
and UO_3364 (O_3364,N_44701,N_40704);
nor UO_3365 (O_3365,N_47764,N_43746);
or UO_3366 (O_3366,N_48952,N_49427);
xor UO_3367 (O_3367,N_42185,N_49617);
nand UO_3368 (O_3368,N_47373,N_43885);
and UO_3369 (O_3369,N_41926,N_40890);
or UO_3370 (O_3370,N_45258,N_44343);
or UO_3371 (O_3371,N_40610,N_47625);
nand UO_3372 (O_3372,N_40480,N_42309);
and UO_3373 (O_3373,N_43625,N_42882);
or UO_3374 (O_3374,N_43984,N_49726);
or UO_3375 (O_3375,N_49261,N_48538);
or UO_3376 (O_3376,N_43511,N_41535);
nand UO_3377 (O_3377,N_45806,N_41556);
nor UO_3378 (O_3378,N_49639,N_42546);
or UO_3379 (O_3379,N_42367,N_46580);
nor UO_3380 (O_3380,N_40364,N_41752);
nand UO_3381 (O_3381,N_41440,N_44181);
nand UO_3382 (O_3382,N_46492,N_43808);
and UO_3383 (O_3383,N_44915,N_42928);
nand UO_3384 (O_3384,N_45601,N_47119);
or UO_3385 (O_3385,N_46239,N_42270);
and UO_3386 (O_3386,N_46173,N_40850);
nor UO_3387 (O_3387,N_46236,N_48131);
and UO_3388 (O_3388,N_47438,N_41069);
and UO_3389 (O_3389,N_43578,N_43650);
and UO_3390 (O_3390,N_40435,N_41416);
and UO_3391 (O_3391,N_41273,N_44845);
or UO_3392 (O_3392,N_45554,N_46331);
nor UO_3393 (O_3393,N_47829,N_42038);
and UO_3394 (O_3394,N_46388,N_42592);
xor UO_3395 (O_3395,N_47372,N_44584);
and UO_3396 (O_3396,N_48115,N_49228);
and UO_3397 (O_3397,N_48810,N_42224);
and UO_3398 (O_3398,N_42237,N_45402);
nand UO_3399 (O_3399,N_41726,N_44035);
nand UO_3400 (O_3400,N_45269,N_46384);
or UO_3401 (O_3401,N_46353,N_49827);
and UO_3402 (O_3402,N_45965,N_44809);
nand UO_3403 (O_3403,N_43644,N_48181);
or UO_3404 (O_3404,N_40047,N_45002);
nor UO_3405 (O_3405,N_42516,N_43363);
nor UO_3406 (O_3406,N_49771,N_42190);
or UO_3407 (O_3407,N_41232,N_41729);
nor UO_3408 (O_3408,N_41093,N_48577);
and UO_3409 (O_3409,N_44408,N_47658);
nand UO_3410 (O_3410,N_45146,N_46792);
or UO_3411 (O_3411,N_42208,N_47747);
xnor UO_3412 (O_3412,N_45136,N_44120);
nor UO_3413 (O_3413,N_48611,N_49181);
nor UO_3414 (O_3414,N_47291,N_41057);
or UO_3415 (O_3415,N_43442,N_49188);
and UO_3416 (O_3416,N_48775,N_45210);
nand UO_3417 (O_3417,N_47121,N_49578);
or UO_3418 (O_3418,N_49623,N_42023);
and UO_3419 (O_3419,N_42475,N_47314);
or UO_3420 (O_3420,N_41737,N_40392);
nand UO_3421 (O_3421,N_46235,N_43651);
nor UO_3422 (O_3422,N_46983,N_43304);
nor UO_3423 (O_3423,N_49871,N_40184);
nor UO_3424 (O_3424,N_43870,N_44410);
or UO_3425 (O_3425,N_42179,N_45270);
nor UO_3426 (O_3426,N_44206,N_48551);
or UO_3427 (O_3427,N_47147,N_46716);
or UO_3428 (O_3428,N_46494,N_48426);
or UO_3429 (O_3429,N_47369,N_43604);
nand UO_3430 (O_3430,N_43390,N_43691);
nand UO_3431 (O_3431,N_44715,N_44733);
nor UO_3432 (O_3432,N_47346,N_46741);
nor UO_3433 (O_3433,N_40670,N_45677);
or UO_3434 (O_3434,N_43387,N_46597);
or UO_3435 (O_3435,N_43523,N_40175);
and UO_3436 (O_3436,N_45217,N_46818);
nor UO_3437 (O_3437,N_48129,N_44165);
nor UO_3438 (O_3438,N_48409,N_43036);
nor UO_3439 (O_3439,N_48072,N_41329);
and UO_3440 (O_3440,N_43136,N_40496);
and UO_3441 (O_3441,N_48122,N_44116);
and UO_3442 (O_3442,N_46038,N_49417);
nand UO_3443 (O_3443,N_42698,N_47135);
and UO_3444 (O_3444,N_43942,N_49430);
and UO_3445 (O_3445,N_45790,N_47951);
and UO_3446 (O_3446,N_46095,N_47535);
and UO_3447 (O_3447,N_49235,N_46598);
nor UO_3448 (O_3448,N_42168,N_43404);
nand UO_3449 (O_3449,N_47757,N_42395);
and UO_3450 (O_3450,N_46051,N_43649);
and UO_3451 (O_3451,N_45470,N_48768);
nor UO_3452 (O_3452,N_46244,N_48932);
xnor UO_3453 (O_3453,N_45147,N_41750);
or UO_3454 (O_3454,N_49010,N_40524);
nand UO_3455 (O_3455,N_48754,N_44240);
nand UO_3456 (O_3456,N_49596,N_49139);
or UO_3457 (O_3457,N_41877,N_47985);
nand UO_3458 (O_3458,N_47621,N_49512);
and UO_3459 (O_3459,N_48324,N_45112);
and UO_3460 (O_3460,N_43450,N_49089);
nand UO_3461 (O_3461,N_45254,N_45511);
nand UO_3462 (O_3462,N_49498,N_47885);
nor UO_3463 (O_3463,N_43325,N_43945);
xor UO_3464 (O_3464,N_47195,N_45265);
and UO_3465 (O_3465,N_49158,N_45489);
xor UO_3466 (O_3466,N_46233,N_46449);
nor UO_3467 (O_3467,N_47936,N_40517);
nand UO_3468 (O_3468,N_42426,N_48570);
xnor UO_3469 (O_3469,N_49799,N_46509);
or UO_3470 (O_3470,N_42841,N_42802);
or UO_3471 (O_3471,N_43631,N_47226);
nor UO_3472 (O_3472,N_46200,N_47964);
nand UO_3473 (O_3473,N_41805,N_42722);
and UO_3474 (O_3474,N_46432,N_49939);
nor UO_3475 (O_3475,N_48274,N_40287);
nand UO_3476 (O_3476,N_46838,N_45141);
nor UO_3477 (O_3477,N_48972,N_47723);
or UO_3478 (O_3478,N_43343,N_40695);
nor UO_3479 (O_3479,N_43251,N_45899);
nand UO_3480 (O_3480,N_48498,N_40497);
or UO_3481 (O_3481,N_41540,N_40293);
or UO_3482 (O_3482,N_44003,N_45382);
or UO_3483 (O_3483,N_46641,N_47763);
xnor UO_3484 (O_3484,N_41253,N_46576);
and UO_3485 (O_3485,N_48535,N_47553);
or UO_3486 (O_3486,N_48087,N_40272);
and UO_3487 (O_3487,N_49493,N_43075);
or UO_3488 (O_3488,N_42213,N_42443);
and UO_3489 (O_3489,N_48177,N_49043);
nor UO_3490 (O_3490,N_43405,N_45821);
nand UO_3491 (O_3491,N_47307,N_43134);
nor UO_3492 (O_3492,N_42102,N_43223);
and UO_3493 (O_3493,N_41558,N_43498);
and UO_3494 (O_3494,N_48958,N_47087);
or UO_3495 (O_3495,N_41487,N_46136);
or UO_3496 (O_3496,N_47313,N_43029);
xnor UO_3497 (O_3497,N_49002,N_43013);
nand UO_3498 (O_3498,N_40417,N_42878);
or UO_3499 (O_3499,N_46033,N_48205);
nor UO_3500 (O_3500,N_48208,N_42275);
xnor UO_3501 (O_3501,N_47537,N_40998);
nand UO_3502 (O_3502,N_48300,N_42659);
or UO_3503 (O_3503,N_40362,N_49420);
or UO_3504 (O_3504,N_41600,N_48412);
and UO_3505 (O_3505,N_48640,N_45388);
nand UO_3506 (O_3506,N_42476,N_44832);
or UO_3507 (O_3507,N_42364,N_41102);
nor UO_3508 (O_3508,N_43038,N_46644);
nand UO_3509 (O_3509,N_41818,N_49712);
and UO_3510 (O_3510,N_46329,N_47882);
nor UO_3511 (O_3511,N_42957,N_45555);
and UO_3512 (O_3512,N_47886,N_48905);
nor UO_3513 (O_3513,N_47281,N_43845);
nor UO_3514 (O_3514,N_46573,N_44423);
nand UO_3515 (O_3515,N_40335,N_40893);
or UO_3516 (O_3516,N_41138,N_48051);
and UO_3517 (O_3517,N_41806,N_44769);
nor UO_3518 (O_3518,N_47528,N_44355);
and UO_3519 (O_3519,N_41866,N_42548);
nor UO_3520 (O_3520,N_48389,N_46370);
nor UO_3521 (O_3521,N_43078,N_40106);
xnor UO_3522 (O_3522,N_44468,N_43812);
and UO_3523 (O_3523,N_41265,N_47264);
and UO_3524 (O_3524,N_47876,N_47009);
and UO_3525 (O_3525,N_47690,N_41967);
nor UO_3526 (O_3526,N_44621,N_40722);
or UO_3527 (O_3527,N_40629,N_49631);
nand UO_3528 (O_3528,N_43165,N_42142);
nand UO_3529 (O_3529,N_40763,N_45035);
and UO_3530 (O_3530,N_47548,N_48862);
nand UO_3531 (O_3531,N_40785,N_44010);
nand UO_3532 (O_3532,N_45557,N_45174);
nand UO_3533 (O_3533,N_49415,N_47163);
nand UO_3534 (O_3534,N_49044,N_40875);
or UO_3535 (O_3535,N_46486,N_44006);
and UO_3536 (O_3536,N_40100,N_40598);
nand UO_3537 (O_3537,N_40765,N_48066);
or UO_3538 (O_3538,N_43860,N_47639);
nand UO_3539 (O_3539,N_43504,N_49409);
nand UO_3540 (O_3540,N_49178,N_45060);
nand UO_3541 (O_3541,N_41160,N_44838);
nand UO_3542 (O_3542,N_44946,N_48320);
nand UO_3543 (O_3543,N_49825,N_42982);
and UO_3544 (O_3544,N_46140,N_42707);
and UO_3545 (O_3545,N_41313,N_43084);
and UO_3546 (O_3546,N_43409,N_40975);
nor UO_3547 (O_3547,N_40398,N_41161);
nor UO_3548 (O_3548,N_49921,N_40711);
nand UO_3549 (O_3549,N_41976,N_46094);
or UO_3550 (O_3550,N_43548,N_40794);
or UO_3551 (O_3551,N_45527,N_49587);
or UO_3552 (O_3552,N_41318,N_40829);
nor UO_3553 (O_3553,N_48245,N_41011);
nor UO_3554 (O_3554,N_40382,N_41020);
or UO_3555 (O_3555,N_43476,N_41925);
nor UO_3556 (O_3556,N_44197,N_49436);
nor UO_3557 (O_3557,N_43121,N_49277);
and UO_3558 (O_3558,N_44974,N_46930);
nand UO_3559 (O_3559,N_47977,N_43377);
or UO_3560 (O_3560,N_40252,N_42838);
nor UO_3561 (O_3561,N_41014,N_45413);
nor UO_3562 (O_3562,N_48020,N_44292);
nand UO_3563 (O_3563,N_41747,N_48419);
nand UO_3564 (O_3564,N_45556,N_46536);
nand UO_3565 (O_3565,N_40673,N_49945);
nand UO_3566 (O_3566,N_45183,N_40839);
nor UO_3567 (O_3567,N_44327,N_43563);
or UO_3568 (O_3568,N_49877,N_43822);
nor UO_3569 (O_3569,N_41279,N_45375);
nor UO_3570 (O_3570,N_40903,N_45369);
nor UO_3571 (O_3571,N_45130,N_49781);
and UO_3572 (O_3572,N_45027,N_41909);
nor UO_3573 (O_3573,N_46989,N_40429);
nor UO_3574 (O_3574,N_43529,N_41283);
and UO_3575 (O_3575,N_44823,N_44052);
xor UO_3576 (O_3576,N_43654,N_40411);
xnor UO_3577 (O_3577,N_42890,N_43127);
nor UO_3578 (O_3578,N_41589,N_44157);
nor UO_3579 (O_3579,N_46616,N_44481);
and UO_3580 (O_3580,N_40075,N_40869);
or UO_3581 (O_3581,N_41103,N_49918);
and UO_3582 (O_3582,N_44195,N_43341);
nor UO_3583 (O_3583,N_45262,N_46219);
nor UO_3584 (O_3584,N_46548,N_45895);
nand UO_3585 (O_3585,N_48113,N_47810);
xor UO_3586 (O_3586,N_47268,N_41081);
or UO_3587 (O_3587,N_48918,N_47215);
and UO_3588 (O_3588,N_43923,N_49275);
and UO_3589 (O_3589,N_47348,N_49374);
or UO_3590 (O_3590,N_46715,N_40571);
nand UO_3591 (O_3591,N_46911,N_44660);
nand UO_3592 (O_3592,N_43603,N_44878);
nand UO_3593 (O_3593,N_43569,N_48908);
and UO_3594 (O_3594,N_47094,N_45846);
or UO_3595 (O_3595,N_45322,N_48436);
and UO_3596 (O_3596,N_45237,N_49563);
and UO_3597 (O_3597,N_45497,N_41190);
nand UO_3598 (O_3598,N_49212,N_43889);
nor UO_3599 (O_3599,N_47315,N_40687);
nand UO_3600 (O_3600,N_41678,N_40739);
or UO_3601 (O_3601,N_44867,N_45084);
nor UO_3602 (O_3602,N_46704,N_48930);
nor UO_3603 (O_3603,N_45769,N_46012);
and UO_3604 (O_3604,N_43820,N_47253);
and UO_3605 (O_3605,N_48308,N_45745);
or UO_3606 (O_3606,N_42798,N_47990);
nand UO_3607 (O_3607,N_45171,N_46778);
nor UO_3608 (O_3608,N_47484,N_42043);
or UO_3609 (O_3609,N_41009,N_43235);
and UO_3610 (O_3610,N_41612,N_46453);
nand UO_3611 (O_3611,N_46473,N_49611);
nor UO_3612 (O_3612,N_48468,N_47330);
xor UO_3613 (O_3613,N_44908,N_46523);
nand UO_3614 (O_3614,N_44576,N_40793);
and UO_3615 (O_3615,N_43558,N_47355);
and UO_3616 (O_3616,N_48742,N_40454);
xor UO_3617 (O_3617,N_40388,N_41597);
xnor UO_3618 (O_3618,N_41856,N_47384);
nor UO_3619 (O_3619,N_49288,N_42863);
nand UO_3620 (O_3620,N_47308,N_43628);
or UO_3621 (O_3621,N_48755,N_48724);
nand UO_3622 (O_3622,N_47730,N_47374);
and UO_3623 (O_3623,N_47130,N_49195);
nand UO_3624 (O_3624,N_42418,N_48467);
xor UO_3625 (O_3625,N_46342,N_47027);
nand UO_3626 (O_3626,N_49987,N_44123);
xnor UO_3627 (O_3627,N_48649,N_42649);
or UO_3628 (O_3628,N_44368,N_47474);
or UO_3629 (O_3629,N_45675,N_46339);
or UO_3630 (O_3630,N_46100,N_41684);
nand UO_3631 (O_3631,N_43330,N_44857);
nand UO_3632 (O_3632,N_40742,N_45567);
nand UO_3633 (O_3633,N_48312,N_46524);
or UO_3634 (O_3634,N_49060,N_44607);
and UO_3635 (O_3635,N_41167,N_40701);
or UO_3636 (O_3636,N_41711,N_46977);
and UO_3637 (O_3637,N_47054,N_43679);
nand UO_3638 (O_3638,N_42433,N_42898);
or UO_3639 (O_3639,N_42169,N_45481);
or UO_3640 (O_3640,N_47020,N_46561);
nand UO_3641 (O_3641,N_47850,N_46825);
nor UO_3642 (O_3642,N_49880,N_46332);
nor UO_3643 (O_3643,N_46797,N_44987);
xnor UO_3644 (O_3644,N_40261,N_45582);
or UO_3645 (O_3645,N_49947,N_49320);
and UO_3646 (O_3646,N_40267,N_44278);
or UO_3647 (O_3647,N_43894,N_45144);
and UO_3648 (O_3648,N_49558,N_44174);
or UO_3649 (O_3649,N_45305,N_40264);
or UO_3650 (O_3650,N_48524,N_47874);
nor UO_3651 (O_3651,N_41094,N_49798);
xnor UO_3652 (O_3652,N_48559,N_42590);
nand UO_3653 (O_3653,N_49893,N_47000);
nand UO_3654 (O_3654,N_46277,N_46021);
nor UO_3655 (O_3655,N_49724,N_44196);
and UO_3656 (O_3656,N_42790,N_43352);
nand UO_3657 (O_3657,N_42413,N_47249);
nand UO_3658 (O_3658,N_40438,N_44899);
nand UO_3659 (O_3659,N_47402,N_43832);
xor UO_3660 (O_3660,N_43275,N_49290);
nor UO_3661 (O_3661,N_40180,N_41326);
and UO_3662 (O_3662,N_43086,N_42130);
nor UO_3663 (O_3663,N_43231,N_45006);
and UO_3664 (O_3664,N_41031,N_48025);
and UO_3665 (O_3665,N_41362,N_44804);
xnor UO_3666 (O_3666,N_45343,N_48523);
and UO_3667 (O_3667,N_48138,N_44058);
nand UO_3668 (O_3668,N_47356,N_49747);
nand UO_3669 (O_3669,N_43867,N_44693);
nand UO_3670 (O_3670,N_49561,N_46574);
and UO_3671 (O_3671,N_49393,N_45394);
xor UO_3672 (O_3672,N_47661,N_45898);
nand UO_3673 (O_3673,N_46723,N_41194);
nor UO_3674 (O_3674,N_46142,N_49536);
nor UO_3675 (O_3675,N_40522,N_43313);
and UO_3676 (O_3676,N_46004,N_45761);
nor UO_3677 (O_3677,N_45902,N_43738);
and UO_3678 (O_3678,N_47532,N_48150);
or UO_3679 (O_3679,N_45428,N_48787);
and UO_3680 (O_3680,N_49363,N_49183);
nor UO_3681 (O_3681,N_45212,N_46184);
xnor UO_3682 (O_3682,N_44651,N_44759);
nor UO_3683 (O_3683,N_43105,N_48686);
and UO_3684 (O_3684,N_44022,N_42087);
nand UO_3685 (O_3685,N_49206,N_45804);
or UO_3686 (O_3686,N_43737,N_47814);
nor UO_3687 (O_3687,N_46885,N_41382);
or UO_3688 (O_3688,N_40955,N_40748);
nor UO_3689 (O_3689,N_41604,N_48194);
xnor UO_3690 (O_3690,N_41331,N_41248);
nand UO_3691 (O_3691,N_48364,N_42817);
and UO_3692 (O_3692,N_43243,N_43101);
nor UO_3693 (O_3693,N_47104,N_43310);
or UO_3694 (O_3694,N_49709,N_43028);
or UO_3695 (O_3695,N_41381,N_40562);
or UO_3696 (O_3696,N_41284,N_40179);
nor UO_3697 (O_3697,N_49477,N_42969);
and UO_3698 (O_3698,N_48222,N_42156);
and UO_3699 (O_3699,N_42823,N_45290);
and UO_3700 (O_3700,N_49063,N_47636);
or UO_3701 (O_3701,N_48534,N_41098);
xor UO_3702 (O_3702,N_42466,N_45779);
nor UO_3703 (O_3703,N_45887,N_49398);
and UO_3704 (O_3704,N_49588,N_40560);
or UO_3705 (O_3705,N_43359,N_44169);
or UO_3706 (O_3706,N_41513,N_43099);
nor UO_3707 (O_3707,N_41927,N_48833);
nand UO_3708 (O_3708,N_43218,N_48352);
xnor UO_3709 (O_3709,N_40712,N_49807);
or UO_3710 (O_3710,N_42403,N_47732);
nor UO_3711 (O_3711,N_45251,N_48244);
nor UO_3712 (O_3712,N_48767,N_41263);
nand UO_3713 (O_3713,N_48258,N_48356);
nand UO_3714 (O_3714,N_40647,N_48216);
nor UO_3715 (O_3715,N_40018,N_41736);
nand UO_3716 (O_3716,N_46648,N_44445);
nor UO_3717 (O_3717,N_42348,N_47501);
nor UO_3718 (O_3718,N_44522,N_47407);
or UO_3719 (O_3719,N_49900,N_42635);
and UO_3720 (O_3720,N_44275,N_45483);
or UO_3721 (O_3721,N_40046,N_44306);
nand UO_3722 (O_3722,N_43505,N_43371);
nor UO_3723 (O_3723,N_45793,N_40221);
nor UO_3724 (O_3724,N_40108,N_49532);
xnor UO_3725 (O_3725,N_47405,N_44382);
and UO_3726 (O_3726,N_44711,N_45974);
nand UO_3727 (O_3727,N_45574,N_46659);
and UO_3728 (O_3728,N_48697,N_48369);
or UO_3729 (O_3729,N_41553,N_40263);
nand UO_3730 (O_3730,N_46990,N_48477);
and UO_3731 (O_3731,N_49076,N_48383);
nand UO_3732 (O_3732,N_49553,N_44657);
nor UO_3733 (O_3733,N_46572,N_45587);
nor UO_3734 (O_3734,N_43816,N_44650);
nand UO_3735 (O_3735,N_46313,N_41999);
or UO_3736 (O_3736,N_43089,N_47327);
and UO_3737 (O_3737,N_40478,N_40508);
nand UO_3738 (O_3738,N_40539,N_43519);
and UO_3739 (O_3739,N_48086,N_40305);
nor UO_3740 (O_3740,N_48034,N_43760);
or UO_3741 (O_3741,N_45326,N_40483);
or UO_3742 (O_3742,N_48501,N_43844);
xnor UO_3743 (O_3743,N_42474,N_47190);
nor UO_3744 (O_3744,N_41512,N_48801);
or UO_3745 (O_3745,N_42473,N_47299);
xnor UO_3746 (O_3746,N_47583,N_47618);
and UO_3747 (O_3747,N_43179,N_48680);
nor UO_3748 (O_3748,N_49170,N_48322);
nor UO_3749 (O_3749,N_48284,N_44521);
nand UO_3750 (O_3750,N_43898,N_49369);
and UO_3751 (O_3751,N_43601,N_44467);
and UO_3752 (O_3752,N_45129,N_42158);
nor UO_3753 (O_3753,N_44039,N_42357);
nor UO_3754 (O_3754,N_49514,N_49733);
nand UO_3755 (O_3755,N_42642,N_44684);
and UO_3756 (O_3756,N_49635,N_47686);
nor UO_3757 (O_3757,N_48831,N_43534);
and UO_3758 (O_3758,N_43345,N_43500);
nor UO_3759 (O_3759,N_49160,N_46290);
nor UO_3760 (O_3760,N_47278,N_48340);
nand UO_3761 (O_3761,N_40176,N_47211);
xnor UO_3762 (O_3762,N_42105,N_44441);
and UO_3763 (O_3763,N_48376,N_44549);
and UO_3764 (O_3764,N_46804,N_43761);
and UO_3765 (O_3765,N_45611,N_49102);
nand UO_3766 (O_3766,N_43635,N_40865);
nor UO_3767 (O_3767,N_45864,N_41649);
nand UO_3768 (O_3768,N_43502,N_41438);
nand UO_3769 (O_3769,N_42409,N_47472);
nor UO_3770 (O_3770,N_41117,N_49120);
nor UO_3771 (O_3771,N_49953,N_41492);
or UO_3772 (O_3772,N_42631,N_49738);
nor UO_3773 (O_3773,N_49479,N_44784);
xnor UO_3774 (O_3774,N_49497,N_43278);
xor UO_3775 (O_3775,N_42712,N_46808);
and UO_3776 (O_3776,N_45487,N_45602);
nor UO_3777 (O_3777,N_41480,N_42171);
nor UO_3778 (O_3778,N_49584,N_44238);
xor UO_3779 (O_3779,N_46618,N_46396);
xnor UO_3780 (O_3780,N_46471,N_49349);
nor UO_3781 (O_3781,N_44364,N_40814);
or UO_3782 (O_3782,N_46460,N_49088);
and UO_3783 (O_3783,N_47401,N_43140);
and UO_3784 (O_3784,N_47578,N_41618);
or UO_3785 (O_3785,N_48760,N_41490);
and UO_3786 (O_3786,N_40316,N_41617);
xnor UO_3787 (O_3787,N_47762,N_43394);
nor UO_3788 (O_3788,N_49521,N_42870);
nand UO_3789 (O_3789,N_40710,N_44542);
nor UO_3790 (O_3790,N_43886,N_43787);
and UO_3791 (O_3791,N_41797,N_47644);
and UO_3792 (O_3792,N_40450,N_45341);
nor UO_3793 (O_3793,N_43033,N_46918);
and UO_3794 (O_3794,N_45001,N_42351);
and UO_3795 (O_3795,N_45429,N_41299);
nor UO_3796 (O_3796,N_43484,N_43872);
nand UO_3797 (O_3797,N_43002,N_45639);
nor UO_3798 (O_3798,N_47478,N_47536);
or UO_3799 (O_3799,N_46034,N_44390);
nand UO_3800 (O_3800,N_47336,N_41266);
nor UO_3801 (O_3801,N_42167,N_40766);
nor UO_3802 (O_3802,N_45755,N_43207);
xnor UO_3803 (O_3803,N_44284,N_41666);
and UO_3804 (O_3804,N_42323,N_41089);
nor UO_3805 (O_3805,N_47620,N_41353);
nand UO_3806 (O_3806,N_45316,N_40708);
and UO_3807 (O_3807,N_45757,N_42795);
or UO_3808 (O_3808,N_47158,N_48917);
xnor UO_3809 (O_3809,N_42953,N_49625);
xnor UO_3810 (O_3810,N_42007,N_48510);
or UO_3811 (O_3811,N_41024,N_42336);
nand UO_3812 (O_3812,N_46557,N_43264);
nand UO_3813 (O_3813,N_44344,N_40042);
or UO_3814 (O_3814,N_43721,N_44188);
xor UO_3815 (O_3815,N_47023,N_43232);
xnor UO_3816 (O_3816,N_46134,N_43788);
or UO_3817 (O_3817,N_42202,N_47607);
nand UO_3818 (O_3818,N_42315,N_46781);
nand UO_3819 (O_3819,N_41297,N_44632);
and UO_3820 (O_3820,N_40721,N_44582);
and UO_3821 (O_3821,N_48105,N_49526);
and UO_3822 (O_3822,N_43912,N_46993);
and UO_3823 (O_3823,N_49863,N_42562);
and UO_3824 (O_3824,N_48180,N_42244);
xor UO_3825 (O_3825,N_46553,N_47486);
xnor UO_3826 (O_3826,N_44569,N_45458);
nor UO_3827 (O_3827,N_46954,N_47049);
nor UO_3828 (O_3828,N_48446,N_49716);
nand UO_3829 (O_3829,N_45533,N_48984);
and UO_3830 (O_3830,N_43108,N_40414);
nor UO_3831 (O_3831,N_41327,N_49452);
nand UO_3832 (O_3832,N_41421,N_40188);
nor UO_3833 (O_3833,N_47828,N_43546);
nand UO_3834 (O_3834,N_45538,N_49816);
nor UO_3835 (O_3835,N_43995,N_45692);
nor UO_3836 (O_3836,N_45358,N_46023);
nor UO_3837 (O_3837,N_46593,N_45252);
nor UO_3838 (O_3838,N_47697,N_45698);
xor UO_3839 (O_3839,N_41727,N_42667);
and UO_3840 (O_3840,N_40534,N_46250);
and UO_3841 (O_3841,N_43850,N_43408);
and UO_3842 (O_3842,N_42906,N_44768);
or UO_3843 (O_3843,N_43293,N_48689);
nand UO_3844 (O_3844,N_46728,N_40090);
nor UO_3845 (O_3845,N_44805,N_42469);
or UO_3846 (O_3846,N_40098,N_48236);
nand UO_3847 (O_3847,N_48638,N_49729);
xor UO_3848 (O_3848,N_42645,N_40370);
xnor UO_3849 (O_3849,N_40770,N_47733);
or UO_3850 (O_3850,N_44994,N_46368);
nand UO_3851 (O_3851,N_45439,N_40400);
nand UO_3852 (O_3852,N_46068,N_49821);
nand UO_3853 (O_3853,N_42752,N_42427);
and UO_3854 (O_3854,N_42803,N_48001);
or UO_3855 (O_3855,N_40044,N_40549);
and UO_3856 (O_3856,N_42770,N_49714);
nand UO_3857 (O_3857,N_41245,N_43263);
nor UO_3858 (O_3858,N_48488,N_49171);
nand UO_3859 (O_3859,N_47900,N_49111);
nor UO_3860 (O_3860,N_44962,N_48028);
nor UO_3861 (O_3861,N_43460,N_40096);
nand UO_3862 (O_3862,N_48197,N_46615);
and UO_3863 (O_3863,N_49672,N_46827);
and UO_3864 (O_3864,N_44512,N_43714);
nor UO_3865 (O_3865,N_43395,N_46014);
and UO_3866 (O_3866,N_47906,N_48881);
or UO_3867 (O_3867,N_42261,N_45673);
nor UO_3868 (O_3868,N_42941,N_47703);
nor UO_3869 (O_3869,N_42338,N_49861);
and UO_3870 (O_3870,N_41048,N_46213);
nand UO_3871 (O_3871,N_40802,N_40380);
or UO_3872 (O_3872,N_42262,N_48741);
or UO_3873 (O_3873,N_47716,N_49801);
and UO_3874 (O_3874,N_40071,N_41817);
nor UO_3875 (O_3875,N_43447,N_45445);
and UO_3876 (O_3876,N_49889,N_41002);
nand UO_3877 (O_3877,N_49668,N_45603);
or UO_3878 (O_3878,N_44509,N_49046);
or UO_3879 (O_3879,N_42855,N_43909);
or UO_3880 (O_3880,N_46785,N_48637);
and UO_3881 (O_3881,N_40087,N_47573);
and UO_3882 (O_3882,N_44579,N_44726);
nor UO_3883 (O_3883,N_49202,N_43226);
or UO_3884 (O_3884,N_41559,N_48102);
or UO_3885 (O_3885,N_49750,N_46320);
or UO_3886 (O_3886,N_40326,N_46441);
or UO_3887 (O_3887,N_42621,N_48506);
nor UO_3888 (O_3888,N_49234,N_45393);
nor UO_3889 (O_3889,N_45260,N_45723);
nand UO_3890 (O_3890,N_40514,N_47782);
nand UO_3891 (O_3891,N_41638,N_43940);
nand UO_3892 (O_3892,N_48088,N_41307);
xor UO_3893 (O_3893,N_41860,N_40094);
and UO_3894 (O_3894,N_40755,N_44714);
xnor UO_3895 (O_3895,N_47460,N_43262);
and UO_3896 (O_3896,N_40294,N_48847);
and UO_3897 (O_3897,N_49260,N_40815);
xnor UO_3898 (O_3898,N_43197,N_45409);
and UO_3899 (O_3899,N_42804,N_43661);
nor UO_3900 (O_3900,N_41240,N_45870);
xnor UO_3901 (O_3901,N_46594,N_45033);
nor UO_3902 (O_3902,N_40535,N_48496);
nand UO_3903 (O_3903,N_48773,N_44357);
nor UO_3904 (O_3904,N_43615,N_47418);
xnor UO_3905 (O_3905,N_44242,N_42289);
nand UO_3906 (O_3906,N_49106,N_42076);
and UO_3907 (O_3907,N_44346,N_44101);
or UO_3908 (O_3908,N_47755,N_46426);
nand UO_3909 (O_3909,N_47458,N_47751);
or UO_3910 (O_3910,N_47752,N_43372);
xnor UO_3911 (O_3911,N_45885,N_41309);
and UO_3912 (O_3912,N_45256,N_48309);
or UO_3913 (O_3913,N_42025,N_44773);
nand UO_3914 (O_3914,N_44271,N_41304);
or UO_3915 (O_3915,N_40349,N_47099);
nand UO_3916 (O_3916,N_47932,N_41951);
and UO_3917 (O_3917,N_49761,N_41135);
nor UO_3918 (O_3918,N_46271,N_40209);
or UO_3919 (O_3919,N_42990,N_49506);
xnor UO_3920 (O_3920,N_42715,N_40807);
nor UO_3921 (O_3921,N_45695,N_47696);
nand UO_3922 (O_3922,N_45640,N_47225);
nand UO_3923 (O_3923,N_40322,N_43607);
and UO_3924 (O_3924,N_49440,N_44953);
or UO_3925 (O_3925,N_49769,N_45120);
nand UO_3926 (O_3926,N_43510,N_42447);
nor UO_3927 (O_3927,N_45879,N_46915);
or UO_3928 (O_3928,N_42264,N_41740);
nand UO_3929 (O_3929,N_47623,N_48160);
and UO_3930 (O_3930,N_48769,N_42815);
nor UO_3931 (O_3931,N_48944,N_49646);
or UO_3932 (O_3932,N_46468,N_40391);
xnor UO_3933 (O_3933,N_44897,N_45679);
or UO_3934 (O_3934,N_45187,N_47653);
or UO_3935 (O_3935,N_40005,N_40374);
nor UO_3936 (O_3936,N_47376,N_44699);
nand UO_3937 (O_3937,N_48272,N_45450);
nor UO_3938 (O_3938,N_43007,N_48147);
nor UO_3939 (O_3939,N_45854,N_43690);
xor UO_3940 (O_3940,N_47159,N_43230);
or UO_3941 (O_3941,N_47028,N_41681);
and UO_3942 (O_3942,N_44675,N_46273);
or UO_3943 (O_3943,N_42650,N_49978);
or UO_3944 (O_3944,N_47818,N_43982);
or UO_3945 (O_3945,N_43452,N_48330);
nand UO_3946 (O_3946,N_45190,N_44496);
nor UO_3947 (O_3947,N_48959,N_42077);
nand UO_3948 (O_3948,N_46839,N_40505);
and UO_3949 (O_3949,N_43133,N_48688);
nor UO_3950 (O_3950,N_46010,N_48043);
xor UO_3951 (O_3951,N_48075,N_48338);
and UO_3952 (O_3952,N_48727,N_49507);
and UO_3953 (O_3953,N_48711,N_49858);
and UO_3954 (O_3954,N_41237,N_41317);
and UO_3955 (O_3955,N_42052,N_40751);
nand UO_3956 (O_3956,N_41296,N_44687);
nor UO_3957 (O_3957,N_44356,N_47561);
nor UO_3958 (O_3958,N_40017,N_49310);
or UO_3959 (O_3959,N_49758,N_41034);
nand UO_3960 (O_3960,N_46114,N_46451);
or UO_3961 (O_3961,N_44620,N_43780);
and UO_3962 (O_3962,N_41940,N_45097);
nand UO_3963 (O_3963,N_46391,N_40196);
or UO_3964 (O_3964,N_47179,N_46048);
and UO_3965 (O_3965,N_49856,N_42099);
or UO_3966 (O_3966,N_44457,N_42633);
or UO_3967 (O_3967,N_44981,N_49049);
and UO_3968 (O_3968,N_41528,N_44047);
or UO_3969 (O_3969,N_41171,N_48821);
or UO_3970 (O_3970,N_44605,N_41682);
and UO_3971 (O_3971,N_42401,N_49238);
nand UO_3972 (O_3972,N_43418,N_46525);
or UO_3973 (O_3973,N_45031,N_41001);
xor UO_3974 (O_3974,N_45381,N_42006);
nor UO_3975 (O_3975,N_42316,N_45861);
nand UO_3976 (O_3976,N_46201,N_43114);
nor UO_3977 (O_3977,N_44472,N_40665);
or UO_3978 (O_3978,N_48290,N_42278);
nor UO_3979 (O_3979,N_43254,N_44446);
nand UO_3980 (O_3980,N_45596,N_44229);
nand UO_3981 (O_3981,N_47812,N_49728);
nor UO_3982 (O_3982,N_49552,N_41267);
or UO_3983 (O_3983,N_40110,N_49701);
and UO_3984 (O_3984,N_46020,N_48583);
and UO_3985 (O_3985,N_47368,N_42616);
or UO_3986 (O_3986,N_49348,N_43814);
nor UO_3987 (O_3987,N_45606,N_46903);
nand UO_3988 (O_3988,N_47858,N_40306);
or UO_3989 (O_3989,N_42731,N_42271);
nor UO_3990 (O_3990,N_44507,N_40375);
nor UO_3991 (O_3991,N_43193,N_44399);
and UO_3992 (O_3992,N_45520,N_48886);
xor UO_3993 (O_3993,N_47236,N_49213);
nand UO_3994 (O_3994,N_41607,N_43180);
nor UO_3995 (O_3995,N_44459,N_48307);
or UO_3996 (O_3996,N_44916,N_40579);
xor UO_3997 (O_3997,N_47298,N_43195);
and UO_3998 (O_3998,N_47220,N_46545);
and UO_3999 (O_3999,N_47637,N_40409);
xor UO_4000 (O_4000,N_47149,N_40758);
nor UO_4001 (O_4001,N_41557,N_48373);
xnor UO_4002 (O_4002,N_43096,N_49433);
nor UO_4003 (O_4003,N_45782,N_44674);
xnor UO_4004 (O_4004,N_49142,N_43730);
xnor UO_4005 (O_4005,N_44040,N_45801);
nand UO_4006 (O_4006,N_46442,N_41021);
nor UO_4007 (O_4007,N_41212,N_47871);
nor UO_4008 (O_4008,N_46653,N_42856);
nand UO_4009 (O_4009,N_45559,N_49058);
or UO_4010 (O_4010,N_47955,N_43606);
and UO_4011 (O_4011,N_45430,N_41789);
and UO_4012 (O_4012,N_46208,N_40443);
nand UO_4013 (O_4013,N_47284,N_48492);
or UO_4014 (O_4014,N_43514,N_47413);
nor UO_4015 (O_4015,N_46975,N_42332);
or UO_4016 (O_4016,N_48193,N_42230);
nor UO_4017 (O_4017,N_44696,N_45949);
nor UO_4018 (O_4018,N_45228,N_49190);
nand UO_4019 (O_4019,N_45038,N_47456);
or UO_4020 (O_4020,N_41292,N_47109);
or UO_4021 (O_4021,N_47194,N_46666);
nor UO_4022 (O_4022,N_43237,N_46727);
and UO_4023 (O_4023,N_42499,N_45700);
nor UO_4024 (O_4024,N_42624,N_43403);
or UO_4025 (O_4025,N_43989,N_44384);
and UO_4026 (O_4026,N_43466,N_44548);
or UO_4027 (O_4027,N_46874,N_46286);
nor UO_4028 (O_4028,N_49255,N_44966);
nand UO_4029 (O_4029,N_44068,N_41985);
and UO_4030 (O_4030,N_47881,N_40581);
nand UO_4031 (O_4031,N_49007,N_48059);
nand UO_4032 (O_4032,N_40377,N_47830);
and UO_4033 (O_4033,N_45535,N_45724);
nand UO_4034 (O_4034,N_47185,N_42708);
xor UO_4035 (O_4035,N_40139,N_43181);
nor UO_4036 (O_4036,N_44203,N_49148);
nand UO_4037 (O_4037,N_45563,N_43991);
nand UO_4038 (O_4038,N_45398,N_46268);
and UO_4039 (O_4039,N_43074,N_47172);
and UO_4040 (O_4040,N_46683,N_49358);
or UO_4041 (O_4041,N_47245,N_43319);
or UO_4042 (O_4042,N_42065,N_44252);
xor UO_4043 (O_4043,N_49492,N_44080);
nor UO_4044 (O_4044,N_47210,N_45412);
and UO_4045 (O_4045,N_44230,N_45189);
and UO_4046 (O_4046,N_49568,N_42000);
nor UO_4047 (O_4047,N_46872,N_48106);
and UO_4048 (O_4048,N_47475,N_46252);
or UO_4049 (O_4049,N_42772,N_45696);
and UO_4050 (O_4050,N_44541,N_48007);
or UO_4051 (O_4051,N_41564,N_47448);
nand UO_4052 (O_4052,N_41839,N_42311);
nor UO_4053 (O_4053,N_44280,N_40885);
and UO_4054 (O_4054,N_43106,N_49708);
or UO_4055 (O_4055,N_49986,N_40754);
nor UO_4056 (O_4056,N_49981,N_40963);
nand UO_4057 (O_4057,N_48283,N_49346);
or UO_4058 (O_4058,N_48202,N_41270);
nor UO_4059 (O_4059,N_49104,N_46029);
nor UO_4060 (O_4060,N_41361,N_46243);
and UO_4061 (O_4061,N_41507,N_45623);
nand UO_4062 (O_4062,N_47988,N_41676);
and UO_4063 (O_4063,N_45955,N_42425);
xor UO_4064 (O_4064,N_46256,N_48866);
or UO_4065 (O_4065,N_40938,N_43731);
or UO_4066 (O_4066,N_44647,N_42834);
nand UO_4067 (O_4067,N_47793,N_44416);
or UO_4068 (O_4068,N_42824,N_41610);
or UO_4069 (O_4069,N_41246,N_44562);
and UO_4070 (O_4070,N_44606,N_41845);
nand UO_4071 (O_4071,N_46844,N_44933);
nand UO_4072 (O_4072,N_49543,N_49303);
or UO_4073 (O_4073,N_48946,N_42284);
or UO_4074 (O_4074,N_47267,N_49074);
and UO_4075 (O_4075,N_46671,N_47131);
nor UO_4076 (O_4076,N_44274,N_41751);
nor UO_4077 (O_4077,N_49930,N_41043);
or UO_4078 (O_4078,N_48133,N_47453);
or UO_4079 (O_4079,N_41308,N_48555);
and UO_4080 (O_4080,N_40023,N_44391);
nor UO_4081 (O_4081,N_46934,N_41532);
or UO_4082 (O_4082,N_46280,N_45838);
nor UO_4083 (O_4083,N_41290,N_49599);
and UO_4084 (O_4084,N_48863,N_42279);
nand UO_4085 (O_4085,N_40329,N_40025);
nor UO_4086 (O_4086,N_46876,N_41702);
or UO_4087 (O_4087,N_42194,N_48061);
and UO_4088 (O_4088,N_45273,N_48661);
or UO_4089 (O_4089,N_42308,N_45287);
nand UO_4090 (O_4090,N_43046,N_48667);
or UO_4091 (O_4091,N_45945,N_45342);
and UO_4092 (O_4092,N_49546,N_46307);
or UO_4093 (O_4093,N_41987,N_44519);
and UO_4094 (O_4094,N_41178,N_47677);
nor UO_4095 (O_4095,N_40644,N_43219);
or UO_4096 (O_4096,N_49690,N_42472);
and UO_4097 (O_4097,N_49593,N_47254);
nand UO_4098 (O_4098,N_46152,N_49067);
nor UO_4099 (O_4099,N_40648,N_47761);
nand UO_4100 (O_4100,N_43189,N_41404);
nor UO_4101 (O_4101,N_44033,N_43458);
xnor UO_4102 (O_4102,N_46341,N_41330);
and UO_4103 (O_4103,N_43283,N_49620);
nor UO_4104 (O_4104,N_43483,N_41000);
nand UO_4105 (O_4105,N_44377,N_44322);
nand UO_4106 (O_4106,N_43931,N_42889);
or UO_4107 (O_4107,N_41142,N_45528);
or UO_4108 (O_4108,N_43030,N_47504);
and UO_4109 (O_4109,N_48995,N_45417);
or UO_4110 (O_4110,N_47041,N_44713);
and UO_4111 (O_4111,N_48532,N_49849);
xnor UO_4112 (O_4112,N_44432,N_41186);
nor UO_4113 (O_4113,N_46056,N_43240);
and UO_4114 (O_4114,N_46571,N_43385);
nor UO_4115 (O_4115,N_41708,N_43602);
xor UO_4116 (O_4116,N_48117,N_46795);
or UO_4117 (O_4117,N_42533,N_44789);
and UO_4118 (O_4118,N_47191,N_47774);
xor UO_4119 (O_4119,N_41659,N_47359);
nand UO_4120 (O_4120,N_47035,N_48176);
nand UO_4121 (O_4121,N_41760,N_49442);
and UO_4122 (O_4122,N_41431,N_41430);
or UO_4123 (O_4123,N_44753,N_44677);
nor UO_4124 (O_4124,N_48789,N_45913);
xnor UO_4125 (O_4125,N_48485,N_46555);
and UO_4126 (O_4126,N_49468,N_44210);
nand UO_4127 (O_4127,N_44479,N_44792);
or UO_4128 (O_4128,N_44248,N_46458);
nor UO_4129 (O_4129,N_46841,N_45318);
nor UO_4130 (O_4130,N_44494,N_49791);
or UO_4131 (O_4131,N_44458,N_47656);
nand UO_4132 (O_4132,N_44882,N_49891);
and UO_4133 (O_4133,N_42971,N_43039);
and UO_4134 (O_4134,N_40068,N_41346);
nor UO_4135 (O_4135,N_40270,N_40477);
nor UO_4136 (O_4136,N_43308,N_47260);
and UO_4137 (O_4137,N_41730,N_42389);
nor UO_4138 (O_4138,N_42600,N_40245);
or UO_4139 (O_4139,N_46498,N_43270);
and UO_4140 (O_4140,N_46397,N_43557);
and UO_4141 (O_4141,N_40891,N_47521);
nor UO_4142 (O_4142,N_45395,N_45613);
nand UO_4143 (O_4143,N_44751,N_43614);
and UO_4144 (O_4144,N_44808,N_49673);
and UO_4145 (O_4145,N_48721,N_44216);
nor UO_4146 (O_4146,N_44618,N_49322);
and UO_4147 (O_4147,N_43162,N_49072);
and UO_4148 (O_4148,N_44951,N_47275);
nand UO_4149 (O_4149,N_40323,N_43015);
nand UO_4150 (O_4150,N_43126,N_42932);
nand UO_4151 (O_4151,N_46757,N_45688);
nor UO_4152 (O_4152,N_47014,N_42959);
nand UO_4153 (O_4153,N_43874,N_46003);
xnor UO_4154 (O_4154,N_49449,N_49676);
or UO_4155 (O_4155,N_47026,N_41635);
nor UO_4156 (O_4156,N_44968,N_47540);
nor UO_4157 (O_4157,N_40191,N_44415);
xor UO_4158 (O_4158,N_46375,N_48044);
and UO_4159 (O_4159,N_44000,N_46180);
nand UO_4160 (O_4160,N_49720,N_47302);
nand UO_4161 (O_4161,N_44880,N_44821);
xor UO_4162 (O_4162,N_46162,N_45990);
and UO_4163 (O_4163,N_47958,N_44227);
nand UO_4164 (O_4164,N_44765,N_44608);
and UO_4165 (O_4165,N_44641,N_45777);
and UO_4166 (O_4166,N_41983,N_41504);
or UO_4167 (O_4167,N_47991,N_48904);
and UO_4168 (O_4168,N_45731,N_40493);
xor UO_4169 (O_4169,N_43985,N_49995);
nand UO_4170 (O_4170,N_42408,N_43759);
or UO_4171 (O_4171,N_45441,N_42468);
or UO_4172 (O_4172,N_40733,N_48192);
xor UO_4173 (O_4173,N_46195,N_40344);
and UO_4174 (O_4174,N_48460,N_42553);
and UO_4175 (O_4175,N_46082,N_46227);
or UO_4176 (O_4176,N_44700,N_48682);
nand UO_4177 (O_4177,N_42069,N_40084);
or UO_4178 (O_4178,N_44145,N_48050);
nor UO_4179 (O_4179,N_47279,N_41181);
nand UO_4180 (O_4180,N_43206,N_48315);
and UO_4181 (O_4181,N_46916,N_45666);
nor UO_4182 (O_4182,N_43562,N_44024);
nor UO_4183 (O_4183,N_40107,N_46390);
nand UO_4184 (O_4184,N_40512,N_41606);
xnor UO_4185 (O_4185,N_48064,N_43622);
nor UO_4186 (O_4186,N_40728,N_45408);
or UO_4187 (O_4187,N_49175,N_46917);
nor UO_4188 (O_4188,N_44060,N_43457);
or UO_4189 (O_4189,N_42840,N_49156);
nor UO_4190 (O_4190,N_49697,N_40225);
nor UO_4191 (O_4191,N_47682,N_49764);
nand UO_4192 (O_4192,N_41448,N_40124);
and UO_4193 (O_4193,N_48794,N_47811);
and UO_4194 (O_4194,N_40633,N_47481);
or UO_4195 (O_4195,N_40993,N_49340);
and UO_4196 (O_4196,N_49576,N_44404);
nand UO_4197 (O_4197,N_47050,N_41294);
nor UO_4198 (O_4198,N_48487,N_49364);
nor UO_4199 (O_4199,N_47389,N_45064);
or UO_4200 (O_4200,N_49429,N_42952);
xnor UO_4201 (O_4201,N_48663,N_40792);
and UO_4202 (O_4202,N_40283,N_43932);
xnor UO_4203 (O_4203,N_44102,N_43191);
nor UO_4204 (O_4204,N_41824,N_42892);
nor UO_4205 (O_4205,N_45005,N_44427);
nand UO_4206 (O_4206,N_43220,N_46065);
and UO_4207 (O_4207,N_44811,N_40960);
xor UO_4208 (O_4208,N_40577,N_48745);
nor UO_4209 (O_4209,N_46980,N_43611);
or UO_4210 (O_4210,N_47144,N_46024);
nand UO_4211 (O_4211,N_47465,N_47952);
and UO_4212 (O_4212,N_48618,N_42963);
nand UO_4213 (O_4213,N_48757,N_43621);
or UO_4214 (O_4214,N_45703,N_45544);
nor UO_4215 (O_4215,N_41384,N_44587);
or UO_4216 (O_4216,N_47692,N_43627);
or UO_4217 (O_4217,N_46600,N_47184);
and UO_4218 (O_4218,N_42676,N_40803);
nand UO_4219 (O_4219,N_44824,N_41301);
and UO_4220 (O_4220,N_46760,N_43282);
or UO_4221 (O_4221,N_46848,N_41966);
or UO_4222 (O_4222,N_45674,N_49135);
nand UO_4223 (O_4223,N_44510,N_46758);
or UO_4224 (O_4224,N_44514,N_41324);
or UO_4225 (O_4225,N_45221,N_44029);
or UO_4226 (O_4226,N_40677,N_40846);
nor UO_4227 (O_4227,N_44766,N_40642);
xor UO_4228 (O_4228,N_46374,N_43953);
and UO_4229 (O_4229,N_44762,N_43589);
nand UO_4230 (O_4230,N_46679,N_42711);
and UO_4231 (O_4231,N_46565,N_41595);
and UO_4232 (O_4232,N_45512,N_43474);
nor UO_4233 (O_4233,N_48988,N_48591);
nor UO_4234 (O_4234,N_44081,N_45011);
and UO_4235 (O_4235,N_45467,N_43296);
nand UO_4236 (O_4236,N_46154,N_48223);
or UO_4237 (O_4237,N_41572,N_44038);
nor UO_4238 (O_4238,N_43185,N_49866);
or UO_4239 (O_4239,N_46098,N_46711);
nor UO_4240 (O_4240,N_44048,N_49925);
or UO_4241 (O_4241,N_48285,N_44635);
and UO_4242 (O_4242,N_40913,N_46389);
and UO_4243 (O_4243,N_42831,N_43441);
xor UO_4244 (O_4244,N_49185,N_42891);
nor UO_4245 (O_4245,N_41661,N_48823);
and UO_4246 (O_4246,N_41838,N_41188);
nor UO_4247 (O_4247,N_43854,N_43402);
nand UO_4248 (O_4248,N_40183,N_40786);
or UO_4249 (O_4249,N_49959,N_41175);
nand UO_4250 (O_4250,N_42782,N_40835);
or UO_4251 (O_4251,N_45819,N_41960);
xor UO_4252 (O_4252,N_43717,N_47843);
nand UO_4253 (O_4253,N_49023,N_43843);
nor UO_4254 (O_4254,N_44475,N_45866);
or UO_4255 (O_4255,N_43398,N_44189);
and UO_4256 (O_4256,N_44558,N_48986);
or UO_4257 (O_4257,N_43353,N_47742);
nand UO_4258 (O_4258,N_45277,N_48772);
and UO_4259 (O_4259,N_41122,N_49615);
and UO_4260 (O_4260,N_46269,N_48509);
and UO_4261 (O_4261,N_40973,N_41672);
nor UO_4262 (O_4262,N_44345,N_42021);
xor UO_4263 (O_4263,N_44243,N_45607);
xor UO_4264 (O_4264,N_48567,N_41686);
nor UO_4265 (O_4265,N_43252,N_46991);
nor UO_4266 (O_4266,N_41462,N_42421);
xor UO_4267 (O_4267,N_40925,N_44820);
and UO_4268 (O_4268,N_44891,N_43963);
nand UO_4269 (O_4269,N_40932,N_40078);
nand UO_4270 (O_4270,N_42778,N_45590);
nor UO_4271 (O_4271,N_41275,N_40873);
nor UO_4272 (O_4272,N_44323,N_40692);
nand UO_4273 (O_4273,N_43198,N_45654);
nor UO_4274 (O_4274,N_45739,N_42534);
nand UO_4275 (O_4275,N_43671,N_40871);
or UO_4276 (O_4276,N_45787,N_49487);
or UO_4277 (O_4277,N_41568,N_40460);
nor UO_4278 (O_4278,N_44983,N_46291);
or UO_4279 (O_4279,N_44168,N_46858);
and UO_4280 (O_4280,N_45346,N_41894);
or UO_4281 (O_4281,N_46146,N_43439);
nand UO_4282 (O_4282,N_41796,N_45397);
nand UO_4283 (O_4283,N_44626,N_46665);
and UO_4284 (O_4284,N_43961,N_40824);
and UO_4285 (O_4285,N_45687,N_44683);
nor UO_4286 (O_4286,N_43533,N_41196);
and UO_4287 (O_4287,N_41671,N_47628);
or UO_4288 (O_4288,N_42743,N_41631);
and UO_4289 (O_4289,N_48630,N_49395);
xnor UO_4290 (O_4290,N_49075,N_44369);
nand UO_4291 (O_4291,N_46507,N_42287);
and UO_4292 (O_4292,N_49725,N_47784);
and UO_4293 (O_4293,N_48439,N_44828);
nor UO_4294 (O_4294,N_41065,N_43713);
or UO_4295 (O_4295,N_49270,N_45659);
or UO_4296 (O_4296,N_44837,N_44253);
and UO_4297 (O_4297,N_43636,N_43535);
and UO_4298 (O_4298,N_40953,N_40159);
and UO_4299 (O_4299,N_40016,N_42786);
xor UO_4300 (O_4300,N_47247,N_42675);
and UO_4301 (O_4301,N_43044,N_47657);
and UO_4302 (O_4302,N_46246,N_46421);
and UO_4303 (O_4303,N_46407,N_48828);
and UO_4304 (O_4304,N_40618,N_42175);
or UO_4305 (O_4305,N_41028,N_48022);
nor UO_4306 (O_4306,N_40366,N_43937);
and UO_4307 (O_4307,N_42946,N_49404);
and UO_4308 (O_4308,N_41971,N_43010);
and UO_4309 (O_4309,N_48459,N_41879);
and UO_4310 (O_4310,N_48306,N_48431);
nand UO_4311 (O_4311,N_47868,N_44830);
nand UO_4312 (O_4312,N_40470,N_41387);
nand UO_4313 (O_4313,N_40437,N_41087);
and UO_4314 (O_4314,N_44862,N_47333);
or UO_4315 (O_4315,N_42949,N_48158);
nand UO_4316 (O_4316,N_41295,N_44070);
nand UO_4317 (O_4317,N_43944,N_42594);
nand UO_4318 (O_4318,N_41460,N_43113);
nor UO_4319 (O_4319,N_46587,N_40631);
nor UO_4320 (O_4320,N_47115,N_45125);
or UO_4321 (O_4321,N_42933,N_43833);
nor UO_4322 (O_4322,N_47611,N_43998);
nor UO_4323 (O_4323,N_41261,N_43686);
and UO_4324 (O_4324,N_41516,N_41200);
and UO_4325 (O_4325,N_46944,N_48145);
or UO_4326 (O_4326,N_40767,N_46931);
or UO_4327 (O_4327,N_43446,N_49308);
nor UO_4328 (O_4328,N_40039,N_48503);
or UO_4329 (O_4329,N_42849,N_41775);
nand UO_4330 (O_4330,N_47675,N_43537);
nand UO_4331 (O_4331,N_48927,N_47705);
nand UO_4332 (O_4332,N_44497,N_43841);
and UO_4333 (O_4333,N_47058,N_44947);
and UO_4334 (O_4334,N_47296,N_48168);
xnor UO_4335 (O_4335,N_41611,N_49012);
or UO_4336 (O_4336,N_42684,N_40197);
or UO_4337 (O_4337,N_46472,N_45432);
or UO_4338 (O_4338,N_41548,N_49538);
nand UO_4339 (O_4339,N_49052,N_49107);
or UO_4340 (O_4340,N_45175,N_42127);
and UO_4341 (O_4341,N_42204,N_47743);
nand UO_4342 (O_4342,N_45331,N_44925);
or UO_4343 (O_4343,N_48991,N_47923);
and UO_4344 (O_4344,N_43344,N_43388);
xnor UO_4345 (O_4345,N_48859,N_44492);
nor UO_4346 (O_4346,N_42560,N_46895);
xnor UO_4347 (O_4347,N_46962,N_44221);
nand UO_4348 (O_4348,N_47257,N_47941);
nor UO_4349 (O_4349,N_49407,N_45513);
or UO_4350 (O_4350,N_40509,N_44852);
or UO_4351 (O_4351,N_44539,N_45158);
nor UO_4352 (O_4352,N_42155,N_43999);
nor UO_4353 (O_4353,N_40014,N_45771);
nand UO_4354 (O_4354,N_44115,N_42745);
and UO_4355 (O_4355,N_49598,N_49327);
nand UO_4356 (O_4356,N_49753,N_40240);
and UO_4357 (O_4357,N_43268,N_49767);
or UO_4358 (O_4358,N_41836,N_45825);
nand UO_4359 (O_4359,N_47139,N_43102);
nand UO_4360 (O_4360,N_43100,N_49670);
xor UO_4361 (O_4361,N_40714,N_40310);
nand UO_4362 (O_4362,N_43076,N_43926);
nand UO_4363 (O_4363,N_48563,N_49454);
and UO_4364 (O_4364,N_41957,N_41881);
nor UO_4365 (O_4365,N_45976,N_41156);
xor UO_4366 (O_4366,N_43712,N_46998);
xnor UO_4367 (O_4367,N_48827,N_47772);
and UO_4368 (O_4368,N_48165,N_47788);
nand UO_4369 (O_4369,N_43634,N_47043);
and UO_4370 (O_4370,N_45932,N_45469);
nor UO_4371 (O_4371,N_45092,N_49389);
xnor UO_4372 (O_4372,N_40566,N_49573);
and UO_4373 (O_4373,N_44055,N_46677);
and UO_4374 (O_4374,N_47549,N_41933);
and UO_4375 (O_4375,N_46742,N_48327);
xnor UO_4376 (O_4376,N_47341,N_46408);
or UO_4377 (O_4377,N_45255,N_45233);
and UO_4378 (O_4378,N_43663,N_45241);
or UO_4379 (O_4379,N_44731,N_44256);
and UO_4380 (O_4380,N_42726,N_43008);
xnor UO_4381 (O_4381,N_40694,N_48564);
xor UO_4382 (O_4382,N_42688,N_48855);
or UO_4383 (O_4383,N_42902,N_41950);
nor UO_4384 (O_4384,N_44944,N_48797);
or UO_4385 (O_4385,N_49748,N_44686);
or UO_4386 (O_4386,N_46447,N_47673);
xnor UO_4387 (O_4387,N_48936,N_40022);
nor UO_4388 (O_4388,N_44665,N_40040);
nand UO_4389 (O_4389,N_40986,N_46856);
nor UO_4390 (O_4390,N_45775,N_43367);
nor UO_4391 (O_4391,N_44051,N_49752);
or UO_4392 (O_4392,N_48805,N_44778);
xor UO_4393 (O_4393,N_42523,N_46684);
or UO_4394 (O_4394,N_49649,N_46942);
or UO_4395 (O_4395,N_42131,N_45629);
and UO_4396 (O_4396,N_43383,N_48965);
nor UO_4397 (O_4397,N_46592,N_46662);
or UO_4398 (O_4398,N_41861,N_43831);
nor UO_4399 (O_4399,N_47072,N_40700);
or UO_4400 (O_4400,N_48199,N_46037);
xnor UO_4401 (O_4401,N_44337,N_47485);
and UO_4402 (O_4402,N_46148,N_47852);
or UO_4403 (O_4403,N_47630,N_49926);
xnor UO_4404 (O_4404,N_41995,N_44147);
and UO_4405 (O_4405,N_45897,N_48081);
nor UO_4406 (O_4406,N_47120,N_45926);
nand UO_4407 (O_4407,N_47970,N_47683);
nand UO_4408 (O_4408,N_43839,N_42086);
nand UO_4409 (O_4409,N_43201,N_48198);
nand UO_4410 (O_4410,N_43164,N_41840);
or UO_4411 (O_4411,N_47199,N_41077);
nand UO_4412 (O_4412,N_43316,N_40597);
nand UO_4413 (O_4413,N_42319,N_49032);
or UO_4414 (O_4414,N_49645,N_46940);
nand UO_4415 (O_4415,N_48672,N_43459);
and UO_4416 (O_4416,N_42041,N_44304);
nor UO_4417 (O_4417,N_45518,N_44113);
and UO_4418 (O_4418,N_44434,N_46007);
nor UO_4419 (O_4419,N_45656,N_45706);
nor UO_4420 (O_4420,N_40921,N_47999);
xor UO_4421 (O_4421,N_41281,N_49432);
nor UO_4422 (O_4422,N_48429,N_46081);
nand UO_4423 (O_4423,N_49603,N_49974);
nand UO_4424 (O_4424,N_49602,N_46015);
nor UO_4425 (O_4425,N_47538,N_48816);
and UO_4426 (O_4426,N_49792,N_46063);
nand UO_4427 (O_4427,N_47983,N_43378);
nand UO_4428 (O_4428,N_49117,N_43356);
or UO_4429 (O_4429,N_45545,N_48659);
and UO_4430 (O_4430,N_41144,N_46156);
or UO_4431 (O_4431,N_49713,N_45181);
nand UO_4432 (O_4432,N_43131,N_46710);
nor UO_4433 (O_4433,N_45386,N_44130);
nor UO_4434 (O_4434,N_47973,N_40821);
nand UO_4435 (O_4435,N_45086,N_41447);
and UO_4436 (O_4436,N_43609,N_41637);
nand UO_4437 (O_4437,N_46088,N_45068);
nor UO_4438 (O_4438,N_44470,N_45943);
and UO_4439 (O_4439,N_48243,N_44781);
xor UO_4440 (O_4440,N_47136,N_49029);
or UO_4441 (O_4441,N_46546,N_49665);
and UO_4442 (O_4442,N_46359,N_40971);
and UO_4443 (O_4443,N_44623,N_41059);
or UO_4444 (O_4444,N_43968,N_43163);
and UO_4445 (O_4445,N_46984,N_42926);
and UO_4446 (O_4446,N_43391,N_42996);
nand UO_4447 (O_4447,N_48432,N_48019);
or UO_4448 (O_4448,N_49999,N_43838);
and UO_4449 (O_4449,N_42247,N_40837);
and UO_4450 (O_4450,N_43461,N_41821);
or UO_4451 (O_4451,N_46626,N_43129);
nor UO_4452 (O_4452,N_46310,N_44430);
or UO_4453 (O_4453,N_45482,N_40654);
and UO_4454 (O_4454,N_41763,N_48508);
or UO_4455 (O_4455,N_44412,N_47753);
and UO_4456 (O_4456,N_45515,N_41131);
or UO_4457 (O_4457,N_44114,N_48602);
nor UO_4458 (O_4458,N_46477,N_40055);
nand UO_4459 (O_4459,N_48759,N_45315);
nand UO_4460 (O_4460,N_40968,N_46732);
nand UO_4461 (O_4461,N_48237,N_40605);
nor UO_4462 (O_4462,N_43790,N_45225);
nand UO_4463 (O_4463,N_41566,N_47837);
or UO_4464 (O_4464,N_42206,N_49469);
and UO_4465 (O_4465,N_43637,N_49189);
nor UO_4466 (O_4466,N_43166,N_48009);
nand UO_4467 (O_4467,N_45053,N_45966);
and UO_4468 (O_4468,N_41911,N_45889);
nor UO_4469 (O_4469,N_40157,N_44295);
xnor UO_4470 (O_4470,N_47011,N_45599);
xor UO_4471 (O_4471,N_46311,N_43848);
nand UO_4472 (O_4472,N_42362,N_48758);
nand UO_4473 (O_4473,N_44333,N_40691);
nor UO_4474 (O_4474,N_42221,N_46958);
and UO_4475 (O_4475,N_42122,N_41907);
or UO_4476 (O_4476,N_42141,N_49675);
or UO_4477 (O_4477,N_42622,N_41233);
or UO_4478 (O_4478,N_44524,N_41624);
and UO_4479 (O_4479,N_40776,N_44932);
nor UO_4480 (O_4480,N_40808,N_44045);
nand UO_4481 (O_4481,N_46305,N_48541);
or UO_4482 (O_4482,N_46901,N_40977);
or UO_4483 (O_4483,N_42724,N_45843);
or UO_4484 (O_4484,N_41921,N_44599);
nand UO_4485 (O_4485,N_45365,N_45134);
nor UO_4486 (O_4486,N_46515,N_46567);
or UO_4487 (O_4487,N_49342,N_43934);
nand UO_4488 (O_4488,N_41835,N_41756);
nand UO_4489 (O_4489,N_48537,N_40956);
nand UO_4490 (O_4490,N_42703,N_47111);
or UO_4491 (O_4491,N_45299,N_49678);
or UO_4492 (O_4492,N_41236,N_43800);
or UO_4493 (O_4493,N_45699,N_44833);
nand UO_4494 (O_4494,N_48765,N_41302);
nor UO_4495 (O_4495,N_41872,N_48418);
xor UO_4496 (O_4496,N_45070,N_41544);
xnor UO_4497 (O_4497,N_45929,N_45459);
or UO_4498 (O_4498,N_42114,N_45089);
nor UO_4499 (O_4499,N_40523,N_46801);
and UO_4500 (O_4500,N_41502,N_43083);
nor UO_4501 (O_4501,N_42779,N_49253);
or UO_4502 (O_4502,N_47766,N_47415);
nand UO_4503 (O_4503,N_48642,N_43723);
or UO_4504 (O_4504,N_40404,N_46393);
nand UO_4505 (O_4505,N_44956,N_45494);
or UO_4506 (O_4506,N_43805,N_44724);
or UO_4507 (O_4507,N_41932,N_42632);
or UO_4508 (O_4508,N_49554,N_43172);
nand UO_4509 (O_4509,N_48634,N_49530);
and UO_4510 (O_4510,N_49273,N_48552);
nor UO_4511 (O_4511,N_40805,N_47638);
nand UO_4512 (O_4512,N_45697,N_46036);
and UO_4513 (O_4513,N_49131,N_49775);
and UO_4514 (O_4514,N_48782,N_44462);
and UO_4515 (O_4515,N_47678,N_43060);
xnor UO_4516 (O_4516,N_45922,N_42976);
xor UO_4517 (O_4517,N_49887,N_48493);
nor UO_4518 (O_4518,N_47600,N_41288);
xnor UO_4519 (O_4519,N_42602,N_46899);
or UO_4520 (O_4520,N_44202,N_48017);
or UO_4521 (O_4521,N_42060,N_47326);
nand UO_4522 (O_4522,N_40168,N_45420);
and UO_4523 (O_4523,N_45831,N_44505);
nor UO_4524 (O_4524,N_46520,N_45848);
nor UO_4525 (O_4525,N_48853,N_48454);
nand UO_4526 (O_4526,N_43000,N_40442);
and UO_4527 (O_4527,N_45019,N_47075);
nor UO_4528 (O_4528,N_48036,N_48291);
nand UO_4529 (O_4529,N_47322,N_43186);
or UO_4530 (O_4530,N_47125,N_46748);
or UO_4531 (O_4531,N_49416,N_49009);
nand UO_4532 (O_4532,N_44783,N_44796);
and UO_4533 (O_4533,N_45722,N_45969);
xor UO_4534 (O_4534,N_40586,N_44419);
xor UO_4535 (O_4535,N_46400,N_49056);
nand UO_4536 (O_4536,N_49674,N_45231);
and UO_4537 (O_4537,N_43698,N_42874);
and UO_4538 (O_4538,N_42495,N_45788);
nand UO_4539 (O_4539,N_42995,N_44393);
nand UO_4540 (O_4540,N_46689,N_46807);
or UO_4541 (O_4541,N_48756,N_46463);
and UO_4542 (O_4542,N_46589,N_45729);
and UO_4543 (O_4543,N_42732,N_46639);
nand UO_4544 (O_4544,N_47534,N_40563);
nor UO_4545 (O_4545,N_41128,N_44332);
nand UO_4546 (O_4546,N_48277,N_41870);
nand UO_4547 (O_4547,N_46935,N_42847);
xnor UO_4548 (O_4548,N_43811,N_48846);
and UO_4549 (O_4549,N_40485,N_48910);
nand UO_4550 (O_4550,N_43720,N_41119);
nor UO_4551 (O_4551,N_49636,N_47473);
and UO_4552 (O_4552,N_41518,N_40151);
nor UO_4553 (O_4553,N_41973,N_42623);
and UO_4554 (O_4554,N_47593,N_44162);
nand UO_4555 (O_4555,N_45826,N_49601);
nor UO_4556 (O_4556,N_45891,N_48213);
nand UO_4557 (O_4557,N_40129,N_40202);
nand UO_4558 (O_4558,N_49078,N_40420);
or UO_4559 (O_4559,N_41842,N_40490);
or UO_4560 (O_4560,N_49894,N_42525);
and UO_4561 (O_4561,N_43574,N_48812);
and UO_4562 (O_4562,N_44026,N_47310);
and UO_4563 (O_4563,N_43299,N_48170);
and UO_4564 (O_4564,N_42973,N_48209);
and UO_4565 (O_4565,N_46209,N_46815);
and UO_4566 (O_4566,N_44309,N_45229);
and UO_4567 (O_4567,N_45573,N_47754);
or UO_4568 (O_4568,N_40054,N_49466);
and UO_4569 (O_4569,N_45616,N_46774);
or UO_4570 (O_4570,N_45050,N_46912);
or UO_4571 (O_4571,N_49326,N_42216);
and UO_4572 (O_4572,N_44553,N_40136);
nand UO_4573 (O_4573,N_47806,N_40230);
or UO_4574 (O_4574,N_43085,N_41432);
and UO_4575 (O_4575,N_45116,N_46440);
and UO_4576 (O_4576,N_40990,N_48703);
nor UO_4577 (O_4577,N_44745,N_46198);
nand UO_4578 (O_4578,N_47447,N_45924);
nor UO_4579 (O_4579,N_40943,N_41762);
nor UO_4580 (O_4580,N_41090,N_48260);
or UO_4581 (O_4581,N_47388,N_46084);
xor UO_4582 (O_4582,N_48267,N_43877);
xnor UO_4583 (O_4583,N_41667,N_44224);
or UO_4584 (O_4584,N_47404,N_42981);
nand UO_4585 (O_4585,N_46454,N_48957);
xor UO_4586 (O_4586,N_42049,N_47452);
nor UO_4587 (O_4587,N_41562,N_47603);
and UO_4588 (O_4588,N_44609,N_40825);
xor UO_4589 (O_4589,N_43006,N_40651);
and UO_4590 (O_4590,N_44478,N_42691);
nand UO_4591 (O_4591,N_42588,N_40285);
and UO_4592 (O_4592,N_46676,N_47443);
nand UO_4593 (O_4593,N_45622,N_49045);
nor UO_4594 (O_4594,N_49703,N_45970);
or UO_4595 (O_4595,N_46611,N_49192);
nand UO_4596 (O_4596,N_44178,N_45406);
and UO_4597 (O_4597,N_44712,N_44991);
and UO_4598 (O_4598,N_45310,N_40819);
and UO_4599 (O_4599,N_45933,N_41123);
nor UO_4600 (O_4600,N_43289,N_40360);
and UO_4601 (O_4601,N_46249,N_45206);
or UO_4602 (O_4602,N_44813,N_44439);
nand UO_4603 (O_4603,N_41205,N_48427);
xnor UO_4604 (O_4604,N_48820,N_41183);
and UO_4605 (O_4605,N_42282,N_43073);
xor UO_4606 (O_4606,N_46737,N_42524);
nor UO_4607 (O_4607,N_47140,N_40521);
nand UO_4608 (O_4608,N_47091,N_46334);
nand UO_4609 (O_4609,N_42811,N_46067);
nor UO_4610 (O_4610,N_40788,N_48746);
nand UO_4611 (O_4611,N_40639,N_40434);
and UO_4612 (O_4612,N_40506,N_42583);
nand UO_4613 (O_4613,N_47916,N_40341);
or UO_4614 (O_4614,N_49017,N_44014);
nand UO_4615 (O_4615,N_47008,N_49702);
nand UO_4616 (O_4616,N_43003,N_44320);
or UO_4617 (O_4617,N_46493,N_49824);
or UO_4618 (O_4618,N_46419,N_41778);
or UO_4619 (O_4619,N_48348,N_42044);
nand UO_4620 (O_4620,N_40531,N_45465);
or UO_4621 (O_4621,N_48654,N_47337);
nor UO_4622 (O_4622,N_40929,N_47077);
nand UO_4623 (O_4623,N_44028,N_46628);
or UO_4624 (O_4624,N_48143,N_40941);
xor UO_4625 (O_4625,N_47188,N_40595);
nand UO_4626 (O_4626,N_43097,N_46232);
and UO_4627 (O_4627,N_44708,N_48031);
or UO_4628 (O_4628,N_42828,N_44059);
or UO_4629 (O_4629,N_44777,N_42153);
xor UO_4630 (O_4630,N_43337,N_48186);
nand UO_4631 (O_4631,N_44057,N_43199);
or UO_4632 (O_4632,N_40621,N_44254);
and UO_4633 (O_4633,N_46177,N_43791);
and UO_4634 (O_4634,N_43639,N_47994);
xor UO_4635 (O_4635,N_48478,N_49653);
nand UO_4636 (O_4636,N_49518,N_45238);
xnor UO_4637 (O_4637,N_46894,N_43031);
or UO_4638 (O_4638,N_41376,N_49634);
nor UO_4639 (O_4639,N_49211,N_46306);
or UO_4640 (O_4640,N_45373,N_43298);
or UO_4641 (O_4641,N_48124,N_41061);
or UO_4642 (O_4642,N_48234,N_41578);
or UO_4643 (O_4643,N_42781,N_42145);
or UO_4644 (O_4644,N_48055,N_43425);
and UO_4645 (O_4645,N_47978,N_41656);
and UO_4646 (O_4646,N_41863,N_47820);
nand UO_4647 (O_4647,N_43704,N_46321);
nand UO_4648 (O_4648,N_44487,N_41150);
nand UO_4649 (O_4649,N_46987,N_49125);
nor UO_4650 (O_4650,N_43559,N_48024);
and UO_4651 (O_4651,N_44289,N_42730);
and UO_4652 (O_4652,N_43852,N_42359);
or UO_4653 (O_4653,N_49669,N_43369);
nor UO_4654 (O_4654,N_44825,N_46178);
or UO_4655 (O_4655,N_43001,N_48270);
and UO_4656 (O_4656,N_49377,N_48391);
and UO_4657 (O_4657,N_45354,N_41859);
nand UO_4658 (O_4658,N_44754,N_43768);
or UO_4659 (O_4659,N_43155,N_41943);
nand UO_4660 (O_4660,N_48639,N_46079);
nand UO_4661 (O_4661,N_47694,N_48648);
nor UO_4662 (O_4662,N_48596,N_47395);
xor UO_4663 (O_4663,N_43979,N_40291);
nand UO_4664 (O_4664,N_47919,N_49174);
nor UO_4665 (O_4665,N_40838,N_47432);
nor UO_4666 (O_4666,N_49878,N_41718);
or UO_4667 (O_4667,N_48483,N_41311);
nor UO_4668 (O_4668,N_46044,N_43485);
or UO_4669 (O_4669,N_49328,N_46657);
nand UO_4670 (O_4670,N_46409,N_47513);
nor UO_4671 (O_4671,N_42884,N_46610);
nand UO_4672 (O_4672,N_41252,N_40256);
nand UO_4673 (O_4673,N_44922,N_43962);
nor UO_4674 (O_4674,N_49037,N_49990);
nor UO_4675 (O_4675,N_49087,N_46976);
and UO_4676 (O_4676,N_46017,N_42085);
or UO_4677 (O_4677,N_41086,N_40313);
and UO_4678 (O_4678,N_47518,N_48313);
xnor UO_4679 (O_4679,N_42192,N_47592);
or UO_4680 (O_4680,N_48720,N_42964);
or UO_4681 (O_4681,N_49179,N_42686);
or UO_4682 (O_4682,N_46806,N_43762);
and UO_4683 (O_4683,N_46429,N_46985);
and UO_4684 (O_4684,N_41316,N_49198);
nor UO_4685 (O_4685,N_48098,N_40706);
and UO_4686 (O_4686,N_40527,N_42353);
nor UO_4687 (O_4687,N_46427,N_48480);
xor UO_4688 (O_4688,N_46344,N_46415);
xor UO_4689 (O_4689,N_43248,N_48456);
nor UO_4690 (O_4690,N_46622,N_44220);
and UO_4691 (O_4691,N_49399,N_46625);
and UO_4692 (O_4692,N_42755,N_42186);
or UO_4693 (O_4693,N_40031,N_40583);
or UO_4694 (O_4694,N_47032,N_43798);
nand UO_4695 (O_4695,N_43556,N_45720);
nand UO_4696 (O_4696,N_47241,N_44682);
nand UO_4697 (O_4697,N_43782,N_44074);
or UO_4698 (O_4698,N_40784,N_43906);
xor UO_4699 (O_4699,N_47779,N_48490);
nand UO_4700 (O_4700,N_44359,N_46923);
nand UO_4701 (O_4701,N_44990,N_45099);
nand UO_4702 (O_4702,N_40999,N_40027);
xnor UO_4703 (O_4703,N_41543,N_44090);
or UO_4704 (O_4704,N_41804,N_49828);
nand UO_4705 (O_4705,N_41486,N_40255);
nor UO_4706 (O_4706,N_48763,N_40895);
and UO_4707 (O_4707,N_42912,N_41162);
and UO_4708 (O_4708,N_40623,N_48444);
or UO_4709 (O_4709,N_49600,N_47777);
nor UO_4710 (O_4710,N_49276,N_44318);
nor UO_4711 (O_4711,N_46218,N_48310);
or UO_4712 (O_4712,N_43381,N_49094);
xnor UO_4713 (O_4713,N_44822,N_42002);
and UO_4714 (O_4714,N_47500,N_46420);
nand UO_4715 (O_4715,N_47617,N_40936);
xnor UO_4716 (O_4716,N_43493,N_45658);
nor UO_4717 (O_4717,N_47903,N_42535);
and UO_4718 (O_4718,N_40369,N_41039);
and UO_4719 (O_4719,N_48798,N_43137);
and UO_4720 (O_4720,N_43065,N_47780);
and UO_4721 (O_4721,N_44287,N_48670);
and UO_4722 (O_4722,N_41406,N_41509);
or UO_4723 (O_4723,N_48417,N_42392);
nand UO_4724 (O_4724,N_45830,N_40214);
xor UO_4725 (O_4725,N_45455,N_43584);
nand UO_4726 (O_4726,N_49274,N_49627);
and UO_4727 (O_4727,N_45748,N_44676);
nand UO_4728 (O_4728,N_49679,N_42780);
or UO_4729 (O_4729,N_42948,N_42629);
or UO_4730 (O_4730,N_44873,N_40307);
xnor UO_4731 (O_4731,N_49372,N_45148);
nand UO_4732 (O_4732,N_45257,N_41575);
nor UO_4733 (O_4733,N_49077,N_41955);
nor UO_4734 (O_4734,N_40596,N_40418);
or UO_4735 (O_4735,N_46512,N_47261);
and UO_4736 (O_4736,N_44403,N_44772);
and UO_4737 (O_4737,N_43695,N_42410);
nand UO_4738 (O_4738,N_45797,N_47334);
nand UO_4739 (O_4739,N_41576,N_43173);
nor UO_4740 (O_4740,N_41478,N_48973);
or UO_4741 (O_4741,N_45330,N_46192);
nor UO_4742 (O_4742,N_47409,N_45728);
and UO_4743 (O_4743,N_41033,N_45815);
and UO_4744 (O_4744,N_43802,N_41491);
and UO_4745 (O_4745,N_42446,N_40844);
or UO_4746 (O_4746,N_49286,N_40675);
xor UO_4747 (O_4747,N_41847,N_49000);
or UO_4748 (O_4748,N_49494,N_43913);
nor UO_4749 (O_4749,N_47240,N_44363);
nand UO_4750 (O_4750,N_48993,N_42465);
or UO_4751 (O_4751,N_43927,N_44923);
and UO_4752 (O_4752,N_44354,N_41496);
nand UO_4753 (O_4753,N_46852,N_41319);
or UO_4754 (O_4754,N_42800,N_43952);
nand UO_4755 (O_4755,N_46860,N_45564);
nand UO_4756 (O_4756,N_42396,N_42071);
and UO_4757 (O_4757,N_41303,N_47632);
or UO_4758 (O_4758,N_47162,N_41355);
nand UO_4759 (O_4759,N_40697,N_48540);
or UO_4760 (O_4760,N_41210,N_46721);
nand UO_4761 (O_4761,N_49345,N_46281);
nand UO_4762 (O_4762,N_46867,N_45157);
nand UO_4763 (O_4763,N_44594,N_41356);
and UO_4764 (O_4764,N_43149,N_46049);
or UO_4765 (O_4765,N_41315,N_46220);
or UO_4766 (O_4766,N_43482,N_47614);
and UO_4767 (O_4767,N_41625,N_48899);
nand UO_4768 (O_4768,N_42822,N_42209);
and UO_4769 (O_4769,N_43212,N_42084);
or UO_4770 (O_4770,N_44788,N_47597);
or UO_4771 (O_4771,N_45516,N_43678);
nor UO_4772 (O_4772,N_43974,N_44008);
or UO_4773 (O_4773,N_42435,N_47795);
xor UO_4774 (O_4774,N_49062,N_46738);
xor UO_4775 (O_4775,N_43309,N_49355);
or UO_4776 (O_4776,N_40422,N_45638);
and UO_4777 (O_4777,N_47295,N_47720);
nand UO_4778 (O_4778,N_49366,N_48398);
nand UO_4779 (O_4779,N_45348,N_49428);
nor UO_4780 (O_4780,N_41218,N_45182);
and UO_4781 (O_4781,N_48774,N_46607);
xnor UO_4782 (O_4782,N_49696,N_45008);
nor UO_4783 (O_4783,N_48547,N_41918);
and UO_4784 (O_4784,N_48302,N_41022);
and UO_4785 (O_4785,N_47398,N_48334);
or UO_4786 (O_4786,N_41615,N_45437);
or UO_4787 (O_4787,N_42658,N_45317);
nor UO_4788 (O_4788,N_44517,N_41642);
or UO_4789 (O_4789,N_49642,N_43617);
and UO_4790 (O_4790,N_43941,N_45278);
nand UO_4791 (O_4791,N_41499,N_40331);
or UO_4792 (O_4792,N_45750,N_46603);
and UO_4793 (O_4793,N_41115,N_40901);
or UO_4794 (O_4794,N_48111,N_41601);
nand UO_4795 (O_4795,N_44370,N_45007);
and UO_4796 (O_4796,N_46831,N_49472);
or UO_4797 (O_4797,N_45957,N_43382);
nand UO_4798 (O_4798,N_48990,N_41127);
and UO_4799 (O_4799,N_46687,N_49071);
nor UO_4800 (O_4800,N_43836,N_44263);
nor UO_4801 (O_4801,N_43277,N_43471);
nand UO_4802 (O_4802,N_44451,N_43132);
or UO_4803 (O_4803,N_44255,N_45643);
and UO_4804 (O_4804,N_40062,N_48299);
xor UO_4805 (O_4805,N_45911,N_49217);
and UO_4806 (O_4806,N_44017,N_44917);
or UO_4807 (O_4807,N_48347,N_47543);
or UO_4808 (O_4808,N_40676,N_42923);
or UO_4809 (O_4809,N_46110,N_49483);
or UO_4810 (O_4810,N_43756,N_46960);
or UO_4811 (O_4811,N_42619,N_48788);
or UO_4812 (O_4812,N_47790,N_42719);
nor UO_4813 (O_4813,N_45923,N_43365);
or UO_4814 (O_4814,N_43286,N_48318);
or UO_4815 (O_4815,N_48981,N_48529);
nor UO_4816 (O_4816,N_45794,N_44139);
xor UO_4817 (O_4817,N_47574,N_47420);
nand UO_4818 (O_4818,N_42879,N_47071);
or UO_4819 (O_4819,N_42027,N_48594);
or UO_4820 (O_4820,N_49200,N_43722);
and UO_4821 (O_4821,N_47114,N_42013);
nor UO_4822 (O_4822,N_41808,N_45662);
and UO_4823 (O_4823,N_44212,N_47208);
or UO_4824 (O_4824,N_49540,N_46073);
or UO_4825 (O_4825,N_47365,N_42057);
and UO_4826 (O_4826,N_44050,N_44367);
nor UO_4827 (O_4827,N_46743,N_41078);
nand UO_4828 (O_4828,N_41411,N_48989);
or UO_4829 (O_4829,N_44204,N_43503);
nand UO_4830 (O_4830,N_40161,N_49193);
and UO_4831 (O_4831,N_40174,N_46761);
nand UO_4832 (O_4832,N_43421,N_48390);
and UO_4833 (O_4833,N_48185,N_48047);
nand UO_4834 (O_4834,N_45503,N_40726);
or UO_4835 (O_4835,N_47320,N_43801);
nor UO_4836 (O_4836,N_43214,N_44883);
xor UO_4837 (O_4837,N_41363,N_43520);
and UO_4838 (O_4838,N_47503,N_48606);
nor UO_4839 (O_4839,N_49165,N_47652);
and UO_4840 (O_4840,N_47166,N_47750);
and UO_4841 (O_4841,N_48200,N_41174);
and UO_4842 (O_4842,N_48375,N_46028);
and UO_4843 (O_4843,N_41394,N_49980);
nand UO_4844 (O_4844,N_45871,N_40772);
or UO_4845 (O_4845,N_49319,N_43868);
nand UO_4846 (O_4846,N_48685,N_48152);
nor UO_4847 (O_4847,N_46075,N_49061);
nor UO_4848 (O_4848,N_47039,N_40339);
and UO_4849 (O_4849,N_40775,N_49463);
nand UO_4850 (O_4850,N_43249,N_48632);
nor UO_4851 (O_4851,N_48228,N_42162);
or UO_4852 (O_4852,N_45685,N_43726);
or UO_4853 (O_4853,N_41766,N_49591);
and UO_4854 (O_4854,N_48922,N_44603);
nor UO_4855 (O_4855,N_40777,N_42478);
nand UO_4856 (O_4856,N_44767,N_49166);
and UO_4857 (O_4857,N_41032,N_47244);
xor UO_4858 (O_4858,N_46499,N_45140);
nor UO_4859 (O_4859,N_45335,N_42471);
nor UO_4860 (O_4860,N_42661,N_46508);
and UO_4861 (O_4861,N_44870,N_41905);
and UO_4862 (O_4862,N_48832,N_43190);
and UO_4863 (O_4863,N_41428,N_48675);
xnor UO_4864 (O_4864,N_40425,N_48869);
and UO_4865 (O_4865,N_48615,N_41004);
or UO_4866 (O_4866,N_46205,N_47577);
nor UO_4867 (O_4867,N_42152,N_45425);
nor UO_4868 (O_4868,N_49140,N_43908);
nor UO_4869 (O_4869,N_44785,N_46921);
nor UO_4870 (O_4870,N_47340,N_43586);
and UO_4871 (O_4871,N_49471,N_49869);
or UO_4872 (O_4872,N_48447,N_43080);
or UO_4873 (O_4873,N_43672,N_40045);
nand UO_4874 (O_4874,N_47331,N_41348);
and UO_4875 (O_4875,N_48985,N_40609);
or UO_4876 (O_4876,N_41358,N_40709);
nor UO_4877 (O_4877,N_44177,N_46725);
or UO_4878 (O_4878,N_43778,N_44285);
or UO_4879 (O_4879,N_48148,N_45630);
nand UO_4880 (O_4880,N_49972,N_42150);
and UO_4881 (O_4881,N_43170,N_44780);
xor UO_4882 (O_4882,N_49802,N_48811);
nand UO_4883 (O_4883,N_47520,N_41064);
nand UO_4884 (O_4884,N_41132,N_42258);
and UO_4885 (O_4885,N_48116,N_49021);
nand UO_4886 (O_4886,N_40908,N_44108);
nand UO_4887 (O_4887,N_48974,N_40553);
nor UO_4888 (O_4888,N_46702,N_43539);
nand UO_4889 (O_4889,N_49296,N_41694);
nand UO_4890 (O_4890,N_48466,N_43022);
or UO_4891 (O_4891,N_41780,N_40982);
nor UO_4892 (O_4892,N_42390,N_48332);
and UO_4893 (O_4893,N_45915,N_47490);
nand UO_4894 (O_4894,N_44749,N_45029);
and UO_4895 (O_4895,N_46234,N_40356);
or UO_4896 (O_4896,N_43435,N_43068);
and UO_4897 (O_4897,N_48793,N_49906);
and UO_4898 (O_4898,N_44325,N_46590);
and UO_4899 (O_4899,N_44456,N_41640);
nand UO_4900 (O_4900,N_41124,N_45114);
nor UO_4901 (O_4901,N_42112,N_47080);
or UO_4902 (O_4902,N_49760,N_45579);
nor UO_4903 (O_4903,N_48229,N_41017);
nand UO_4904 (O_4904,N_47556,N_46466);
and UO_4905 (O_4905,N_43669,N_41179);
and UO_4906 (O_4906,N_46229,N_46821);
nand UO_4907 (O_4907,N_46647,N_42893);
xnor UO_4908 (O_4908,N_41650,N_47277);
nand UO_4909 (O_4909,N_42042,N_41900);
xnor UO_4910 (O_4910,N_42531,N_48732);
or UO_4911 (O_4911,N_45169,N_40190);
nand UO_4912 (O_4912,N_45917,N_44748);
and UO_4913 (O_4913,N_43317,N_46837);
nor UO_4914 (O_4914,N_47606,N_46215);
and UO_4915 (O_4915,N_48141,N_49783);
and UO_4916 (O_4916,N_45045,N_42674);
and UO_4917 (O_4917,N_44756,N_43881);
or UO_4918 (O_4918,N_48357,N_46315);
and UO_4919 (O_4919,N_49375,N_49204);
nand UO_4920 (O_4920,N_46656,N_44563);
or UO_4921 (O_4921,N_47915,N_49048);
or UO_4922 (O_4922,N_47863,N_49221);
and UO_4923 (O_4923,N_42371,N_46174);
nor UO_4924 (O_4924,N_49967,N_46999);
or UO_4925 (O_4925,N_45118,N_42491);
and UO_4926 (O_4926,N_44643,N_49441);
xnor UO_4927 (O_4927,N_48400,N_44819);
and UO_4928 (O_4928,N_43138,N_47633);
xnor UO_4929 (O_4929,N_47835,N_46401);
nor UO_4930 (O_4930,N_41498,N_47419);
and UO_4931 (O_4931,N_48967,N_44531);
or UO_4932 (O_4932,N_49652,N_45892);
and UO_4933 (O_4933,N_42075,N_47137);
and UO_4934 (O_4934,N_49284,N_47966);
and UO_4935 (O_4935,N_41573,N_45507);
nor UO_4936 (O_4936,N_40282,N_46430);
and UO_4937 (O_4937,N_42723,N_44940);
and UO_4938 (O_4938,N_45842,N_45813);
or UO_4939 (O_4939,N_45542,N_43773);
and UO_4940 (O_4940,N_46558,N_44634);
nand UO_4941 (O_4941,N_44290,N_46582);
nand UO_4942 (O_4942,N_46637,N_47219);
and UO_4943 (O_4943,N_41906,N_48609);
or UO_4944 (O_4944,N_42290,N_42965);
xor UO_4945 (O_4945,N_46920,N_44771);
or UO_4946 (O_4946,N_49034,N_42125);
xor UO_4947 (O_4947,N_46035,N_45073);
nand UO_4948 (O_4948,N_40049,N_47318);
and UO_4949 (O_4949,N_42010,N_42480);
or UO_4950 (O_4950,N_49692,N_45122);
nand UO_4951 (O_4951,N_46811,N_42111);
nand UO_4952 (O_4952,N_40826,N_46833);
nor UO_4953 (O_4953,N_42327,N_41464);
and UO_4954 (O_4954,N_48600,N_49351);
or UO_4955 (O_4955,N_48636,N_49112);
nor UO_4956 (O_4956,N_48287,N_40915);
nor UO_4957 (O_4957,N_42544,N_41998);
nor UO_4958 (O_4958,N_41068,N_43401);
and UO_4959 (O_4959,N_49888,N_46226);
and UO_4960 (O_4960,N_43035,N_43141);
and UO_4961 (O_4961,N_42502,N_44518);
and UO_4962 (O_4962,N_40729,N_44072);
or UO_4963 (O_4963,N_45044,N_46772);
and UO_4964 (O_4964,N_49564,N_45767);
nor UO_4965 (O_4965,N_49912,N_46719);
nor UO_4966 (O_4966,N_43389,N_43901);
nor UO_4967 (O_4967,N_44324,N_45681);
and UO_4968 (O_4968,N_40298,N_45303);
and UO_4969 (O_4969,N_41100,N_45710);
and UO_4970 (O_4970,N_40830,N_40440);
nand UO_4971 (O_4971,N_44219,N_44739);
and UO_4972 (O_4972,N_45672,N_44380);
xor UO_4973 (O_4973,N_42873,N_48750);
or UO_4974 (O_4974,N_49064,N_49510);
nand UO_4975 (O_4975,N_49057,N_43724);
nand UO_4976 (O_4976,N_41701,N_42598);
nor UO_4977 (O_4977,N_44338,N_49387);
nand UO_4978 (O_4978,N_47997,N_43287);
xor UO_4979 (O_4979,N_43360,N_44150);
nor UO_4980 (O_4980,N_44672,N_43049);
nand UO_4981 (O_4981,N_47495,N_44970);
nand UO_4982 (O_4982,N_46182,N_43581);
nand UO_4983 (O_4983,N_42484,N_49954);
nor UO_4984 (O_4984,N_46053,N_40614);
and UO_4985 (O_4985,N_41242,N_45707);
or UO_4986 (O_4986,N_48934,N_42913);
nor UO_4987 (O_4987,N_44205,N_41592);
xnor UO_4988 (O_4988,N_40845,N_49850);
nand UO_4989 (O_4989,N_43125,N_48403);
nor UO_4990 (O_4990,N_48997,N_44483);
nand UO_4991 (O_4991,N_46357,N_46878);
nand UO_4992 (O_4992,N_47889,N_43496);
and UO_4993 (O_4993,N_49035,N_46779);
xor UO_4994 (O_4994,N_47129,N_41552);
and UO_4995 (O_4995,N_40812,N_46470);
or UO_4996 (O_4996,N_44037,N_49647);
nor UO_4997 (O_4997,N_44580,N_47862);
and UO_4998 (O_4998,N_46601,N_46187);
nand UO_4999 (O_4999,N_45852,N_47238);
endmodule