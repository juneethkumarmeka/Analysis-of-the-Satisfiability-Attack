module basic_500_3000_500_5_levels_2xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_281,In_404);
and U1 (N_1,In_351,In_269);
nand U2 (N_2,In_102,In_438);
or U3 (N_3,In_59,In_324);
or U4 (N_4,In_284,In_148);
and U5 (N_5,In_424,In_412);
nor U6 (N_6,In_239,In_110);
or U7 (N_7,In_235,In_464);
nand U8 (N_8,In_211,In_330);
or U9 (N_9,In_48,In_334);
nor U10 (N_10,In_21,In_302);
or U11 (N_11,In_264,In_497);
or U12 (N_12,In_232,In_46);
or U13 (N_13,In_210,In_278);
nand U14 (N_14,In_309,In_405);
or U15 (N_15,In_119,In_203);
and U16 (N_16,In_73,In_267);
nor U17 (N_17,In_9,In_230);
or U18 (N_18,In_172,In_47);
or U19 (N_19,In_494,In_435);
nor U20 (N_20,In_123,In_447);
and U21 (N_21,In_261,In_234);
or U22 (N_22,In_190,In_87);
and U23 (N_23,In_157,In_384);
nor U24 (N_24,In_250,In_33);
nor U25 (N_25,In_456,In_204);
nand U26 (N_26,In_331,In_376);
nor U27 (N_27,In_255,In_275);
and U28 (N_28,In_104,In_4);
or U29 (N_29,In_368,In_429);
nor U30 (N_30,In_150,In_94);
nor U31 (N_31,In_256,In_365);
nor U32 (N_32,In_38,In_249);
and U33 (N_33,In_214,In_205);
nand U34 (N_34,In_348,In_373);
or U35 (N_35,In_30,In_332);
or U36 (N_36,In_175,In_98);
nand U37 (N_37,In_292,In_370);
and U38 (N_38,In_470,In_403);
or U39 (N_39,In_137,In_51);
nor U40 (N_40,In_116,In_446);
nand U41 (N_41,In_485,In_359);
and U42 (N_42,In_27,In_481);
nor U43 (N_43,In_53,In_316);
nor U44 (N_44,In_147,In_294);
nand U45 (N_45,In_377,In_92);
nand U46 (N_46,In_71,In_493);
nor U47 (N_47,In_76,In_186);
and U48 (N_48,In_188,In_286);
or U49 (N_49,In_222,In_12);
and U50 (N_50,In_430,In_22);
or U51 (N_51,In_455,In_483);
or U52 (N_52,In_419,In_138);
nand U53 (N_53,In_374,In_69);
or U54 (N_54,In_372,In_260);
and U55 (N_55,In_262,In_346);
or U56 (N_56,In_417,In_224);
and U57 (N_57,In_364,In_496);
xnor U58 (N_58,In_390,In_469);
or U59 (N_59,In_304,In_454);
or U60 (N_60,In_449,In_81);
and U61 (N_61,In_398,In_149);
or U62 (N_62,In_13,In_167);
and U63 (N_63,In_171,In_174);
and U64 (N_64,In_215,In_333);
or U65 (N_65,In_245,In_194);
nor U66 (N_66,In_460,In_335);
nand U67 (N_67,In_144,In_476);
or U68 (N_68,In_162,In_307);
and U69 (N_69,In_233,In_380);
nor U70 (N_70,In_451,In_431);
nand U71 (N_71,In_236,In_375);
and U72 (N_72,In_158,In_37);
xnor U73 (N_73,In_58,In_296);
and U74 (N_74,In_289,In_246);
nand U75 (N_75,In_421,In_313);
and U76 (N_76,In_479,In_314);
nand U77 (N_77,In_401,In_442);
nor U78 (N_78,In_42,In_213);
nand U79 (N_79,In_347,In_107);
and U80 (N_80,In_394,In_487);
and U81 (N_81,In_461,In_11);
nor U82 (N_82,In_322,In_279);
or U83 (N_83,In_410,In_77);
or U84 (N_84,In_128,In_237);
nand U85 (N_85,In_121,In_40);
nand U86 (N_86,In_89,In_29);
and U87 (N_87,In_60,In_32);
xnor U88 (N_88,In_274,In_399);
or U89 (N_89,In_432,In_299);
nand U90 (N_90,In_66,In_135);
or U91 (N_91,In_474,In_96);
and U92 (N_92,In_221,In_463);
and U93 (N_93,In_385,In_25);
nor U94 (N_94,In_450,In_181);
or U95 (N_95,In_68,In_78);
or U96 (N_96,In_407,In_409);
nor U97 (N_97,In_413,In_218);
nor U98 (N_98,In_329,In_82);
or U99 (N_99,In_393,In_56);
nand U100 (N_100,In_341,In_423);
and U101 (N_101,In_379,In_103);
and U102 (N_102,In_342,In_400);
nand U103 (N_103,In_273,In_337);
nand U104 (N_104,In_439,In_306);
nor U105 (N_105,In_295,In_349);
or U106 (N_106,In_179,In_276);
and U107 (N_107,In_416,In_259);
nor U108 (N_108,In_223,In_160);
nor U109 (N_109,In_226,In_139);
nor U110 (N_110,In_343,In_391);
nor U111 (N_111,In_36,In_23);
nor U112 (N_112,In_195,In_231);
and U113 (N_113,In_257,In_445);
nand U114 (N_114,In_193,In_18);
nor U115 (N_115,In_287,In_358);
and U116 (N_116,In_491,In_145);
and U117 (N_117,In_434,In_344);
and U118 (N_118,In_65,In_219);
and U119 (N_119,In_108,In_441);
nand U120 (N_120,In_143,In_206);
nor U121 (N_121,In_124,In_253);
xnor U122 (N_122,In_39,In_64);
or U123 (N_123,In_122,In_14);
nand U124 (N_124,In_254,In_305);
nand U125 (N_125,In_371,In_406);
nand U126 (N_126,In_244,In_184);
nor U127 (N_127,In_270,In_425);
or U128 (N_128,In_489,In_345);
nand U129 (N_129,In_85,In_217);
or U130 (N_130,In_197,In_15);
nor U131 (N_131,In_319,In_24);
and U132 (N_132,In_166,In_49);
and U133 (N_133,In_177,In_387);
nand U134 (N_134,In_420,In_315);
nand U135 (N_135,In_99,In_452);
nand U136 (N_136,In_339,In_207);
or U137 (N_137,In_482,In_310);
or U138 (N_138,In_422,In_288);
nor U139 (N_139,In_62,In_31);
or U140 (N_140,In_202,In_84);
nand U141 (N_141,In_132,In_72);
nor U142 (N_142,In_468,In_325);
nand U143 (N_143,In_475,In_303);
xnor U144 (N_144,In_159,In_114);
nor U145 (N_145,In_402,In_152);
or U146 (N_146,In_1,In_176);
nor U147 (N_147,In_75,In_228);
or U148 (N_148,In_378,In_396);
nor U149 (N_149,In_318,In_251);
and U150 (N_150,In_198,In_208);
and U151 (N_151,In_361,In_473);
or U152 (N_152,In_43,In_41);
and U153 (N_153,In_155,In_74);
xnor U154 (N_154,In_408,In_83);
nand U155 (N_155,In_227,In_354);
or U156 (N_156,In_388,In_185);
nand U157 (N_157,In_86,In_252);
nand U158 (N_158,In_20,In_282);
or U159 (N_159,In_101,In_352);
or U160 (N_160,In_216,In_353);
nor U161 (N_161,In_2,In_277);
and U162 (N_162,In_52,In_178);
nor U163 (N_163,In_290,In_247);
or U164 (N_164,In_133,In_165);
or U165 (N_165,In_467,In_8);
and U166 (N_166,In_297,In_453);
xor U167 (N_167,In_258,In_67);
nand U168 (N_168,In_19,In_243);
nand U169 (N_169,In_495,In_57);
nor U170 (N_170,In_486,In_115);
or U171 (N_171,In_285,In_444);
or U172 (N_172,In_283,In_383);
nor U173 (N_173,In_180,In_240);
nand U174 (N_174,In_161,In_189);
and U175 (N_175,In_28,In_477);
nand U176 (N_176,In_490,In_50);
nor U177 (N_177,In_142,In_268);
nor U178 (N_178,In_118,In_300);
or U179 (N_179,In_386,In_301);
nand U180 (N_180,In_168,In_201);
nand U181 (N_181,In_326,In_112);
nor U182 (N_182,In_88,In_321);
xnor U183 (N_183,In_266,In_126);
and U184 (N_184,In_323,In_411);
nand U185 (N_185,In_338,In_170);
nand U186 (N_186,In_105,In_428);
or U187 (N_187,In_366,In_462);
nor U188 (N_188,In_169,In_3);
nor U189 (N_189,In_111,In_16);
and U190 (N_190,In_5,In_153);
nor U191 (N_191,In_26,In_478);
nor U192 (N_192,In_311,In_492);
nand U193 (N_193,In_196,In_173);
nor U194 (N_194,In_357,In_17);
nor U195 (N_195,In_355,In_443);
and U196 (N_196,In_472,In_106);
nor U197 (N_197,In_134,In_238);
nand U198 (N_198,In_440,In_54);
and U199 (N_199,In_127,In_272);
or U200 (N_200,In_209,In_97);
nor U201 (N_201,In_164,In_437);
nand U202 (N_202,In_280,In_360);
and U203 (N_203,In_136,In_248);
nand U204 (N_204,In_488,In_298);
and U205 (N_205,In_7,In_381);
and U206 (N_206,In_225,In_6);
or U207 (N_207,In_340,In_100);
or U208 (N_208,In_436,In_44);
xnor U209 (N_209,In_93,In_480);
or U210 (N_210,In_414,In_395);
and U211 (N_211,In_156,In_308);
nand U212 (N_212,In_242,In_163);
nor U213 (N_213,In_392,In_55);
nand U214 (N_214,In_187,In_90);
nand U215 (N_215,In_459,In_293);
nand U216 (N_216,In_350,In_458);
nor U217 (N_217,In_466,In_45);
and U218 (N_218,In_448,In_320);
and U219 (N_219,In_192,In_369);
or U220 (N_220,In_498,In_182);
nand U221 (N_221,In_327,In_389);
nor U222 (N_222,In_312,In_120);
nor U223 (N_223,In_79,In_140);
or U224 (N_224,In_10,In_117);
nand U225 (N_225,In_0,In_418);
nor U226 (N_226,In_212,In_199);
and U227 (N_227,In_362,In_426);
and U228 (N_228,In_356,In_229);
or U229 (N_229,In_125,In_415);
nand U230 (N_230,In_397,In_457);
or U231 (N_231,In_95,In_317);
nor U232 (N_232,In_336,In_484);
nor U233 (N_233,In_146,In_291);
nor U234 (N_234,In_183,In_382);
or U235 (N_235,In_433,In_271);
and U236 (N_236,In_220,In_113);
or U237 (N_237,In_328,In_427);
nand U238 (N_238,In_130,In_80);
nand U239 (N_239,In_367,In_63);
nand U240 (N_240,In_151,In_471);
or U241 (N_241,In_154,In_499);
and U242 (N_242,In_265,In_109);
xor U243 (N_243,In_263,In_465);
nor U244 (N_244,In_191,In_61);
nand U245 (N_245,In_91,In_200);
or U246 (N_246,In_141,In_363);
or U247 (N_247,In_131,In_70);
and U248 (N_248,In_35,In_129);
nor U249 (N_249,In_241,In_34);
and U250 (N_250,In_51,In_87);
xor U251 (N_251,In_18,In_318);
or U252 (N_252,In_475,In_307);
nor U253 (N_253,In_438,In_300);
nor U254 (N_254,In_37,In_207);
nand U255 (N_255,In_477,In_76);
or U256 (N_256,In_268,In_37);
nor U257 (N_257,In_132,In_447);
or U258 (N_258,In_469,In_83);
and U259 (N_259,In_448,In_300);
nand U260 (N_260,In_151,In_449);
or U261 (N_261,In_17,In_119);
and U262 (N_262,In_74,In_445);
or U263 (N_263,In_180,In_309);
or U264 (N_264,In_37,In_48);
nor U265 (N_265,In_345,In_453);
or U266 (N_266,In_172,In_362);
and U267 (N_267,In_480,In_347);
nand U268 (N_268,In_204,In_231);
nor U269 (N_269,In_273,In_192);
and U270 (N_270,In_193,In_100);
nor U271 (N_271,In_232,In_416);
and U272 (N_272,In_202,In_423);
or U273 (N_273,In_41,In_376);
and U274 (N_274,In_165,In_344);
nor U275 (N_275,In_140,In_238);
nor U276 (N_276,In_165,In_175);
nor U277 (N_277,In_471,In_331);
nand U278 (N_278,In_109,In_123);
and U279 (N_279,In_218,In_476);
xnor U280 (N_280,In_111,In_203);
xor U281 (N_281,In_6,In_326);
and U282 (N_282,In_375,In_147);
nor U283 (N_283,In_112,In_496);
or U284 (N_284,In_93,In_0);
or U285 (N_285,In_413,In_179);
and U286 (N_286,In_26,In_242);
or U287 (N_287,In_197,In_163);
and U288 (N_288,In_173,In_200);
nor U289 (N_289,In_498,In_334);
nand U290 (N_290,In_352,In_43);
and U291 (N_291,In_349,In_174);
nand U292 (N_292,In_18,In_419);
and U293 (N_293,In_37,In_395);
nand U294 (N_294,In_30,In_490);
and U295 (N_295,In_161,In_142);
or U296 (N_296,In_485,In_114);
nor U297 (N_297,In_366,In_372);
nand U298 (N_298,In_282,In_73);
nor U299 (N_299,In_139,In_140);
and U300 (N_300,In_252,In_204);
and U301 (N_301,In_20,In_399);
nor U302 (N_302,In_124,In_307);
nand U303 (N_303,In_191,In_468);
nor U304 (N_304,In_454,In_142);
or U305 (N_305,In_240,In_40);
nand U306 (N_306,In_39,In_140);
nor U307 (N_307,In_120,In_355);
and U308 (N_308,In_360,In_81);
or U309 (N_309,In_458,In_315);
or U310 (N_310,In_380,In_221);
or U311 (N_311,In_61,In_202);
and U312 (N_312,In_228,In_26);
nor U313 (N_313,In_174,In_366);
and U314 (N_314,In_349,In_355);
xnor U315 (N_315,In_489,In_153);
and U316 (N_316,In_189,In_455);
or U317 (N_317,In_105,In_487);
nor U318 (N_318,In_405,In_320);
nor U319 (N_319,In_421,In_465);
nor U320 (N_320,In_191,In_24);
or U321 (N_321,In_422,In_63);
nand U322 (N_322,In_391,In_137);
and U323 (N_323,In_453,In_427);
nand U324 (N_324,In_376,In_245);
and U325 (N_325,In_480,In_478);
and U326 (N_326,In_265,In_464);
nand U327 (N_327,In_24,In_437);
or U328 (N_328,In_425,In_464);
or U329 (N_329,In_81,In_103);
and U330 (N_330,In_240,In_405);
nor U331 (N_331,In_243,In_117);
nand U332 (N_332,In_38,In_233);
nand U333 (N_333,In_385,In_331);
or U334 (N_334,In_462,In_223);
nor U335 (N_335,In_484,In_173);
nor U336 (N_336,In_8,In_162);
nor U337 (N_337,In_269,In_106);
and U338 (N_338,In_26,In_216);
nor U339 (N_339,In_242,In_491);
or U340 (N_340,In_372,In_87);
or U341 (N_341,In_383,In_347);
and U342 (N_342,In_112,In_176);
or U343 (N_343,In_295,In_86);
and U344 (N_344,In_90,In_234);
and U345 (N_345,In_335,In_311);
and U346 (N_346,In_498,In_224);
nand U347 (N_347,In_416,In_421);
and U348 (N_348,In_443,In_81);
nor U349 (N_349,In_70,In_215);
and U350 (N_350,In_219,In_185);
and U351 (N_351,In_469,In_464);
nand U352 (N_352,In_206,In_309);
and U353 (N_353,In_106,In_448);
or U354 (N_354,In_497,In_489);
xnor U355 (N_355,In_214,In_372);
nand U356 (N_356,In_328,In_204);
nor U357 (N_357,In_396,In_195);
nand U358 (N_358,In_228,In_176);
and U359 (N_359,In_188,In_497);
nand U360 (N_360,In_484,In_37);
nor U361 (N_361,In_488,In_443);
nand U362 (N_362,In_336,In_450);
nand U363 (N_363,In_124,In_189);
and U364 (N_364,In_127,In_402);
xnor U365 (N_365,In_97,In_355);
xnor U366 (N_366,In_469,In_457);
nand U367 (N_367,In_201,In_219);
and U368 (N_368,In_247,In_149);
or U369 (N_369,In_248,In_96);
or U370 (N_370,In_393,In_443);
nand U371 (N_371,In_26,In_372);
or U372 (N_372,In_442,In_246);
and U373 (N_373,In_91,In_361);
or U374 (N_374,In_83,In_284);
and U375 (N_375,In_229,In_240);
nor U376 (N_376,In_354,In_7);
nor U377 (N_377,In_384,In_317);
nor U378 (N_378,In_475,In_363);
or U379 (N_379,In_171,In_412);
or U380 (N_380,In_434,In_49);
and U381 (N_381,In_427,In_342);
nor U382 (N_382,In_395,In_19);
and U383 (N_383,In_161,In_439);
nor U384 (N_384,In_91,In_98);
nand U385 (N_385,In_63,In_492);
nand U386 (N_386,In_207,In_283);
and U387 (N_387,In_428,In_330);
nor U388 (N_388,In_85,In_194);
nor U389 (N_389,In_44,In_380);
nor U390 (N_390,In_227,In_443);
nor U391 (N_391,In_167,In_372);
and U392 (N_392,In_426,In_420);
nor U393 (N_393,In_213,In_388);
nor U394 (N_394,In_165,In_7);
nand U395 (N_395,In_308,In_213);
or U396 (N_396,In_380,In_253);
nand U397 (N_397,In_434,In_395);
and U398 (N_398,In_202,In_304);
nand U399 (N_399,In_409,In_257);
nor U400 (N_400,In_171,In_68);
nand U401 (N_401,In_16,In_377);
and U402 (N_402,In_38,In_269);
or U403 (N_403,In_310,In_389);
or U404 (N_404,In_237,In_131);
or U405 (N_405,In_139,In_167);
xor U406 (N_406,In_156,In_218);
nor U407 (N_407,In_26,In_386);
nor U408 (N_408,In_54,In_405);
and U409 (N_409,In_163,In_127);
nor U410 (N_410,In_142,In_26);
nor U411 (N_411,In_362,In_485);
nand U412 (N_412,In_305,In_96);
nor U413 (N_413,In_202,In_421);
or U414 (N_414,In_233,In_413);
and U415 (N_415,In_465,In_308);
nand U416 (N_416,In_164,In_285);
and U417 (N_417,In_474,In_410);
nand U418 (N_418,In_391,In_322);
nor U419 (N_419,In_247,In_243);
or U420 (N_420,In_114,In_298);
nand U421 (N_421,In_303,In_444);
nand U422 (N_422,In_111,In_168);
nand U423 (N_423,In_134,In_182);
nand U424 (N_424,In_421,In_426);
xor U425 (N_425,In_100,In_336);
nand U426 (N_426,In_477,In_436);
and U427 (N_427,In_114,In_167);
nand U428 (N_428,In_339,In_186);
nor U429 (N_429,In_498,In_362);
nand U430 (N_430,In_234,In_176);
or U431 (N_431,In_53,In_139);
nor U432 (N_432,In_293,In_72);
or U433 (N_433,In_455,In_410);
nand U434 (N_434,In_83,In_29);
or U435 (N_435,In_242,In_328);
and U436 (N_436,In_122,In_217);
nor U437 (N_437,In_118,In_156);
nand U438 (N_438,In_344,In_191);
nand U439 (N_439,In_203,In_67);
nand U440 (N_440,In_358,In_373);
nor U441 (N_441,In_369,In_485);
nand U442 (N_442,In_471,In_189);
and U443 (N_443,In_438,In_123);
and U444 (N_444,In_71,In_414);
xor U445 (N_445,In_397,In_491);
nor U446 (N_446,In_44,In_435);
nand U447 (N_447,In_464,In_334);
nor U448 (N_448,In_313,In_285);
nor U449 (N_449,In_322,In_455);
or U450 (N_450,In_125,In_244);
or U451 (N_451,In_279,In_243);
xnor U452 (N_452,In_129,In_303);
and U453 (N_453,In_41,In_254);
nand U454 (N_454,In_147,In_362);
or U455 (N_455,In_309,In_257);
xnor U456 (N_456,In_390,In_266);
or U457 (N_457,In_54,In_156);
or U458 (N_458,In_116,In_403);
or U459 (N_459,In_496,In_123);
xor U460 (N_460,In_334,In_51);
nor U461 (N_461,In_315,In_77);
or U462 (N_462,In_305,In_238);
nor U463 (N_463,In_374,In_76);
and U464 (N_464,In_203,In_422);
nand U465 (N_465,In_323,In_70);
and U466 (N_466,In_370,In_165);
nor U467 (N_467,In_74,In_307);
nor U468 (N_468,In_113,In_18);
nand U469 (N_469,In_315,In_142);
or U470 (N_470,In_166,In_386);
and U471 (N_471,In_210,In_346);
and U472 (N_472,In_136,In_192);
nor U473 (N_473,In_239,In_5);
and U474 (N_474,In_448,In_416);
and U475 (N_475,In_41,In_299);
nand U476 (N_476,In_295,In_141);
or U477 (N_477,In_152,In_325);
nand U478 (N_478,In_170,In_76);
nor U479 (N_479,In_207,In_295);
and U480 (N_480,In_166,In_448);
and U481 (N_481,In_179,In_303);
xnor U482 (N_482,In_216,In_492);
nand U483 (N_483,In_75,In_250);
and U484 (N_484,In_331,In_39);
nor U485 (N_485,In_250,In_484);
or U486 (N_486,In_407,In_248);
and U487 (N_487,In_13,In_76);
nand U488 (N_488,In_317,In_170);
or U489 (N_489,In_200,In_458);
xnor U490 (N_490,In_473,In_45);
and U491 (N_491,In_243,In_338);
nor U492 (N_492,In_484,In_497);
or U493 (N_493,In_452,In_200);
nand U494 (N_494,In_319,In_25);
and U495 (N_495,In_129,In_265);
nor U496 (N_496,In_358,In_344);
or U497 (N_497,In_276,In_50);
nand U498 (N_498,In_94,In_393);
nor U499 (N_499,In_440,In_324);
nand U500 (N_500,In_479,In_267);
nand U501 (N_501,In_37,In_22);
or U502 (N_502,In_50,In_14);
nand U503 (N_503,In_413,In_151);
nor U504 (N_504,In_409,In_295);
and U505 (N_505,In_491,In_77);
and U506 (N_506,In_151,In_294);
or U507 (N_507,In_412,In_229);
nand U508 (N_508,In_98,In_421);
nor U509 (N_509,In_160,In_43);
nor U510 (N_510,In_496,In_278);
or U511 (N_511,In_127,In_128);
nand U512 (N_512,In_238,In_404);
and U513 (N_513,In_89,In_73);
and U514 (N_514,In_187,In_284);
or U515 (N_515,In_146,In_64);
nor U516 (N_516,In_147,In_327);
and U517 (N_517,In_177,In_354);
nor U518 (N_518,In_162,In_3);
or U519 (N_519,In_275,In_125);
and U520 (N_520,In_215,In_290);
nor U521 (N_521,In_248,In_300);
nor U522 (N_522,In_239,In_343);
or U523 (N_523,In_318,In_330);
nor U524 (N_524,In_173,In_234);
and U525 (N_525,In_112,In_430);
or U526 (N_526,In_393,In_9);
nor U527 (N_527,In_346,In_97);
nor U528 (N_528,In_359,In_131);
and U529 (N_529,In_399,In_150);
nand U530 (N_530,In_348,In_328);
nand U531 (N_531,In_170,In_23);
nand U532 (N_532,In_200,In_389);
nand U533 (N_533,In_301,In_244);
nor U534 (N_534,In_7,In_146);
nand U535 (N_535,In_360,In_484);
nand U536 (N_536,In_133,In_33);
or U537 (N_537,In_131,In_415);
nor U538 (N_538,In_49,In_56);
or U539 (N_539,In_202,In_151);
and U540 (N_540,In_287,In_473);
xor U541 (N_541,In_322,In_373);
nand U542 (N_542,In_36,In_367);
and U543 (N_543,In_16,In_125);
nand U544 (N_544,In_276,In_460);
and U545 (N_545,In_460,In_96);
and U546 (N_546,In_435,In_377);
nor U547 (N_547,In_235,In_432);
nand U548 (N_548,In_114,In_170);
nand U549 (N_549,In_470,In_51);
or U550 (N_550,In_18,In_150);
xor U551 (N_551,In_10,In_323);
nor U552 (N_552,In_31,In_442);
or U553 (N_553,In_171,In_490);
and U554 (N_554,In_179,In_401);
nand U555 (N_555,In_468,In_273);
and U556 (N_556,In_175,In_230);
nor U557 (N_557,In_327,In_431);
nor U558 (N_558,In_475,In_406);
nand U559 (N_559,In_265,In_312);
nand U560 (N_560,In_147,In_128);
nand U561 (N_561,In_62,In_246);
or U562 (N_562,In_297,In_283);
and U563 (N_563,In_154,In_492);
and U564 (N_564,In_128,In_386);
or U565 (N_565,In_447,In_466);
and U566 (N_566,In_398,In_464);
nand U567 (N_567,In_369,In_187);
nand U568 (N_568,In_7,In_424);
and U569 (N_569,In_336,In_422);
or U570 (N_570,In_338,In_301);
or U571 (N_571,In_244,In_44);
and U572 (N_572,In_403,In_392);
and U573 (N_573,In_110,In_199);
and U574 (N_574,In_483,In_144);
or U575 (N_575,In_211,In_203);
or U576 (N_576,In_33,In_239);
nand U577 (N_577,In_342,In_478);
or U578 (N_578,In_266,In_165);
nand U579 (N_579,In_80,In_303);
nor U580 (N_580,In_274,In_359);
nand U581 (N_581,In_181,In_7);
nand U582 (N_582,In_83,In_154);
and U583 (N_583,In_183,In_292);
or U584 (N_584,In_409,In_486);
nor U585 (N_585,In_416,In_489);
nand U586 (N_586,In_274,In_126);
and U587 (N_587,In_420,In_249);
nand U588 (N_588,In_238,In_333);
nor U589 (N_589,In_44,In_249);
or U590 (N_590,In_270,In_192);
and U591 (N_591,In_71,In_428);
nand U592 (N_592,In_447,In_272);
nand U593 (N_593,In_13,In_116);
and U594 (N_594,In_322,In_286);
nand U595 (N_595,In_239,In_242);
nand U596 (N_596,In_342,In_73);
nor U597 (N_597,In_20,In_297);
and U598 (N_598,In_155,In_224);
nand U599 (N_599,In_287,In_403);
and U600 (N_600,N_62,N_325);
or U601 (N_601,N_371,N_243);
xor U602 (N_602,N_218,N_203);
nand U603 (N_603,N_156,N_435);
and U604 (N_604,N_335,N_3);
nor U605 (N_605,N_564,N_63);
nor U606 (N_606,N_37,N_186);
or U607 (N_607,N_567,N_278);
nand U608 (N_608,N_282,N_460);
nand U609 (N_609,N_554,N_493);
nand U610 (N_610,N_254,N_94);
and U611 (N_611,N_221,N_569);
and U612 (N_612,N_195,N_78);
nor U613 (N_613,N_418,N_2);
nor U614 (N_614,N_125,N_486);
or U615 (N_615,N_369,N_303);
and U616 (N_616,N_330,N_14);
and U617 (N_617,N_134,N_197);
nor U618 (N_618,N_235,N_449);
and U619 (N_619,N_455,N_210);
nor U620 (N_620,N_531,N_226);
and U621 (N_621,N_196,N_321);
nand U622 (N_622,N_59,N_160);
nand U623 (N_623,N_273,N_92);
nor U624 (N_624,N_316,N_255);
or U625 (N_625,N_318,N_399);
nor U626 (N_626,N_523,N_236);
nand U627 (N_627,N_121,N_309);
nor U628 (N_628,N_437,N_337);
and U629 (N_629,N_154,N_495);
nand U630 (N_630,N_597,N_144);
and U631 (N_631,N_205,N_208);
and U632 (N_632,N_110,N_367);
and U633 (N_633,N_136,N_188);
and U634 (N_634,N_301,N_490);
nor U635 (N_635,N_66,N_18);
or U636 (N_636,N_485,N_185);
nor U637 (N_637,N_389,N_474);
nand U638 (N_638,N_151,N_40);
nor U639 (N_639,N_377,N_64);
or U640 (N_640,N_133,N_572);
or U641 (N_641,N_99,N_15);
or U642 (N_642,N_350,N_191);
and U643 (N_643,N_5,N_329);
nor U644 (N_644,N_406,N_122);
nor U645 (N_645,N_198,N_171);
nor U646 (N_646,N_117,N_7);
nor U647 (N_647,N_539,N_39);
and U648 (N_648,N_322,N_311);
nand U649 (N_649,N_223,N_44);
nand U650 (N_650,N_349,N_417);
nand U651 (N_651,N_155,N_428);
nor U652 (N_652,N_376,N_576);
nor U653 (N_653,N_281,N_469);
and U654 (N_654,N_147,N_300);
and U655 (N_655,N_142,N_310);
nor U656 (N_656,N_484,N_343);
nor U657 (N_657,N_542,N_512);
nand U658 (N_658,N_6,N_192);
nand U659 (N_659,N_555,N_323);
and U660 (N_660,N_585,N_28);
or U661 (N_661,N_275,N_314);
nor U662 (N_662,N_217,N_114);
or U663 (N_663,N_81,N_24);
and U664 (N_664,N_274,N_519);
and U665 (N_665,N_100,N_42);
nor U666 (N_666,N_375,N_126);
and U667 (N_667,N_279,N_283);
or U668 (N_668,N_494,N_17);
nand U669 (N_669,N_116,N_97);
or U670 (N_670,N_219,N_390);
or U671 (N_671,N_550,N_387);
nand U672 (N_672,N_295,N_527);
nor U673 (N_673,N_170,N_204);
nor U674 (N_674,N_292,N_391);
nand U675 (N_675,N_368,N_21);
or U676 (N_676,N_287,N_517);
nand U677 (N_677,N_286,N_510);
nand U678 (N_678,N_332,N_70);
nand U679 (N_679,N_194,N_556);
and U680 (N_680,N_159,N_544);
xnor U681 (N_681,N_161,N_416);
and U682 (N_682,N_294,N_241);
nor U683 (N_683,N_260,N_363);
or U684 (N_684,N_558,N_138);
xnor U685 (N_685,N_344,N_130);
nand U686 (N_686,N_73,N_302);
or U687 (N_687,N_454,N_338);
xor U688 (N_688,N_49,N_583);
nor U689 (N_689,N_384,N_423);
nand U690 (N_690,N_450,N_67);
nor U691 (N_691,N_34,N_521);
xor U692 (N_692,N_482,N_596);
xnor U693 (N_693,N_71,N_563);
nor U694 (N_694,N_380,N_361);
and U695 (N_695,N_552,N_157);
or U696 (N_696,N_489,N_187);
nand U697 (N_697,N_307,N_346);
nand U698 (N_698,N_11,N_30);
nor U699 (N_699,N_357,N_497);
nand U700 (N_700,N_320,N_16);
nand U701 (N_701,N_355,N_271);
or U702 (N_702,N_87,N_448);
or U703 (N_703,N_46,N_89);
and U704 (N_704,N_119,N_297);
nor U705 (N_705,N_127,N_465);
nand U706 (N_706,N_19,N_386);
nand U707 (N_707,N_445,N_319);
or U708 (N_708,N_143,N_20);
nor U709 (N_709,N_393,N_200);
xnor U710 (N_710,N_249,N_421);
nor U711 (N_711,N_169,N_31);
nor U712 (N_712,N_559,N_52);
or U713 (N_713,N_258,N_193);
nor U714 (N_714,N_265,N_43);
nand U715 (N_715,N_348,N_57);
and U716 (N_716,N_439,N_324);
and U717 (N_717,N_457,N_534);
or U718 (N_718,N_93,N_207);
nor U719 (N_719,N_591,N_108);
or U720 (N_720,N_545,N_408);
nor U721 (N_721,N_199,N_83);
and U722 (N_722,N_333,N_353);
nand U723 (N_723,N_22,N_85);
nand U724 (N_724,N_181,N_214);
nor U725 (N_725,N_587,N_443);
or U726 (N_726,N_296,N_586);
and U727 (N_727,N_359,N_86);
nor U728 (N_728,N_526,N_141);
or U729 (N_729,N_299,N_411);
nand U730 (N_730,N_502,N_250);
and U731 (N_731,N_268,N_543);
or U732 (N_732,N_263,N_549);
or U733 (N_733,N_464,N_269);
nand U734 (N_734,N_366,N_50);
or U735 (N_735,N_483,N_284);
or U736 (N_736,N_446,N_381);
or U737 (N_737,N_392,N_398);
and U738 (N_738,N_440,N_182);
nand U739 (N_739,N_267,N_315);
nand U740 (N_740,N_341,N_546);
nor U741 (N_741,N_364,N_209);
or U742 (N_742,N_436,N_225);
and U743 (N_743,N_475,N_277);
or U744 (N_744,N_397,N_29);
nor U745 (N_745,N_132,N_331);
or U746 (N_746,N_358,N_588);
or U747 (N_747,N_261,N_478);
and U748 (N_748,N_84,N_354);
or U749 (N_749,N_74,N_77);
or U750 (N_750,N_480,N_431);
and U751 (N_751,N_352,N_342);
nand U752 (N_752,N_266,N_491);
and U753 (N_753,N_360,N_237);
and U754 (N_754,N_153,N_470);
nand U755 (N_755,N_553,N_253);
or U756 (N_756,N_162,N_365);
and U757 (N_757,N_163,N_115);
or U758 (N_758,N_290,N_164);
nand U759 (N_759,N_202,N_405);
and U760 (N_760,N_106,N_592);
nand U761 (N_761,N_167,N_492);
nor U762 (N_762,N_538,N_75);
nand U763 (N_763,N_415,N_540);
or U764 (N_764,N_312,N_444);
or U765 (N_765,N_257,N_424);
nor U766 (N_766,N_173,N_506);
nand U767 (N_767,N_95,N_574);
and U768 (N_768,N_581,N_288);
nand U769 (N_769,N_109,N_48);
nand U770 (N_770,N_242,N_396);
and U771 (N_771,N_120,N_234);
nor U772 (N_772,N_407,N_165);
nand U773 (N_773,N_463,N_13);
nor U774 (N_774,N_180,N_272);
or U775 (N_775,N_238,N_178);
or U776 (N_776,N_533,N_479);
and U777 (N_777,N_252,N_68);
and U778 (N_778,N_579,N_370);
nor U779 (N_779,N_334,N_129);
nand U780 (N_780,N_26,N_262);
nor U781 (N_781,N_584,N_36);
xor U782 (N_782,N_378,N_224);
nand U783 (N_783,N_251,N_230);
and U784 (N_784,N_308,N_441);
or U785 (N_785,N_404,N_524);
nand U786 (N_786,N_498,N_453);
nand U787 (N_787,N_240,N_245);
nand U788 (N_788,N_211,N_433);
and U789 (N_789,N_25,N_537);
nor U790 (N_790,N_351,N_189);
or U791 (N_791,N_58,N_427);
or U792 (N_792,N_174,N_575);
or U793 (N_793,N_500,N_206);
nor U794 (N_794,N_551,N_516);
nor U795 (N_795,N_213,N_442);
nor U796 (N_796,N_327,N_520);
or U797 (N_797,N_462,N_379);
nand U798 (N_798,N_54,N_228);
nand U799 (N_799,N_566,N_91);
and U800 (N_800,N_104,N_90);
nand U801 (N_801,N_298,N_82);
or U802 (N_802,N_56,N_201);
nor U803 (N_803,N_573,N_507);
nand U804 (N_804,N_69,N_80);
and U805 (N_805,N_216,N_413);
or U806 (N_806,N_113,N_562);
and U807 (N_807,N_9,N_65);
nor U808 (N_808,N_340,N_12);
and U809 (N_809,N_179,N_471);
and U810 (N_810,N_458,N_79);
nand U811 (N_811,N_131,N_246);
or U812 (N_812,N_256,N_432);
nor U813 (N_813,N_112,N_103);
or U814 (N_814,N_326,N_313);
xor U815 (N_815,N_45,N_145);
and U816 (N_816,N_222,N_503);
or U817 (N_817,N_468,N_598);
nand U818 (N_818,N_426,N_33);
nor U819 (N_819,N_72,N_347);
and U820 (N_820,N_373,N_146);
and U821 (N_821,N_102,N_152);
and U822 (N_822,N_47,N_536);
nor U823 (N_823,N_96,N_305);
nor U824 (N_824,N_451,N_459);
or U825 (N_825,N_402,N_434);
or U826 (N_826,N_582,N_304);
nand U827 (N_827,N_425,N_403);
nand U828 (N_828,N_589,N_515);
and U829 (N_829,N_420,N_514);
or U830 (N_830,N_528,N_61);
and U831 (N_831,N_395,N_477);
and U832 (N_832,N_525,N_76);
nand U833 (N_833,N_183,N_388);
or U834 (N_834,N_577,N_55);
nand U835 (N_835,N_150,N_530);
nand U836 (N_836,N_233,N_259);
nand U837 (N_837,N_128,N_8);
nand U838 (N_838,N_247,N_101);
nand U839 (N_839,N_32,N_38);
or U840 (N_840,N_372,N_105);
or U841 (N_841,N_422,N_306);
or U842 (N_842,N_60,N_496);
nand U843 (N_843,N_1,N_362);
nor U844 (N_844,N_565,N_98);
nor U845 (N_845,N_410,N_229);
nor U846 (N_846,N_487,N_149);
nand U847 (N_847,N_476,N_509);
nor U848 (N_848,N_548,N_345);
nor U849 (N_849,N_176,N_599);
or U850 (N_850,N_289,N_231);
and U851 (N_851,N_456,N_264);
xnor U852 (N_852,N_467,N_473);
or U853 (N_853,N_560,N_0);
or U854 (N_854,N_148,N_419);
nand U855 (N_855,N_123,N_532);
and U856 (N_856,N_212,N_53);
or U857 (N_857,N_578,N_438);
and U858 (N_858,N_168,N_328);
or U859 (N_859,N_140,N_414);
and U860 (N_860,N_336,N_41);
or U861 (N_861,N_27,N_293);
or U862 (N_862,N_518,N_35);
or U863 (N_863,N_547,N_430);
nand U864 (N_864,N_374,N_190);
and U865 (N_865,N_594,N_522);
nor U866 (N_866,N_400,N_401);
and U867 (N_867,N_385,N_232);
and U868 (N_868,N_447,N_571);
nand U869 (N_869,N_124,N_175);
nand U870 (N_870,N_137,N_529);
and U871 (N_871,N_481,N_590);
nor U872 (N_872,N_383,N_317);
and U873 (N_873,N_452,N_394);
xor U874 (N_874,N_382,N_227);
or U875 (N_875,N_535,N_248);
and U876 (N_876,N_595,N_88);
or U877 (N_877,N_429,N_244);
nor U878 (N_878,N_139,N_501);
nand U879 (N_879,N_276,N_111);
and U880 (N_880,N_172,N_280);
and U881 (N_881,N_499,N_461);
and U882 (N_882,N_508,N_10);
or U883 (N_883,N_561,N_580);
and U884 (N_884,N_166,N_4);
or U885 (N_885,N_513,N_135);
or U886 (N_886,N_291,N_51);
nand U887 (N_887,N_568,N_215);
nand U888 (N_888,N_505,N_356);
nor U889 (N_889,N_466,N_339);
and U890 (N_890,N_270,N_412);
and U891 (N_891,N_541,N_158);
and U892 (N_892,N_570,N_488);
nand U893 (N_893,N_511,N_118);
nor U894 (N_894,N_239,N_504);
nor U895 (N_895,N_409,N_177);
and U896 (N_896,N_107,N_23);
nand U897 (N_897,N_472,N_285);
or U898 (N_898,N_593,N_557);
or U899 (N_899,N_220,N_184);
and U900 (N_900,N_145,N_467);
nor U901 (N_901,N_53,N_390);
nand U902 (N_902,N_195,N_520);
and U903 (N_903,N_199,N_518);
and U904 (N_904,N_287,N_290);
nor U905 (N_905,N_185,N_236);
and U906 (N_906,N_554,N_46);
or U907 (N_907,N_428,N_115);
nand U908 (N_908,N_466,N_271);
xnor U909 (N_909,N_535,N_407);
nand U910 (N_910,N_10,N_592);
and U911 (N_911,N_314,N_15);
nor U912 (N_912,N_518,N_457);
and U913 (N_913,N_498,N_193);
or U914 (N_914,N_91,N_436);
and U915 (N_915,N_334,N_53);
nor U916 (N_916,N_60,N_116);
xnor U917 (N_917,N_25,N_243);
nand U918 (N_918,N_39,N_273);
xor U919 (N_919,N_441,N_238);
and U920 (N_920,N_351,N_367);
nand U921 (N_921,N_339,N_340);
or U922 (N_922,N_336,N_365);
and U923 (N_923,N_350,N_119);
nor U924 (N_924,N_81,N_349);
nor U925 (N_925,N_481,N_586);
nand U926 (N_926,N_399,N_73);
or U927 (N_927,N_497,N_35);
nand U928 (N_928,N_259,N_479);
nor U929 (N_929,N_262,N_462);
xor U930 (N_930,N_218,N_422);
nand U931 (N_931,N_374,N_206);
and U932 (N_932,N_434,N_208);
and U933 (N_933,N_40,N_12);
or U934 (N_934,N_201,N_507);
and U935 (N_935,N_416,N_144);
or U936 (N_936,N_109,N_266);
nand U937 (N_937,N_145,N_300);
nand U938 (N_938,N_67,N_378);
nand U939 (N_939,N_562,N_306);
and U940 (N_940,N_239,N_329);
nor U941 (N_941,N_147,N_67);
nor U942 (N_942,N_367,N_67);
nor U943 (N_943,N_435,N_99);
or U944 (N_944,N_47,N_483);
nor U945 (N_945,N_51,N_513);
or U946 (N_946,N_353,N_2);
nand U947 (N_947,N_157,N_154);
nand U948 (N_948,N_65,N_586);
xnor U949 (N_949,N_503,N_152);
nand U950 (N_950,N_229,N_292);
or U951 (N_951,N_189,N_212);
nand U952 (N_952,N_408,N_110);
nor U953 (N_953,N_573,N_365);
nand U954 (N_954,N_440,N_273);
or U955 (N_955,N_530,N_15);
or U956 (N_956,N_125,N_387);
nor U957 (N_957,N_398,N_117);
or U958 (N_958,N_162,N_97);
nand U959 (N_959,N_112,N_462);
nand U960 (N_960,N_115,N_443);
and U961 (N_961,N_592,N_217);
or U962 (N_962,N_121,N_314);
or U963 (N_963,N_198,N_551);
nor U964 (N_964,N_17,N_381);
nand U965 (N_965,N_222,N_203);
and U966 (N_966,N_595,N_420);
nand U967 (N_967,N_508,N_468);
or U968 (N_968,N_524,N_6);
nand U969 (N_969,N_21,N_511);
nor U970 (N_970,N_135,N_313);
and U971 (N_971,N_119,N_69);
nand U972 (N_972,N_115,N_590);
nand U973 (N_973,N_335,N_77);
nand U974 (N_974,N_95,N_271);
or U975 (N_975,N_261,N_292);
nor U976 (N_976,N_4,N_158);
nand U977 (N_977,N_45,N_258);
or U978 (N_978,N_252,N_400);
or U979 (N_979,N_104,N_64);
nor U980 (N_980,N_131,N_284);
or U981 (N_981,N_31,N_417);
and U982 (N_982,N_401,N_182);
or U983 (N_983,N_123,N_149);
or U984 (N_984,N_155,N_580);
nor U985 (N_985,N_1,N_69);
and U986 (N_986,N_459,N_195);
or U987 (N_987,N_93,N_176);
nand U988 (N_988,N_75,N_231);
or U989 (N_989,N_52,N_326);
nor U990 (N_990,N_37,N_503);
nand U991 (N_991,N_67,N_422);
and U992 (N_992,N_85,N_562);
nor U993 (N_993,N_24,N_310);
or U994 (N_994,N_140,N_360);
or U995 (N_995,N_202,N_575);
and U996 (N_996,N_188,N_445);
or U997 (N_997,N_28,N_90);
or U998 (N_998,N_478,N_423);
and U999 (N_999,N_89,N_458);
nor U1000 (N_1000,N_277,N_29);
nor U1001 (N_1001,N_146,N_440);
and U1002 (N_1002,N_499,N_226);
nor U1003 (N_1003,N_151,N_272);
nor U1004 (N_1004,N_395,N_203);
or U1005 (N_1005,N_365,N_150);
nor U1006 (N_1006,N_265,N_47);
or U1007 (N_1007,N_376,N_310);
nor U1008 (N_1008,N_312,N_79);
and U1009 (N_1009,N_564,N_187);
nand U1010 (N_1010,N_180,N_337);
nor U1011 (N_1011,N_78,N_13);
nand U1012 (N_1012,N_489,N_318);
or U1013 (N_1013,N_496,N_587);
nor U1014 (N_1014,N_559,N_316);
or U1015 (N_1015,N_202,N_101);
or U1016 (N_1016,N_120,N_518);
or U1017 (N_1017,N_69,N_470);
nor U1018 (N_1018,N_134,N_494);
and U1019 (N_1019,N_557,N_575);
or U1020 (N_1020,N_411,N_215);
nand U1021 (N_1021,N_488,N_413);
or U1022 (N_1022,N_536,N_306);
nor U1023 (N_1023,N_438,N_293);
xor U1024 (N_1024,N_570,N_374);
and U1025 (N_1025,N_35,N_196);
xor U1026 (N_1026,N_7,N_448);
nand U1027 (N_1027,N_272,N_383);
nand U1028 (N_1028,N_30,N_274);
or U1029 (N_1029,N_35,N_267);
or U1030 (N_1030,N_538,N_173);
nor U1031 (N_1031,N_562,N_586);
nor U1032 (N_1032,N_418,N_209);
or U1033 (N_1033,N_25,N_200);
nor U1034 (N_1034,N_392,N_321);
nor U1035 (N_1035,N_184,N_86);
and U1036 (N_1036,N_70,N_397);
or U1037 (N_1037,N_397,N_142);
and U1038 (N_1038,N_30,N_363);
and U1039 (N_1039,N_291,N_581);
nand U1040 (N_1040,N_196,N_447);
and U1041 (N_1041,N_308,N_241);
and U1042 (N_1042,N_275,N_172);
or U1043 (N_1043,N_205,N_453);
or U1044 (N_1044,N_79,N_392);
nor U1045 (N_1045,N_278,N_228);
or U1046 (N_1046,N_162,N_114);
nand U1047 (N_1047,N_394,N_457);
nand U1048 (N_1048,N_255,N_438);
nor U1049 (N_1049,N_4,N_208);
nor U1050 (N_1050,N_294,N_543);
nor U1051 (N_1051,N_166,N_147);
nor U1052 (N_1052,N_532,N_135);
nor U1053 (N_1053,N_478,N_465);
and U1054 (N_1054,N_129,N_509);
or U1055 (N_1055,N_431,N_38);
nand U1056 (N_1056,N_439,N_381);
or U1057 (N_1057,N_573,N_394);
or U1058 (N_1058,N_266,N_97);
and U1059 (N_1059,N_371,N_119);
nand U1060 (N_1060,N_586,N_14);
or U1061 (N_1061,N_578,N_528);
nand U1062 (N_1062,N_305,N_213);
and U1063 (N_1063,N_392,N_34);
or U1064 (N_1064,N_140,N_366);
nor U1065 (N_1065,N_207,N_277);
and U1066 (N_1066,N_72,N_209);
and U1067 (N_1067,N_374,N_412);
or U1068 (N_1068,N_351,N_406);
nor U1069 (N_1069,N_258,N_140);
or U1070 (N_1070,N_53,N_567);
and U1071 (N_1071,N_131,N_145);
nor U1072 (N_1072,N_102,N_432);
and U1073 (N_1073,N_71,N_385);
nor U1074 (N_1074,N_537,N_393);
nand U1075 (N_1075,N_158,N_494);
nor U1076 (N_1076,N_274,N_13);
and U1077 (N_1077,N_2,N_447);
or U1078 (N_1078,N_148,N_527);
nand U1079 (N_1079,N_297,N_595);
or U1080 (N_1080,N_231,N_180);
nor U1081 (N_1081,N_128,N_223);
or U1082 (N_1082,N_117,N_433);
nand U1083 (N_1083,N_157,N_279);
nand U1084 (N_1084,N_138,N_177);
nand U1085 (N_1085,N_518,N_398);
or U1086 (N_1086,N_482,N_586);
nand U1087 (N_1087,N_18,N_95);
nor U1088 (N_1088,N_479,N_427);
or U1089 (N_1089,N_77,N_503);
or U1090 (N_1090,N_423,N_32);
nor U1091 (N_1091,N_582,N_79);
nand U1092 (N_1092,N_181,N_248);
nand U1093 (N_1093,N_169,N_468);
or U1094 (N_1094,N_576,N_233);
or U1095 (N_1095,N_172,N_334);
and U1096 (N_1096,N_589,N_177);
or U1097 (N_1097,N_29,N_592);
or U1098 (N_1098,N_254,N_314);
or U1099 (N_1099,N_181,N_324);
nor U1100 (N_1100,N_409,N_148);
and U1101 (N_1101,N_367,N_143);
and U1102 (N_1102,N_284,N_518);
or U1103 (N_1103,N_285,N_433);
nor U1104 (N_1104,N_8,N_219);
and U1105 (N_1105,N_90,N_165);
nor U1106 (N_1106,N_150,N_181);
and U1107 (N_1107,N_34,N_371);
or U1108 (N_1108,N_340,N_289);
nand U1109 (N_1109,N_241,N_1);
or U1110 (N_1110,N_317,N_265);
or U1111 (N_1111,N_480,N_49);
or U1112 (N_1112,N_121,N_490);
or U1113 (N_1113,N_260,N_304);
nand U1114 (N_1114,N_103,N_433);
nand U1115 (N_1115,N_324,N_60);
nor U1116 (N_1116,N_44,N_215);
or U1117 (N_1117,N_290,N_476);
or U1118 (N_1118,N_20,N_270);
nand U1119 (N_1119,N_22,N_78);
and U1120 (N_1120,N_400,N_269);
and U1121 (N_1121,N_433,N_112);
nor U1122 (N_1122,N_103,N_193);
and U1123 (N_1123,N_401,N_448);
or U1124 (N_1124,N_242,N_464);
nand U1125 (N_1125,N_82,N_187);
or U1126 (N_1126,N_520,N_537);
and U1127 (N_1127,N_139,N_62);
nand U1128 (N_1128,N_307,N_319);
and U1129 (N_1129,N_126,N_321);
and U1130 (N_1130,N_266,N_39);
or U1131 (N_1131,N_273,N_296);
nand U1132 (N_1132,N_372,N_299);
and U1133 (N_1133,N_142,N_157);
and U1134 (N_1134,N_345,N_429);
nand U1135 (N_1135,N_482,N_218);
or U1136 (N_1136,N_561,N_296);
nand U1137 (N_1137,N_338,N_360);
nand U1138 (N_1138,N_420,N_135);
nor U1139 (N_1139,N_307,N_334);
xnor U1140 (N_1140,N_264,N_322);
nand U1141 (N_1141,N_479,N_403);
and U1142 (N_1142,N_0,N_526);
or U1143 (N_1143,N_506,N_76);
nor U1144 (N_1144,N_354,N_489);
and U1145 (N_1145,N_282,N_190);
nand U1146 (N_1146,N_411,N_11);
nor U1147 (N_1147,N_49,N_174);
or U1148 (N_1148,N_223,N_545);
nand U1149 (N_1149,N_47,N_25);
xnor U1150 (N_1150,N_87,N_112);
or U1151 (N_1151,N_73,N_229);
nand U1152 (N_1152,N_88,N_32);
nor U1153 (N_1153,N_192,N_297);
or U1154 (N_1154,N_538,N_239);
or U1155 (N_1155,N_565,N_250);
nand U1156 (N_1156,N_586,N_351);
or U1157 (N_1157,N_284,N_419);
nor U1158 (N_1158,N_97,N_548);
and U1159 (N_1159,N_23,N_114);
nor U1160 (N_1160,N_528,N_410);
or U1161 (N_1161,N_78,N_407);
and U1162 (N_1162,N_12,N_566);
or U1163 (N_1163,N_234,N_198);
and U1164 (N_1164,N_24,N_535);
nand U1165 (N_1165,N_453,N_87);
nor U1166 (N_1166,N_276,N_424);
and U1167 (N_1167,N_529,N_131);
or U1168 (N_1168,N_475,N_583);
and U1169 (N_1169,N_438,N_360);
nor U1170 (N_1170,N_30,N_569);
and U1171 (N_1171,N_81,N_285);
or U1172 (N_1172,N_221,N_22);
or U1173 (N_1173,N_169,N_297);
and U1174 (N_1174,N_202,N_582);
and U1175 (N_1175,N_453,N_251);
nor U1176 (N_1176,N_329,N_382);
and U1177 (N_1177,N_186,N_527);
nor U1178 (N_1178,N_532,N_352);
and U1179 (N_1179,N_104,N_146);
nand U1180 (N_1180,N_572,N_29);
and U1181 (N_1181,N_374,N_429);
nor U1182 (N_1182,N_597,N_557);
xnor U1183 (N_1183,N_439,N_193);
nand U1184 (N_1184,N_217,N_344);
nand U1185 (N_1185,N_514,N_117);
and U1186 (N_1186,N_89,N_291);
and U1187 (N_1187,N_17,N_179);
and U1188 (N_1188,N_427,N_516);
nand U1189 (N_1189,N_367,N_52);
or U1190 (N_1190,N_206,N_172);
and U1191 (N_1191,N_344,N_147);
or U1192 (N_1192,N_346,N_439);
nor U1193 (N_1193,N_192,N_126);
xor U1194 (N_1194,N_253,N_213);
or U1195 (N_1195,N_323,N_110);
or U1196 (N_1196,N_298,N_365);
and U1197 (N_1197,N_196,N_267);
nand U1198 (N_1198,N_7,N_222);
nor U1199 (N_1199,N_309,N_143);
nand U1200 (N_1200,N_1132,N_778);
nor U1201 (N_1201,N_749,N_1086);
and U1202 (N_1202,N_1120,N_966);
nand U1203 (N_1203,N_787,N_738);
xor U1204 (N_1204,N_1034,N_1020);
or U1205 (N_1205,N_620,N_1139);
nand U1206 (N_1206,N_854,N_1031);
nand U1207 (N_1207,N_1138,N_970);
nor U1208 (N_1208,N_607,N_630);
or U1209 (N_1209,N_1036,N_955);
or U1210 (N_1210,N_691,N_1134);
and U1211 (N_1211,N_1012,N_818);
xnor U1212 (N_1212,N_763,N_654);
nand U1213 (N_1213,N_640,N_1094);
xnor U1214 (N_1214,N_1124,N_940);
xnor U1215 (N_1215,N_1005,N_1111);
nor U1216 (N_1216,N_884,N_781);
nor U1217 (N_1217,N_1194,N_926);
nor U1218 (N_1218,N_887,N_931);
nor U1219 (N_1219,N_1071,N_904);
nand U1220 (N_1220,N_725,N_1142);
nor U1221 (N_1221,N_605,N_776);
and U1222 (N_1222,N_706,N_711);
or U1223 (N_1223,N_1015,N_611);
nand U1224 (N_1224,N_784,N_921);
nor U1225 (N_1225,N_1079,N_1003);
nand U1226 (N_1226,N_1008,N_1114);
nor U1227 (N_1227,N_680,N_879);
nand U1228 (N_1228,N_1040,N_897);
or U1229 (N_1229,N_1144,N_855);
nand U1230 (N_1230,N_899,N_824);
and U1231 (N_1231,N_1004,N_646);
and U1232 (N_1232,N_650,N_1032);
nor U1233 (N_1233,N_658,N_1191);
nor U1234 (N_1234,N_718,N_726);
and U1235 (N_1235,N_865,N_750);
nand U1236 (N_1236,N_610,N_950);
nand U1237 (N_1237,N_746,N_1149);
or U1238 (N_1238,N_1055,N_633);
nand U1239 (N_1239,N_810,N_700);
nand U1240 (N_1240,N_1126,N_615);
or U1241 (N_1241,N_846,N_626);
nor U1242 (N_1242,N_965,N_715);
nor U1243 (N_1243,N_877,N_687);
and U1244 (N_1244,N_734,N_1123);
and U1245 (N_1245,N_668,N_869);
nor U1246 (N_1246,N_894,N_771);
nor U1247 (N_1247,N_1053,N_802);
or U1248 (N_1248,N_1076,N_934);
and U1249 (N_1249,N_624,N_1140);
or U1250 (N_1250,N_989,N_831);
nor U1251 (N_1251,N_864,N_649);
or U1252 (N_1252,N_785,N_1048);
nor U1253 (N_1253,N_914,N_881);
and U1254 (N_1254,N_696,N_883);
nor U1255 (N_1255,N_1164,N_760);
and U1256 (N_1256,N_1065,N_937);
or U1257 (N_1257,N_740,N_808);
nand U1258 (N_1258,N_975,N_1029);
nand U1259 (N_1259,N_1074,N_617);
nand U1260 (N_1260,N_983,N_948);
nor U1261 (N_1261,N_1033,N_722);
or U1262 (N_1262,N_1181,N_827);
nand U1263 (N_1263,N_839,N_666);
nand U1264 (N_1264,N_604,N_898);
and U1265 (N_1265,N_905,N_916);
nor U1266 (N_1266,N_1007,N_751);
or U1267 (N_1267,N_1168,N_920);
or U1268 (N_1268,N_856,N_803);
nand U1269 (N_1269,N_930,N_944);
nand U1270 (N_1270,N_821,N_1006);
nor U1271 (N_1271,N_1022,N_782);
and U1272 (N_1272,N_951,N_647);
nand U1273 (N_1273,N_768,N_728);
xor U1274 (N_1274,N_942,N_1150);
nor U1275 (N_1275,N_1121,N_967);
nand U1276 (N_1276,N_1063,N_878);
or U1277 (N_1277,N_848,N_999);
nor U1278 (N_1278,N_1098,N_1171);
nor U1279 (N_1279,N_952,N_1105);
and U1280 (N_1280,N_741,N_851);
or U1281 (N_1281,N_1078,N_1131);
nor U1282 (N_1282,N_789,N_713);
nor U1283 (N_1283,N_1064,N_632);
nand U1284 (N_1284,N_1070,N_912);
or U1285 (N_1285,N_835,N_608);
and U1286 (N_1286,N_699,N_621);
nor U1287 (N_1287,N_1195,N_695);
and U1288 (N_1288,N_913,N_1162);
or U1289 (N_1289,N_1185,N_1046);
nand U1290 (N_1290,N_703,N_823);
nand U1291 (N_1291,N_1147,N_843);
nand U1292 (N_1292,N_755,N_1179);
or U1293 (N_1293,N_670,N_758);
nor U1294 (N_1294,N_1002,N_797);
nand U1295 (N_1295,N_1042,N_963);
nor U1296 (N_1296,N_1092,N_659);
and U1297 (N_1297,N_1133,N_1173);
nand U1298 (N_1298,N_903,N_1192);
nand U1299 (N_1299,N_1155,N_775);
nand U1300 (N_1300,N_689,N_790);
or U1301 (N_1301,N_769,N_686);
and U1302 (N_1302,N_1082,N_1095);
or U1303 (N_1303,N_719,N_978);
and U1304 (N_1304,N_956,N_1077);
nand U1305 (N_1305,N_709,N_745);
or U1306 (N_1306,N_669,N_688);
nor U1307 (N_1307,N_1050,N_892);
nand U1308 (N_1308,N_601,N_1057);
nand U1309 (N_1309,N_932,N_836);
nor U1310 (N_1310,N_941,N_1001);
or U1311 (N_1311,N_925,N_900);
nor U1312 (N_1312,N_761,N_938);
xor U1313 (N_1313,N_623,N_1068);
xor U1314 (N_1314,N_627,N_902);
nor U1315 (N_1315,N_988,N_667);
nor U1316 (N_1316,N_643,N_794);
and U1317 (N_1317,N_795,N_1051);
or U1318 (N_1318,N_1159,N_739);
nand U1319 (N_1319,N_1027,N_862);
nor U1320 (N_1320,N_1073,N_890);
nor U1321 (N_1321,N_886,N_1136);
or U1322 (N_1322,N_716,N_1069);
or U1323 (N_1323,N_697,N_1030);
nand U1324 (N_1324,N_679,N_1058);
nand U1325 (N_1325,N_857,N_1117);
or U1326 (N_1326,N_743,N_960);
nor U1327 (N_1327,N_830,N_685);
nand U1328 (N_1328,N_1067,N_805);
and U1329 (N_1329,N_1096,N_602);
nor U1330 (N_1330,N_1160,N_662);
nor U1331 (N_1331,N_1026,N_850);
nand U1332 (N_1332,N_663,N_1148);
nand U1333 (N_1333,N_870,N_859);
and U1334 (N_1334,N_777,N_801);
nor U1335 (N_1335,N_664,N_874);
and U1336 (N_1336,N_1080,N_759);
nand U1337 (N_1337,N_655,N_733);
nor U1338 (N_1338,N_1169,N_1197);
and U1339 (N_1339,N_1128,N_765);
nor U1340 (N_1340,N_928,N_1177);
and U1341 (N_1341,N_1054,N_1125);
nand U1342 (N_1342,N_917,N_799);
nor U1343 (N_1343,N_901,N_1180);
or U1344 (N_1344,N_1024,N_815);
or U1345 (N_1345,N_858,N_683);
nand U1346 (N_1346,N_773,N_1170);
and U1347 (N_1347,N_1011,N_1175);
or U1348 (N_1348,N_677,N_705);
nand U1349 (N_1349,N_923,N_1045);
nand U1350 (N_1350,N_910,N_1104);
and U1351 (N_1351,N_653,N_652);
xnor U1352 (N_1352,N_1018,N_949);
and U1353 (N_1353,N_964,N_1059);
or U1354 (N_1354,N_729,N_1172);
nand U1355 (N_1355,N_993,N_845);
and U1356 (N_1356,N_717,N_710);
or U1357 (N_1357,N_834,N_796);
nor U1358 (N_1358,N_1044,N_701);
and U1359 (N_1359,N_698,N_863);
and U1360 (N_1360,N_994,N_1025);
nor U1361 (N_1361,N_1129,N_1178);
nor U1362 (N_1362,N_682,N_644);
nand U1363 (N_1363,N_748,N_1166);
xnor U1364 (N_1364,N_1188,N_987);
nand U1365 (N_1365,N_1112,N_958);
nand U1366 (N_1366,N_651,N_1130);
or U1367 (N_1367,N_919,N_968);
and U1368 (N_1368,N_1083,N_1107);
nand U1369 (N_1369,N_969,N_935);
and U1370 (N_1370,N_906,N_603);
nand U1371 (N_1371,N_840,N_1101);
nand U1372 (N_1372,N_806,N_723);
or U1373 (N_1373,N_1119,N_674);
nand U1374 (N_1374,N_635,N_833);
or U1375 (N_1375,N_798,N_1088);
nand U1376 (N_1376,N_1061,N_832);
nand U1377 (N_1377,N_995,N_866);
and U1378 (N_1378,N_614,N_645);
nand U1379 (N_1379,N_690,N_1081);
and U1380 (N_1380,N_816,N_754);
or U1381 (N_1381,N_1113,N_976);
and U1382 (N_1382,N_720,N_849);
and U1383 (N_1383,N_996,N_707);
and U1384 (N_1384,N_756,N_1010);
or U1385 (N_1385,N_1103,N_882);
and U1386 (N_1386,N_811,N_661);
nand U1387 (N_1387,N_1021,N_961);
or U1388 (N_1388,N_673,N_612);
xor U1389 (N_1389,N_929,N_619);
nand U1390 (N_1390,N_636,N_979);
nor U1391 (N_1391,N_998,N_731);
nand U1392 (N_1392,N_753,N_1122);
nor U1393 (N_1393,N_730,N_852);
nand U1394 (N_1394,N_984,N_939);
or U1395 (N_1395,N_671,N_986);
or U1396 (N_1396,N_1176,N_1049);
and U1397 (N_1397,N_1154,N_812);
or U1398 (N_1398,N_997,N_767);
or U1399 (N_1399,N_1151,N_957);
and U1400 (N_1400,N_954,N_860);
nor U1401 (N_1401,N_953,N_1085);
and U1402 (N_1402,N_911,N_973);
nor U1403 (N_1403,N_888,N_793);
nand U1404 (N_1404,N_762,N_712);
nor U1405 (N_1405,N_631,N_681);
or U1406 (N_1406,N_837,N_1127);
nor U1407 (N_1407,N_817,N_809);
nor U1408 (N_1408,N_1047,N_1153);
or U1409 (N_1409,N_665,N_786);
or U1410 (N_1410,N_1158,N_1198);
or U1411 (N_1411,N_628,N_1167);
nand U1412 (N_1412,N_774,N_1141);
or U1413 (N_1413,N_742,N_1099);
nand U1414 (N_1414,N_804,N_962);
nor U1415 (N_1415,N_838,N_676);
or U1416 (N_1416,N_1183,N_1187);
or U1417 (N_1417,N_873,N_1075);
nor U1418 (N_1418,N_1062,N_981);
nand U1419 (N_1419,N_1163,N_1017);
and U1420 (N_1420,N_947,N_842);
nor U1421 (N_1421,N_638,N_772);
or U1422 (N_1422,N_1090,N_724);
nand U1423 (N_1423,N_639,N_841);
nand U1424 (N_1424,N_820,N_692);
or U1425 (N_1425,N_992,N_1190);
or U1426 (N_1426,N_1087,N_972);
or U1427 (N_1427,N_1093,N_1102);
and U1428 (N_1428,N_1110,N_1115);
and U1429 (N_1429,N_684,N_828);
and U1430 (N_1430,N_946,N_945);
and U1431 (N_1431,N_1072,N_918);
nand U1432 (N_1432,N_800,N_744);
and U1433 (N_1433,N_609,N_1052);
nand U1434 (N_1434,N_1084,N_1043);
and U1435 (N_1435,N_1041,N_637);
or U1436 (N_1436,N_1035,N_844);
or U1437 (N_1437,N_985,N_927);
or U1438 (N_1438,N_737,N_1039);
or U1439 (N_1439,N_814,N_896);
nor U1440 (N_1440,N_708,N_1193);
or U1441 (N_1441,N_1089,N_829);
or U1442 (N_1442,N_885,N_732);
and U1443 (N_1443,N_694,N_788);
nand U1444 (N_1444,N_766,N_907);
and U1445 (N_1445,N_1028,N_924);
and U1446 (N_1446,N_893,N_1000);
and U1447 (N_1447,N_915,N_727);
nor U1448 (N_1448,N_895,N_1182);
xnor U1449 (N_1449,N_678,N_672);
nand U1450 (N_1450,N_922,N_959);
or U1451 (N_1451,N_1016,N_641);
nand U1452 (N_1452,N_936,N_770);
or U1453 (N_1453,N_1184,N_1143);
or U1454 (N_1454,N_622,N_1023);
nor U1455 (N_1455,N_714,N_933);
and U1456 (N_1456,N_822,N_752);
nor U1457 (N_1457,N_813,N_1109);
or U1458 (N_1458,N_1165,N_1060);
or U1459 (N_1459,N_974,N_826);
or U1460 (N_1460,N_1116,N_1100);
nand U1461 (N_1461,N_1145,N_1157);
nor U1462 (N_1462,N_1135,N_656);
nand U1463 (N_1463,N_943,N_1019);
and U1464 (N_1464,N_660,N_779);
and U1465 (N_1465,N_634,N_606);
nor U1466 (N_1466,N_1066,N_747);
and U1467 (N_1467,N_618,N_867);
nor U1468 (N_1468,N_1013,N_1038);
nand U1469 (N_1469,N_980,N_648);
or U1470 (N_1470,N_1199,N_1091);
nand U1471 (N_1471,N_704,N_693);
nor U1472 (N_1472,N_642,N_991);
nand U1473 (N_1473,N_1186,N_657);
and U1474 (N_1474,N_675,N_909);
or U1475 (N_1475,N_971,N_1161);
or U1476 (N_1476,N_853,N_1196);
nor U1477 (N_1477,N_735,N_1037);
or U1478 (N_1478,N_629,N_625);
nor U1479 (N_1479,N_889,N_891);
xor U1480 (N_1480,N_990,N_1014);
nand U1481 (N_1481,N_908,N_1106);
and U1482 (N_1482,N_880,N_807);
nand U1483 (N_1483,N_868,N_757);
and U1484 (N_1484,N_616,N_783);
or U1485 (N_1485,N_1174,N_1146);
and U1486 (N_1486,N_1156,N_1137);
and U1487 (N_1487,N_875,N_861);
nand U1488 (N_1488,N_871,N_819);
or U1489 (N_1489,N_702,N_1097);
xnor U1490 (N_1490,N_764,N_721);
and U1491 (N_1491,N_613,N_600);
nor U1492 (N_1492,N_1189,N_1118);
nor U1493 (N_1493,N_780,N_847);
or U1494 (N_1494,N_977,N_736);
nor U1495 (N_1495,N_1009,N_1152);
nand U1496 (N_1496,N_792,N_982);
nor U1497 (N_1497,N_791,N_876);
and U1498 (N_1498,N_1108,N_872);
or U1499 (N_1499,N_1056,N_825);
nor U1500 (N_1500,N_723,N_964);
nand U1501 (N_1501,N_1023,N_895);
nor U1502 (N_1502,N_783,N_685);
and U1503 (N_1503,N_1075,N_610);
and U1504 (N_1504,N_690,N_1083);
nand U1505 (N_1505,N_794,N_1016);
nand U1506 (N_1506,N_755,N_1104);
nand U1507 (N_1507,N_970,N_931);
and U1508 (N_1508,N_701,N_1145);
nand U1509 (N_1509,N_1177,N_766);
or U1510 (N_1510,N_896,N_1085);
nand U1511 (N_1511,N_812,N_647);
nand U1512 (N_1512,N_673,N_905);
and U1513 (N_1513,N_937,N_1051);
or U1514 (N_1514,N_752,N_1110);
or U1515 (N_1515,N_1199,N_619);
nor U1516 (N_1516,N_860,N_671);
or U1517 (N_1517,N_669,N_1111);
nand U1518 (N_1518,N_781,N_702);
and U1519 (N_1519,N_1016,N_686);
or U1520 (N_1520,N_1042,N_923);
and U1521 (N_1521,N_685,N_687);
and U1522 (N_1522,N_1188,N_601);
and U1523 (N_1523,N_1037,N_945);
nor U1524 (N_1524,N_1196,N_1118);
nand U1525 (N_1525,N_1094,N_980);
and U1526 (N_1526,N_708,N_1116);
nor U1527 (N_1527,N_1069,N_973);
or U1528 (N_1528,N_1150,N_932);
nand U1529 (N_1529,N_910,N_895);
nor U1530 (N_1530,N_931,N_1166);
and U1531 (N_1531,N_1069,N_938);
nor U1532 (N_1532,N_676,N_1010);
nand U1533 (N_1533,N_1034,N_995);
or U1534 (N_1534,N_1021,N_1166);
xnor U1535 (N_1535,N_786,N_1034);
or U1536 (N_1536,N_1012,N_1118);
or U1537 (N_1537,N_1152,N_1057);
and U1538 (N_1538,N_919,N_804);
nor U1539 (N_1539,N_637,N_1054);
nand U1540 (N_1540,N_1069,N_832);
or U1541 (N_1541,N_932,N_793);
nand U1542 (N_1542,N_680,N_698);
or U1543 (N_1543,N_876,N_635);
or U1544 (N_1544,N_1064,N_799);
nor U1545 (N_1545,N_951,N_1096);
and U1546 (N_1546,N_1068,N_628);
nor U1547 (N_1547,N_639,N_1071);
and U1548 (N_1548,N_616,N_872);
nor U1549 (N_1549,N_934,N_964);
and U1550 (N_1550,N_909,N_663);
and U1551 (N_1551,N_1161,N_905);
nor U1552 (N_1552,N_637,N_1124);
and U1553 (N_1553,N_861,N_1122);
or U1554 (N_1554,N_766,N_846);
xnor U1555 (N_1555,N_601,N_860);
and U1556 (N_1556,N_1173,N_776);
and U1557 (N_1557,N_705,N_1092);
nor U1558 (N_1558,N_783,N_891);
and U1559 (N_1559,N_744,N_869);
and U1560 (N_1560,N_796,N_737);
nand U1561 (N_1561,N_861,N_934);
or U1562 (N_1562,N_853,N_848);
nand U1563 (N_1563,N_1040,N_613);
nor U1564 (N_1564,N_921,N_1157);
nand U1565 (N_1565,N_1073,N_1004);
nand U1566 (N_1566,N_612,N_727);
and U1567 (N_1567,N_662,N_603);
or U1568 (N_1568,N_1045,N_628);
and U1569 (N_1569,N_720,N_1108);
nor U1570 (N_1570,N_902,N_724);
nand U1571 (N_1571,N_1076,N_688);
nor U1572 (N_1572,N_1013,N_1153);
nand U1573 (N_1573,N_869,N_754);
nand U1574 (N_1574,N_1010,N_1095);
or U1575 (N_1575,N_1030,N_1047);
nor U1576 (N_1576,N_777,N_804);
and U1577 (N_1577,N_715,N_733);
and U1578 (N_1578,N_838,N_1100);
nand U1579 (N_1579,N_662,N_1131);
and U1580 (N_1580,N_1192,N_777);
and U1581 (N_1581,N_779,N_902);
and U1582 (N_1582,N_1131,N_626);
nand U1583 (N_1583,N_936,N_634);
nand U1584 (N_1584,N_1161,N_791);
and U1585 (N_1585,N_949,N_1107);
nand U1586 (N_1586,N_1168,N_944);
or U1587 (N_1587,N_1135,N_1061);
or U1588 (N_1588,N_723,N_866);
nor U1589 (N_1589,N_1123,N_1138);
or U1590 (N_1590,N_1122,N_1139);
nand U1591 (N_1591,N_939,N_750);
or U1592 (N_1592,N_914,N_707);
or U1593 (N_1593,N_1151,N_948);
or U1594 (N_1594,N_997,N_991);
nand U1595 (N_1595,N_1067,N_781);
or U1596 (N_1596,N_884,N_876);
or U1597 (N_1597,N_994,N_1090);
nor U1598 (N_1598,N_960,N_803);
or U1599 (N_1599,N_1001,N_720);
and U1600 (N_1600,N_885,N_797);
xnor U1601 (N_1601,N_1090,N_632);
nand U1602 (N_1602,N_869,N_686);
nor U1603 (N_1603,N_715,N_735);
nand U1604 (N_1604,N_799,N_866);
or U1605 (N_1605,N_842,N_1195);
nor U1606 (N_1606,N_748,N_1029);
or U1607 (N_1607,N_861,N_809);
nor U1608 (N_1608,N_900,N_918);
nor U1609 (N_1609,N_923,N_681);
nor U1610 (N_1610,N_1015,N_1116);
and U1611 (N_1611,N_804,N_958);
or U1612 (N_1612,N_674,N_939);
xnor U1613 (N_1613,N_1019,N_691);
nor U1614 (N_1614,N_614,N_797);
nor U1615 (N_1615,N_934,N_1188);
or U1616 (N_1616,N_1003,N_733);
nor U1617 (N_1617,N_755,N_891);
nor U1618 (N_1618,N_751,N_1000);
and U1619 (N_1619,N_1011,N_1055);
nand U1620 (N_1620,N_899,N_768);
nand U1621 (N_1621,N_1020,N_655);
and U1622 (N_1622,N_844,N_1142);
or U1623 (N_1623,N_889,N_1092);
or U1624 (N_1624,N_847,N_613);
nor U1625 (N_1625,N_1031,N_628);
or U1626 (N_1626,N_1104,N_800);
or U1627 (N_1627,N_764,N_993);
nand U1628 (N_1628,N_981,N_1060);
and U1629 (N_1629,N_730,N_1193);
nand U1630 (N_1630,N_901,N_666);
or U1631 (N_1631,N_1185,N_955);
or U1632 (N_1632,N_1029,N_611);
and U1633 (N_1633,N_1150,N_1137);
or U1634 (N_1634,N_823,N_926);
nor U1635 (N_1635,N_757,N_1066);
and U1636 (N_1636,N_1112,N_690);
and U1637 (N_1637,N_1176,N_1037);
and U1638 (N_1638,N_1111,N_1035);
and U1639 (N_1639,N_769,N_914);
nor U1640 (N_1640,N_1158,N_1097);
nor U1641 (N_1641,N_922,N_886);
nor U1642 (N_1642,N_1004,N_738);
or U1643 (N_1643,N_817,N_1154);
nor U1644 (N_1644,N_1091,N_1189);
nand U1645 (N_1645,N_1185,N_755);
or U1646 (N_1646,N_741,N_1019);
and U1647 (N_1647,N_611,N_1005);
xor U1648 (N_1648,N_1037,N_1050);
nor U1649 (N_1649,N_727,N_773);
nand U1650 (N_1650,N_1068,N_670);
and U1651 (N_1651,N_672,N_1127);
and U1652 (N_1652,N_1163,N_1180);
and U1653 (N_1653,N_882,N_1025);
nand U1654 (N_1654,N_979,N_1132);
and U1655 (N_1655,N_634,N_886);
nor U1656 (N_1656,N_1049,N_765);
nand U1657 (N_1657,N_710,N_1067);
and U1658 (N_1658,N_1061,N_987);
xor U1659 (N_1659,N_906,N_994);
nor U1660 (N_1660,N_876,N_1104);
nor U1661 (N_1661,N_1161,N_605);
or U1662 (N_1662,N_843,N_723);
nor U1663 (N_1663,N_1155,N_676);
nand U1664 (N_1664,N_1129,N_1168);
or U1665 (N_1665,N_819,N_794);
nor U1666 (N_1666,N_1034,N_1196);
nand U1667 (N_1667,N_1139,N_1164);
nand U1668 (N_1668,N_789,N_777);
or U1669 (N_1669,N_1051,N_1176);
xor U1670 (N_1670,N_1062,N_866);
nor U1671 (N_1671,N_871,N_996);
and U1672 (N_1672,N_884,N_618);
or U1673 (N_1673,N_1149,N_858);
and U1674 (N_1674,N_1196,N_1172);
nand U1675 (N_1675,N_1165,N_997);
nand U1676 (N_1676,N_878,N_1023);
nand U1677 (N_1677,N_696,N_1169);
nand U1678 (N_1678,N_1155,N_1062);
nor U1679 (N_1679,N_862,N_1094);
nand U1680 (N_1680,N_973,N_1095);
xor U1681 (N_1681,N_1165,N_943);
or U1682 (N_1682,N_1086,N_699);
and U1683 (N_1683,N_745,N_825);
nor U1684 (N_1684,N_932,N_902);
or U1685 (N_1685,N_1030,N_1100);
or U1686 (N_1686,N_791,N_1109);
xnor U1687 (N_1687,N_1179,N_905);
or U1688 (N_1688,N_705,N_949);
and U1689 (N_1689,N_983,N_903);
or U1690 (N_1690,N_1031,N_647);
and U1691 (N_1691,N_752,N_986);
and U1692 (N_1692,N_1145,N_815);
xnor U1693 (N_1693,N_931,N_747);
or U1694 (N_1694,N_771,N_1163);
nor U1695 (N_1695,N_697,N_742);
nand U1696 (N_1696,N_672,N_1139);
nor U1697 (N_1697,N_634,N_909);
nor U1698 (N_1698,N_811,N_721);
xnor U1699 (N_1699,N_1156,N_650);
nor U1700 (N_1700,N_1169,N_616);
nor U1701 (N_1701,N_839,N_713);
nand U1702 (N_1702,N_762,N_931);
nor U1703 (N_1703,N_1027,N_744);
and U1704 (N_1704,N_645,N_904);
or U1705 (N_1705,N_846,N_1145);
nand U1706 (N_1706,N_832,N_1032);
and U1707 (N_1707,N_971,N_1148);
nor U1708 (N_1708,N_814,N_627);
or U1709 (N_1709,N_1031,N_829);
and U1710 (N_1710,N_751,N_1166);
nor U1711 (N_1711,N_707,N_773);
or U1712 (N_1712,N_669,N_676);
nor U1713 (N_1713,N_922,N_621);
and U1714 (N_1714,N_948,N_1071);
nor U1715 (N_1715,N_1143,N_1004);
nor U1716 (N_1716,N_616,N_1142);
and U1717 (N_1717,N_1160,N_813);
nand U1718 (N_1718,N_724,N_1154);
nand U1719 (N_1719,N_714,N_800);
nor U1720 (N_1720,N_1070,N_814);
nand U1721 (N_1721,N_781,N_1180);
and U1722 (N_1722,N_1044,N_862);
or U1723 (N_1723,N_602,N_1174);
nor U1724 (N_1724,N_786,N_848);
and U1725 (N_1725,N_1054,N_729);
nor U1726 (N_1726,N_829,N_682);
nor U1727 (N_1727,N_962,N_1172);
nor U1728 (N_1728,N_600,N_687);
and U1729 (N_1729,N_982,N_743);
or U1730 (N_1730,N_834,N_1102);
or U1731 (N_1731,N_730,N_832);
nand U1732 (N_1732,N_1094,N_1057);
nand U1733 (N_1733,N_946,N_1190);
or U1734 (N_1734,N_920,N_884);
nor U1735 (N_1735,N_780,N_705);
and U1736 (N_1736,N_861,N_999);
and U1737 (N_1737,N_758,N_1089);
and U1738 (N_1738,N_669,N_989);
or U1739 (N_1739,N_692,N_633);
or U1740 (N_1740,N_877,N_1103);
or U1741 (N_1741,N_674,N_637);
nor U1742 (N_1742,N_771,N_1048);
and U1743 (N_1743,N_1055,N_643);
nor U1744 (N_1744,N_1013,N_1129);
or U1745 (N_1745,N_1094,N_1145);
nor U1746 (N_1746,N_842,N_837);
or U1747 (N_1747,N_1027,N_753);
or U1748 (N_1748,N_762,N_960);
and U1749 (N_1749,N_707,N_927);
and U1750 (N_1750,N_961,N_1173);
nor U1751 (N_1751,N_780,N_870);
nand U1752 (N_1752,N_772,N_1152);
or U1753 (N_1753,N_1087,N_1083);
nand U1754 (N_1754,N_832,N_851);
and U1755 (N_1755,N_925,N_604);
or U1756 (N_1756,N_677,N_805);
or U1757 (N_1757,N_1179,N_803);
or U1758 (N_1758,N_612,N_926);
nor U1759 (N_1759,N_1063,N_800);
or U1760 (N_1760,N_1189,N_607);
xnor U1761 (N_1761,N_704,N_835);
and U1762 (N_1762,N_1168,N_829);
and U1763 (N_1763,N_722,N_1056);
nor U1764 (N_1764,N_812,N_686);
or U1765 (N_1765,N_806,N_1008);
nand U1766 (N_1766,N_1100,N_822);
and U1767 (N_1767,N_722,N_1164);
nor U1768 (N_1768,N_1012,N_946);
nor U1769 (N_1769,N_1134,N_613);
or U1770 (N_1770,N_730,N_985);
nand U1771 (N_1771,N_696,N_1089);
nand U1772 (N_1772,N_761,N_1004);
and U1773 (N_1773,N_748,N_1099);
nor U1774 (N_1774,N_983,N_1027);
and U1775 (N_1775,N_802,N_1177);
or U1776 (N_1776,N_826,N_737);
nand U1777 (N_1777,N_1153,N_895);
nor U1778 (N_1778,N_880,N_922);
and U1779 (N_1779,N_663,N_1157);
nor U1780 (N_1780,N_1090,N_1076);
and U1781 (N_1781,N_1193,N_677);
nand U1782 (N_1782,N_1052,N_1146);
nor U1783 (N_1783,N_888,N_1048);
nand U1784 (N_1784,N_1092,N_1173);
nand U1785 (N_1785,N_764,N_883);
nor U1786 (N_1786,N_975,N_1112);
and U1787 (N_1787,N_1093,N_978);
nand U1788 (N_1788,N_649,N_741);
nor U1789 (N_1789,N_1032,N_1104);
and U1790 (N_1790,N_1049,N_1156);
nor U1791 (N_1791,N_1125,N_1090);
or U1792 (N_1792,N_691,N_866);
and U1793 (N_1793,N_854,N_944);
nand U1794 (N_1794,N_1133,N_931);
nand U1795 (N_1795,N_873,N_630);
or U1796 (N_1796,N_1146,N_926);
and U1797 (N_1797,N_965,N_857);
or U1798 (N_1798,N_765,N_942);
or U1799 (N_1799,N_770,N_960);
and U1800 (N_1800,N_1330,N_1228);
and U1801 (N_1801,N_1664,N_1625);
and U1802 (N_1802,N_1491,N_1763);
or U1803 (N_1803,N_1390,N_1743);
or U1804 (N_1804,N_1547,N_1518);
or U1805 (N_1805,N_1497,N_1787);
and U1806 (N_1806,N_1741,N_1509);
or U1807 (N_1807,N_1654,N_1736);
or U1808 (N_1808,N_1663,N_1474);
nand U1809 (N_1809,N_1325,N_1733);
nand U1810 (N_1810,N_1519,N_1289);
or U1811 (N_1811,N_1582,N_1363);
or U1812 (N_1812,N_1710,N_1404);
nor U1813 (N_1813,N_1453,N_1378);
nand U1814 (N_1814,N_1515,N_1340);
or U1815 (N_1815,N_1224,N_1521);
nand U1816 (N_1816,N_1621,N_1255);
nor U1817 (N_1817,N_1237,N_1308);
nor U1818 (N_1818,N_1788,N_1797);
or U1819 (N_1819,N_1775,N_1220);
nor U1820 (N_1820,N_1760,N_1600);
nor U1821 (N_1821,N_1402,N_1719);
and U1822 (N_1822,N_1571,N_1717);
xor U1823 (N_1823,N_1370,N_1494);
and U1824 (N_1824,N_1799,N_1245);
nand U1825 (N_1825,N_1752,N_1534);
and U1826 (N_1826,N_1414,N_1688);
or U1827 (N_1827,N_1704,N_1669);
nor U1828 (N_1828,N_1352,N_1498);
nand U1829 (N_1829,N_1400,N_1606);
nor U1830 (N_1830,N_1348,N_1268);
or U1831 (N_1831,N_1292,N_1681);
nand U1832 (N_1832,N_1619,N_1326);
nor U1833 (N_1833,N_1631,N_1251);
and U1834 (N_1834,N_1342,N_1336);
xor U1835 (N_1835,N_1248,N_1304);
nor U1836 (N_1836,N_1589,N_1581);
nand U1837 (N_1837,N_1495,N_1371);
xor U1838 (N_1838,N_1607,N_1670);
nand U1839 (N_1839,N_1761,N_1679);
and U1840 (N_1840,N_1266,N_1791);
nand U1841 (N_1841,N_1381,N_1332);
or U1842 (N_1842,N_1367,N_1707);
nand U1843 (N_1843,N_1483,N_1529);
and U1844 (N_1844,N_1323,N_1272);
nand U1845 (N_1845,N_1240,N_1588);
nand U1846 (N_1846,N_1629,N_1662);
nor U1847 (N_1847,N_1290,N_1790);
nand U1848 (N_1848,N_1299,N_1466);
and U1849 (N_1849,N_1723,N_1243);
nand U1850 (N_1850,N_1481,N_1226);
or U1851 (N_1851,N_1208,N_1559);
nor U1852 (N_1852,N_1410,N_1614);
or U1853 (N_1853,N_1744,N_1615);
nand U1854 (N_1854,N_1555,N_1227);
nand U1855 (N_1855,N_1746,N_1617);
nor U1856 (N_1856,N_1257,N_1201);
nor U1857 (N_1857,N_1409,N_1317);
nor U1858 (N_1858,N_1734,N_1722);
nor U1859 (N_1859,N_1644,N_1278);
and U1860 (N_1860,N_1527,N_1433);
nand U1861 (N_1861,N_1469,N_1305);
nor U1862 (N_1862,N_1210,N_1673);
nand U1863 (N_1863,N_1467,N_1503);
nand U1864 (N_1864,N_1449,N_1658);
nor U1865 (N_1865,N_1238,N_1471);
and U1866 (N_1866,N_1680,N_1270);
or U1867 (N_1867,N_1488,N_1353);
and U1868 (N_1868,N_1484,N_1345);
nand U1869 (N_1869,N_1458,N_1705);
nor U1870 (N_1870,N_1451,N_1781);
and U1871 (N_1871,N_1701,N_1375);
or U1872 (N_1872,N_1700,N_1379);
nor U1873 (N_1873,N_1568,N_1319);
or U1874 (N_1874,N_1321,N_1429);
or U1875 (N_1875,N_1695,N_1421);
nand U1876 (N_1876,N_1706,N_1630);
nor U1877 (N_1877,N_1398,N_1362);
or U1878 (N_1878,N_1464,N_1612);
and U1879 (N_1879,N_1261,N_1508);
or U1880 (N_1880,N_1372,N_1230);
nor U1881 (N_1881,N_1649,N_1253);
or U1882 (N_1882,N_1528,N_1496);
or U1883 (N_1883,N_1768,N_1720);
and U1884 (N_1884,N_1616,N_1712);
and U1885 (N_1885,N_1597,N_1206);
nor U1886 (N_1886,N_1563,N_1611);
or U1887 (N_1887,N_1287,N_1737);
nor U1888 (N_1888,N_1748,N_1273);
nor U1889 (N_1889,N_1213,N_1252);
xor U1890 (N_1890,N_1401,N_1728);
nor U1891 (N_1891,N_1640,N_1281);
and U1892 (N_1892,N_1215,N_1329);
xor U1893 (N_1893,N_1694,N_1267);
nor U1894 (N_1894,N_1393,N_1553);
or U1895 (N_1895,N_1526,N_1396);
nor U1896 (N_1896,N_1641,N_1324);
and U1897 (N_1897,N_1794,N_1338);
and U1898 (N_1898,N_1279,N_1301);
and U1899 (N_1899,N_1460,N_1485);
nand U1900 (N_1900,N_1558,N_1686);
or U1901 (N_1901,N_1668,N_1575);
or U1902 (N_1902,N_1277,N_1373);
nand U1903 (N_1903,N_1356,N_1677);
and U1904 (N_1904,N_1718,N_1294);
nor U1905 (N_1905,N_1351,N_1693);
and U1906 (N_1906,N_1647,N_1260);
or U1907 (N_1907,N_1387,N_1523);
nand U1908 (N_1908,N_1696,N_1740);
and U1909 (N_1909,N_1365,N_1595);
nand U1910 (N_1910,N_1546,N_1234);
nand U1911 (N_1911,N_1296,N_1542);
and U1912 (N_1912,N_1377,N_1275);
nand U1913 (N_1913,N_1507,N_1425);
or U1914 (N_1914,N_1535,N_1236);
nand U1915 (N_1915,N_1666,N_1209);
and U1916 (N_1916,N_1682,N_1514);
and U1917 (N_1917,N_1417,N_1572);
and U1918 (N_1918,N_1730,N_1388);
nor U1919 (N_1919,N_1601,N_1544);
nor U1920 (N_1920,N_1359,N_1759);
and U1921 (N_1921,N_1415,N_1477);
nand U1922 (N_1922,N_1636,N_1231);
or U1923 (N_1923,N_1239,N_1754);
nand U1924 (N_1924,N_1620,N_1276);
nand U1925 (N_1925,N_1347,N_1697);
nand U1926 (N_1926,N_1422,N_1506);
or U1927 (N_1927,N_1316,N_1739);
nor U1928 (N_1928,N_1298,N_1596);
and U1929 (N_1929,N_1357,N_1328);
and U1930 (N_1930,N_1235,N_1403);
or U1931 (N_1931,N_1628,N_1386);
or U1932 (N_1932,N_1242,N_1432);
nor U1933 (N_1933,N_1532,N_1713);
nor U1934 (N_1934,N_1786,N_1282);
xor U1935 (N_1935,N_1285,N_1436);
nor U1936 (N_1936,N_1447,N_1397);
nor U1937 (N_1937,N_1702,N_1703);
nor U1938 (N_1938,N_1566,N_1205);
nand U1939 (N_1939,N_1286,N_1511);
nand U1940 (N_1940,N_1557,N_1594);
or U1941 (N_1941,N_1627,N_1764);
and U1942 (N_1942,N_1750,N_1510);
nand U1943 (N_1943,N_1683,N_1309);
and U1944 (N_1944,N_1776,N_1556);
nand U1945 (N_1945,N_1691,N_1455);
nor U1946 (N_1946,N_1318,N_1490);
nand U1947 (N_1947,N_1747,N_1709);
and U1948 (N_1948,N_1531,N_1462);
nand U1949 (N_1949,N_1366,N_1653);
or U1950 (N_1950,N_1525,N_1618);
and U1951 (N_1951,N_1549,N_1214);
nand U1952 (N_1952,N_1633,N_1598);
or U1953 (N_1953,N_1283,N_1482);
nor U1954 (N_1954,N_1755,N_1771);
or U1955 (N_1955,N_1470,N_1376);
nor U1956 (N_1956,N_1424,N_1445);
or U1957 (N_1957,N_1465,N_1420);
and U1958 (N_1958,N_1576,N_1322);
nor U1959 (N_1959,N_1711,N_1291);
and U1960 (N_1960,N_1284,N_1602);
and U1961 (N_1961,N_1554,N_1479);
xor U1962 (N_1962,N_1431,N_1461);
nand U1963 (N_1963,N_1419,N_1655);
nor U1964 (N_1964,N_1623,N_1346);
nor U1965 (N_1965,N_1335,N_1472);
nor U1966 (N_1966,N_1729,N_1590);
and U1967 (N_1967,N_1573,N_1492);
and U1968 (N_1968,N_1341,N_1624);
and U1969 (N_1969,N_1232,N_1217);
and U1970 (N_1970,N_1473,N_1605);
nor U1971 (N_1971,N_1692,N_1293);
nor U1972 (N_1972,N_1638,N_1533);
or U1973 (N_1973,N_1721,N_1468);
nor U1974 (N_1974,N_1676,N_1463);
or U1975 (N_1975,N_1650,N_1726);
or U1976 (N_1976,N_1603,N_1574);
and U1977 (N_1977,N_1349,N_1307);
and U1978 (N_1978,N_1735,N_1263);
or U1979 (N_1979,N_1541,N_1264);
and U1980 (N_1980,N_1408,N_1334);
and U1981 (N_1981,N_1225,N_1350);
nand U1982 (N_1982,N_1500,N_1698);
or U1983 (N_1983,N_1552,N_1667);
or U1984 (N_1984,N_1203,N_1502);
and U1985 (N_1985,N_1678,N_1756);
nor U1986 (N_1986,N_1265,N_1580);
or U1987 (N_1987,N_1459,N_1312);
or U1988 (N_1988,N_1407,N_1383);
and U1989 (N_1989,N_1758,N_1774);
nor U1990 (N_1990,N_1586,N_1779);
nand U1991 (N_1991,N_1648,N_1592);
nand U1992 (N_1992,N_1297,N_1643);
xnor U1993 (N_1993,N_1565,N_1645);
or U1994 (N_1994,N_1456,N_1395);
nand U1995 (N_1995,N_1274,N_1742);
and U1996 (N_1996,N_1689,N_1331);
nor U1997 (N_1997,N_1499,N_1646);
nand U1998 (N_1998,N_1548,N_1657);
or U1999 (N_1999,N_1738,N_1724);
nand U2000 (N_2000,N_1249,N_1480);
and U2001 (N_2001,N_1785,N_1344);
or U2002 (N_2002,N_1651,N_1604);
or U2003 (N_2003,N_1584,N_1457);
and U2004 (N_2004,N_1295,N_1577);
and U2005 (N_2005,N_1725,N_1765);
or U2006 (N_2006,N_1212,N_1382);
nand U2007 (N_2007,N_1258,N_1652);
and U2008 (N_2008,N_1418,N_1306);
and U2009 (N_2009,N_1454,N_1536);
or U2010 (N_2010,N_1504,N_1540);
or U2011 (N_2011,N_1200,N_1512);
nor U2012 (N_2012,N_1244,N_1216);
nand U2013 (N_2013,N_1610,N_1241);
nor U2014 (N_2014,N_1441,N_1784);
and U2015 (N_2015,N_1745,N_1690);
and U2016 (N_2016,N_1218,N_1777);
nand U2017 (N_2017,N_1570,N_1204);
or U2018 (N_2018,N_1635,N_1310);
nand U2019 (N_2019,N_1637,N_1579);
and U2020 (N_2020,N_1384,N_1405);
and U2021 (N_2021,N_1358,N_1661);
nand U2022 (N_2022,N_1280,N_1626);
nand U2023 (N_2023,N_1254,N_1438);
nor U2024 (N_2024,N_1608,N_1444);
and U2025 (N_2025,N_1639,N_1769);
or U2026 (N_2026,N_1360,N_1674);
and U2027 (N_2027,N_1476,N_1406);
xnor U2028 (N_2028,N_1440,N_1505);
nor U2029 (N_2029,N_1583,N_1770);
nand U2030 (N_2030,N_1439,N_1524);
or U2031 (N_2031,N_1684,N_1659);
or U2032 (N_2032,N_1551,N_1369);
nor U2033 (N_2033,N_1632,N_1355);
nor U2034 (N_2034,N_1793,N_1427);
and U2035 (N_2035,N_1762,N_1543);
nand U2036 (N_2036,N_1487,N_1223);
or U2037 (N_2037,N_1560,N_1766);
nor U2038 (N_2038,N_1778,N_1246);
nand U2039 (N_2039,N_1434,N_1591);
nor U2040 (N_2040,N_1368,N_1300);
or U2041 (N_2041,N_1314,N_1798);
nand U2042 (N_2042,N_1399,N_1430);
or U2043 (N_2043,N_1364,N_1354);
nand U2044 (N_2044,N_1561,N_1327);
nor U2045 (N_2045,N_1339,N_1538);
and U2046 (N_2046,N_1671,N_1416);
and U2047 (N_2047,N_1672,N_1437);
xnor U2048 (N_2048,N_1675,N_1259);
nor U2049 (N_2049,N_1391,N_1796);
or U2050 (N_2050,N_1380,N_1562);
and U2051 (N_2051,N_1520,N_1685);
and U2052 (N_2052,N_1564,N_1250);
and U2053 (N_2053,N_1302,N_1207);
nand U2054 (N_2054,N_1385,N_1578);
or U2055 (N_2055,N_1714,N_1545);
nor U2056 (N_2056,N_1392,N_1343);
nand U2057 (N_2057,N_1780,N_1320);
and U2058 (N_2058,N_1789,N_1426);
nand U2059 (N_2059,N_1530,N_1749);
and U2060 (N_2060,N_1262,N_1256);
nand U2061 (N_2061,N_1550,N_1613);
nand U2062 (N_2062,N_1585,N_1716);
nor U2063 (N_2063,N_1219,N_1229);
and U2064 (N_2064,N_1715,N_1448);
nor U2065 (N_2065,N_1428,N_1537);
xnor U2066 (N_2066,N_1757,N_1374);
or U2067 (N_2067,N_1642,N_1599);
nand U2068 (N_2068,N_1475,N_1269);
nand U2069 (N_2069,N_1795,N_1516);
nand U2070 (N_2070,N_1288,N_1446);
and U2071 (N_2071,N_1731,N_1699);
nor U2072 (N_2072,N_1435,N_1656);
nand U2073 (N_2073,N_1708,N_1783);
nor U2074 (N_2074,N_1452,N_1315);
xnor U2075 (N_2075,N_1634,N_1222);
and U2076 (N_2076,N_1333,N_1247);
nor U2077 (N_2077,N_1501,N_1442);
and U2078 (N_2078,N_1567,N_1609);
or U2079 (N_2079,N_1450,N_1513);
or U2080 (N_2080,N_1271,N_1303);
nand U2081 (N_2081,N_1337,N_1687);
nor U2082 (N_2082,N_1569,N_1792);
nand U2083 (N_2083,N_1478,N_1539);
or U2084 (N_2084,N_1413,N_1493);
xnor U2085 (N_2085,N_1522,N_1489);
nand U2086 (N_2086,N_1411,N_1622);
nor U2087 (N_2087,N_1593,N_1202);
and U2088 (N_2088,N_1211,N_1767);
xor U2089 (N_2089,N_1443,N_1233);
or U2090 (N_2090,N_1727,N_1423);
nor U2091 (N_2091,N_1221,N_1412);
and U2092 (N_2092,N_1660,N_1394);
or U2093 (N_2093,N_1751,N_1389);
nor U2094 (N_2094,N_1773,N_1517);
nor U2095 (N_2095,N_1782,N_1753);
xnor U2096 (N_2096,N_1732,N_1361);
nor U2097 (N_2097,N_1311,N_1587);
nor U2098 (N_2098,N_1665,N_1486);
nor U2099 (N_2099,N_1313,N_1772);
nand U2100 (N_2100,N_1333,N_1574);
xor U2101 (N_2101,N_1549,N_1550);
and U2102 (N_2102,N_1702,N_1418);
nor U2103 (N_2103,N_1495,N_1379);
nand U2104 (N_2104,N_1307,N_1529);
or U2105 (N_2105,N_1646,N_1563);
and U2106 (N_2106,N_1715,N_1619);
nor U2107 (N_2107,N_1661,N_1662);
or U2108 (N_2108,N_1567,N_1683);
and U2109 (N_2109,N_1428,N_1280);
or U2110 (N_2110,N_1289,N_1369);
and U2111 (N_2111,N_1430,N_1796);
nor U2112 (N_2112,N_1413,N_1697);
nand U2113 (N_2113,N_1710,N_1789);
nor U2114 (N_2114,N_1787,N_1592);
xor U2115 (N_2115,N_1446,N_1328);
or U2116 (N_2116,N_1621,N_1379);
and U2117 (N_2117,N_1574,N_1499);
nor U2118 (N_2118,N_1380,N_1674);
or U2119 (N_2119,N_1418,N_1576);
nor U2120 (N_2120,N_1302,N_1524);
and U2121 (N_2121,N_1413,N_1452);
nor U2122 (N_2122,N_1341,N_1760);
or U2123 (N_2123,N_1784,N_1339);
and U2124 (N_2124,N_1645,N_1743);
nand U2125 (N_2125,N_1290,N_1738);
nand U2126 (N_2126,N_1779,N_1575);
or U2127 (N_2127,N_1547,N_1441);
nor U2128 (N_2128,N_1398,N_1411);
nor U2129 (N_2129,N_1677,N_1681);
nor U2130 (N_2130,N_1557,N_1791);
nand U2131 (N_2131,N_1336,N_1698);
and U2132 (N_2132,N_1528,N_1684);
or U2133 (N_2133,N_1430,N_1618);
nor U2134 (N_2134,N_1310,N_1284);
or U2135 (N_2135,N_1529,N_1546);
nor U2136 (N_2136,N_1668,N_1796);
nand U2137 (N_2137,N_1440,N_1261);
nor U2138 (N_2138,N_1619,N_1754);
nor U2139 (N_2139,N_1561,N_1530);
and U2140 (N_2140,N_1623,N_1339);
nor U2141 (N_2141,N_1567,N_1637);
or U2142 (N_2142,N_1540,N_1626);
and U2143 (N_2143,N_1418,N_1610);
or U2144 (N_2144,N_1357,N_1414);
nor U2145 (N_2145,N_1333,N_1400);
nand U2146 (N_2146,N_1449,N_1415);
nor U2147 (N_2147,N_1496,N_1786);
nand U2148 (N_2148,N_1286,N_1627);
and U2149 (N_2149,N_1558,N_1512);
and U2150 (N_2150,N_1546,N_1241);
and U2151 (N_2151,N_1365,N_1549);
nand U2152 (N_2152,N_1480,N_1625);
nor U2153 (N_2153,N_1545,N_1641);
nand U2154 (N_2154,N_1494,N_1528);
or U2155 (N_2155,N_1279,N_1777);
or U2156 (N_2156,N_1664,N_1235);
nor U2157 (N_2157,N_1358,N_1492);
nor U2158 (N_2158,N_1670,N_1709);
nor U2159 (N_2159,N_1605,N_1782);
and U2160 (N_2160,N_1372,N_1572);
or U2161 (N_2161,N_1441,N_1256);
or U2162 (N_2162,N_1217,N_1401);
nor U2163 (N_2163,N_1775,N_1432);
or U2164 (N_2164,N_1318,N_1300);
nand U2165 (N_2165,N_1673,N_1666);
or U2166 (N_2166,N_1509,N_1503);
nand U2167 (N_2167,N_1561,N_1246);
nor U2168 (N_2168,N_1491,N_1217);
or U2169 (N_2169,N_1325,N_1638);
xor U2170 (N_2170,N_1497,N_1502);
nor U2171 (N_2171,N_1682,N_1739);
nor U2172 (N_2172,N_1246,N_1479);
or U2173 (N_2173,N_1411,N_1479);
or U2174 (N_2174,N_1431,N_1271);
nor U2175 (N_2175,N_1321,N_1548);
nor U2176 (N_2176,N_1788,N_1494);
or U2177 (N_2177,N_1450,N_1546);
nor U2178 (N_2178,N_1398,N_1520);
nor U2179 (N_2179,N_1364,N_1394);
and U2180 (N_2180,N_1340,N_1570);
nor U2181 (N_2181,N_1715,N_1352);
nor U2182 (N_2182,N_1611,N_1746);
and U2183 (N_2183,N_1454,N_1256);
nand U2184 (N_2184,N_1575,N_1656);
or U2185 (N_2185,N_1368,N_1467);
and U2186 (N_2186,N_1592,N_1306);
nand U2187 (N_2187,N_1503,N_1473);
or U2188 (N_2188,N_1538,N_1799);
nor U2189 (N_2189,N_1571,N_1379);
nand U2190 (N_2190,N_1227,N_1533);
nor U2191 (N_2191,N_1388,N_1386);
or U2192 (N_2192,N_1287,N_1270);
nor U2193 (N_2193,N_1427,N_1595);
nor U2194 (N_2194,N_1270,N_1368);
or U2195 (N_2195,N_1239,N_1383);
and U2196 (N_2196,N_1794,N_1392);
nand U2197 (N_2197,N_1474,N_1682);
nand U2198 (N_2198,N_1527,N_1749);
nand U2199 (N_2199,N_1706,N_1739);
or U2200 (N_2200,N_1378,N_1563);
and U2201 (N_2201,N_1652,N_1500);
nor U2202 (N_2202,N_1515,N_1711);
nor U2203 (N_2203,N_1310,N_1769);
nor U2204 (N_2204,N_1605,N_1735);
and U2205 (N_2205,N_1639,N_1260);
nor U2206 (N_2206,N_1319,N_1231);
nand U2207 (N_2207,N_1284,N_1757);
nand U2208 (N_2208,N_1431,N_1622);
and U2209 (N_2209,N_1476,N_1459);
nor U2210 (N_2210,N_1664,N_1576);
and U2211 (N_2211,N_1487,N_1709);
or U2212 (N_2212,N_1701,N_1615);
nand U2213 (N_2213,N_1544,N_1384);
nand U2214 (N_2214,N_1755,N_1305);
or U2215 (N_2215,N_1588,N_1429);
and U2216 (N_2216,N_1701,N_1260);
nand U2217 (N_2217,N_1593,N_1429);
and U2218 (N_2218,N_1543,N_1374);
nor U2219 (N_2219,N_1571,N_1249);
or U2220 (N_2220,N_1492,N_1692);
and U2221 (N_2221,N_1455,N_1286);
nor U2222 (N_2222,N_1600,N_1353);
xnor U2223 (N_2223,N_1544,N_1707);
and U2224 (N_2224,N_1779,N_1692);
or U2225 (N_2225,N_1492,N_1738);
nand U2226 (N_2226,N_1263,N_1622);
or U2227 (N_2227,N_1205,N_1248);
nor U2228 (N_2228,N_1724,N_1246);
nand U2229 (N_2229,N_1596,N_1294);
and U2230 (N_2230,N_1554,N_1269);
nand U2231 (N_2231,N_1343,N_1446);
nor U2232 (N_2232,N_1583,N_1699);
nand U2233 (N_2233,N_1394,N_1792);
nand U2234 (N_2234,N_1439,N_1235);
xor U2235 (N_2235,N_1638,N_1589);
nor U2236 (N_2236,N_1797,N_1538);
and U2237 (N_2237,N_1459,N_1789);
and U2238 (N_2238,N_1595,N_1397);
nand U2239 (N_2239,N_1330,N_1260);
nor U2240 (N_2240,N_1596,N_1721);
and U2241 (N_2241,N_1382,N_1409);
and U2242 (N_2242,N_1470,N_1581);
nand U2243 (N_2243,N_1452,N_1766);
or U2244 (N_2244,N_1287,N_1409);
nand U2245 (N_2245,N_1579,N_1686);
and U2246 (N_2246,N_1577,N_1493);
nor U2247 (N_2247,N_1755,N_1230);
nand U2248 (N_2248,N_1721,N_1237);
nand U2249 (N_2249,N_1307,N_1745);
or U2250 (N_2250,N_1288,N_1608);
and U2251 (N_2251,N_1360,N_1578);
nand U2252 (N_2252,N_1754,N_1521);
or U2253 (N_2253,N_1333,N_1503);
and U2254 (N_2254,N_1275,N_1257);
nor U2255 (N_2255,N_1277,N_1707);
nand U2256 (N_2256,N_1635,N_1261);
xor U2257 (N_2257,N_1634,N_1684);
nand U2258 (N_2258,N_1716,N_1243);
nor U2259 (N_2259,N_1357,N_1382);
xor U2260 (N_2260,N_1389,N_1404);
nand U2261 (N_2261,N_1639,N_1559);
or U2262 (N_2262,N_1444,N_1320);
and U2263 (N_2263,N_1258,N_1763);
nand U2264 (N_2264,N_1303,N_1735);
nor U2265 (N_2265,N_1778,N_1482);
and U2266 (N_2266,N_1380,N_1508);
or U2267 (N_2267,N_1696,N_1544);
nor U2268 (N_2268,N_1315,N_1619);
or U2269 (N_2269,N_1246,N_1679);
or U2270 (N_2270,N_1607,N_1423);
and U2271 (N_2271,N_1521,N_1638);
nand U2272 (N_2272,N_1590,N_1569);
and U2273 (N_2273,N_1781,N_1457);
and U2274 (N_2274,N_1724,N_1354);
nor U2275 (N_2275,N_1295,N_1492);
and U2276 (N_2276,N_1462,N_1694);
nand U2277 (N_2277,N_1344,N_1679);
or U2278 (N_2278,N_1584,N_1375);
and U2279 (N_2279,N_1736,N_1333);
nor U2280 (N_2280,N_1474,N_1652);
or U2281 (N_2281,N_1438,N_1627);
nor U2282 (N_2282,N_1382,N_1645);
and U2283 (N_2283,N_1218,N_1390);
and U2284 (N_2284,N_1459,N_1337);
and U2285 (N_2285,N_1388,N_1538);
and U2286 (N_2286,N_1532,N_1670);
nor U2287 (N_2287,N_1264,N_1512);
and U2288 (N_2288,N_1264,N_1726);
and U2289 (N_2289,N_1296,N_1754);
nand U2290 (N_2290,N_1663,N_1291);
and U2291 (N_2291,N_1276,N_1360);
nor U2292 (N_2292,N_1608,N_1582);
nand U2293 (N_2293,N_1303,N_1399);
nand U2294 (N_2294,N_1690,N_1556);
and U2295 (N_2295,N_1521,N_1317);
and U2296 (N_2296,N_1554,N_1533);
or U2297 (N_2297,N_1761,N_1791);
and U2298 (N_2298,N_1490,N_1653);
nor U2299 (N_2299,N_1462,N_1397);
xor U2300 (N_2300,N_1779,N_1644);
or U2301 (N_2301,N_1619,N_1617);
and U2302 (N_2302,N_1273,N_1330);
or U2303 (N_2303,N_1512,N_1463);
or U2304 (N_2304,N_1516,N_1413);
and U2305 (N_2305,N_1795,N_1404);
nand U2306 (N_2306,N_1368,N_1748);
nand U2307 (N_2307,N_1392,N_1737);
nor U2308 (N_2308,N_1519,N_1565);
or U2309 (N_2309,N_1378,N_1348);
and U2310 (N_2310,N_1439,N_1752);
and U2311 (N_2311,N_1534,N_1568);
nand U2312 (N_2312,N_1612,N_1728);
and U2313 (N_2313,N_1306,N_1355);
or U2314 (N_2314,N_1770,N_1402);
xnor U2315 (N_2315,N_1413,N_1556);
or U2316 (N_2316,N_1799,N_1567);
nor U2317 (N_2317,N_1584,N_1494);
or U2318 (N_2318,N_1286,N_1446);
nor U2319 (N_2319,N_1727,N_1677);
nand U2320 (N_2320,N_1415,N_1469);
nand U2321 (N_2321,N_1523,N_1399);
or U2322 (N_2322,N_1791,N_1244);
nand U2323 (N_2323,N_1328,N_1736);
and U2324 (N_2324,N_1209,N_1285);
nor U2325 (N_2325,N_1247,N_1562);
xor U2326 (N_2326,N_1638,N_1688);
or U2327 (N_2327,N_1681,N_1635);
or U2328 (N_2328,N_1300,N_1490);
nor U2329 (N_2329,N_1205,N_1297);
or U2330 (N_2330,N_1477,N_1271);
and U2331 (N_2331,N_1777,N_1250);
nor U2332 (N_2332,N_1232,N_1796);
or U2333 (N_2333,N_1653,N_1249);
and U2334 (N_2334,N_1371,N_1541);
and U2335 (N_2335,N_1637,N_1389);
and U2336 (N_2336,N_1351,N_1465);
nand U2337 (N_2337,N_1304,N_1399);
nor U2338 (N_2338,N_1209,N_1647);
and U2339 (N_2339,N_1591,N_1342);
nand U2340 (N_2340,N_1718,N_1636);
or U2341 (N_2341,N_1688,N_1450);
nor U2342 (N_2342,N_1740,N_1216);
nand U2343 (N_2343,N_1316,N_1636);
or U2344 (N_2344,N_1565,N_1675);
and U2345 (N_2345,N_1531,N_1754);
nor U2346 (N_2346,N_1694,N_1395);
nor U2347 (N_2347,N_1323,N_1560);
xor U2348 (N_2348,N_1217,N_1439);
nand U2349 (N_2349,N_1220,N_1245);
nand U2350 (N_2350,N_1378,N_1373);
nand U2351 (N_2351,N_1378,N_1210);
nor U2352 (N_2352,N_1228,N_1289);
nor U2353 (N_2353,N_1726,N_1275);
or U2354 (N_2354,N_1646,N_1511);
or U2355 (N_2355,N_1744,N_1584);
and U2356 (N_2356,N_1486,N_1287);
nor U2357 (N_2357,N_1666,N_1671);
nor U2358 (N_2358,N_1343,N_1769);
and U2359 (N_2359,N_1263,N_1494);
nor U2360 (N_2360,N_1686,N_1780);
xor U2361 (N_2361,N_1624,N_1387);
nor U2362 (N_2362,N_1712,N_1794);
or U2363 (N_2363,N_1366,N_1598);
and U2364 (N_2364,N_1726,N_1686);
nor U2365 (N_2365,N_1609,N_1612);
nand U2366 (N_2366,N_1647,N_1255);
nor U2367 (N_2367,N_1296,N_1478);
xor U2368 (N_2368,N_1731,N_1297);
and U2369 (N_2369,N_1240,N_1466);
nand U2370 (N_2370,N_1250,N_1305);
xnor U2371 (N_2371,N_1582,N_1689);
or U2372 (N_2372,N_1513,N_1661);
nor U2373 (N_2373,N_1216,N_1695);
nor U2374 (N_2374,N_1501,N_1255);
xor U2375 (N_2375,N_1429,N_1637);
nor U2376 (N_2376,N_1540,N_1373);
or U2377 (N_2377,N_1430,N_1466);
and U2378 (N_2378,N_1346,N_1668);
or U2379 (N_2379,N_1778,N_1658);
or U2380 (N_2380,N_1413,N_1484);
and U2381 (N_2381,N_1566,N_1293);
nor U2382 (N_2382,N_1677,N_1582);
or U2383 (N_2383,N_1336,N_1728);
nand U2384 (N_2384,N_1371,N_1266);
nor U2385 (N_2385,N_1790,N_1373);
nor U2386 (N_2386,N_1593,N_1656);
nor U2387 (N_2387,N_1409,N_1274);
and U2388 (N_2388,N_1530,N_1578);
nor U2389 (N_2389,N_1264,N_1413);
or U2390 (N_2390,N_1795,N_1736);
nor U2391 (N_2391,N_1511,N_1446);
and U2392 (N_2392,N_1771,N_1414);
and U2393 (N_2393,N_1456,N_1610);
or U2394 (N_2394,N_1467,N_1369);
nor U2395 (N_2395,N_1437,N_1436);
or U2396 (N_2396,N_1426,N_1331);
nor U2397 (N_2397,N_1695,N_1685);
or U2398 (N_2398,N_1524,N_1664);
nor U2399 (N_2399,N_1210,N_1405);
and U2400 (N_2400,N_1874,N_2381);
nand U2401 (N_2401,N_1827,N_2255);
nand U2402 (N_2402,N_2075,N_2174);
nor U2403 (N_2403,N_2093,N_2288);
nand U2404 (N_2404,N_2248,N_1949);
or U2405 (N_2405,N_2217,N_1810);
or U2406 (N_2406,N_2136,N_2098);
nor U2407 (N_2407,N_2146,N_1844);
or U2408 (N_2408,N_2399,N_1987);
nand U2409 (N_2409,N_1910,N_2163);
nor U2410 (N_2410,N_2230,N_2392);
or U2411 (N_2411,N_1903,N_2150);
nand U2412 (N_2412,N_1935,N_2005);
nor U2413 (N_2413,N_2040,N_1954);
or U2414 (N_2414,N_2173,N_2127);
nor U2415 (N_2415,N_1826,N_2006);
nand U2416 (N_2416,N_2322,N_1963);
nand U2417 (N_2417,N_2316,N_1957);
and U2418 (N_2418,N_1973,N_2167);
and U2419 (N_2419,N_2170,N_1851);
and U2420 (N_2420,N_2188,N_2056);
and U2421 (N_2421,N_1882,N_1988);
and U2422 (N_2422,N_2083,N_2176);
or U2423 (N_2423,N_1905,N_2063);
or U2424 (N_2424,N_2222,N_2292);
or U2425 (N_2425,N_1815,N_1929);
and U2426 (N_2426,N_1822,N_2303);
or U2427 (N_2427,N_2268,N_1962);
xnor U2428 (N_2428,N_2192,N_2315);
nor U2429 (N_2429,N_1863,N_2311);
or U2430 (N_2430,N_1971,N_2007);
and U2431 (N_2431,N_2317,N_1921);
and U2432 (N_2432,N_1816,N_2319);
nor U2433 (N_2433,N_2291,N_1912);
nand U2434 (N_2434,N_2210,N_2215);
and U2435 (N_2435,N_1833,N_2226);
or U2436 (N_2436,N_1952,N_2211);
nand U2437 (N_2437,N_1937,N_2385);
and U2438 (N_2438,N_1809,N_2280);
and U2439 (N_2439,N_2221,N_2344);
and U2440 (N_2440,N_2143,N_2364);
nor U2441 (N_2441,N_2369,N_1968);
nand U2442 (N_2442,N_2356,N_2131);
or U2443 (N_2443,N_1848,N_2086);
nor U2444 (N_2444,N_2139,N_2122);
or U2445 (N_2445,N_2106,N_2335);
nand U2446 (N_2446,N_2240,N_2123);
nand U2447 (N_2447,N_2147,N_2087);
and U2448 (N_2448,N_2144,N_1950);
nand U2449 (N_2449,N_2142,N_1852);
nor U2450 (N_2450,N_1996,N_1944);
or U2451 (N_2451,N_2012,N_2051);
nor U2452 (N_2452,N_1993,N_2084);
nor U2453 (N_2453,N_2391,N_1958);
and U2454 (N_2454,N_1881,N_2134);
nor U2455 (N_2455,N_1840,N_2237);
nor U2456 (N_2456,N_2297,N_2029);
or U2457 (N_2457,N_2293,N_1974);
or U2458 (N_2458,N_1884,N_2074);
or U2459 (N_2459,N_2125,N_2080);
or U2460 (N_2460,N_2341,N_2002);
or U2461 (N_2461,N_2299,N_1823);
nor U2462 (N_2462,N_2078,N_2193);
and U2463 (N_2463,N_1857,N_1893);
nor U2464 (N_2464,N_2042,N_2371);
nand U2465 (N_2465,N_2151,N_2333);
xor U2466 (N_2466,N_1934,N_1946);
nand U2467 (N_2467,N_2037,N_2104);
and U2468 (N_2468,N_1837,N_2031);
nand U2469 (N_2469,N_2201,N_1967);
or U2470 (N_2470,N_2312,N_1897);
or U2471 (N_2471,N_1859,N_2039);
nor U2472 (N_2472,N_2017,N_2236);
and U2473 (N_2473,N_1972,N_1861);
and U2474 (N_2474,N_1834,N_1832);
or U2475 (N_2475,N_2105,N_2102);
or U2476 (N_2476,N_2015,N_1831);
nand U2477 (N_2477,N_2388,N_1866);
nor U2478 (N_2478,N_2383,N_2013);
nor U2479 (N_2479,N_2300,N_2234);
nand U2480 (N_2480,N_2379,N_2153);
nand U2481 (N_2481,N_2032,N_1803);
nor U2482 (N_2482,N_2332,N_2099);
nor U2483 (N_2483,N_2091,N_2286);
nand U2484 (N_2484,N_1875,N_1924);
nor U2485 (N_2485,N_2185,N_2137);
and U2486 (N_2486,N_2362,N_2119);
nor U2487 (N_2487,N_2004,N_2145);
and U2488 (N_2488,N_1915,N_2314);
and U2489 (N_2489,N_1941,N_2320);
or U2490 (N_2490,N_2008,N_2073);
or U2491 (N_2491,N_1800,N_1867);
or U2492 (N_2492,N_1979,N_1943);
nand U2493 (N_2493,N_2169,N_2393);
and U2494 (N_2494,N_2339,N_2380);
nand U2495 (N_2495,N_2160,N_1932);
or U2496 (N_2496,N_2057,N_1983);
and U2497 (N_2497,N_1936,N_2090);
nand U2498 (N_2498,N_2289,N_1825);
nor U2499 (N_2499,N_2273,N_1821);
nor U2500 (N_2500,N_1830,N_1985);
or U2501 (N_2501,N_2269,N_1911);
or U2502 (N_2502,N_1870,N_1933);
nor U2503 (N_2503,N_2378,N_2081);
and U2504 (N_2504,N_2166,N_2306);
nor U2505 (N_2505,N_2296,N_2329);
nor U2506 (N_2506,N_2347,N_2359);
nor U2507 (N_2507,N_2020,N_2115);
or U2508 (N_2508,N_2065,N_1913);
or U2509 (N_2509,N_1843,N_1853);
nand U2510 (N_2510,N_2249,N_2103);
and U2511 (N_2511,N_2338,N_2281);
nand U2512 (N_2512,N_1918,N_1969);
or U2513 (N_2513,N_2313,N_1824);
and U2514 (N_2514,N_1938,N_1953);
or U2515 (N_2515,N_2187,N_2373);
nor U2516 (N_2516,N_2244,N_2178);
nand U2517 (N_2517,N_2271,N_1845);
nand U2518 (N_2518,N_2172,N_1819);
nor U2519 (N_2519,N_2116,N_2054);
or U2520 (N_2520,N_2113,N_1898);
nor U2521 (N_2521,N_2366,N_2257);
or U2522 (N_2522,N_2328,N_2181);
xnor U2523 (N_2523,N_2390,N_1980);
or U2524 (N_2524,N_1876,N_1838);
nand U2525 (N_2525,N_2377,N_1871);
and U2526 (N_2526,N_2001,N_2034);
nor U2527 (N_2527,N_2070,N_2171);
nor U2528 (N_2528,N_2047,N_2206);
and U2529 (N_2529,N_2168,N_2274);
and U2530 (N_2530,N_1854,N_2016);
nor U2531 (N_2531,N_2374,N_1899);
or U2532 (N_2532,N_1978,N_1966);
nand U2533 (N_2533,N_1923,N_2183);
or U2534 (N_2534,N_2395,N_2128);
nand U2535 (N_2535,N_2294,N_2219);
and U2536 (N_2536,N_1970,N_2228);
nor U2537 (N_2537,N_2350,N_1812);
nor U2538 (N_2538,N_1801,N_2245);
nand U2539 (N_2539,N_1849,N_2129);
nor U2540 (N_2540,N_2052,N_1892);
and U2541 (N_2541,N_1886,N_2101);
and U2542 (N_2542,N_2355,N_2033);
and U2543 (N_2543,N_2071,N_2241);
nor U2544 (N_2544,N_1961,N_1909);
nand U2545 (N_2545,N_1916,N_2055);
nand U2546 (N_2546,N_2049,N_2207);
nand U2547 (N_2547,N_2233,N_2044);
nor U2548 (N_2548,N_2024,N_1907);
nor U2549 (N_2549,N_1880,N_2212);
nor U2550 (N_2550,N_1989,N_2096);
or U2551 (N_2551,N_2256,N_1990);
nand U2552 (N_2552,N_2307,N_2041);
and U2553 (N_2553,N_2301,N_2154);
or U2554 (N_2554,N_2331,N_1991);
and U2555 (N_2555,N_2179,N_2066);
and U2556 (N_2556,N_1900,N_1856);
xor U2557 (N_2557,N_2360,N_1804);
or U2558 (N_2558,N_2100,N_2357);
and U2559 (N_2559,N_1942,N_2097);
and U2560 (N_2560,N_1839,N_1885);
or U2561 (N_2561,N_2229,N_2191);
and U2562 (N_2562,N_2214,N_2326);
nand U2563 (N_2563,N_1960,N_2111);
nor U2564 (N_2564,N_2260,N_2345);
or U2565 (N_2565,N_2323,N_1928);
and U2566 (N_2566,N_2209,N_1872);
nor U2567 (N_2567,N_2023,N_2223);
nor U2568 (N_2568,N_2365,N_2177);
nand U2569 (N_2569,N_2351,N_2067);
and U2570 (N_2570,N_1914,N_1939);
or U2571 (N_2571,N_2022,N_1965);
and U2572 (N_2572,N_2082,N_2343);
nand U2573 (N_2573,N_1975,N_2336);
or U2574 (N_2574,N_2019,N_1891);
nand U2575 (N_2575,N_2069,N_1890);
nor U2576 (N_2576,N_2130,N_2048);
nor U2577 (N_2577,N_2107,N_2352);
nand U2578 (N_2578,N_2277,N_2003);
or U2579 (N_2579,N_1865,N_2318);
or U2580 (N_2580,N_1922,N_2059);
or U2581 (N_2581,N_2224,N_1889);
and U2582 (N_2582,N_1864,N_2198);
nand U2583 (N_2583,N_2018,N_2035);
or U2584 (N_2584,N_2158,N_2050);
or U2585 (N_2585,N_1945,N_1806);
nor U2586 (N_2586,N_2284,N_1877);
or U2587 (N_2587,N_2009,N_2349);
nor U2588 (N_2588,N_2021,N_2372);
and U2589 (N_2589,N_2194,N_1917);
nor U2590 (N_2590,N_2064,N_2076);
nor U2591 (N_2591,N_1926,N_2200);
nor U2592 (N_2592,N_2060,N_2156);
nor U2593 (N_2593,N_2302,N_2354);
nand U2594 (N_2594,N_2164,N_2072);
nor U2595 (N_2595,N_2165,N_2186);
nor U2596 (N_2596,N_1895,N_2367);
and U2597 (N_2597,N_1858,N_2304);
nand U2598 (N_2598,N_2327,N_1998);
nand U2599 (N_2599,N_2259,N_1887);
or U2600 (N_2600,N_2218,N_1850);
nor U2601 (N_2601,N_1896,N_2028);
nor U2602 (N_2602,N_2085,N_2014);
nand U2603 (N_2603,N_2384,N_1836);
or U2604 (N_2604,N_2197,N_2253);
nor U2605 (N_2605,N_2267,N_1818);
nand U2606 (N_2606,N_2348,N_1894);
or U2607 (N_2607,N_2225,N_2308);
and U2608 (N_2608,N_1805,N_1919);
and U2609 (N_2609,N_2295,N_2199);
or U2610 (N_2610,N_2000,N_2298);
or U2611 (N_2611,N_2045,N_1802);
or U2612 (N_2612,N_1927,N_2276);
nor U2613 (N_2613,N_2272,N_2305);
nand U2614 (N_2614,N_2309,N_2278);
nor U2615 (N_2615,N_2375,N_2262);
nand U2616 (N_2616,N_2068,N_1940);
and U2617 (N_2617,N_2148,N_2114);
or U2618 (N_2618,N_2025,N_2398);
and U2619 (N_2619,N_1842,N_2196);
or U2620 (N_2620,N_2011,N_2370);
and U2621 (N_2621,N_2283,N_2232);
nor U2622 (N_2622,N_2095,N_2337);
xor U2623 (N_2623,N_2118,N_1869);
and U2624 (N_2624,N_2263,N_2152);
and U2625 (N_2625,N_1948,N_1902);
nor U2626 (N_2626,N_2133,N_1873);
or U2627 (N_2627,N_2112,N_1808);
nand U2628 (N_2628,N_2252,N_1994);
nand U2629 (N_2629,N_2157,N_2342);
nand U2630 (N_2630,N_2132,N_2243);
or U2631 (N_2631,N_2046,N_2246);
and U2632 (N_2632,N_1951,N_2062);
nor U2633 (N_2633,N_2346,N_2202);
or U2634 (N_2634,N_2030,N_1984);
and U2635 (N_2635,N_2138,N_2058);
nor U2636 (N_2636,N_2155,N_1999);
nor U2637 (N_2637,N_1977,N_2275);
nor U2638 (N_2638,N_2204,N_2149);
nand U2639 (N_2639,N_1813,N_2368);
nor U2640 (N_2640,N_2387,N_2108);
and U2641 (N_2641,N_2135,N_2140);
nor U2642 (N_2642,N_1829,N_2266);
nor U2643 (N_2643,N_2089,N_1982);
or U2644 (N_2644,N_2353,N_1868);
and U2645 (N_2645,N_1981,N_2238);
or U2646 (N_2646,N_2340,N_2189);
nand U2647 (N_2647,N_2358,N_2325);
nor U2648 (N_2648,N_2094,N_1879);
nor U2649 (N_2649,N_2036,N_2264);
nor U2650 (N_2650,N_2126,N_2361);
nand U2651 (N_2651,N_2389,N_2027);
or U2652 (N_2652,N_2386,N_2180);
or U2653 (N_2653,N_2110,N_1920);
nand U2654 (N_2654,N_2261,N_2053);
nand U2655 (N_2655,N_1811,N_2258);
or U2656 (N_2656,N_1817,N_2285);
nor U2657 (N_2657,N_2287,N_2043);
or U2658 (N_2658,N_1906,N_2279);
and U2659 (N_2659,N_2208,N_1841);
nand U2660 (N_2660,N_2250,N_2231);
nor U2661 (N_2661,N_1986,N_1992);
nand U2662 (N_2662,N_2109,N_1860);
and U2663 (N_2663,N_2120,N_2010);
nand U2664 (N_2664,N_2216,N_2270);
nor U2665 (N_2665,N_2038,N_2227);
or U2666 (N_2666,N_2321,N_2121);
and U2667 (N_2667,N_1855,N_2061);
nor U2668 (N_2668,N_2184,N_2363);
nor U2669 (N_2669,N_2251,N_1997);
nor U2670 (N_2670,N_1995,N_2247);
and U2671 (N_2671,N_2117,N_2382);
nor U2672 (N_2672,N_1862,N_1820);
and U2673 (N_2673,N_2182,N_2310);
xnor U2674 (N_2674,N_2396,N_1828);
and U2675 (N_2675,N_1930,N_2190);
and U2676 (N_2676,N_2282,N_2159);
nand U2677 (N_2677,N_2394,N_2397);
and U2678 (N_2678,N_1814,N_1955);
nor U2679 (N_2679,N_1807,N_2077);
or U2680 (N_2680,N_2203,N_1878);
nor U2681 (N_2681,N_1888,N_2330);
nor U2682 (N_2682,N_1959,N_1846);
xnor U2683 (N_2683,N_2254,N_2092);
or U2684 (N_2684,N_1901,N_2162);
or U2685 (N_2685,N_2205,N_2242);
and U2686 (N_2686,N_2324,N_1847);
or U2687 (N_2687,N_1956,N_2026);
or U2688 (N_2688,N_1964,N_2195);
and U2689 (N_2689,N_2141,N_1931);
nor U2690 (N_2690,N_2220,N_1883);
nor U2691 (N_2691,N_2213,N_2376);
or U2692 (N_2692,N_2161,N_2334);
nor U2693 (N_2693,N_2175,N_1925);
nand U2694 (N_2694,N_2290,N_1947);
nor U2695 (N_2695,N_2239,N_2235);
and U2696 (N_2696,N_1976,N_2124);
and U2697 (N_2697,N_1835,N_2079);
nand U2698 (N_2698,N_2265,N_2088);
nand U2699 (N_2699,N_1908,N_1904);
and U2700 (N_2700,N_2186,N_2246);
nor U2701 (N_2701,N_1801,N_2306);
and U2702 (N_2702,N_2164,N_2285);
and U2703 (N_2703,N_2032,N_2354);
nor U2704 (N_2704,N_1859,N_2375);
and U2705 (N_2705,N_2241,N_1956);
or U2706 (N_2706,N_1859,N_2094);
or U2707 (N_2707,N_1983,N_1939);
nand U2708 (N_2708,N_2375,N_2084);
and U2709 (N_2709,N_2357,N_2169);
nor U2710 (N_2710,N_2065,N_2165);
or U2711 (N_2711,N_2393,N_2204);
or U2712 (N_2712,N_2080,N_1917);
nor U2713 (N_2713,N_2370,N_1975);
and U2714 (N_2714,N_1816,N_2304);
nand U2715 (N_2715,N_2106,N_2243);
nand U2716 (N_2716,N_2232,N_2214);
or U2717 (N_2717,N_2391,N_2154);
or U2718 (N_2718,N_2222,N_2221);
and U2719 (N_2719,N_2049,N_2161);
or U2720 (N_2720,N_2063,N_2023);
or U2721 (N_2721,N_2211,N_2162);
and U2722 (N_2722,N_1963,N_2116);
and U2723 (N_2723,N_1810,N_1886);
nor U2724 (N_2724,N_1885,N_2105);
nand U2725 (N_2725,N_2027,N_1808);
nand U2726 (N_2726,N_1978,N_1892);
or U2727 (N_2727,N_2125,N_2273);
nand U2728 (N_2728,N_2221,N_2179);
nand U2729 (N_2729,N_2004,N_2390);
and U2730 (N_2730,N_2166,N_2334);
or U2731 (N_2731,N_2018,N_1937);
nand U2732 (N_2732,N_1986,N_1810);
and U2733 (N_2733,N_1806,N_1813);
or U2734 (N_2734,N_2241,N_1892);
and U2735 (N_2735,N_2133,N_1800);
nor U2736 (N_2736,N_1844,N_2095);
or U2737 (N_2737,N_1943,N_2019);
nand U2738 (N_2738,N_1820,N_2205);
and U2739 (N_2739,N_2385,N_1824);
nor U2740 (N_2740,N_1938,N_2268);
and U2741 (N_2741,N_2212,N_1971);
nand U2742 (N_2742,N_2231,N_2232);
and U2743 (N_2743,N_2290,N_1967);
nor U2744 (N_2744,N_1815,N_1857);
or U2745 (N_2745,N_2143,N_2112);
nor U2746 (N_2746,N_2226,N_2272);
nand U2747 (N_2747,N_2045,N_2282);
nand U2748 (N_2748,N_2303,N_2211);
and U2749 (N_2749,N_1991,N_1883);
and U2750 (N_2750,N_2238,N_2151);
and U2751 (N_2751,N_2223,N_2099);
nand U2752 (N_2752,N_2280,N_1873);
nor U2753 (N_2753,N_1844,N_1943);
or U2754 (N_2754,N_2197,N_2123);
nor U2755 (N_2755,N_1922,N_2046);
and U2756 (N_2756,N_2228,N_2182);
nand U2757 (N_2757,N_2150,N_2120);
xor U2758 (N_2758,N_1841,N_1936);
and U2759 (N_2759,N_2376,N_2158);
and U2760 (N_2760,N_2234,N_1856);
nand U2761 (N_2761,N_2018,N_1978);
or U2762 (N_2762,N_2159,N_2237);
and U2763 (N_2763,N_2111,N_2021);
nand U2764 (N_2764,N_1929,N_2352);
and U2765 (N_2765,N_2039,N_1877);
or U2766 (N_2766,N_1995,N_2088);
and U2767 (N_2767,N_1929,N_2270);
or U2768 (N_2768,N_1961,N_2103);
nand U2769 (N_2769,N_2140,N_2250);
nand U2770 (N_2770,N_1993,N_1916);
and U2771 (N_2771,N_1984,N_2315);
or U2772 (N_2772,N_2332,N_1806);
nand U2773 (N_2773,N_1950,N_2262);
nor U2774 (N_2774,N_1815,N_2237);
or U2775 (N_2775,N_2382,N_2006);
or U2776 (N_2776,N_2365,N_1909);
or U2777 (N_2777,N_1885,N_1921);
nand U2778 (N_2778,N_1876,N_2131);
nor U2779 (N_2779,N_2084,N_2044);
nand U2780 (N_2780,N_1849,N_1949);
nor U2781 (N_2781,N_1882,N_2288);
or U2782 (N_2782,N_2270,N_2318);
or U2783 (N_2783,N_1834,N_2064);
and U2784 (N_2784,N_2317,N_1869);
nand U2785 (N_2785,N_2118,N_2051);
nand U2786 (N_2786,N_2048,N_2102);
or U2787 (N_2787,N_1828,N_2065);
nor U2788 (N_2788,N_2161,N_1802);
nor U2789 (N_2789,N_2292,N_2052);
or U2790 (N_2790,N_2391,N_2224);
or U2791 (N_2791,N_1900,N_2049);
nor U2792 (N_2792,N_1949,N_2045);
nor U2793 (N_2793,N_2294,N_2372);
and U2794 (N_2794,N_2279,N_2144);
nand U2795 (N_2795,N_1873,N_1975);
nor U2796 (N_2796,N_2248,N_2178);
nor U2797 (N_2797,N_2100,N_1861);
or U2798 (N_2798,N_1956,N_2345);
or U2799 (N_2799,N_1890,N_1822);
and U2800 (N_2800,N_1991,N_2138);
nor U2801 (N_2801,N_2042,N_2051);
or U2802 (N_2802,N_1909,N_1808);
nor U2803 (N_2803,N_1943,N_2175);
or U2804 (N_2804,N_2154,N_2291);
or U2805 (N_2805,N_1915,N_2127);
nand U2806 (N_2806,N_2214,N_2310);
nand U2807 (N_2807,N_2145,N_2076);
and U2808 (N_2808,N_2169,N_1909);
nand U2809 (N_2809,N_1963,N_1909);
and U2810 (N_2810,N_2280,N_2096);
nor U2811 (N_2811,N_2272,N_2066);
nand U2812 (N_2812,N_2289,N_1952);
nor U2813 (N_2813,N_2014,N_2218);
nand U2814 (N_2814,N_1915,N_2174);
nor U2815 (N_2815,N_2250,N_2091);
and U2816 (N_2816,N_1967,N_2327);
or U2817 (N_2817,N_2187,N_2005);
nand U2818 (N_2818,N_2129,N_1939);
and U2819 (N_2819,N_2020,N_2053);
and U2820 (N_2820,N_1816,N_1838);
nand U2821 (N_2821,N_2153,N_1819);
nor U2822 (N_2822,N_2308,N_2334);
or U2823 (N_2823,N_1803,N_1869);
nand U2824 (N_2824,N_1995,N_2215);
xor U2825 (N_2825,N_1833,N_2306);
nand U2826 (N_2826,N_1942,N_2006);
or U2827 (N_2827,N_2007,N_2278);
nand U2828 (N_2828,N_1982,N_1885);
nand U2829 (N_2829,N_2155,N_1858);
and U2830 (N_2830,N_1814,N_2287);
or U2831 (N_2831,N_2083,N_2188);
or U2832 (N_2832,N_2236,N_2155);
or U2833 (N_2833,N_1814,N_2143);
or U2834 (N_2834,N_2130,N_2197);
and U2835 (N_2835,N_2013,N_1994);
nor U2836 (N_2836,N_1913,N_2207);
nand U2837 (N_2837,N_2015,N_1843);
nor U2838 (N_2838,N_2277,N_2091);
and U2839 (N_2839,N_1956,N_2351);
nand U2840 (N_2840,N_1928,N_2331);
or U2841 (N_2841,N_2177,N_1933);
nor U2842 (N_2842,N_2193,N_2092);
or U2843 (N_2843,N_1999,N_2363);
or U2844 (N_2844,N_2319,N_2002);
and U2845 (N_2845,N_1935,N_2331);
nor U2846 (N_2846,N_2289,N_1914);
nor U2847 (N_2847,N_1848,N_2162);
nor U2848 (N_2848,N_1923,N_2101);
nor U2849 (N_2849,N_2130,N_1863);
nand U2850 (N_2850,N_2113,N_2160);
nor U2851 (N_2851,N_2065,N_1914);
or U2852 (N_2852,N_1976,N_1852);
nor U2853 (N_2853,N_1863,N_2160);
or U2854 (N_2854,N_2177,N_2332);
or U2855 (N_2855,N_2331,N_1913);
and U2856 (N_2856,N_2244,N_2186);
nand U2857 (N_2857,N_2012,N_1989);
or U2858 (N_2858,N_1935,N_2378);
nand U2859 (N_2859,N_2176,N_2374);
nand U2860 (N_2860,N_1830,N_2150);
xnor U2861 (N_2861,N_1865,N_2189);
and U2862 (N_2862,N_1967,N_1974);
or U2863 (N_2863,N_1886,N_2163);
nand U2864 (N_2864,N_2173,N_2385);
and U2865 (N_2865,N_2294,N_2172);
nand U2866 (N_2866,N_2210,N_2199);
or U2867 (N_2867,N_2006,N_1954);
or U2868 (N_2868,N_1909,N_2296);
nor U2869 (N_2869,N_2226,N_2077);
nor U2870 (N_2870,N_2260,N_1879);
and U2871 (N_2871,N_2243,N_2114);
or U2872 (N_2872,N_2020,N_2040);
and U2873 (N_2873,N_2339,N_2255);
or U2874 (N_2874,N_2231,N_1929);
or U2875 (N_2875,N_1863,N_2065);
nor U2876 (N_2876,N_2155,N_2148);
nand U2877 (N_2877,N_2045,N_1966);
and U2878 (N_2878,N_1843,N_2149);
nand U2879 (N_2879,N_2197,N_2020);
or U2880 (N_2880,N_1851,N_2088);
and U2881 (N_2881,N_1948,N_2373);
nand U2882 (N_2882,N_2078,N_2083);
or U2883 (N_2883,N_1833,N_2346);
and U2884 (N_2884,N_1981,N_2215);
nand U2885 (N_2885,N_1859,N_2002);
and U2886 (N_2886,N_2026,N_2192);
nand U2887 (N_2887,N_2311,N_2075);
nor U2888 (N_2888,N_1855,N_2127);
nor U2889 (N_2889,N_2013,N_2328);
or U2890 (N_2890,N_1998,N_2138);
or U2891 (N_2891,N_2024,N_2019);
or U2892 (N_2892,N_2351,N_2083);
and U2893 (N_2893,N_2073,N_1838);
nand U2894 (N_2894,N_2161,N_2138);
nand U2895 (N_2895,N_1829,N_1929);
nor U2896 (N_2896,N_2170,N_1977);
or U2897 (N_2897,N_2200,N_1841);
and U2898 (N_2898,N_1857,N_1945);
nor U2899 (N_2899,N_2084,N_2235);
nand U2900 (N_2900,N_2360,N_2224);
or U2901 (N_2901,N_1808,N_1809);
or U2902 (N_2902,N_2348,N_1968);
and U2903 (N_2903,N_2167,N_2162);
nor U2904 (N_2904,N_1808,N_1839);
nand U2905 (N_2905,N_1901,N_2279);
nor U2906 (N_2906,N_2071,N_2228);
xor U2907 (N_2907,N_1944,N_2366);
nand U2908 (N_2908,N_2278,N_1951);
or U2909 (N_2909,N_2365,N_2327);
nor U2910 (N_2910,N_2102,N_2017);
nor U2911 (N_2911,N_2207,N_2074);
nand U2912 (N_2912,N_2320,N_1979);
nor U2913 (N_2913,N_2180,N_2103);
nor U2914 (N_2914,N_1801,N_2117);
nand U2915 (N_2915,N_1913,N_2057);
and U2916 (N_2916,N_2021,N_1806);
nand U2917 (N_2917,N_1873,N_2075);
nor U2918 (N_2918,N_2258,N_1829);
or U2919 (N_2919,N_2099,N_2179);
nor U2920 (N_2920,N_1815,N_1841);
nand U2921 (N_2921,N_2379,N_1987);
and U2922 (N_2922,N_2057,N_2123);
nand U2923 (N_2923,N_1822,N_2171);
and U2924 (N_2924,N_1891,N_2248);
and U2925 (N_2925,N_2276,N_1811);
or U2926 (N_2926,N_1937,N_2297);
nor U2927 (N_2927,N_1866,N_2379);
and U2928 (N_2928,N_2158,N_1905);
nand U2929 (N_2929,N_2000,N_2195);
and U2930 (N_2930,N_2167,N_2081);
and U2931 (N_2931,N_2299,N_2314);
nor U2932 (N_2932,N_1846,N_1984);
nand U2933 (N_2933,N_2155,N_2084);
nand U2934 (N_2934,N_2130,N_2034);
or U2935 (N_2935,N_2146,N_1970);
nand U2936 (N_2936,N_1921,N_2292);
or U2937 (N_2937,N_1804,N_2362);
nor U2938 (N_2938,N_2248,N_2029);
or U2939 (N_2939,N_2009,N_2207);
or U2940 (N_2940,N_1808,N_2354);
and U2941 (N_2941,N_2283,N_2307);
or U2942 (N_2942,N_1900,N_2267);
nand U2943 (N_2943,N_2280,N_1863);
nand U2944 (N_2944,N_2206,N_2356);
or U2945 (N_2945,N_1888,N_1875);
nand U2946 (N_2946,N_2371,N_2007);
and U2947 (N_2947,N_1953,N_2342);
or U2948 (N_2948,N_1983,N_1936);
and U2949 (N_2949,N_2113,N_1806);
or U2950 (N_2950,N_1845,N_1817);
nor U2951 (N_2951,N_1994,N_2086);
or U2952 (N_2952,N_2365,N_2333);
or U2953 (N_2953,N_1988,N_2038);
nor U2954 (N_2954,N_1915,N_1877);
and U2955 (N_2955,N_2329,N_2142);
and U2956 (N_2956,N_1841,N_1809);
nand U2957 (N_2957,N_2351,N_1903);
nor U2958 (N_2958,N_2239,N_1833);
xnor U2959 (N_2959,N_2380,N_2399);
or U2960 (N_2960,N_2225,N_1962);
nand U2961 (N_2961,N_1978,N_2044);
nand U2962 (N_2962,N_1989,N_2356);
or U2963 (N_2963,N_1908,N_1990);
nand U2964 (N_2964,N_1810,N_2054);
nand U2965 (N_2965,N_2386,N_2126);
nor U2966 (N_2966,N_2399,N_1890);
or U2967 (N_2967,N_1850,N_2391);
nor U2968 (N_2968,N_2304,N_1872);
and U2969 (N_2969,N_2380,N_1943);
and U2970 (N_2970,N_1990,N_1904);
or U2971 (N_2971,N_2189,N_2134);
nor U2972 (N_2972,N_2223,N_1983);
or U2973 (N_2973,N_2249,N_2105);
nor U2974 (N_2974,N_2076,N_2071);
nor U2975 (N_2975,N_2160,N_2322);
or U2976 (N_2976,N_1938,N_2277);
nand U2977 (N_2977,N_2176,N_1854);
nor U2978 (N_2978,N_2043,N_2201);
or U2979 (N_2979,N_2323,N_2230);
xor U2980 (N_2980,N_2110,N_1983);
and U2981 (N_2981,N_2075,N_2176);
and U2982 (N_2982,N_2120,N_1813);
xor U2983 (N_2983,N_1954,N_2251);
and U2984 (N_2984,N_2335,N_2338);
nor U2985 (N_2985,N_2301,N_2121);
nand U2986 (N_2986,N_1826,N_1874);
and U2987 (N_2987,N_2108,N_1982);
nor U2988 (N_2988,N_2183,N_2331);
nand U2989 (N_2989,N_2041,N_1890);
nand U2990 (N_2990,N_2311,N_2219);
nor U2991 (N_2991,N_2211,N_2066);
or U2992 (N_2992,N_2289,N_1974);
nand U2993 (N_2993,N_1887,N_2167);
nor U2994 (N_2994,N_1976,N_2099);
or U2995 (N_2995,N_1902,N_2039);
and U2996 (N_2996,N_1917,N_2393);
nand U2997 (N_2997,N_2010,N_2278);
and U2998 (N_2998,N_2265,N_2068);
nor U2999 (N_2999,N_1875,N_2191);
nand UO_0 (O_0,N_2911,N_2539);
xnor UO_1 (O_1,N_2966,N_2444);
xor UO_2 (O_2,N_2897,N_2989);
nor UO_3 (O_3,N_2418,N_2504);
or UO_4 (O_4,N_2459,N_2685);
or UO_5 (O_5,N_2657,N_2781);
nor UO_6 (O_6,N_2864,N_2667);
and UO_7 (O_7,N_2853,N_2973);
and UO_8 (O_8,N_2754,N_2970);
or UO_9 (O_9,N_2651,N_2465);
or UO_10 (O_10,N_2585,N_2799);
nand UO_11 (O_11,N_2600,N_2936);
nand UO_12 (O_12,N_2728,N_2818);
or UO_13 (O_13,N_2987,N_2684);
nor UO_14 (O_14,N_2785,N_2437);
nand UO_15 (O_15,N_2851,N_2934);
or UO_16 (O_16,N_2944,N_2976);
and UO_17 (O_17,N_2741,N_2500);
nor UO_18 (O_18,N_2790,N_2972);
nand UO_19 (O_19,N_2784,N_2968);
nor UO_20 (O_20,N_2903,N_2647);
or UO_21 (O_21,N_2886,N_2681);
and UO_22 (O_22,N_2695,N_2601);
nor UO_23 (O_23,N_2527,N_2889);
and UO_24 (O_24,N_2672,N_2922);
nand UO_25 (O_25,N_2674,N_2965);
nand UO_26 (O_26,N_2845,N_2740);
nor UO_27 (O_27,N_2501,N_2505);
and UO_28 (O_28,N_2863,N_2919);
xor UO_29 (O_29,N_2441,N_2718);
xor UO_30 (O_30,N_2478,N_2920);
nor UO_31 (O_31,N_2562,N_2708);
nand UO_32 (O_32,N_2964,N_2872);
nor UO_33 (O_33,N_2727,N_2443);
nor UO_34 (O_34,N_2883,N_2469);
or UO_35 (O_35,N_2737,N_2570);
nor UO_36 (O_36,N_2795,N_2991);
nor UO_37 (O_37,N_2400,N_2438);
nand UO_38 (O_38,N_2706,N_2524);
and UO_39 (O_39,N_2683,N_2884);
nor UO_40 (O_40,N_2617,N_2619);
or UO_41 (O_41,N_2419,N_2658);
nor UO_42 (O_42,N_2963,N_2560);
or UO_43 (O_43,N_2497,N_2519);
and UO_44 (O_44,N_2645,N_2630);
and UO_45 (O_45,N_2756,N_2850);
and UO_46 (O_46,N_2981,N_2486);
and UO_47 (O_47,N_2468,N_2719);
and UO_48 (O_48,N_2530,N_2881);
and UO_49 (O_49,N_2548,N_2557);
or UO_50 (O_50,N_2646,N_2440);
and UO_51 (O_51,N_2652,N_2520);
nor UO_52 (O_52,N_2638,N_2753);
nand UO_53 (O_53,N_2580,N_2875);
or UO_54 (O_54,N_2885,N_2536);
or UO_55 (O_55,N_2542,N_2910);
nand UO_56 (O_56,N_2528,N_2545);
or UO_57 (O_57,N_2602,N_2406);
nand UO_58 (O_58,N_2430,N_2711);
or UO_59 (O_59,N_2434,N_2534);
nand UO_60 (O_60,N_2742,N_2415);
and UO_61 (O_61,N_2916,N_2703);
nor UO_62 (O_62,N_2767,N_2757);
nor UO_63 (O_63,N_2531,N_2957);
xnor UO_64 (O_64,N_2788,N_2538);
nand UO_65 (O_65,N_2893,N_2868);
or UO_66 (O_66,N_2618,N_2961);
nor UO_67 (O_67,N_2848,N_2955);
and UO_68 (O_68,N_2447,N_2631);
or UO_69 (O_69,N_2834,N_2787);
nor UO_70 (O_70,N_2947,N_2458);
and UO_71 (O_71,N_2852,N_2840);
nor UO_72 (O_72,N_2694,N_2643);
and UO_73 (O_73,N_2938,N_2496);
or UO_74 (O_74,N_2523,N_2661);
nor UO_75 (O_75,N_2690,N_2994);
nor UO_76 (O_76,N_2898,N_2584);
nand UO_77 (O_77,N_2763,N_2629);
nand UO_78 (O_78,N_2417,N_2574);
nand UO_79 (O_79,N_2993,N_2857);
nor UO_80 (O_80,N_2825,N_2907);
nor UO_81 (O_81,N_2675,N_2791);
and UO_82 (O_82,N_2554,N_2710);
nand UO_83 (O_83,N_2641,N_2571);
and UO_84 (O_84,N_2828,N_2621);
nor UO_85 (O_85,N_2773,N_2827);
nor UO_86 (O_86,N_2770,N_2482);
and UO_87 (O_87,N_2516,N_2862);
and UO_88 (O_88,N_2591,N_2759);
nor UO_89 (O_89,N_2954,N_2768);
nand UO_90 (O_90,N_2452,N_2697);
or UO_91 (O_91,N_2755,N_2449);
or UO_92 (O_92,N_2564,N_2462);
or UO_93 (O_93,N_2945,N_2448);
nor UO_94 (O_94,N_2926,N_2810);
nor UO_95 (O_95,N_2783,N_2854);
and UO_96 (O_96,N_2593,N_2698);
nor UO_97 (O_97,N_2456,N_2809);
xor UO_98 (O_98,N_2635,N_2822);
nand UO_99 (O_99,N_2811,N_2775);
nor UO_100 (O_100,N_2717,N_2603);
nand UO_101 (O_101,N_2990,N_2807);
and UO_102 (O_102,N_2779,N_2569);
nand UO_103 (O_103,N_2833,N_2835);
nor UO_104 (O_104,N_2761,N_2928);
nor UO_105 (O_105,N_2623,N_2701);
and UO_106 (O_106,N_2942,N_2529);
and UO_107 (O_107,N_2606,N_2561);
nor UO_108 (O_108,N_2669,N_2817);
or UO_109 (O_109,N_2613,N_2436);
and UO_110 (O_110,N_2992,N_2874);
or UO_111 (O_111,N_2549,N_2867);
nor UO_112 (O_112,N_2655,N_2581);
nand UO_113 (O_113,N_2550,N_2626);
and UO_114 (O_114,N_2432,N_2654);
nor UO_115 (O_115,N_2464,N_2939);
nand UO_116 (O_116,N_2512,N_2743);
nor UO_117 (O_117,N_2691,N_2582);
and UO_118 (O_118,N_2442,N_2507);
or UO_119 (O_119,N_2454,N_2900);
or UO_120 (O_120,N_2533,N_2838);
and UO_121 (O_121,N_2460,N_2410);
or UO_122 (O_122,N_2772,N_2566);
nand UO_123 (O_123,N_2481,N_2769);
nand UO_124 (O_124,N_2878,N_2403);
or UO_125 (O_125,N_2480,N_2943);
or UO_126 (O_126,N_2579,N_2849);
and UO_127 (O_127,N_2793,N_2814);
or UO_128 (O_128,N_2747,N_2721);
or UO_129 (O_129,N_2611,N_2586);
and UO_130 (O_130,N_2988,N_2625);
and UO_131 (O_131,N_2917,N_2677);
and UO_132 (O_132,N_2909,N_2639);
or UO_133 (O_133,N_2762,N_2433);
and UO_134 (O_134,N_2723,N_2877);
or UO_135 (O_135,N_2680,N_2633);
nor UO_136 (O_136,N_2485,N_2855);
or UO_137 (O_137,N_2426,N_2477);
nand UO_138 (O_138,N_2982,N_2563);
and UO_139 (O_139,N_2429,N_2950);
nor UO_140 (O_140,N_2746,N_2842);
or UO_141 (O_141,N_2535,N_2587);
nor UO_142 (O_142,N_2826,N_2699);
or UO_143 (O_143,N_2590,N_2979);
or UO_144 (O_144,N_2820,N_2899);
nor UO_145 (O_145,N_2732,N_2543);
nand UO_146 (O_146,N_2595,N_2472);
or UO_147 (O_147,N_2904,N_2882);
and UO_148 (O_148,N_2998,N_2607);
nor UO_149 (O_149,N_2521,N_2515);
nand UO_150 (O_150,N_2688,N_2511);
nor UO_151 (O_151,N_2748,N_2656);
nand UO_152 (O_152,N_2659,N_2873);
nand UO_153 (O_153,N_2896,N_2503);
nor UO_154 (O_154,N_2673,N_2952);
nor UO_155 (O_155,N_2856,N_2764);
or UO_156 (O_156,N_2766,N_2876);
and UO_157 (O_157,N_2627,N_2402);
and UO_158 (O_158,N_2887,N_2765);
or UO_159 (O_159,N_2514,N_2610);
nand UO_160 (O_160,N_2622,N_2905);
nand UO_161 (O_161,N_2782,N_2941);
xor UO_162 (O_162,N_2517,N_2662);
nor UO_163 (O_163,N_2730,N_2803);
and UO_164 (O_164,N_2594,N_2847);
nor UO_165 (O_165,N_2423,N_2713);
xnor UO_166 (O_166,N_2975,N_2986);
nand UO_167 (O_167,N_2522,N_2498);
nand UO_168 (O_168,N_2445,N_2453);
or UO_169 (O_169,N_2751,N_2455);
nor UO_170 (O_170,N_2598,N_2700);
nor UO_171 (O_171,N_2880,N_2632);
nor UO_172 (O_172,N_2792,N_2971);
and UO_173 (O_173,N_2490,N_2760);
and UO_174 (O_174,N_2439,N_2984);
and UO_175 (O_175,N_2494,N_2771);
and UO_176 (O_176,N_2537,N_2744);
or UO_177 (O_177,N_2890,N_2815);
nand UO_178 (O_178,N_2612,N_2650);
nor UO_179 (O_179,N_2526,N_2914);
and UO_180 (O_180,N_2461,N_2935);
and UO_181 (O_181,N_2518,N_2640);
and UO_182 (O_182,N_2861,N_2604);
and UO_183 (O_183,N_2615,N_2686);
or UO_184 (O_184,N_2802,N_2865);
or UO_185 (O_185,N_2745,N_2642);
or UO_186 (O_186,N_2451,N_2474);
or UO_187 (O_187,N_2555,N_2892);
and UO_188 (O_188,N_2953,N_2932);
and UO_189 (O_189,N_2409,N_2692);
nor UO_190 (O_190,N_2552,N_2556);
or UO_191 (O_191,N_2404,N_2412);
nor UO_192 (O_192,N_2491,N_2806);
and UO_193 (O_193,N_2467,N_2843);
and UO_194 (O_194,N_2891,N_2565);
nand UO_195 (O_195,N_2575,N_2479);
and UO_196 (O_196,N_2484,N_2836);
nor UO_197 (O_197,N_2962,N_2525);
and UO_198 (O_198,N_2821,N_2588);
and UO_199 (O_199,N_2546,N_2949);
xor UO_200 (O_200,N_2636,N_2805);
and UO_201 (O_201,N_2797,N_2724);
nor UO_202 (O_202,N_2715,N_2421);
or UO_203 (O_203,N_2411,N_2752);
nand UO_204 (O_204,N_2830,N_2502);
and UO_205 (O_205,N_2804,N_2463);
nor UO_206 (O_206,N_2510,N_2999);
nand UO_207 (O_207,N_2733,N_2902);
or UO_208 (O_208,N_2918,N_2985);
nand UO_209 (O_209,N_2435,N_2649);
nor UO_210 (O_210,N_2794,N_2407);
nor UO_211 (O_211,N_2860,N_2653);
or UO_212 (O_212,N_2660,N_2492);
and UO_213 (O_213,N_2476,N_2424);
and UO_214 (O_214,N_2405,N_2726);
and UO_215 (O_215,N_2725,N_2596);
and UO_216 (O_216,N_2506,N_2679);
or UO_217 (O_217,N_2906,N_2705);
and UO_218 (O_218,N_2413,N_2933);
or UO_219 (O_219,N_2967,N_2508);
and UO_220 (O_220,N_2997,N_2774);
xor UO_221 (O_221,N_2888,N_2839);
or UO_222 (O_222,N_2731,N_2509);
nor UO_223 (O_223,N_2578,N_2977);
nor UO_224 (O_224,N_2837,N_2644);
nand UO_225 (O_225,N_2996,N_2614);
or UO_226 (O_226,N_2583,N_2895);
or UO_227 (O_227,N_2983,N_2457);
or UO_228 (O_228,N_2824,N_2832);
nor UO_229 (O_229,N_2473,N_2894);
or UO_230 (O_230,N_2712,N_2758);
and UO_231 (O_231,N_2866,N_2446);
xor UO_232 (O_232,N_2929,N_2951);
or UO_233 (O_233,N_2930,N_2634);
or UO_234 (O_234,N_2577,N_2609);
and UO_235 (O_235,N_2568,N_2678);
nand UO_236 (O_236,N_2995,N_2978);
and UO_237 (O_237,N_2925,N_2665);
nand UO_238 (O_238,N_2924,N_2869);
or UO_239 (O_239,N_2913,N_2841);
nand UO_240 (O_240,N_2414,N_2738);
xor UO_241 (O_241,N_2846,N_2736);
and UO_242 (O_242,N_2716,N_2682);
nor UO_243 (O_243,N_2558,N_2475);
or UO_244 (O_244,N_2722,N_2819);
or UO_245 (O_245,N_2470,N_2671);
and UO_246 (O_246,N_2599,N_2696);
nand UO_247 (O_247,N_2450,N_2551);
or UO_248 (O_248,N_2714,N_2734);
nor UO_249 (O_249,N_2616,N_2663);
nor UO_250 (O_250,N_2489,N_2796);
and UO_251 (O_251,N_2670,N_2471);
xnor UO_252 (O_252,N_2547,N_2420);
nand UO_253 (O_253,N_2958,N_2488);
or UO_254 (O_254,N_2425,N_2693);
or UO_255 (O_255,N_2573,N_2901);
or UO_256 (O_256,N_2422,N_2823);
nand UO_257 (O_257,N_2927,N_2707);
or UO_258 (O_258,N_2592,N_2720);
or UO_259 (O_259,N_2844,N_2493);
nor UO_260 (O_260,N_2960,N_2915);
nor UO_261 (O_261,N_2750,N_2813);
nand UO_262 (O_262,N_2923,N_2879);
and UO_263 (O_263,N_2567,N_2605);
and UO_264 (O_264,N_2946,N_2749);
nand UO_265 (O_265,N_2739,N_2798);
nand UO_266 (O_266,N_2709,N_2401);
nor UO_267 (O_267,N_2912,N_2648);
nor UO_268 (O_268,N_2553,N_2931);
nor UO_269 (O_269,N_2637,N_2483);
xor UO_270 (O_270,N_2544,N_2676);
nand UO_271 (O_271,N_2940,N_2801);
nand UO_272 (O_272,N_2541,N_2666);
nor UO_273 (O_273,N_2589,N_2816);
nor UO_274 (O_274,N_2664,N_2702);
nor UO_275 (O_275,N_2948,N_2974);
nor UO_276 (O_276,N_2735,N_2466);
or UO_277 (O_277,N_2959,N_2831);
and UO_278 (O_278,N_2704,N_2808);
nand UO_279 (O_279,N_2871,N_2540);
or UO_280 (O_280,N_2870,N_2487);
and UO_281 (O_281,N_2495,N_2858);
or UO_282 (O_282,N_2668,N_2532);
or UO_283 (O_283,N_2777,N_2780);
nor UO_284 (O_284,N_2800,N_2829);
nor UO_285 (O_285,N_2576,N_2729);
nand UO_286 (O_286,N_2956,N_2608);
and UO_287 (O_287,N_2921,N_2628);
nand UO_288 (O_288,N_2499,N_2620);
nand UO_289 (O_289,N_2786,N_2431);
or UO_290 (O_290,N_2812,N_2559);
nand UO_291 (O_291,N_2408,N_2908);
nor UO_292 (O_292,N_2572,N_2687);
or UO_293 (O_293,N_2689,N_2427);
nand UO_294 (O_294,N_2969,N_2859);
nor UO_295 (O_295,N_2937,N_2776);
nand UO_296 (O_296,N_2597,N_2980);
nand UO_297 (O_297,N_2789,N_2624);
and UO_298 (O_298,N_2778,N_2513);
nor UO_299 (O_299,N_2428,N_2416);
nor UO_300 (O_300,N_2415,N_2743);
nor UO_301 (O_301,N_2861,N_2813);
nand UO_302 (O_302,N_2911,N_2507);
or UO_303 (O_303,N_2565,N_2833);
nand UO_304 (O_304,N_2843,N_2525);
nor UO_305 (O_305,N_2631,N_2431);
or UO_306 (O_306,N_2511,N_2991);
nand UO_307 (O_307,N_2473,N_2810);
and UO_308 (O_308,N_2632,N_2526);
and UO_309 (O_309,N_2459,N_2841);
or UO_310 (O_310,N_2537,N_2476);
and UO_311 (O_311,N_2786,N_2824);
and UO_312 (O_312,N_2967,N_2554);
and UO_313 (O_313,N_2546,N_2867);
and UO_314 (O_314,N_2916,N_2931);
xor UO_315 (O_315,N_2497,N_2479);
nand UO_316 (O_316,N_2720,N_2956);
nand UO_317 (O_317,N_2544,N_2788);
or UO_318 (O_318,N_2967,N_2861);
nor UO_319 (O_319,N_2880,N_2794);
and UO_320 (O_320,N_2653,N_2442);
and UO_321 (O_321,N_2699,N_2776);
or UO_322 (O_322,N_2747,N_2895);
nand UO_323 (O_323,N_2725,N_2910);
and UO_324 (O_324,N_2733,N_2486);
and UO_325 (O_325,N_2660,N_2682);
nor UO_326 (O_326,N_2682,N_2948);
nand UO_327 (O_327,N_2955,N_2775);
and UO_328 (O_328,N_2505,N_2793);
nor UO_329 (O_329,N_2615,N_2585);
nor UO_330 (O_330,N_2722,N_2915);
or UO_331 (O_331,N_2437,N_2751);
or UO_332 (O_332,N_2830,N_2537);
nand UO_333 (O_333,N_2518,N_2725);
nand UO_334 (O_334,N_2734,N_2726);
nor UO_335 (O_335,N_2447,N_2409);
xnor UO_336 (O_336,N_2523,N_2828);
and UO_337 (O_337,N_2796,N_2851);
or UO_338 (O_338,N_2604,N_2669);
nand UO_339 (O_339,N_2889,N_2560);
and UO_340 (O_340,N_2809,N_2584);
nor UO_341 (O_341,N_2758,N_2411);
or UO_342 (O_342,N_2469,N_2713);
nor UO_343 (O_343,N_2658,N_2724);
or UO_344 (O_344,N_2947,N_2510);
nand UO_345 (O_345,N_2893,N_2593);
nor UO_346 (O_346,N_2866,N_2539);
or UO_347 (O_347,N_2458,N_2985);
nor UO_348 (O_348,N_2574,N_2818);
or UO_349 (O_349,N_2633,N_2799);
nor UO_350 (O_350,N_2431,N_2425);
nor UO_351 (O_351,N_2669,N_2989);
nand UO_352 (O_352,N_2646,N_2577);
nand UO_353 (O_353,N_2882,N_2533);
and UO_354 (O_354,N_2981,N_2968);
nand UO_355 (O_355,N_2843,N_2665);
nand UO_356 (O_356,N_2718,N_2917);
nor UO_357 (O_357,N_2592,N_2481);
nand UO_358 (O_358,N_2966,N_2602);
nor UO_359 (O_359,N_2790,N_2976);
nor UO_360 (O_360,N_2978,N_2568);
nor UO_361 (O_361,N_2991,N_2461);
nand UO_362 (O_362,N_2575,N_2938);
nand UO_363 (O_363,N_2854,N_2589);
nor UO_364 (O_364,N_2720,N_2760);
and UO_365 (O_365,N_2643,N_2824);
or UO_366 (O_366,N_2723,N_2849);
nand UO_367 (O_367,N_2447,N_2487);
or UO_368 (O_368,N_2862,N_2530);
nand UO_369 (O_369,N_2636,N_2957);
xor UO_370 (O_370,N_2794,N_2813);
nor UO_371 (O_371,N_2533,N_2535);
nand UO_372 (O_372,N_2986,N_2484);
or UO_373 (O_373,N_2678,N_2919);
and UO_374 (O_374,N_2915,N_2930);
nand UO_375 (O_375,N_2768,N_2836);
nor UO_376 (O_376,N_2904,N_2556);
and UO_377 (O_377,N_2896,N_2764);
nand UO_378 (O_378,N_2755,N_2901);
or UO_379 (O_379,N_2444,N_2841);
xor UO_380 (O_380,N_2968,N_2503);
nand UO_381 (O_381,N_2748,N_2498);
or UO_382 (O_382,N_2681,N_2835);
and UO_383 (O_383,N_2503,N_2827);
or UO_384 (O_384,N_2788,N_2554);
nand UO_385 (O_385,N_2826,N_2881);
or UO_386 (O_386,N_2813,N_2836);
or UO_387 (O_387,N_2590,N_2883);
and UO_388 (O_388,N_2856,N_2925);
nand UO_389 (O_389,N_2880,N_2922);
nand UO_390 (O_390,N_2700,N_2781);
and UO_391 (O_391,N_2652,N_2490);
nor UO_392 (O_392,N_2846,N_2508);
nand UO_393 (O_393,N_2837,N_2554);
or UO_394 (O_394,N_2874,N_2665);
or UO_395 (O_395,N_2955,N_2970);
nand UO_396 (O_396,N_2470,N_2544);
or UO_397 (O_397,N_2708,N_2783);
and UO_398 (O_398,N_2997,N_2496);
nand UO_399 (O_399,N_2959,N_2781);
or UO_400 (O_400,N_2675,N_2508);
nand UO_401 (O_401,N_2520,N_2466);
nor UO_402 (O_402,N_2939,N_2519);
or UO_403 (O_403,N_2809,N_2592);
or UO_404 (O_404,N_2644,N_2784);
and UO_405 (O_405,N_2923,N_2421);
nand UO_406 (O_406,N_2477,N_2638);
nand UO_407 (O_407,N_2702,N_2419);
nand UO_408 (O_408,N_2970,N_2597);
or UO_409 (O_409,N_2629,N_2940);
nor UO_410 (O_410,N_2870,N_2532);
nand UO_411 (O_411,N_2645,N_2556);
nand UO_412 (O_412,N_2575,N_2993);
and UO_413 (O_413,N_2895,N_2901);
nor UO_414 (O_414,N_2878,N_2923);
nand UO_415 (O_415,N_2711,N_2642);
and UO_416 (O_416,N_2775,N_2708);
nand UO_417 (O_417,N_2612,N_2971);
and UO_418 (O_418,N_2873,N_2433);
nor UO_419 (O_419,N_2752,N_2558);
and UO_420 (O_420,N_2668,N_2596);
nor UO_421 (O_421,N_2689,N_2706);
nor UO_422 (O_422,N_2996,N_2976);
or UO_423 (O_423,N_2638,N_2504);
and UO_424 (O_424,N_2934,N_2706);
or UO_425 (O_425,N_2502,N_2725);
or UO_426 (O_426,N_2986,N_2948);
nand UO_427 (O_427,N_2645,N_2566);
nor UO_428 (O_428,N_2496,N_2574);
nand UO_429 (O_429,N_2632,N_2696);
nor UO_430 (O_430,N_2794,N_2471);
nor UO_431 (O_431,N_2453,N_2879);
or UO_432 (O_432,N_2819,N_2970);
and UO_433 (O_433,N_2791,N_2961);
nand UO_434 (O_434,N_2480,N_2605);
nor UO_435 (O_435,N_2512,N_2948);
nor UO_436 (O_436,N_2692,N_2842);
nand UO_437 (O_437,N_2781,N_2603);
and UO_438 (O_438,N_2791,N_2946);
nand UO_439 (O_439,N_2778,N_2887);
or UO_440 (O_440,N_2885,N_2836);
nor UO_441 (O_441,N_2851,N_2793);
nand UO_442 (O_442,N_2418,N_2850);
nor UO_443 (O_443,N_2789,N_2696);
or UO_444 (O_444,N_2806,N_2557);
or UO_445 (O_445,N_2525,N_2769);
nor UO_446 (O_446,N_2622,N_2890);
nor UO_447 (O_447,N_2564,N_2662);
nand UO_448 (O_448,N_2792,N_2435);
and UO_449 (O_449,N_2569,N_2775);
nand UO_450 (O_450,N_2548,N_2731);
nand UO_451 (O_451,N_2448,N_2524);
nand UO_452 (O_452,N_2596,N_2424);
nand UO_453 (O_453,N_2856,N_2563);
or UO_454 (O_454,N_2476,N_2597);
xnor UO_455 (O_455,N_2979,N_2861);
and UO_456 (O_456,N_2586,N_2857);
and UO_457 (O_457,N_2496,N_2855);
nor UO_458 (O_458,N_2484,N_2894);
nor UO_459 (O_459,N_2467,N_2502);
nor UO_460 (O_460,N_2621,N_2755);
nor UO_461 (O_461,N_2430,N_2520);
or UO_462 (O_462,N_2953,N_2885);
or UO_463 (O_463,N_2532,N_2563);
and UO_464 (O_464,N_2535,N_2476);
nor UO_465 (O_465,N_2695,N_2553);
nand UO_466 (O_466,N_2599,N_2619);
nor UO_467 (O_467,N_2638,N_2654);
nand UO_468 (O_468,N_2653,N_2762);
and UO_469 (O_469,N_2984,N_2936);
or UO_470 (O_470,N_2514,N_2570);
and UO_471 (O_471,N_2883,N_2609);
nor UO_472 (O_472,N_2773,N_2587);
or UO_473 (O_473,N_2802,N_2805);
or UO_474 (O_474,N_2651,N_2776);
and UO_475 (O_475,N_2748,N_2863);
nand UO_476 (O_476,N_2705,N_2676);
and UO_477 (O_477,N_2771,N_2697);
or UO_478 (O_478,N_2963,N_2506);
nand UO_479 (O_479,N_2592,N_2660);
xnor UO_480 (O_480,N_2544,N_2947);
nand UO_481 (O_481,N_2412,N_2634);
and UO_482 (O_482,N_2739,N_2514);
xnor UO_483 (O_483,N_2753,N_2431);
and UO_484 (O_484,N_2903,N_2723);
nand UO_485 (O_485,N_2999,N_2526);
nand UO_486 (O_486,N_2785,N_2757);
and UO_487 (O_487,N_2795,N_2629);
nand UO_488 (O_488,N_2620,N_2835);
nor UO_489 (O_489,N_2772,N_2933);
nor UO_490 (O_490,N_2840,N_2401);
and UO_491 (O_491,N_2455,N_2622);
nand UO_492 (O_492,N_2992,N_2462);
or UO_493 (O_493,N_2548,N_2576);
or UO_494 (O_494,N_2894,N_2621);
and UO_495 (O_495,N_2448,N_2854);
and UO_496 (O_496,N_2468,N_2995);
or UO_497 (O_497,N_2864,N_2650);
and UO_498 (O_498,N_2664,N_2553);
nand UO_499 (O_499,N_2892,N_2767);
endmodule