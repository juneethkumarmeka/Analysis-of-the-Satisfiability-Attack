module basic_5000_50000_5000_25_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
or U0 (N_0,In_2774,In_4535);
nand U1 (N_1,In_2490,In_213);
nor U2 (N_2,In_1941,In_861);
xnor U3 (N_3,In_2660,In_4805);
xnor U4 (N_4,In_730,In_4741);
nand U5 (N_5,In_3220,In_4892);
or U6 (N_6,In_4485,In_2676);
or U7 (N_7,In_4197,In_510);
or U8 (N_8,In_160,In_2870);
and U9 (N_9,In_4942,In_3489);
nor U10 (N_10,In_181,In_3057);
nand U11 (N_11,In_1672,In_1559);
nor U12 (N_12,In_663,In_4771);
and U13 (N_13,In_4593,In_2250);
xor U14 (N_14,In_4159,In_1150);
nand U15 (N_15,In_4876,In_4281);
nand U16 (N_16,In_2419,In_1304);
nand U17 (N_17,In_505,In_1533);
nand U18 (N_18,In_790,In_561);
or U19 (N_19,In_2692,In_4732);
xnor U20 (N_20,In_4763,In_2390);
and U21 (N_21,In_1510,In_3235);
and U22 (N_22,In_3447,In_954);
nor U23 (N_23,In_4565,In_3246);
nand U24 (N_24,In_2518,In_865);
xor U25 (N_25,In_2000,In_1200);
xor U26 (N_26,In_3405,In_1957);
xor U27 (N_27,In_3641,In_203);
nor U28 (N_28,In_3066,In_190);
nand U29 (N_29,In_1347,In_174);
or U30 (N_30,In_3393,In_302);
nand U31 (N_31,In_224,In_1246);
nand U32 (N_32,In_1903,In_4868);
xor U33 (N_33,In_2929,In_4486);
xor U34 (N_34,In_66,In_1290);
xnor U35 (N_35,In_1016,In_284);
or U36 (N_36,In_3963,In_4389);
xnor U37 (N_37,In_1373,In_4970);
or U38 (N_38,In_73,In_4765);
or U39 (N_39,In_4304,In_2127);
or U40 (N_40,In_765,In_4896);
and U41 (N_41,In_703,In_2142);
nor U42 (N_42,In_4110,In_1588);
xnor U43 (N_43,In_2824,In_175);
and U44 (N_44,In_3889,In_642);
and U45 (N_45,In_432,In_4267);
and U46 (N_46,In_111,In_1499);
nand U47 (N_47,In_3098,In_1942);
or U48 (N_48,In_4540,In_3189);
and U49 (N_49,In_1963,In_110);
nor U50 (N_50,In_1688,In_4716);
and U51 (N_51,In_231,In_3542);
nor U52 (N_52,In_2222,In_2117);
nor U53 (N_53,In_451,In_4012);
nand U54 (N_54,In_1766,In_4826);
nand U55 (N_55,In_1974,In_3179);
xnor U56 (N_56,In_4562,In_4632);
nor U57 (N_57,In_3031,In_3032);
nor U58 (N_58,In_1561,In_2878);
xnor U59 (N_59,In_3941,In_2916);
xnor U60 (N_60,In_953,In_3910);
and U61 (N_61,In_273,In_3666);
and U62 (N_62,In_4794,In_454);
and U63 (N_63,In_4994,In_2011);
nand U64 (N_64,In_2778,In_4891);
nor U65 (N_65,In_4909,In_2082);
nand U66 (N_66,In_1548,In_341);
nor U67 (N_67,In_1949,In_4627);
xor U68 (N_68,In_1118,In_4835);
or U69 (N_69,In_2183,In_4974);
nor U70 (N_70,In_2372,In_4704);
nor U71 (N_71,In_1295,In_3525);
nor U72 (N_72,In_4548,In_1564);
nand U73 (N_73,In_4167,In_3712);
and U74 (N_74,In_134,In_4407);
or U75 (N_75,In_3343,In_21);
nor U76 (N_76,In_325,In_1115);
and U77 (N_77,In_1123,In_4984);
xnor U78 (N_78,In_3109,In_1946);
nor U79 (N_79,In_4405,In_1686);
or U80 (N_80,In_4599,In_4946);
nand U81 (N_81,In_408,In_2963);
nand U82 (N_82,In_3578,In_4039);
nor U83 (N_83,In_3852,In_1569);
or U84 (N_84,In_2683,In_564);
or U85 (N_85,In_35,In_3789);
or U86 (N_86,In_715,In_4662);
nor U87 (N_87,In_2513,In_742);
nand U88 (N_88,In_2242,In_1212);
xor U89 (N_89,In_2131,In_4708);
and U90 (N_90,In_4682,In_344);
or U91 (N_91,In_4888,In_3243);
xnor U92 (N_92,In_4742,In_1233);
or U93 (N_93,In_2861,In_4262);
nor U94 (N_94,In_726,In_2704);
nor U95 (N_95,In_4426,In_4388);
xor U96 (N_96,In_1558,In_1959);
nor U97 (N_97,In_2087,In_1495);
and U98 (N_98,In_3947,In_138);
and U99 (N_99,In_2305,In_452);
nor U100 (N_100,In_3239,In_3352);
and U101 (N_101,In_1267,In_1969);
nor U102 (N_102,In_1129,In_3142);
xor U103 (N_103,In_4484,In_4014);
and U104 (N_104,In_792,In_2693);
xnor U105 (N_105,In_1802,In_4344);
nand U106 (N_106,In_1813,In_166);
xnor U107 (N_107,In_3307,In_4506);
xnor U108 (N_108,In_4639,In_3194);
and U109 (N_109,In_1114,In_2874);
or U110 (N_110,In_1448,In_2610);
or U111 (N_111,In_412,In_2926);
xnor U112 (N_112,In_2327,In_2005);
or U113 (N_113,In_4218,In_3378);
nor U114 (N_114,In_1216,In_3533);
and U115 (N_115,In_4057,In_1798);
nand U116 (N_116,In_1932,In_2915);
xnor U117 (N_117,In_617,In_938);
xor U118 (N_118,In_1539,In_550);
and U119 (N_119,In_3135,In_2418);
and U120 (N_120,In_3391,In_2709);
xor U121 (N_121,In_128,In_2149);
nor U122 (N_122,In_2954,In_3455);
xnor U123 (N_123,In_533,In_1687);
nor U124 (N_124,In_930,In_1536);
or U125 (N_125,In_2734,In_2323);
nor U126 (N_126,In_2401,In_1498);
and U127 (N_127,In_1938,In_3071);
xnor U128 (N_128,In_655,In_3012);
nor U129 (N_129,In_973,In_3281);
nand U130 (N_130,In_3065,In_1742);
or U131 (N_131,In_3959,In_2066);
nand U132 (N_132,In_2231,In_1286);
nand U133 (N_133,In_3260,In_4071);
nor U134 (N_134,In_1836,In_1840);
nor U135 (N_135,In_3736,In_4203);
nand U136 (N_136,In_4550,In_72);
nor U137 (N_137,In_2900,In_3100);
nand U138 (N_138,In_4130,In_976);
nor U139 (N_139,In_1426,In_2135);
nor U140 (N_140,In_4859,In_1215);
or U141 (N_141,In_4224,In_754);
nand U142 (N_142,In_3492,In_363);
xnor U143 (N_143,In_1638,In_3766);
xnor U144 (N_144,In_3161,In_60);
or U145 (N_145,In_415,In_1505);
nand U146 (N_146,In_1477,In_2852);
nand U147 (N_147,In_1833,In_4236);
nor U148 (N_148,In_4033,In_3844);
xor U149 (N_149,In_3141,In_1240);
xnor U150 (N_150,In_4529,In_2735);
or U151 (N_151,In_3017,In_4844);
nand U152 (N_152,In_4427,In_631);
or U153 (N_153,In_1772,In_1827);
nor U154 (N_154,In_2786,In_4710);
and U155 (N_155,In_3070,In_154);
xor U156 (N_156,In_4748,In_2634);
and U157 (N_157,In_4144,In_3202);
nand U158 (N_158,In_4059,In_3210);
xor U159 (N_159,In_4845,In_4425);
nand U160 (N_160,In_2985,In_4040);
xor U161 (N_161,In_568,In_4079);
xor U162 (N_162,In_3322,In_3565);
nand U163 (N_163,In_724,In_991);
and U164 (N_164,In_1951,In_3116);
and U165 (N_165,In_4368,In_1829);
xnor U166 (N_166,In_4920,In_1610);
xor U167 (N_167,In_3277,In_3458);
nand U168 (N_168,In_33,In_1665);
xor U169 (N_169,In_1487,In_1762);
nand U170 (N_170,In_3150,In_1668);
nor U171 (N_171,In_3536,In_643);
nand U172 (N_172,In_2883,In_3512);
or U173 (N_173,In_95,In_4754);
or U174 (N_174,In_878,In_4);
xnor U175 (N_175,In_3808,In_4515);
and U176 (N_176,In_2072,In_43);
nand U177 (N_177,In_4557,In_404);
and U178 (N_178,In_1245,In_1079);
nand U179 (N_179,In_3932,In_2485);
nand U180 (N_180,In_4701,In_4596);
or U181 (N_181,In_4969,In_4229);
nor U182 (N_182,In_3511,In_4923);
and U183 (N_183,In_588,In_1484);
nor U184 (N_184,In_3462,In_3681);
xnor U185 (N_185,In_4310,In_301);
xnor U186 (N_186,In_600,In_984);
or U187 (N_187,In_579,In_4044);
xnor U188 (N_188,In_4465,In_3154);
and U189 (N_189,In_4105,In_3242);
nand U190 (N_190,In_96,In_2188);
nand U191 (N_191,In_558,In_42);
nor U192 (N_192,In_4987,In_3807);
nor U193 (N_193,In_3625,In_4201);
xor U194 (N_194,In_842,In_3203);
xnor U195 (N_195,In_2342,In_4204);
nand U196 (N_196,In_1884,In_2393);
nand U197 (N_197,In_3845,In_3323);
nor U198 (N_198,In_2218,In_3927);
or U199 (N_199,In_4966,In_4968);
and U200 (N_200,In_556,In_628);
nor U201 (N_201,In_3521,In_2541);
nor U202 (N_202,In_2351,In_2416);
or U203 (N_203,In_4069,In_1117);
and U204 (N_204,In_3174,In_1193);
nand U205 (N_205,In_534,In_1977);
xor U206 (N_206,In_4861,In_1526);
nor U207 (N_207,In_565,In_3482);
nor U208 (N_208,In_4660,In_4193);
xor U209 (N_209,In_3309,In_4017);
and U210 (N_210,In_1708,In_601);
or U211 (N_211,In_312,In_4330);
nor U212 (N_212,In_1981,In_2946);
xor U213 (N_213,In_4037,In_4125);
nor U214 (N_214,In_2332,In_710);
or U215 (N_215,In_581,In_4084);
nand U216 (N_216,In_1001,In_3073);
xor U217 (N_217,In_908,In_319);
xor U218 (N_218,In_654,In_3812);
nand U219 (N_219,In_398,In_2320);
xnor U220 (N_220,In_3125,In_1392);
nor U221 (N_221,In_3048,In_2456);
nand U222 (N_222,In_3782,In_4703);
nand U223 (N_223,In_3774,In_996);
nand U224 (N_224,In_13,In_4364);
or U225 (N_225,In_1305,In_2803);
and U226 (N_226,In_2615,In_92);
nand U227 (N_227,In_2220,In_3158);
xor U228 (N_228,In_4433,In_477);
nor U229 (N_229,In_833,In_1219);
nand U230 (N_230,In_1275,In_1489);
nor U231 (N_231,In_3600,In_2088);
xor U232 (N_232,In_1741,In_941);
or U233 (N_233,In_909,In_2689);
xor U234 (N_234,In_4509,In_488);
or U235 (N_235,In_1650,In_3215);
nor U236 (N_236,In_1624,In_4996);
nor U237 (N_237,In_4603,In_468);
or U238 (N_238,In_1707,In_4027);
nand U239 (N_239,In_3706,In_2367);
nand U240 (N_240,In_622,In_2442);
nor U241 (N_241,In_2528,In_2617);
or U242 (N_242,In_1675,In_4695);
or U243 (N_243,In_3701,In_2132);
and U244 (N_244,In_989,In_2801);
nor U245 (N_245,In_3185,In_1756);
xnor U246 (N_246,In_808,In_3524);
xnor U247 (N_247,In_1660,In_1398);
and U248 (N_248,In_2046,In_3126);
nand U249 (N_249,In_2715,In_883);
nor U250 (N_250,In_1481,In_937);
nor U251 (N_251,In_2007,In_801);
and U252 (N_252,In_4434,In_2873);
or U253 (N_253,In_725,In_1594);
and U254 (N_254,In_444,In_649);
xor U255 (N_255,In_3919,In_2821);
and U256 (N_256,In_1099,In_1980);
or U257 (N_257,In_1158,In_2204);
or U258 (N_258,In_4463,In_3561);
nor U259 (N_259,In_3668,In_1352);
nor U260 (N_260,In_2872,In_4683);
or U261 (N_261,In_504,In_2172);
nand U262 (N_262,In_233,In_1080);
nand U263 (N_263,In_3629,In_4808);
and U264 (N_264,In_2221,In_2882);
xor U265 (N_265,In_4537,In_1256);
and U266 (N_266,In_4643,In_3897);
or U267 (N_267,In_618,In_557);
and U268 (N_268,In_38,In_2616);
nand U269 (N_269,In_3218,In_590);
xnor U270 (N_270,In_689,In_193);
nor U271 (N_271,In_3571,In_1435);
and U272 (N_272,In_2487,In_3764);
or U273 (N_273,In_2939,In_3716);
nor U274 (N_274,In_3484,In_3016);
nor U275 (N_275,In_1143,In_4390);
or U276 (N_276,In_791,In_1783);
xor U277 (N_277,In_3157,In_3957);
and U278 (N_278,In_3357,In_1655);
xor U279 (N_279,In_2414,In_2607);
nor U280 (N_280,In_1621,In_1329);
nor U281 (N_281,In_783,In_2802);
xor U282 (N_282,In_1272,In_4099);
or U283 (N_283,In_380,In_2094);
and U284 (N_284,In_604,In_4782);
xnor U285 (N_285,In_553,In_2745);
nand U286 (N_286,In_1933,In_1050);
or U287 (N_287,In_971,In_212);
nand U288 (N_288,In_2879,In_4688);
and U289 (N_289,In_2769,In_104);
nand U290 (N_290,In_1844,In_4823);
xor U291 (N_291,In_4962,In_3693);
or U292 (N_292,In_1371,In_2090);
and U293 (N_293,In_3193,In_370);
nand U294 (N_294,In_1796,In_364);
or U295 (N_295,In_3900,In_1341);
nor U296 (N_296,In_4690,In_3232);
or U297 (N_297,In_3181,In_100);
or U298 (N_298,In_3334,In_1644);
nor U299 (N_299,In_1464,In_3652);
and U300 (N_300,In_3702,In_3597);
xor U301 (N_301,In_4792,In_2421);
xnor U302 (N_302,In_1449,In_491);
or U303 (N_303,In_3086,In_1051);
and U304 (N_304,In_2105,In_3035);
nand U305 (N_305,In_2399,In_2428);
or U306 (N_306,In_4739,In_4553);
xnor U307 (N_307,In_2259,In_2994);
xnor U308 (N_308,In_1091,In_769);
or U309 (N_309,In_1557,In_1750);
xnor U310 (N_310,In_3544,In_4349);
nor U311 (N_311,In_2101,In_3167);
nor U312 (N_312,In_4004,In_2848);
nand U313 (N_313,In_3560,In_205);
nor U314 (N_314,In_3172,In_986);
xor U315 (N_315,In_1178,In_536);
nand U316 (N_316,In_2590,In_3251);
or U317 (N_317,In_2891,In_3526);
xnor U318 (N_318,In_1088,In_799);
nand U319 (N_319,In_308,In_409);
nand U320 (N_320,In_247,In_3984);
nor U321 (N_321,In_830,In_4856);
nor U322 (N_322,In_220,In_50);
and U323 (N_323,In_320,In_2316);
xor U324 (N_324,In_260,In_4293);
nand U325 (N_325,In_2405,In_4897);
or U326 (N_326,In_4761,In_3926);
xor U327 (N_327,In_3691,In_775);
or U328 (N_328,In_1623,In_3199);
and U329 (N_329,In_875,In_4294);
nor U330 (N_330,In_2196,In_2533);
xnor U331 (N_331,In_2261,In_90);
and U332 (N_332,In_2168,In_137);
and U333 (N_333,In_1478,In_161);
nand U334 (N_334,In_414,In_47);
xnor U335 (N_335,In_3383,In_3865);
or U336 (N_336,In_841,In_2628);
xnor U337 (N_337,In_2760,In_4881);
xor U338 (N_338,In_3553,In_4104);
or U339 (N_339,In_2136,In_3420);
nor U340 (N_340,In_2458,In_3392);
xor U341 (N_341,In_4787,In_2677);
nand U342 (N_342,In_3052,In_854);
or U343 (N_343,In_4939,In_2568);
or U344 (N_344,In_3505,In_1622);
xor U345 (N_345,In_3358,In_3087);
xnor U346 (N_346,In_1599,In_4572);
nor U347 (N_347,In_4722,In_3440);
nand U348 (N_348,In_3223,In_276);
nand U349 (N_349,In_179,In_2104);
nand U350 (N_350,In_3513,In_4519);
or U351 (N_351,In_2181,In_1474);
nor U352 (N_352,In_2850,In_1364);
nand U353 (N_353,In_4948,In_4614);
or U354 (N_354,In_3964,In_1389);
xor U355 (N_355,In_2252,In_143);
and U356 (N_356,In_1731,In_419);
nand U357 (N_357,In_1411,In_4827);
nor U358 (N_358,In_1652,In_2353);
xor U359 (N_359,In_734,In_4882);
or U360 (N_360,In_2571,In_3345);
and U361 (N_361,In_1345,In_695);
nand U362 (N_362,In_3463,In_3248);
or U363 (N_363,In_4395,In_956);
xor U364 (N_364,In_8,In_3833);
nor U365 (N_365,In_3403,In_3213);
nand U366 (N_366,In_2762,In_674);
xor U367 (N_367,In_4333,In_658);
nand U368 (N_368,In_1704,In_2678);
or U369 (N_369,In_787,In_2018);
xnor U370 (N_370,In_241,In_3617);
nand U371 (N_371,In_1094,In_3424);
nor U372 (N_372,In_3282,In_1175);
or U373 (N_373,In_4534,In_1547);
nand U374 (N_374,In_3990,In_4290);
or U375 (N_375,In_4610,In_3559);
or U376 (N_376,In_292,In_4691);
nor U377 (N_377,In_1460,In_2482);
or U378 (N_378,In_1319,In_11);
and U379 (N_379,In_3911,In_321);
and U380 (N_380,In_1683,In_4905);
nor U381 (N_381,In_294,In_632);
or U382 (N_382,In_4146,In_2161);
nor U383 (N_383,In_4865,In_3822);
nand U384 (N_384,In_1281,In_1021);
and U385 (N_385,In_1191,In_3953);
or U386 (N_386,In_4259,In_2956);
nor U387 (N_387,In_2731,In_2603);
and U388 (N_388,In_1238,In_1823);
or U389 (N_389,In_2549,In_108);
nand U390 (N_390,In_3880,In_2996);
nand U391 (N_391,In_3648,In_2927);
xor U392 (N_392,In_771,In_1689);
xnor U393 (N_393,In_1887,In_4006);
or U394 (N_394,In_4833,In_2065);
nor U395 (N_395,In_3955,In_3022);
or U396 (N_396,In_3175,In_1553);
and U397 (N_397,In_4331,In_117);
or U398 (N_398,In_91,In_4337);
nor U399 (N_399,In_744,In_2842);
and U400 (N_400,In_3139,In_3754);
and U401 (N_401,In_3208,In_1537);
nand U402 (N_402,In_2322,In_4480);
nand U403 (N_403,In_2108,In_267);
nor U404 (N_404,In_3201,In_322);
or U405 (N_405,In_1781,In_1111);
and U406 (N_406,In_24,In_4371);
nor U407 (N_407,In_1615,In_3972);
and U408 (N_408,In_1424,In_2349);
and U409 (N_409,In_159,In_2256);
and U410 (N_410,In_493,In_4589);
xor U411 (N_411,In_3237,In_2903);
or U412 (N_412,In_229,In_4119);
nor U413 (N_413,In_1112,In_1782);
xor U414 (N_414,In_1493,In_2575);
nor U415 (N_415,In_677,In_3169);
nand U416 (N_416,In_2448,In_2373);
or U417 (N_417,In_1183,In_7);
xor U418 (N_418,In_2701,In_2730);
nand U419 (N_419,In_2404,In_3615);
and U420 (N_420,In_4212,In_1078);
or U421 (N_421,In_4047,In_862);
and U422 (N_422,In_3234,In_3620);
nor U423 (N_423,In_3662,In_3661);
nand U424 (N_424,In_2712,In_2667);
nor U425 (N_425,In_913,In_1882);
and U426 (N_426,In_167,In_2481);
xor U427 (N_427,In_2566,In_3187);
or U428 (N_428,In_2649,In_599);
nor U429 (N_429,In_1181,In_3831);
and U430 (N_430,In_1375,In_1948);
nor U431 (N_431,In_4776,In_3388);
nand U432 (N_432,In_3084,In_2330);
nor U433 (N_433,In_1230,In_1223);
or U434 (N_434,In_1832,In_1144);
or U435 (N_435,In_3456,In_2656);
or U436 (N_436,In_442,In_1595);
nand U437 (N_437,In_2889,In_4579);
xor U438 (N_438,In_2306,In_1788);
or U439 (N_439,In_53,In_3450);
or U440 (N_440,In_3399,In_2158);
or U441 (N_441,In_2284,In_2647);
nor U442 (N_442,In_196,In_2641);
nand U443 (N_443,In_4911,In_639);
and U444 (N_444,In_1298,In_4080);
xnor U445 (N_445,In_876,In_3504);
and U446 (N_446,In_79,In_3532);
or U447 (N_447,In_1086,In_3397);
nand U448 (N_448,In_3614,In_3777);
or U449 (N_449,In_2999,In_424);
nor U450 (N_450,In_4820,In_1755);
nand U451 (N_451,In_3847,In_1355);
and U452 (N_452,In_465,In_4789);
and U453 (N_453,In_4286,In_157);
xor U454 (N_454,In_687,In_3832);
nor U455 (N_455,In_484,In_4387);
nor U456 (N_456,In_1972,In_805);
nand U457 (N_457,In_4957,In_1254);
nand U458 (N_458,In_957,In_317);
and U459 (N_459,In_3912,In_1578);
or U460 (N_460,In_848,In_4437);
nor U461 (N_461,In_1771,In_2075);
nor U462 (N_462,In_4258,In_2097);
nand U463 (N_463,In_54,In_4618);
xnor U464 (N_464,In_3421,In_4185);
xnor U465 (N_465,In_3138,In_1470);
or U466 (N_466,In_4490,In_1242);
xnor U467 (N_467,In_1761,In_2292);
nand U468 (N_468,In_4421,In_1868);
and U469 (N_469,In_2076,In_4800);
nor U470 (N_470,In_2394,In_2074);
nand U471 (N_471,In_136,In_1330);
or U472 (N_472,In_4903,In_2800);
nor U473 (N_473,In_745,In_4275);
and U474 (N_474,In_4001,In_2720);
nand U475 (N_475,In_1459,In_4809);
or U476 (N_476,In_4680,In_2278);
and U477 (N_477,In_4539,In_3030);
nor U478 (N_478,In_2875,In_2860);
nand U479 (N_479,In_3800,In_4738);
xnor U480 (N_480,In_2589,In_1812);
and U481 (N_481,In_4450,In_3036);
or U482 (N_482,In_4947,In_1185);
nor U483 (N_483,In_4819,In_4894);
nor U484 (N_484,In_2546,In_3904);
xor U485 (N_485,In_1285,In_4278);
or U486 (N_486,In_4992,In_1187);
nand U487 (N_487,In_4462,In_3163);
and U488 (N_488,In_2558,In_767);
or U489 (N_489,In_4577,In_3933);
or U490 (N_490,In_1611,In_3222);
nand U491 (N_491,In_2449,In_4210);
xnor U492 (N_492,In_3688,In_188);
and U493 (N_493,In_3453,In_44);
nand U494 (N_494,In_2832,In_3209);
or U495 (N_495,In_3594,In_4009);
and U496 (N_496,In_4875,In_1930);
nor U497 (N_497,In_2780,In_3806);
or U498 (N_498,In_439,In_3628);
nor U499 (N_499,In_4842,In_3770);
nor U500 (N_500,In_122,In_812);
nor U501 (N_501,In_4343,In_4678);
nor U502 (N_502,In_2344,In_4404);
nand U503 (N_503,In_4273,In_4724);
nor U504 (N_504,In_3180,In_3680);
or U505 (N_505,In_1726,In_526);
xnor U506 (N_506,In_1502,In_1584);
xor U507 (N_507,In_339,In_1306);
or U508 (N_508,In_925,In_4309);
nand U509 (N_509,In_3864,In_4482);
xor U510 (N_510,In_2992,In_2846);
or U511 (N_511,In_4220,In_2896);
and U512 (N_512,In_3105,In_3316);
and U513 (N_513,In_2671,In_1596);
xnor U514 (N_514,In_2425,In_215);
and U515 (N_515,In_4366,In_2455);
and U516 (N_516,In_2744,In_192);
or U517 (N_517,In_4325,In_389);
xnor U518 (N_518,In_4336,In_459);
or U519 (N_519,In_1702,In_4569);
nor U520 (N_520,In_2480,In_2417);
nand U521 (N_521,In_171,In_2548);
nand U522 (N_522,In_944,In_3305);
xor U523 (N_523,In_713,In_1432);
and U524 (N_524,In_2947,In_3233);
or U525 (N_525,In_1962,In_1433);
nand U526 (N_526,In_311,In_4908);
and U527 (N_527,In_4731,In_1934);
or U528 (N_528,In_4866,In_383);
nor U529 (N_529,In_2391,In_3460);
xor U530 (N_530,In_2974,In_1857);
nor U531 (N_531,In_3520,In_4661);
and U532 (N_532,In_978,In_1579);
and U533 (N_533,In_2206,In_348);
and U534 (N_534,In_4062,In_1437);
nor U535 (N_535,In_1989,In_3534);
xor U536 (N_536,In_2049,In_1430);
nor U537 (N_537,In_2343,In_4452);
nor U538 (N_538,In_4757,In_4502);
or U539 (N_539,In_1024,In_3500);
or U540 (N_540,In_3756,In_3278);
or U541 (N_541,In_3651,In_3224);
nor U542 (N_542,In_2907,In_1785);
nand U543 (N_543,In_388,In_2489);
and U544 (N_544,In_1363,In_2569);
nor U545 (N_545,In_2134,In_4192);
xor U546 (N_546,In_4148,In_4638);
or U547 (N_547,In_3667,In_3670);
nor U548 (N_548,In_4234,In_661);
nand U549 (N_549,In_3514,In_3940);
nor U550 (N_550,In_3074,In_297);
or U551 (N_551,In_1737,In_1401);
xor U552 (N_552,In_4993,In_1912);
xnor U553 (N_553,In_4063,In_306);
xnor U554 (N_554,In_3009,In_690);
and U555 (N_555,In_182,In_2822);
nand U556 (N_556,In_4166,In_3147);
and U557 (N_557,In_4586,In_2496);
and U558 (N_558,In_3414,In_3759);
nor U559 (N_559,In_3313,In_4772);
nand U560 (N_560,In_684,In_293);
nor U561 (N_561,In_2329,In_2737);
or U562 (N_562,In_1406,In_1542);
nor U563 (N_563,In_3360,In_4604);
or U564 (N_564,In_74,In_3747);
and U565 (N_565,In_3751,In_443);
xor U566 (N_566,In_966,In_3021);
xnor U567 (N_567,In_3675,In_1780);
nand U568 (N_568,In_2140,In_4752);
nor U569 (N_569,In_2396,In_2950);
xor U570 (N_570,In_2570,In_4533);
and U571 (N_571,In_4737,In_426);
xnor U572 (N_572,In_2945,In_2733);
and U573 (N_573,In_3936,In_1047);
xor U574 (N_574,In_3739,In_4283);
nand U575 (N_575,In_1864,In_4620);
and U576 (N_576,In_3211,In_1148);
nand U577 (N_577,In_3710,In_2039);
nand U578 (N_578,In_4653,In_3804);
xnor U579 (N_579,In_4124,In_3905);
or U580 (N_580,In_41,In_3370);
xor U581 (N_581,In_4971,In_1670);
nand U582 (N_582,In_2053,In_4913);
nor U583 (N_583,In_647,In_1247);
nor U584 (N_584,In_4338,In_1945);
xor U585 (N_585,In_2207,In_1444);
nor U586 (N_586,In_3840,In_4838);
nand U587 (N_587,In_1067,In_1501);
or U588 (N_588,In_4313,In_225);
xor U589 (N_589,In_255,In_3551);
xnor U590 (N_590,In_1469,In_2044);
nor U591 (N_591,In_531,In_1855);
nor U592 (N_592,In_2299,In_347);
nand U593 (N_593,In_1572,In_2970);
xor U594 (N_594,In_2620,In_1849);
nor U595 (N_595,In_3301,In_1475);
and U596 (N_596,In_2336,In_3892);
or U597 (N_597,In_4931,In_4516);
and U598 (N_598,In_1312,In_4141);
nor U599 (N_599,In_3607,In_2863);
xnor U600 (N_600,In_4246,In_2186);
nor U601 (N_601,In_2348,In_1408);
nand U602 (N_602,In_461,In_798);
nand U603 (N_603,In_4982,In_4112);
or U604 (N_604,In_1831,In_2768);
and U605 (N_605,In_2658,In_549);
xor U606 (N_606,In_1083,In_3920);
nor U607 (N_607,In_1872,In_3761);
and U608 (N_608,In_1236,In_2215);
nand U609 (N_609,In_929,In_2901);
or U610 (N_610,In_3624,In_2602);
and U611 (N_611,In_2029,In_3395);
xnor U612 (N_612,In_1262,In_226);
or U613 (N_613,In_3929,In_1482);
xnor U614 (N_614,In_1473,In_1388);
nor U615 (N_615,In_2017,In_1715);
nand U616 (N_616,In_3530,In_1879);
and U617 (N_617,In_766,In_3999);
and U618 (N_618,In_3925,In_1643);
or U619 (N_619,In_261,In_2721);
nor U620 (N_620,In_2093,In_55);
and U621 (N_621,In_4750,In_2577);
xnor U622 (N_622,In_2625,In_3165);
and U623 (N_623,In_3027,In_3335);
or U624 (N_624,In_1661,In_2395);
and U625 (N_625,In_2529,In_384);
nand U626 (N_626,In_4231,In_435);
xnor U627 (N_627,In_4779,In_919);
and U628 (N_628,In_75,In_1077);
xnor U629 (N_629,In_3881,In_646);
or U630 (N_630,In_3682,In_1084);
xor U631 (N_631,In_3726,In_3993);
nor U632 (N_632,In_970,In_704);
or U633 (N_633,In_3471,In_2914);
and U634 (N_634,In_4116,In_2202);
or U635 (N_635,In_3939,In_1425);
and U636 (N_636,In_1563,In_1639);
nor U637 (N_637,In_968,In_2103);
xnor U638 (N_638,In_3058,In_4302);
xnor U639 (N_639,In_666,In_702);
xor U640 (N_640,In_1461,In_4142);
nor U641 (N_641,In_1131,In_2420);
or U642 (N_642,In_1431,In_2829);
or U643 (N_643,In_1324,In_3742);
nor U644 (N_644,In_1328,In_4798);
nor U645 (N_645,In_3679,In_3669);
nor U646 (N_646,In_4853,In_34);
and U647 (N_647,In_3937,In_368);
nand U648 (N_648,In_3871,In_2048);
or U649 (N_649,In_614,In_1005);
nand U650 (N_650,In_1378,In_2194);
nor U651 (N_651,In_893,In_3366);
xor U652 (N_652,In_4301,In_4934);
or U653 (N_653,In_4209,In_4658);
xnor U654 (N_654,In_4904,In_3523);
or U655 (N_655,In_1335,In_185);
or U656 (N_656,In_1224,In_3110);
nor U657 (N_657,In_40,In_4219);
nand U658 (N_658,In_2739,In_1180);
and U659 (N_659,In_4065,In_63);
or U660 (N_660,In_786,In_139);
nand U661 (N_661,In_4785,In_2378);
or U662 (N_662,In_668,In_3946);
xor U663 (N_663,In_1141,In_2851);
and U664 (N_664,In_1747,In_1713);
and U665 (N_665,In_3801,In_1800);
nand U666 (N_666,In_4895,In_2700);
and U667 (N_667,In_918,In_2233);
or U668 (N_668,In_2376,In_1897);
nand U669 (N_669,In_3433,In_340);
nor U670 (N_670,In_527,In_2806);
and U671 (N_671,In_3406,In_3332);
xnor U672 (N_672,In_4106,In_1241);
xor U673 (N_673,In_2714,In_2652);
nor U674 (N_674,In_223,In_2064);
nor U675 (N_675,In_258,In_2201);
and U676 (N_676,In_1574,In_1803);
xor U677 (N_677,In_2200,In_1387);
nor U678 (N_678,In_3697,In_625);
xnor U679 (N_679,In_3118,In_2387);
or U680 (N_680,In_816,In_1468);
nand U681 (N_681,In_4518,In_420);
xnor U682 (N_682,In_1751,In_1116);
xor U683 (N_683,In_337,In_4177);
xnor U684 (N_684,In_2655,In_3229);
and U685 (N_685,In_4617,In_3997);
nor U686 (N_686,In_1087,In_3286);
nand U687 (N_687,In_88,In_264);
and U688 (N_688,In_3621,In_3091);
or U689 (N_689,In_2169,In_4979);
nand U690 (N_690,In_1861,In_4855);
or U691 (N_691,In_3374,In_2574);
nand U692 (N_692,In_2813,In_586);
or U693 (N_693,In_2581,In_2717);
nor U694 (N_694,In_3639,In_2642);
xor U695 (N_695,In_4641,In_2047);
nor U696 (N_696,In_3671,In_410);
or U697 (N_697,In_4667,In_3318);
and U698 (N_698,In_3296,In_3271);
nand U699 (N_699,In_4213,In_1586);
and U700 (N_700,In_1858,In_814);
nand U701 (N_701,In_3882,In_3732);
or U702 (N_702,In_2380,In_4291);
xor U703 (N_703,In_2636,In_4114);
nand U704 (N_704,In_3499,In_2325);
or U705 (N_705,In_2887,In_457);
and U706 (N_706,In_1232,In_507);
nor U707 (N_707,In_2973,In_3596);
or U708 (N_708,In_1636,In_2562);
nand U709 (N_709,In_2785,In_234);
nand U710 (N_710,In_548,In_3762);
and U711 (N_711,In_4476,In_1839);
xnor U712 (N_712,In_2032,In_2171);
or U713 (N_713,In_4332,In_2723);
nor U714 (N_714,In_1002,In_153);
nand U715 (N_715,In_272,In_3288);
or U716 (N_716,In_1824,In_4428);
nand U717 (N_717,In_756,In_48);
xnor U718 (N_718,In_3212,In_2270);
xor U719 (N_719,In_1598,In_2255);
nand U720 (N_720,In_1189,In_1774);
nor U721 (N_721,In_4964,In_1429);
and U722 (N_722,In_4928,In_940);
nor U723 (N_723,In_2118,In_3351);
nor U724 (N_724,In_2531,In_4817);
and U725 (N_725,In_2273,In_2503);
nand U726 (N_726,In_2251,In_4613);
and U727 (N_727,In_1348,In_78);
or U728 (N_728,In_977,In_2137);
and U729 (N_729,In_3115,In_4060);
nand U730 (N_730,In_4702,In_2068);
nor U731 (N_731,In_3315,In_1905);
nor U732 (N_732,In_2454,In_2272);
and U733 (N_733,In_1013,In_2732);
and U734 (N_734,In_2965,In_4164);
xor U735 (N_735,In_2210,In_743);
or U736 (N_736,In_2228,In_3830);
nor U737 (N_737,In_1380,In_2461);
nor U738 (N_738,In_45,In_1108);
xnor U739 (N_739,In_2457,In_2178);
xor U740 (N_740,In_3298,In_1327);
or U741 (N_741,In_934,In_4097);
nand U742 (N_742,In_4296,In_2573);
xor U743 (N_743,In_502,In_1452);
or U744 (N_744,In_2234,In_3290);
xnor U745 (N_745,In_3319,In_3276);
nand U746 (N_746,In_269,In_3744);
and U747 (N_747,In_1010,In_2952);
and U748 (N_748,In_4431,In_3598);
and U749 (N_749,In_2479,In_2612);
or U750 (N_750,In_274,In_3548);
nand U751 (N_751,In_3468,In_2346);
nor U752 (N_752,In_4788,In_3934);
nor U753 (N_753,In_892,In_3292);
xnor U754 (N_754,In_2051,In_1544);
xnor U755 (N_755,In_3545,In_3431);
or U756 (N_756,In_4824,In_300);
nand U757 (N_757,In_4651,In_1835);
xnor U758 (N_758,In_4329,In_4172);
or U759 (N_759,In_2708,In_836);
and U760 (N_760,In_4580,In_467);
or U761 (N_761,In_4816,In_530);
and U762 (N_762,In_784,In_4886);
xor U763 (N_763,In_169,In_540);
and U764 (N_764,In_1873,In_4030);
xor U765 (N_765,In_3059,In_4976);
nand U766 (N_766,In_3572,In_3502);
nor U767 (N_767,In_3295,In_1808);
xor U768 (N_768,In_3856,In_4663);
xor U769 (N_769,In_3384,In_405);
xor U770 (N_770,In_289,In_3061);
and U771 (N_771,In_49,In_4901);
nand U772 (N_772,In_248,In_1918);
or U773 (N_773,In_4570,In_126);
xor U774 (N_774,In_888,In_4128);
and U775 (N_775,In_1205,In_795);
nand U776 (N_776,In_4378,In_809);
or U777 (N_777,In_4415,In_2643);
nor U778 (N_778,In_3386,In_969);
nand U779 (N_779,In_353,In_2141);
nand U780 (N_780,In_4692,In_105);
or U781 (N_781,In_141,In_2354);
nor U782 (N_782,In_3884,In_2925);
nor U783 (N_783,In_2159,In_3587);
nand U784 (N_784,In_3369,In_4015);
nand U785 (N_785,In_2995,In_4268);
nand U786 (N_786,In_667,In_2237);
xnor U787 (N_787,In_3878,In_2818);
or U788 (N_788,In_3978,In_1757);
and U789 (N_789,In_3969,In_515);
nand U790 (N_790,In_916,In_1681);
or U791 (N_791,In_567,In_194);
and U792 (N_792,In_2654,In_4318);
nor U793 (N_793,In_4940,In_4883);
nor U794 (N_794,In_1645,In_692);
or U795 (N_795,In_1732,In_3654);
or U796 (N_796,In_1679,In_3184);
nor U797 (N_797,In_3973,In_4893);
and U798 (N_798,In_164,In_4151);
xnor U799 (N_799,In_2892,In_972);
nand U800 (N_800,In_4085,In_1421);
xnor U801 (N_801,In_1260,In_1278);
xnor U802 (N_802,In_4673,In_2587);
and U803 (N_803,In_1703,In_547);
nor U804 (N_804,In_3033,In_4072);
or U805 (N_805,In_3348,In_939);
nor U806 (N_806,In_3394,In_3449);
nor U807 (N_807,In_2934,In_4791);
xor U808 (N_808,In_3200,In_4409);
xnor U809 (N_809,In_2670,In_2124);
nor U810 (N_810,In_3013,In_603);
xnor U811 (N_811,In_3914,In_3028);
and U812 (N_812,In_2583,In_2217);
and U813 (N_813,In_235,In_221);
or U814 (N_814,In_3122,In_596);
or U815 (N_815,In_4869,In_871);
or U816 (N_816,In_2070,In_1562);
nand U817 (N_817,In_1369,In_4573);
or U818 (N_818,In_921,In_3687);
nor U819 (N_819,In_897,In_4649);
or U820 (N_820,In_4054,In_629);
nand U821 (N_821,In_2182,In_4541);
or U822 (N_822,In_3007,In_1540);
xnor U823 (N_823,In_2165,In_2563);
and U824 (N_824,In_2223,In_4630);
or U825 (N_825,In_1825,In_2111);
nor U826 (N_826,In_2675,In_3746);
or U827 (N_827,In_806,In_3930);
xnor U828 (N_828,In_1073,In_4423);
or U829 (N_829,In_5,In_2028);
and U830 (N_830,In_835,In_304);
or U831 (N_831,In_1320,In_2742);
or U832 (N_832,In_4804,In_2424);
nand U833 (N_833,In_382,In_793);
and U834 (N_834,In_2435,In_503);
nand U835 (N_835,In_10,In_2580);
and U836 (N_836,In_1454,In_521);
and U837 (N_837,In_4851,In_3769);
and U838 (N_838,In_3988,In_2514);
nand U839 (N_839,In_315,In_1695);
nand U840 (N_840,In_3101,In_634);
and U841 (N_841,In_3540,In_752);
nand U842 (N_842,In_163,In_4242);
nand U843 (N_843,In_495,In_3300);
xnor U844 (N_844,In_4380,In_2679);
or U845 (N_845,In_2943,In_2116);
nor U846 (N_846,In_872,In_4384);
nand U847 (N_847,In_2958,In_4362);
nand U848 (N_848,In_208,In_3906);
or U849 (N_849,In_839,In_2951);
nor U850 (N_850,In_2645,In_1582);
or U851 (N_851,In_863,In_4288);
nor U852 (N_852,In_1607,In_3974);
nor U853 (N_853,In_2287,In_620);
nor U854 (N_854,In_316,In_2091);
xor U855 (N_855,In_2451,In_338);
xor U856 (N_856,In_2967,In_2246);
nand U857 (N_857,In_1534,In_377);
nand U858 (N_858,In_3547,In_1883);
nor U859 (N_859,In_4353,In_2584);
and U860 (N_860,In_3622,In_32);
nand U861 (N_861,In_3231,In_3510);
nand U862 (N_862,In_4832,In_4121);
nor U863 (N_863,In_1147,In_3259);
nor U864 (N_864,In_1826,In_3151);
xor U865 (N_865,In_2880,In_3968);
xor U866 (N_866,In_3217,In_4795);
and U867 (N_867,In_3003,In_2844);
nand U868 (N_868,In_3554,In_3333);
xnor U869 (N_869,In_4102,In_204);
or U870 (N_870,In_2002,In_1692);
nor U871 (N_871,In_195,In_2987);
nand U872 (N_872,In_3992,In_4696);
nor U873 (N_873,In_4032,In_3563);
nand U874 (N_874,In_3778,In_1273);
nand U875 (N_875,In_529,In_3809);
nand U876 (N_876,In_3784,In_165);
and U877 (N_877,In_4126,In_1443);
nor U878 (N_878,In_3851,In_3987);
and U879 (N_879,In_2979,In_3507);
nand U880 (N_880,In_1032,In_555);
and U881 (N_881,In_232,In_4023);
and U882 (N_882,In_2031,In_3020);
nand U883 (N_883,In_3176,In_3310);
nor U884 (N_884,In_3917,In_4810);
and U885 (N_885,In_1927,In_2550);
nand U886 (N_886,In_1908,In_249);
or U887 (N_887,In_2084,In_4616);
nand U888 (N_888,In_3304,In_1609);
or U889 (N_889,In_4163,In_1852);
xnor U890 (N_890,In_2497,In_4075);
or U891 (N_891,In_721,In_2793);
xnor U892 (N_892,In_845,In_2523);
or U893 (N_893,In_1280,In_4298);
nor U894 (N_894,In_1799,In_4467);
xnor U895 (N_895,In_385,In_2572);
nor U896 (N_896,In_4306,In_711);
and U897 (N_897,In_4807,In_997);
nor U898 (N_898,In_1075,In_3569);
nor U899 (N_899,In_3478,In_2781);
xnor U900 (N_900,In_4312,In_4311);
nor U901 (N_901,In_1819,In_2212);
nor U902 (N_902,In_359,In_2726);
nand U903 (N_903,In_598,In_2190);
or U904 (N_904,In_332,In_2552);
and U905 (N_905,In_4127,In_2904);
nand U906 (N_906,In_3872,In_3236);
or U907 (N_907,In_4778,In_2619);
and U908 (N_908,In_4640,In_4402);
nor U909 (N_909,In_2521,In_2983);
nor U910 (N_910,In_2016,In_2369);
nand U911 (N_911,In_1249,In_4418);
or U912 (N_912,In_1954,In_509);
or U913 (N_913,In_2756,In_15);
and U914 (N_914,In_2639,In_4361);
nor U915 (N_915,In_2176,In_3344);
and U916 (N_916,In_3114,In_4668);
nor U917 (N_917,In_83,In_1374);
and U918 (N_918,In_4507,In_882);
or U919 (N_919,In_2604,In_1126);
nand U920 (N_920,In_295,In_1637);
and U921 (N_921,In_3131,In_3811);
xnor U922 (N_922,In_3121,In_821);
and U923 (N_923,In_626,In_3401);
nor U924 (N_924,In_1924,In_656);
or U925 (N_925,In_1530,In_2400);
xnor U926 (N_926,In_3473,In_751);
nor U927 (N_927,In_1659,In_290);
and U928 (N_928,In_3991,In_2928);
nand U929 (N_929,In_4365,In_4215);
and U930 (N_930,In_4871,In_4191);
and U931 (N_931,In_3901,In_146);
xor U932 (N_932,In_1729,In_902);
or U933 (N_933,In_2443,In_1445);
xnor U934 (N_934,In_4342,In_4315);
xor U935 (N_935,In_3869,In_587);
nor U936 (N_936,In_3270,In_2540);
xor U937 (N_937,In_1199,In_2682);
nand U938 (N_938,In_979,In_1538);
xnor U939 (N_939,In_943,In_27);
xor U940 (N_940,In_492,In_361);
nor U941 (N_941,In_1311,In_4852);
nand U942 (N_942,In_2452,In_2908);
or U943 (N_943,In_4953,In_4147);
and U944 (N_944,In_2069,In_873);
xnor U945 (N_945,In_4890,In_3144);
or U946 (N_946,In_2794,In_2314);
or U947 (N_947,In_1467,In_709);
xor U948 (N_948,In_4591,In_1251);
xor U949 (N_949,In_1936,In_4879);
and U950 (N_950,In_1915,In_1049);
nand U951 (N_951,In_2765,In_429);
xnor U952 (N_952,In_4173,In_1722);
xnor U953 (N_953,In_4556,In_3501);
nor U954 (N_954,In_4900,In_1874);
nor U955 (N_955,In_1931,In_506);
or U956 (N_956,In_995,In_4777);
nand U957 (N_957,In_2705,In_4634);
nand U958 (N_958,In_2192,In_464);
or U959 (N_959,In_2716,In_2890);
and U960 (N_960,In_4744,In_524);
nand U961 (N_961,In_378,In_764);
xor U962 (N_962,In_4885,In_1152);
or U963 (N_963,In_3149,In_2027);
xnor U964 (N_964,In_4150,In_3891);
xnor U965 (N_965,In_4607,In_2160);
and U966 (N_966,In_3496,In_728);
nand U967 (N_967,In_1284,In_3459);
nor U968 (N_968,In_2633,In_818);
and U969 (N_969,In_1739,In_4140);
and U970 (N_970,In_4305,In_345);
nor U971 (N_971,In_1003,In_369);
xor U972 (N_972,In_4686,In_2784);
or U973 (N_973,In_4605,In_3760);
xnor U974 (N_974,In_3592,In_4441);
nor U975 (N_975,In_2412,In_960);
nor U976 (N_976,In_4180,In_2894);
nand U977 (N_977,In_3538,In_4773);
nor U978 (N_978,In_828,In_3466);
or U979 (N_979,In_4289,In_29);
or U980 (N_980,In_4100,In_3986);
nor U981 (N_981,In_1662,In_1511);
nor U982 (N_982,In_1476,In_3467);
xor U983 (N_983,In_2467,In_2506);
nor U984 (N_984,In_731,In_4951);
xnor U985 (N_985,In_2290,In_4740);
and U986 (N_986,In_391,In_4359);
and U987 (N_987,In_2795,In_662);
nand U988 (N_988,In_3367,In_3183);
or U989 (N_989,In_2809,In_113);
nor U990 (N_990,In_4326,In_860);
nand U991 (N_991,In_3633,In_1520);
and U992 (N_992,In_572,In_4492);
nand U993 (N_993,In_575,In_982);
nor U994 (N_994,In_1923,In_4292);
xor U995 (N_995,In_637,In_4264);
nor U996 (N_996,In_4115,In_1647);
nand U997 (N_997,In_3078,In_4373);
xor U998 (N_998,In_1580,In_4098);
xnor U999 (N_999,In_1653,In_3132);
xor U1000 (N_1000,In_3376,In_3935);
nor U1001 (N_1001,In_3314,In_4002);
nand U1002 (N_1002,In_176,In_1550);
xor U1003 (N_1003,In_4927,In_2447);
and U1004 (N_1004,In_849,In_3247);
xor U1005 (N_1005,In_4372,In_2304);
xnor U1006 (N_1006,In_4035,In_4120);
xnor U1007 (N_1007,In_4412,In_2691);
or U1008 (N_1008,In_4972,In_3642);
nand U1009 (N_1009,In_3866,In_2668);
nand U1010 (N_1010,In_3015,In_178);
nor U1011 (N_1011,In_1308,In_3197);
and U1012 (N_1012,In_1666,In_3043);
nor U1013 (N_1013,In_1581,In_645);
nor U1014 (N_1014,In_469,In_3045);
nor U1015 (N_1015,In_4043,In_2500);
xnor U1016 (N_1016,In_2003,In_3609);
xor U1017 (N_1017,In_2269,In_2279);
xor U1018 (N_1018,In_4780,In_180);
and U1019 (N_1019,In_4189,In_2013);
or U1020 (N_1020,In_3665,In_2334);
nor U1021 (N_1021,In_1419,In_3646);
or U1022 (N_1022,In_3133,In_716);
or U1023 (N_1023,In_211,In_3214);
or U1024 (N_1024,In_1410,In_3724);
nor U1025 (N_1025,In_1875,In_3752);
xnor U1026 (N_1026,In_2980,In_129);
nor U1027 (N_1027,In_1853,In_1307);
and U1028 (N_1028,In_1603,In_4675);
or U1029 (N_1029,In_2113,In_1956);
and U1030 (N_1030,In_2096,In_4991);
nand U1031 (N_1031,In_2360,In_4153);
xor U1032 (N_1032,In_481,In_3415);
xor U1033 (N_1033,In_4588,In_3857);
or U1034 (N_1034,In_4019,In_4483);
xor U1035 (N_1035,In_3379,In_4759);
or U1036 (N_1036,In_4376,In_992);
xnor U1037 (N_1037,In_2197,In_1769);
or U1038 (N_1038,In_2450,In_4392);
and U1039 (N_1039,In_4276,In_254);
nand U1040 (N_1040,In_1935,In_2164);
nor U1041 (N_1041,In_4265,In_1877);
or U1042 (N_1042,In_582,In_974);
nand U1043 (N_1043,In_4408,In_2488);
or U1044 (N_1044,In_1656,In_358);
xnor U1045 (N_1045,In_2015,In_4677);
nand U1046 (N_1046,In_993,In_508);
xnor U1047 (N_1047,In_93,In_1480);
nor U1048 (N_1048,In_998,In_585);
nor U1049 (N_1049,In_1282,In_2133);
xnor U1050 (N_1050,In_1039,In_539);
or U1051 (N_1051,In_4790,In_2754);
and U1052 (N_1052,In_2446,In_3755);
nand U1053 (N_1053,In_3416,In_2060);
and U1054 (N_1054,In_1685,In_4160);
xor U1055 (N_1055,In_2998,In_739);
nand U1056 (N_1056,In_3166,In_4854);
nor U1057 (N_1057,In_638,In_4626);
and U1058 (N_1058,In_3096,In_3887);
or U1059 (N_1059,In_2606,In_733);
nand U1060 (N_1060,In_3303,In_1929);
nor U1061 (N_1061,In_4200,In_1037);
or U1062 (N_1062,In_4394,In_1361);
and U1063 (N_1063,In_2179,In_4749);
and U1064 (N_1064,In_1673,In_1519);
xor U1065 (N_1065,In_4847,In_2240);
nand U1066 (N_1066,In_1377,In_760);
xnor U1067 (N_1067,In_714,In_1059);
nand U1068 (N_1068,In_544,In_2532);
nor U1069 (N_1069,In_2333,In_777);
nand U1070 (N_1070,In_76,In_4092);
and U1071 (N_1071,In_1198,In_1625);
nand U1072 (N_1072,In_778,In_3264);
and U1073 (N_1073,In_2770,In_486);
xnor U1074 (N_1074,In_3385,In_1516);
xnor U1075 (N_1075,In_3275,In_4135);
nor U1076 (N_1076,In_4453,In_1350);
nand U1077 (N_1077,In_3837,In_1587);
xnor U1078 (N_1078,In_4107,In_2637);
xnor U1079 (N_1079,In_3630,In_2236);
nor U1080 (N_1080,In_3757,In_4566);
and U1081 (N_1081,In_1863,In_1043);
or U1082 (N_1082,In_1358,In_3674);
and U1083 (N_1083,In_1031,In_494);
xor U1084 (N_1084,In_788,In_2960);
xor U1085 (N_1085,In_376,In_3338);
and U1086 (N_1086,In_551,In_472);
or U1087 (N_1087,In_2187,In_1368);
xor U1088 (N_1088,In_4202,In_2905);
nand U1089 (N_1089,In_844,In_686);
and U1090 (N_1090,In_2440,In_4513);
and U1091 (N_1091,In_2071,In_4666);
nand U1092 (N_1092,In_4959,In_4611);
nand U1093 (N_1093,In_3916,In_2544);
xnor U1094 (N_1094,In_2504,In_4468);
or U1095 (N_1095,In_1462,In_2431);
or U1096 (N_1096,In_758,In_4307);
nand U1097 (N_1097,In_1294,In_2696);
nand U1098 (N_1098,In_2814,In_4424);
and U1099 (N_1099,In_1940,In_2632);
or U1100 (N_1100,In_4581,In_3023);
or U1101 (N_1101,In_4517,In_2820);
xnor U1102 (N_1102,In_474,In_1314);
xnor U1103 (N_1103,In_3686,In_3170);
xor U1104 (N_1104,In_3626,In_3267);
or U1105 (N_1105,In_4530,In_4949);
xor U1106 (N_1106,In_4806,In_1492);
and U1107 (N_1107,In_2154,In_59);
nand U1108 (N_1108,In_437,In_1109);
nand U1109 (N_1109,In_351,In_4528);
nor U1110 (N_1110,In_1814,In_19);
nand U1111 (N_1111,In_1268,In_3943);
nand U1112 (N_1112,In_3527,In_1301);
xnor U1113 (N_1113,In_4055,In_1056);
nor U1114 (N_1114,In_2484,In_1630);
nand U1115 (N_1115,In_450,In_2989);
or U1116 (N_1116,In_12,In_560);
xor U1117 (N_1117,In_2472,In_3975);
nand U1118 (N_1118,In_2624,In_4590);
and U1119 (N_1119,In_3336,In_1736);
and U1120 (N_1120,In_846,In_891);
nand U1121 (N_1121,In_106,In_4007);
xnor U1122 (N_1122,In_3452,In_2249);
and U1123 (N_1123,In_3436,In_3439);
or U1124 (N_1124,In_3272,In_3001);
or U1125 (N_1125,In_4628,In_4357);
or U1126 (N_1126,In_2441,In_3143);
nand U1127 (N_1127,In_374,In_1289);
nand U1128 (N_1128,In_2138,In_3464);
nor U1129 (N_1129,In_1370,In_1628);
or U1130 (N_1130,In_1237,In_1626);
nand U1131 (N_1131,In_2808,In_914);
nor U1132 (N_1132,In_3539,In_2122);
xnor U1133 (N_1133,In_1743,In_4910);
or U1134 (N_1134,In_3694,In_142);
nand U1135 (N_1135,In_201,In_700);
nor U1136 (N_1136,In_1514,In_1053);
and U1137 (N_1137,In_4665,In_3823);
nor U1138 (N_1138,In_448,In_3191);
and U1139 (N_1139,In_4058,In_1446);
xor U1140 (N_1140,In_1395,In_4073);
or U1141 (N_1141,In_4170,In_3324);
nor U1142 (N_1142,In_2586,In_1265);
and U1143 (N_1143,In_563,In_3727);
or U1144 (N_1144,In_4873,In_1057);
nand U1145 (N_1145,In_1407,In_2492);
xor U1146 (N_1146,In_2684,In_949);
nor U1147 (N_1147,In_112,In_2662);
nand U1148 (N_1148,In_4912,In_3794);
nor U1149 (N_1149,In_2635,In_2486);
nand U1150 (N_1150,In_266,In_2107);
xnor U1151 (N_1151,In_2898,In_4508);
nor U1152 (N_1152,In_453,In_4633);
nand U1153 (N_1153,In_2789,In_1965);
or U1154 (N_1154,In_4815,In_1869);
xnor U1155 (N_1155,In_3494,In_1195);
and U1156 (N_1156,In_4320,In_2198);
and U1157 (N_1157,In_1991,In_1993);
nand U1158 (N_1158,In_669,In_1913);
nand U1159 (N_1159,In_1512,In_1221);
or U1160 (N_1160,In_2067,In_4917);
or U1161 (N_1161,In_2056,In_4818);
or U1162 (N_1162,In_3094,In_785);
or U1163 (N_1163,In_3254,In_1420);
or U1164 (N_1164,In_2886,In_3079);
nand U1165 (N_1165,In_323,In_4198);
nand U1166 (N_1166,In_3543,In_4096);
nand U1167 (N_1167,In_901,In_2972);
xnor U1168 (N_1168,In_1999,In_2507);
nor U1169 (N_1169,In_2997,In_811);
or U1170 (N_1170,In_1317,In_2403);
or U1171 (N_1171,In_4317,In_3570);
nor U1172 (N_1172,In_4230,In_4026);
and U1173 (N_1173,In_313,In_2466);
or U1174 (N_1174,In_2324,In_2356);
nor U1175 (N_1175,In_4078,In_3961);
xnor U1176 (N_1176,In_1381,In_1818);
or U1177 (N_1177,In_2505,In_2300);
and U1178 (N_1178,In_2139,In_3838);
nand U1179 (N_1179,In_1841,In_2906);
nand U1180 (N_1180,In_879,In_1450);
nor U1181 (N_1181,In_1992,In_1837);
nor U1182 (N_1182,In_2033,In_1677);
and U1183 (N_1183,In_183,In_107);
and U1184 (N_1184,In_84,In_2285);
nand U1185 (N_1185,In_4878,In_2576);
and U1186 (N_1186,In_184,In_605);
nand U1187 (N_1187,In_2166,In_3599);
or U1188 (N_1188,In_4053,In_4419);
xnor U1189 (N_1189,In_770,In_4571);
and U1190 (N_1190,In_3741,In_2163);
nor U1191 (N_1191,In_3256,In_1717);
nor U1192 (N_1192,In_1998,In_4717);
xor U1193 (N_1193,In_2340,In_3268);
or U1194 (N_1194,In_4117,In_2527);
or U1195 (N_1195,In_885,In_3263);
or U1196 (N_1196,In_298,In_3262);
nor U1197 (N_1197,In_1418,In_4358);
xor U1198 (N_1198,In_1202,In_3308);
nand U1199 (N_1199,In_1438,In_1);
xor U1200 (N_1200,In_2476,In_2783);
or U1201 (N_1201,In_303,In_4050);
xor U1202 (N_1202,In_1714,In_4796);
or U1203 (N_1203,In_2597,In_3942);
nand U1204 (N_1204,In_3112,In_3164);
nand U1205 (N_1205,In_1953,In_4545);
nor U1206 (N_1206,In_3522,In_4645);
or U1207 (N_1207,In_2957,In_1845);
and U1208 (N_1208,In_3442,In_1515);
nor U1209 (N_1209,In_514,In_773);
and U1210 (N_1210,In_4430,In_3080);
nand U1211 (N_1211,In_3647,In_2358);
xnor U1212 (N_1212,In_2153,In_2579);
xnor U1213 (N_1213,In_1428,In_2433);
or U1214 (N_1214,In_4600,In_2386);
and U1215 (N_1215,In_4352,In_2713);
or U1216 (N_1216,In_3047,In_4095);
xnor U1217 (N_1217,In_155,In_4475);
nor U1218 (N_1218,In_1784,In_4656);
nor U1219 (N_1219,In_4082,In_1211);
nand U1220 (N_1220,In_4685,In_4436);
xnor U1221 (N_1221,In_2697,In_1033);
nand U1222 (N_1222,In_1218,In_1577);
nor U1223 (N_1223,In_1871,In_1876);
and U1224 (N_1224,In_2203,In_287);
and U1225 (N_1225,In_4887,In_1518);
or U1226 (N_1226,In_2977,In_4225);
or U1227 (N_1227,In_3618,In_4322);
nand U1228 (N_1228,In_2767,In_1186);
nor U1229 (N_1229,In_1699,In_750);
and U1230 (N_1230,In_1192,In_3451);
and U1231 (N_1231,In_94,In_1807);
or U1232 (N_1232,In_271,In_1372);
and U1233 (N_1233,In_947,In_3053);
or U1234 (N_1234,In_4245,In_395);
or U1235 (N_1235,In_490,In_1227);
nor U1236 (N_1236,In_4355,In_1276);
or U1237 (N_1237,In_3948,In_2812);
and U1238 (N_1238,In_1154,In_1566);
nand U1239 (N_1239,In_4042,In_4472);
xnor U1240 (N_1240,In_4377,In_3567);
nor U1241 (N_1241,In_4712,In_898);
and U1242 (N_1242,In_3994,In_2881);
xnor U1243 (N_1243,In_2537,In_1177);
xor U1244 (N_1244,In_1173,In_4194);
nand U1245 (N_1245,In_3328,In_4401);
nand U1246 (N_1246,In_3695,In_2748);
and U1247 (N_1247,In_4367,In_1015);
xnor U1248 (N_1248,In_3075,In_3064);
or U1249 (N_1249,In_2078,In_4621);
nand U1250 (N_1250,In_1235,In_1222);
nor U1251 (N_1251,In_3798,In_431);
or U1252 (N_1252,In_314,In_4478);
or U1253 (N_1253,In_2805,In_2752);
and U1254 (N_1254,In_2130,In_1507);
or U1255 (N_1255,In_318,In_3870);
nand U1256 (N_1256,In_4186,In_4783);
nand U1257 (N_1257,In_1719,In_3162);
or U1258 (N_1258,In_4719,In_2508);
or U1259 (N_1259,In_2623,In_333);
xor U1260 (N_1260,In_1220,In_877);
xor U1261 (N_1261,In_4733,In_2465);
xnor U1262 (N_1262,In_1706,In_4646);
nand U1263 (N_1263,In_2605,In_2185);
nor U1264 (N_1264,In_2375,In_449);
or U1265 (N_1265,In_4837,In_1102);
nor U1266 (N_1266,In_933,In_983);
nor U1267 (N_1267,In_3055,In_3457);
or U1268 (N_1268,In_1684,In_2729);
and U1269 (N_1269,In_4849,In_4723);
or U1270 (N_1270,In_2244,In_4088);
or U1271 (N_1271,In_4786,In_4676);
and U1272 (N_1272,In_1340,In_4625);
or U1273 (N_1273,In_4860,In_476);
nor U1274 (N_1274,In_39,In_62);
and U1275 (N_1275,In_1110,In_1740);
and U1276 (N_1276,In_511,In_1921);
nor U1277 (N_1277,In_2510,In_3952);
xnor U1278 (N_1278,In_4228,In_3849);
nor U1279 (N_1279,In_430,In_1551);
nand U1280 (N_1280,In_3171,In_4829);
nor U1281 (N_1281,In_4877,In_407);
xor U1282 (N_1282,In_3603,In_4263);
nor U1283 (N_1283,In_0,In_612);
xor U1284 (N_1284,In_4700,In_440);
xnor U1285 (N_1285,In_4279,In_3409);
or U1286 (N_1286,In_2341,In_238);
xnor U1287 (N_1287,In_1231,In_2564);
xnor U1288 (N_1288,In_1257,In_4489);
nand U1289 (N_1289,In_1342,In_3102);
xor U1290 (N_1290,In_2811,In_390);
and U1291 (N_1291,In_1174,In_4340);
or U1292 (N_1292,In_889,In_810);
and U1293 (N_1293,In_3465,In_3576);
xnor U1294 (N_1294,In_37,In_2241);
or U1295 (N_1295,In_4937,In_1878);
nand U1296 (N_1296,In_1365,In_1848);
and U1297 (N_1297,In_3038,In_3776);
nand U1298 (N_1298,In_1763,In_2749);
xor U1299 (N_1299,In_4029,In_4575);
and U1300 (N_1300,In_198,In_2699);
or U1301 (N_1301,In_4303,In_1071);
or U1302 (N_1302,In_2710,In_3895);
and U1303 (N_1303,In_4360,In_3795);
and U1304 (N_1304,In_1632,In_1310);
and U1305 (N_1305,In_584,In_4028);
and U1306 (N_1306,In_1014,In_4766);
nor U1307 (N_1307,In_2853,In_1076);
or U1308 (N_1308,In_2640,In_583);
or U1309 (N_1309,In_2430,In_1453);
and U1310 (N_1310,In_1157,In_1354);
and U1311 (N_1311,In_4233,In_1034);
xor U1312 (N_1312,In_4277,In_23);
or U1313 (N_1313,In_3979,In_3299);
nand U1314 (N_1314,In_2309,In_3443);
and U1315 (N_1315,In_1620,In_3788);
or U1316 (N_1316,In_4444,In_2685);
nand U1317 (N_1317,In_4935,In_988);
and U1318 (N_1318,In_965,In_6);
nor U1319 (N_1319,In_4083,In_3632);
nor U1320 (N_1320,In_3643,In_2553);
and U1321 (N_1321,In_387,In_1982);
or U1322 (N_1322,In_3796,In_170);
nor U1323 (N_1323,In_2966,In_1964);
xor U1324 (N_1324,In_1436,In_4764);
nand U1325 (N_1325,In_3339,In_4615);
xor U1326 (N_1326,In_2941,In_1590);
nor U1327 (N_1327,In_3029,In_4335);
and U1328 (N_1328,In_1955,In_30);
or U1329 (N_1329,In_2771,In_1288);
nor U1330 (N_1330,In_3041,In_1744);
or U1331 (N_1331,In_2557,In_4801);
xnor U1332 (N_1332,In_4587,In_535);
or U1333 (N_1333,In_4187,In_813);
and U1334 (N_1334,In_4076,In_4902);
and U1335 (N_1335,In_46,In_3590);
and U1336 (N_1336,In_1817,In_1061);
nor U1337 (N_1337,In_3274,In_2816);
and U1338 (N_1338,In_2933,In_1795);
xnor U1339 (N_1339,In_1122,In_36);
and U1340 (N_1340,In_1069,In_2459);
nor U1341 (N_1341,In_763,In_4091);
xnor U1342 (N_1342,In_942,In_3412);
xor U1343 (N_1343,In_3518,In_135);
nor U1344 (N_1344,In_4179,In_3497);
or U1345 (N_1345,In_2427,In_2397);
xor U1346 (N_1346,In_421,In_3026);
nand U1347 (N_1347,In_2054,In_1124);
nor U1348 (N_1348,In_1752,In_1491);
and U1349 (N_1349,In_3396,In_4709);
or U1350 (N_1350,In_1465,In_4542);
or U1351 (N_1351,In_2526,In_3446);
and U1352 (N_1352,In_1134,In_3039);
and U1353 (N_1353,In_4232,In_1820);
nor U1354 (N_1354,In_4207,In_4235);
nor U1355 (N_1355,In_1095,In_3034);
xor U1356 (N_1356,In_4872,In_3818);
nand U1357 (N_1357,In_4784,In_782);
or U1358 (N_1358,In_1894,In_2688);
nor U1359 (N_1359,In_1081,In_3410);
xnor U1360 (N_1360,In_3985,In_2148);
nor U1361 (N_1361,In_1570,In_3155);
xor U1362 (N_1362,In_3054,In_2384);
nor U1363 (N_1363,In_4932,In_2247);
and U1364 (N_1364,In_2988,In_569);
xor U1365 (N_1365,In_352,In_3951);
xor U1366 (N_1366,In_2867,In_425);
nand U1367 (N_1367,In_1593,In_525);
and U1368 (N_1368,In_3325,In_2843);
xnor U1369 (N_1369,In_1764,In_2897);
and U1370 (N_1370,In_4559,In_4950);
or U1371 (N_1371,In_2516,In_3894);
and U1372 (N_1372,In_951,In_3454);
xor U1373 (N_1373,In_4867,In_2275);
nor U1374 (N_1374,In_2289,In_4118);
nand U1375 (N_1375,In_2,In_1911);
xor U1376 (N_1376,In_3103,In_1376);
nor U1377 (N_1377,In_2831,In_3287);
nor U1378 (N_1378,In_688,In_2940);
xnor U1379 (N_1379,In_1027,In_246);
nor U1380 (N_1380,In_3285,In_4999);
or U1381 (N_1381,In_2899,In_2893);
and U1382 (N_1382,In_2037,In_641);
and U1383 (N_1383,In_4880,In_922);
or U1384 (N_1384,In_542,In_3863);
or U1385 (N_1385,In_2319,In_3606);
or U1386 (N_1386,In_3195,In_4655);
nor U1387 (N_1387,In_3550,In_3330);
xnor U1388 (N_1388,In_2779,In_580);
nand U1389 (N_1389,In_4256,In_4351);
nor U1390 (N_1390,In_1128,In_1724);
xnor U1391 (N_1391,In_327,In_2079);
and U1392 (N_1392,In_4555,In_127);
nand U1393 (N_1393,In_4730,In_2707);
nor U1394 (N_1394,In_1346,In_4282);
nor U1395 (N_1395,In_1127,In_2157);
nor U1396 (N_1396,In_3279,In_2836);
nand U1397 (N_1397,In_3711,In_1164);
and U1398 (N_1398,In_1880,In_219);
and U1399 (N_1399,In_4363,In_2773);
and U1400 (N_1400,In_268,In_56);
nand U1401 (N_1401,In_3354,In_4500);
or U1402 (N_1402,In_1529,In_3014);
xor U1403 (N_1403,In_1442,In_148);
and U1404 (N_1404,In_2439,In_1721);
nor U1405 (N_1405,In_4965,In_4511);
nand U1406 (N_1406,In_2363,In_3915);
or U1407 (N_1407,In_4514,In_3799);
and U1408 (N_1408,In_4036,In_1146);
xnor U1409 (N_1409,In_1163,In_4447);
nand U1410 (N_1410,In_2764,In_3938);
nor U1411 (N_1411,In_3828,In_2525);
and U1412 (N_1412,In_466,In_4720);
nor U1413 (N_1413,In_4523,In_366);
or U1414 (N_1414,In_1440,In_4385);
nand U1415 (N_1415,In_2931,In_1263);
xor U1416 (N_1416,In_2810,In_3709);
xor U1417 (N_1417,In_1213,In_2885);
xor U1418 (N_1418,In_827,In_4149);
or U1419 (N_1419,In_3006,In_4558);
or U1420 (N_1420,In_2902,In_227);
and U1421 (N_1421,In_1718,In_4698);
and U1422 (N_1422,In_3476,In_1571);
and U1423 (N_1423,In_2243,In_471);
nor U1424 (N_1424,In_4398,In_2990);
xnor U1425 (N_1425,In_4158,In_3854);
or U1426 (N_1426,In_1063,In_252);
xnor U1427 (N_1427,In_3134,In_1343);
nand U1428 (N_1428,In_2024,In_2038);
and U1429 (N_1429,In_3729,In_4494);
or U1430 (N_1430,In_3971,In_1503);
or U1431 (N_1431,In_4753,In_3153);
nor U1432 (N_1432,In_4295,In_4978);
or U1433 (N_1433,In_1866,In_4321);
and U1434 (N_1434,In_335,In_3676);
or U1435 (N_1435,In_3743,In_4347);
xnor U1436 (N_1436,In_2522,In_3160);
or U1437 (N_1437,In_2423,In_1296);
nand U1438 (N_1438,In_2193,In_762);
nand U1439 (N_1439,In_1860,In_1315);
nor U1440 (N_1440,In_589,In_3931);
nand U1441 (N_1441,In_3612,In_1156);
nand U1442 (N_1442,In_487,In_732);
nor U1443 (N_1443,In_1483,In_3740);
xor U1444 (N_1444,In_4457,In_3283);
nor U1445 (N_1445,In_2115,In_2283);
nand U1446 (N_1446,In_4205,In_3331);
nor U1447 (N_1447,In_1890,In_3273);
or U1448 (N_1448,In_4501,In_2477);
xor U1449 (N_1449,In_591,In_931);
or U1450 (N_1450,In_952,In_3786);
xor U1451 (N_1451,In_4726,In_1975);
nand U1452 (N_1452,In_987,In_2174);
xnor U1453 (N_1453,In_4348,In_927);
nand U1454 (N_1454,In_4397,In_4495);
xor U1455 (N_1455,In_3371,In_2949);
xor U1456 (N_1456,In_1028,In_1029);
or U1457 (N_1457,In_4520,In_2189);
nand U1458 (N_1458,In_2725,In_3350);
or U1459 (N_1459,In_907,In_3685);
nor U1460 (N_1460,In_2254,In_101);
nand U1461 (N_1461,In_2368,In_1528);
and U1462 (N_1462,In_354,In_3441);
nor U1463 (N_1463,In_3728,In_2561);
xor U1464 (N_1464,In_1667,In_4938);
xor U1465 (N_1465,In_652,In_832);
nand U1466 (N_1466,In_2578,In_3042);
nor U1467 (N_1467,In_3924,In_615);
xor U1468 (N_1468,In_3958,In_3883);
nand U1469 (N_1469,In_2948,In_71);
nor U1470 (N_1470,In_576,In_2993);
nand U1471 (N_1471,In_1171,In_2498);
xor U1472 (N_1472,In_3470,In_1504);
nor U1473 (N_1473,In_328,In_3867);
or U1474 (N_1474,In_2209,In_3861);
nor U1475 (N_1475,In_1810,In_2297);
xnor U1476 (N_1476,In_3241,In_4066);
or U1477 (N_1477,In_4374,In_3779);
or U1478 (N_1478,In_910,In_1135);
nor U1479 (N_1479,In_1054,In_4382);
or U1480 (N_1480,In_719,In_749);
and U1481 (N_1481,In_2536,In_3062);
nor U1482 (N_1482,In_2542,In_3593);
or U1483 (N_1483,In_1606,In_2592);
or U1484 (N_1484,In_4056,In_2517);
nor U1485 (N_1485,In_4211,In_2058);
nand U1486 (N_1486,In_1549,In_152);
and U1487 (N_1487,In_1634,In_4936);
nor U1488 (N_1488,In_1776,In_1834);
nand U1489 (N_1489,In_1787,In_3346);
and U1490 (N_1490,In_3498,In_2008);
and U1491 (N_1491,In_3577,In_1971);
nor U1492 (N_1492,In_4863,In_1691);
nor U1493 (N_1493,In_671,In_736);
and U1494 (N_1494,In_1264,In_4413);
and U1495 (N_1495,In_1101,In_1300);
nand U1496 (N_1496,In_210,In_2291);
and U1497 (N_1497,In_3719,In_2622);
nor U1498 (N_1498,In_2792,In_2147);
nand U1499 (N_1499,In_3555,In_1093);
xnor U1500 (N_1500,In_2753,In_1456);
nand U1501 (N_1501,In_1008,In_1234);
nor U1502 (N_1502,In_4195,In_2534);
and U1503 (N_1503,In_1142,In_2511);
nand U1504 (N_1504,In_3579,In_3575);
xnor U1505 (N_1505,In_1770,In_4527);
nand U1506 (N_1506,In_2286,In_1618);
xnor U1507 (N_1507,In_1916,In_1417);
xor U1508 (N_1508,In_3398,In_1760);
xnor U1509 (N_1509,In_2493,In_3148);
xnor U1510 (N_1510,In_1682,In_2364);
or U1511 (N_1511,In_3753,In_1248);
nor U1512 (N_1512,In_2357,In_735);
nand U1513 (N_1513,In_1865,In_857);
or U1514 (N_1514,In_4619,In_1413);
and U1515 (N_1515,In_3359,In_1394);
and U1516 (N_1516,In_1333,In_1206);
nand U1517 (N_1517,In_4090,In_2335);
or U1518 (N_1518,In_4123,In_1944);
xnor U1519 (N_1519,In_3037,In_613);
or U1520 (N_1520,In_3095,In_566);
nand U1521 (N_1521,In_4497,In_2282);
and U1522 (N_1522,In_2857,In_2672);
and U1523 (N_1523,In_2755,In_4995);
or U1524 (N_1524,In_2545,In_67);
and U1525 (N_1525,In_2180,In_2919);
nor U1526 (N_1526,In_4671,In_3839);
nand U1527 (N_1527,In_880,In_4241);
nand U1528 (N_1528,In_346,In_2175);
nor U1529 (N_1529,In_1026,In_119);
or U1530 (N_1530,In_1830,In_2010);
nor U1531 (N_1531,In_2337,In_1983);
nor U1532 (N_1532,In_1966,In_2519);
nor U1533 (N_1533,In_562,In_3472);
nor U1534 (N_1534,In_1385,In_932);
and U1535 (N_1535,In_3750,In_3956);
nand U1536 (N_1536,In_501,In_3610);
and U1537 (N_1537,In_499,In_1292);
xnor U1538 (N_1538,In_2788,In_1663);
xor U1539 (N_1539,In_3280,In_9);
nand U1540 (N_1540,In_3219,In_4755);
or U1541 (N_1541,In_2869,In_768);
nor U1542 (N_1542,In_4477,In_950);
and U1543 (N_1543,In_3699,In_3178);
and U1544 (N_1544,In_4802,In_3556);
xnor U1545 (N_1545,In_3010,In_3516);
or U1546 (N_1546,In_676,In_4918);
xor U1547 (N_1547,In_151,In_279);
and U1548 (N_1548,In_3040,In_394);
nand U1549 (N_1549,In_2235,In_1497);
nor U1550 (N_1550,In_1427,In_3432);
xnor U1551 (N_1551,In_2501,In_717);
and U1552 (N_1552,In_747,In_2173);
or U1553 (N_1553,In_3745,In_4583);
nand U1554 (N_1554,In_3337,In_1040);
nor U1555 (N_1555,In_1228,In_4446);
and U1556 (N_1556,In_2274,In_200);
nor U1557 (N_1557,In_3611,In_1403);
or U1558 (N_1558,In_3771,In_4825);
and U1559 (N_1559,In_2338,In_2930);
or U1560 (N_1560,In_237,In_4945);
nand U1561 (N_1561,In_1804,In_653);
or U1562 (N_1562,In_2746,In_4369);
xor U1563 (N_1563,In_4943,In_1161);
xor U1564 (N_1564,In_61,In_1384);
or U1565 (N_1565,In_124,In_4261);
nand U1566 (N_1566,In_1167,In_2520);
or U1567 (N_1567,In_2776,In_4300);
nor U1568 (N_1568,In_3802,In_1169);
nand U1569 (N_1569,In_1011,In_4980);
or U1570 (N_1570,In_1412,In_2621);
or U1571 (N_1571,In_3902,In_2862);
nor U1572 (N_1572,In_2152,In_2392);
nor U1573 (N_1573,In_961,In_1754);
and U1574 (N_1574,In_3790,In_2618);
nand U1575 (N_1575,In_3803,In_4341);
nor U1576 (N_1576,In_3960,In_1846);
or U1577 (N_1577,In_2614,In_904);
nand U1578 (N_1578,In_3106,In_2014);
xor U1579 (N_1579,In_3876,In_291);
and U1580 (N_1580,In_2199,In_1576);
and U1581 (N_1581,In_3763,In_672);
nor U1582 (N_1582,In_280,In_2426);
and U1583 (N_1583,In_1517,In_1044);
nand U1584 (N_1584,In_2982,In_3445);
or U1585 (N_1585,In_3772,In_3692);
or U1586 (N_1586,In_1952,In_1383);
and U1587 (N_1587,In_737,In_4199);
or U1588 (N_1588,In_2837,In_3245);
or U1589 (N_1589,In_554,In_2266);
and U1590 (N_1590,In_2463,In_2986);
and U1591 (N_1591,In_847,In_270);
and U1592 (N_1592,In_4960,In_815);
and U1593 (N_1593,In_4052,In_4799);
nand U1594 (N_1594,In_4602,In_1597);
nand U1595 (N_1595,In_826,In_1705);
or U1596 (N_1596,In_3225,In_2798);
nor U1597 (N_1597,In_3461,In_537);
nand U1598 (N_1598,In_633,In_3493);
xor U1599 (N_1599,In_3320,In_2938);
nand U1600 (N_1600,In_3970,In_2080);
nand U1601 (N_1601,In_2828,In_69);
and U1602 (N_1602,In_3004,In_1471);
and U1603 (N_1603,In_4188,In_485);
and U1604 (N_1604,In_3581,In_1334);
nand U1605 (N_1605,In_869,In_3877);
nand U1606 (N_1606,In_3340,In_4429);
nor U1607 (N_1607,In_3361,In_4274);
xor U1608 (N_1608,In_4459,In_4955);
and U1609 (N_1609,In_1279,In_4907);
nor U1610 (N_1610,In_3349,In_3437);
nor U1611 (N_1611,In_2817,In_3190);
or U1612 (N_1612,In_3589,In_3725);
nand U1613 (N_1613,In_1391,In_4440);
and U1614 (N_1614,In_4239,In_3557);
and U1615 (N_1615,In_3093,In_1627);
nand U1616 (N_1616,In_571,In_441);
nor U1617 (N_1617,In_659,In_1259);
and U1618 (N_1618,In_1036,In_2389);
nor U1619 (N_1619,In_975,In_1847);
and U1620 (N_1620,In_3738,In_3705);
nor U1621 (N_1621,In_1379,In_4839);
nor U1622 (N_1622,In_4181,In_4944);
nand U1623 (N_1623,In_528,In_4287);
nor U1624 (N_1624,In_2081,In_4089);
xor U1625 (N_1625,In_4707,In_4498);
xor U1626 (N_1626,In_538,In_3049);
xnor U1627 (N_1627,In_3108,In_4919);
xnor U1628 (N_1628,In_755,In_4493);
xor U1629 (N_1629,In_4456,In_1463);
or U1630 (N_1630,In_399,In_4113);
nand U1631 (N_1631,In_4470,In_3635);
xnor U1632 (N_1632,In_197,In_797);
nor U1633 (N_1633,In_355,In_1575);
xnor U1634 (N_1634,In_2613,In_130);
nor U1635 (N_1635,In_2638,In_2509);
xor U1636 (N_1636,In_3111,In_4094);
xnor U1637 (N_1637,In_2876,In_4206);
xor U1638 (N_1638,In_379,In_3207);
nand U1639 (N_1639,In_3515,In_4830);
nor U1640 (N_1640,In_4323,In_371);
or U1641 (N_1641,In_2690,In_114);
or U1642 (N_1642,In_3145,In_400);
or U1643 (N_1643,In_4182,In_4157);
or U1644 (N_1644,In_2706,In_2436);
xor U1645 (N_1645,In_1556,In_2432);
xnor U1646 (N_1646,In_3663,In_1455);
xor U1647 (N_1647,In_397,In_4841);
xor U1648 (N_1648,In_917,In_3825);
nor U1649 (N_1649,In_1633,In_2681);
and U1650 (N_1650,In_1950,In_4131);
or U1651 (N_1651,In_1693,In_3503);
or U1652 (N_1652,In_2659,In_4774);
and U1653 (N_1653,In_3312,In_456);
nor U1654 (N_1654,In_611,In_3546);
or U1655 (N_1655,In_222,In_2295);
nand U1656 (N_1656,In_1506,In_4108);
nand U1657 (N_1657,In_3252,In_2077);
and U1658 (N_1658,In_2009,In_4734);
nor U1659 (N_1659,In_1850,In_3734);
or U1660 (N_1660,In_3306,In_4963);
and U1661 (N_1661,In_2177,In_522);
nor U1662 (N_1662,In_1085,In_1132);
xor U1663 (N_1663,In_4642,In_707);
nor U1664 (N_1664,In_4449,In_2219);
nor U1665 (N_1665,In_1806,In_4381);
nand U1666 (N_1666,In_3198,In_253);
or U1667 (N_1667,In_1159,In_1210);
xnor U1668 (N_1668,In_2195,In_3566);
or U1669 (N_1669,In_935,In_3266);
nand U1670 (N_1670,In_324,In_1546);
or U1671 (N_1671,In_4422,In_2001);
and U1672 (N_1672,In_89,In_2722);
nor U1673 (N_1673,In_1856,In_4247);
nand U1674 (N_1674,In_2371,In_2539);
xnor U1675 (N_1675,In_1019,In_1791);
nor U1676 (N_1676,In_1255,In_285);
and U1677 (N_1677,In_4608,In_3085);
nor U1678 (N_1678,In_746,In_2129);
or U1679 (N_1679,In_2718,In_1100);
nor U1680 (N_1680,In_3873,In_3664);
nor U1681 (N_1681,In_4024,In_3813);
and U1682 (N_1682,In_4184,In_4399);
or U1683 (N_1683,In_4226,In_3820);
and U1684 (N_1684,In_3082,In_4647);
xnor U1685 (N_1685,In_1404,In_87);
nor U1686 (N_1686,In_2106,In_162);
nor U1687 (N_1687,In_4375,In_1842);
xor U1688 (N_1688,In_1106,In_277);
nor U1689 (N_1689,In_228,In_817);
and U1690 (N_1690,In_881,In_4176);
nor U1691 (N_1691,In_3090,In_3411);
and U1692 (N_1692,In_532,In_896);
nand U1693 (N_1693,In_500,In_948);
or U1694 (N_1694,In_2248,In_2835);
nor U1695 (N_1695,In_2191,In_3269);
and U1696 (N_1696,In_1997,In_1447);
and U1697 (N_1697,In_4143,In_804);
nor U1698 (N_1698,In_2402,In_4469);
nor U1699 (N_1699,In_906,In_3815);
xor U1700 (N_1700,In_4396,In_2061);
nor U1701 (N_1701,In_1616,In_381);
nor U1702 (N_1702,In_1828,In_115);
nand U1703 (N_1703,In_1035,In_2702);
xor U1704 (N_1704,In_635,In_3474);
nand U1705 (N_1705,In_2307,In_4986);
and U1706 (N_1706,In_1360,In_2345);
nor U1707 (N_1707,In_2317,In_4846);
and U1708 (N_1708,In_1472,In_1604);
nand U1709 (N_1709,In_2942,In_2471);
or U1710 (N_1710,In_870,In_3558);
and U1711 (N_1711,In_3469,In_1619);
nor U1712 (N_1712,In_2673,In_3081);
or U1713 (N_1713,In_4814,In_2599);
or U1714 (N_1714,In_1250,In_2410);
nand U1715 (N_1715,In_3430,In_1486);
and U1716 (N_1716,In_3238,In_1889);
and U1717 (N_1717,In_3356,In_4531);
and U1718 (N_1718,In_2089,In_4155);
or U1719 (N_1719,In_4250,In_1527);
or U1720 (N_1720,In_1690,In_4227);
nand U1721 (N_1721,In_416,In_3257);
or U1722 (N_1722,In_964,In_58);
nor U1723 (N_1723,In_523,In_1137);
nor U1724 (N_1724,In_2339,In_3419);
and U1725 (N_1725,In_2694,In_403);
nor U1726 (N_1726,In_670,In_1020);
or U1727 (N_1727,In_3434,In_3205);
nand U1728 (N_1728,In_2932,In_1201);
and U1729 (N_1729,In_2328,In_545);
and U1730 (N_1730,In_1786,In_2922);
xnor U1731 (N_1731,In_3529,In_4914);
or U1732 (N_1732,In_2747,In_3417);
nor U1733 (N_1733,In_3879,In_3982);
nand U1734 (N_1734,In_3616,In_2937);
nand U1735 (N_1735,In_305,In_1025);
or U1736 (N_1736,In_2964,In_4010);
nand U1737 (N_1737,In_1004,In_3487);
nand U1738 (N_1738,In_218,In_2777);
nand U1739 (N_1739,In_1727,In_4601);
or U1740 (N_1740,In_1121,In_3583);
nand U1741 (N_1741,In_2600,In_1985);
and U1742 (N_1742,In_173,In_3826);
nor U1743 (N_1743,In_3819,In_3829);
xnor U1744 (N_1744,In_4455,In_1573);
xnor U1745 (N_1745,In_2750,In_1243);
nor U1746 (N_1746,In_3683,In_1096);
xor U1747 (N_1747,In_4086,In_3850);
nand U1748 (N_1748,In_3535,In_496);
and U1749 (N_1749,In_2313,In_623);
nor U1750 (N_1750,In_1065,In_2849);
nand U1751 (N_1751,In_2975,In_1439);
xor U1752 (N_1752,In_4956,In_436);
and U1753 (N_1753,In_2347,In_2276);
xor U1754 (N_1754,In_3067,In_4168);
or U1755 (N_1755,In_2738,In_2955);
nor U1756 (N_1756,In_1960,In_2535);
or U1757 (N_1757,In_3893,In_3903);
and U1758 (N_1758,In_4898,In_3810);
or U1759 (N_1759,In_753,In_3595);
and U1760 (N_1760,In_3289,In_512);
and U1761 (N_1761,In_3342,In_4693);
nor U1762 (N_1762,In_3640,In_2263);
or U1763 (N_1763,In_2530,In_2281);
or U1764 (N_1764,In_1303,In_1734);
nor U1765 (N_1765,In_3425,In_920);
and U1766 (N_1766,In_1767,In_1568);
nand U1767 (N_1767,In_4346,In_4152);
xor U1768 (N_1768,In_386,In_4736);
nor U1769 (N_1769,In_1899,In_2588);
or U1770 (N_1770,In_3382,In_3076);
xnor U1771 (N_1771,In_1996,In_334);
nand U1772 (N_1772,In_3659,In_874);
xnor U1773 (N_1773,In_4674,In_2230);
nand U1774 (N_1774,In_2365,In_2799);
xnor U1775 (N_1775,In_796,In_3704);
nand U1776 (N_1776,In_1758,In_3690);
xor U1777 (N_1777,In_4547,In_1082);
and U1778 (N_1778,In_209,In_3913);
or U1779 (N_1779,In_3949,In_3128);
or U1780 (N_1780,In_779,In_4922);
xnor U1781 (N_1781,In_928,In_1277);
and U1782 (N_1782,In_2110,In_2698);
and U1783 (N_1783,In_2740,In_2772);
nand U1784 (N_1784,In_2944,In_2935);
nor U1785 (N_1785,In_884,In_2043);
xor U1786 (N_1786,In_824,In_1321);
nand U1787 (N_1787,In_18,In_1509);
xor U1788 (N_1788,In_2543,In_3258);
and U1789 (N_1789,In_3177,In_2611);
xnor U1790 (N_1790,In_1007,In_3775);
xor U1791 (N_1791,In_1555,In_4216);
xor U1792 (N_1792,In_4623,In_4175);
xor U1793 (N_1793,In_803,In_619);
or U1794 (N_1794,In_1023,In_393);
xnor U1795 (N_1795,In_2023,In_2766);
or U1796 (N_1796,In_3737,In_3703);
nor U1797 (N_1797,In_168,In_681);
nand U1798 (N_1798,In_2827,In_3168);
nor U1799 (N_1799,In_1409,In_446);
nand U1800 (N_1800,In_3549,In_1168);
nand U1801 (N_1801,In_1048,In_3848);
nor U1802 (N_1802,In_3836,In_3653);
and U1803 (N_1803,In_1902,In_4074);
and U1804 (N_1804,In_1434,In_4924);
and U1805 (N_1805,In_2468,In_3068);
nand U1806 (N_1806,In_513,In_2512);
and U1807 (N_1807,In_118,In_837);
and U1808 (N_1808,In_4568,In_3092);
or U1809 (N_1809,In_1302,In_1188);
nor U1810 (N_1810,In_4473,In_3221);
nor U1811 (N_1811,In_4735,In_4812);
or U1812 (N_1812,In_594,In_4930);
nand U1813 (N_1813,In_4679,In_4051);
xor U1814 (N_1814,In_3072,In_1893);
or U1815 (N_1815,In_82,In_4967);
nand U1816 (N_1816,In_963,In_3791);
xor U1817 (N_1817,In_3582,In_4248);
or U1818 (N_1818,In_1541,In_4252);
nor U1819 (N_1819,In_262,In_2626);
and U1820 (N_1820,In_3714,In_2627);
or U1821 (N_1821,In_3402,In_1745);
or U1822 (N_1822,In_2470,In_438);
or U1823 (N_1823,In_2413,In_263);
or U1824 (N_1824,In_4797,In_147);
xnor U1825 (N_1825,In_780,In_1239);
nor U1826 (N_1826,In_1336,In_3637);
nand U1827 (N_1827,In_1759,In_866);
or U1828 (N_1828,In_288,In_3568);
or U1829 (N_1829,In_3921,In_1390);
nand U1830 (N_1830,In_4551,In_4319);
or U1831 (N_1831,In_2004,In_2355);
or U1832 (N_1832,In_1978,In_665);
and U1833 (N_1833,In_4612,In_1513);
nand U1834 (N_1834,In_3051,In_4916);
xnor U1835 (N_1835,In_1179,In_3429);
and U1836 (N_1836,In_1405,In_1988);
xor U1837 (N_1837,In_1402,In_2167);
nand U1838 (N_1838,In_4584,In_2884);
or U1839 (N_1839,In_4760,In_3842);
or U1840 (N_1840,In_4775,In_1815);
xnor U1841 (N_1841,In_3019,In_923);
and U1842 (N_1842,In_4445,In_3817);
and U1843 (N_1843,In_2022,In_3684);
and U1844 (N_1844,In_2567,In_4393);
and U1845 (N_1845,In_899,In_4162);
nor U1846 (N_1846,In_1886,In_1811);
or U1847 (N_1847,In_2961,In_2429);
nor U1848 (N_1848,In_1125,In_1822);
nor U1849 (N_1849,In_3240,In_3980);
xor U1850 (N_1850,In_3846,In_2063);
nand U1851 (N_1851,In_2877,In_64);
nand U1852 (N_1852,In_1792,In_1821);
and U1853 (N_1853,In_2661,In_1423);
nor U1854 (N_1854,In_3855,In_1697);
nor U1855 (N_1855,In_4977,In_3050);
and U1856 (N_1856,In_834,In_1749);
nor U1857 (N_1857,In_2083,In_372);
xnor U1858 (N_1858,In_1535,In_4101);
and U1859 (N_1859,In_3656,In_2895);
or U1860 (N_1860,In_1017,In_3749);
xor U1861 (N_1861,In_1331,In_2155);
and U1862 (N_1862,In_660,In_1521);
and U1863 (N_1863,In_1103,In_206);
xnor U1864 (N_1864,In_3341,In_2473);
nand U1865 (N_1865,In_2025,In_1698);
xor U1866 (N_1866,In_1859,In_1145);
xor U1867 (N_1867,In_3156,In_1712);
nor U1868 (N_1868,In_2034,In_1490);
xor U1869 (N_1869,In_2050,In_2383);
nand U1870 (N_1870,In_1917,In_4578);
and U1871 (N_1871,In_2409,In_2026);
xor U1872 (N_1872,In_3644,In_2761);
nand U1873 (N_1873,In_3928,In_2991);
nor U1874 (N_1874,In_470,In_1694);
nor U1875 (N_1875,In_202,In_216);
and U1876 (N_1876,In_2680,In_630);
nor U1877 (N_1877,In_1984,In_2560);
and U1878 (N_1878,In_3631,In_2312);
xnor U1879 (N_1879,In_1922,In_624);
xor U1880 (N_1880,In_2422,In_3950);
nand U1881 (N_1881,In_1052,In_1600);
or U1882 (N_1882,In_3989,In_1545);
xor U1883 (N_1883,In_1939,In_3069);
and U1884 (N_1884,In_3700,In_4451);
xor U1885 (N_1885,In_1926,In_3230);
nor U1886 (N_1886,In_367,In_4087);
xor U1887 (N_1887,In_186,In_4266);
nor U1888 (N_1888,In_3645,In_705);
and U1889 (N_1889,In_4174,In_693);
nand U1890 (N_1890,In_422,In_4921);
xor U1891 (N_1891,In_4420,In_1190);
or U1892 (N_1892,In_3475,In_852);
or U1893 (N_1893,In_158,In_4758);
xnor U1894 (N_1894,In_4442,In_3113);
and U1895 (N_1895,In_4715,In_1746);
or U1896 (N_1896,In_2743,In_2856);
xnor U1897 (N_1897,In_3730,In_959);
nor U1898 (N_1898,In_2630,In_1382);
nand U1899 (N_1899,In_4510,In_3718);
xnor U1900 (N_1900,In_1338,In_4958);
nand U1901 (N_1901,In_473,In_4546);
nand U1902 (N_1902,In_3491,In_2815);
and U1903 (N_1903,In_3721,In_4038);
or U1904 (N_1904,In_4481,In_2920);
nand U1905 (N_1905,In_2208,In_4609);
and U1906 (N_1906,In_3302,In_738);
and U1907 (N_1907,In_2921,In_820);
nor U1908 (N_1908,In_3860,In_4889);
nor U1909 (N_1909,In_4416,In_2170);
and U1910 (N_1910,In_4836,In_774);
and U1911 (N_1911,In_3011,In_4496);
and U1912 (N_1912,In_3588,In_4718);
nand U1913 (N_1913,In_417,In_4522);
or U1914 (N_1914,In_4487,In_2310);
and U1915 (N_1915,In_1107,In_70);
or U1916 (N_1916,In_3506,In_4650);
and U1917 (N_1917,In_102,In_3124);
nor U1918 (N_1918,In_283,In_2524);
xnor U1919 (N_1919,In_3591,In_3908);
nor U1920 (N_1920,In_2019,In_4354);
xor U1921 (N_1921,In_4237,In_1457);
nand U1922 (N_1922,In_1400,In_489);
nor U1923 (N_1923,In_3326,In_411);
xor U1924 (N_1924,In_480,In_4512);
nand U1925 (N_1925,In_4020,In_125);
and U1926 (N_1926,In_2302,In_3427);
nand U1927 (N_1927,In_3186,In_4684);
xnor U1928 (N_1928,In_2112,In_985);
nor U1929 (N_1929,In_4000,In_2758);
nor U1930 (N_1930,In_1676,In_2918);
or U1931 (N_1931,In_275,In_3317);
xor U1932 (N_1932,In_4048,In_1270);
or U1933 (N_1933,In_1775,In_4706);
nor U1934 (N_1934,In_3657,In_329);
xor U1935 (N_1935,In_1042,In_3173);
nor U1936 (N_1936,In_1000,In_1332);
nor U1937 (N_1937,In_4339,In_683);
and U1938 (N_1938,In_2224,In_1055);
nor U1939 (N_1939,In_2464,In_1748);
nor U1940 (N_1940,In_1779,In_2585);
xor U1941 (N_1941,In_1362,In_781);
or U1942 (N_1942,In_1961,In_1194);
nor U1943 (N_1943,In_3008,In_4714);
or U1944 (N_1944,In_2257,In_2303);
nand U1945 (N_1945,In_2582,In_3841);
or U1946 (N_1946,In_1062,In_3060);
nand U1947 (N_1947,In_1649,In_156);
nor U1948 (N_1948,In_2859,In_1207);
and U1949 (N_1949,In_4769,In_4254);
nor U1950 (N_1950,In_2326,In_1318);
nor U1951 (N_1951,In_4552,In_1214);
nor U1952 (N_1952,In_4070,In_4864);
or U1953 (N_1953,In_3723,In_2855);
nand U1954 (N_1954,In_3793,In_1973);
and U1955 (N_1955,In_4768,In_1130);
xor U1956 (N_1956,In_1060,In_3715);
and U1957 (N_1957,In_3909,In_3083);
or U1958 (N_1958,In_1217,In_375);
xor U1959 (N_1959,In_3389,In_31);
and U1960 (N_1960,In_541,In_794);
or U1961 (N_1961,In_1901,In_3485);
and U1962 (N_1962,In_4093,In_4045);
nor U1963 (N_1963,In_800,In_3380);
xor U1964 (N_1964,In_3768,In_307);
xor U1965 (N_1965,In_4822,In_4221);
xnor U1966 (N_1966,In_2547,In_1133);
or U1967 (N_1967,In_1479,In_741);
and U1968 (N_1968,In_1266,In_4874);
and U1969 (N_1969,In_2787,In_1678);
nand U1970 (N_1970,In_706,In_3765);
xor U1971 (N_1971,In_3689,In_2631);
xnor U1972 (N_1972,In_4461,In_2591);
and U1973 (N_1973,In_926,In_123);
and U1974 (N_1974,In_1592,In_4933);
or U1975 (N_1975,In_4751,In_2388);
and U1976 (N_1976,In_761,In_2554);
xnor U1977 (N_1977,In_396,In_250);
or U1978 (N_1978,In_1773,In_3966);
and U1979 (N_1979,In_675,In_4644);
nor U1980 (N_1980,In_4356,In_3962);
and U1981 (N_1981,In_3368,In_4657);
and U1982 (N_1982,In_2978,In_2264);
xnor U1983 (N_1983,In_1357,In_1523);
nand U1984 (N_1984,In_682,In_4954);
and U1985 (N_1985,In_2366,In_3531);
nor U1986 (N_1986,In_1641,In_1943);
nand U1987 (N_1987,In_2791,In_1451);
and U1988 (N_1988,In_191,In_1919);
and U1989 (N_1989,In_4400,In_3787);
nand U1990 (N_1990,In_1366,In_543);
or U1991 (N_1991,In_4013,In_3448);
nor U1992 (N_1992,In_3407,In_2959);
nor U1993 (N_1993,In_1937,In_4165);
and U1994 (N_1994,In_2156,In_4137);
or U1995 (N_1995,In_1196,In_851);
xnor U1996 (N_1996,In_2969,In_1291);
nand U1997 (N_1997,In_4831,In_4410);
nand U1998 (N_1998,In_172,In_1797);
nor U1999 (N_1999,In_1968,In_2042);
nand U2000 (N_2000,N_1525,In_2775);
nor U2001 (N_2001,In_1967,In_4488);
xor U2002 (N_2002,N_977,N_1242);
xnor U2003 (N_2003,N_1324,N_972);
nor U2004 (N_2004,In_2830,In_3188);
nand U2005 (N_2005,N_1118,N_1553);
nand U2006 (N_2006,In_2953,N_1070);
and U2007 (N_2007,N_1057,N_1277);
xnor U2008 (N_2008,N_1496,N_416);
xnor U2009 (N_2009,In_3373,N_34);
or U2010 (N_2010,N_21,In_3390);
or U2011 (N_2011,In_4762,In_2213);
xnor U2012 (N_2012,In_673,N_1948);
nand U2013 (N_2013,N_1020,N_1790);
nor U2014 (N_2014,N_1532,In_2608);
or U2015 (N_2015,In_3182,In_3613);
or U2016 (N_2016,In_2565,N_671);
nor U2017 (N_2017,N_843,N_1292);
xor U2018 (N_2018,N_1212,N_1391);
xor U2019 (N_2019,In_1070,In_2086);
or U2020 (N_2020,N_1715,N_285);
and U2021 (N_2021,N_1643,In_4654);
nand U2022 (N_2022,N_1008,N_779);
and U2023 (N_2023,N_1741,N_704);
xor U2024 (N_2024,N_591,In_144);
nand U2025 (N_2025,N_952,N_507);
and U2026 (N_2026,N_407,N_1869);
nand U2027 (N_2027,N_903,In_77);
and U2028 (N_2028,N_697,N_1484);
nand U2029 (N_2029,N_753,N_1755);
nor U2030 (N_2030,N_1540,In_458);
nor U2031 (N_2031,N_83,In_1532);
nor U2032 (N_2032,N_1076,N_598);
nand U2033 (N_2033,N_600,N_1241);
and U2034 (N_2034,N_1,N_1421);
nand U2035 (N_2035,In_25,N_1920);
xnor U2036 (N_2036,In_2823,In_3658);
xor U2037 (N_2037,In_1166,In_1297);
and U2038 (N_2038,N_320,In_1608);
and U2039 (N_2039,N_35,In_2143);
xnor U2040 (N_2040,In_4466,N_831);
and U2041 (N_2041,In_4269,N_1021);
and U2042 (N_2042,N_1125,N_1883);
xnor U2043 (N_2043,N_1996,N_1162);
and U2044 (N_2044,N_1139,In_2909);
nor U2045 (N_2045,In_895,N_851);
and U2046 (N_2046,N_1402,N_794);
xnor U2047 (N_2047,N_913,N_867);
nand U2048 (N_2048,N_383,N_1624);
and U2049 (N_2049,In_4925,N_1739);
nand U2050 (N_2050,N_1602,In_1805);
and U2051 (N_2051,N_1301,N_1264);
nor U2052 (N_2052,In_2782,N_795);
and U2053 (N_2053,N_933,N_681);
xor U2054 (N_2054,N_1059,In_789);
nor U2055 (N_2055,In_1068,N_1583);
and U2056 (N_2056,N_220,In_1104);
and U2057 (N_2057,N_338,In_2445);
nand U2058 (N_2058,N_822,N_1669);
and U2059 (N_2059,In_3843,N_1718);
nor U2060 (N_2060,N_839,In_4103);
xnor U2061 (N_2061,N_1219,In_4906);
xnor U2062 (N_2062,N_907,In_1269);
nand U2063 (N_2063,N_608,In_855);
or U2064 (N_2064,N_520,N_374);
xor U2065 (N_2065,In_423,N_752);
xor U2066 (N_2066,N_1198,N_1792);
nand U2067 (N_2067,In_4637,N_1375);
or U2068 (N_2068,In_4008,N_1362);
xnor U2069 (N_2069,N_1877,N_1133);
nor U2070 (N_2070,N_773,N_723);
nor U2071 (N_2071,In_3119,In_2041);
or U2072 (N_2072,N_748,In_80);
and U2073 (N_2073,In_4988,N_882);
xnor U2074 (N_2074,N_1810,In_2040);
or U2075 (N_2075,In_4793,N_1904);
nand U2076 (N_2076,N_175,N_1510);
or U2077 (N_2077,N_833,N_1440);
or U2078 (N_2078,In_3954,N_574);
nor U2079 (N_2079,N_70,N_844);
xor U2080 (N_2080,In_1862,N_615);
nand U2081 (N_2081,N_1243,N_1007);
nor U2082 (N_2082,N_1685,In_1182);
nand U2083 (N_2083,N_1462,N_620);
or U2084 (N_2084,N_64,In_2062);
nand U2085 (N_2085,N_841,N_309);
xor U2086 (N_2086,In_2648,N_206);
or U2087 (N_2087,N_1982,N_514);
or U2088 (N_2088,N_1803,N_891);
xnor U2089 (N_2089,In_2216,N_363);
xnor U2090 (N_2090,In_2976,In_831);
nor U2091 (N_2091,N_1594,In_592);
nor U2092 (N_2092,N_151,N_1272);
xnor U2093 (N_2093,In_1646,N_1121);
or U2094 (N_2094,N_1665,N_18);
and U2095 (N_2095,N_1706,N_1597);
nor U2096 (N_2096,In_3117,N_1922);
or U2097 (N_2097,In_2757,In_696);
xor U2098 (N_2098,N_17,In_1393);
and U2099 (N_2099,N_858,In_657);
nand U2100 (N_2100,N_1040,In_86);
nor U2101 (N_2101,N_1795,In_2245);
or U2102 (N_2102,N_85,N_1742);
xor U2103 (N_2103,N_989,N_193);
xor U2104 (N_2104,In_3981,In_1253);
and U2105 (N_2105,N_1774,N_20);
xor U2106 (N_2106,N_1379,N_1932);
or U2107 (N_2107,In_3097,N_787);
or U2108 (N_2108,In_4448,N_108);
nor U2109 (N_2109,In_1226,In_447);
or U2110 (N_2110,N_483,In_1155);
or U2111 (N_2111,In_3480,In_2145);
and U2112 (N_2112,N_1545,N_234);
or U2113 (N_2113,N_266,In_3660);
xnor U2114 (N_2114,In_2059,N_842);
xnor U2115 (N_2115,N_394,N_216);
nand U2116 (N_2116,N_498,N_605);
nor U2117 (N_2117,In_14,N_1122);
nor U2118 (N_2118,In_694,N_864);
nand U2119 (N_2119,In_433,N_1854);
nand U2120 (N_2120,N_1963,In_4308);
or U2121 (N_2121,N_1182,N_735);
nor U2122 (N_2122,N_862,N_966);
and U2123 (N_2123,In_3638,N_1991);
or U2124 (N_2124,N_1200,N_838);
or U2125 (N_2125,N_393,In_894);
xnor U2126 (N_2126,N_88,N_1295);
nand U2127 (N_2127,N_321,N_627);
or U2128 (N_2128,In_2144,N_496);
or U2129 (N_2129,N_1989,N_525);
and U2130 (N_2130,In_3321,In_1552);
nand U2131 (N_2131,N_1546,N_744);
nand U2132 (N_2132,N_378,In_4350);
nand U2133 (N_2133,N_602,N_810);
nand U2134 (N_2134,In_1738,In_1325);
and U2135 (N_2135,In_4648,N_1754);
or U2136 (N_2136,N_550,N_37);
xnor U2137 (N_2137,N_428,N_306);
nand U2138 (N_2138,In_2398,N_1926);
and U2139 (N_2139,N_226,In_4021);
xor U2140 (N_2140,In_4622,N_865);
or U2141 (N_2141,N_12,In_772);
nand U2142 (N_2142,N_1082,N_144);
nand U2143 (N_2143,N_96,In_1119);
and U2144 (N_2144,N_478,In_4272);
or U2145 (N_2145,In_2494,N_1183);
xor U2146 (N_2146,N_273,In_3136);
xor U2147 (N_2147,N_521,N_1247);
nand U2148 (N_2148,N_352,In_2664);
and U2149 (N_2149,N_800,In_4989);
nor U2150 (N_2150,N_275,In_678);
or U2151 (N_2151,In_4129,In_20);
or U2152 (N_2152,N_596,N_249);
and U2153 (N_2153,In_4432,In_1066);
nor U2154 (N_2154,N_1717,N_1766);
and U2155 (N_2155,In_4582,In_1006);
nand U2156 (N_2156,N_1584,N_1923);
nor U2157 (N_2157,N_229,In_256);
nand U2158 (N_2158,N_476,N_364);
and U2159 (N_2159,N_1073,N_481);
or U2160 (N_2160,N_887,N_1666);
or U2161 (N_2161,N_946,N_641);
nor U2162 (N_2162,N_424,N_1734);
xor U2163 (N_2163,N_180,In_518);
or U2164 (N_2164,N_1526,N_876);
xor U2165 (N_2165,N_1966,N_869);
and U2166 (N_2166,N_1001,N_329);
nor U2167 (N_2167,In_4025,In_4379);
nand U2168 (N_2168,N_1498,In_1870);
nor U2169 (N_2169,N_1935,N_1335);
or U2170 (N_2170,N_75,N_207);
nand U2171 (N_2171,N_1617,In_2162);
nand U2172 (N_2172,N_1763,N_1671);
xnor U2173 (N_2173,In_4196,In_1881);
nor U2174 (N_2174,N_1684,N_1651);
and U2175 (N_2175,In_1585,N_917);
xor U2176 (N_2176,In_1309,N_272);
nand U2177 (N_2177,N_472,N_656);
and U2178 (N_2178,N_1676,N_182);
or U2179 (N_2179,N_590,N_1645);
nand U2180 (N_2180,In_2098,N_1165);
xnor U2181 (N_2181,N_432,N_1449);
nor U2182 (N_2182,In_2331,In_4222);
xor U2183 (N_2183,N_1945,N_1056);
nor U2184 (N_2184,In_1041,N_71);
or U2185 (N_2185,N_1163,In_2092);
nand U2186 (N_2186,In_1735,N_1796);
and U2187 (N_2187,N_613,N_1481);
and U2188 (N_2188,N_1675,N_1899);
nand U2189 (N_2189,N_1314,In_463);
xor U2190 (N_2190,N_1644,N_1039);
and U2191 (N_2191,In_2858,In_1367);
xor U2192 (N_2192,In_4821,In_3586);
or U2193 (N_2193,N_818,N_1354);
and U2194 (N_2194,N_1610,N_48);
xor U2195 (N_2195,N_1824,N_201);
or U2196 (N_2196,N_804,N_429);
nand U2197 (N_2197,In_1778,N_927);
nand U2198 (N_2198,N_616,N_43);
or U2199 (N_2199,N_1010,N_1129);
nor U2200 (N_2200,N_1144,N_883);
xor U2201 (N_2201,In_1098,N_323);
and U2202 (N_2202,N_72,N_1063);
or U2203 (N_2203,N_420,In_4862);
or U2204 (N_2204,In_1046,N_390);
xor U2205 (N_2205,N_541,N_80);
and U2206 (N_2206,N_1290,N_1975);
or U2207 (N_2207,In_4238,N_1760);
xnor U2208 (N_2208,N_1099,N_668);
nand U2209 (N_2209,In_1986,In_3375);
or U2210 (N_2210,In_3923,N_1471);
nand U2211 (N_2211,N_633,N_1045);
nand U2212 (N_2212,N_1090,N_198);
nor U2213 (N_2213,N_1841,In_242);
nor U2214 (N_2214,N_1522,N_1579);
xor U2215 (N_2215,In_3255,N_1343);
nand U2216 (N_2216,N_850,In_3945);
nor U2217 (N_2217,N_1155,N_1972);
and U2218 (N_2218,In_3422,N_951);
nor U2219 (N_2219,N_1246,N_1486);
or U2220 (N_2220,N_1901,N_421);
nor U2221 (N_2221,N_1033,In_1162);
nor U2222 (N_2222,In_478,N_1042);
xor U2223 (N_2223,N_1918,N_170);
nand U2224 (N_2224,In_4504,In_1723);
or U2225 (N_2225,N_1327,In_3767);
or U2226 (N_2226,N_205,N_1523);
and U2227 (N_2227,In_999,N_1960);
nor U2228 (N_2228,N_65,N_1848);
and U2229 (N_2229,In_4081,In_1252);
xor U2230 (N_2230,N_662,N_1613);
and U2231 (N_2231,N_1515,N_1764);
nand U2232 (N_2232,N_1323,In_1508);
nor U2233 (N_2233,N_988,N_857);
or U2234 (N_2234,In_2012,N_1470);
or U2235 (N_2235,N_943,N_1424);
nand U2236 (N_2236,In_3077,N_836);
nand U2237 (N_2237,N_204,In_4705);
or U2238 (N_2238,In_1466,In_3228);
and U2239 (N_2239,N_1611,N_1184);
nand U2240 (N_2240,In_4345,N_533);
nor U2241 (N_2241,In_4458,N_1022);
nor U2242 (N_2242,In_1160,N_425);
and U2243 (N_2243,In_2839,N_196);
nand U2244 (N_2244,In_2434,N_629);
and U2245 (N_2245,In_2913,N_592);
or U2246 (N_2246,N_1363,N_403);
or U2247 (N_2247,N_895,N_202);
and U2248 (N_2248,N_1800,In_4985);
or U2249 (N_2249,N_1957,N_149);
and U2250 (N_2250,In_2385,N_1320);
nor U2251 (N_2251,N_1776,N_1917);
nor U2252 (N_2252,N_322,N_1003);
and U2253 (N_2253,In_945,N_1979);
nand U2254 (N_2254,In_2609,N_1322);
or U2255 (N_2255,N_1539,In_859);
or U2256 (N_2256,N_141,N_209);
and U2257 (N_2257,N_1655,N_1887);
or U2258 (N_2258,In_418,N_189);
nand U2259 (N_2259,N_1307,In_2121);
xor U2260 (N_2260,N_926,N_1652);
or U2261 (N_2261,In_520,In_1730);
nor U2262 (N_2262,N_1697,In_4840);
xnor U2263 (N_2263,N_1708,N_333);
nand U2264 (N_2264,N_1068,N_1618);
or U2265 (N_2265,N_859,In_3104);
nor U2266 (N_2266,In_2379,N_547);
xnor U2267 (N_2267,N_1709,N_1358);
xor U2268 (N_2268,N_106,N_1822);
nand U2269 (N_2269,In_133,N_1194);
and U2270 (N_2270,N_1037,N_15);
nand U2271 (N_2271,N_132,N_1973);
and U2272 (N_2272,N_689,In_356);
and U2273 (N_2273,N_1128,N_655);
nand U2274 (N_2274,In_4636,N_350);
and U2275 (N_2275,In_1208,In_3249);
nand U2276 (N_2276,N_975,In_850);
xor U2277 (N_2277,In_4711,N_117);
or U2278 (N_2278,N_601,N_799);
and U2279 (N_2279,N_461,N_480);
nor U2280 (N_2280,N_1101,N_938);
nor U2281 (N_2281,N_1171,N_1479);
nor U2282 (N_2282,N_297,In_16);
or U2283 (N_2283,N_86,In_4672);
nor U2284 (N_2284,In_4132,N_556);
xor U2285 (N_2285,In_3486,N_287);
nor U2286 (N_2286,In_905,In_2229);
xor U2287 (N_2287,In_4460,N_734);
nor U2288 (N_2288,N_1113,In_1299);
and U2289 (N_2289,N_906,N_994);
and U2290 (N_2290,N_1662,N_1124);
nand U2291 (N_2291,In_2593,N_715);
and U2292 (N_2292,N_243,N_431);
nand U2293 (N_2293,N_958,N_712);
nor U2294 (N_2294,N_118,In_1064);
and U2295 (N_2295,N_1779,In_4694);
nor U2296 (N_2296,N_1293,In_3636);
nand U2297 (N_2297,N_1572,In_4138);
xor U2298 (N_2298,N_218,N_462);
or U2299 (N_2299,N_409,N_560);
nor U2300 (N_2300,N_852,N_729);
xor U2301 (N_2301,N_1952,N_1160);
nor U2302 (N_2302,N_1062,N_240);
and U2303 (N_2303,N_411,N_194);
nor U2304 (N_2304,In_967,N_1338);
and U2305 (N_2305,N_484,N_1825);
and U2306 (N_2306,In_606,In_748);
nor U2307 (N_2307,N_1844,N_241);
and U2308 (N_2308,N_49,N_1938);
xnor U2309 (N_2309,N_1051,In_3899);
xnor U2310 (N_2310,In_2444,N_1980);
nor U2311 (N_2311,N_545,N_1149);
or U2312 (N_2312,N_1340,In_3890);
nor U2313 (N_2313,N_875,N_588);
xnor U2314 (N_2314,In_823,N_1360);
and U2315 (N_2315,In_2538,N_423);
or U2316 (N_2316,N_371,In_2184);
xnor U2317 (N_2317,In_1170,In_1022);
or U2318 (N_2318,N_185,In_3044);
and U2319 (N_2319,N_1209,In_1642);
nand U2320 (N_2320,N_1970,N_522);
or U2321 (N_2321,N_1521,N_344);
or U2322 (N_2322,N_255,N_1456);
nand U2323 (N_2323,N_99,In_1925);
nand U2324 (N_2324,In_3353,N_730);
nand U2325 (N_2325,In_1531,N_1458);
or U2326 (N_2326,N_1131,In_1138);
or U2327 (N_2327,N_747,N_1403);
or U2328 (N_2328,N_97,N_485);
and U2329 (N_2329,N_7,In_838);
xnor U2330 (N_2330,N_1649,In_2460);
and U2331 (N_2331,N_1081,N_1890);
nor U2332 (N_2332,N_1262,N_1053);
xor U2333 (N_2333,N_731,N_583);
or U2334 (N_2334,N_1312,N_1574);
and U2335 (N_2335,N_282,In_214);
nand U2336 (N_2336,N_22,N_419);
and U2337 (N_2337,In_685,N_1965);
nor U2338 (N_2338,N_683,N_1705);
nand U2339 (N_2339,In_2361,N_725);
or U2340 (N_2340,N_1691,N_1758);
nand U2341 (N_2341,N_1164,N_860);
or U2342 (N_2342,In_552,N_1761);
nand U2343 (N_2343,In_4574,In_4003);
nand U2344 (N_2344,N_1370,N_1048);
nor U2345 (N_2345,In_4316,In_3976);
nor U2346 (N_2346,In_887,N_1808);
or U2347 (N_2347,In_2239,N_1030);
nor U2348 (N_2348,In_4161,In_3821);
xor U2349 (N_2349,N_879,N_1944);
nor U2350 (N_2350,N_147,In_3479);
and U2351 (N_2351,N_488,N_1964);
nand U2352 (N_2352,N_768,N_1104);
nand U2353 (N_2353,In_140,N_801);
nor U2354 (N_2354,N_918,In_2759);
xnor U2355 (N_2355,N_1298,In_4848);
or U2356 (N_2356,In_4169,N_642);
or U2357 (N_2357,In_3089,N_469);
or U2358 (N_2358,N_1564,N_174);
xnor U2359 (N_2359,N_617,N_781);
and U2360 (N_2360,N_854,N_1940);
nor U2361 (N_2361,N_1527,In_4770);
nor U2362 (N_2362,N_295,N_274);
or U2363 (N_2363,In_729,In_3408);
and U2364 (N_2364,N_817,N_967);
xnor U2365 (N_2365,N_1223,N_1388);
nand U2366 (N_2366,N_1900,In_2912);
xor U2367 (N_2367,In_2483,N_1596);
nor U2368 (N_2368,In_4324,N_25);
nor U2369 (N_2369,In_4260,In_2126);
nor U2370 (N_2370,In_4133,N_1680);
nor U2371 (N_2371,N_203,In_1337);
or U2372 (N_2372,N_1429,N_1703);
or U2373 (N_2373,N_826,In_4016);
nor U2374 (N_2374,N_181,N_985);
nand U2375 (N_2375,N_912,N_46);
xnor U2376 (N_2376,N_1927,In_4383);
and U2377 (N_2377,N_1018,N_871);
nor U2378 (N_2378,N_1078,In_4670);
xnor U2379 (N_2379,N_232,N_279);
and U2380 (N_2380,In_2727,In_1322);
or U2381 (N_2381,In_336,N_1993);
xor U2382 (N_2382,N_1276,In_3490);
nor U2383 (N_2383,N_1988,N_1411);
and U2384 (N_2384,In_2438,In_2262);
and U2385 (N_2385,N_422,In_819);
xnor U2386 (N_2386,In_2833,N_1064);
nand U2387 (N_2387,N_292,N_55);
nor U2388 (N_2388,N_1269,N_1404);
nand U2389 (N_2389,N_31,In_1204);
or U2390 (N_2390,N_1495,N_1336);
and U2391 (N_2391,N_1942,N_761);
xnor U2392 (N_2392,In_3418,N_1749);
xor U2393 (N_2393,N_1573,N_370);
and U2394 (N_2394,In_2695,N_1011);
nand U2395 (N_2395,N_962,In_1422);
nand U2396 (N_2396,N_540,N_1263);
xnor U2397 (N_2397,N_1413,N_1002);
xor U2398 (N_2398,N_1308,N_700);
nand U2399 (N_2399,In_4689,N_314);
and U2400 (N_2400,N_707,In_4271);
nor U2401 (N_2401,In_4297,In_3619);
nand U2402 (N_2402,In_4811,N_1491);
xnor U2403 (N_2403,In_299,In_2686);
and U2404 (N_2404,N_283,N_176);
and U2405 (N_2405,N_1156,In_3627);
nand U2406 (N_2406,N_502,N_714);
or U2407 (N_2407,In_3063,In_2321);
nor U2408 (N_2408,N_524,N_1633);
xor U2409 (N_2409,N_1505,N_1580);
nand U2410 (N_2410,N_1864,N_1444);
and U2411 (N_2411,N_349,N_150);
or U2412 (N_2412,N_1519,N_1647);
or U2413 (N_2413,N_919,N_1317);
nand U2414 (N_2414,N_331,N_1568);
nand U2415 (N_2415,N_1170,N_1346);
or U2416 (N_2416,In_2151,In_2035);
and U2417 (N_2417,N_1700,N_1216);
nand U2418 (N_2418,N_1488,In_4526);
nor U2419 (N_2419,N_98,In_2724);
nor U2420 (N_2420,N_580,In_52);
nor U2421 (N_2421,N_1382,N_1248);
xnor U2422 (N_2422,N_928,N_1225);
xnor U2423 (N_2423,In_679,N_1853);
and U2424 (N_2424,In_1648,N_920);
xnor U2425 (N_2425,N_1032,N_1821);
or U2426 (N_2426,N_1809,N_1968);
xnor U2427 (N_2427,In_602,N_257);
nor U2428 (N_2428,In_2657,N_1934);
nand U2429 (N_2429,In_116,N_1892);
nand U2430 (N_2430,N_1772,In_2763);
nand U2431 (N_2431,In_1386,In_740);
and U2432 (N_2432,N_1193,N_1047);
nand U2433 (N_2433,N_1398,N_1028);
nand U2434 (N_2434,In_236,N_442);
xor U2435 (N_2435,N_120,In_3311);
and U2436 (N_2436,In_3284,In_1316);
nor U2437 (N_2437,N_1017,N_763);
or U2438 (N_2438,In_3000,N_610);
nor U2439 (N_2439,N_1366,N_1091);
and U2440 (N_2440,N_231,N_1386);
and U2441 (N_2441,N_1218,N_1740);
and U2442 (N_2442,In_4997,N_1454);
nand U2443 (N_2443,In_1674,In_3365);
or U2444 (N_2444,In_4629,N_1357);
nor U2445 (N_2445,N_1773,In_1612);
nand U2446 (N_2446,In_244,N_152);
or U2447 (N_2447,N_1214,N_1482);
xnor U2448 (N_2448,N_848,N_577);
xnor U2449 (N_2449,In_2910,N_1635);
xor U2450 (N_2450,N_1369,N_573);
nand U2451 (N_2451,N_1547,In_4975);
nand U2452 (N_2452,N_335,In_2045);
nand U2453 (N_2453,In_1113,N_1467);
nand U2454 (N_2454,In_2020,N_355);
nor U2455 (N_2455,In_4952,N_1304);
nand U2456 (N_2456,In_2099,In_2382);
or U2457 (N_2457,N_1704,N_1559);
and U2458 (N_2458,N_780,In_3859);
nand U2459 (N_2459,N_1348,N_1497);
nand U2460 (N_2460,N_1215,N_1681);
nor U2461 (N_2461,In_3717,N_827);
nand U2462 (N_2462,In_1801,N_1771);
nand U2463 (N_2463,N_143,In_3435);
nand U2464 (N_2464,N_1696,N_1674);
and U2465 (N_2465,N_166,N_415);
nand U2466 (N_2466,In_722,N_376);
and U2467 (N_2467,In_4597,N_911);
nand U2468 (N_2468,N_1985,In_3773);
xor U2469 (N_2469,In_994,N_1513);
xor U2470 (N_2470,N_640,N_549);
or U2471 (N_2471,In_1018,N_1374);
nor U2472 (N_2472,In_1777,In_2556);
nand U2473 (N_2473,N_1911,In_903);
and U2474 (N_2474,N_1603,N_1043);
xnor U2475 (N_2475,N_1607,In_2301);
nor U2476 (N_2476,In_4299,In_4022);
xnor U2477 (N_2477,In_1914,In_608);
xor U2478 (N_2478,In_4858,In_1012);
and U2479 (N_2479,N_1959,In_1614);
nor U2480 (N_2480,N_1998,N_1150);
xnor U2481 (N_2481,In_4208,In_1359);
nand U2482 (N_2482,N_1813,N_740);
or U2483 (N_2483,N_1392,N_384);
or U2484 (N_2484,In_1313,In_4031);
or U2485 (N_2485,N_1106,In_3713);
nor U2486 (N_2486,In_1349,In_4064);
and U2487 (N_2487,N_578,N_1541);
xnor U2488 (N_2488,N_467,N_13);
nor U2489 (N_2489,N_585,In_150);
xnor U2490 (N_2490,N_116,N_705);
nand U2491 (N_2491,N_1520,In_4576);
xnor U2492 (N_2492,N_536,N_953);
nand U2493 (N_2493,N_892,N_1981);
nor U2494 (N_2494,N_304,In_4767);
nor U2495 (N_2495,N_492,N_955);
or U2496 (N_2496,N_1016,N_372);
nor U2497 (N_2497,N_1098,N_789);
and U2498 (N_2498,N_126,N_1721);
and U2499 (N_2499,N_1937,N_1514);
nor U2500 (N_2500,N_1849,N_131);
nand U2501 (N_2501,N_819,N_1279);
nor U2502 (N_2502,In_1149,N_769);
xnor U2503 (N_2503,N_299,In_3005);
nand U2504 (N_2504,In_3835,N_1228);
and U2505 (N_2505,N_439,N_957);
nand U2506 (N_2506,N_745,N_345);
nor U2507 (N_2507,N_941,N_674);
nand U2508 (N_2508,N_1085,N_219);
nor U2509 (N_2509,N_426,N_1977);
and U2510 (N_2510,N_1055,N_1060);
nor U2511 (N_2511,In_3634,In_2551);
nand U2512 (N_2512,N_238,N_1648);
nand U2513 (N_2513,N_1035,N_1087);
or U2514 (N_2514,N_1138,N_135);
and U2515 (N_2515,In_3996,N_1619);
nand U2516 (N_2516,N_140,N_1229);
nand U2517 (N_2517,N_1552,N_1722);
and U2518 (N_2518,N_91,N_910);
xnor U2519 (N_2519,N_264,In_3792);
and U2520 (N_2520,N_638,In_1287);
nand U2521 (N_2521,In_3797,In_1090);
nand U2522 (N_2522,In_257,N_1600);
nor U2523 (N_2523,In_3291,In_4721);
and U2524 (N_2524,N_1616,In_727);
xor U2525 (N_2525,In_2936,In_2595);
or U2526 (N_2526,In_3244,In_2125);
nor U2527 (N_2527,N_535,N_445);
nor U2528 (N_2528,N_538,N_802);
and U2529 (N_2529,In_3580,In_4257);
nand U2530 (N_2530,N_929,In_3362);
and U2531 (N_2531,In_829,In_1669);
nor U2532 (N_2532,N_1902,In_1543);
nand U2533 (N_2533,In_759,N_1589);
nor U2534 (N_2534,N_386,N_1837);
nor U2535 (N_2535,In_3608,N_1058);
nand U2536 (N_2536,In_4243,N_778);
nand U2537 (N_2537,In_2288,N_318);
and U2538 (N_2538,N_1332,N_1884);
or U2539 (N_2539,N_1356,N_1297);
nand U2540 (N_2540,N_334,N_652);
xor U2541 (N_2541,N_223,In_3025);
and U2542 (N_2542,N_1720,In_2646);
nand U2543 (N_2543,N_513,In_4781);
nand U2544 (N_2544,In_1928,N_122);
nor U2545 (N_2545,N_1640,N_1191);
xor U2546 (N_2546,N_1211,In_2594);
and U2547 (N_2547,In_4981,N_888);
nand U2548 (N_2548,N_1406,N_45);
nand U2549 (N_2549,In_1888,N_288);
xor U2550 (N_2550,N_868,In_3347);
nand U2551 (N_2551,N_1423,In_4983);
or U2552 (N_2552,In_1496,N_308);
nand U2553 (N_2553,N_317,In_2350);
xor U2554 (N_2554,In_1987,In_958);
xnor U2555 (N_2555,In_1140,In_2651);
nor U2556 (N_2556,N_452,N_366);
nor U2557 (N_2557,In_4828,In_2057);
xnor U2558 (N_2558,In_2085,N_1956);
or U2559 (N_2559,In_1635,In_1225);
xnor U2560 (N_2560,N_183,N_1895);
nand U2561 (N_2561,N_1251,N_1507);
xor U2562 (N_2562,N_109,N_1818);
nor U2563 (N_2563,N_1141,N_1736);
and U2564 (N_2564,In_392,In_4464);
xor U2565 (N_2565,In_627,In_3698);
nand U2566 (N_2566,N_448,In_2370);
and U2567 (N_2567,N_581,In_2362);
and U2568 (N_2568,N_1244,N_1537);
nand U2569 (N_2569,In_330,N_1548);
xor U2570 (N_2570,In_3204,In_4567);
and U2571 (N_2571,N_965,N_250);
nand U2572 (N_2572,N_706,N_1236);
and U2573 (N_2573,In_462,In_840);
xor U2574 (N_2574,In_3123,N_717);
or U2575 (N_2575,In_3896,N_298);
nand U2576 (N_2576,N_217,N_703);
nor U2577 (N_2577,N_743,In_776);
and U2578 (N_2578,N_1180,N_258);
nand U2579 (N_2579,N_1732,N_1457);
nand U2580 (N_2580,N_1416,N_1955);
and U2581 (N_2581,In_497,N_482);
and U2582 (N_2582,N_1562,N_945);
and U2583 (N_2583,N_1460,N_1339);
and U2584 (N_2584,N_1373,N_495);
or U2585 (N_2585,N_1426,N_66);
or U2586 (N_2586,N_512,In_4713);
xor U2587 (N_2587,In_4681,In_2917);
nor U2588 (N_2588,N_1281,N_1560);
nor U2589 (N_2589,N_1252,In_65);
xor U2590 (N_2590,N_102,N_1582);
nand U2591 (N_2591,N_1157,N_554);
and U2592 (N_2592,N_459,N_1650);
xnor U2593 (N_2593,N_1756,In_4077);
nor U2594 (N_2594,N_1105,In_4850);
xnor U2595 (N_2595,N_1330,In_4134);
or U2596 (N_2596,In_2030,N_1536);
nor U2597 (N_2597,N_67,N_1023);
and U2598 (N_2598,N_1757,In_4631);
and U2599 (N_2599,N_1504,In_867);
nand U2600 (N_2600,N_1833,In_2807);
and U2601 (N_2601,In_2598,N_294);
nand U2602 (N_2602,In_2719,N_1176);
xor U2603 (N_2603,N_94,N_1593);
nor U2604 (N_2604,N_1827,N_1679);
nor U2605 (N_2605,N_726,N_1832);
and U2606 (N_2606,N_808,N_832);
and U2607 (N_2607,In_265,N_632);
or U2608 (N_2608,N_1302,N_248);
nor U2609 (N_2609,N_828,In_3056);
nand U2610 (N_2610,N_280,In_3426);
nand U2611 (N_2611,N_1907,In_2826);
and U2612 (N_2612,In_4183,N_1201);
and U2613 (N_2613,N_499,In_4870);
and U2614 (N_2614,N_1802,N_26);
or U2615 (N_2615,N_688,N_1112);
nand U2616 (N_2616,N_77,In_3573);
or U2617 (N_2617,In_4240,N_1192);
xor U2618 (N_2618,N_971,N_687);
nand U2619 (N_2619,N_146,N_1478);
nor U2620 (N_2620,In_3965,N_1857);
or U2621 (N_2621,In_1970,N_1342);
nand U2622 (N_2622,N_746,N_834);
nor U2623 (N_2623,N_1433,In_2381);
xnor U2624 (N_2624,N_1609,N_1512);
nor U2625 (N_2625,In_3677,N_636);
and U2626 (N_2626,N_1100,N_557);
nor U2627 (N_2627,N_145,In_4595);
and U2628 (N_2628,In_4635,N_727);
nand U2629 (N_2629,N_1983,N_693);
and U2630 (N_2630,N_664,N_1217);
and U2631 (N_2631,N_909,N_1797);
or U2632 (N_2632,N_1516,N_68);
and U2633 (N_2633,In_1009,N_1142);
xnor U2634 (N_2634,In_3444,N_1783);
nor U2635 (N_2635,N_1786,N_1750);
xor U2636 (N_2636,N_658,N_438);
nor U2637 (N_2637,In_3400,N_1284);
and U2638 (N_2638,In_3481,In_2834);
and U2639 (N_2639,In_3707,In_4438);
nand U2640 (N_2640,N_1041,In_2055);
xnor U2641 (N_2641,N_1178,N_103);
and U2642 (N_2642,In_4727,In_4491);
or U2643 (N_2643,N_168,N_296);
nand U2644 (N_2644,N_1341,In_1900);
and U2645 (N_2645,In_2073,In_1229);
or U2646 (N_2646,N_508,N_346);
nor U2647 (N_2647,N_881,N_1601);
xnor U2648 (N_2648,In_2437,N_501);
nor U2649 (N_2649,In_616,N_922);
and U2650 (N_2650,N_1949,N_58);
xor U2651 (N_2651,N_263,N_1031);
and U2652 (N_2652,N_670,In_1768);
nand U2653 (N_2653,N_982,N_961);
or U2654 (N_2654,N_1639,In_68);
nand U2655 (N_2655,In_3495,In_3868);
xnor U2656 (N_2656,N_1604,N_1843);
xor U2657 (N_2657,In_3564,In_402);
xnor U2658 (N_2658,N_1046,In_1885);
or U2659 (N_2659,N_1143,N_950);
xnor U2660 (N_2660,N_807,In_4391);
or U2661 (N_2661,N_1220,N_1326);
and U2662 (N_2662,In_2238,N_1699);
nand U2663 (N_2663,N_121,N_466);
and U2664 (N_2664,N_1588,N_129);
or U2665 (N_2665,N_1350,N_1769);
or U2666 (N_2666,N_1511,In_3602);
or U2667 (N_2667,N_1310,N_1693);
xnor U2668 (N_2668,N_1422,N_119);
or U2669 (N_2669,In_259,N_1524);
xor U2670 (N_2670,N_1364,N_1557);
nor U2671 (N_2671,N_195,N_305);
xnor U2672 (N_2672,In_2271,In_3552);
xnor U2673 (N_2673,In_1909,N_1663);
nor U2674 (N_2674,N_465,N_1102);
or U2675 (N_2675,N_925,N_978);
nor U2676 (N_2676,N_289,N_1453);
or U2677 (N_2677,In_4564,In_1640);
xor U2678 (N_2678,In_189,N_5);
nand U2679 (N_2679,In_1074,N_1441);
nand U2680 (N_2680,N_1014,N_267);
and U2681 (N_2681,N_1490,In_3364);
and U2682 (N_2682,N_1865,In_3977);
nor U2683 (N_2683,N_1551,N_924);
nand U2684 (N_2684,In_856,In_4699);
xor U2685 (N_2685,N_1296,N_410);
nand U2686 (N_2686,In_2109,N_1492);
and U2687 (N_2687,In_2971,N_1412);
nand U2688 (N_2688,In_230,N_38);
and U2689 (N_2689,N_1381,N_1227);
or U2690 (N_2690,N_1024,N_1166);
or U2691 (N_2691,N_1543,In_4285);
and U2692 (N_2692,N_637,N_534);
nand U2693 (N_2693,In_145,N_1856);
nand U2694 (N_2694,In_4505,In_4005);
nand U2695 (N_2695,In_3099,In_3816);
or U2696 (N_2696,N_347,N_1401);
nor U2697 (N_2697,In_2819,N_265);
nand U2698 (N_2698,In_570,N_1906);
nor U2699 (N_2699,N_1443,N_1565);
xnor U2700 (N_2700,N_127,In_3585);
nand U2701 (N_2701,In_4280,In_609);
xor U2702 (N_2702,N_1765,N_1563);
and U2703 (N_2703,In_4687,N_537);
xnor U2704 (N_2704,N_654,N_312);
xnor U2705 (N_2705,N_474,N_1427);
nor U2706 (N_2706,N_253,In_4049);
and U2707 (N_2707,In_4998,N_1745);
and U2708 (N_2708,N_570,In_1696);
or U2709 (N_2709,N_1599,In_3758);
xor U2710 (N_2710,N_1414,N_1019);
xor U2711 (N_2711,N_1659,N_277);
xor U2712 (N_2712,N_506,In_3785);
or U2713 (N_2713,In_2911,N_449);
nor U2714 (N_2714,N_54,N_417);
nor U2715 (N_2715,N_934,N_1474);
nand U2716 (N_2716,In_1038,In_2825);
nand U2717 (N_2717,N_983,N_1469);
nand U2718 (N_2718,N_365,N_1632);
nand U2719 (N_2719,N_30,N_192);
nor U2720 (N_2720,In_4669,In_1711);
xnor U2721 (N_2721,N_464,In_4544);
xor U2722 (N_2722,In_1753,N_1107);
nand U2723 (N_2723,N_1908,N_489);
or U2724 (N_2724,In_2495,N_1054);
or U2725 (N_2725,In_4223,N_369);
nand U2726 (N_2726,In_664,N_172);
xor U2727 (N_2727,In_3731,N_1352);
nand U2728 (N_2728,N_1701,N_53);
or U2729 (N_2729,N_1384,N_643);
nor U2730 (N_2730,N_1189,N_214);
and U2731 (N_2731,N_359,N_754);
nor U2732 (N_2732,N_156,N_1726);
or U2733 (N_2733,N_1161,N_491);
and U2734 (N_2734,N_916,In_807);
nor U2735 (N_2735,N_648,N_1661);
and U2736 (N_2736,N_1862,N_900);
nor U2737 (N_2737,In_699,N_187);
and U2738 (N_2738,N_1120,N_433);
xor U2739 (N_2739,N_1367,N_1493);
and U2740 (N_2740,In_955,N_1746);
or U2741 (N_2741,N_623,N_682);
xor U2742 (N_2742,N_1238,N_1418);
or U2743 (N_2743,N_647,N_756);
or U2744 (N_2744,In_296,N_1393);
or U2745 (N_2745,In_1030,In_4411);
or U2746 (N_2746,N_142,N_247);
xnor U2747 (N_2747,In_4136,In_4743);
and U2748 (N_2748,N_380,N_1530);
and U2749 (N_2749,In_251,N_1874);
nand U2750 (N_2750,N_101,N_1733);
nor U2751 (N_2751,N_191,N_377);
xnor U2752 (N_2752,In_4652,N_1775);
xnor U2753 (N_2753,N_1465,N_1044);
and U2754 (N_2754,N_659,N_1785);
or U2755 (N_2755,In_132,N_1318);
nor U2756 (N_2756,N_870,N_1485);
xor U2757 (N_2757,N_351,In_3541);
nand U2758 (N_2758,N_631,In_17);
or U2759 (N_2759,In_1209,In_1895);
or U2760 (N_2760,N_976,In_1664);
and U2761 (N_2761,N_772,N_1816);
and U2762 (N_2762,In_691,N_1836);
and U2763 (N_2763,N_24,In_1680);
and U2764 (N_2764,N_755,In_4474);
xor U2765 (N_2765,N_923,N_89);
and U2766 (N_2766,N_1305,N_29);
xnor U2767 (N_2767,N_1627,N_1285);
nand U2768 (N_2768,N_1815,In_26);
nor U2769 (N_2769,In_2741,N_1919);
xor U2770 (N_2770,N_1451,In_2406);
and U2771 (N_2771,N_269,N_1377);
nor U2772 (N_2772,In_2294,In_1654);
xor U2773 (N_2773,N_1108,N_1172);
and U2774 (N_2774,N_62,N_1029);
nor U2775 (N_2775,In_498,N_937);
or U2776 (N_2776,In_640,N_1345);
xnor U2777 (N_2777,N_1930,In_360);
and U2778 (N_2778,In_1867,N_87);
or U2779 (N_2779,N_1079,N_1567);
and U2780 (N_2780,N_1554,N_39);
xor U2781 (N_2781,N_739,N_1188);
nand U2782 (N_2782,N_475,N_1576);
or U2783 (N_2783,In_1396,N_992);
nor U2784 (N_2784,N_330,N_1159);
xnor U2785 (N_2785,N_1590,N_1634);
nor U2786 (N_2786,In_2601,In_1522);
xor U2787 (N_2787,In_2100,N_548);
and U2788 (N_2788,N_1061,N_1383);
or U2789 (N_2789,N_609,N_539);
nand U2790 (N_2790,N_1863,N_357);
nor U2791 (N_2791,N_902,N_1751);
xor U2792 (N_2792,N_944,N_784);
nand U2793 (N_2793,N_1408,N_398);
and U2794 (N_2794,N_1870,N_399);
and U2795 (N_2795,In_4454,In_1339);
nor U2796 (N_2796,N_1210,In_2415);
xor U2797 (N_2797,N_1397,N_1743);
nand U2798 (N_2798,In_4386,N_1788);
xnor U2799 (N_2799,N_1365,In_3);
or U2800 (N_2800,In_3046,N_698);
and U2801 (N_2801,N_391,In_4746);
nor U2802 (N_2802,N_1206,N_447);
nor U2803 (N_2803,N_1199,In_4253);
nand U2804 (N_2804,N_1049,N_785);
xor U2805 (N_2805,N_1658,N_665);
xor U2806 (N_2806,In_4697,In_864);
xnor U2807 (N_2807,N_565,N_1517);
and U2808 (N_2808,N_980,N_1621);
xnor U2809 (N_2809,In_1589,N_1325);
nor U2810 (N_2810,In_4549,N_1415);
nand U2811 (N_2811,In_644,N_1265);
xor U2812 (N_2812,In_3088,In_2128);
or U2813 (N_2813,N_1974,N_1894);
and U2814 (N_2814,N_1767,In_1283);
and U2815 (N_2815,In_1092,In_1560);
nor U2816 (N_2816,N_531,N_1958);
and U2817 (N_2817,In_2804,In_3517);
nor U2818 (N_2818,N_1811,N_702);
and U2819 (N_2819,N_1347,N_1657);
nor U2820 (N_2820,N_1678,In_281);
xor U2821 (N_2821,N_974,N_215);
or U2822 (N_2822,N_993,N_760);
nor U2823 (N_2823,N_1313,N_885);
xnor U2824 (N_2824,In_2095,N_878);
nor U2825 (N_2825,N_1677,N_1328);
and U2826 (N_2826,In_1701,In_4664);
nor U2827 (N_2827,In_2653,N_1446);
nand U2828 (N_2828,In_3196,In_822);
or U2829 (N_2829,N_646,N_1866);
and U2830 (N_2830,N_1909,In_4843);
nand U2831 (N_2831,N_767,N_1213);
nor U2832 (N_2832,N_813,N_1103);
nand U2833 (N_2833,N_1893,In_980);
nor U2834 (N_2834,N_709,N_395);
or U2835 (N_2835,N_1595,N_155);
nand U2836 (N_2836,In_2469,In_4334);
or U2837 (N_2837,N_1807,N_562);
nor U2838 (N_2838,N_1394,In_1293);
nand U2839 (N_2839,N_1828,In_4536);
and U2840 (N_2840,N_434,N_1036);
nor U2841 (N_2841,N_889,In_3250);
xnor U2842 (N_2842,N_311,In_2703);
nand U2843 (N_2843,N_792,N_737);
or U2844 (N_2844,N_228,N_1494);
nor U2845 (N_2845,In_3574,N_138);
xnor U2846 (N_2846,N_1066,N_1855);
nor U2847 (N_2847,N_856,N_1280);
or U2848 (N_2848,N_1185,N_1196);
nand U2849 (N_2849,In_2666,N_235);
nand U2850 (N_2850,In_4156,N_1258);
xor U2851 (N_2851,N_105,N_1829);
xor U2852 (N_2852,In_697,N_28);
and U2853 (N_2853,N_354,In_57);
and U2854 (N_2854,N_1707,N_914);
nand U2855 (N_2855,In_3605,N_516);
nand U2856 (N_2856,In_2293,N_750);
and U2857 (N_2857,N_582,N_1385);
and U2858 (N_2858,N_1725,N_1646);
and U2859 (N_2859,N_278,In_2841);
xor U2860 (N_2860,In_3483,N_339);
and U2861 (N_2861,In_2211,In_3623);
xor U2862 (N_2862,In_1097,In_3327);
and U2863 (N_2863,N_158,N_811);
xor U2864 (N_2864,N_684,N_3);
and U2865 (N_2865,N_587,N_666);
and U2866 (N_2866,N_1748,N_543);
or U2867 (N_2867,In_85,N_1729);
nand U2868 (N_2868,N_1889,In_2644);
or U2869 (N_2869,In_3874,In_2962);
or U2870 (N_2870,In_1197,N_759);
nand U2871 (N_2871,In_2258,N_327);
nand U2872 (N_2872,In_757,In_4171);
xor U2873 (N_2873,N_1093,In_483);
nand U2874 (N_2874,N_586,In_1906);
xnor U2875 (N_2875,N_1034,N_657);
nor U2876 (N_2876,N_1067,In_1920);
nand U2877 (N_2877,N_148,In_2790);
xor U2878 (N_2878,N_388,In_4403);
xor U2879 (N_2879,In_1720,In_3024);
nand U2880 (N_2880,N_766,N_771);
nand U2881 (N_2881,N_1239,In_597);
nand U2882 (N_2882,N_457,In_2374);
or U2883 (N_2883,N_1804,In_427);
xor U2884 (N_2884,N_1875,N_873);
nor U2885 (N_2885,N_1094,In_4190);
nand U2886 (N_2886,In_4217,N_1770);
nand U2887 (N_2887,In_1658,N_1939);
and U2888 (N_2888,In_4990,N_470);
and U2889 (N_2889,N_336,In_636);
nor U2890 (N_2890,In_3253,N_1910);
nor U2891 (N_2891,N_1791,In_4499);
or U2892 (N_2892,N_1027,N_1605);
nor U2893 (N_2893,N_1835,In_1356);
xnor U2894 (N_2894,N_1842,N_1954);
or U2895 (N_2895,N_210,N_134);
and U2896 (N_2896,N_1331,N_847);
xor U2897 (N_2897,N_1561,In_4745);
nand U2898 (N_2898,N_1291,N_1995);
nand U2899 (N_2899,N_348,In_2280);
xor U2900 (N_2900,N_61,In_3387);
xor U2901 (N_2901,N_1234,In_3995);
xnor U2902 (N_2902,In_3107,N_1175);
xor U2903 (N_2903,N_775,N_1585);
or U2904 (N_2904,N_123,N_517);
or U2905 (N_2905,N_1834,N_815);
and U2906 (N_2906,In_4915,N_614);
nand U2907 (N_2907,In_109,In_1441);
nand U2908 (N_2908,In_2838,N_1782);
nand U2909 (N_2909,N_381,In_1979);
nor U2910 (N_2910,N_1396,N_1506);
xnor U2911 (N_2911,N_1888,N_1135);
xor U2912 (N_2912,N_1762,N_1425);
nor U2913 (N_2913,In_4803,N_1787);
nand U2914 (N_2914,N_260,In_4926);
or U2915 (N_2915,N_1656,N_463);
nor U2916 (N_2916,N_1095,In_1151);
or U2917 (N_2917,N_1378,N_504);
or U2918 (N_2918,N_1876,In_3137);
nor U2919 (N_2919,N_1924,N_1629);
nor U2920 (N_2920,In_2232,N_1306);
nor U2921 (N_2921,N_261,N_1929);
xor U2922 (N_2922,N_1410,N_222);
nand U2923 (N_2923,N_42,N_1197);
and U2924 (N_2924,N_893,N_1738);
nand U2925 (N_2925,N_1867,In_3519);
nand U2926 (N_2926,In_2669,In_1896);
xor U2927 (N_2927,N_1879,In_1976);
nand U2928 (N_2928,In_802,In_2268);
nor U2929 (N_2929,In_1994,N_451);
nand U2930 (N_2930,N_1089,N_268);
xor U2931 (N_2931,N_1913,In_2515);
xnor U2932 (N_2932,N_412,In_3780);
nor U2933 (N_2933,In_610,N_1882);
xor U2934 (N_2934,In_4756,N_1683);
nor U2935 (N_2935,N_1168,N_782);
nand U2936 (N_2936,N_1071,N_340);
nand U2937 (N_2937,N_1092,N_1283);
or U2938 (N_2938,In_4061,In_2728);
and U2939 (N_2939,In_2650,N_1151);
or U2940 (N_2940,In_4214,N_1287);
nor U2941 (N_2941,In_720,N_188);
nand U2942 (N_2942,N_110,N_1673);
and U2943 (N_2943,N_960,N_530);
and U2944 (N_2944,N_1694,In_2796);
xor U2945 (N_2945,N_368,In_4560);
or U2946 (N_2946,N_315,N_373);
and U2947 (N_2947,In_1136,N_382);
and U2948 (N_2948,N_713,N_675);
or U2949 (N_2949,N_1181,N_270);
or U2950 (N_2950,In_4154,In_3297);
or U2951 (N_2951,N_1275,In_1458);
xor U2952 (N_2952,N_367,N_849);
and U2953 (N_2953,In_2407,N_360);
or U2954 (N_2954,N_1123,N_959);
or U2955 (N_2955,In_1794,In_2736);
nor U2956 (N_2956,N_686,N_1273);
nor U2957 (N_2957,N_1253,In_3261);
xnor U2958 (N_2958,N_1793,In_3404);
nor U2959 (N_2959,In_2359,N_200);
nor U2960 (N_2960,N_1075,N_628);
xor U2961 (N_2961,N_63,In_1601);
nand U2962 (N_2962,In_2052,In_2267);
nand U2963 (N_2963,N_1052,N_387);
xor U2964 (N_2964,In_3720,N_313);
or U2965 (N_2965,N_1851,N_10);
or U2966 (N_2966,N_1177,In_1733);
nor U2967 (N_2967,In_2036,N_527);
nor U2968 (N_2968,N_1747,N_1231);
nand U2969 (N_2969,N_173,N_515);
nor U2970 (N_2970,N_1466,N_361);
xnor U2971 (N_2971,N_901,N_128);
and U2972 (N_2972,N_1472,N_1147);
or U2973 (N_2973,N_809,In_97);
nor U2974 (N_2974,In_593,In_309);
xor U2975 (N_2975,In_546,N_51);
nand U2976 (N_2976,In_2265,N_1830);
nand U2977 (N_2977,N_1730,N_1550);
xor U2978 (N_2978,In_2968,N_1969);
and U2979 (N_2979,In_3329,N_1925);
nand U2980 (N_2980,In_4067,N_1083);
xnor U2981 (N_2981,N_6,N_1903);
xor U2982 (N_2982,In_2888,N_353);
xor U2983 (N_2983,N_619,In_362);
and U2984 (N_2984,N_36,N_806);
and U2985 (N_2985,N_1724,N_167);
and U2986 (N_2986,N_1282,N_825);
nand U2987 (N_2987,In_2923,N_93);
and U2988 (N_2988,N_991,N_1950);
xor U2989 (N_2989,N_230,In_574);
or U2990 (N_2990,In_2226,In_4111);
xnor U2991 (N_2991,N_1987,N_1084);
or U2992 (N_2992,N_19,N_1476);
and U2993 (N_2993,In_4439,N_1303);
nor U2994 (N_2994,N_332,In_2146);
xor U2995 (N_2995,N_1814,N_749);
xor U2996 (N_2996,In_2663,N_1636);
xor U2997 (N_2997,N_673,N_589);
or U2998 (N_2998,In_1120,N_1806);
and U2999 (N_2999,N_1716,N_1591);
or U3000 (N_3000,N_137,N_435);
xor U3001 (N_3001,N_896,N_1026);
nand U3002 (N_3002,N_964,N_1946);
or U3003 (N_3003,N_1407,In_1617);
xnor U3004 (N_3004,N_798,N_718);
nor U3005 (N_3005,N_1372,In_1165);
nor U3006 (N_3006,N_553,N_2);
nor U3007 (N_3007,N_212,N_1420);
nand U3008 (N_3008,N_1962,N_1753);
nand U3009 (N_3009,In_1274,In_1789);
or U3010 (N_3010,N_904,N_1390);
nor U3011 (N_3011,N_1670,N_73);
and U3012 (N_3012,In_1613,N_1626);
nor U3013 (N_3013,In_2854,N_401);
or U3014 (N_3014,N_1208,N_699);
nand U3015 (N_3015,In_4725,In_3853);
and U3016 (N_3016,In_4813,N_1847);
xnor U3017 (N_3017,N_224,N_113);
nor U3018 (N_3018,In_245,In_2411);
nand U3019 (N_3019,N_979,N_1260);
xor U3020 (N_3020,N_803,N_1951);
nand U3021 (N_3021,N_319,In_4417);
xor U3022 (N_3022,In_103,N_741);
or U3023 (N_3023,N_728,N_139);
or U3024 (N_3024,N_777,In_3722);
xor U3025 (N_3025,N_774,N_1933);
and U3026 (N_3026,In_3293,N_1990);
xor U3027 (N_3027,In_3922,N_50);
nand U3028 (N_3028,In_4139,In_3967);
and U3029 (N_3029,N_1137,In_650);
or U3030 (N_3030,N_271,In_886);
xnor U3031 (N_3031,In_131,In_3735);
nand U3032 (N_3032,N_1127,In_3983);
or U3033 (N_3033,N_1447,N_667);
and U3034 (N_3034,N_855,In_4857);
nand U3035 (N_3035,N_1799,N_1723);
nor U3036 (N_3036,N_890,In_3655);
nand U3037 (N_3037,N_1419,N_494);
and U3038 (N_3038,N_1976,In_3918);
and U3039 (N_3039,N_184,In_4941);
xnor U3040 (N_3040,N_651,In_3377);
or U3041 (N_3041,In_1629,N_233);
and U3042 (N_3042,In_1139,In_4018);
or U3043 (N_3043,N_1558,In_1891);
nor U3044 (N_3044,In_121,N_1838);
nand U3045 (N_3045,N_680,N_1232);
nand U3046 (N_3046,N_1873,N_115);
nand U3047 (N_3047,N_1625,In_3372);
and U3048 (N_3048,N_400,N_300);
and U3049 (N_3049,In_1907,In_22);
xnor U3050 (N_3050,In_2296,N_497);
xnor U3051 (N_3051,In_3508,N_1013);
xor U3052 (N_3052,In_365,N_1654);
nand U3053 (N_3053,N_711,In_4521);
and U3054 (N_3054,N_621,N_1337);
and U3055 (N_3055,N_52,In_1525);
nand U3056 (N_3056,In_1809,N_604);
and U3057 (N_3057,N_342,N_324);
and U3058 (N_3058,N_197,In_4443);
and U3059 (N_3059,In_1176,In_890);
or U3060 (N_3060,N_82,N_343);
and U3061 (N_3061,In_2311,N_567);
xor U3062 (N_3062,N_1140,In_1203);
nand U3063 (N_3063,In_1089,N_939);
or U3064 (N_3064,In_2475,N_100);
or U3065 (N_3065,N_84,N_996);
nand U3066 (N_3066,In_3120,N_783);
xor U3067 (N_3067,N_546,N_1300);
nand U3068 (N_3068,In_4328,N_404);
nor U3069 (N_3069,N_935,In_3130);
nor U3070 (N_3070,In_2555,N_1221);
or U3071 (N_3071,In_2868,In_2227);
and U3072 (N_3072,N_921,N_362);
nor U3073 (N_3073,N_33,In_1725);
and U3074 (N_3074,N_236,N_644);
nand U3075 (N_3075,N_1682,In_1898);
or U3076 (N_3076,N_1461,N_47);
nor U3077 (N_3077,In_723,In_1765);
and U3078 (N_3078,N_1202,N_1689);
xnor U3079 (N_3079,N_611,N_1464);
or U3080 (N_3080,N_1556,N_1698);
or U3081 (N_3081,N_1417,N_1620);
or U3082 (N_3082,In_4606,In_4538);
xnor U3083 (N_3083,N_1598,In_595);
nand U3084 (N_3084,N_1050,In_4729);
xnor U3085 (N_3085,N_677,N_1614);
or U3086 (N_3086,N_898,N_816);
xnor U3087 (N_3087,N_1148,N_56);
or U3088 (N_3088,N_213,N_990);
nor U3089 (N_3089,N_114,N_1333);
xor U3090 (N_3090,N_1387,In_4973);
and U3091 (N_3091,In_843,N_1688);
and U3092 (N_3092,In_2318,In_3650);
nor U3093 (N_3093,N_259,N_1921);
or U3094 (N_3094,In_1415,N_454);
nand U3095 (N_3095,N_532,N_528);
xor U3096 (N_3096,N_225,In_981);
xor U3097 (N_3097,In_3601,N_256);
xor U3098 (N_3098,N_1784,N_899);
or U3099 (N_3099,N_618,In_4406);
xor U3100 (N_3100,In_1892,N_1136);
and U3101 (N_3101,N_446,N_1850);
nor U3102 (N_3102,In_434,N_1267);
xnor U3103 (N_3103,N_450,N_78);
nand U3104 (N_3104,N_1179,In_2277);
nand U3105 (N_3105,N_162,N_625);
nor U3106 (N_3106,In_2491,N_597);
and U3107 (N_3107,N_584,In_3206);
or U3108 (N_3108,N_742,N_1798);
or U3109 (N_3109,In_2225,In_3216);
nor U3110 (N_3110,N_458,In_3898);
nor U3111 (N_3111,In_81,N_956);
nor U3112 (N_3112,N_11,In_460);
and U3113 (N_3113,In_517,N_738);
and U3114 (N_3114,N_69,In_3438);
and U3115 (N_3115,N_1628,N_1115);
nor U3116 (N_3116,N_1096,In_1261);
nor U3117 (N_3117,N_1173,In_475);
xor U3118 (N_3118,N_1664,N_1805);
nand U3119 (N_3119,In_3678,N_987);
and U3120 (N_3120,N_1480,N_1111);
nor U3121 (N_3121,N_639,In_4370);
or U3122 (N_3122,N_1622,N_1710);
or U3123 (N_3123,In_342,In_911);
or U3124 (N_3124,In_1591,N_227);
nand U3125 (N_3125,N_1351,N_1831);
and U3126 (N_3126,In_3381,In_4479);
or U3127 (N_3127,N_969,N_92);
or U3128 (N_3128,N_375,N_846);
or U3129 (N_3129,N_1077,N_60);
nand U3130 (N_3130,N_797,N_358);
nor U3131 (N_3131,N_104,N_41);
xnor U3132 (N_3132,N_551,N_626);
nor U3133 (N_3133,N_634,N_561);
nor U3134 (N_3134,N_1608,N_1852);
and U3135 (N_3135,N_511,In_3363);
nand U3136 (N_3136,N_493,N_1534);
xnor U3137 (N_3137,In_1838,In_278);
xnor U3138 (N_3138,N_208,In_1105);
xnor U3139 (N_3139,N_1270,N_1569);
nor U3140 (N_3140,N_1207,In_3858);
xnor U3141 (N_3141,In_3159,N_290);
nand U3142 (N_3142,N_1780,N_1255);
nand U3143 (N_3143,N_905,In_331);
nor U3144 (N_3144,N_487,N_786);
nand U3145 (N_3145,N_441,In_1488);
or U3146 (N_3146,N_1713,N_456);
xor U3147 (N_3147,N_635,In_3824);
nand U3148 (N_3148,In_1567,N_490);
and U3149 (N_3149,N_1268,N_337);
xor U3150 (N_3150,N_239,In_936);
nand U3151 (N_3151,N_14,In_2866);
nand U3152 (N_3152,N_1174,N_874);
nand U3153 (N_3153,N_1376,N_1445);
or U3154 (N_3154,N_427,N_1254);
and U3155 (N_3155,N_1868,N_1502);
nand U3156 (N_3156,N_163,N_973);
xor U3157 (N_3157,N_1329,N_694);
or U3158 (N_3158,In_286,In_1058);
or U3159 (N_3159,N_1069,N_254);
nand U3160 (N_3160,N_1978,N_1334);
nand U3161 (N_3161,N_931,In_1657);
or U3162 (N_3162,In_177,In_3604);
nor U3163 (N_3163,N_95,In_4624);
xor U3164 (N_3164,In_573,N_1380);
nand U3165 (N_3165,N_1581,N_1109);
nand U3166 (N_3166,N_1984,N_823);
and U3167 (N_3167,N_563,N_884);
nand U3168 (N_3168,N_765,In_708);
nor U3169 (N_3169,N_1463,In_4178);
xor U3170 (N_3170,N_866,In_1709);
or U3171 (N_3171,In_401,N_861);
nand U3172 (N_3172,In_4594,N_1499);
and U3173 (N_3173,N_649,N_1344);
or U3174 (N_3174,N_1368,N_1735);
xnor U3175 (N_3175,In_900,In_1716);
nor U3176 (N_3176,N_1587,In_1990);
nor U3177 (N_3177,N_915,In_1554);
or U3178 (N_3178,In_4145,In_2453);
or U3179 (N_3179,In_3649,N_606);
nor U3180 (N_3180,N_1881,N_1672);
nor U3181 (N_3181,N_57,In_2499);
nand U3182 (N_3182,In_2871,N_1905);
and U3183 (N_3183,N_1431,N_1395);
xnor U3184 (N_3184,In_3152,In_217);
nand U3185 (N_3185,N_1475,N_721);
and U3186 (N_3186,N_326,N_1878);
nand U3187 (N_3187,N_1690,N_1912);
xor U3188 (N_3188,N_1311,N_630);
nand U3189 (N_3189,N_947,In_2687);
nand U3190 (N_3190,N_1931,N_1439);
nand U3191 (N_3191,In_577,In_3886);
or U3192 (N_3192,N_408,N_9);
or U3193 (N_3193,N_453,N_770);
or U3194 (N_3194,N_1986,In_479);
nand U3195 (N_3195,N_1826,In_946);
nor U3196 (N_3196,In_2502,N_341);
xnor U3197 (N_3197,N_663,In_149);
nand U3198 (N_3198,N_1119,N_886);
nand U3199 (N_3199,N_897,N_758);
nor U3200 (N_3200,N_1190,N_1240);
and U3201 (N_3201,N_276,N_396);
xnor U3202 (N_3202,In_3834,N_1503);
and U3203 (N_3203,N_1468,In_1851);
or U3204 (N_3204,N_1667,N_1501);
xor U3205 (N_3205,N_406,In_3733);
xor U3206 (N_3206,In_1258,N_1928);
or U3207 (N_3207,N_1994,N_936);
and U3208 (N_3208,In_1326,In_621);
xor U3209 (N_3209,N_593,N_970);
or U3210 (N_3210,N_27,In_3294);
and U3211 (N_3211,N_1886,N_1153);
nand U3212 (N_3212,In_2462,N_1126);
and U3213 (N_3213,N_1086,In_2298);
nor U3214 (N_3214,In_1500,N_940);
xnor U3215 (N_3215,In_1045,N_701);
xor U3216 (N_3216,In_712,N_821);
nor U3217 (N_3217,N_685,N_1631);
nor U3218 (N_3218,In_4314,N_1286);
or U3219 (N_3219,N_963,N_1294);
nor U3220 (N_3220,N_523,N_579);
nor U3221 (N_3221,N_1535,N_301);
xnor U3222 (N_3222,N_1278,N_595);
or U3223 (N_3223,N_477,In_578);
and U3224 (N_3224,N_814,In_962);
nor U3225 (N_3225,In_2114,N_1158);
nor U3226 (N_3226,N_776,N_716);
or U3227 (N_3227,N_997,N_1134);
or U3228 (N_3228,N_1915,N_645);
and U3229 (N_3229,In_406,N_133);
or U3230 (N_3230,In_1790,N_1222);
or U3231 (N_3231,N_1897,N_244);
nor U3232 (N_3232,In_1153,In_3907);
or U3233 (N_3233,N_473,In_3814);
nor U3234 (N_3234,In_2377,N_281);
and U3235 (N_3235,In_853,N_552);
nor U3236 (N_3236,In_2214,N_1006);
xor U3237 (N_3237,N_1555,In_4251);
xor U3238 (N_3238,N_696,N_1080);
xor U3239 (N_3239,N_1768,N_164);
xor U3240 (N_3240,N_402,N_690);
nand U3241 (N_3241,In_1793,N_169);
nor U3242 (N_3242,In_1816,N_880);
or U3243 (N_3243,N_607,N_1668);
and U3244 (N_3244,N_310,In_4543);
and U3245 (N_3245,N_16,N_708);
nand U3246 (N_3246,N_612,In_3888);
or U3247 (N_3247,N_405,In_3192);
and U3248 (N_3248,N_1936,N_1509);
or U3249 (N_3249,N_1167,In_1524);
or U3250 (N_3250,In_2102,N_653);
and U3251 (N_3251,N_1714,N_1638);
xor U3252 (N_3252,In_2751,N_221);
nor U3253 (N_3253,N_303,In_482);
and U3254 (N_3254,In_2315,N_1473);
and U3255 (N_3255,N_1256,In_2865);
xnor U3256 (N_3256,In_2924,N_397);
and U3257 (N_3257,N_211,N_1235);
xnor U3258 (N_3258,N_1152,N_444);
nand U3259 (N_3259,In_99,In_4249);
xor U3260 (N_3260,N_385,In_3355);
nand U3261 (N_3261,N_1660,N_328);
and U3262 (N_3262,In_1172,N_1943);
or U3263 (N_3263,N_59,N_1508);
nand U3264 (N_3264,N_1437,N_178);
or U3265 (N_3265,N_179,N_1321);
xnor U3266 (N_3266,N_845,N_555);
nand U3267 (N_3267,N_526,N_1612);
or U3268 (N_3268,In_3265,N_1389);
xnor U3269 (N_3269,In_701,N_695);
nor U3270 (N_3270,In_3509,N_1744);
and U3271 (N_3271,N_479,N_999);
or U3272 (N_3272,In_651,N_692);
xor U3273 (N_3273,N_1592,N_252);
or U3274 (N_3274,In_1910,N_1839);
or U3275 (N_3275,N_190,N_1615);
nand U3276 (N_3276,N_1400,In_4554);
nand U3277 (N_3277,N_44,In_4046);
nand U3278 (N_3278,N_572,In_4899);
xor U3279 (N_3279,N_1692,In_2629);
and U3280 (N_3280,N_1203,In_2478);
or U3281 (N_3281,In_349,N_112);
xor U3282 (N_3282,N_1409,N_40);
nand U3283 (N_3283,N_1637,N_440);
nand U3284 (N_3284,N_853,N_1169);
xnor U3285 (N_3285,In_199,In_4255);
nor U3286 (N_3286,N_1261,In_3227);
xor U3287 (N_3287,N_468,N_720);
nor U3288 (N_3288,In_2981,N_32);
or U3289 (N_3289,In_2205,N_1891);
nand U3290 (N_3290,N_1459,N_111);
or U3291 (N_3291,N_518,In_187);
xor U3292 (N_3292,In_1494,In_282);
or U3293 (N_3293,N_1997,N_599);
or U3294 (N_3294,In_4728,N_1250);
nand U3295 (N_3295,N_1947,In_3875);
nor U3296 (N_3296,In_343,In_1344);
and U3297 (N_3297,In_1843,In_2006);
and U3298 (N_3298,N_1428,N_1230);
nor U3299 (N_3299,In_4327,N_1578);
nor U3300 (N_3300,In_3562,N_8);
nor U3301 (N_3301,In_912,N_1871);
or U3302 (N_3302,N_793,N_1777);
and U3303 (N_3303,N_471,N_1531);
or U3304 (N_3304,In_326,N_79);
and U3305 (N_3305,In_3140,N_186);
and U3306 (N_3306,In_2797,In_373);
nor U3307 (N_3307,N_1916,N_437);
or U3308 (N_3308,N_751,In_1353);
xor U3309 (N_3309,N_1355,N_733);
xnor U3310 (N_3310,In_2253,In_1710);
or U3311 (N_3311,N_1025,N_559);
nor U3312 (N_3312,N_1038,In_4884);
xnor U3313 (N_3313,In_1700,N_1299);
nor U3314 (N_3314,N_679,In_3584);
and U3315 (N_3315,N_672,N_1434);
or U3316 (N_3316,In_4284,N_130);
and U3317 (N_3317,In_858,N_1819);
xnor U3318 (N_3318,N_1359,In_3748);
nor U3319 (N_3319,N_1846,In_4414);
and U3320 (N_3320,In_2123,N_153);
xnor U3321 (N_3321,In_3129,N_1145);
xor U3322 (N_3322,N_4,N_930);
nor U3323 (N_3323,N_1941,In_4563);
and U3324 (N_3324,In_413,N_1566);
xnor U3325 (N_3325,N_710,N_1992);
nor U3326 (N_3326,N_1731,N_136);
xor U3327 (N_3327,N_1801,In_243);
nor U3328 (N_3328,N_840,N_1885);
or U3329 (N_3329,N_1898,N_1533);
nor U3330 (N_3330,N_1110,In_516);
and U3331 (N_3331,N_1999,In_2120);
nand U3332 (N_3332,In_1854,In_240);
and U3333 (N_3333,N_1204,N_571);
and U3334 (N_3334,In_4270,N_877);
and U3335 (N_3335,N_1737,In_4598);
xor U3336 (N_3336,N_460,In_2021);
or U3337 (N_3337,In_718,N_932);
and U3338 (N_3338,In_51,N_719);
and U3339 (N_3339,In_3781,N_171);
xnor U3340 (N_3340,In_607,In_3018);
or U3341 (N_3341,In_868,N_1448);
nor U3342 (N_3342,In_4747,N_1823);
nand U3343 (N_3343,In_445,In_4471);
and U3344 (N_3344,In_4525,N_948);
and U3345 (N_3345,N_1000,N_894);
nor U3346 (N_3346,N_455,N_161);
xnor U3347 (N_3347,N_316,N_23);
nor U3348 (N_3348,In_3127,N_1130);
nand U3349 (N_3349,In_2845,N_1529);
nor U3350 (N_3350,N_291,N_246);
xor U3351 (N_3351,N_1349,In_1244);
and U3352 (N_3352,N_1712,In_4122);
nor U3353 (N_3353,N_1430,N_486);
or U3354 (N_3354,In_4435,In_4109);
and U3355 (N_3355,N_1872,N_722);
or U3356 (N_3356,N_1450,N_1518);
and U3357 (N_3357,N_1759,In_350);
nand U3358 (N_3358,In_4524,N_160);
and U3359 (N_3359,N_509,In_3413);
and U3360 (N_3360,In_2840,In_2847);
or U3361 (N_3361,In_2596,N_791);
nor U3362 (N_3362,In_1904,In_1583);
xnor U3363 (N_3363,In_1184,N_307);
or U3364 (N_3364,In_4041,N_661);
and U3365 (N_3365,N_1544,N_805);
nor U3366 (N_3366,N_669,N_1812);
nor U3367 (N_3367,In_1072,N_1249);
xnor U3368 (N_3368,In_680,N_1074);
and U3369 (N_3369,N_519,In_1416);
or U3370 (N_3370,N_529,N_418);
and U3371 (N_3371,In_2308,In_120);
xor U3372 (N_3372,In_310,N_1778);
nand U3373 (N_3373,N_245,In_4503);
xor U3374 (N_3374,N_1004,N_1623);
nor U3375 (N_3375,In_3146,N_1752);
or U3376 (N_3376,In_455,N_568);
nor U3377 (N_3377,N_1226,In_1728);
nand U3378 (N_3378,N_566,In_1485);
nand U3379 (N_3379,In_1351,In_28);
xor U3380 (N_3380,N_154,In_98);
and U3381 (N_3381,N_1186,N_1088);
nand U3382 (N_3382,N_1319,In_3428);
and U3383 (N_3383,N_1586,In_698);
nand U3384 (N_3384,N_594,N_736);
xnor U3385 (N_3385,N_1233,N_829);
and U3386 (N_3386,N_1728,In_2474);
nand U3387 (N_3387,In_2119,N_76);
nand U3388 (N_3388,N_356,N_762);
or U3389 (N_3389,N_430,N_981);
and U3390 (N_3390,In_559,In_2711);
or U3391 (N_3391,N_1789,N_1309);
nand U3392 (N_3392,N_1781,N_542);
nand U3393 (N_3393,In_1399,N_1187);
or U3394 (N_3394,In_3537,N_392);
xnor U3395 (N_3395,In_1671,N_1117);
and U3396 (N_3396,N_1858,N_1794);
xor U3397 (N_3397,N_1687,N_1653);
and U3398 (N_3398,In_4592,N_1967);
nor U3399 (N_3399,N_1953,N_678);
xnor U3400 (N_3400,N_1570,N_436);
nor U3401 (N_3401,N_1005,N_1914);
xnor U3402 (N_3402,N_1489,In_1397);
or U3403 (N_3403,N_443,N_1487);
or U3404 (N_3404,N_564,N_1245);
nand U3405 (N_3405,N_1361,In_1565);
xor U3406 (N_3406,In_4011,N_1880);
nor U3407 (N_3407,N_1500,N_1271);
or U3408 (N_3408,In_3672,N_796);
and U3409 (N_3409,N_732,N_691);
xor U3410 (N_3410,In_3488,N_872);
and U3411 (N_3411,In_4929,N_1146);
nand U3412 (N_3412,N_1528,N_650);
and U3413 (N_3413,N_764,N_724);
nand U3414 (N_3414,In_990,N_1860);
nor U3415 (N_3415,N_1686,N_1436);
or U3416 (N_3416,N_1642,N_1971);
and U3417 (N_3417,N_820,N_558);
and U3418 (N_3418,N_812,In_4659);
nor U3419 (N_3419,In_4561,N_1538);
and U3420 (N_3420,In_4961,N_251);
or U3421 (N_3421,In_3805,In_2260);
nor U3422 (N_3422,N_177,N_1961);
and U3423 (N_3423,In_207,In_2674);
or U3424 (N_3424,In_825,In_2559);
and U3425 (N_3425,N_159,N_576);
and U3426 (N_3426,N_1861,N_863);
nand U3427 (N_3427,N_90,N_1257);
or U3428 (N_3428,N_1630,N_1399);
nor U3429 (N_3429,N_284,N_676);
and U3430 (N_3430,N_603,In_3002);
or U3431 (N_3431,N_1711,In_519);
nand U3432 (N_3432,N_1315,N_503);
and U3433 (N_3433,N_325,N_107);
or U3434 (N_3434,N_1065,N_1154);
nor U3435 (N_3435,In_3862,N_389);
nor U3436 (N_3436,N_824,N_1432);
nand U3437 (N_3437,In_1323,N_1817);
or U3438 (N_3438,N_286,N_74);
nor U3439 (N_3439,N_1452,N_165);
xor U3440 (N_3440,N_1483,N_984);
xnor U3441 (N_3441,In_4244,N_1289);
nand U3442 (N_3442,N_830,In_1414);
and U3443 (N_3443,N_1224,N_1195);
nand U3444 (N_3444,N_1702,N_379);
xor U3445 (N_3445,In_1271,N_199);
nor U3446 (N_3446,N_1015,In_915);
nor U3447 (N_3447,N_1012,In_1602);
xor U3448 (N_3448,N_1820,N_544);
nand U3449 (N_3449,N_1266,N_757);
and U3450 (N_3450,N_157,N_1259);
xnor U3451 (N_3451,N_1542,N_1353);
and U3452 (N_3452,In_924,In_4068);
nand U3453 (N_3453,In_1605,In_3885);
or U3454 (N_3454,N_1009,In_1631);
xnor U3455 (N_3455,In_1995,In_2665);
and U3456 (N_3456,N_569,N_1438);
nand U3457 (N_3457,N_1577,N_908);
or U3458 (N_3458,N_1442,N_1132);
xor U3459 (N_3459,N_413,N_1205);
or U3460 (N_3460,N_1571,N_986);
and U3461 (N_3461,N_262,N_1727);
nor U3462 (N_3462,N_1274,N_1575);
and U3463 (N_3463,N_302,N_510);
or U3464 (N_3464,N_505,In_4034);
nand U3465 (N_3465,N_949,In_1947);
xnor U3466 (N_3466,In_3783,In_357);
nor U3467 (N_3467,N_835,In_3423);
nand U3468 (N_3468,In_4834,N_1316);
nor U3469 (N_3469,In_2352,N_1371);
nand U3470 (N_3470,N_1859,In_3827);
nand U3471 (N_3471,N_125,N_1237);
nand U3472 (N_3472,In_3696,N_942);
xor U3473 (N_3473,N_1896,N_968);
and U3474 (N_3474,N_622,In_3226);
xor U3475 (N_3475,In_4585,In_3528);
nor U3476 (N_3476,N_1549,In_3944);
xor U3477 (N_3477,N_1288,N_1072);
nand U3478 (N_3478,In_3998,N_124);
and U3479 (N_3479,N_1405,In_648);
nor U3480 (N_3480,In_2984,N_414);
nand U3481 (N_3481,N_1845,N_1097);
nand U3482 (N_3482,N_1840,N_0);
nand U3483 (N_3483,N_1641,N_1116);
and U3484 (N_3484,In_1958,N_660);
nor U3485 (N_3485,N_1455,N_837);
or U3486 (N_3486,In_3673,In_239);
and U3487 (N_3487,N_81,N_575);
nand U3488 (N_3488,N_500,N_1477);
or U3489 (N_3489,N_954,N_293);
xor U3490 (N_3490,N_998,N_790);
nor U3491 (N_3491,N_1695,N_242);
xor U3492 (N_3492,N_995,In_3708);
xnor U3493 (N_3493,N_1435,In_2408);
xor U3494 (N_3494,In_2864,N_1606);
and U3495 (N_3495,N_788,N_237);
or U3496 (N_3496,In_1651,In_2150);
or U3497 (N_3497,In_428,N_1719);
nand U3498 (N_3498,In_3477,N_624);
or U3499 (N_3499,In_4532,N_1114);
xnor U3500 (N_3500,N_419,N_1831);
nand U3501 (N_3501,N_1683,N_1817);
or U3502 (N_3502,N_1657,N_500);
or U3503 (N_3503,N_1431,N_1228);
xor U3504 (N_3504,N_697,In_1500);
and U3505 (N_3505,N_318,N_932);
or U3506 (N_3506,N_1273,N_259);
nor U3507 (N_3507,N_375,N_950);
xor U3508 (N_3508,N_1884,In_2555);
nand U3509 (N_3509,In_4858,N_485);
xor U3510 (N_3510,N_371,N_317);
nor U3511 (N_3511,In_3063,N_733);
nor U3512 (N_3512,N_1502,In_3649);
nand U3513 (N_3513,N_583,In_1648);
xor U3514 (N_3514,In_1710,In_2629);
nand U3515 (N_3515,N_481,N_204);
nand U3516 (N_3516,N_1099,In_4929);
or U3517 (N_3517,N_1905,N_1740);
nand U3518 (N_3518,In_2321,N_1268);
and U3519 (N_3519,N_1338,N_1476);
or U3520 (N_3520,N_668,In_2910);
nor U3521 (N_3521,In_3678,In_657);
or U3522 (N_3522,N_1491,N_1097);
xor U3523 (N_3523,N_1500,N_1169);
or U3524 (N_3524,N_1154,N_1841);
nor U3525 (N_3525,N_1503,N_1701);
and U3526 (N_3526,N_1596,N_1508);
nor U3527 (N_3527,In_2741,In_3885);
nand U3528 (N_3528,N_1713,N_1239);
xnor U3529 (N_3529,In_4438,In_1244);
nor U3530 (N_3530,In_4728,N_148);
or U3531 (N_3531,N_916,In_4770);
nor U3532 (N_3532,N_449,N_592);
xnor U3533 (N_3533,N_1543,N_1535);
xor U3534 (N_3534,N_1328,N_1695);
xnor U3535 (N_3535,N_1017,N_474);
nor U3536 (N_3536,N_1098,In_4592);
nor U3537 (N_3537,N_932,In_593);
nand U3538 (N_3538,In_103,In_20);
or U3539 (N_3539,N_1571,N_1744);
and U3540 (N_3540,N_327,N_1752);
or U3541 (N_3541,N_573,N_226);
nor U3542 (N_3542,N_247,N_1749);
xnor U3543 (N_3543,N_945,N_688);
or U3544 (N_3544,N_723,N_1441);
nand U3545 (N_3545,In_17,N_1056);
xor U3546 (N_3546,N_1066,In_772);
or U3547 (N_3547,N_429,N_1965);
nor U3548 (N_3548,N_527,N_1532);
xnor U3549 (N_3549,N_816,In_1651);
xor U3550 (N_3550,In_1657,In_97);
nand U3551 (N_3551,In_2267,N_726);
nor U3552 (N_3552,N_1773,N_1606);
or U3553 (N_3553,N_1785,N_1655);
nand U3554 (N_3554,N_1550,In_2757);
nor U3555 (N_3555,N_1989,In_3773);
nor U3556 (N_3556,N_963,In_57);
xnor U3557 (N_3557,In_4941,N_934);
xnor U3558 (N_3558,N_1995,N_1338);
and U3559 (N_3559,In_1496,In_1092);
or U3560 (N_3560,N_143,N_382);
nand U3561 (N_3561,N_1925,N_797);
nand U3562 (N_3562,N_350,N_1827);
nor U3563 (N_3563,N_299,N_1476);
nand U3564 (N_3564,N_26,N_1758);
nand U3565 (N_3565,N_1096,N_1576);
nor U3566 (N_3566,In_4223,In_4249);
nor U3567 (N_3567,In_2398,In_4705);
nand U3568 (N_3568,In_2695,N_1753);
and U3569 (N_3569,N_1991,N_62);
nand U3570 (N_3570,N_1567,In_365);
and U3571 (N_3571,N_1464,N_596);
or U3572 (N_3572,N_1721,N_581);
and U3573 (N_3573,In_1313,In_664);
and U3574 (N_3574,N_566,N_1643);
or U3575 (N_3575,N_1306,In_644);
nand U3576 (N_3576,In_2864,N_1418);
xnor U3577 (N_3577,N_1234,In_3655);
and U3578 (N_3578,In_3426,N_1687);
xnor U3579 (N_3579,N_1043,N_341);
nand U3580 (N_3580,N_840,N_1799);
or U3581 (N_3581,N_132,N_1932);
xnor U3582 (N_3582,N_417,In_1466);
and U3583 (N_3583,In_2984,N_1889);
nor U3584 (N_3584,In_2917,In_3495);
or U3585 (N_3585,N_1689,In_2268);
or U3586 (N_3586,N_1706,In_2385);
and U3587 (N_3587,In_4068,In_2311);
nor U3588 (N_3588,N_835,N_978);
or U3589 (N_3589,In_546,N_1006);
and U3590 (N_3590,N_1758,N_89);
or U3591 (N_3591,In_3123,N_886);
or U3592 (N_3592,N_39,In_4595);
nor U3593 (N_3593,In_4327,N_1840);
nor U3594 (N_3594,N_1682,N_718);
or U3595 (N_3595,N_390,N_1471);
nand U3596 (N_3596,In_2551,N_273);
and U3597 (N_3597,In_2741,In_1891);
nand U3598 (N_3598,N_103,In_4504);
xor U3599 (N_3599,N_759,In_967);
and U3600 (N_3600,In_1359,N_61);
nor U3601 (N_3601,N_1082,In_3377);
nand U3602 (N_3602,N_377,N_613);
xor U3603 (N_3603,In_701,N_1344);
nand U3604 (N_3604,N_1842,N_75);
or U3605 (N_3605,N_1480,In_900);
xnor U3606 (N_3606,N_812,N_232);
or U3607 (N_3607,N_482,N_1890);
xnor U3608 (N_3608,N_969,In_2838);
or U3609 (N_3609,In_357,N_911);
nand U3610 (N_3610,N_386,In_1651);
and U3611 (N_3611,In_1326,In_2144);
or U3612 (N_3612,N_1014,In_4694);
nor U3613 (N_3613,N_1270,N_384);
or U3614 (N_3614,N_153,N_334);
nand U3615 (N_3615,N_1693,In_1399);
nand U3616 (N_3616,N_1031,N_1845);
or U3617 (N_3617,N_1007,N_1159);
nor U3618 (N_3618,N_1995,In_1166);
or U3619 (N_3619,N_1550,N_108);
nor U3620 (N_3620,In_1589,N_340);
or U3621 (N_3621,N_576,N_376);
and U3622 (N_3622,In_593,N_753);
nand U3623 (N_3623,N_1110,N_1739);
nand U3624 (N_3624,In_1359,In_4077);
and U3625 (N_3625,N_1328,N_1874);
nand U3626 (N_3626,N_1424,N_520);
nor U3627 (N_3627,N_1317,N_471);
xnor U3628 (N_3628,N_64,N_287);
nor U3629 (N_3629,In_4122,In_2644);
xnor U3630 (N_3630,N_1992,N_195);
nand U3631 (N_3631,N_595,In_4280);
or U3632 (N_3632,N_1488,In_144);
nor U3633 (N_3633,In_1987,N_1273);
and U3634 (N_3634,N_714,N_1886);
xnor U3635 (N_3635,N_940,N_721);
and U3636 (N_3636,In_2495,In_2854);
nand U3637 (N_3637,In_85,In_4031);
xor U3638 (N_3638,N_1821,In_1851);
or U3639 (N_3639,N_975,N_349);
xor U3640 (N_3640,N_171,In_4681);
nor U3641 (N_3641,N_1099,In_482);
nor U3642 (N_3642,N_241,N_1756);
nand U3643 (N_3643,In_357,In_3528);
or U3644 (N_3644,N_1770,N_556);
nand U3645 (N_3645,N_389,N_1528);
and U3646 (N_3646,N_1752,N_1995);
nand U3647 (N_3647,N_296,N_284);
or U3648 (N_3648,N_863,N_1767);
nor U3649 (N_3649,N_1385,N_379);
or U3650 (N_3650,N_393,N_656);
xnor U3651 (N_3651,N_214,N_1049);
nand U3652 (N_3652,N_818,In_819);
xor U3653 (N_3653,N_676,N_231);
nor U3654 (N_3654,In_592,N_470);
and U3655 (N_3655,In_2150,In_967);
nand U3656 (N_3656,In_570,N_1644);
xor U3657 (N_3657,In_2775,N_674);
nor U3658 (N_3658,N_1148,N_467);
xor U3659 (N_3659,N_384,In_759);
or U3660 (N_3660,In_299,N_1995);
xnor U3661 (N_3661,In_3327,In_3063);
and U3662 (N_3662,N_1374,N_800);
or U3663 (N_3663,In_230,N_836);
xnor U3664 (N_3664,N_756,In_4654);
nand U3665 (N_3665,In_3541,N_508);
nor U3666 (N_3666,N_1667,N_202);
nor U3667 (N_3667,N_419,In_2045);
nor U3668 (N_3668,N_92,N_1334);
xor U3669 (N_3669,N_1213,In_4406);
or U3670 (N_3670,In_3918,N_562);
nand U3671 (N_3671,N_112,N_1761);
nor U3672 (N_3672,N_158,In_1113);
or U3673 (N_3673,In_3152,N_1936);
and U3674 (N_3674,N_1977,N_1546);
nand U3675 (N_3675,N_115,N_271);
nor U3676 (N_3676,In_99,N_1803);
nor U3677 (N_3677,N_744,N_290);
nor U3678 (N_3678,In_2971,N_1669);
or U3679 (N_3679,N_262,In_607);
and U3680 (N_3680,N_1742,In_4705);
nor U3681 (N_3681,In_4034,In_2123);
or U3682 (N_3682,In_2099,In_1605);
nor U3683 (N_3683,In_2445,N_612);
nor U3684 (N_3684,N_1372,N_247);
or U3685 (N_3685,N_522,N_983);
xor U3686 (N_3686,N_796,N_40);
xnor U3687 (N_3687,In_427,In_4747);
xor U3688 (N_3688,N_673,N_1958);
xnor U3689 (N_3689,In_1176,N_1435);
nand U3690 (N_3690,N_1137,N_577);
nand U3691 (N_3691,N_785,In_3552);
xnor U3692 (N_3692,N_27,In_1422);
and U3693 (N_3693,N_1029,In_610);
and U3694 (N_3694,N_1425,In_1508);
and U3695 (N_3695,N_1087,N_446);
and U3696 (N_3696,N_711,N_865);
or U3697 (N_3697,N_92,N_460);
xor U3698 (N_3698,N_1231,In_245);
xor U3699 (N_3699,N_305,In_3965);
and U3700 (N_3700,N_654,In_3552);
or U3701 (N_3701,N_628,N_1958);
nor U3702 (N_3702,N_36,N_1347);
and U3703 (N_3703,N_1625,N_1050);
and U3704 (N_3704,N_1760,N_1985);
nor U3705 (N_3705,N_176,N_1558);
nor U3706 (N_3706,In_3375,In_2406);
or U3707 (N_3707,In_1778,In_4269);
xor U3708 (N_3708,In_3483,N_1761);
and U3709 (N_3709,N_1772,N_1924);
xnor U3710 (N_3710,N_668,N_1963);
nor U3711 (N_3711,N_1280,In_4064);
xnor U3712 (N_3712,In_2462,N_1192);
or U3713 (N_3713,In_2126,N_1883);
xor U3714 (N_3714,In_636,N_1274);
nor U3715 (N_3715,In_2598,N_1522);
and U3716 (N_3716,N_1249,N_148);
and U3717 (N_3717,N_1047,N_1844);
and U3718 (N_3718,N_329,N_1501);
and U3719 (N_3719,N_1960,N_326);
and U3720 (N_3720,In_4134,In_330);
xnor U3721 (N_3721,N_216,N_1800);
xor U3722 (N_3722,N_1650,In_4746);
xnor U3723 (N_3723,N_464,N_1286);
nor U3724 (N_3724,In_1651,N_568);
xnor U3725 (N_3725,N_764,N_261);
nand U3726 (N_3726,In_4756,N_1750);
nor U3727 (N_3727,In_150,In_867);
nor U3728 (N_3728,N_1318,In_3995);
xnor U3729 (N_3729,N_1316,N_1270);
and U3730 (N_3730,N_412,N_426);
xor U3731 (N_3731,In_608,In_1648);
or U3732 (N_3732,N_762,N_1817);
or U3733 (N_3733,N_69,N_779);
nand U3734 (N_3734,N_694,N_908);
and U3735 (N_3735,N_623,N_1656);
and U3736 (N_3736,N_1668,N_1652);
and U3737 (N_3737,In_4081,N_1451);
nor U3738 (N_3738,N_1026,In_68);
and U3739 (N_3739,N_900,N_1398);
nor U3740 (N_3740,In_2162,N_892);
and U3741 (N_3741,In_4196,In_2724);
and U3742 (N_3742,N_1706,N_258);
or U3743 (N_3743,N_1383,In_2352);
or U3744 (N_3744,N_1475,N_1354);
or U3745 (N_3745,N_1663,In_2687);
nor U3746 (N_3746,In_498,N_821);
and U3747 (N_3747,In_2438,N_1135);
nor U3748 (N_3748,N_1981,In_4448);
xor U3749 (N_3749,N_159,N_1728);
nand U3750 (N_3750,N_727,N_647);
nand U3751 (N_3751,N_730,N_1899);
nor U3752 (N_3752,In_4543,N_1767);
and U3753 (N_3753,In_2225,In_3088);
xnor U3754 (N_3754,N_1288,N_984);
or U3755 (N_3755,N_174,N_1698);
nor U3756 (N_3756,N_408,N_1770);
or U3757 (N_3757,In_2834,N_469);
or U3758 (N_3758,N_235,In_2909);
nand U3759 (N_3759,N_231,N_1171);
xor U3760 (N_3760,N_1017,In_1316);
nand U3761 (N_3761,N_1737,N_896);
nand U3762 (N_3762,In_1485,N_419);
or U3763 (N_3763,In_4521,N_918);
and U3764 (N_3764,N_696,In_1359);
or U3765 (N_3765,N_1848,N_181);
xor U3766 (N_3766,N_1897,N_1451);
xnor U3767 (N_3767,N_545,N_1035);
nand U3768 (N_3768,N_810,N_129);
nor U3769 (N_3769,In_257,N_895);
or U3770 (N_3770,N_1776,N_770);
and U3771 (N_3771,N_471,N_691);
xor U3772 (N_3772,N_966,N_351);
or U3773 (N_3773,N_170,N_927);
nand U3774 (N_3774,N_1697,N_892);
or U3775 (N_3775,N_1473,N_267);
and U3776 (N_3776,N_88,N_669);
and U3777 (N_3777,N_658,N_964);
and U3778 (N_3778,In_4544,In_1197);
and U3779 (N_3779,N_191,N_1067);
xnor U3780 (N_3780,N_735,N_1);
nand U3781 (N_3781,In_150,In_3821);
xor U3782 (N_3782,N_1406,N_627);
nor U3783 (N_3783,N_1213,N_1829);
and U3784 (N_3784,In_3362,In_1337);
nand U3785 (N_3785,N_1326,N_1180);
xnor U3786 (N_3786,In_2298,In_2055);
xor U3787 (N_3787,In_3284,N_1748);
nor U3788 (N_3788,N_1804,N_1761);
nor U3789 (N_3789,N_179,N_1001);
or U3790 (N_3790,N_1415,N_1034);
nand U3791 (N_3791,N_222,N_648);
and U3792 (N_3792,In_2059,N_1992);
and U3793 (N_3793,N_991,N_951);
xor U3794 (N_3794,N_1968,In_2663);
xor U3795 (N_3795,N_499,N_341);
nand U3796 (N_3796,N_932,N_1352);
or U3797 (N_3797,N_1841,N_618);
or U3798 (N_3798,In_1605,In_214);
nor U3799 (N_3799,N_267,In_1006);
and U3800 (N_3800,N_1539,N_85);
xor U3801 (N_3801,In_4479,N_293);
or U3802 (N_3802,N_1265,N_1391);
nand U3803 (N_3803,N_597,N_77);
xor U3804 (N_3804,N_1929,N_190);
and U3805 (N_3805,N_358,In_1730);
nand U3806 (N_3806,N_1666,N_938);
xnor U3807 (N_3807,N_697,In_1642);
and U3808 (N_3808,N_362,In_1184);
and U3809 (N_3809,N_1690,N_656);
xnor U3810 (N_3810,N_1440,N_811);
and U3811 (N_3811,N_140,N_1989);
and U3812 (N_3812,N_598,N_952);
nand U3813 (N_3813,In_2012,N_4);
or U3814 (N_3814,N_1901,In_856);
and U3815 (N_3815,N_1056,N_1936);
or U3816 (N_3816,N_743,In_3698);
nand U3817 (N_3817,N_1300,N_446);
nand U3818 (N_3818,In_3018,N_1544);
or U3819 (N_3819,N_1878,In_2385);
or U3820 (N_3820,In_4471,In_4543);
nor U3821 (N_3821,N_216,In_831);
xor U3822 (N_3822,N_1901,N_937);
xnor U3823 (N_3823,N_1342,N_749);
or U3824 (N_3824,N_319,N_1713);
nor U3825 (N_3825,N_1028,N_1363);
xor U3826 (N_3826,N_721,In_4803);
nor U3827 (N_3827,N_520,N_123);
nor U3828 (N_3828,N_1576,N_81);
xor U3829 (N_3829,N_209,N_95);
nand U3830 (N_3830,In_3977,N_1434);
nand U3831 (N_3831,N_1187,In_712);
or U3832 (N_3832,N_902,N_41);
and U3833 (N_3833,N_571,N_1008);
nor U3834 (N_3834,N_193,N_645);
nand U3835 (N_3835,N_121,N_1956);
nor U3836 (N_3836,In_1524,N_361);
and U3837 (N_3837,In_2381,N_120);
nand U3838 (N_3838,N_1921,N_618);
and U3839 (N_3839,In_4018,In_4721);
nand U3840 (N_3840,N_403,In_4848);
or U3841 (N_3841,N_1068,In_4998);
nor U3842 (N_3842,N_342,In_3584);
nand U3843 (N_3843,N_1557,N_11);
xor U3844 (N_3844,N_90,In_3495);
and U3845 (N_3845,In_4664,In_3418);
nand U3846 (N_3846,N_782,In_2411);
nor U3847 (N_3847,N_1038,In_2381);
xor U3848 (N_3848,N_87,N_120);
or U3849 (N_3849,N_458,In_2917);
or U3850 (N_3850,In_3204,N_993);
and U3851 (N_3851,In_3373,N_975);
xnor U3852 (N_3852,In_602,In_4068);
xor U3853 (N_3853,N_1378,N_1779);
or U3854 (N_3854,N_1527,In_3438);
or U3855 (N_3855,N_1016,N_336);
or U3856 (N_3856,In_829,N_646);
nor U3857 (N_3857,N_1671,N_1519);
xnor U3858 (N_3858,N_200,N_1287);
or U3859 (N_3859,In_2109,N_483);
and U3860 (N_3860,N_454,N_866);
or U3861 (N_3861,N_950,In_4435);
and U3862 (N_3862,N_1461,N_1641);
and U3863 (N_3863,N_209,In_694);
and U3864 (N_3864,N_245,N_1988);
and U3865 (N_3865,In_16,N_506);
xnor U3866 (N_3866,In_3,N_1102);
nand U3867 (N_3867,N_584,In_4848);
and U3868 (N_3868,N_1577,N_275);
or U3869 (N_3869,N_817,N_1013);
or U3870 (N_3870,N_971,In_2434);
xor U3871 (N_3871,In_2035,N_687);
nand U3872 (N_3872,N_1140,In_1414);
or U3873 (N_3873,In_2686,N_1632);
nor U3874 (N_3874,N_258,N_1608);
xor U3875 (N_3875,N_1920,In_2120);
xnor U3876 (N_3876,N_688,N_1319);
or U3877 (N_3877,In_1184,N_1841);
or U3878 (N_3878,N_1279,In_2268);
xor U3879 (N_3879,N_1864,N_368);
or U3880 (N_3880,N_269,N_1699);
nor U3881 (N_3881,N_685,In_1906);
nor U3882 (N_3882,In_609,N_1730);
nor U3883 (N_3883,In_3967,In_609);
xnor U3884 (N_3884,In_4525,In_2445);
nor U3885 (N_3885,N_1602,In_3046);
and U3886 (N_3886,N_654,N_1444);
xnor U3887 (N_3887,N_24,N_696);
nand U3888 (N_3888,N_747,N_89);
nor U3889 (N_3889,N_440,N_605);
nand U3890 (N_3890,N_1862,N_1149);
nand U3891 (N_3891,N_1920,In_3552);
xnor U3892 (N_3892,N_744,N_1168);
nor U3893 (N_3893,N_1186,N_1399);
nand U3894 (N_3894,N_1394,N_772);
and U3895 (N_3895,N_1533,In_3995);
nand U3896 (N_3896,N_819,N_1196);
nand U3897 (N_3897,N_60,In_4636);
nand U3898 (N_3898,N_272,N_948);
or U3899 (N_3899,In_3605,In_2216);
nor U3900 (N_3900,In_1613,N_415);
xor U3901 (N_3901,N_759,In_3874);
xor U3902 (N_3902,N_1547,N_964);
nor U3903 (N_3903,In_177,N_1087);
nand U3904 (N_3904,In_4103,In_4781);
nor U3905 (N_3905,In_2724,In_3423);
or U3906 (N_3906,N_1478,N_935);
and U3907 (N_3907,In_3981,N_1328);
and U3908 (N_3908,N_1232,N_1572);
or U3909 (N_3909,In_4929,N_284);
xor U3910 (N_3910,N_1488,N_448);
xnor U3911 (N_3911,In_3297,In_2911);
and U3912 (N_3912,In_4636,In_4081);
or U3913 (N_3913,N_1826,In_239);
and U3914 (N_3914,In_4016,N_1010);
xnor U3915 (N_3915,In_4983,N_911);
xor U3916 (N_3916,N_200,N_841);
nor U3917 (N_3917,N_1883,In_900);
or U3918 (N_3918,N_621,N_1213);
or U3919 (N_3919,N_1739,In_3783);
nand U3920 (N_3920,In_3363,In_4770);
nand U3921 (N_3921,N_1349,N_1304);
nor U3922 (N_3922,N_1592,N_1434);
or U3923 (N_3923,N_689,N_1434);
nand U3924 (N_3924,N_629,N_828);
nand U3925 (N_3925,N_97,In_1325);
nor U3926 (N_3926,In_4582,In_3509);
or U3927 (N_3927,In_4435,N_1274);
nor U3928 (N_3928,In_4713,In_1500);
or U3929 (N_3929,N_34,In_4973);
nand U3930 (N_3930,In_3483,N_1);
xnor U3931 (N_3931,N_1814,N_1107);
xor U3932 (N_3932,N_141,N_1340);
nor U3933 (N_3933,N_775,N_553);
nand U3934 (N_3934,In_3605,In_4314);
nand U3935 (N_3935,N_1797,N_310);
nand U3936 (N_3936,N_1204,N_188);
nand U3937 (N_3937,In_570,N_1588);
and U3938 (N_3938,N_1067,N_138);
and U3939 (N_3939,In_1253,N_1084);
and U3940 (N_3940,In_3783,N_729);
xnor U3941 (N_3941,N_1022,In_214);
xor U3942 (N_3942,N_1174,N_1188);
or U3943 (N_3943,N_576,In_3373);
nor U3944 (N_3944,N_1470,In_2888);
or U3945 (N_3945,N_1695,In_2294);
xor U3946 (N_3946,N_1178,In_4438);
and U3947 (N_3947,N_1268,N_1931);
nand U3948 (N_3948,N_1568,N_756);
xor U3949 (N_3949,N_1386,In_2407);
nand U3950 (N_3950,N_949,N_670);
xor U3951 (N_3951,N_437,N_1965);
and U3952 (N_3952,N_1069,N_687);
or U3953 (N_3953,N_508,N_1589);
nand U3954 (N_3954,N_1686,In_577);
and U3955 (N_3955,N_843,N_1357);
xor U3956 (N_3956,In_145,N_1884);
nand U3957 (N_3957,N_662,N_485);
nand U3958 (N_3958,N_1204,In_1648);
nor U3959 (N_3959,In_256,In_2216);
or U3960 (N_3960,N_811,N_55);
and U3961 (N_3961,N_1807,N_1923);
or U3962 (N_3962,N_756,In_4915);
xor U3963 (N_3963,N_1422,In_4223);
or U3964 (N_3964,In_4840,N_56);
nor U3965 (N_3965,N_745,In_1658);
nor U3966 (N_3966,N_1963,In_2128);
nand U3967 (N_3967,N_242,N_1796);
and U3968 (N_3968,In_855,N_1654);
nand U3969 (N_3969,In_3152,N_1138);
xor U3970 (N_3970,In_4624,N_1506);
xor U3971 (N_3971,In_1892,N_645);
or U3972 (N_3972,In_1979,N_1295);
and U3973 (N_3973,In_1591,N_312);
nand U3974 (N_3974,In_1728,N_498);
and U3975 (N_3975,In_4061,In_1170);
or U3976 (N_3976,N_1829,In_1316);
or U3977 (N_3977,N_847,In_3918);
xor U3978 (N_3978,N_232,In_2437);
or U3979 (N_3979,In_2041,In_616);
or U3980 (N_3980,In_3119,In_3495);
or U3981 (N_3981,N_653,In_3977);
and U3982 (N_3982,In_1768,In_4411);
and U3983 (N_3983,N_754,In_1208);
or U3984 (N_3984,In_2006,N_786);
nand U3985 (N_3985,N_1804,In_3196);
xnor U3986 (N_3986,N_1888,N_222);
nand U3987 (N_3987,N_1547,N_1071);
and U3988 (N_3988,N_661,In_980);
nand U3989 (N_3989,In_3907,N_105);
and U3990 (N_3990,N_1598,In_2359);
and U3991 (N_3991,In_1287,N_536);
xnor U3992 (N_3992,N_1875,In_1710);
nand U3993 (N_3993,In_65,In_4077);
nor U3994 (N_3994,N_535,N_251);
nor U3995 (N_3995,N_261,N_126);
nor U3996 (N_3996,N_347,In_199);
and U3997 (N_3997,N_1673,N_919);
xnor U3998 (N_3998,In_3862,N_52);
nor U3999 (N_3999,N_1694,N_1858);
nor U4000 (N_4000,N_2408,N_2503);
xnor U4001 (N_4001,N_2181,N_2369);
or U4002 (N_4002,N_2627,N_2763);
nand U4003 (N_4003,N_2151,N_3043);
and U4004 (N_4004,N_2126,N_2402);
or U4005 (N_4005,N_2283,N_3110);
or U4006 (N_4006,N_3204,N_3594);
xnor U4007 (N_4007,N_3459,N_3544);
xor U4008 (N_4008,N_2226,N_2866);
or U4009 (N_4009,N_3305,N_3163);
and U4010 (N_4010,N_3773,N_3453);
xnor U4011 (N_4011,N_2237,N_3994);
and U4012 (N_4012,N_3018,N_2939);
nand U4013 (N_4013,N_3705,N_3801);
and U4014 (N_4014,N_2812,N_3216);
nor U4015 (N_4015,N_3091,N_2919);
and U4016 (N_4016,N_3455,N_2212);
xor U4017 (N_4017,N_2047,N_2403);
and U4018 (N_4018,N_2242,N_3959);
xor U4019 (N_4019,N_2593,N_2642);
or U4020 (N_4020,N_3001,N_2329);
or U4021 (N_4021,N_2365,N_2757);
and U4022 (N_4022,N_2167,N_2896);
nor U4023 (N_4023,N_2509,N_2028);
nand U4024 (N_4024,N_3527,N_3341);
nor U4025 (N_4025,N_3424,N_2304);
xor U4026 (N_4026,N_3000,N_3514);
nor U4027 (N_4027,N_3239,N_2565);
and U4028 (N_4028,N_3462,N_2613);
and U4029 (N_4029,N_3195,N_3402);
nor U4030 (N_4030,N_2094,N_3167);
xor U4031 (N_4031,N_3268,N_2779);
nand U4032 (N_4032,N_3059,N_2506);
or U4033 (N_4033,N_2364,N_2920);
or U4034 (N_4034,N_3991,N_2159);
or U4035 (N_4035,N_2837,N_2204);
xor U4036 (N_4036,N_2698,N_2886);
or U4037 (N_4037,N_3207,N_2451);
nor U4038 (N_4038,N_2394,N_3966);
nand U4039 (N_4039,N_2325,N_3182);
and U4040 (N_4040,N_3736,N_3480);
and U4041 (N_4041,N_2553,N_2822);
and U4042 (N_4042,N_2649,N_2046);
xor U4043 (N_4043,N_3977,N_2287);
nor U4044 (N_4044,N_3869,N_2589);
nor U4045 (N_4045,N_2623,N_2755);
xor U4046 (N_4046,N_3866,N_2820);
or U4047 (N_4047,N_2495,N_3232);
and U4048 (N_4048,N_2907,N_2505);
nand U4049 (N_4049,N_2860,N_2806);
nand U4050 (N_4050,N_2307,N_3580);
or U4051 (N_4051,N_3283,N_2691);
or U4052 (N_4052,N_2770,N_2834);
or U4053 (N_4053,N_2957,N_3130);
xor U4054 (N_4054,N_3771,N_3115);
nand U4055 (N_4055,N_3039,N_3149);
and U4056 (N_4056,N_3800,N_3924);
xor U4057 (N_4057,N_2268,N_3260);
nor U4058 (N_4058,N_2074,N_2359);
xor U4059 (N_4059,N_3523,N_2303);
xor U4060 (N_4060,N_3982,N_3882);
nor U4061 (N_4061,N_2174,N_3682);
xnor U4062 (N_4062,N_3999,N_2780);
nand U4063 (N_4063,N_3088,N_3905);
xnor U4064 (N_4064,N_2945,N_2153);
nand U4065 (N_4065,N_2580,N_3593);
and U4066 (N_4066,N_2625,N_3992);
nand U4067 (N_4067,N_2290,N_2192);
nand U4068 (N_4068,N_3577,N_3567);
nor U4069 (N_4069,N_3666,N_3900);
nor U4070 (N_4070,N_2946,N_3173);
nor U4071 (N_4071,N_3152,N_3299);
nor U4072 (N_4072,N_3484,N_2319);
nand U4073 (N_4073,N_3011,N_3450);
and U4074 (N_4074,N_3121,N_3243);
nor U4075 (N_4075,N_2500,N_2578);
nor U4076 (N_4076,N_2947,N_3443);
xor U4077 (N_4077,N_2677,N_3019);
nor U4078 (N_4078,N_2670,N_2768);
or U4079 (N_4079,N_2390,N_2607);
or U4080 (N_4080,N_3409,N_2692);
nor U4081 (N_4081,N_3660,N_2801);
or U4082 (N_4082,N_2327,N_2760);
xor U4083 (N_4083,N_2299,N_2169);
or U4084 (N_4084,N_2416,N_2221);
nor U4085 (N_4085,N_3553,N_2111);
or U4086 (N_4086,N_2023,N_2342);
and U4087 (N_4087,N_3472,N_2675);
nand U4088 (N_4088,N_3194,N_2977);
nor U4089 (N_4089,N_2955,N_3368);
nor U4090 (N_4090,N_2051,N_2889);
or U4091 (N_4091,N_2350,N_3744);
nor U4092 (N_4092,N_3072,N_3071);
and U4093 (N_4093,N_3143,N_2731);
or U4094 (N_4094,N_2586,N_2893);
nand U4095 (N_4095,N_3828,N_2256);
or U4096 (N_4096,N_2213,N_3451);
nor U4097 (N_4097,N_3735,N_2743);
nand U4098 (N_4098,N_3360,N_3141);
and U4099 (N_4099,N_2699,N_2784);
or U4100 (N_4100,N_3648,N_2421);
nor U4101 (N_4101,N_3494,N_2324);
nand U4102 (N_4102,N_2452,N_2116);
or U4103 (N_4103,N_3791,N_2210);
nor U4104 (N_4104,N_2838,N_2217);
nand U4105 (N_4105,N_2693,N_2229);
and U4106 (N_4106,N_3270,N_2869);
nor U4107 (N_4107,N_2783,N_3821);
xor U4108 (N_4108,N_2037,N_3281);
or U4109 (N_4109,N_2078,N_3813);
xnor U4110 (N_4110,N_3090,N_3551);
nor U4111 (N_4111,N_2962,N_3411);
nor U4112 (N_4112,N_2720,N_2152);
or U4113 (N_4113,N_2469,N_2845);
nor U4114 (N_4114,N_3350,N_3016);
nand U4115 (N_4115,N_3668,N_2571);
xnor U4116 (N_4116,N_3199,N_2224);
xor U4117 (N_4117,N_2292,N_2133);
nor U4118 (N_4118,N_2695,N_3446);
nand U4119 (N_4119,N_2501,N_3502);
and U4120 (N_4120,N_2070,N_2227);
xnor U4121 (N_4121,N_2483,N_2923);
nor U4122 (N_4122,N_2308,N_2234);
nand U4123 (N_4123,N_2913,N_2983);
or U4124 (N_4124,N_2712,N_3498);
or U4125 (N_4125,N_2218,N_2246);
xor U4126 (N_4126,N_3843,N_3838);
xor U4127 (N_4127,N_2828,N_2826);
nand U4128 (N_4128,N_3908,N_2877);
and U4129 (N_4129,N_3790,N_2902);
and U4130 (N_4130,N_2027,N_3844);
and U4131 (N_4131,N_2665,N_3321);
and U4132 (N_4132,N_3324,N_3868);
nand U4133 (N_4133,N_3511,N_2008);
nand U4134 (N_4134,N_3720,N_2568);
and U4135 (N_4135,N_3234,N_2089);
xor U4136 (N_4136,N_3903,N_2663);
nor U4137 (N_4137,N_3947,N_2278);
or U4138 (N_4138,N_2482,N_2778);
nand U4139 (N_4139,N_2414,N_2895);
or U4140 (N_4140,N_2117,N_3665);
or U4141 (N_4141,N_2824,N_2848);
nor U4142 (N_4142,N_2658,N_2015);
nor U4143 (N_4143,N_2379,N_3541);
xor U4144 (N_4144,N_2740,N_3265);
or U4145 (N_4145,N_3425,N_3343);
nor U4146 (N_4146,N_2924,N_3670);
or U4147 (N_4147,N_2805,N_2633);
and U4148 (N_4148,N_3871,N_3520);
nand U4149 (N_4149,N_3249,N_2569);
nand U4150 (N_4150,N_2448,N_3953);
and U4151 (N_4151,N_3747,N_2567);
nand U4152 (N_4152,N_2796,N_2711);
nor U4153 (N_4153,N_2534,N_2121);
nor U4154 (N_4154,N_3269,N_2953);
or U4155 (N_4155,N_2943,N_3228);
and U4156 (N_4156,N_2411,N_3925);
nand U4157 (N_4157,N_3189,N_3898);
or U4158 (N_4158,N_3608,N_2185);
and U4159 (N_4159,N_2135,N_2491);
nand U4160 (N_4160,N_2171,N_2279);
nand U4161 (N_4161,N_3555,N_3236);
xnor U4162 (N_4162,N_2526,N_2125);
and U4163 (N_4163,N_2499,N_2694);
xor U4164 (N_4164,N_2490,N_3561);
nor U4165 (N_4165,N_3427,N_2422);
and U4166 (N_4166,N_2005,N_2372);
nand U4167 (N_4167,N_3897,N_3183);
or U4168 (N_4168,N_3622,N_2425);
nand U4169 (N_4169,N_3217,N_2404);
nand U4170 (N_4170,N_3598,N_2540);
xnor U4171 (N_4171,N_2487,N_2198);
nor U4172 (N_4172,N_3979,N_2407);
or U4173 (N_4173,N_2459,N_2925);
and U4174 (N_4174,N_3848,N_3146);
nand U4175 (N_4175,N_3873,N_3487);
and U4176 (N_4176,N_3614,N_3308);
nor U4177 (N_4177,N_2428,N_3406);
nor U4178 (N_4178,N_3175,N_2258);
nor U4179 (N_4179,N_2678,N_3342);
nor U4180 (N_4180,N_3403,N_3361);
and U4181 (N_4181,N_3857,N_3050);
xnor U4182 (N_4182,N_2614,N_2131);
nor U4183 (N_4183,N_2892,N_2274);
nand U4184 (N_4184,N_3086,N_2441);
and U4185 (N_4185,N_2039,N_2315);
nand U4186 (N_4186,N_2998,N_3082);
nand U4187 (N_4187,N_2392,N_3595);
or U4188 (N_4188,N_3714,N_3917);
xor U4189 (N_4189,N_3267,N_2944);
and U4190 (N_4190,N_3884,N_3394);
and U4191 (N_4191,N_3279,N_3205);
and U4192 (N_4192,N_2478,N_3762);
and U4193 (N_4193,N_3988,N_2249);
and U4194 (N_4194,N_3878,N_3677);
xnor U4195 (N_4195,N_3069,N_3290);
or U4196 (N_4196,N_3809,N_3437);
nand U4197 (N_4197,N_3272,N_2208);
nor U4198 (N_4198,N_3847,N_3395);
xor U4199 (N_4199,N_3079,N_3726);
and U4200 (N_4200,N_3004,N_3300);
nor U4201 (N_4201,N_3392,N_2053);
and U4202 (N_4202,N_3795,N_2044);
and U4203 (N_4203,N_3646,N_3027);
or U4204 (N_4204,N_2050,N_3775);
nand U4205 (N_4205,N_2163,N_3597);
or U4206 (N_4206,N_3811,N_2930);
and U4207 (N_4207,N_2343,N_2137);
nand U4208 (N_4208,N_3123,N_3635);
nor U4209 (N_4209,N_2492,N_2069);
nand U4210 (N_4210,N_3683,N_3533);
xnor U4211 (N_4211,N_2366,N_3231);
and U4212 (N_4212,N_3763,N_2259);
and U4213 (N_4213,N_3688,N_2465);
or U4214 (N_4214,N_3074,N_2684);
xor U4215 (N_4215,N_3255,N_2062);
nor U4216 (N_4216,N_2852,N_2751);
nand U4217 (N_4217,N_3081,N_2918);
and U4218 (N_4218,N_2965,N_3824);
and U4219 (N_4219,N_2240,N_2143);
nor U4220 (N_4220,N_2466,N_2543);
nand U4221 (N_4221,N_2029,N_2538);
nand U4222 (N_4222,N_3995,N_2297);
or U4223 (N_4223,N_3565,N_2244);
nand U4224 (N_4224,N_3700,N_3631);
nor U4225 (N_4225,N_2759,N_2401);
and U4226 (N_4226,N_2436,N_2864);
or U4227 (N_4227,N_2427,N_2903);
and U4228 (N_4228,N_2030,N_3754);
nor U4229 (N_4229,N_2187,N_3799);
xnor U4230 (N_4230,N_3549,N_2898);
and U4231 (N_4231,N_3781,N_2055);
or U4232 (N_4232,N_2929,N_2904);
nand U4233 (N_4233,N_3417,N_3637);
and U4234 (N_4234,N_3345,N_2724);
and U4235 (N_4235,N_3226,N_2238);
and U4236 (N_4236,N_3398,N_3960);
nor U4237 (N_4237,N_3535,N_2064);
xnor U4238 (N_4238,N_2042,N_3061);
nor U4239 (N_4239,N_2537,N_3766);
xor U4240 (N_4240,N_3929,N_3056);
and U4241 (N_4241,N_3296,N_2621);
or U4242 (N_4242,N_3547,N_2622);
or U4243 (N_4243,N_2606,N_3349);
or U4244 (N_4244,N_2197,N_2874);
nor U4245 (N_4245,N_3812,N_2950);
nand U4246 (N_4246,N_3554,N_2849);
or U4247 (N_4247,N_2093,N_3574);
nor U4248 (N_4248,N_3471,N_2114);
and U4249 (N_4249,N_2188,N_2917);
nor U4250 (N_4250,N_3522,N_3332);
xor U4251 (N_4251,N_3788,N_3951);
xnor U4252 (N_4252,N_3859,N_3264);
and U4253 (N_4253,N_3853,N_3083);
nor U4254 (N_4254,N_3385,N_2437);
or U4255 (N_4255,N_3619,N_2827);
xor U4256 (N_4256,N_2858,N_3060);
xnor U4257 (N_4257,N_3213,N_2179);
nor U4258 (N_4258,N_2433,N_3664);
nand U4259 (N_4259,N_3286,N_3174);
xnor U4260 (N_4260,N_2150,N_3495);
or U4261 (N_4261,N_3085,N_3315);
nand U4262 (N_4262,N_2843,N_2815);
and U4263 (N_4263,N_3919,N_2970);
nor U4264 (N_4264,N_3669,N_2979);
nand U4265 (N_4265,N_3302,N_3331);
and U4266 (N_4266,N_2548,N_2563);
and U4267 (N_4267,N_2257,N_2371);
and U4268 (N_4268,N_3954,N_2009);
and U4269 (N_4269,N_2672,N_2104);
or U4270 (N_4270,N_2486,N_3662);
nor U4271 (N_4271,N_2986,N_2254);
or U4272 (N_4272,N_3414,N_3944);
and U4273 (N_4273,N_3629,N_3005);
nand U4274 (N_4274,N_2875,N_2583);
nor U4275 (N_4275,N_3126,N_2635);
xnor U4276 (N_4276,N_2921,N_2758);
and U4277 (N_4277,N_3038,N_3576);
or U4278 (N_4278,N_3250,N_3815);
nor U4279 (N_4279,N_3891,N_3021);
or U4280 (N_4280,N_2850,N_2338);
or U4281 (N_4281,N_3109,N_3002);
nand U4282 (N_4282,N_2034,N_2588);
nor U4283 (N_4283,N_2656,N_2611);
or U4284 (N_4284,N_2475,N_3147);
xor U4285 (N_4285,N_2901,N_3024);
xnor U4286 (N_4286,N_2870,N_3928);
nand U4287 (N_4287,N_2739,N_3707);
xor U4288 (N_4288,N_2032,N_2142);
xor U4289 (N_4289,N_2887,N_2453);
nor U4290 (N_4290,N_3972,N_2652);
or U4291 (N_4291,N_3499,N_2400);
and U4292 (N_4292,N_2219,N_3877);
nor U4293 (N_4293,N_3568,N_2443);
or U4294 (N_4294,N_3185,N_3320);
and U4295 (N_4295,N_3783,N_2952);
nand U4296 (N_4296,N_3317,N_2000);
nand U4297 (N_4297,N_2630,N_3470);
or U4298 (N_4298,N_3990,N_3628);
or U4299 (N_4299,N_2967,N_3710);
xor U4300 (N_4300,N_3952,N_3641);
nand U4301 (N_4301,N_3823,N_3810);
xor U4302 (N_4302,N_2629,N_2761);
nor U4303 (N_4303,N_2271,N_3491);
xnor U4304 (N_4304,N_2086,N_3201);
and U4305 (N_4305,N_2239,N_2141);
or U4306 (N_4306,N_3894,N_2510);
xnor U4307 (N_4307,N_2512,N_3846);
and U4308 (N_4308,N_3372,N_2080);
and U4309 (N_4309,N_3263,N_2134);
or U4310 (N_4310,N_2288,N_3640);
and U4311 (N_4311,N_3077,N_3609);
xor U4312 (N_4312,N_3041,N_2103);
and U4313 (N_4313,N_2281,N_2582);
and U4314 (N_4314,N_3776,N_3772);
and U4315 (N_4315,N_2738,N_2183);
nand U4316 (N_4316,N_2682,N_3620);
nand U4317 (N_4317,N_3760,N_3508);
nand U4318 (N_4318,N_3486,N_2429);
xnor U4319 (N_4319,N_2595,N_2581);
nor U4320 (N_4320,N_3093,N_3068);
and U4321 (N_4321,N_3557,N_3507);
or U4322 (N_4322,N_2576,N_2241);
nor U4323 (N_4323,N_2651,N_3337);
and U4324 (N_4324,N_2781,N_3465);
nor U4325 (N_4325,N_3923,N_3626);
nand U4326 (N_4326,N_2749,N_2992);
and U4327 (N_4327,N_2599,N_2835);
and U4328 (N_4328,N_3131,N_2518);
nor U4329 (N_4329,N_2912,N_3055);
or U4330 (N_4330,N_2666,N_2881);
nand U4331 (N_4331,N_3856,N_2194);
and U4332 (N_4332,N_3280,N_2270);
and U4333 (N_4333,N_3684,N_3311);
xor U4334 (N_4334,N_2648,N_2585);
and U4335 (N_4335,N_3503,N_3464);
and U4336 (N_4336,N_2012,N_2277);
or U4337 (N_4337,N_3095,N_3833);
or U4338 (N_4338,N_2211,N_2742);
xor U4339 (N_4339,N_2559,N_3901);
xor U4340 (N_4340,N_2847,N_3984);
nor U4341 (N_4341,N_3896,N_3934);
nor U4342 (N_4342,N_2940,N_3671);
nor U4343 (N_4343,N_3330,N_3753);
xnor U4344 (N_4344,N_3616,N_2332);
or U4345 (N_4345,N_3732,N_2098);
nor U4346 (N_4346,N_2430,N_3571);
and U4347 (N_4347,N_3266,N_3556);
and U4348 (N_4348,N_3135,N_3841);
or U4349 (N_4349,N_3657,N_3780);
or U4350 (N_4350,N_3344,N_3393);
and U4351 (N_4351,N_3731,N_3906);
or U4352 (N_4352,N_3017,N_3757);
and U4353 (N_4353,N_2233,N_2148);
and U4354 (N_4354,N_3063,N_2871);
nor U4355 (N_4355,N_3240,N_3652);
nor U4356 (N_4356,N_3764,N_2832);
nor U4357 (N_4357,N_2190,N_2247);
and U4358 (N_4358,N_3474,N_2667);
xnor U4359 (N_4359,N_2113,N_3940);
nand U4360 (N_4360,N_2120,N_2976);
xor U4361 (N_4361,N_2890,N_3530);
or U4362 (N_4362,N_2508,N_2293);
and U4363 (N_4363,N_3310,N_3113);
nor U4364 (N_4364,N_2426,N_3307);
or U4365 (N_4365,N_3927,N_2591);
xnor U4366 (N_4366,N_2146,N_2434);
or U4367 (N_4367,N_2145,N_2147);
nand U4368 (N_4368,N_2022,N_2232);
or U4369 (N_4369,N_3180,N_2792);
and U4370 (N_4370,N_2091,N_3448);
and U4371 (N_4371,N_3165,N_3981);
and U4372 (N_4372,N_2255,N_3111);
or U4373 (N_4373,N_3687,N_2320);
and U4374 (N_4374,N_2322,N_3383);
nand U4375 (N_4375,N_3604,N_3301);
nor U4376 (N_4376,N_3108,N_3492);
nand U4377 (N_4377,N_3872,N_3118);
or U4378 (N_4378,N_2767,N_2865);
xnor U4379 (N_4379,N_3158,N_2790);
xnor U4380 (N_4380,N_2942,N_3980);
nor U4381 (N_4381,N_3220,N_3161);
nor U4382 (N_4382,N_3209,N_2624);
nand U4383 (N_4383,N_2689,N_2096);
and U4384 (N_4384,N_2765,N_3798);
and U4385 (N_4385,N_3340,N_3410);
xnor U4386 (N_4386,N_2982,N_3658);
or U4387 (N_4387,N_2054,N_2200);
and U4388 (N_4388,N_2574,N_2418);
and U4389 (N_4389,N_2498,N_3475);
xnor U4390 (N_4390,N_2937,N_3329);
xor U4391 (N_4391,N_3262,N_2215);
nand U4392 (N_4392,N_2052,N_3151);
or U4393 (N_4393,N_2747,N_2019);
and U4394 (N_4394,N_3193,N_2417);
nor U4395 (N_4395,N_3627,N_3052);
nand U4396 (N_4396,N_2730,N_3367);
nor U4397 (N_4397,N_2162,N_3238);
or U4398 (N_4398,N_2377,N_2470);
nor U4399 (N_4399,N_3718,N_2284);
nand U4400 (N_4400,N_3883,N_3663);
nand U4401 (N_4401,N_2594,N_2802);
nor U4402 (N_4402,N_2529,N_2524);
or U4403 (N_4403,N_3701,N_3770);
or U4404 (N_4404,N_2076,N_2173);
nand U4405 (N_4405,N_2934,N_3560);
nand U4406 (N_4406,N_2230,N_2991);
and U4407 (N_4407,N_2097,N_3933);
xnor U4408 (N_4408,N_2590,N_2248);
xnor U4409 (N_4409,N_2741,N_3588);
and U4410 (N_4410,N_3765,N_3117);
or U4411 (N_4411,N_3945,N_3440);
and U4412 (N_4412,N_2798,N_2049);
nor U4413 (N_4413,N_3371,N_3287);
xor U4414 (N_4414,N_3012,N_2951);
and U4415 (N_4415,N_3501,N_2024);
nor U4416 (N_4416,N_2603,N_2857);
and U4417 (N_4417,N_2650,N_3755);
or U4418 (N_4418,N_3040,N_3137);
nor U4419 (N_4419,N_3741,N_3950);
nor U4420 (N_4420,N_2880,N_2260);
and U4421 (N_4421,N_2683,N_2931);
or U4422 (N_4422,N_2811,N_3820);
or U4423 (N_4423,N_2885,N_2803);
nand U4424 (N_4424,N_3029,N_2963);
xnor U4425 (N_4425,N_3642,N_2729);
nor U4426 (N_4426,N_2419,N_3046);
nand U4427 (N_4427,N_3469,N_3221);
and U4428 (N_4428,N_3352,N_3087);
nand U4429 (N_4429,N_3322,N_3603);
xnor U4430 (N_4430,N_2696,N_2669);
or U4431 (N_4431,N_3862,N_3515);
and U4432 (N_4432,N_2357,N_2017);
nor U4433 (N_4433,N_2384,N_2549);
or U4434 (N_4434,N_2791,N_3759);
nand U4435 (N_4435,N_2175,N_3025);
nor U4436 (N_4436,N_3822,N_3191);
and U4437 (N_4437,N_3997,N_2984);
nand U4438 (N_4438,N_2207,N_3478);
xnor U4439 (N_4439,N_2618,N_3415);
or U4440 (N_4440,N_3605,N_2846);
or U4441 (N_4441,N_3696,N_2455);
xor U4442 (N_4442,N_2620,N_2804);
or U4443 (N_4443,N_3778,N_2385);
nand U4444 (N_4444,N_2557,N_2602);
and U4445 (N_4445,N_3080,N_3654);
xnor U4446 (N_4446,N_3690,N_3454);
and U4447 (N_4447,N_2960,N_3558);
or U4448 (N_4448,N_3479,N_3548);
nand U4449 (N_4449,N_2494,N_3035);
or U4450 (N_4450,N_3697,N_2476);
nor U4451 (N_4451,N_3030,N_3653);
nor U4452 (N_4452,N_3374,N_2196);
nor U4453 (N_4453,N_3084,N_3888);
and U4454 (N_4454,N_2285,N_3965);
and U4455 (N_4455,N_3792,N_3887);
xnor U4456 (N_4456,N_3463,N_3139);
or U4457 (N_4457,N_2844,N_3336);
or U4458 (N_4458,N_3739,N_2861);
xnor U4459 (N_4459,N_2380,N_2410);
xor U4460 (N_4460,N_3390,N_3309);
xnor U4461 (N_4461,N_3543,N_2671);
nand U4462 (N_4462,N_3699,N_3124);
or U4463 (N_4463,N_3659,N_2573);
nor U4464 (N_4464,N_2993,N_3719);
or U4465 (N_4465,N_3806,N_2467);
xnor U4466 (N_4466,N_2214,N_3623);
xnor U4467 (N_4467,N_3254,N_3391);
and U4468 (N_4468,N_3566,N_3845);
or U4469 (N_4469,N_2966,N_2598);
or U4470 (N_4470,N_2922,N_3733);
nor U4471 (N_4471,N_2617,N_3876);
xor U4472 (N_4472,N_3667,N_2106);
or U4473 (N_4473,N_2818,N_2507);
nand U4474 (N_4474,N_3051,N_2109);
nand U4475 (N_4475,N_3839,N_2286);
xnor U4476 (N_4476,N_3203,N_3721);
nand U4477 (N_4477,N_2128,N_3633);
xor U4478 (N_4478,N_2444,N_3456);
xor U4479 (N_4479,N_2166,N_2555);
nand U4480 (N_4480,N_3819,N_2535);
and U4481 (N_4481,N_3916,N_3192);
nor U4482 (N_4482,N_3282,N_3273);
and U4483 (N_4483,N_2737,N_3400);
nand U4484 (N_4484,N_3211,N_3840);
nand U4485 (N_4485,N_3186,N_3439);
xor U4486 (N_4486,N_2964,N_2178);
or U4487 (N_4487,N_3607,N_2033);
nand U4488 (N_4488,N_3832,N_2272);
and U4489 (N_4489,N_3006,N_2048);
nand U4490 (N_4490,N_3497,N_2978);
nand U4491 (N_4491,N_2915,N_3334);
or U4492 (N_4492,N_3829,N_3673);
and U4493 (N_4493,N_2996,N_2891);
and U4494 (N_4494,N_3986,N_2788);
and U4495 (N_4495,N_3693,N_2514);
and U4496 (N_4496,N_2859,N_2361);
xnor U4497 (N_4497,N_3284,N_3023);
or U4498 (N_4498,N_3170,N_2531);
nand U4499 (N_4499,N_3230,N_3145);
and U4500 (N_4500,N_2488,N_3674);
xor U4501 (N_4501,N_3949,N_2136);
and U4502 (N_4502,N_3550,N_3210);
or U4503 (N_4503,N_3902,N_2605);
nor U4504 (N_4504,N_2084,N_3737);
xor U4505 (N_4505,N_3793,N_2634);
or U4506 (N_4506,N_2138,N_3154);
and U4507 (N_4507,N_2854,N_3681);
nor U4508 (N_4508,N_2867,N_3421);
xor U4509 (N_4509,N_3401,N_2036);
nand U4510 (N_4510,N_3242,N_2685);
nand U4511 (N_4511,N_2330,N_2300);
and U4512 (N_4512,N_3325,N_2018);
and U4513 (N_4513,N_2352,N_3893);
xor U4514 (N_4514,N_2252,N_2201);
xnor U4515 (N_4515,N_3094,N_3187);
and U4516 (N_4516,N_2819,N_3441);
xnor U4517 (N_4517,N_3278,N_3399);
and U4518 (N_4518,N_2225,N_2273);
nand U4519 (N_4519,N_3157,N_2713);
nor U4520 (N_4520,N_2095,N_2551);
nor U4521 (N_4521,N_3886,N_3516);
or U4522 (N_4522,N_3303,N_2245);
xnor U4523 (N_4523,N_2673,N_3767);
and U4524 (N_4524,N_3785,N_2092);
or U4525 (N_4525,N_2243,N_2753);
nand U4526 (N_4526,N_2063,N_2423);
and U4527 (N_4527,N_2206,N_2172);
or U4528 (N_4528,N_3789,N_3971);
nand U4529 (N_4529,N_3911,N_3461);
xnor U4530 (N_4530,N_2552,N_3506);
nand U4531 (N_4531,N_2517,N_2446);
or U4532 (N_4532,N_3519,N_2745);
nor U4533 (N_4533,N_2645,N_2539);
or U4534 (N_4534,N_3937,N_2703);
nor U4535 (N_4535,N_2561,N_3746);
nand U4536 (N_4536,N_3214,N_2335);
or U4537 (N_4537,N_2697,N_3140);
nor U4538 (N_4538,N_2522,N_2202);
or U4539 (N_4539,N_2310,N_2527);
xor U4540 (N_4540,N_2472,N_2406);
nand U4541 (N_4541,N_3202,N_2071);
nor U4542 (N_4542,N_3407,N_3431);
nor U4543 (N_4543,N_2013,N_3524);
and U4544 (N_4544,N_2839,N_3067);
xor U4545 (N_4545,N_2251,N_2102);
or U4546 (N_4546,N_3672,N_3711);
or U4547 (N_4547,N_3500,N_3351);
xor U4548 (N_4548,N_2941,N_3430);
and U4549 (N_4549,N_2504,N_2727);
nor U4550 (N_4550,N_2575,N_2958);
xor U4551 (N_4551,N_2123,N_3874);
nand U4552 (N_4552,N_2059,N_2715);
and U4553 (N_4553,N_3970,N_3138);
or U4554 (N_4554,N_2415,N_3589);
nor U4555 (N_4555,N_3326,N_3724);
or U4556 (N_4556,N_3036,N_3858);
and U4557 (N_4557,N_3473,N_2932);
xnor U4558 (N_4558,N_3851,N_2600);
and U4559 (N_4559,N_2807,N_3802);
nand U4560 (N_4560,N_3517,N_2750);
xor U4561 (N_4561,N_2914,N_2676);
and U4562 (N_4562,N_2519,N_2087);
or U4563 (N_4563,N_3104,N_3606);
or U4564 (N_4564,N_3007,N_3837);
and U4565 (N_4565,N_2776,N_2717);
nor U4566 (N_4566,N_3176,N_3127);
or U4567 (N_4567,N_2628,N_3133);
and U4568 (N_4568,N_2442,N_3615);
xor U4569 (N_4569,N_3476,N_2949);
nand U4570 (N_4570,N_2139,N_2662);
or U4571 (N_4571,N_2708,N_3910);
nand U4572 (N_4572,N_3826,N_2808);
nand U4573 (N_4573,N_3366,N_2821);
nand U4574 (N_4574,N_3375,N_3184);
xor U4575 (N_4575,N_3388,N_3397);
nor U4576 (N_4576,N_3679,N_3935);
and U4577 (N_4577,N_3235,N_2735);
nand U4578 (N_4578,N_3122,N_3978);
xor U4579 (N_4579,N_3618,N_2910);
nor U4580 (N_4580,N_3166,N_3245);
xor U4581 (N_4581,N_2668,N_2170);
and U4582 (N_4582,N_2987,N_3488);
or U4583 (N_4583,N_3196,N_3709);
xor U4584 (N_4584,N_2936,N_2688);
or U4585 (N_4585,N_2956,N_3136);
and U4586 (N_4586,N_2800,N_2916);
and U4587 (N_4587,N_3420,N_3066);
nand U4588 (N_4588,N_3751,N_2773);
nand U4589 (N_4589,N_3382,N_3879);
or U4590 (N_4590,N_3768,N_3259);
or U4591 (N_4591,N_2789,N_2664);
or U4592 (N_4592,N_3749,N_2115);
nor U4593 (N_4593,N_2626,N_3532);
nand U4594 (N_4594,N_2349,N_2370);
and U4595 (N_4595,N_2261,N_3546);
or U4596 (N_4596,N_3485,N_3698);
xor U4597 (N_4597,N_2840,N_3323);
nand U4598 (N_4598,N_3579,N_3346);
xnor U4599 (N_4599,N_3967,N_2067);
xor U4600 (N_4600,N_3630,N_3962);
nand U4601 (N_4601,N_2702,N_3099);
and U4602 (N_4602,N_2579,N_3769);
nand U4603 (N_4603,N_2309,N_3252);
nor U4604 (N_4604,N_2640,N_3153);
xor U4605 (N_4605,N_3695,N_2317);
nand U4606 (N_4606,N_3958,N_3251);
nor U4607 (N_4607,N_2995,N_3132);
or U4608 (N_4608,N_2440,N_3298);
xor U4609 (N_4609,N_2326,N_2836);
and U4610 (N_4610,N_2726,N_3429);
xor U4611 (N_4611,N_3804,N_2530);
and U4612 (N_4612,N_3694,N_2389);
nor U4613 (N_4613,N_2521,N_2816);
xnor U4614 (N_4614,N_2236,N_2331);
nand U4615 (N_4615,N_3229,N_3570);
and U4616 (N_4616,N_2746,N_3661);
and U4617 (N_4617,N_2182,N_3020);
xnor U4618 (N_4618,N_2105,N_2432);
or U4619 (N_4619,N_3941,N_2653);
nor U4620 (N_4620,N_2108,N_3581);
nor U4621 (N_4621,N_2291,N_3738);
or U4622 (N_4622,N_2449,N_2609);
nor U4623 (N_4623,N_2347,N_2295);
xor U4624 (N_4624,N_2644,N_2516);
nor U4625 (N_4625,N_2112,N_3521);
and U4626 (N_4626,N_2637,N_3787);
or U4627 (N_4627,N_2168,N_2968);
or U4628 (N_4628,N_3428,N_2345);
nor U4629 (N_4629,N_2340,N_2935);
nor U4630 (N_4630,N_2489,N_2313);
xnor U4631 (N_4631,N_2961,N_2068);
and U4632 (N_4632,N_3293,N_3904);
or U4633 (N_4633,N_3457,N_2707);
and U4634 (N_4634,N_2040,N_3587);
nand U4635 (N_4635,N_3525,N_2679);
and U4636 (N_4636,N_3223,N_2399);
nor U4637 (N_4637,N_2262,N_3729);
and U4638 (N_4638,N_2748,N_2556);
nor U4639 (N_4639,N_2831,N_2542);
xor U4640 (N_4640,N_3973,N_2420);
xnor U4641 (N_4641,N_2157,N_2100);
xor U4642 (N_4642,N_2906,N_3477);
xnor U4643 (N_4643,N_3482,N_3335);
or U4644 (N_4644,N_3356,N_3150);
or U4645 (N_4645,N_2681,N_3075);
and U4646 (N_4646,N_3651,N_2795);
or U4647 (N_4647,N_3033,N_2165);
xor U4648 (N_4648,N_3922,N_3188);
nor U4649 (N_4649,N_3014,N_2829);
nor U4650 (N_4650,N_3010,N_2714);
or U4651 (N_4651,N_2496,N_2458);
nor U4652 (N_4652,N_3867,N_2316);
xnor U4653 (N_4653,N_2025,N_2344);
xor U4654 (N_4654,N_3316,N_2657);
or U4655 (N_4655,N_3022,N_3827);
xor U4656 (N_4656,N_2853,N_3803);
or U4657 (N_4657,N_3513,N_2382);
nand U4658 (N_4658,N_2777,N_2909);
and U4659 (N_4659,N_2119,N_3423);
xnor U4660 (N_4660,N_3722,N_2754);
and U4661 (N_4661,N_2177,N_3304);
or U4662 (N_4662,N_2376,N_3354);
and U4663 (N_4663,N_2280,N_3215);
and U4664 (N_4664,N_3129,N_3713);
xnor U4665 (N_4665,N_3172,N_2716);
and U4666 (N_4666,N_3042,N_2596);
xor U4667 (N_4667,N_3818,N_2367);
nor U4668 (N_4668,N_3197,N_2266);
xor U4669 (N_4669,N_2358,N_2043);
and U4670 (N_4670,N_2659,N_2368);
xor U4671 (N_4671,N_2306,N_2341);
xnor U4672 (N_4672,N_2336,N_3509);
nand U4673 (N_4673,N_3948,N_3489);
or U4674 (N_4674,N_3106,N_2775);
and U4675 (N_4675,N_2354,N_3932);
nor U4676 (N_4676,N_3889,N_3155);
xor U4677 (N_4677,N_2541,N_2888);
nand U4678 (N_4678,N_2122,N_3834);
xnor U4679 (N_4679,N_2072,N_2413);
nor U4680 (N_4680,N_2038,N_2431);
xnor U4681 (N_4681,N_3212,N_3582);
xnor U4682 (N_4682,N_3575,N_2480);
nand U4683 (N_4683,N_3706,N_2075);
xor U4684 (N_4684,N_3936,N_2954);
and U4685 (N_4685,N_2782,N_3956);
or U4686 (N_4686,N_3160,N_2734);
or U4687 (N_4687,N_3881,N_2736);
nand U4688 (N_4688,N_3836,N_2267);
or U4689 (N_4689,N_2099,N_3435);
and U4690 (N_4690,N_3975,N_2638);
xnor U4691 (N_4691,N_2969,N_2842);
and U4692 (N_4692,N_2294,N_3387);
nand U4693 (N_4693,N_2184,N_2610);
nand U4694 (N_4694,N_3545,N_3599);
and U4695 (N_4695,N_3128,N_3294);
nand U4696 (N_4696,N_2985,N_2328);
xnor U4697 (N_4697,N_3675,N_3708);
and U4698 (N_4698,N_3434,N_2938);
xnor U4699 (N_4699,N_3297,N_3880);
nand U4700 (N_4700,N_3253,N_3353);
xnor U4701 (N_4701,N_3291,N_3416);
nor U4702 (N_4702,N_2823,N_3632);
and U4703 (N_4703,N_3227,N_2057);
and U4704 (N_4704,N_3998,N_3742);
nor U4705 (N_4705,N_3073,N_3842);
nor U4706 (N_4706,N_3946,N_2981);
nor U4707 (N_4707,N_2786,N_3433);
or U4708 (N_4708,N_2546,N_3377);
or U4709 (N_4709,N_2269,N_2523);
nor U4710 (N_4710,N_3976,N_2554);
nand U4711 (N_4711,N_3655,N_3365);
and U4712 (N_4712,N_3285,N_3730);
nor U4713 (N_4713,N_3169,N_2810);
or U4714 (N_4714,N_3444,N_3028);
nor U4715 (N_4715,N_2686,N_2655);
nand U4716 (N_4716,N_3008,N_3328);
xor U4717 (N_4717,N_2817,N_2460);
xor U4718 (N_4718,N_2863,N_3643);
or U4719 (N_4719,N_3396,N_2774);
and U4720 (N_4720,N_3241,N_2771);
nor U4721 (N_4721,N_3092,N_2186);
or U4722 (N_4722,N_3483,N_2337);
nand U4723 (N_4723,N_3849,N_3333);
nand U4724 (N_4724,N_3466,N_3034);
or U4725 (N_4725,N_3339,N_2073);
or U4726 (N_4726,N_3258,N_2339);
xnor U4727 (N_4727,N_3601,N_2592);
nor U4728 (N_4728,N_2894,N_2547);
or U4729 (N_4729,N_2545,N_2700);
or U4730 (N_4730,N_2014,N_2191);
or U4731 (N_4731,N_3717,N_3913);
nor U4732 (N_4732,N_3357,N_3037);
nor U4733 (N_4733,N_2474,N_2438);
nor U4734 (N_4734,N_2158,N_2457);
nor U4735 (N_4735,N_2641,N_2118);
or U4736 (N_4736,N_3144,N_3621);
nor U4737 (N_4737,N_2725,N_2604);
nor U4738 (N_4738,N_3363,N_3678);
and U4739 (N_4739,N_2560,N_3638);
nor U4740 (N_4740,N_3179,N_3850);
nand U4741 (N_4741,N_3452,N_3989);
or U4742 (N_4742,N_2060,N_3704);
or U4743 (N_4743,N_2701,N_3584);
and U4744 (N_4744,N_3572,N_3779);
xnor U4745 (N_4745,N_2719,N_3370);
and U4746 (N_4746,N_3277,N_2011);
xor U4747 (N_4747,N_2189,N_2639);
nor U4748 (N_4748,N_3600,N_3054);
and U4749 (N_4749,N_3993,N_3625);
or U4750 (N_4750,N_3752,N_2209);
and U4751 (N_4751,N_3064,N_2878);
and U4752 (N_4752,N_3274,N_3338);
or U4753 (N_4753,N_3512,N_2830);
xnor U4754 (N_4754,N_2463,N_2066);
xor U4755 (N_4755,N_3490,N_2723);
nand U4756 (N_4756,N_3467,N_2513);
xnor U4757 (N_4757,N_3915,N_2710);
nor U4758 (N_4758,N_3920,N_3078);
and U4759 (N_4759,N_3134,N_2532);
nand U4760 (N_4760,N_3931,N_3355);
xor U4761 (N_4761,N_2841,N_3208);
nor U4762 (N_4762,N_2045,N_3358);
and U4763 (N_4763,N_3885,N_3918);
or U4764 (N_4764,N_3168,N_3105);
and U4765 (N_4765,N_3376,N_3938);
nand U4766 (N_4766,N_2544,N_2654);
xor U4767 (N_4767,N_3445,N_2001);
nand U4768 (N_4768,N_2156,N_2462);
xnor U4769 (N_4769,N_2756,N_2536);
xor U4770 (N_4770,N_3716,N_3758);
nand U4771 (N_4771,N_3817,N_2289);
nand U4772 (N_4772,N_3009,N_2035);
nor U4773 (N_4773,N_2876,N_3743);
nor U4774 (N_4774,N_3447,N_2031);
nor U4775 (N_4775,N_3529,N_3943);
xnor U4776 (N_4776,N_2020,N_2471);
and U4777 (N_4777,N_2680,N_2477);
nand U4778 (N_4778,N_2926,N_2797);
nand U4779 (N_4779,N_2321,N_2140);
nor U4780 (N_4780,N_2375,N_2002);
xor U4781 (N_4781,N_3244,N_2132);
and U4782 (N_4782,N_3860,N_3432);
nor U4783 (N_4783,N_3750,N_3057);
nor U4784 (N_4784,N_2705,N_2799);
nand U4785 (N_4785,N_2809,N_3685);
and U4786 (N_4786,N_2597,N_3295);
or U4787 (N_4787,N_3542,N_2722);
xor U4788 (N_4788,N_3369,N_3171);
or U4789 (N_4789,N_3219,N_2264);
nor U4790 (N_4790,N_3624,N_3112);
nor U4791 (N_4791,N_2447,N_2928);
or U4792 (N_4792,N_3996,N_3493);
xnor U4793 (N_4793,N_3939,N_3070);
nand U4794 (N_4794,N_3048,N_2333);
xor U4795 (N_4795,N_3777,N_2643);
xnor U4796 (N_4796,N_2479,N_3003);
and U4797 (N_4797,N_3289,N_3964);
or U4798 (N_4798,N_3359,N_3539);
and U4799 (N_4799,N_3875,N_3190);
nor U4800 (N_4800,N_3552,N_2883);
and U4801 (N_4801,N_3957,N_2373);
or U4802 (N_4802,N_2296,N_3926);
nand U4803 (N_4803,N_3246,N_2228);
and U4804 (N_4804,N_3830,N_3107);
xor U4805 (N_4805,N_3865,N_3098);
nor U4806 (N_4806,N_3225,N_2176);
and U4807 (N_4807,N_3617,N_2149);
xor U4808 (N_4808,N_3748,N_3639);
nor U4809 (N_4809,N_2199,N_3120);
nand U4810 (N_4810,N_2395,N_3611);
and U4811 (N_4811,N_3206,N_3814);
and U4812 (N_4812,N_2127,N_2856);
xor U4813 (N_4813,N_3426,N_2456);
nor U4814 (N_4814,N_3419,N_2010);
nor U4815 (N_4815,N_3103,N_3712);
xnor U4816 (N_4816,N_3049,N_2409);
xnor U4817 (N_4817,N_2520,N_3691);
nor U4818 (N_4818,N_3985,N_3504);
xor U4819 (N_4819,N_3536,N_2461);
and U4820 (N_4820,N_2124,N_3727);
xnor U4821 (N_4821,N_3895,N_2793);
nor U4822 (N_4822,N_3058,N_3728);
or U4823 (N_4823,N_3256,N_3045);
or U4824 (N_4824,N_3612,N_3348);
or U4825 (N_4825,N_2203,N_2253);
xor U4826 (N_4826,N_2250,N_2882);
nor U4827 (N_4827,N_2769,N_3378);
nand U4828 (N_4828,N_3518,N_2525);
nand U4829 (N_4829,N_3044,N_2314);
and U4830 (N_4830,N_2107,N_2762);
nor U4831 (N_4831,N_3796,N_2744);
xnor U4832 (N_4832,N_3583,N_3969);
and U4833 (N_4833,N_3076,N_3181);
or U4834 (N_4834,N_3676,N_2584);
or U4835 (N_4835,N_3854,N_2424);
nand U4836 (N_4836,N_2674,N_3692);
nand U4837 (N_4837,N_2997,N_2721);
nand U4838 (N_4838,N_2908,N_3408);
nand U4839 (N_4839,N_2265,N_2612);
nand U4840 (N_4840,N_3101,N_3386);
or U4841 (N_4841,N_2718,N_3218);
nand U4842 (N_4842,N_2616,N_3610);
nor U4843 (N_4843,N_2387,N_3805);
nand U4844 (N_4844,N_2787,N_2481);
nor U4845 (N_4845,N_3405,N_3686);
xor U4846 (N_4846,N_2079,N_2660);
xor U4847 (N_4847,N_3224,N_2083);
and U4848 (N_4848,N_2301,N_3870);
nor U4849 (N_4849,N_2223,N_3047);
nor U4850 (N_4850,N_2129,N_2709);
and U4851 (N_4851,N_2473,N_3963);
nor U4852 (N_4852,N_3288,N_2687);
nor U4853 (N_4853,N_2388,N_3380);
nand U4854 (N_4854,N_2356,N_3292);
and U4855 (N_4855,N_3689,N_2275);
xnor U4856 (N_4856,N_3404,N_2383);
or U4857 (N_4857,N_3119,N_2374);
nand U4858 (N_4858,N_3591,N_2999);
or U4859 (N_4859,N_3634,N_3364);
nor U4860 (N_4860,N_2195,N_2454);
nor U4861 (N_4861,N_3510,N_2110);
xnor U4862 (N_4862,N_2511,N_3233);
and U4863 (N_4863,N_2814,N_3590);
xor U4864 (N_4864,N_2994,N_3373);
and U4865 (N_4865,N_3930,N_3636);
nor U4866 (N_4866,N_2334,N_3955);
nor U4867 (N_4867,N_3247,N_2772);
and U4868 (N_4868,N_3968,N_3418);
and U4869 (N_4869,N_3200,N_2562);
nand U4870 (N_4870,N_2391,N_2220);
nand U4871 (N_4871,N_2007,N_2090);
xnor U4872 (N_4872,N_3563,N_3592);
xnor U4873 (N_4873,N_2263,N_3053);
nand U4874 (N_4874,N_2231,N_3178);
and U4875 (N_4875,N_2899,N_3987);
nand U4876 (N_4876,N_2405,N_3065);
nor U4877 (N_4877,N_3312,N_2081);
or U4878 (N_4878,N_3125,N_3596);
nand U4879 (N_4879,N_3313,N_2647);
and U4880 (N_4880,N_3531,N_3013);
nor U4881 (N_4881,N_2515,N_2989);
and U4882 (N_4882,N_3526,N_3573);
xor U4883 (N_4883,N_3864,N_2794);
nor U4884 (N_4884,N_2733,N_2975);
or U4885 (N_4885,N_2412,N_3156);
or U4886 (N_4886,N_3974,N_3237);
nor U4887 (N_4887,N_2378,N_3089);
or U4888 (N_4888,N_2615,N_2785);
or U4889 (N_4889,N_3389,N_3761);
nor U4890 (N_4890,N_2905,N_3540);
nand U4891 (N_4891,N_3794,N_3909);
nand U4892 (N_4892,N_3914,N_3436);
nor U4893 (N_4893,N_3032,N_3026);
nor U4894 (N_4894,N_2933,N_3102);
and U4895 (N_4895,N_3680,N_3578);
xnor U4896 (N_4896,N_2397,N_3422);
xor U4897 (N_4897,N_2386,N_2276);
nand U4898 (N_4898,N_3961,N_2646);
or U4899 (N_4899,N_3159,N_2927);
xnor U4900 (N_4900,N_3831,N_3031);
nand U4901 (N_4901,N_3528,N_2144);
and U4902 (N_4902,N_3645,N_2348);
and U4903 (N_4903,N_2398,N_2570);
nor U4904 (N_4904,N_2766,N_3276);
or U4905 (N_4905,N_2872,N_3808);
xor U4906 (N_4906,N_2825,N_3379);
xor U4907 (N_4907,N_3890,N_2077);
xnor U4908 (N_4908,N_2311,N_3413);
and U4909 (N_4909,N_2041,N_2897);
and U4910 (N_4910,N_3097,N_2533);
nand U4911 (N_4911,N_2085,N_2608);
nand U4912 (N_4912,N_2312,N_3569);
or U4913 (N_4913,N_3458,N_3505);
nor U4914 (N_4914,N_2180,N_2282);
xor U4915 (N_4915,N_3460,N_3899);
nand U4916 (N_4916,N_2435,N_2363);
nand U4917 (N_4917,N_2393,N_3861);
and U4918 (N_4918,N_3412,N_2193);
xnor U4919 (N_4919,N_3096,N_2004);
or U4920 (N_4920,N_3347,N_3983);
or U4921 (N_4921,N_2305,N_2558);
nand U4922 (N_4922,N_3725,N_2061);
xor U4923 (N_4923,N_3774,N_2728);
nor U4924 (N_4924,N_3602,N_3807);
nand U4925 (N_4925,N_3892,N_3723);
or U4926 (N_4926,N_2528,N_3114);
or U4927 (N_4927,N_2381,N_2990);
nand U4928 (N_4928,N_2351,N_2155);
nor U4929 (N_4929,N_2065,N_2318);
xor U4930 (N_4930,N_3222,N_2298);
xnor U4931 (N_4931,N_3562,N_2631);
nor U4932 (N_4932,N_2851,N_3585);
nor U4933 (N_4933,N_3816,N_3784);
xnor U4934 (N_4934,N_2636,N_2450);
and U4935 (N_4935,N_3481,N_2572);
and U4936 (N_4936,N_2464,N_2302);
nor U4937 (N_4937,N_2362,N_2235);
and U4938 (N_4938,N_3537,N_2003);
or U4939 (N_4939,N_2959,N_2497);
or U4940 (N_4940,N_3586,N_2550);
and U4941 (N_4941,N_3703,N_3644);
xor U4942 (N_4942,N_3142,N_3449);
xnor U4943 (N_4943,N_2632,N_2704);
and U4944 (N_4944,N_3468,N_2566);
nor U4945 (N_4945,N_3907,N_2813);
or U4946 (N_4946,N_2130,N_3786);
and U4947 (N_4947,N_2154,N_2058);
nor U4948 (N_4948,N_2833,N_3306);
or U4949 (N_4949,N_3015,N_2016);
nor U4950 (N_4950,N_2972,N_3745);
and U4951 (N_4951,N_2764,N_2101);
xnor U4952 (N_4952,N_2587,N_2161);
or U4953 (N_4953,N_3198,N_3564);
xor U4954 (N_4954,N_2862,N_3650);
xor U4955 (N_4955,N_3148,N_3271);
nor U4956 (N_4956,N_3942,N_3715);
and U4957 (N_4957,N_2732,N_2056);
or U4958 (N_4958,N_2360,N_3649);
nand U4959 (N_4959,N_2661,N_2160);
and U4960 (N_4960,N_3362,N_2346);
nand U4961 (N_4961,N_2082,N_3261);
or U4962 (N_4962,N_2088,N_3863);
xor U4963 (N_4963,N_2601,N_2690);
nor U4964 (N_4964,N_3921,N_2445);
nand U4965 (N_4965,N_3257,N_2988);
or U4966 (N_4966,N_3855,N_3613);
nor U4967 (N_4967,N_2493,N_2971);
xor U4968 (N_4968,N_2900,N_2884);
or U4969 (N_4969,N_3756,N_3100);
nor U4970 (N_4970,N_2868,N_2396);
or U4971 (N_4971,N_3116,N_3314);
xnor U4972 (N_4972,N_3062,N_3438);
or U4973 (N_4973,N_2873,N_2026);
nand U4974 (N_4974,N_2323,N_2502);
xor U4975 (N_4975,N_3656,N_2855);
nor U4976 (N_4976,N_2353,N_3797);
and U4977 (N_4977,N_3702,N_3740);
and U4978 (N_4978,N_3384,N_3442);
xnor U4979 (N_4979,N_3647,N_2216);
nor U4980 (N_4980,N_2484,N_2205);
nor U4981 (N_4981,N_2164,N_2006);
nand U4982 (N_4982,N_3835,N_2619);
and U4983 (N_4983,N_3534,N_3734);
and U4984 (N_4984,N_2752,N_2948);
or U4985 (N_4985,N_3162,N_3912);
nor U4986 (N_4986,N_2564,N_2355);
nor U4987 (N_4987,N_3248,N_3381);
and U4988 (N_4988,N_3559,N_2577);
and U4989 (N_4989,N_2980,N_3852);
nand U4990 (N_4990,N_2485,N_3318);
nor U4991 (N_4991,N_2222,N_2973);
nor U4992 (N_4992,N_3177,N_3319);
or U4993 (N_4993,N_3538,N_2879);
or U4994 (N_4994,N_3164,N_2468);
or U4995 (N_4995,N_2706,N_2021);
nand U4996 (N_4996,N_3275,N_3782);
xor U4997 (N_4997,N_2911,N_2439);
and U4998 (N_4998,N_2974,N_3825);
or U4999 (N_4999,N_3496,N_3327);
xnor U5000 (N_5000,N_2021,N_2803);
nand U5001 (N_5001,N_2131,N_3401);
nand U5002 (N_5002,N_2271,N_3527);
nand U5003 (N_5003,N_2693,N_3999);
nand U5004 (N_5004,N_2176,N_3063);
nand U5005 (N_5005,N_2560,N_2921);
nand U5006 (N_5006,N_3732,N_3874);
or U5007 (N_5007,N_2669,N_3938);
xnor U5008 (N_5008,N_2927,N_2733);
nor U5009 (N_5009,N_3818,N_3695);
xor U5010 (N_5010,N_2954,N_2756);
nand U5011 (N_5011,N_2794,N_3576);
nor U5012 (N_5012,N_2391,N_3999);
or U5013 (N_5013,N_3652,N_3854);
or U5014 (N_5014,N_2806,N_3786);
xor U5015 (N_5015,N_2871,N_3411);
nor U5016 (N_5016,N_3303,N_2867);
and U5017 (N_5017,N_2873,N_3559);
or U5018 (N_5018,N_3763,N_2893);
xor U5019 (N_5019,N_3891,N_2524);
nor U5020 (N_5020,N_2283,N_3394);
xor U5021 (N_5021,N_2486,N_3225);
or U5022 (N_5022,N_2811,N_2493);
or U5023 (N_5023,N_2096,N_2781);
xor U5024 (N_5024,N_3151,N_2260);
nand U5025 (N_5025,N_2185,N_3685);
or U5026 (N_5026,N_3143,N_3343);
nand U5027 (N_5027,N_2208,N_2830);
nand U5028 (N_5028,N_3675,N_3042);
xor U5029 (N_5029,N_2297,N_2103);
nor U5030 (N_5030,N_3325,N_3129);
and U5031 (N_5031,N_2643,N_3143);
or U5032 (N_5032,N_3216,N_2776);
or U5033 (N_5033,N_3803,N_2717);
and U5034 (N_5034,N_3732,N_2265);
nor U5035 (N_5035,N_2842,N_2497);
and U5036 (N_5036,N_2634,N_2466);
nand U5037 (N_5037,N_3689,N_3429);
nor U5038 (N_5038,N_2610,N_3310);
nand U5039 (N_5039,N_3147,N_3447);
nand U5040 (N_5040,N_2334,N_3914);
nand U5041 (N_5041,N_2002,N_2647);
or U5042 (N_5042,N_3350,N_3542);
nand U5043 (N_5043,N_3968,N_3062);
xnor U5044 (N_5044,N_2997,N_2943);
nand U5045 (N_5045,N_2827,N_2784);
or U5046 (N_5046,N_2909,N_2414);
nand U5047 (N_5047,N_3909,N_2605);
xnor U5048 (N_5048,N_3086,N_3825);
nand U5049 (N_5049,N_2436,N_2262);
nor U5050 (N_5050,N_3034,N_3127);
nor U5051 (N_5051,N_2714,N_2054);
and U5052 (N_5052,N_2062,N_2470);
xnor U5053 (N_5053,N_3666,N_2063);
nor U5054 (N_5054,N_2669,N_2709);
and U5055 (N_5055,N_3953,N_2670);
nor U5056 (N_5056,N_2701,N_3326);
nor U5057 (N_5057,N_3491,N_3514);
or U5058 (N_5058,N_3070,N_3194);
nand U5059 (N_5059,N_2119,N_3405);
xor U5060 (N_5060,N_3164,N_3152);
xor U5061 (N_5061,N_2441,N_2207);
or U5062 (N_5062,N_2385,N_3712);
and U5063 (N_5063,N_3152,N_2570);
nor U5064 (N_5064,N_2628,N_3307);
or U5065 (N_5065,N_2753,N_3007);
and U5066 (N_5066,N_2536,N_3149);
or U5067 (N_5067,N_3881,N_3150);
or U5068 (N_5068,N_3067,N_3796);
and U5069 (N_5069,N_2655,N_3507);
or U5070 (N_5070,N_3231,N_2942);
nor U5071 (N_5071,N_3220,N_2428);
xnor U5072 (N_5072,N_3694,N_3986);
or U5073 (N_5073,N_2236,N_2177);
nand U5074 (N_5074,N_2364,N_2752);
nor U5075 (N_5075,N_3866,N_3285);
xnor U5076 (N_5076,N_3914,N_3650);
xnor U5077 (N_5077,N_2345,N_2196);
xor U5078 (N_5078,N_3284,N_2019);
or U5079 (N_5079,N_3907,N_3470);
nand U5080 (N_5080,N_3886,N_2693);
and U5081 (N_5081,N_2011,N_2547);
nor U5082 (N_5082,N_3122,N_2770);
nand U5083 (N_5083,N_2766,N_2246);
or U5084 (N_5084,N_3707,N_2040);
and U5085 (N_5085,N_2995,N_3461);
nor U5086 (N_5086,N_2572,N_2705);
nand U5087 (N_5087,N_2178,N_2821);
and U5088 (N_5088,N_2404,N_3650);
xor U5089 (N_5089,N_2296,N_2275);
or U5090 (N_5090,N_2848,N_3820);
nand U5091 (N_5091,N_3530,N_3748);
nand U5092 (N_5092,N_2762,N_3422);
nor U5093 (N_5093,N_2351,N_3948);
nor U5094 (N_5094,N_3875,N_3755);
xnor U5095 (N_5095,N_3034,N_3706);
and U5096 (N_5096,N_3114,N_3972);
nand U5097 (N_5097,N_3342,N_3957);
nor U5098 (N_5098,N_3143,N_3209);
or U5099 (N_5099,N_2414,N_3434);
xor U5100 (N_5100,N_3934,N_3963);
nand U5101 (N_5101,N_2738,N_2817);
xor U5102 (N_5102,N_2441,N_2657);
nand U5103 (N_5103,N_3380,N_3939);
xor U5104 (N_5104,N_3586,N_3489);
nor U5105 (N_5105,N_2062,N_2785);
or U5106 (N_5106,N_3420,N_2912);
nand U5107 (N_5107,N_2466,N_2118);
nor U5108 (N_5108,N_2635,N_2805);
xor U5109 (N_5109,N_3222,N_2347);
and U5110 (N_5110,N_3275,N_3945);
nand U5111 (N_5111,N_3479,N_2025);
xnor U5112 (N_5112,N_2357,N_3390);
and U5113 (N_5113,N_3353,N_3119);
or U5114 (N_5114,N_3974,N_3402);
nor U5115 (N_5115,N_2042,N_2971);
nor U5116 (N_5116,N_3272,N_3217);
and U5117 (N_5117,N_2433,N_3512);
or U5118 (N_5118,N_2950,N_2340);
nor U5119 (N_5119,N_2830,N_2886);
and U5120 (N_5120,N_3149,N_3860);
and U5121 (N_5121,N_2776,N_2349);
or U5122 (N_5122,N_2822,N_2139);
xor U5123 (N_5123,N_3098,N_3983);
nor U5124 (N_5124,N_2940,N_2943);
nor U5125 (N_5125,N_2004,N_2397);
or U5126 (N_5126,N_2724,N_2395);
xnor U5127 (N_5127,N_2277,N_2306);
or U5128 (N_5128,N_2549,N_3456);
or U5129 (N_5129,N_3121,N_3546);
nand U5130 (N_5130,N_3502,N_2414);
and U5131 (N_5131,N_3799,N_3559);
nand U5132 (N_5132,N_2827,N_3642);
or U5133 (N_5133,N_2743,N_3122);
and U5134 (N_5134,N_2143,N_3071);
or U5135 (N_5135,N_2908,N_3696);
and U5136 (N_5136,N_2362,N_3612);
and U5137 (N_5137,N_2751,N_3940);
nor U5138 (N_5138,N_3797,N_2940);
nor U5139 (N_5139,N_2592,N_3452);
and U5140 (N_5140,N_2512,N_3563);
and U5141 (N_5141,N_3771,N_3016);
and U5142 (N_5142,N_3827,N_2633);
nand U5143 (N_5143,N_2569,N_3379);
or U5144 (N_5144,N_3422,N_2710);
and U5145 (N_5145,N_2760,N_3226);
nor U5146 (N_5146,N_2188,N_3851);
xor U5147 (N_5147,N_2663,N_3138);
and U5148 (N_5148,N_3307,N_2430);
nand U5149 (N_5149,N_2305,N_2805);
or U5150 (N_5150,N_2860,N_2311);
or U5151 (N_5151,N_2077,N_2254);
or U5152 (N_5152,N_2075,N_3372);
and U5153 (N_5153,N_2159,N_2981);
xnor U5154 (N_5154,N_2287,N_2995);
nand U5155 (N_5155,N_2435,N_3817);
or U5156 (N_5156,N_3382,N_2046);
and U5157 (N_5157,N_3081,N_2250);
nand U5158 (N_5158,N_3991,N_3765);
or U5159 (N_5159,N_3055,N_3849);
xor U5160 (N_5160,N_3384,N_2134);
nand U5161 (N_5161,N_2511,N_3133);
nand U5162 (N_5162,N_2715,N_3181);
xnor U5163 (N_5163,N_2583,N_2521);
or U5164 (N_5164,N_2610,N_3017);
or U5165 (N_5165,N_3711,N_2108);
xnor U5166 (N_5166,N_2348,N_3129);
nand U5167 (N_5167,N_3672,N_2625);
and U5168 (N_5168,N_2191,N_3980);
xor U5169 (N_5169,N_3187,N_3505);
and U5170 (N_5170,N_2155,N_2731);
or U5171 (N_5171,N_3118,N_2077);
nand U5172 (N_5172,N_3239,N_2241);
or U5173 (N_5173,N_3188,N_3046);
xnor U5174 (N_5174,N_2237,N_3992);
nand U5175 (N_5175,N_3067,N_3824);
nor U5176 (N_5176,N_2028,N_3832);
xnor U5177 (N_5177,N_3236,N_2935);
or U5178 (N_5178,N_3375,N_3944);
nand U5179 (N_5179,N_3309,N_3496);
or U5180 (N_5180,N_3130,N_2215);
and U5181 (N_5181,N_2001,N_2158);
nor U5182 (N_5182,N_2285,N_3138);
and U5183 (N_5183,N_2062,N_3784);
nand U5184 (N_5184,N_3027,N_2088);
xor U5185 (N_5185,N_3954,N_2279);
or U5186 (N_5186,N_2965,N_3194);
xor U5187 (N_5187,N_2829,N_3709);
or U5188 (N_5188,N_3383,N_2209);
xor U5189 (N_5189,N_3124,N_2019);
nor U5190 (N_5190,N_3271,N_2229);
xnor U5191 (N_5191,N_2718,N_2562);
and U5192 (N_5192,N_3293,N_2902);
nand U5193 (N_5193,N_2787,N_2520);
nand U5194 (N_5194,N_2140,N_3877);
or U5195 (N_5195,N_2772,N_3926);
or U5196 (N_5196,N_3614,N_3138);
nand U5197 (N_5197,N_3525,N_3885);
and U5198 (N_5198,N_3853,N_2532);
or U5199 (N_5199,N_2593,N_3563);
nor U5200 (N_5200,N_2815,N_2585);
nand U5201 (N_5201,N_2305,N_2532);
nor U5202 (N_5202,N_2467,N_2527);
nand U5203 (N_5203,N_3134,N_2949);
nand U5204 (N_5204,N_2576,N_2388);
and U5205 (N_5205,N_2563,N_3177);
or U5206 (N_5206,N_3568,N_2863);
nor U5207 (N_5207,N_3296,N_2863);
and U5208 (N_5208,N_2300,N_3607);
nor U5209 (N_5209,N_3860,N_3803);
nor U5210 (N_5210,N_2039,N_3862);
and U5211 (N_5211,N_2316,N_3712);
or U5212 (N_5212,N_2055,N_2113);
nand U5213 (N_5213,N_3458,N_2582);
nand U5214 (N_5214,N_3146,N_3395);
xor U5215 (N_5215,N_2366,N_3695);
and U5216 (N_5216,N_2596,N_2015);
xnor U5217 (N_5217,N_3032,N_3060);
nand U5218 (N_5218,N_2014,N_2551);
nand U5219 (N_5219,N_3640,N_2611);
and U5220 (N_5220,N_2417,N_2830);
and U5221 (N_5221,N_3935,N_2934);
xnor U5222 (N_5222,N_3327,N_3393);
xnor U5223 (N_5223,N_2371,N_3482);
nor U5224 (N_5224,N_2916,N_3714);
xnor U5225 (N_5225,N_3147,N_2566);
or U5226 (N_5226,N_3977,N_3382);
xor U5227 (N_5227,N_3912,N_2180);
nor U5228 (N_5228,N_3185,N_2908);
or U5229 (N_5229,N_3509,N_2618);
nor U5230 (N_5230,N_3990,N_3939);
nand U5231 (N_5231,N_3999,N_3567);
nand U5232 (N_5232,N_2084,N_2279);
and U5233 (N_5233,N_2023,N_2012);
nand U5234 (N_5234,N_2233,N_2427);
nor U5235 (N_5235,N_2464,N_3637);
nand U5236 (N_5236,N_3093,N_2156);
nand U5237 (N_5237,N_3055,N_2736);
and U5238 (N_5238,N_3039,N_2346);
nand U5239 (N_5239,N_3341,N_2088);
nand U5240 (N_5240,N_3170,N_2330);
xor U5241 (N_5241,N_3145,N_3532);
and U5242 (N_5242,N_2547,N_3482);
or U5243 (N_5243,N_2416,N_3854);
or U5244 (N_5244,N_2887,N_2144);
nor U5245 (N_5245,N_2578,N_3643);
nor U5246 (N_5246,N_3246,N_3824);
nand U5247 (N_5247,N_3083,N_3862);
xnor U5248 (N_5248,N_2057,N_3964);
xor U5249 (N_5249,N_3237,N_3072);
or U5250 (N_5250,N_2576,N_2789);
nand U5251 (N_5251,N_3140,N_3538);
nor U5252 (N_5252,N_2209,N_2050);
nand U5253 (N_5253,N_3312,N_3051);
or U5254 (N_5254,N_2921,N_2614);
nand U5255 (N_5255,N_2448,N_3466);
nor U5256 (N_5256,N_2941,N_3632);
xor U5257 (N_5257,N_3976,N_3322);
or U5258 (N_5258,N_2089,N_2774);
nor U5259 (N_5259,N_2488,N_3784);
nor U5260 (N_5260,N_3843,N_2912);
nor U5261 (N_5261,N_3176,N_2114);
nand U5262 (N_5262,N_3071,N_3861);
nand U5263 (N_5263,N_3509,N_3939);
and U5264 (N_5264,N_3738,N_2196);
nor U5265 (N_5265,N_3641,N_3788);
xnor U5266 (N_5266,N_2959,N_3747);
or U5267 (N_5267,N_2614,N_3681);
xor U5268 (N_5268,N_3324,N_2713);
or U5269 (N_5269,N_3368,N_2979);
and U5270 (N_5270,N_2872,N_3558);
xnor U5271 (N_5271,N_2485,N_3089);
nand U5272 (N_5272,N_2206,N_3607);
xor U5273 (N_5273,N_2567,N_2101);
or U5274 (N_5274,N_3941,N_2803);
and U5275 (N_5275,N_3497,N_2019);
or U5276 (N_5276,N_3347,N_3473);
nor U5277 (N_5277,N_3811,N_2174);
xnor U5278 (N_5278,N_2561,N_2017);
xnor U5279 (N_5279,N_3306,N_3660);
or U5280 (N_5280,N_3923,N_3834);
nor U5281 (N_5281,N_3042,N_2841);
xnor U5282 (N_5282,N_3687,N_3928);
xnor U5283 (N_5283,N_2817,N_2538);
xnor U5284 (N_5284,N_3217,N_2347);
and U5285 (N_5285,N_2341,N_2362);
nor U5286 (N_5286,N_3064,N_3589);
xnor U5287 (N_5287,N_3044,N_3166);
or U5288 (N_5288,N_3094,N_2951);
nand U5289 (N_5289,N_3479,N_3350);
xor U5290 (N_5290,N_3237,N_3170);
xnor U5291 (N_5291,N_2170,N_2444);
nand U5292 (N_5292,N_2046,N_2129);
and U5293 (N_5293,N_3187,N_2164);
and U5294 (N_5294,N_3217,N_2657);
and U5295 (N_5295,N_3335,N_2910);
and U5296 (N_5296,N_2865,N_2495);
nor U5297 (N_5297,N_3621,N_2010);
nor U5298 (N_5298,N_3854,N_3975);
nor U5299 (N_5299,N_2576,N_2478);
nor U5300 (N_5300,N_3575,N_2163);
nor U5301 (N_5301,N_2074,N_3155);
nor U5302 (N_5302,N_2700,N_3710);
or U5303 (N_5303,N_2864,N_2561);
nor U5304 (N_5304,N_2034,N_2330);
or U5305 (N_5305,N_3863,N_3998);
nor U5306 (N_5306,N_2545,N_2119);
xnor U5307 (N_5307,N_2968,N_2540);
or U5308 (N_5308,N_2829,N_3127);
nor U5309 (N_5309,N_3550,N_2210);
nand U5310 (N_5310,N_2433,N_3414);
xnor U5311 (N_5311,N_2386,N_2992);
nor U5312 (N_5312,N_3025,N_2846);
nand U5313 (N_5313,N_3904,N_3664);
xnor U5314 (N_5314,N_2184,N_3683);
or U5315 (N_5315,N_3978,N_2947);
nor U5316 (N_5316,N_3269,N_3993);
xor U5317 (N_5317,N_3476,N_3743);
nor U5318 (N_5318,N_3759,N_2958);
and U5319 (N_5319,N_3073,N_3950);
nand U5320 (N_5320,N_3419,N_3023);
or U5321 (N_5321,N_2059,N_3263);
or U5322 (N_5322,N_3945,N_3299);
xor U5323 (N_5323,N_3594,N_3712);
or U5324 (N_5324,N_3926,N_3054);
nor U5325 (N_5325,N_2811,N_2609);
or U5326 (N_5326,N_2474,N_2684);
nand U5327 (N_5327,N_3988,N_2634);
xnor U5328 (N_5328,N_3985,N_3474);
and U5329 (N_5329,N_3723,N_3463);
nand U5330 (N_5330,N_3197,N_3024);
xor U5331 (N_5331,N_2627,N_3766);
and U5332 (N_5332,N_3535,N_3527);
nand U5333 (N_5333,N_3247,N_2014);
or U5334 (N_5334,N_2806,N_3239);
xnor U5335 (N_5335,N_3649,N_2004);
nand U5336 (N_5336,N_3036,N_2207);
and U5337 (N_5337,N_3728,N_3977);
nor U5338 (N_5338,N_2171,N_2760);
or U5339 (N_5339,N_3244,N_3077);
nor U5340 (N_5340,N_2488,N_2287);
xor U5341 (N_5341,N_3953,N_2581);
xor U5342 (N_5342,N_2320,N_3895);
xnor U5343 (N_5343,N_2706,N_2275);
xor U5344 (N_5344,N_3727,N_2889);
nor U5345 (N_5345,N_3486,N_3363);
nand U5346 (N_5346,N_3211,N_2503);
xnor U5347 (N_5347,N_3792,N_3824);
or U5348 (N_5348,N_2329,N_3150);
nor U5349 (N_5349,N_3926,N_3913);
and U5350 (N_5350,N_2713,N_2740);
nand U5351 (N_5351,N_3546,N_2249);
or U5352 (N_5352,N_2344,N_2469);
xnor U5353 (N_5353,N_2018,N_3158);
xor U5354 (N_5354,N_3327,N_3186);
nand U5355 (N_5355,N_2826,N_2468);
or U5356 (N_5356,N_2919,N_3162);
nand U5357 (N_5357,N_2115,N_3662);
nand U5358 (N_5358,N_3965,N_2991);
and U5359 (N_5359,N_2641,N_2362);
nor U5360 (N_5360,N_3433,N_3746);
xor U5361 (N_5361,N_2667,N_2466);
xor U5362 (N_5362,N_2626,N_3963);
xor U5363 (N_5363,N_2708,N_2410);
xnor U5364 (N_5364,N_2729,N_3909);
nor U5365 (N_5365,N_2567,N_3020);
xor U5366 (N_5366,N_2137,N_2141);
nor U5367 (N_5367,N_2315,N_2599);
and U5368 (N_5368,N_3893,N_2402);
or U5369 (N_5369,N_2828,N_2515);
xor U5370 (N_5370,N_3852,N_3387);
and U5371 (N_5371,N_3798,N_3757);
nor U5372 (N_5372,N_3852,N_2647);
nor U5373 (N_5373,N_2589,N_2820);
and U5374 (N_5374,N_2839,N_3285);
nand U5375 (N_5375,N_3540,N_2102);
and U5376 (N_5376,N_3631,N_2384);
and U5377 (N_5377,N_2336,N_3536);
xor U5378 (N_5378,N_3834,N_3098);
or U5379 (N_5379,N_3774,N_2611);
and U5380 (N_5380,N_3951,N_2187);
xnor U5381 (N_5381,N_3801,N_2322);
xnor U5382 (N_5382,N_3477,N_2971);
or U5383 (N_5383,N_2169,N_2912);
nand U5384 (N_5384,N_3863,N_3444);
nor U5385 (N_5385,N_3896,N_2965);
or U5386 (N_5386,N_2469,N_3344);
or U5387 (N_5387,N_3396,N_2244);
nor U5388 (N_5388,N_2128,N_3484);
xor U5389 (N_5389,N_2108,N_3542);
or U5390 (N_5390,N_3598,N_2931);
or U5391 (N_5391,N_2080,N_3903);
or U5392 (N_5392,N_2593,N_2242);
nand U5393 (N_5393,N_3007,N_3138);
or U5394 (N_5394,N_2358,N_3060);
and U5395 (N_5395,N_2904,N_3035);
nor U5396 (N_5396,N_2541,N_3038);
nand U5397 (N_5397,N_3604,N_3681);
and U5398 (N_5398,N_3002,N_2315);
nand U5399 (N_5399,N_3196,N_3458);
or U5400 (N_5400,N_2366,N_2864);
nand U5401 (N_5401,N_3620,N_3799);
or U5402 (N_5402,N_3285,N_3664);
nor U5403 (N_5403,N_3957,N_2644);
nor U5404 (N_5404,N_3399,N_3612);
xnor U5405 (N_5405,N_2325,N_2078);
nand U5406 (N_5406,N_3115,N_2472);
xnor U5407 (N_5407,N_2502,N_2320);
or U5408 (N_5408,N_3271,N_2095);
and U5409 (N_5409,N_2460,N_2974);
or U5410 (N_5410,N_3997,N_3929);
or U5411 (N_5411,N_2982,N_2977);
nor U5412 (N_5412,N_2265,N_3052);
or U5413 (N_5413,N_2236,N_2382);
nor U5414 (N_5414,N_3708,N_2789);
or U5415 (N_5415,N_3928,N_2451);
or U5416 (N_5416,N_3732,N_3367);
or U5417 (N_5417,N_2970,N_2505);
and U5418 (N_5418,N_2224,N_3916);
or U5419 (N_5419,N_2774,N_2278);
nor U5420 (N_5420,N_2618,N_3256);
or U5421 (N_5421,N_3980,N_2349);
nor U5422 (N_5422,N_2074,N_3228);
xor U5423 (N_5423,N_3845,N_3890);
and U5424 (N_5424,N_3181,N_2735);
nand U5425 (N_5425,N_3914,N_3385);
and U5426 (N_5426,N_2925,N_3627);
nand U5427 (N_5427,N_2486,N_2645);
nand U5428 (N_5428,N_2258,N_3408);
nand U5429 (N_5429,N_3313,N_3254);
nand U5430 (N_5430,N_3951,N_3933);
nor U5431 (N_5431,N_2616,N_3604);
and U5432 (N_5432,N_3196,N_2413);
xnor U5433 (N_5433,N_2556,N_3188);
and U5434 (N_5434,N_3971,N_2078);
xnor U5435 (N_5435,N_3634,N_3488);
nor U5436 (N_5436,N_3497,N_2202);
nand U5437 (N_5437,N_2896,N_2979);
nor U5438 (N_5438,N_2489,N_3093);
and U5439 (N_5439,N_2410,N_3790);
or U5440 (N_5440,N_2038,N_3693);
and U5441 (N_5441,N_3173,N_2090);
and U5442 (N_5442,N_2903,N_2932);
and U5443 (N_5443,N_2767,N_2378);
xnor U5444 (N_5444,N_2646,N_3328);
and U5445 (N_5445,N_2798,N_3038);
or U5446 (N_5446,N_3873,N_2433);
nor U5447 (N_5447,N_3695,N_2671);
nor U5448 (N_5448,N_3753,N_3303);
or U5449 (N_5449,N_3953,N_2488);
xor U5450 (N_5450,N_2029,N_2064);
nand U5451 (N_5451,N_2104,N_3621);
nor U5452 (N_5452,N_2489,N_2749);
xnor U5453 (N_5453,N_3764,N_3309);
and U5454 (N_5454,N_3768,N_2862);
and U5455 (N_5455,N_2480,N_3974);
nor U5456 (N_5456,N_2069,N_2140);
nand U5457 (N_5457,N_3958,N_3695);
xnor U5458 (N_5458,N_2304,N_2039);
and U5459 (N_5459,N_2585,N_3092);
and U5460 (N_5460,N_2848,N_3736);
and U5461 (N_5461,N_2630,N_2390);
and U5462 (N_5462,N_2358,N_2570);
and U5463 (N_5463,N_3628,N_2929);
nand U5464 (N_5464,N_2688,N_2573);
xnor U5465 (N_5465,N_2907,N_3805);
xor U5466 (N_5466,N_3051,N_2694);
and U5467 (N_5467,N_3282,N_3219);
xor U5468 (N_5468,N_3691,N_2662);
or U5469 (N_5469,N_2067,N_2863);
nand U5470 (N_5470,N_3740,N_2734);
or U5471 (N_5471,N_2605,N_3325);
or U5472 (N_5472,N_3217,N_3860);
and U5473 (N_5473,N_3418,N_3500);
or U5474 (N_5474,N_3309,N_3021);
xor U5475 (N_5475,N_3298,N_3066);
nand U5476 (N_5476,N_2466,N_2121);
nand U5477 (N_5477,N_2285,N_3927);
and U5478 (N_5478,N_2637,N_2427);
or U5479 (N_5479,N_2280,N_2964);
or U5480 (N_5480,N_3335,N_2075);
nand U5481 (N_5481,N_2724,N_2620);
nor U5482 (N_5482,N_3044,N_2112);
nor U5483 (N_5483,N_2686,N_2222);
nand U5484 (N_5484,N_3817,N_2619);
nor U5485 (N_5485,N_2308,N_2373);
xor U5486 (N_5486,N_2474,N_2607);
nor U5487 (N_5487,N_3439,N_2242);
nand U5488 (N_5488,N_3577,N_3106);
xor U5489 (N_5489,N_3207,N_3377);
nor U5490 (N_5490,N_2757,N_2389);
xor U5491 (N_5491,N_3552,N_3767);
or U5492 (N_5492,N_2674,N_3669);
nand U5493 (N_5493,N_3822,N_2296);
xnor U5494 (N_5494,N_3247,N_3658);
nor U5495 (N_5495,N_2570,N_3194);
nor U5496 (N_5496,N_2152,N_3480);
nor U5497 (N_5497,N_3879,N_3072);
or U5498 (N_5498,N_3362,N_3111);
or U5499 (N_5499,N_3544,N_3765);
xnor U5500 (N_5500,N_2555,N_2601);
or U5501 (N_5501,N_2537,N_2578);
nor U5502 (N_5502,N_3368,N_2553);
nor U5503 (N_5503,N_3037,N_3360);
nor U5504 (N_5504,N_3607,N_2870);
nand U5505 (N_5505,N_2645,N_3456);
nor U5506 (N_5506,N_2343,N_3226);
and U5507 (N_5507,N_2042,N_3284);
nand U5508 (N_5508,N_3739,N_3578);
or U5509 (N_5509,N_3871,N_2272);
xnor U5510 (N_5510,N_3972,N_3522);
nand U5511 (N_5511,N_3401,N_2773);
or U5512 (N_5512,N_2935,N_3363);
or U5513 (N_5513,N_3429,N_2209);
nor U5514 (N_5514,N_2595,N_3132);
xnor U5515 (N_5515,N_2285,N_3454);
or U5516 (N_5516,N_3164,N_2259);
nand U5517 (N_5517,N_2523,N_3992);
nand U5518 (N_5518,N_3157,N_3327);
nand U5519 (N_5519,N_2037,N_3853);
nand U5520 (N_5520,N_3900,N_2880);
and U5521 (N_5521,N_2300,N_3850);
or U5522 (N_5522,N_2110,N_2269);
and U5523 (N_5523,N_3745,N_2102);
xnor U5524 (N_5524,N_2615,N_2410);
or U5525 (N_5525,N_2322,N_2415);
nor U5526 (N_5526,N_2209,N_3034);
nand U5527 (N_5527,N_3400,N_2208);
and U5528 (N_5528,N_2514,N_3313);
nand U5529 (N_5529,N_2786,N_2860);
or U5530 (N_5530,N_2982,N_2661);
or U5531 (N_5531,N_3994,N_2247);
nor U5532 (N_5532,N_3693,N_2950);
and U5533 (N_5533,N_3686,N_2896);
or U5534 (N_5534,N_2202,N_2219);
or U5535 (N_5535,N_3572,N_3287);
or U5536 (N_5536,N_2162,N_2441);
xor U5537 (N_5537,N_2080,N_3771);
and U5538 (N_5538,N_3748,N_2707);
and U5539 (N_5539,N_3203,N_3645);
nor U5540 (N_5540,N_2354,N_3744);
and U5541 (N_5541,N_2089,N_2519);
and U5542 (N_5542,N_2555,N_2149);
xor U5543 (N_5543,N_3509,N_3721);
and U5544 (N_5544,N_2528,N_2924);
xnor U5545 (N_5545,N_2648,N_3748);
nor U5546 (N_5546,N_3754,N_2697);
or U5547 (N_5547,N_2816,N_3327);
xor U5548 (N_5548,N_2921,N_3350);
nand U5549 (N_5549,N_3551,N_3725);
and U5550 (N_5550,N_2016,N_3997);
and U5551 (N_5551,N_3257,N_2332);
xor U5552 (N_5552,N_3867,N_3240);
or U5553 (N_5553,N_2205,N_2047);
nand U5554 (N_5554,N_2604,N_2481);
or U5555 (N_5555,N_3321,N_2305);
xnor U5556 (N_5556,N_2165,N_3508);
nor U5557 (N_5557,N_2166,N_2730);
xnor U5558 (N_5558,N_2235,N_2052);
and U5559 (N_5559,N_2805,N_3313);
and U5560 (N_5560,N_3720,N_2715);
or U5561 (N_5561,N_2945,N_3692);
or U5562 (N_5562,N_3530,N_3832);
nand U5563 (N_5563,N_2384,N_3219);
nor U5564 (N_5564,N_3640,N_3876);
xor U5565 (N_5565,N_3488,N_3612);
and U5566 (N_5566,N_2984,N_2517);
nor U5567 (N_5567,N_3179,N_3231);
and U5568 (N_5568,N_2303,N_2363);
or U5569 (N_5569,N_3882,N_2486);
nor U5570 (N_5570,N_2516,N_2816);
nand U5571 (N_5571,N_2357,N_2854);
nand U5572 (N_5572,N_3804,N_2192);
nor U5573 (N_5573,N_2461,N_3257);
xor U5574 (N_5574,N_2259,N_3992);
nand U5575 (N_5575,N_2431,N_3141);
xor U5576 (N_5576,N_3567,N_2582);
or U5577 (N_5577,N_3309,N_2445);
xnor U5578 (N_5578,N_2672,N_3324);
nor U5579 (N_5579,N_3667,N_3709);
or U5580 (N_5580,N_2831,N_3259);
and U5581 (N_5581,N_2703,N_2687);
and U5582 (N_5582,N_2462,N_2696);
nand U5583 (N_5583,N_2893,N_3499);
nor U5584 (N_5584,N_3507,N_2481);
nand U5585 (N_5585,N_3584,N_2240);
or U5586 (N_5586,N_3958,N_2896);
or U5587 (N_5587,N_3088,N_3707);
nor U5588 (N_5588,N_2022,N_2003);
and U5589 (N_5589,N_2709,N_3596);
nand U5590 (N_5590,N_3453,N_2952);
nor U5591 (N_5591,N_2471,N_3089);
nand U5592 (N_5592,N_2794,N_2823);
and U5593 (N_5593,N_3809,N_2497);
or U5594 (N_5594,N_2910,N_2103);
nor U5595 (N_5595,N_2925,N_2327);
nor U5596 (N_5596,N_2680,N_3742);
xor U5597 (N_5597,N_3989,N_2527);
xnor U5598 (N_5598,N_2476,N_2181);
nand U5599 (N_5599,N_2149,N_2129);
nor U5600 (N_5600,N_3512,N_3841);
xor U5601 (N_5601,N_2759,N_2113);
and U5602 (N_5602,N_3272,N_2824);
or U5603 (N_5603,N_2302,N_3397);
and U5604 (N_5604,N_2078,N_3032);
and U5605 (N_5605,N_2202,N_2727);
xnor U5606 (N_5606,N_3713,N_3470);
or U5607 (N_5607,N_3023,N_3302);
and U5608 (N_5608,N_2307,N_2221);
xor U5609 (N_5609,N_2217,N_3552);
xnor U5610 (N_5610,N_2785,N_2365);
or U5611 (N_5611,N_2704,N_2524);
xnor U5612 (N_5612,N_2069,N_2977);
nand U5613 (N_5613,N_3016,N_3602);
nor U5614 (N_5614,N_3923,N_3855);
and U5615 (N_5615,N_2474,N_3619);
and U5616 (N_5616,N_3619,N_2437);
or U5617 (N_5617,N_3955,N_2052);
nand U5618 (N_5618,N_2652,N_3461);
and U5619 (N_5619,N_2799,N_2347);
xnor U5620 (N_5620,N_2613,N_3565);
and U5621 (N_5621,N_2345,N_2601);
and U5622 (N_5622,N_2878,N_2112);
or U5623 (N_5623,N_3500,N_2604);
nand U5624 (N_5624,N_2624,N_2068);
or U5625 (N_5625,N_2880,N_2007);
nor U5626 (N_5626,N_2821,N_2779);
or U5627 (N_5627,N_3784,N_2669);
nor U5628 (N_5628,N_2013,N_2532);
and U5629 (N_5629,N_2101,N_2952);
xnor U5630 (N_5630,N_2451,N_2571);
nor U5631 (N_5631,N_2881,N_2410);
and U5632 (N_5632,N_2683,N_3502);
xor U5633 (N_5633,N_3590,N_2101);
nor U5634 (N_5634,N_3395,N_2453);
and U5635 (N_5635,N_2194,N_3763);
or U5636 (N_5636,N_3007,N_3539);
nand U5637 (N_5637,N_3192,N_2670);
or U5638 (N_5638,N_2967,N_3390);
nand U5639 (N_5639,N_3499,N_2278);
or U5640 (N_5640,N_3320,N_3256);
and U5641 (N_5641,N_3693,N_3127);
nand U5642 (N_5642,N_3599,N_2274);
and U5643 (N_5643,N_2044,N_2460);
or U5644 (N_5644,N_3258,N_2461);
xor U5645 (N_5645,N_2582,N_3254);
or U5646 (N_5646,N_3125,N_2794);
and U5647 (N_5647,N_3110,N_2414);
xnor U5648 (N_5648,N_2064,N_2362);
and U5649 (N_5649,N_2550,N_3529);
and U5650 (N_5650,N_2150,N_2064);
nor U5651 (N_5651,N_2581,N_2735);
or U5652 (N_5652,N_3042,N_2732);
nor U5653 (N_5653,N_2335,N_3427);
xor U5654 (N_5654,N_3627,N_3209);
nor U5655 (N_5655,N_2908,N_2459);
xnor U5656 (N_5656,N_3496,N_3016);
xor U5657 (N_5657,N_2747,N_2661);
nand U5658 (N_5658,N_2684,N_2391);
nor U5659 (N_5659,N_3025,N_3983);
xor U5660 (N_5660,N_2283,N_2995);
nand U5661 (N_5661,N_2993,N_3325);
or U5662 (N_5662,N_3730,N_3313);
and U5663 (N_5663,N_3589,N_2084);
or U5664 (N_5664,N_3194,N_3124);
nor U5665 (N_5665,N_3244,N_3389);
or U5666 (N_5666,N_3737,N_3082);
xnor U5667 (N_5667,N_2582,N_3554);
nand U5668 (N_5668,N_2893,N_2071);
nor U5669 (N_5669,N_2285,N_3239);
xnor U5670 (N_5670,N_2843,N_3848);
and U5671 (N_5671,N_2647,N_3194);
and U5672 (N_5672,N_3954,N_3923);
or U5673 (N_5673,N_3293,N_2948);
nor U5674 (N_5674,N_2238,N_3643);
nor U5675 (N_5675,N_2612,N_3626);
nor U5676 (N_5676,N_3432,N_3217);
or U5677 (N_5677,N_3499,N_2545);
nor U5678 (N_5678,N_2109,N_2613);
and U5679 (N_5679,N_2927,N_3338);
or U5680 (N_5680,N_3712,N_3376);
nor U5681 (N_5681,N_2612,N_3254);
xor U5682 (N_5682,N_2022,N_3278);
or U5683 (N_5683,N_2361,N_3597);
nor U5684 (N_5684,N_2012,N_2299);
and U5685 (N_5685,N_3198,N_3154);
xor U5686 (N_5686,N_3638,N_2753);
nand U5687 (N_5687,N_2235,N_2453);
and U5688 (N_5688,N_3014,N_2352);
nand U5689 (N_5689,N_2670,N_3907);
xor U5690 (N_5690,N_2724,N_3843);
nor U5691 (N_5691,N_3877,N_3635);
xnor U5692 (N_5692,N_3913,N_3643);
nor U5693 (N_5693,N_2060,N_2484);
nor U5694 (N_5694,N_3649,N_2434);
or U5695 (N_5695,N_2745,N_2465);
and U5696 (N_5696,N_3626,N_2978);
or U5697 (N_5697,N_2181,N_2359);
nor U5698 (N_5698,N_2378,N_2771);
or U5699 (N_5699,N_2929,N_3287);
or U5700 (N_5700,N_3477,N_2974);
and U5701 (N_5701,N_2504,N_2796);
xor U5702 (N_5702,N_3023,N_3726);
or U5703 (N_5703,N_3409,N_3798);
or U5704 (N_5704,N_2966,N_3718);
nand U5705 (N_5705,N_2641,N_3260);
nor U5706 (N_5706,N_3984,N_3454);
or U5707 (N_5707,N_3738,N_3387);
nand U5708 (N_5708,N_3248,N_2219);
xor U5709 (N_5709,N_2070,N_3774);
nor U5710 (N_5710,N_3601,N_3383);
and U5711 (N_5711,N_2814,N_2965);
xnor U5712 (N_5712,N_3290,N_3726);
and U5713 (N_5713,N_3200,N_3839);
nand U5714 (N_5714,N_3032,N_3519);
and U5715 (N_5715,N_2968,N_3636);
and U5716 (N_5716,N_3297,N_2150);
and U5717 (N_5717,N_3041,N_2504);
nand U5718 (N_5718,N_3048,N_3398);
or U5719 (N_5719,N_3608,N_3948);
xor U5720 (N_5720,N_3051,N_3300);
nand U5721 (N_5721,N_3579,N_3648);
or U5722 (N_5722,N_2036,N_2222);
or U5723 (N_5723,N_3019,N_2277);
xnor U5724 (N_5724,N_3833,N_3861);
nor U5725 (N_5725,N_3771,N_3014);
or U5726 (N_5726,N_2219,N_2100);
and U5727 (N_5727,N_3165,N_3859);
nor U5728 (N_5728,N_3332,N_2986);
or U5729 (N_5729,N_2203,N_3707);
xor U5730 (N_5730,N_3033,N_3374);
and U5731 (N_5731,N_3558,N_3244);
or U5732 (N_5732,N_3041,N_2158);
nand U5733 (N_5733,N_2061,N_2502);
xnor U5734 (N_5734,N_2955,N_2900);
nand U5735 (N_5735,N_2064,N_2879);
nand U5736 (N_5736,N_2481,N_3240);
or U5737 (N_5737,N_2357,N_3138);
xnor U5738 (N_5738,N_3638,N_2297);
or U5739 (N_5739,N_3114,N_3695);
nand U5740 (N_5740,N_2149,N_3905);
xnor U5741 (N_5741,N_3830,N_2458);
and U5742 (N_5742,N_2762,N_2576);
xor U5743 (N_5743,N_3569,N_2264);
nand U5744 (N_5744,N_2629,N_3214);
nor U5745 (N_5745,N_3575,N_3574);
xor U5746 (N_5746,N_2087,N_3192);
and U5747 (N_5747,N_3129,N_2343);
nand U5748 (N_5748,N_2826,N_3530);
nand U5749 (N_5749,N_3853,N_3026);
xnor U5750 (N_5750,N_3918,N_2909);
xnor U5751 (N_5751,N_2830,N_2817);
and U5752 (N_5752,N_3107,N_3443);
xor U5753 (N_5753,N_3385,N_2790);
or U5754 (N_5754,N_2068,N_3085);
nor U5755 (N_5755,N_3374,N_2786);
and U5756 (N_5756,N_2218,N_2594);
or U5757 (N_5757,N_2979,N_2468);
nand U5758 (N_5758,N_2358,N_3540);
or U5759 (N_5759,N_3126,N_3297);
and U5760 (N_5760,N_3406,N_3877);
and U5761 (N_5761,N_2183,N_2135);
or U5762 (N_5762,N_2567,N_2876);
nor U5763 (N_5763,N_3257,N_2459);
nand U5764 (N_5764,N_3994,N_2578);
or U5765 (N_5765,N_3303,N_3689);
and U5766 (N_5766,N_3904,N_2688);
nor U5767 (N_5767,N_2843,N_2134);
and U5768 (N_5768,N_3455,N_2281);
and U5769 (N_5769,N_2775,N_3059);
xnor U5770 (N_5770,N_2836,N_2416);
nand U5771 (N_5771,N_2559,N_2310);
or U5772 (N_5772,N_3247,N_3979);
xor U5773 (N_5773,N_3487,N_2071);
and U5774 (N_5774,N_3342,N_2845);
xor U5775 (N_5775,N_2631,N_2103);
or U5776 (N_5776,N_2867,N_3383);
nor U5777 (N_5777,N_2728,N_3720);
nor U5778 (N_5778,N_3000,N_3587);
xor U5779 (N_5779,N_3715,N_2452);
xnor U5780 (N_5780,N_3889,N_2692);
or U5781 (N_5781,N_2282,N_3353);
nand U5782 (N_5782,N_2719,N_2399);
xnor U5783 (N_5783,N_3210,N_2777);
and U5784 (N_5784,N_3233,N_3659);
xnor U5785 (N_5785,N_2985,N_2843);
nand U5786 (N_5786,N_2988,N_3673);
or U5787 (N_5787,N_3921,N_3370);
nand U5788 (N_5788,N_3473,N_3710);
or U5789 (N_5789,N_2623,N_2304);
nor U5790 (N_5790,N_3795,N_2337);
and U5791 (N_5791,N_3030,N_3888);
and U5792 (N_5792,N_2082,N_3362);
or U5793 (N_5793,N_2608,N_3770);
or U5794 (N_5794,N_3644,N_3795);
and U5795 (N_5795,N_3657,N_3892);
or U5796 (N_5796,N_3321,N_3732);
nand U5797 (N_5797,N_3550,N_2470);
and U5798 (N_5798,N_2903,N_3411);
nor U5799 (N_5799,N_2857,N_2337);
or U5800 (N_5800,N_2993,N_2486);
nand U5801 (N_5801,N_2474,N_2457);
xnor U5802 (N_5802,N_2119,N_2420);
nor U5803 (N_5803,N_3883,N_3446);
or U5804 (N_5804,N_3618,N_3840);
or U5805 (N_5805,N_2905,N_2461);
and U5806 (N_5806,N_2527,N_2438);
and U5807 (N_5807,N_2887,N_2720);
and U5808 (N_5808,N_3572,N_3737);
nand U5809 (N_5809,N_3193,N_3007);
xnor U5810 (N_5810,N_2532,N_3259);
or U5811 (N_5811,N_3974,N_3716);
xor U5812 (N_5812,N_2900,N_3696);
xor U5813 (N_5813,N_2740,N_3298);
nand U5814 (N_5814,N_3542,N_2050);
and U5815 (N_5815,N_3816,N_2659);
nor U5816 (N_5816,N_3823,N_2736);
nand U5817 (N_5817,N_2472,N_2029);
and U5818 (N_5818,N_3325,N_2583);
xor U5819 (N_5819,N_2673,N_3729);
or U5820 (N_5820,N_2289,N_2142);
and U5821 (N_5821,N_3137,N_2319);
and U5822 (N_5822,N_2958,N_2520);
and U5823 (N_5823,N_2154,N_3184);
nand U5824 (N_5824,N_2475,N_3252);
xor U5825 (N_5825,N_2041,N_2300);
nor U5826 (N_5826,N_2953,N_2617);
xnor U5827 (N_5827,N_2810,N_2034);
nand U5828 (N_5828,N_2253,N_3528);
nand U5829 (N_5829,N_2520,N_3108);
or U5830 (N_5830,N_2474,N_3300);
xnor U5831 (N_5831,N_2586,N_2023);
nand U5832 (N_5832,N_2928,N_2606);
or U5833 (N_5833,N_2015,N_2651);
nor U5834 (N_5834,N_2495,N_2608);
and U5835 (N_5835,N_2480,N_3143);
xnor U5836 (N_5836,N_3773,N_2831);
and U5837 (N_5837,N_2803,N_3527);
nand U5838 (N_5838,N_3702,N_2799);
nand U5839 (N_5839,N_3838,N_3277);
nand U5840 (N_5840,N_3742,N_3476);
xor U5841 (N_5841,N_2724,N_2470);
and U5842 (N_5842,N_3576,N_3044);
xor U5843 (N_5843,N_3692,N_2134);
xor U5844 (N_5844,N_2996,N_3519);
or U5845 (N_5845,N_3456,N_3319);
nor U5846 (N_5846,N_3723,N_3184);
nor U5847 (N_5847,N_3268,N_2941);
and U5848 (N_5848,N_2950,N_2784);
nor U5849 (N_5849,N_3949,N_3244);
and U5850 (N_5850,N_2031,N_3678);
xnor U5851 (N_5851,N_2377,N_2429);
nand U5852 (N_5852,N_2529,N_2319);
and U5853 (N_5853,N_2182,N_2557);
or U5854 (N_5854,N_2484,N_3238);
or U5855 (N_5855,N_2522,N_2730);
or U5856 (N_5856,N_3344,N_3693);
nand U5857 (N_5857,N_2913,N_3948);
xnor U5858 (N_5858,N_2377,N_2740);
nand U5859 (N_5859,N_3612,N_3863);
or U5860 (N_5860,N_2584,N_3326);
and U5861 (N_5861,N_3403,N_3383);
xor U5862 (N_5862,N_2651,N_2667);
and U5863 (N_5863,N_3488,N_3769);
nor U5864 (N_5864,N_2721,N_3737);
and U5865 (N_5865,N_3368,N_3605);
nor U5866 (N_5866,N_2354,N_3474);
and U5867 (N_5867,N_3997,N_2990);
nor U5868 (N_5868,N_3993,N_2898);
xor U5869 (N_5869,N_3015,N_3182);
nand U5870 (N_5870,N_3733,N_3765);
or U5871 (N_5871,N_2402,N_3738);
xnor U5872 (N_5872,N_2214,N_2720);
or U5873 (N_5873,N_2074,N_3407);
nand U5874 (N_5874,N_3106,N_2982);
nor U5875 (N_5875,N_3664,N_3069);
xnor U5876 (N_5876,N_3908,N_3989);
nand U5877 (N_5877,N_3105,N_3076);
nand U5878 (N_5878,N_2141,N_2652);
nor U5879 (N_5879,N_3541,N_2681);
nand U5880 (N_5880,N_2383,N_3392);
xor U5881 (N_5881,N_2584,N_3763);
nor U5882 (N_5882,N_3381,N_2084);
or U5883 (N_5883,N_3089,N_3442);
and U5884 (N_5884,N_3013,N_3262);
or U5885 (N_5885,N_2428,N_3401);
and U5886 (N_5886,N_3194,N_3000);
nand U5887 (N_5887,N_2095,N_2891);
and U5888 (N_5888,N_3641,N_3189);
nor U5889 (N_5889,N_3806,N_3911);
xnor U5890 (N_5890,N_3223,N_3715);
or U5891 (N_5891,N_2764,N_2075);
or U5892 (N_5892,N_3872,N_3658);
nor U5893 (N_5893,N_3480,N_3367);
or U5894 (N_5894,N_3720,N_2054);
or U5895 (N_5895,N_3844,N_2300);
xnor U5896 (N_5896,N_3505,N_2158);
nand U5897 (N_5897,N_2731,N_2487);
nand U5898 (N_5898,N_2696,N_2210);
nand U5899 (N_5899,N_2166,N_3267);
or U5900 (N_5900,N_2066,N_3957);
and U5901 (N_5901,N_2330,N_3680);
xnor U5902 (N_5902,N_3036,N_2978);
xnor U5903 (N_5903,N_3798,N_2408);
nand U5904 (N_5904,N_2920,N_2444);
xor U5905 (N_5905,N_3099,N_3321);
nor U5906 (N_5906,N_3935,N_2753);
nor U5907 (N_5907,N_3719,N_2972);
nand U5908 (N_5908,N_3058,N_3646);
or U5909 (N_5909,N_2303,N_2274);
xnor U5910 (N_5910,N_2354,N_2067);
nor U5911 (N_5911,N_2315,N_3767);
or U5912 (N_5912,N_3608,N_3730);
and U5913 (N_5913,N_2213,N_2952);
xor U5914 (N_5914,N_3066,N_2328);
or U5915 (N_5915,N_3070,N_3525);
xnor U5916 (N_5916,N_2618,N_3852);
and U5917 (N_5917,N_3623,N_2393);
xnor U5918 (N_5918,N_3945,N_3964);
nor U5919 (N_5919,N_3864,N_2198);
nor U5920 (N_5920,N_3355,N_3704);
nor U5921 (N_5921,N_3532,N_2734);
and U5922 (N_5922,N_3130,N_3898);
xor U5923 (N_5923,N_3558,N_2113);
nor U5924 (N_5924,N_3030,N_2143);
nand U5925 (N_5925,N_3563,N_3336);
nand U5926 (N_5926,N_3811,N_3397);
nand U5927 (N_5927,N_2137,N_3228);
xnor U5928 (N_5928,N_2296,N_2472);
xor U5929 (N_5929,N_2856,N_2504);
nand U5930 (N_5930,N_3642,N_3186);
nor U5931 (N_5931,N_2458,N_2355);
xnor U5932 (N_5932,N_2718,N_2224);
nand U5933 (N_5933,N_3128,N_3056);
xnor U5934 (N_5934,N_2573,N_2095);
nor U5935 (N_5935,N_2054,N_3003);
xnor U5936 (N_5936,N_2639,N_3615);
nor U5937 (N_5937,N_3489,N_3762);
or U5938 (N_5938,N_2932,N_2038);
and U5939 (N_5939,N_2432,N_2610);
nand U5940 (N_5940,N_2479,N_2340);
xnor U5941 (N_5941,N_3642,N_3577);
or U5942 (N_5942,N_3760,N_3134);
nand U5943 (N_5943,N_2698,N_3627);
and U5944 (N_5944,N_3716,N_2782);
nor U5945 (N_5945,N_2307,N_3454);
and U5946 (N_5946,N_3652,N_2128);
or U5947 (N_5947,N_2640,N_2938);
xor U5948 (N_5948,N_2163,N_2577);
or U5949 (N_5949,N_2268,N_2746);
xor U5950 (N_5950,N_2696,N_3867);
and U5951 (N_5951,N_3152,N_3796);
and U5952 (N_5952,N_3036,N_3230);
and U5953 (N_5953,N_2344,N_3352);
nand U5954 (N_5954,N_3991,N_2411);
or U5955 (N_5955,N_2814,N_2703);
and U5956 (N_5956,N_2253,N_3252);
xnor U5957 (N_5957,N_2391,N_3185);
and U5958 (N_5958,N_2479,N_2232);
nand U5959 (N_5959,N_2590,N_2980);
or U5960 (N_5960,N_3154,N_2862);
xor U5961 (N_5961,N_2470,N_2183);
nand U5962 (N_5962,N_3791,N_3154);
xor U5963 (N_5963,N_3688,N_3062);
nor U5964 (N_5964,N_2029,N_3119);
nand U5965 (N_5965,N_2438,N_3673);
or U5966 (N_5966,N_2966,N_2362);
nand U5967 (N_5967,N_3454,N_2310);
or U5968 (N_5968,N_3890,N_3288);
nand U5969 (N_5969,N_2456,N_3554);
and U5970 (N_5970,N_2481,N_2778);
and U5971 (N_5971,N_3920,N_2913);
nor U5972 (N_5972,N_3585,N_3659);
xnor U5973 (N_5973,N_2968,N_2350);
and U5974 (N_5974,N_2531,N_2551);
xor U5975 (N_5975,N_2655,N_3211);
xnor U5976 (N_5976,N_2525,N_3865);
xor U5977 (N_5977,N_2011,N_2602);
xnor U5978 (N_5978,N_3844,N_3431);
nand U5979 (N_5979,N_2662,N_3770);
and U5980 (N_5980,N_3141,N_3251);
nand U5981 (N_5981,N_2359,N_3513);
nor U5982 (N_5982,N_2652,N_3991);
nor U5983 (N_5983,N_3914,N_3855);
nand U5984 (N_5984,N_3404,N_2150);
or U5985 (N_5985,N_3396,N_2400);
xor U5986 (N_5986,N_2896,N_3187);
nor U5987 (N_5987,N_3753,N_3386);
or U5988 (N_5988,N_3597,N_3460);
or U5989 (N_5989,N_3687,N_2493);
xor U5990 (N_5990,N_3047,N_3161);
nor U5991 (N_5991,N_2850,N_2079);
xnor U5992 (N_5992,N_3561,N_2177);
or U5993 (N_5993,N_3571,N_3678);
nor U5994 (N_5994,N_3684,N_2660);
xnor U5995 (N_5995,N_2482,N_3549);
or U5996 (N_5996,N_2054,N_2570);
or U5997 (N_5997,N_2692,N_3923);
and U5998 (N_5998,N_3956,N_2726);
and U5999 (N_5999,N_2569,N_2948);
and U6000 (N_6000,N_4103,N_4354);
and U6001 (N_6001,N_4301,N_5135);
nand U6002 (N_6002,N_5014,N_4950);
or U6003 (N_6003,N_4138,N_5813);
xnor U6004 (N_6004,N_4848,N_5031);
and U6005 (N_6005,N_4704,N_4619);
nand U6006 (N_6006,N_4483,N_5217);
nor U6007 (N_6007,N_5733,N_5743);
xnor U6008 (N_6008,N_4226,N_4441);
and U6009 (N_6009,N_4062,N_4465);
or U6010 (N_6010,N_4426,N_5313);
and U6011 (N_6011,N_5554,N_5245);
nand U6012 (N_6012,N_4931,N_5249);
and U6013 (N_6013,N_4575,N_4146);
xor U6014 (N_6014,N_5248,N_4785);
nand U6015 (N_6015,N_4231,N_5696);
and U6016 (N_6016,N_5271,N_4476);
or U6017 (N_6017,N_4596,N_4529);
nor U6018 (N_6018,N_4321,N_5358);
nand U6019 (N_6019,N_5586,N_5240);
or U6020 (N_6020,N_5516,N_4431);
xnor U6021 (N_6021,N_4816,N_5747);
nor U6022 (N_6022,N_4825,N_4257);
nand U6023 (N_6023,N_4292,N_4063);
nand U6024 (N_6024,N_4627,N_5418);
xor U6025 (N_6025,N_4054,N_4938);
xor U6026 (N_6026,N_5151,N_4453);
nand U6027 (N_6027,N_4568,N_5609);
nand U6028 (N_6028,N_5835,N_4173);
nand U6029 (N_6029,N_5417,N_4872);
or U6030 (N_6030,N_5209,N_4290);
xnor U6031 (N_6031,N_5081,N_4068);
nor U6032 (N_6032,N_4571,N_5889);
nand U6033 (N_6033,N_5004,N_4428);
nor U6034 (N_6034,N_4709,N_4207);
or U6035 (N_6035,N_5080,N_5264);
xnor U6036 (N_6036,N_4444,N_4884);
nand U6037 (N_6037,N_4224,N_5930);
nand U6038 (N_6038,N_5875,N_5924);
nor U6039 (N_6039,N_4688,N_5472);
and U6040 (N_6040,N_5578,N_5452);
nand U6041 (N_6041,N_5369,N_5092);
xor U6042 (N_6042,N_4873,N_5295);
and U6043 (N_6043,N_4693,N_4936);
nor U6044 (N_6044,N_4202,N_4663);
or U6045 (N_6045,N_5167,N_5337);
nand U6046 (N_6046,N_5778,N_5037);
nand U6047 (N_6047,N_4576,N_4748);
or U6048 (N_6048,N_5508,N_5323);
or U6049 (N_6049,N_4573,N_4554);
nor U6050 (N_6050,N_5289,N_5117);
nand U6051 (N_6051,N_4674,N_4332);
or U6052 (N_6052,N_5048,N_5247);
nor U6053 (N_6053,N_4863,N_4020);
xor U6054 (N_6054,N_5684,N_5128);
and U6055 (N_6055,N_5792,N_4253);
and U6056 (N_6056,N_5726,N_5635);
and U6057 (N_6057,N_4752,N_4451);
and U6058 (N_6058,N_4157,N_5690);
xnor U6059 (N_6059,N_4864,N_4588);
or U6060 (N_6060,N_5562,N_5277);
nor U6061 (N_6061,N_5978,N_5728);
or U6062 (N_6062,N_4996,N_4605);
nand U6063 (N_6063,N_5294,N_5102);
and U6064 (N_6064,N_4920,N_5234);
and U6065 (N_6065,N_5995,N_5707);
xnor U6066 (N_6066,N_5285,N_4548);
or U6067 (N_6067,N_5156,N_5502);
and U6068 (N_6068,N_5238,N_4985);
or U6069 (N_6069,N_5618,N_4843);
or U6070 (N_6070,N_5364,N_5598);
or U6071 (N_6071,N_5398,N_5841);
and U6072 (N_6072,N_5492,N_4788);
and U6073 (N_6073,N_5612,N_4701);
and U6074 (N_6074,N_5071,N_4763);
xor U6075 (N_6075,N_4512,N_4502);
nand U6076 (N_6076,N_4448,N_5212);
xnor U6077 (N_6077,N_5720,N_5711);
nand U6078 (N_6078,N_5695,N_5381);
xnor U6079 (N_6079,N_4600,N_4417);
nor U6080 (N_6080,N_5730,N_4654);
nor U6081 (N_6081,N_4632,N_4021);
and U6082 (N_6082,N_5632,N_5988);
and U6083 (N_6083,N_4880,N_5438);
or U6084 (N_6084,N_5574,N_5393);
or U6085 (N_6085,N_4239,N_5959);
xnor U6086 (N_6086,N_4587,N_4683);
and U6087 (N_6087,N_5994,N_4361);
or U6088 (N_6088,N_4655,N_4852);
nor U6089 (N_6089,N_4245,N_5310);
xor U6090 (N_6090,N_4589,N_5833);
nand U6091 (N_6091,N_5363,N_4120);
nor U6092 (N_6092,N_4800,N_5172);
nor U6093 (N_6093,N_4133,N_5488);
nor U6094 (N_6094,N_5410,N_4932);
xor U6095 (N_6095,N_4064,N_5231);
or U6096 (N_6096,N_5246,N_5675);
and U6097 (N_6097,N_4498,N_4810);
xnor U6098 (N_6098,N_4877,N_4993);
xor U6099 (N_6099,N_4408,N_5282);
nand U6100 (N_6100,N_4601,N_5573);
nand U6101 (N_6101,N_5493,N_5126);
or U6102 (N_6102,N_4539,N_4425);
nand U6103 (N_6103,N_5713,N_4486);
xnor U6104 (N_6104,N_4187,N_5577);
nor U6105 (N_6105,N_5397,N_4044);
nor U6106 (N_6106,N_4255,N_5170);
and U6107 (N_6107,N_5811,N_4939);
nand U6108 (N_6108,N_4339,N_5750);
or U6109 (N_6109,N_4598,N_4343);
xnor U6110 (N_6110,N_4637,N_4527);
and U6111 (N_6111,N_4492,N_5845);
nor U6112 (N_6112,N_5773,N_4190);
or U6113 (N_6113,N_4506,N_5769);
xor U6114 (N_6114,N_4188,N_4553);
xnor U6115 (N_6115,N_4610,N_5718);
and U6116 (N_6116,N_5885,N_4040);
or U6117 (N_6117,N_5288,N_4925);
xor U6118 (N_6118,N_5342,N_4928);
or U6119 (N_6119,N_4052,N_5592);
nand U6120 (N_6120,N_4849,N_4764);
or U6121 (N_6121,N_4724,N_4489);
nand U6122 (N_6122,N_5570,N_5389);
and U6123 (N_6123,N_4208,N_4930);
nand U6124 (N_6124,N_5098,N_4842);
xnor U6125 (N_6125,N_5022,N_5878);
nand U6126 (N_6126,N_4046,N_4907);
or U6127 (N_6127,N_5680,N_5453);
xnor U6128 (N_6128,N_5340,N_5274);
or U6129 (N_6129,N_5341,N_5872);
or U6130 (N_6130,N_4404,N_4283);
xor U6131 (N_6131,N_4243,N_5049);
or U6132 (N_6132,N_5040,N_5893);
nor U6133 (N_6133,N_5668,N_5515);
xor U6134 (N_6134,N_5704,N_4914);
nand U6135 (N_6135,N_5162,N_5205);
and U6136 (N_6136,N_5464,N_4656);
or U6137 (N_6137,N_4707,N_5806);
and U6138 (N_6138,N_5854,N_4369);
nand U6139 (N_6139,N_4978,N_4983);
nor U6140 (N_6140,N_5332,N_5350);
or U6141 (N_6141,N_4429,N_4703);
nand U6142 (N_6142,N_4944,N_4813);
or U6143 (N_6143,N_4533,N_5531);
nor U6144 (N_6144,N_4186,N_5512);
nor U6145 (N_6145,N_5146,N_5280);
nor U6146 (N_6146,N_4114,N_5585);
nor U6147 (N_6147,N_4557,N_4591);
nand U6148 (N_6148,N_5401,N_4935);
nand U6149 (N_6149,N_5386,N_5977);
nor U6150 (N_6150,N_5185,N_4771);
nor U6151 (N_6151,N_5859,N_4413);
nand U6152 (N_6152,N_5178,N_5634);
and U6153 (N_6153,N_4664,N_5682);
nand U6154 (N_6154,N_5252,N_4593);
or U6155 (N_6155,N_4463,N_4370);
and U6156 (N_6156,N_5458,N_4574);
nor U6157 (N_6157,N_5907,N_5745);
nand U6158 (N_6158,N_4711,N_5347);
nor U6159 (N_6159,N_4334,N_5106);
or U6160 (N_6160,N_4201,N_4182);
or U6161 (N_6161,N_4549,N_5915);
nand U6162 (N_6162,N_5874,N_5537);
xnor U6163 (N_6163,N_4324,N_5015);
or U6164 (N_6164,N_5858,N_5793);
xor U6165 (N_6165,N_4858,N_5463);
or U6166 (N_6166,N_4160,N_5032);
and U6167 (N_6167,N_5055,N_5072);
or U6168 (N_6168,N_4639,N_5933);
nor U6169 (N_6169,N_5853,N_5108);
xnor U6170 (N_6170,N_5630,N_5519);
nand U6171 (N_6171,N_4302,N_4437);
nor U6172 (N_6172,N_5287,N_4738);
or U6173 (N_6173,N_4464,N_4795);
nand U6174 (N_6174,N_5557,N_4172);
or U6175 (N_6175,N_5912,N_4875);
xnor U6176 (N_6176,N_4633,N_5949);
xnor U6177 (N_6177,N_5073,N_5758);
nand U6178 (N_6178,N_5569,N_4244);
nor U6179 (N_6179,N_5767,N_5074);
nand U6180 (N_6180,N_4113,N_4143);
xor U6181 (N_6181,N_5955,N_4047);
or U6182 (N_6182,N_4288,N_4027);
or U6183 (N_6183,N_5385,N_5936);
xnor U6184 (N_6184,N_5931,N_5154);
nand U6185 (N_6185,N_4341,N_5681);
or U6186 (N_6186,N_4101,N_4176);
nand U6187 (N_6187,N_5088,N_4168);
nor U6188 (N_6188,N_5132,N_5714);
or U6189 (N_6189,N_4325,N_5239);
xor U6190 (N_6190,N_4058,N_4434);
and U6191 (N_6191,N_4670,N_5651);
nand U6192 (N_6192,N_5993,N_5474);
nand U6193 (N_6193,N_4127,N_5535);
or U6194 (N_6194,N_5625,N_5960);
nand U6195 (N_6195,N_5378,N_5286);
nand U6196 (N_6196,N_4070,N_5201);
nor U6197 (N_6197,N_4956,N_4974);
nand U6198 (N_6198,N_4005,N_4728);
or U6199 (N_6199,N_4712,N_5867);
xnor U6200 (N_6200,N_4085,N_5517);
xor U6201 (N_6201,N_5065,N_5593);
nor U6202 (N_6202,N_5655,N_4254);
nand U6203 (N_6203,N_4261,N_5383);
and U6204 (N_6204,N_4487,N_4997);
nand U6205 (N_6205,N_4668,N_5000);
nor U6206 (N_6206,N_4505,N_4350);
or U6207 (N_6207,N_4640,N_5921);
nand U6208 (N_6208,N_4107,N_5021);
nor U6209 (N_6209,N_5789,N_5673);
or U6210 (N_6210,N_5171,N_4802);
and U6211 (N_6211,N_5270,N_5660);
nor U6212 (N_6212,N_4147,N_4870);
and U6213 (N_6213,N_5199,N_4280);
nor U6214 (N_6214,N_4616,N_5965);
nor U6215 (N_6215,N_4841,N_5173);
and U6216 (N_6216,N_5650,N_4910);
nand U6217 (N_6217,N_5862,N_4720);
nor U6218 (N_6218,N_5616,N_4937);
and U6219 (N_6219,N_4384,N_4756);
nor U6220 (N_6220,N_5153,N_4310);
nor U6221 (N_6221,N_5339,N_4178);
and U6222 (N_6222,N_5432,N_4647);
xor U6223 (N_6223,N_4999,N_5365);
xor U6224 (N_6224,N_5975,N_4091);
nand U6225 (N_6225,N_4584,N_5045);
and U6226 (N_6226,N_4789,N_4879);
nor U6227 (N_6227,N_4761,N_4791);
and U6228 (N_6228,N_5572,N_4272);
nor U6229 (N_6229,N_5211,N_5888);
and U6230 (N_6230,N_5552,N_4374);
or U6231 (N_6231,N_5964,N_4990);
nand U6232 (N_6232,N_5250,N_5206);
or U6233 (N_6233,N_4913,N_5388);
nor U6234 (N_6234,N_4909,N_4328);
xnor U6235 (N_6235,N_4976,N_5953);
or U6236 (N_6236,N_4890,N_4561);
and U6237 (N_6237,N_5213,N_4866);
xnor U6238 (N_6238,N_4395,N_5105);
xor U6239 (N_6239,N_4900,N_4626);
nand U6240 (N_6240,N_5068,N_5429);
nand U6241 (N_6241,N_4965,N_5085);
nor U6242 (N_6242,N_4675,N_4973);
xnor U6243 (N_6243,N_5445,N_5605);
nor U6244 (N_6244,N_5896,N_4439);
or U6245 (N_6245,N_5198,N_4811);
and U6246 (N_6246,N_4089,N_5320);
and U6247 (N_6247,N_4525,N_4820);
nand U6248 (N_6248,N_4216,N_5780);
nor U6249 (N_6249,N_5740,N_5158);
and U6250 (N_6250,N_4170,N_4916);
and U6251 (N_6251,N_5372,N_4195);
nand U6252 (N_6252,N_5717,N_5749);
nor U6253 (N_6253,N_4689,N_5497);
or U6254 (N_6254,N_5599,N_4203);
xor U6255 (N_6255,N_5678,N_4926);
nor U6256 (N_6256,N_4003,N_5805);
nand U6257 (N_6257,N_5615,N_4097);
nor U6258 (N_6258,N_5812,N_4697);
xor U6259 (N_6259,N_5791,N_5543);
or U6260 (N_6260,N_4482,N_4346);
xnor U6261 (N_6261,N_4686,N_4340);
nand U6262 (N_6262,N_4962,N_4002);
xor U6263 (N_6263,N_4776,N_4475);
or U6264 (N_6264,N_4679,N_4555);
and U6265 (N_6265,N_4037,N_4406);
xnor U6266 (N_6266,N_5118,N_5958);
and U6267 (N_6267,N_4676,N_4594);
and U6268 (N_6268,N_4887,N_4941);
nor U6269 (N_6269,N_5373,N_4702);
nand U6270 (N_6270,N_4358,N_5189);
nand U6271 (N_6271,N_4353,N_5788);
xor U6272 (N_6272,N_4380,N_5762);
or U6273 (N_6273,N_4660,N_4570);
xor U6274 (N_6274,N_5708,N_5734);
xnor U6275 (N_6275,N_4634,N_5620);
or U6276 (N_6276,N_5215,N_4268);
nor U6277 (N_6277,N_4758,N_4139);
nand U6278 (N_6278,N_4236,N_4387);
and U6279 (N_6279,N_5722,N_4249);
xnor U6280 (N_6280,N_5428,N_4644);
or U6281 (N_6281,N_4893,N_4391);
nand U6282 (N_6282,N_5403,N_5224);
xnor U6283 (N_6283,N_4414,N_4577);
nand U6284 (N_6284,N_5104,N_4322);
or U6285 (N_6285,N_5175,N_4958);
or U6286 (N_6286,N_5402,N_5269);
xnor U6287 (N_6287,N_4899,N_5043);
xor U6288 (N_6288,N_5525,N_4171);
nand U6289 (N_6289,N_5529,N_4443);
and U6290 (N_6290,N_4508,N_5989);
xnor U6291 (N_6291,N_5943,N_4242);
xnor U6292 (N_6292,N_5265,N_5737);
nor U6293 (N_6293,N_5276,N_4356);
and U6294 (N_6294,N_4572,N_5099);
nand U6295 (N_6295,N_4278,N_4184);
xnor U6296 (N_6296,N_4912,N_4213);
or U6297 (N_6297,N_5775,N_5882);
and U6298 (N_6298,N_5894,N_5705);
and U6299 (N_6299,N_5404,N_4327);
xor U6300 (N_6300,N_4081,N_5984);
nor U6301 (N_6301,N_5870,N_4599);
xnor U6302 (N_6302,N_4049,N_5140);
nand U6303 (N_6303,N_4102,N_4264);
xnor U6304 (N_6304,N_5563,N_4499);
xnor U6305 (N_6305,N_4263,N_4342);
and U6306 (N_6306,N_4750,N_5507);
nor U6307 (N_6307,N_5446,N_4410);
nand U6308 (N_6308,N_4876,N_5909);
nand U6309 (N_6309,N_5380,N_5584);
and U6310 (N_6310,N_5305,N_4725);
xor U6311 (N_6311,N_5476,N_4294);
xor U6312 (N_6312,N_5093,N_4917);
nand U6313 (N_6313,N_5054,N_4844);
xnor U6314 (N_6314,N_5603,N_5887);
nor U6315 (N_6315,N_5691,N_5848);
or U6316 (N_6316,N_5091,N_5868);
or U6317 (N_6317,N_5110,N_5763);
xnor U6318 (N_6318,N_4981,N_4645);
nor U6319 (N_6319,N_4377,N_5028);
xnor U6320 (N_6320,N_4716,N_5968);
nand U6321 (N_6321,N_5186,N_4155);
nand U6322 (N_6322,N_4747,N_5024);
or U6323 (N_6323,N_5631,N_5840);
nor U6324 (N_6324,N_5130,N_4969);
or U6325 (N_6325,N_5601,N_4753);
nand U6326 (N_6326,N_4164,N_4765);
nor U6327 (N_6327,N_5371,N_4613);
nand U6328 (N_6328,N_5555,N_5127);
and U6329 (N_6329,N_4017,N_5657);
or U6330 (N_6330,N_5384,N_4421);
xnor U6331 (N_6331,N_4034,N_4351);
xor U6332 (N_6332,N_5374,N_5430);
and U6333 (N_6333,N_5216,N_4951);
or U6334 (N_6334,N_5075,N_5647);
or U6335 (N_6335,N_5544,N_4381);
or U6336 (N_6336,N_4528,N_4450);
nand U6337 (N_6337,N_5884,N_5470);
and U6338 (N_6338,N_5541,N_4167);
and U6339 (N_6339,N_4766,N_5168);
nand U6340 (N_6340,N_5416,N_4478);
and U6341 (N_6341,N_5376,N_4726);
nand U6342 (N_6342,N_4635,N_4218);
nor U6343 (N_6343,N_5712,N_4995);
xor U6344 (N_6344,N_5799,N_4082);
xnor U6345 (N_6345,N_4181,N_4135);
and U6346 (N_6346,N_5278,N_4851);
nor U6347 (N_6347,N_5222,N_5451);
or U6348 (N_6348,N_5083,N_5422);
or U6349 (N_6349,N_4982,N_4156);
and U6350 (N_6350,N_5308,N_4717);
nand U6351 (N_6351,N_5917,N_5348);
nor U6352 (N_6352,N_4485,N_4882);
or U6353 (N_6353,N_5619,N_5210);
nand U6354 (N_6354,N_4388,N_5467);
and U6355 (N_6355,N_5129,N_5606);
xnor U6356 (N_6356,N_5735,N_4927);
nor U6357 (N_6357,N_5116,N_5257);
and U6358 (N_6358,N_4745,N_5957);
nand U6359 (N_6359,N_4488,N_4401);
and U6360 (N_6360,N_5732,N_5768);
xor U6361 (N_6361,N_4611,N_5700);
nand U6362 (N_6362,N_5152,N_5942);
nand U6363 (N_6363,N_5659,N_5662);
or U6364 (N_6364,N_5319,N_4886);
nand U6365 (N_6365,N_4620,N_5672);
nand U6366 (N_6366,N_4241,N_5610);
or U6367 (N_6367,N_4579,N_5941);
xor U6368 (N_6368,N_4162,N_5351);
nand U6369 (N_6369,N_5851,N_5361);
xor U6370 (N_6370,N_5200,N_5897);
and U6371 (N_6371,N_5654,N_4379);
and U6372 (N_6372,N_5078,N_5594);
xnor U6373 (N_6373,N_5621,N_4442);
or U6374 (N_6374,N_4045,N_5640);
nor U6375 (N_6375,N_5765,N_4713);
and U6376 (N_6376,N_5084,N_5456);
nor U6377 (N_6377,N_4298,N_4519);
or U6378 (N_6378,N_4768,N_5639);
nor U6379 (N_6379,N_4977,N_4817);
or U6380 (N_6380,N_5483,N_4824);
xnor U6381 (N_6381,N_5665,N_4558);
xor U6382 (N_6382,N_5298,N_5785);
or U6383 (N_6383,N_4744,N_4372);
nor U6384 (N_6384,N_5094,N_5473);
xor U6385 (N_6385,N_4865,N_4636);
nand U6386 (N_6386,N_4830,N_4023);
and U6387 (N_6387,N_5122,N_4335);
nor U6388 (N_6388,N_4531,N_5827);
and U6389 (N_6389,N_5008,N_4667);
xor U6390 (N_6390,N_5952,N_4892);
xnor U6391 (N_6391,N_5898,N_5880);
nor U6392 (N_6392,N_4087,N_4193);
nand U6393 (N_6393,N_5992,N_5809);
nand U6394 (N_6394,N_5499,N_4603);
nor U6395 (N_6395,N_5336,N_5546);
xor U6396 (N_6396,N_4311,N_4940);
or U6397 (N_6397,N_4347,N_4737);
or U6398 (N_6398,N_5437,N_4095);
or U6399 (N_6399,N_4397,N_4299);
or U6400 (N_6400,N_4467,N_5677);
nor U6401 (N_6401,N_5149,N_5772);
nand U6402 (N_6402,N_4859,N_4457);
nor U6403 (N_6403,N_4905,N_5795);
and U6404 (N_6404,N_5596,N_5967);
xor U6405 (N_6405,N_5804,N_4007);
xnor U6406 (N_6406,N_4125,N_4234);
nor U6407 (N_6407,N_5455,N_4303);
and U6408 (N_6408,N_5136,N_5831);
or U6409 (N_6409,N_4191,N_5946);
xnor U6410 (N_6410,N_4966,N_5913);
nor U6411 (N_6411,N_5645,N_5739);
or U6412 (N_6412,N_5561,N_4869);
or U6413 (N_6413,N_4612,N_5935);
nand U6414 (N_6414,N_5814,N_4142);
or U6415 (N_6415,N_5038,N_4206);
nor U6416 (N_6416,N_4032,N_5727);
and U6417 (N_6417,N_5808,N_5395);
xnor U6418 (N_6418,N_4780,N_5399);
nor U6419 (N_6419,N_5834,N_5932);
or U6420 (N_6420,N_4894,N_5617);
nand U6421 (N_6421,N_4200,N_4080);
nor U6422 (N_6422,N_4772,N_4790);
and U6423 (N_6423,N_5522,N_4832);
xor U6424 (N_6424,N_4411,N_4069);
xor U6425 (N_6425,N_4694,N_4386);
xnor U6426 (N_6426,N_4608,N_5316);
nor U6427 (N_6427,N_5487,N_4862);
or U6428 (N_6428,N_4727,N_5566);
or U6429 (N_6429,N_4530,N_5643);
xor U6430 (N_6430,N_5477,N_5017);
and U6431 (N_6431,N_4651,N_4390);
nor U6432 (N_6432,N_4375,N_4210);
and U6433 (N_6433,N_4371,N_5018);
and U6434 (N_6434,N_4602,N_4757);
and U6435 (N_6435,N_5580,N_5521);
nand U6436 (N_6436,N_5821,N_5147);
nand U6437 (N_6437,N_4071,N_5160);
or U6438 (N_6438,N_4315,N_4933);
or U6439 (N_6439,N_5462,N_4345);
and U6440 (N_6440,N_4104,N_5802);
nand U6441 (N_6441,N_4992,N_4128);
nand U6442 (N_6442,N_5721,N_5836);
and U6443 (N_6443,N_5818,N_4535);
nor U6444 (N_6444,N_5759,N_5484);
or U6445 (N_6445,N_4698,N_5044);
xnor U6446 (N_6446,N_4883,N_4084);
xor U6447 (N_6447,N_4316,N_4118);
or U6448 (N_6448,N_5237,N_5387);
nor U6449 (N_6449,N_5095,N_4874);
or U6450 (N_6450,N_5220,N_5176);
nor U6451 (N_6451,N_5050,N_5797);
or U6452 (N_6452,N_4653,N_4050);
xor U6453 (N_6453,N_4398,N_4440);
or U6454 (N_6454,N_5442,N_4806);
xor U6455 (N_6455,N_4673,N_5689);
or U6456 (N_6456,N_4742,N_4036);
nor U6457 (N_6457,N_4722,N_5019);
or U6458 (N_6458,N_4355,N_4497);
xnor U6459 (N_6459,N_5545,N_5981);
and U6460 (N_6460,N_5548,N_4378);
nor U6461 (N_6461,N_5783,N_5670);
nand U6462 (N_6462,N_4396,N_5971);
and U6463 (N_6463,N_4053,N_5489);
xor U6464 (N_6464,N_4915,N_4400);
nand U6465 (N_6465,N_5279,N_5301);
nor U6466 (N_6466,N_4556,N_5419);
or U6467 (N_6467,N_5194,N_4043);
nand U6468 (N_6468,N_4854,N_5180);
or U6469 (N_6469,N_4552,N_5891);
xnor U6470 (N_6470,N_5608,N_5653);
and U6471 (N_6471,N_4964,N_4165);
nor U6472 (N_6472,N_5998,N_4714);
nor U6473 (N_6473,N_5622,N_5724);
and U6474 (N_6474,N_4331,N_5796);
nand U6475 (N_6475,N_5039,N_5774);
and U6476 (N_6476,N_5330,N_4215);
or U6477 (N_6477,N_4534,N_4592);
and U6478 (N_6478,N_5159,N_4551);
and U6479 (N_6479,N_4407,N_5318);
or U6480 (N_6480,N_5284,N_5261);
or U6481 (N_6481,N_5823,N_4296);
and U6482 (N_6482,N_5303,N_4337);
nor U6483 (N_6483,N_5852,N_4831);
nand U6484 (N_6484,N_5839,N_5699);
and U6485 (N_6485,N_5435,N_4086);
nand U6486 (N_6486,N_4898,N_5627);
xnor U6487 (N_6487,N_4061,N_4814);
nand U6488 (N_6488,N_4083,N_5536);
or U6489 (N_6489,N_5856,N_5235);
nor U6490 (N_6490,N_4661,N_5847);
or U6491 (N_6491,N_5877,N_4222);
and U6492 (N_6492,N_5746,N_4265);
nor U6493 (N_6493,N_5766,N_4902);
or U6494 (N_6494,N_4491,N_4798);
and U6495 (N_6495,N_4389,N_5436);
or U6496 (N_6496,N_4057,N_5272);
and U6497 (N_6497,N_4129,N_4088);
nand U6498 (N_6498,N_4718,N_4246);
xor U6499 (N_6499,N_4520,N_4818);
nor U6500 (N_6500,N_5113,N_4819);
xor U6501 (N_6501,N_4537,N_4897);
and U6502 (N_6502,N_5002,N_5177);
nand U6503 (N_6503,N_5534,N_4060);
nand U6504 (N_6504,N_5475,N_4077);
xnor U6505 (N_6505,N_5131,N_4274);
or U6506 (N_6506,N_5688,N_5029);
nand U6507 (N_6507,N_4319,N_4889);
xor U6508 (N_6508,N_4908,N_5549);
xor U6509 (N_6509,N_5709,N_4685);
or U6510 (N_6510,N_5142,N_4782);
or U6511 (N_6511,N_5307,N_4793);
and U6512 (N_6512,N_4710,N_4116);
nor U6513 (N_6513,N_5524,N_4666);
or U6514 (N_6514,N_4896,N_5409);
nor U6515 (N_6515,N_4364,N_5425);
nor U6516 (N_6516,N_4625,N_4154);
and U6517 (N_6517,N_4775,N_4019);
nand U6518 (N_6518,N_5925,N_4987);
and U6519 (N_6519,N_5648,N_4452);
xor U6520 (N_6520,N_4011,N_4008);
or U6521 (N_6521,N_4059,N_4629);
nor U6522 (N_6522,N_4500,N_4117);
and U6523 (N_6523,N_5326,N_5001);
xor U6524 (N_6524,N_4001,N_5057);
or U6525 (N_6525,N_4252,N_5676);
and U6526 (N_6526,N_5034,N_5214);
xnor U6527 (N_6527,N_4305,N_4262);
or U6528 (N_6528,N_4991,N_5207);
nand U6529 (N_6529,N_5010,N_4778);
or U6530 (N_6530,N_4422,N_5020);
or U6531 (N_6531,N_5685,N_5633);
or U6532 (N_6532,N_5985,N_4433);
nand U6533 (N_6533,N_5667,N_4111);
nand U6534 (N_6534,N_4198,N_4079);
or U6535 (N_6535,N_4881,N_5077);
nand U6536 (N_6536,N_4947,N_4163);
nor U6537 (N_6537,N_5838,N_5354);
nand U6538 (N_6538,N_5391,N_5011);
and U6539 (N_6539,N_5460,N_5103);
or U6540 (N_6540,N_4075,N_5583);
nor U6541 (N_6541,N_4462,N_5311);
nor U6542 (N_6542,N_5581,N_4496);
or U6543 (N_6543,N_5697,N_5459);
nor U6544 (N_6544,N_4177,N_4247);
or U6545 (N_6545,N_4623,N_5916);
and U6546 (N_6546,N_5963,N_5299);
or U6547 (N_6547,N_4652,N_4403);
nor U6548 (N_6548,N_4638,N_4860);
nand U6549 (N_6549,N_5161,N_4029);
or U6550 (N_6550,N_5703,N_4828);
or U6551 (N_6551,N_4269,N_4669);
or U6552 (N_6552,N_4855,N_5830);
nand U6553 (N_6553,N_4291,N_4871);
or U6554 (N_6554,N_5182,N_5902);
and U6555 (N_6555,N_5575,N_5962);
xor U6556 (N_6556,N_4110,N_5243);
or U6557 (N_6557,N_5973,N_5390);
xnor U6558 (N_6558,N_4065,N_4318);
nor U6559 (N_6559,N_4681,N_4929);
or U6560 (N_6560,N_5613,N_4615);
or U6561 (N_6561,N_5803,N_5413);
nor U6562 (N_6562,N_5777,N_5064);
and U6563 (N_6563,N_5514,N_5658);
nand U6564 (N_6564,N_4151,N_5926);
or U6565 (N_6565,N_5324,N_5315);
or U6566 (N_6566,N_4169,N_4888);
xor U6567 (N_6567,N_4955,N_5412);
nand U6568 (N_6568,N_4412,N_5748);
nand U6569 (N_6569,N_5503,N_5485);
or U6570 (N_6570,N_5871,N_4516);
and U6571 (N_6571,N_5754,N_5466);
and U6572 (N_6572,N_5741,N_4509);
nand U6573 (N_6573,N_4098,N_4330);
or U6574 (N_6574,N_4056,N_4317);
xnor U6575 (N_6575,N_5646,N_5974);
and U6576 (N_6576,N_5855,N_5355);
or U6577 (N_6577,N_4368,N_5671);
nor U6578 (N_6578,N_5776,N_5300);
or U6579 (N_6579,N_5910,N_5112);
xor U6580 (N_6580,N_4479,N_5023);
or U6581 (N_6581,N_4751,N_5600);
nand U6582 (N_6582,N_5565,N_5863);
and U6583 (N_6583,N_4643,N_5951);
xor U6584 (N_6584,N_4779,N_4562);
nand U6585 (N_6585,N_5377,N_4856);
or U6586 (N_6586,N_4237,N_5693);
nand U6587 (N_6587,N_5155,N_4363);
nand U6588 (N_6588,N_4066,N_4734);
nor U6589 (N_6589,N_5009,N_5923);
xnor U6590 (N_6590,N_4141,N_4150);
and U6591 (N_6591,N_5559,N_5553);
nand U6592 (N_6592,N_5293,N_5191);
and U6593 (N_6593,N_5496,N_5196);
and U6594 (N_6594,N_4799,N_4705);
nand U6595 (N_6595,N_5661,N_4590);
xnor U6596 (N_6596,N_4166,N_4423);
xnor U6597 (N_6597,N_4980,N_5753);
and U6598 (N_6598,N_4474,N_5256);
and U6599 (N_6599,N_4924,N_5138);
or U6600 (N_6600,N_4867,N_4197);
xnor U6601 (N_6601,N_5567,N_5550);
or U6602 (N_6602,N_4687,N_4826);
nand U6603 (N_6603,N_4031,N_4901);
or U6604 (N_6604,N_5498,N_4821);
nand U6605 (N_6605,N_4267,N_4333);
xor U6606 (N_6606,N_5725,N_5761);
or U6607 (N_6607,N_4022,N_5331);
nand U6608 (N_6608,N_5333,N_5431);
and U6609 (N_6609,N_5558,N_4606);
or U6610 (N_6610,N_5547,N_4642);
xnor U6611 (N_6611,N_4259,N_5986);
or U6612 (N_6612,N_4749,N_4837);
and U6613 (N_6613,N_4484,N_4682);
and U6614 (N_6614,N_5070,N_5251);
nor U6615 (N_6615,N_4631,N_5454);
nor U6616 (N_6616,N_4025,N_4953);
xor U6617 (N_6617,N_5291,N_5900);
or U6618 (N_6618,N_5850,N_5174);
nand U6619 (N_6619,N_5461,N_4628);
nand U6620 (N_6620,N_4131,N_4180);
or U6621 (N_6621,N_4979,N_4994);
and U6622 (N_6622,N_4739,N_5204);
nand U6623 (N_6623,N_5228,N_5701);
and U6624 (N_6624,N_5060,N_4494);
nand U6625 (N_6625,N_5815,N_5405);
and U6626 (N_6626,N_5538,N_5945);
xor U6627 (N_6627,N_4233,N_5268);
nor U6628 (N_6628,N_5597,N_5066);
or U6629 (N_6629,N_5327,N_4521);
or U6630 (N_6630,N_4942,N_4258);
or U6631 (N_6631,N_4836,N_5511);
and U6632 (N_6632,N_4582,N_5426);
nor U6633 (N_6633,N_4219,N_4460);
nand U6634 (N_6634,N_5742,N_4878);
nand U6635 (N_6635,N_4174,N_4517);
nand U6636 (N_6636,N_4998,N_4706);
nand U6637 (N_6637,N_4809,N_5642);
nor U6638 (N_6638,N_4550,N_4649);
nor U6639 (N_6639,N_5861,N_5523);
nand U6640 (N_6640,N_4100,N_4402);
xor U6641 (N_6641,N_5542,N_4336);
nand U6642 (N_6642,N_5229,N_5589);
and U6643 (N_6643,N_4093,N_5423);
xor U6644 (N_6644,N_5490,N_5447);
nor U6645 (N_6645,N_4074,N_4731);
and U6646 (N_6646,N_4048,N_4123);
or U6647 (N_6647,N_5306,N_5520);
and U6648 (N_6648,N_5312,N_4284);
xor U6649 (N_6649,N_5035,N_4677);
nand U6650 (N_6650,N_5047,N_5976);
nand U6651 (N_6651,N_5226,N_5764);
or U6652 (N_6652,N_5527,N_4471);
nor U6653 (N_6653,N_4657,N_4846);
xnor U6654 (N_6654,N_4038,N_5757);
nor U6655 (N_6655,N_4349,N_5532);
and U6656 (N_6656,N_4861,N_5408);
xnor U6657 (N_6657,N_4250,N_4194);
nor U6658 (N_6658,N_5996,N_4122);
nand U6659 (N_6659,N_4140,N_5604);
xnor U6660 (N_6660,N_5370,N_5781);
xnor U6661 (N_6661,N_5914,N_4416);
nor U6662 (N_6662,N_5349,N_5934);
and U6663 (N_6663,N_4134,N_5819);
and U6664 (N_6664,N_5491,N_5669);
nor U6665 (N_6665,N_5346,N_4746);
xnor U6666 (N_6666,N_5267,N_5947);
nand U6667 (N_6667,N_4159,N_5786);
nor U6668 (N_6668,N_5687,N_4891);
and U6669 (N_6669,N_5281,N_5241);
or U6670 (N_6670,N_5571,N_4895);
nand U6671 (N_6671,N_5134,N_5302);
xor U6672 (N_6672,N_4903,N_5407);
or U6673 (N_6673,N_4595,N_5053);
and U6674 (N_6674,N_4823,N_4671);
and U6675 (N_6675,N_5842,N_4199);
nand U6676 (N_6676,N_4781,N_5006);
nand U6677 (N_6677,N_4523,N_5375);
nor U6678 (N_6678,N_5837,N_5101);
nor U6679 (N_6679,N_4546,N_4812);
xnor U6680 (N_6680,N_4511,N_5067);
nor U6681 (N_6681,N_4835,N_5937);
xnor U6682 (N_6682,N_5736,N_5056);
and U6683 (N_6683,N_5879,N_4338);
nand U6684 (N_6684,N_5061,N_5283);
or U6685 (N_6685,N_4228,N_4563);
xnor U6686 (N_6686,N_5233,N_5263);
nand U6687 (N_6687,N_4024,N_4076);
nor U6688 (N_6688,N_5297,N_5790);
xnor U6689 (N_6689,N_4000,N_4158);
nor U6690 (N_6690,N_5096,N_4109);
xnor U6691 (N_6691,N_5551,N_5663);
or U6692 (N_6692,N_4470,N_5335);
and U6693 (N_6693,N_5424,N_4567);
or U6694 (N_6694,N_4149,N_5367);
xor U6695 (N_6695,N_5920,N_4136);
or U6696 (N_6696,N_5328,N_4559);
nor U6697 (N_6697,N_5787,N_5702);
nand U6698 (N_6698,N_5752,N_4648);
nor U6699 (N_6699,N_4446,N_4921);
nand U6700 (N_6700,N_4108,N_5273);
nor U6701 (N_6701,N_5449,N_4490);
and U6702 (N_6702,N_5345,N_4204);
or U6703 (N_6703,N_4853,N_4121);
or U6704 (N_6704,N_5706,N_4192);
nor U6705 (N_6705,N_5007,N_5016);
and U6706 (N_6706,N_5779,N_5133);
nor U6707 (N_6707,N_5208,N_5844);
nand U6708 (N_6708,N_4906,N_4459);
or U6709 (N_6709,N_4106,N_5729);
and U6710 (N_6710,N_5392,N_5664);
xnor U6711 (N_6711,N_4329,N_5190);
or U6712 (N_6712,N_5927,N_4845);
and U6713 (N_6713,N_5782,N_4042);
nand U6714 (N_6714,N_5148,N_5242);
or U6715 (N_6715,N_5560,N_4565);
nor U6716 (N_6716,N_5119,N_4013);
xor U6717 (N_6717,N_4986,N_5353);
nor U6718 (N_6718,N_5362,N_4641);
or U6719 (N_6719,N_5090,N_4312);
and U6720 (N_6720,N_5188,N_4217);
or U6721 (N_6721,N_4544,N_5564);
or U6722 (N_6722,N_5114,N_4314);
nor U6723 (N_6723,N_4468,N_5869);
and U6724 (N_6724,N_4526,N_4586);
or U6725 (N_6725,N_5611,N_4769);
nor U6726 (N_6726,N_4251,N_4954);
and U6727 (N_6727,N_5794,N_5181);
xnor U6728 (N_6728,N_4473,N_5255);
and U6729 (N_6729,N_4240,N_4960);
xor U6730 (N_6730,N_5012,N_4039);
or U6731 (N_6731,N_5292,N_4659);
nor U6732 (N_6732,N_4607,N_5987);
or U6733 (N_6733,N_4545,N_4266);
and U6734 (N_6734,N_4275,N_4919);
or U6735 (N_6735,N_4822,N_5443);
xor U6736 (N_6736,N_5825,N_4055);
nand U6737 (N_6737,N_5026,N_4767);
nor U6738 (N_6738,N_4922,N_4295);
or U6739 (N_6739,N_4540,N_4229);
xor U6740 (N_6740,N_4033,N_5069);
or U6741 (N_6741,N_5183,N_5760);
nand U6742 (N_6742,N_4196,N_5343);
nor U6743 (N_6743,N_5163,N_5997);
nor U6744 (N_6744,N_5980,N_4495);
or U6745 (N_6745,N_4580,N_4365);
nand U6746 (N_6746,N_5832,N_4904);
nand U6747 (N_6747,N_4566,N_5686);
or U6748 (N_6748,N_5482,N_5798);
or U6749 (N_6749,N_5539,N_5042);
xnor U6750 (N_6750,N_4466,N_4362);
nand U6751 (N_6751,N_4300,N_5225);
xor U6752 (N_6752,N_4420,N_5179);
xor U6753 (N_6753,N_4418,N_5005);
and U6754 (N_6754,N_5595,N_4409);
xor U6755 (N_6755,N_5415,N_5540);
xor U6756 (N_6756,N_5873,N_5956);
and U6757 (N_6757,N_5590,N_5800);
or U6758 (N_6758,N_5036,N_5883);
and U6759 (N_6759,N_5807,N_4923);
or U6760 (N_6760,N_4392,N_5607);
or U6761 (N_6761,N_4857,N_5100);
and U6762 (N_6762,N_4918,N_4130);
nand U6763 (N_6763,N_5556,N_5195);
xnor U6764 (N_6764,N_4755,N_5500);
xnor U6765 (N_6765,N_4153,N_4092);
or U6766 (N_6766,N_4721,N_5258);
nand U6767 (N_6767,N_5359,N_4096);
nor U6768 (N_6768,N_4513,N_4868);
nor U6769 (N_6769,N_5314,N_5439);
nor U6770 (N_6770,N_4051,N_5528);
and U6771 (N_6771,N_4323,N_5334);
xor U6772 (N_6772,N_5193,N_5694);
nand U6773 (N_6773,N_4456,N_5046);
or U6774 (N_6774,N_4665,N_5820);
nand U6775 (N_6775,N_4622,N_4715);
or U6776 (N_6776,N_5624,N_5969);
xnor U6777 (N_6777,N_5892,N_5411);
nor U6778 (N_6778,N_4105,N_5457);
and U6779 (N_6779,N_4393,N_5058);
or U6780 (N_6780,N_5638,N_5382);
or U6781 (N_6781,N_5829,N_5504);
or U6782 (N_6782,N_4436,N_5082);
xor U6783 (N_6783,N_4366,N_4609);
or U6784 (N_6784,N_4030,N_4522);
nand U6785 (N_6785,N_4840,N_4438);
and U6786 (N_6786,N_4352,N_4383);
or U6787 (N_6787,N_4009,N_5895);
nand U6788 (N_6788,N_5866,N_4695);
nand U6789 (N_6789,N_4126,N_5698);
nand U6790 (N_6790,N_4137,N_4394);
nor U6791 (N_6791,N_5427,N_4289);
or U6792 (N_6792,N_4367,N_5360);
and U6793 (N_6793,N_4399,N_4850);
and U6794 (N_6794,N_5079,N_4560);
nor U6795 (N_6795,N_5115,N_5325);
or U6796 (N_6796,N_5157,N_4984);
xor U6797 (N_6797,N_4376,N_5506);
xnor U6798 (N_6798,N_4515,N_4493);
nand U6799 (N_6799,N_5513,N_5232);
nor U6800 (N_6800,N_4597,N_5579);
xor U6801 (N_6801,N_5479,N_5296);
xor U6802 (N_6802,N_4971,N_5141);
nand U6803 (N_6803,N_5903,N_4501);
or U6804 (N_6804,N_4012,N_4834);
or U6805 (N_6805,N_4617,N_5486);
nand U6806 (N_6806,N_4943,N_5990);
xnor U6807 (N_6807,N_4542,N_4455);
xnor U6808 (N_6808,N_4304,N_4730);
nor U6809 (N_6809,N_5904,N_4743);
and U6810 (N_6810,N_4359,N_5368);
nand U6811 (N_6811,N_4430,N_4803);
nor U6812 (N_6812,N_4232,N_4124);
xnor U6813 (N_6813,N_4691,N_5860);
xor U6814 (N_6814,N_4684,N_4010);
nand U6815 (N_6815,N_4307,N_5123);
and U6816 (N_6816,N_4078,N_4989);
xor U6817 (N_6817,N_4957,N_4975);
and U6818 (N_6818,N_5003,N_4967);
nand U6819 (N_6819,N_5197,N_5202);
nand U6820 (N_6820,N_5928,N_4805);
nand U6821 (N_6821,N_5145,N_5719);
nor U6822 (N_6822,N_4119,N_4696);
and U6823 (N_6823,N_4672,N_4449);
or U6824 (N_6824,N_5013,N_4792);
nand U6825 (N_6825,N_4796,N_4680);
nand U6826 (N_6826,N_4405,N_4016);
nor U6827 (N_6827,N_4326,N_4297);
xnor U6828 (N_6828,N_5683,N_4248);
or U6829 (N_6829,N_5121,N_4223);
or U6830 (N_6830,N_4435,N_5063);
nand U6831 (N_6831,N_5919,N_4018);
or U6832 (N_6832,N_4293,N_5107);
nor U6833 (N_6833,N_4839,N_5614);
or U6834 (N_6834,N_5120,N_4729);
nor U6835 (N_6835,N_5886,N_4740);
or U6836 (N_6836,N_4432,N_5656);
and U6837 (N_6837,N_5881,N_5076);
nor U6838 (N_6838,N_4773,N_4145);
and U6839 (N_6839,N_5244,N_5999);
or U6840 (N_6840,N_4949,N_4277);
xor U6841 (N_6841,N_4690,N_5716);
or U6842 (N_6842,N_5471,N_4161);
nand U6843 (N_6843,N_5518,N_4604);
nor U6844 (N_6844,N_4564,N_4630);
nand U6845 (N_6845,N_4209,N_5400);
nor U6846 (N_6846,N_5505,N_5203);
xor U6847 (N_6847,N_4741,N_5187);
nor U6848 (N_6848,N_5169,N_5469);
nand U6849 (N_6849,N_4238,N_4759);
nor U6850 (N_6850,N_5582,N_4313);
nor U6851 (N_6851,N_5922,N_4225);
nand U6852 (N_6852,N_4760,N_4735);
nor U6853 (N_6853,N_5321,N_5938);
xnor U6854 (N_6854,N_4281,N_4183);
nand U6855 (N_6855,N_5450,N_4833);
nand U6856 (N_6856,N_4481,N_5715);
xor U6857 (N_6857,N_4815,N_5991);
nor U6858 (N_6858,N_4072,N_4230);
nand U6859 (N_6859,N_5817,N_4504);
nor U6860 (N_6860,N_5030,N_4952);
nand U6861 (N_6861,N_4946,N_5236);
xor U6862 (N_6862,N_4662,N_4970);
and U6863 (N_6863,N_4348,N_4447);
nor U6864 (N_6864,N_4004,N_5810);
nor U6865 (N_6865,N_5674,N_5139);
or U6866 (N_6866,N_4614,N_4279);
xor U6867 (N_6867,N_4320,N_4235);
nand U6868 (N_6868,N_4469,N_5843);
nand U6869 (N_6869,N_4569,N_5770);
nor U6870 (N_6870,N_5744,N_5530);
nor U6871 (N_6871,N_5219,N_5822);
nor U6872 (N_6872,N_5262,N_4285);
xnor U6873 (N_6873,N_4212,N_4543);
or U6874 (N_6874,N_4621,N_5899);
nor U6875 (N_6875,N_5025,N_5602);
nor U6876 (N_6876,N_4536,N_4189);
and U6877 (N_6877,N_5164,N_5033);
nor U6878 (N_6878,N_4185,N_4510);
and U6879 (N_6879,N_5929,N_5501);
and U6880 (N_6880,N_5344,N_5143);
xnor U6881 (N_6881,N_4309,N_5379);
nor U6882 (N_6882,N_5509,N_5259);
xor U6883 (N_6883,N_4132,N_5441);
nand U6884 (N_6884,N_4911,N_4026);
and U6885 (N_6885,N_5940,N_5192);
nand U6886 (N_6886,N_5510,N_5051);
nand U6887 (N_6887,N_5109,N_5576);
nand U6888 (N_6888,N_5865,N_4678);
and U6889 (N_6889,N_4099,N_5918);
nor U6890 (N_6890,N_5637,N_4445);
nand U6891 (N_6891,N_5679,N_5970);
nand U6892 (N_6892,N_4538,N_4035);
xnor U6893 (N_6893,N_4507,N_4961);
nor U6894 (N_6894,N_5588,N_4959);
xor U6895 (N_6895,N_4041,N_5876);
and U6896 (N_6896,N_4461,N_5731);
or U6897 (N_6897,N_4427,N_4754);
and U6898 (N_6898,N_5309,N_5223);
and U6899 (N_6899,N_4658,N_5052);
xnor U6900 (N_6900,N_5901,N_4306);
or U6901 (N_6901,N_4373,N_4205);
nand U6902 (N_6902,N_5253,N_4700);
nand U6903 (N_6903,N_4692,N_4807);
or U6904 (N_6904,N_5890,N_4073);
or U6905 (N_6905,N_5771,N_4829);
or U6906 (N_6906,N_5433,N_4708);
xor U6907 (N_6907,N_5911,N_4424);
xnor U6908 (N_6908,N_5828,N_5948);
or U6909 (N_6909,N_5751,N_4286);
xnor U6910 (N_6910,N_5448,N_5979);
nor U6911 (N_6911,N_4518,N_5982);
and U6912 (N_6912,N_5628,N_5352);
nor U6913 (N_6913,N_5420,N_5801);
nor U6914 (N_6914,N_5166,N_5954);
or U6915 (N_6915,N_4723,N_4736);
nand U6916 (N_6916,N_4211,N_5137);
and U6917 (N_6917,N_4360,N_5317);
xor U6918 (N_6918,N_4847,N_5480);
and U6919 (N_6919,N_5649,N_5961);
nand U6920 (N_6920,N_4015,N_5421);
nor U6921 (N_6921,N_5440,N_4804);
and U6922 (N_6922,N_5444,N_5906);
xor U6923 (N_6923,N_5260,N_5396);
xnor U6924 (N_6924,N_5111,N_5568);
and U6925 (N_6925,N_4006,N_5481);
nand U6926 (N_6926,N_4945,N_4624);
xor U6927 (N_6927,N_4344,N_4968);
nand U6928 (N_6928,N_5086,N_5494);
xnor U6929 (N_6929,N_4774,N_4733);
or U6930 (N_6930,N_5059,N_5738);
nor U6931 (N_6931,N_5950,N_5644);
or U6932 (N_6932,N_5710,N_4458);
and U6933 (N_6933,N_4148,N_5125);
nand U6934 (N_6934,N_5227,N_4972);
nor U6935 (N_6935,N_5641,N_4472);
xnor U6936 (N_6936,N_5652,N_5414);
nor U6937 (N_6937,N_4273,N_4179);
xor U6938 (N_6938,N_4287,N_4934);
nor U6939 (N_6939,N_4112,N_5356);
and U6940 (N_6940,N_4948,N_5097);
xor U6941 (N_6941,N_5144,N_4583);
or U6942 (N_6942,N_4650,N_5972);
and U6943 (N_6943,N_5322,N_4221);
or U6944 (N_6944,N_4419,N_5591);
or U6945 (N_6945,N_4514,N_5755);
and U6946 (N_6946,N_4787,N_5864);
and U6947 (N_6947,N_5756,N_4090);
nand U6948 (N_6948,N_4524,N_4308);
nand U6949 (N_6949,N_4028,N_5150);
and U6950 (N_6950,N_4699,N_5784);
nor U6951 (N_6951,N_4585,N_5636);
and U6952 (N_6952,N_5329,N_4094);
xnor U6953 (N_6953,N_4503,N_5230);
or U6954 (N_6954,N_4271,N_5304);
and U6955 (N_6955,N_4786,N_4276);
or U6956 (N_6956,N_5905,N_5623);
nor U6957 (N_6957,N_5087,N_4801);
nand U6958 (N_6958,N_4227,N_4578);
or U6959 (N_6959,N_4797,N_5434);
or U6960 (N_6960,N_5495,N_4885);
and U6961 (N_6961,N_4357,N_5629);
nand U6962 (N_6962,N_5983,N_5478);
nor U6963 (N_6963,N_4220,N_5406);
or U6964 (N_6964,N_4454,N_5027);
nand U6965 (N_6965,N_5062,N_5184);
xor U6966 (N_6966,N_4541,N_4762);
or U6967 (N_6967,N_5826,N_5124);
xnor U6968 (N_6968,N_5849,N_5366);
nand U6969 (N_6969,N_4808,N_4646);
xor U6970 (N_6970,N_4152,N_5221);
nor U6971 (N_6971,N_4777,N_5394);
or U6972 (N_6972,N_4719,N_4014);
nor U6973 (N_6973,N_4827,N_5533);
or U6974 (N_6974,N_4770,N_4732);
nand U6975 (N_6975,N_5468,N_4547);
nand U6976 (N_6976,N_4415,N_5944);
or U6977 (N_6977,N_5338,N_4067);
nor U6978 (N_6978,N_5908,N_5275);
nor U6979 (N_6979,N_5824,N_5966);
or U6980 (N_6980,N_4794,N_5626);
nor U6981 (N_6981,N_4480,N_5254);
nand U6982 (N_6982,N_4144,N_5357);
or U6983 (N_6983,N_4532,N_4270);
or U6984 (N_6984,N_5089,N_4282);
nand U6985 (N_6985,N_4838,N_5266);
xnor U6986 (N_6986,N_4783,N_4618);
nand U6987 (N_6987,N_4115,N_5692);
xnor U6988 (N_6988,N_5816,N_4385);
and U6989 (N_6989,N_4988,N_5218);
and U6990 (N_6990,N_4175,N_5041);
nor U6991 (N_6991,N_4477,N_5465);
nor U6992 (N_6992,N_4256,N_5857);
xor U6993 (N_6993,N_5939,N_4784);
and U6994 (N_6994,N_5723,N_5587);
nand U6995 (N_6995,N_5846,N_5526);
and U6996 (N_6996,N_4214,N_5290);
or U6997 (N_6997,N_4382,N_4963);
nand U6998 (N_6998,N_4260,N_4581);
xnor U6999 (N_6999,N_5666,N_5165);
nor U7000 (N_7000,N_4039,N_5453);
xor U7001 (N_7001,N_5119,N_4923);
nor U7002 (N_7002,N_5353,N_5024);
nor U7003 (N_7003,N_5275,N_4047);
nand U7004 (N_7004,N_4321,N_4288);
nor U7005 (N_7005,N_4736,N_4973);
nand U7006 (N_7006,N_4156,N_5861);
xnor U7007 (N_7007,N_4759,N_5364);
and U7008 (N_7008,N_5394,N_4191);
nand U7009 (N_7009,N_4917,N_4312);
and U7010 (N_7010,N_4175,N_4380);
xor U7011 (N_7011,N_4413,N_5568);
or U7012 (N_7012,N_5591,N_4920);
or U7013 (N_7013,N_4728,N_4163);
or U7014 (N_7014,N_5241,N_4979);
nor U7015 (N_7015,N_4284,N_5751);
xnor U7016 (N_7016,N_5812,N_4231);
nor U7017 (N_7017,N_5155,N_5798);
and U7018 (N_7018,N_4251,N_4078);
and U7019 (N_7019,N_5983,N_5902);
or U7020 (N_7020,N_4618,N_4801);
nor U7021 (N_7021,N_5662,N_4646);
or U7022 (N_7022,N_4393,N_5520);
or U7023 (N_7023,N_4045,N_5215);
xor U7024 (N_7024,N_4045,N_5769);
nand U7025 (N_7025,N_5171,N_4728);
xnor U7026 (N_7026,N_5264,N_5657);
or U7027 (N_7027,N_5389,N_5280);
xnor U7028 (N_7028,N_4447,N_4905);
nor U7029 (N_7029,N_4306,N_4226);
or U7030 (N_7030,N_4306,N_5982);
or U7031 (N_7031,N_5541,N_4259);
nand U7032 (N_7032,N_4741,N_4125);
and U7033 (N_7033,N_5422,N_4073);
xor U7034 (N_7034,N_4425,N_5512);
nor U7035 (N_7035,N_5991,N_5266);
xnor U7036 (N_7036,N_5294,N_4621);
or U7037 (N_7037,N_4917,N_4952);
and U7038 (N_7038,N_5820,N_5238);
and U7039 (N_7039,N_4631,N_5481);
nor U7040 (N_7040,N_5361,N_5654);
and U7041 (N_7041,N_5562,N_5785);
nor U7042 (N_7042,N_4951,N_4573);
xor U7043 (N_7043,N_5829,N_4383);
and U7044 (N_7044,N_5041,N_5473);
nor U7045 (N_7045,N_4502,N_5836);
nor U7046 (N_7046,N_5929,N_5199);
and U7047 (N_7047,N_4099,N_4743);
and U7048 (N_7048,N_4210,N_5302);
or U7049 (N_7049,N_5439,N_4531);
and U7050 (N_7050,N_4184,N_4156);
nor U7051 (N_7051,N_4642,N_4429);
xor U7052 (N_7052,N_4071,N_5843);
and U7053 (N_7053,N_4765,N_4616);
nand U7054 (N_7054,N_4035,N_5449);
and U7055 (N_7055,N_4107,N_5095);
or U7056 (N_7056,N_4535,N_5707);
nor U7057 (N_7057,N_5269,N_4871);
nor U7058 (N_7058,N_4683,N_5522);
xnor U7059 (N_7059,N_4964,N_5830);
xnor U7060 (N_7060,N_4730,N_4521);
nand U7061 (N_7061,N_5928,N_5365);
or U7062 (N_7062,N_4660,N_4149);
nor U7063 (N_7063,N_4513,N_5393);
and U7064 (N_7064,N_5749,N_5950);
and U7065 (N_7065,N_5588,N_5071);
nor U7066 (N_7066,N_5576,N_4725);
or U7067 (N_7067,N_5398,N_5095);
nor U7068 (N_7068,N_5487,N_5678);
and U7069 (N_7069,N_5906,N_4424);
xnor U7070 (N_7070,N_4459,N_5154);
xor U7071 (N_7071,N_4696,N_5702);
xor U7072 (N_7072,N_4738,N_5258);
nor U7073 (N_7073,N_5650,N_4869);
nand U7074 (N_7074,N_4405,N_5803);
nor U7075 (N_7075,N_4527,N_5063);
nor U7076 (N_7076,N_5736,N_4021);
nand U7077 (N_7077,N_5405,N_5982);
nand U7078 (N_7078,N_5535,N_4480);
nand U7079 (N_7079,N_5749,N_5316);
nand U7080 (N_7080,N_4589,N_5620);
nand U7081 (N_7081,N_4177,N_4046);
nand U7082 (N_7082,N_4580,N_4766);
nor U7083 (N_7083,N_4297,N_5444);
and U7084 (N_7084,N_5255,N_4854);
and U7085 (N_7085,N_5912,N_5913);
nand U7086 (N_7086,N_4160,N_4360);
xnor U7087 (N_7087,N_5637,N_5659);
nand U7088 (N_7088,N_4179,N_5827);
and U7089 (N_7089,N_5621,N_4259);
nand U7090 (N_7090,N_5876,N_5779);
and U7091 (N_7091,N_4266,N_4578);
xnor U7092 (N_7092,N_4512,N_4184);
nor U7093 (N_7093,N_5588,N_5422);
and U7094 (N_7094,N_5452,N_5210);
xnor U7095 (N_7095,N_5359,N_4412);
nor U7096 (N_7096,N_4282,N_5262);
and U7097 (N_7097,N_4285,N_5343);
or U7098 (N_7098,N_4699,N_5876);
and U7099 (N_7099,N_5232,N_5723);
nand U7100 (N_7100,N_5793,N_4825);
nor U7101 (N_7101,N_4162,N_4485);
nand U7102 (N_7102,N_5991,N_5358);
and U7103 (N_7103,N_5684,N_4103);
nor U7104 (N_7104,N_5601,N_4452);
nor U7105 (N_7105,N_5453,N_4473);
xnor U7106 (N_7106,N_5430,N_5413);
and U7107 (N_7107,N_4214,N_5068);
or U7108 (N_7108,N_4782,N_5947);
nand U7109 (N_7109,N_4821,N_4326);
or U7110 (N_7110,N_5036,N_4321);
nor U7111 (N_7111,N_4673,N_5359);
and U7112 (N_7112,N_4975,N_4086);
nand U7113 (N_7113,N_4699,N_5363);
or U7114 (N_7114,N_5229,N_4800);
and U7115 (N_7115,N_4997,N_5821);
nor U7116 (N_7116,N_4300,N_5001);
xnor U7117 (N_7117,N_5100,N_4621);
xnor U7118 (N_7118,N_5082,N_4704);
nand U7119 (N_7119,N_4220,N_5690);
xor U7120 (N_7120,N_4336,N_5599);
nand U7121 (N_7121,N_4042,N_4050);
nor U7122 (N_7122,N_4038,N_5455);
nand U7123 (N_7123,N_5795,N_5127);
nor U7124 (N_7124,N_5065,N_5098);
or U7125 (N_7125,N_5842,N_5230);
and U7126 (N_7126,N_4025,N_5402);
nor U7127 (N_7127,N_5077,N_5830);
and U7128 (N_7128,N_4930,N_4205);
nor U7129 (N_7129,N_5436,N_4092);
and U7130 (N_7130,N_4430,N_4318);
xor U7131 (N_7131,N_5362,N_5513);
or U7132 (N_7132,N_5342,N_5055);
xnor U7133 (N_7133,N_5636,N_4662);
or U7134 (N_7134,N_4439,N_5659);
xnor U7135 (N_7135,N_4626,N_5634);
xor U7136 (N_7136,N_4051,N_4765);
and U7137 (N_7137,N_4675,N_5981);
nor U7138 (N_7138,N_5878,N_4203);
nand U7139 (N_7139,N_4294,N_4408);
nand U7140 (N_7140,N_5031,N_5440);
or U7141 (N_7141,N_4939,N_4923);
or U7142 (N_7142,N_4990,N_5032);
and U7143 (N_7143,N_4773,N_5168);
or U7144 (N_7144,N_5127,N_4850);
xor U7145 (N_7145,N_5418,N_5953);
and U7146 (N_7146,N_5361,N_5925);
nand U7147 (N_7147,N_5157,N_4338);
xor U7148 (N_7148,N_4023,N_4814);
nand U7149 (N_7149,N_4626,N_5959);
nand U7150 (N_7150,N_4048,N_5084);
nand U7151 (N_7151,N_4486,N_4531);
and U7152 (N_7152,N_4070,N_4283);
nor U7153 (N_7153,N_4125,N_4071);
nor U7154 (N_7154,N_4939,N_4128);
xnor U7155 (N_7155,N_4774,N_4369);
nand U7156 (N_7156,N_5335,N_5256);
nor U7157 (N_7157,N_5106,N_5437);
and U7158 (N_7158,N_4919,N_4383);
or U7159 (N_7159,N_4595,N_5870);
or U7160 (N_7160,N_4337,N_4741);
xor U7161 (N_7161,N_4374,N_5462);
nor U7162 (N_7162,N_5645,N_5510);
nor U7163 (N_7163,N_5275,N_4452);
xnor U7164 (N_7164,N_5863,N_5695);
nor U7165 (N_7165,N_5008,N_5468);
nand U7166 (N_7166,N_4533,N_5318);
nor U7167 (N_7167,N_4221,N_4636);
and U7168 (N_7168,N_4702,N_4645);
nand U7169 (N_7169,N_5224,N_4734);
nand U7170 (N_7170,N_5996,N_4563);
nand U7171 (N_7171,N_4861,N_5074);
nand U7172 (N_7172,N_5757,N_5414);
xnor U7173 (N_7173,N_4268,N_4692);
nor U7174 (N_7174,N_5795,N_5386);
or U7175 (N_7175,N_4954,N_4476);
nand U7176 (N_7176,N_4468,N_4994);
nor U7177 (N_7177,N_5170,N_5938);
and U7178 (N_7178,N_5475,N_4931);
or U7179 (N_7179,N_5383,N_4915);
xnor U7180 (N_7180,N_5594,N_5961);
nand U7181 (N_7181,N_5055,N_4939);
nand U7182 (N_7182,N_4144,N_5674);
nor U7183 (N_7183,N_5792,N_4355);
nand U7184 (N_7184,N_4376,N_4424);
and U7185 (N_7185,N_5806,N_5724);
and U7186 (N_7186,N_4313,N_4060);
or U7187 (N_7187,N_4178,N_5564);
nand U7188 (N_7188,N_4816,N_4529);
nand U7189 (N_7189,N_5370,N_5473);
nor U7190 (N_7190,N_5897,N_5097);
nor U7191 (N_7191,N_4839,N_5961);
nor U7192 (N_7192,N_4956,N_5127);
and U7193 (N_7193,N_4892,N_4389);
and U7194 (N_7194,N_4046,N_4186);
xor U7195 (N_7195,N_4311,N_5257);
xor U7196 (N_7196,N_4738,N_4197);
and U7197 (N_7197,N_4825,N_5896);
nand U7198 (N_7198,N_5926,N_5908);
and U7199 (N_7199,N_4971,N_5859);
or U7200 (N_7200,N_5932,N_5730);
or U7201 (N_7201,N_4762,N_5722);
nor U7202 (N_7202,N_5341,N_5462);
nor U7203 (N_7203,N_4659,N_4438);
nand U7204 (N_7204,N_5506,N_5632);
xor U7205 (N_7205,N_4507,N_4096);
nand U7206 (N_7206,N_4689,N_4819);
or U7207 (N_7207,N_4340,N_4816);
xnor U7208 (N_7208,N_5362,N_4060);
nand U7209 (N_7209,N_4759,N_4406);
and U7210 (N_7210,N_4761,N_4151);
nor U7211 (N_7211,N_5212,N_5291);
nor U7212 (N_7212,N_4867,N_4730);
nand U7213 (N_7213,N_4617,N_4077);
and U7214 (N_7214,N_5590,N_4472);
nand U7215 (N_7215,N_4153,N_5759);
or U7216 (N_7216,N_5421,N_5294);
and U7217 (N_7217,N_5728,N_4507);
nand U7218 (N_7218,N_4100,N_5634);
nand U7219 (N_7219,N_5983,N_4734);
and U7220 (N_7220,N_5211,N_4521);
xor U7221 (N_7221,N_5957,N_4993);
nor U7222 (N_7222,N_4196,N_5788);
nor U7223 (N_7223,N_5667,N_5142);
xnor U7224 (N_7224,N_4664,N_4331);
or U7225 (N_7225,N_5587,N_5672);
nor U7226 (N_7226,N_4597,N_5488);
nand U7227 (N_7227,N_4038,N_4583);
nor U7228 (N_7228,N_4229,N_4335);
and U7229 (N_7229,N_4165,N_4445);
and U7230 (N_7230,N_4497,N_5831);
nor U7231 (N_7231,N_5990,N_4965);
or U7232 (N_7232,N_4750,N_4918);
and U7233 (N_7233,N_5571,N_5229);
nor U7234 (N_7234,N_4964,N_5800);
nand U7235 (N_7235,N_5996,N_5257);
or U7236 (N_7236,N_5485,N_5024);
nor U7237 (N_7237,N_4030,N_4150);
xnor U7238 (N_7238,N_5114,N_5051);
xnor U7239 (N_7239,N_5566,N_5275);
nand U7240 (N_7240,N_5416,N_5082);
or U7241 (N_7241,N_4168,N_5476);
and U7242 (N_7242,N_4731,N_5772);
nor U7243 (N_7243,N_5907,N_4215);
nor U7244 (N_7244,N_4117,N_5690);
nor U7245 (N_7245,N_5804,N_5757);
xor U7246 (N_7246,N_5106,N_5407);
and U7247 (N_7247,N_4656,N_4119);
and U7248 (N_7248,N_4648,N_4146);
and U7249 (N_7249,N_5759,N_4069);
or U7250 (N_7250,N_5612,N_4124);
or U7251 (N_7251,N_4271,N_4583);
nand U7252 (N_7252,N_5707,N_5533);
nand U7253 (N_7253,N_4885,N_4118);
nand U7254 (N_7254,N_4429,N_4225);
xnor U7255 (N_7255,N_5440,N_4394);
xor U7256 (N_7256,N_5010,N_4739);
or U7257 (N_7257,N_5741,N_5686);
nand U7258 (N_7258,N_4355,N_5629);
xor U7259 (N_7259,N_4542,N_5933);
nor U7260 (N_7260,N_5343,N_5543);
nor U7261 (N_7261,N_5365,N_5205);
or U7262 (N_7262,N_4371,N_4946);
nor U7263 (N_7263,N_5412,N_4468);
and U7264 (N_7264,N_4760,N_4278);
xor U7265 (N_7265,N_4738,N_5064);
nor U7266 (N_7266,N_4411,N_5139);
or U7267 (N_7267,N_4767,N_5850);
nor U7268 (N_7268,N_5535,N_4739);
xnor U7269 (N_7269,N_4671,N_5885);
xnor U7270 (N_7270,N_4659,N_4523);
or U7271 (N_7271,N_4092,N_5176);
and U7272 (N_7272,N_4734,N_4075);
nor U7273 (N_7273,N_5675,N_5884);
nand U7274 (N_7274,N_4144,N_4087);
nand U7275 (N_7275,N_4822,N_5253);
nand U7276 (N_7276,N_4642,N_5401);
or U7277 (N_7277,N_4101,N_5631);
nand U7278 (N_7278,N_4447,N_5640);
nor U7279 (N_7279,N_4417,N_5035);
nand U7280 (N_7280,N_4686,N_4327);
xor U7281 (N_7281,N_4746,N_4702);
nor U7282 (N_7282,N_5095,N_5075);
or U7283 (N_7283,N_5394,N_4516);
nand U7284 (N_7284,N_4376,N_5175);
nand U7285 (N_7285,N_4593,N_4135);
and U7286 (N_7286,N_5493,N_5286);
xnor U7287 (N_7287,N_4389,N_5196);
or U7288 (N_7288,N_4707,N_4613);
xnor U7289 (N_7289,N_4506,N_4471);
xnor U7290 (N_7290,N_5487,N_4707);
xnor U7291 (N_7291,N_4813,N_5228);
or U7292 (N_7292,N_5800,N_5324);
or U7293 (N_7293,N_5857,N_4170);
xnor U7294 (N_7294,N_4472,N_4833);
or U7295 (N_7295,N_4575,N_4572);
and U7296 (N_7296,N_4164,N_5435);
or U7297 (N_7297,N_4445,N_4662);
and U7298 (N_7298,N_5847,N_4151);
nand U7299 (N_7299,N_5087,N_4091);
nor U7300 (N_7300,N_5633,N_4380);
nand U7301 (N_7301,N_4692,N_4389);
nand U7302 (N_7302,N_5248,N_4162);
and U7303 (N_7303,N_4158,N_5191);
and U7304 (N_7304,N_5112,N_5010);
nor U7305 (N_7305,N_4491,N_5931);
nor U7306 (N_7306,N_4836,N_5267);
nor U7307 (N_7307,N_5356,N_5917);
nor U7308 (N_7308,N_5225,N_5357);
nand U7309 (N_7309,N_4373,N_5938);
and U7310 (N_7310,N_5750,N_4408);
nor U7311 (N_7311,N_4945,N_5729);
nor U7312 (N_7312,N_5982,N_4536);
nand U7313 (N_7313,N_5043,N_4603);
and U7314 (N_7314,N_4442,N_4702);
nand U7315 (N_7315,N_5737,N_4307);
xor U7316 (N_7316,N_4728,N_4276);
and U7317 (N_7317,N_5333,N_4508);
or U7318 (N_7318,N_4605,N_5627);
nand U7319 (N_7319,N_4871,N_5767);
nor U7320 (N_7320,N_4379,N_5241);
nand U7321 (N_7321,N_4041,N_4080);
nand U7322 (N_7322,N_5740,N_5076);
and U7323 (N_7323,N_4407,N_4770);
xnor U7324 (N_7324,N_5122,N_5316);
xor U7325 (N_7325,N_4594,N_5922);
and U7326 (N_7326,N_5128,N_4720);
or U7327 (N_7327,N_4748,N_4714);
or U7328 (N_7328,N_5174,N_4817);
and U7329 (N_7329,N_4771,N_5509);
xor U7330 (N_7330,N_4372,N_4599);
or U7331 (N_7331,N_5907,N_4821);
or U7332 (N_7332,N_5122,N_4498);
or U7333 (N_7333,N_4050,N_4066);
nand U7334 (N_7334,N_5195,N_4520);
and U7335 (N_7335,N_4618,N_4687);
xor U7336 (N_7336,N_5077,N_4625);
nand U7337 (N_7337,N_4675,N_4891);
or U7338 (N_7338,N_5907,N_4629);
and U7339 (N_7339,N_5754,N_5706);
xnor U7340 (N_7340,N_4489,N_5791);
and U7341 (N_7341,N_4870,N_5667);
xnor U7342 (N_7342,N_5755,N_4977);
and U7343 (N_7343,N_4891,N_4829);
or U7344 (N_7344,N_4739,N_5799);
nand U7345 (N_7345,N_5098,N_4185);
nand U7346 (N_7346,N_4665,N_5043);
nor U7347 (N_7347,N_5839,N_4843);
nand U7348 (N_7348,N_4190,N_5707);
nor U7349 (N_7349,N_5271,N_4588);
nor U7350 (N_7350,N_5859,N_4126);
and U7351 (N_7351,N_5682,N_4399);
nor U7352 (N_7352,N_5253,N_4236);
or U7353 (N_7353,N_4970,N_4500);
nand U7354 (N_7354,N_5717,N_4533);
or U7355 (N_7355,N_5554,N_4844);
or U7356 (N_7356,N_5798,N_5189);
nor U7357 (N_7357,N_5876,N_5571);
nand U7358 (N_7358,N_4239,N_4847);
and U7359 (N_7359,N_5271,N_5101);
nand U7360 (N_7360,N_4932,N_4033);
and U7361 (N_7361,N_5322,N_4298);
xor U7362 (N_7362,N_5846,N_4394);
nor U7363 (N_7363,N_4684,N_5342);
xnor U7364 (N_7364,N_4141,N_4474);
and U7365 (N_7365,N_4798,N_5457);
and U7366 (N_7366,N_5634,N_4857);
nand U7367 (N_7367,N_4243,N_5622);
or U7368 (N_7368,N_5585,N_5237);
xnor U7369 (N_7369,N_5108,N_5139);
nand U7370 (N_7370,N_4837,N_4107);
and U7371 (N_7371,N_4244,N_5254);
or U7372 (N_7372,N_4441,N_4681);
and U7373 (N_7373,N_5164,N_4955);
and U7374 (N_7374,N_5643,N_4923);
xnor U7375 (N_7375,N_5324,N_4121);
nor U7376 (N_7376,N_5072,N_5442);
and U7377 (N_7377,N_5150,N_4250);
or U7378 (N_7378,N_5048,N_5903);
nand U7379 (N_7379,N_4361,N_5232);
xor U7380 (N_7380,N_4866,N_4135);
nand U7381 (N_7381,N_5132,N_4695);
and U7382 (N_7382,N_5609,N_5184);
nor U7383 (N_7383,N_5383,N_4508);
and U7384 (N_7384,N_4160,N_5956);
and U7385 (N_7385,N_5225,N_4695);
xnor U7386 (N_7386,N_4883,N_4367);
xor U7387 (N_7387,N_5613,N_5677);
nor U7388 (N_7388,N_4621,N_5641);
nor U7389 (N_7389,N_5131,N_5695);
nand U7390 (N_7390,N_4635,N_4905);
nand U7391 (N_7391,N_5601,N_5154);
nand U7392 (N_7392,N_5426,N_5676);
nand U7393 (N_7393,N_5833,N_5723);
and U7394 (N_7394,N_5485,N_4246);
nor U7395 (N_7395,N_5788,N_5449);
or U7396 (N_7396,N_5871,N_4376);
and U7397 (N_7397,N_4894,N_4541);
xor U7398 (N_7398,N_5380,N_5377);
nand U7399 (N_7399,N_5337,N_5335);
and U7400 (N_7400,N_5962,N_5228);
and U7401 (N_7401,N_5457,N_5205);
and U7402 (N_7402,N_4492,N_4232);
or U7403 (N_7403,N_5307,N_4891);
xnor U7404 (N_7404,N_5820,N_5960);
nand U7405 (N_7405,N_4609,N_5959);
nand U7406 (N_7406,N_4885,N_4568);
nor U7407 (N_7407,N_5978,N_4938);
and U7408 (N_7408,N_5312,N_5819);
nand U7409 (N_7409,N_5373,N_5579);
nor U7410 (N_7410,N_5326,N_4241);
nor U7411 (N_7411,N_5886,N_4622);
or U7412 (N_7412,N_4290,N_4434);
and U7413 (N_7413,N_5603,N_5117);
nand U7414 (N_7414,N_5140,N_5502);
and U7415 (N_7415,N_5995,N_4047);
or U7416 (N_7416,N_4249,N_5264);
nor U7417 (N_7417,N_5821,N_5080);
xor U7418 (N_7418,N_4512,N_4255);
and U7419 (N_7419,N_5968,N_5427);
nor U7420 (N_7420,N_5588,N_4315);
nor U7421 (N_7421,N_5643,N_5881);
and U7422 (N_7422,N_5413,N_4504);
or U7423 (N_7423,N_4514,N_4063);
nand U7424 (N_7424,N_5356,N_5507);
nor U7425 (N_7425,N_5248,N_5563);
xnor U7426 (N_7426,N_5468,N_5987);
xnor U7427 (N_7427,N_5452,N_4903);
or U7428 (N_7428,N_4471,N_4687);
and U7429 (N_7429,N_5457,N_5266);
xor U7430 (N_7430,N_4695,N_5850);
xnor U7431 (N_7431,N_5503,N_5976);
nor U7432 (N_7432,N_4708,N_4655);
or U7433 (N_7433,N_4696,N_5700);
and U7434 (N_7434,N_4004,N_5666);
nand U7435 (N_7435,N_4065,N_4257);
nor U7436 (N_7436,N_4600,N_5466);
xor U7437 (N_7437,N_5446,N_5930);
or U7438 (N_7438,N_4089,N_5263);
and U7439 (N_7439,N_5182,N_4884);
xnor U7440 (N_7440,N_4614,N_4226);
nor U7441 (N_7441,N_4699,N_4663);
or U7442 (N_7442,N_5682,N_4460);
nor U7443 (N_7443,N_5918,N_4897);
nand U7444 (N_7444,N_4427,N_4065);
or U7445 (N_7445,N_4332,N_5735);
or U7446 (N_7446,N_5179,N_4229);
nor U7447 (N_7447,N_4385,N_5540);
xnor U7448 (N_7448,N_4112,N_5857);
xnor U7449 (N_7449,N_4566,N_4950);
xor U7450 (N_7450,N_4871,N_4746);
and U7451 (N_7451,N_4804,N_4213);
xnor U7452 (N_7452,N_4261,N_5855);
nand U7453 (N_7453,N_4649,N_5972);
or U7454 (N_7454,N_4076,N_5323);
xnor U7455 (N_7455,N_4982,N_4514);
nor U7456 (N_7456,N_5110,N_5356);
nand U7457 (N_7457,N_4685,N_4831);
nor U7458 (N_7458,N_5043,N_4288);
nor U7459 (N_7459,N_4556,N_4893);
xnor U7460 (N_7460,N_4381,N_4798);
nand U7461 (N_7461,N_4672,N_5109);
or U7462 (N_7462,N_5698,N_5082);
nor U7463 (N_7463,N_5556,N_4464);
nor U7464 (N_7464,N_4183,N_4382);
nand U7465 (N_7465,N_4984,N_4762);
and U7466 (N_7466,N_4810,N_5550);
xor U7467 (N_7467,N_5966,N_5400);
and U7468 (N_7468,N_4385,N_4016);
nor U7469 (N_7469,N_5943,N_4350);
nor U7470 (N_7470,N_4897,N_5245);
xor U7471 (N_7471,N_4426,N_5822);
xor U7472 (N_7472,N_5843,N_4534);
nor U7473 (N_7473,N_4195,N_5467);
xor U7474 (N_7474,N_4891,N_5024);
nor U7475 (N_7475,N_4212,N_5759);
nor U7476 (N_7476,N_5757,N_5425);
nor U7477 (N_7477,N_4333,N_4720);
or U7478 (N_7478,N_4656,N_4824);
nand U7479 (N_7479,N_5226,N_4723);
nand U7480 (N_7480,N_4767,N_5241);
nor U7481 (N_7481,N_5526,N_5430);
xnor U7482 (N_7482,N_4048,N_4570);
nor U7483 (N_7483,N_4420,N_5997);
nor U7484 (N_7484,N_5468,N_4756);
or U7485 (N_7485,N_5971,N_4880);
nand U7486 (N_7486,N_4083,N_4175);
and U7487 (N_7487,N_4523,N_5460);
nand U7488 (N_7488,N_4688,N_5270);
nor U7489 (N_7489,N_5711,N_5828);
nand U7490 (N_7490,N_5629,N_4494);
xnor U7491 (N_7491,N_5562,N_4755);
nor U7492 (N_7492,N_4792,N_4819);
or U7493 (N_7493,N_4938,N_5944);
or U7494 (N_7494,N_4190,N_4083);
nand U7495 (N_7495,N_5209,N_5983);
nand U7496 (N_7496,N_4787,N_5231);
xor U7497 (N_7497,N_5512,N_4789);
or U7498 (N_7498,N_4066,N_5876);
or U7499 (N_7499,N_5751,N_4441);
nor U7500 (N_7500,N_4220,N_4723);
xor U7501 (N_7501,N_5535,N_4295);
xnor U7502 (N_7502,N_5978,N_5805);
xor U7503 (N_7503,N_5690,N_5059);
xnor U7504 (N_7504,N_4858,N_4288);
xnor U7505 (N_7505,N_5492,N_4098);
nand U7506 (N_7506,N_5041,N_4089);
nand U7507 (N_7507,N_4486,N_4520);
nor U7508 (N_7508,N_5499,N_5034);
nand U7509 (N_7509,N_5020,N_4950);
and U7510 (N_7510,N_5742,N_5077);
xnor U7511 (N_7511,N_5874,N_4212);
nor U7512 (N_7512,N_5168,N_5568);
nor U7513 (N_7513,N_4823,N_5533);
nand U7514 (N_7514,N_5625,N_5779);
nand U7515 (N_7515,N_5658,N_4384);
or U7516 (N_7516,N_5022,N_5458);
nand U7517 (N_7517,N_4881,N_4267);
or U7518 (N_7518,N_4980,N_5846);
xor U7519 (N_7519,N_5712,N_4908);
or U7520 (N_7520,N_5801,N_5660);
or U7521 (N_7521,N_4069,N_4072);
xor U7522 (N_7522,N_5669,N_5865);
or U7523 (N_7523,N_4824,N_5999);
or U7524 (N_7524,N_5754,N_4076);
xor U7525 (N_7525,N_5515,N_4170);
nand U7526 (N_7526,N_4948,N_5375);
nand U7527 (N_7527,N_4345,N_4294);
nor U7528 (N_7528,N_5081,N_5821);
or U7529 (N_7529,N_4324,N_5612);
xnor U7530 (N_7530,N_5425,N_4986);
nand U7531 (N_7531,N_4208,N_5052);
nor U7532 (N_7532,N_4659,N_5337);
nor U7533 (N_7533,N_5027,N_5516);
and U7534 (N_7534,N_5883,N_5154);
nand U7535 (N_7535,N_5075,N_5793);
or U7536 (N_7536,N_4187,N_5580);
or U7537 (N_7537,N_5679,N_4649);
or U7538 (N_7538,N_5235,N_5319);
or U7539 (N_7539,N_4134,N_5061);
and U7540 (N_7540,N_4368,N_5007);
and U7541 (N_7541,N_5134,N_5036);
or U7542 (N_7542,N_4948,N_5179);
xor U7543 (N_7543,N_4019,N_5490);
xor U7544 (N_7544,N_5959,N_4862);
xnor U7545 (N_7545,N_5774,N_4072);
or U7546 (N_7546,N_4660,N_4146);
nor U7547 (N_7547,N_5909,N_4312);
nor U7548 (N_7548,N_4962,N_5244);
or U7549 (N_7549,N_4413,N_5146);
or U7550 (N_7550,N_4386,N_5841);
and U7551 (N_7551,N_5504,N_4647);
or U7552 (N_7552,N_5828,N_4725);
nand U7553 (N_7553,N_4425,N_4581);
xor U7554 (N_7554,N_5196,N_4903);
nand U7555 (N_7555,N_4796,N_5082);
xor U7556 (N_7556,N_4621,N_4480);
xnor U7557 (N_7557,N_5115,N_4433);
or U7558 (N_7558,N_4384,N_5567);
or U7559 (N_7559,N_5679,N_5543);
and U7560 (N_7560,N_4423,N_5546);
xor U7561 (N_7561,N_4027,N_5477);
xnor U7562 (N_7562,N_5673,N_4027);
xnor U7563 (N_7563,N_4689,N_5420);
xor U7564 (N_7564,N_4676,N_4895);
nor U7565 (N_7565,N_4905,N_5504);
or U7566 (N_7566,N_4234,N_5054);
and U7567 (N_7567,N_5649,N_5342);
nand U7568 (N_7568,N_5291,N_4859);
nand U7569 (N_7569,N_5219,N_5679);
nand U7570 (N_7570,N_5907,N_4245);
or U7571 (N_7571,N_4526,N_5902);
and U7572 (N_7572,N_5750,N_5748);
and U7573 (N_7573,N_4175,N_4206);
or U7574 (N_7574,N_4950,N_4723);
and U7575 (N_7575,N_4590,N_5365);
nor U7576 (N_7576,N_5817,N_4745);
nor U7577 (N_7577,N_5693,N_5400);
xor U7578 (N_7578,N_4617,N_5950);
and U7579 (N_7579,N_5324,N_4941);
xnor U7580 (N_7580,N_5483,N_4499);
xor U7581 (N_7581,N_5951,N_5144);
or U7582 (N_7582,N_4987,N_4716);
or U7583 (N_7583,N_4816,N_4184);
xnor U7584 (N_7584,N_5442,N_4823);
nor U7585 (N_7585,N_5019,N_4379);
and U7586 (N_7586,N_5429,N_5820);
and U7587 (N_7587,N_4481,N_4279);
or U7588 (N_7588,N_5004,N_4816);
and U7589 (N_7589,N_4459,N_5528);
xnor U7590 (N_7590,N_5214,N_4746);
nand U7591 (N_7591,N_4903,N_4314);
nand U7592 (N_7592,N_4559,N_4738);
or U7593 (N_7593,N_5401,N_5152);
nand U7594 (N_7594,N_5880,N_4419);
nand U7595 (N_7595,N_5694,N_5857);
or U7596 (N_7596,N_4590,N_5009);
xnor U7597 (N_7597,N_5481,N_5809);
nand U7598 (N_7598,N_5693,N_4508);
and U7599 (N_7599,N_4350,N_4712);
nor U7600 (N_7600,N_4676,N_4043);
or U7601 (N_7601,N_5513,N_4254);
xor U7602 (N_7602,N_5055,N_5046);
or U7603 (N_7603,N_4753,N_4387);
xnor U7604 (N_7604,N_5107,N_4046);
nor U7605 (N_7605,N_5002,N_4375);
and U7606 (N_7606,N_5956,N_4679);
or U7607 (N_7607,N_4732,N_4769);
xnor U7608 (N_7608,N_4532,N_4726);
and U7609 (N_7609,N_4909,N_4530);
nor U7610 (N_7610,N_4158,N_4774);
nor U7611 (N_7611,N_5739,N_5535);
nor U7612 (N_7612,N_5790,N_4983);
or U7613 (N_7613,N_4386,N_4589);
xnor U7614 (N_7614,N_5520,N_4051);
or U7615 (N_7615,N_5035,N_5881);
and U7616 (N_7616,N_5380,N_5927);
nand U7617 (N_7617,N_5146,N_4561);
xor U7618 (N_7618,N_4891,N_4373);
or U7619 (N_7619,N_4441,N_4994);
xor U7620 (N_7620,N_4562,N_5468);
and U7621 (N_7621,N_4720,N_5559);
nand U7622 (N_7622,N_5630,N_5109);
and U7623 (N_7623,N_5114,N_4065);
nand U7624 (N_7624,N_4351,N_5003);
and U7625 (N_7625,N_4010,N_4385);
nor U7626 (N_7626,N_5639,N_4503);
nor U7627 (N_7627,N_5850,N_5177);
and U7628 (N_7628,N_4748,N_5870);
nand U7629 (N_7629,N_4259,N_4576);
or U7630 (N_7630,N_4834,N_4825);
nor U7631 (N_7631,N_5714,N_4062);
or U7632 (N_7632,N_4232,N_4786);
xor U7633 (N_7633,N_4315,N_4560);
xor U7634 (N_7634,N_4822,N_4030);
and U7635 (N_7635,N_4115,N_5709);
xnor U7636 (N_7636,N_5483,N_4504);
or U7637 (N_7637,N_4743,N_5852);
and U7638 (N_7638,N_5008,N_5883);
nor U7639 (N_7639,N_5423,N_5645);
and U7640 (N_7640,N_5672,N_4969);
xor U7641 (N_7641,N_5790,N_4007);
and U7642 (N_7642,N_4839,N_4276);
or U7643 (N_7643,N_5952,N_4751);
nor U7644 (N_7644,N_4708,N_4725);
or U7645 (N_7645,N_5018,N_5436);
xnor U7646 (N_7646,N_5449,N_5721);
or U7647 (N_7647,N_5714,N_4060);
or U7648 (N_7648,N_5207,N_5416);
xnor U7649 (N_7649,N_5853,N_5306);
and U7650 (N_7650,N_4942,N_4971);
nor U7651 (N_7651,N_4467,N_4632);
nand U7652 (N_7652,N_4720,N_5499);
nand U7653 (N_7653,N_5558,N_4720);
nand U7654 (N_7654,N_5576,N_5821);
nor U7655 (N_7655,N_5698,N_4933);
nand U7656 (N_7656,N_4780,N_5606);
nand U7657 (N_7657,N_4579,N_5231);
and U7658 (N_7658,N_4401,N_5021);
or U7659 (N_7659,N_4694,N_4942);
or U7660 (N_7660,N_4022,N_5185);
nor U7661 (N_7661,N_4863,N_5797);
nand U7662 (N_7662,N_5689,N_4242);
or U7663 (N_7663,N_4231,N_4357);
nor U7664 (N_7664,N_5640,N_5092);
nor U7665 (N_7665,N_5710,N_4474);
nor U7666 (N_7666,N_4995,N_4864);
xnor U7667 (N_7667,N_4703,N_4414);
xnor U7668 (N_7668,N_5535,N_4714);
xnor U7669 (N_7669,N_4065,N_5978);
xor U7670 (N_7670,N_4601,N_4616);
xor U7671 (N_7671,N_5481,N_4360);
nor U7672 (N_7672,N_4740,N_4232);
or U7673 (N_7673,N_5871,N_4350);
nand U7674 (N_7674,N_4234,N_4673);
or U7675 (N_7675,N_5498,N_4054);
xor U7676 (N_7676,N_5590,N_5058);
xnor U7677 (N_7677,N_4741,N_5347);
xnor U7678 (N_7678,N_5276,N_4686);
and U7679 (N_7679,N_4412,N_4928);
nand U7680 (N_7680,N_5391,N_4576);
nand U7681 (N_7681,N_4122,N_5139);
nor U7682 (N_7682,N_4261,N_4220);
nor U7683 (N_7683,N_5470,N_4542);
and U7684 (N_7684,N_5214,N_5761);
or U7685 (N_7685,N_5602,N_5073);
or U7686 (N_7686,N_5707,N_5667);
or U7687 (N_7687,N_5938,N_5952);
or U7688 (N_7688,N_5435,N_4988);
nor U7689 (N_7689,N_5451,N_5329);
and U7690 (N_7690,N_4023,N_4072);
xor U7691 (N_7691,N_5800,N_4664);
nand U7692 (N_7692,N_5317,N_4385);
nand U7693 (N_7693,N_4066,N_5792);
xnor U7694 (N_7694,N_5035,N_5106);
and U7695 (N_7695,N_4421,N_4919);
and U7696 (N_7696,N_5031,N_4596);
nand U7697 (N_7697,N_5550,N_5736);
nand U7698 (N_7698,N_4529,N_5870);
xor U7699 (N_7699,N_5635,N_4350);
and U7700 (N_7700,N_4406,N_4651);
nand U7701 (N_7701,N_5931,N_5605);
nor U7702 (N_7702,N_4713,N_4959);
xnor U7703 (N_7703,N_5094,N_4940);
xor U7704 (N_7704,N_5417,N_5332);
nand U7705 (N_7705,N_5140,N_4978);
xor U7706 (N_7706,N_5705,N_5389);
nor U7707 (N_7707,N_5613,N_4982);
and U7708 (N_7708,N_5342,N_5966);
nor U7709 (N_7709,N_5687,N_4948);
or U7710 (N_7710,N_4264,N_5796);
nand U7711 (N_7711,N_4435,N_4965);
nor U7712 (N_7712,N_5166,N_5992);
nor U7713 (N_7713,N_5074,N_4757);
nor U7714 (N_7714,N_4866,N_5340);
or U7715 (N_7715,N_4186,N_5363);
xor U7716 (N_7716,N_4691,N_5212);
and U7717 (N_7717,N_5855,N_5858);
xnor U7718 (N_7718,N_5654,N_4097);
xnor U7719 (N_7719,N_4362,N_4099);
and U7720 (N_7720,N_4576,N_4973);
nand U7721 (N_7721,N_4022,N_5202);
or U7722 (N_7722,N_4856,N_4954);
and U7723 (N_7723,N_4485,N_4188);
or U7724 (N_7724,N_5157,N_4560);
nand U7725 (N_7725,N_4656,N_4814);
nand U7726 (N_7726,N_4658,N_5562);
nand U7727 (N_7727,N_5122,N_5857);
nand U7728 (N_7728,N_4758,N_4577);
nor U7729 (N_7729,N_4443,N_4532);
nor U7730 (N_7730,N_4968,N_4567);
nor U7731 (N_7731,N_4893,N_5268);
and U7732 (N_7732,N_5228,N_4298);
nand U7733 (N_7733,N_4304,N_5773);
nand U7734 (N_7734,N_4239,N_5290);
nor U7735 (N_7735,N_5864,N_5554);
or U7736 (N_7736,N_4296,N_4721);
and U7737 (N_7737,N_5827,N_5510);
or U7738 (N_7738,N_5886,N_5706);
xnor U7739 (N_7739,N_5285,N_4894);
nor U7740 (N_7740,N_5332,N_4397);
xnor U7741 (N_7741,N_5619,N_4094);
and U7742 (N_7742,N_4302,N_4523);
nand U7743 (N_7743,N_5554,N_5856);
or U7744 (N_7744,N_4060,N_5640);
xnor U7745 (N_7745,N_4381,N_4734);
or U7746 (N_7746,N_5576,N_5152);
or U7747 (N_7747,N_5670,N_5675);
nor U7748 (N_7748,N_5366,N_5002);
and U7749 (N_7749,N_5802,N_5948);
or U7750 (N_7750,N_5398,N_4873);
and U7751 (N_7751,N_5954,N_4548);
nand U7752 (N_7752,N_4981,N_4312);
nand U7753 (N_7753,N_4926,N_4765);
xnor U7754 (N_7754,N_4351,N_4750);
and U7755 (N_7755,N_4789,N_5672);
nand U7756 (N_7756,N_5108,N_4944);
or U7757 (N_7757,N_4885,N_5829);
nor U7758 (N_7758,N_5012,N_5935);
xnor U7759 (N_7759,N_4604,N_5916);
xnor U7760 (N_7760,N_4524,N_4684);
xnor U7761 (N_7761,N_4120,N_4597);
and U7762 (N_7762,N_5427,N_5966);
or U7763 (N_7763,N_5259,N_4539);
or U7764 (N_7764,N_4226,N_5897);
nor U7765 (N_7765,N_4412,N_4775);
xor U7766 (N_7766,N_5586,N_4344);
or U7767 (N_7767,N_5276,N_4877);
nor U7768 (N_7768,N_5155,N_5305);
xnor U7769 (N_7769,N_4377,N_5863);
nor U7770 (N_7770,N_5422,N_5791);
xor U7771 (N_7771,N_5750,N_4610);
or U7772 (N_7772,N_5958,N_4577);
nor U7773 (N_7773,N_4581,N_4716);
nand U7774 (N_7774,N_5487,N_5603);
nor U7775 (N_7775,N_4539,N_5590);
and U7776 (N_7776,N_5859,N_4848);
nor U7777 (N_7777,N_4132,N_4871);
or U7778 (N_7778,N_5294,N_5562);
or U7779 (N_7779,N_4387,N_5600);
and U7780 (N_7780,N_4263,N_5593);
nand U7781 (N_7781,N_5741,N_4247);
xnor U7782 (N_7782,N_5739,N_5042);
xnor U7783 (N_7783,N_4215,N_5768);
nor U7784 (N_7784,N_4974,N_4689);
and U7785 (N_7785,N_4785,N_5298);
xor U7786 (N_7786,N_4258,N_5513);
nor U7787 (N_7787,N_5533,N_5879);
nand U7788 (N_7788,N_4837,N_4899);
nand U7789 (N_7789,N_5188,N_4285);
nor U7790 (N_7790,N_5551,N_4319);
nand U7791 (N_7791,N_4147,N_5171);
nor U7792 (N_7792,N_4717,N_5202);
and U7793 (N_7793,N_4008,N_4046);
nor U7794 (N_7794,N_4380,N_5582);
nor U7795 (N_7795,N_5258,N_4548);
nand U7796 (N_7796,N_5813,N_5772);
xor U7797 (N_7797,N_4232,N_4040);
or U7798 (N_7798,N_4512,N_5365);
xnor U7799 (N_7799,N_4784,N_4408);
nor U7800 (N_7800,N_5890,N_4675);
xor U7801 (N_7801,N_5588,N_4942);
or U7802 (N_7802,N_4443,N_4979);
xnor U7803 (N_7803,N_5563,N_5545);
nand U7804 (N_7804,N_4474,N_4681);
or U7805 (N_7805,N_5362,N_5939);
nand U7806 (N_7806,N_5764,N_5121);
or U7807 (N_7807,N_5887,N_5561);
and U7808 (N_7808,N_5184,N_5710);
nand U7809 (N_7809,N_5744,N_4497);
nand U7810 (N_7810,N_5006,N_4182);
xnor U7811 (N_7811,N_4702,N_4203);
or U7812 (N_7812,N_5972,N_4362);
nor U7813 (N_7813,N_4305,N_5892);
nor U7814 (N_7814,N_4325,N_4402);
nand U7815 (N_7815,N_5228,N_4041);
nor U7816 (N_7816,N_4137,N_4138);
nor U7817 (N_7817,N_5322,N_4492);
nor U7818 (N_7818,N_5078,N_5918);
xnor U7819 (N_7819,N_4823,N_5890);
and U7820 (N_7820,N_4411,N_4296);
or U7821 (N_7821,N_5546,N_5184);
nand U7822 (N_7822,N_4294,N_5792);
nand U7823 (N_7823,N_5194,N_4000);
and U7824 (N_7824,N_5521,N_4000);
and U7825 (N_7825,N_5471,N_5804);
nor U7826 (N_7826,N_4570,N_5368);
and U7827 (N_7827,N_4692,N_4171);
nand U7828 (N_7828,N_5600,N_5114);
or U7829 (N_7829,N_4763,N_5323);
and U7830 (N_7830,N_4450,N_5900);
and U7831 (N_7831,N_5526,N_5001);
and U7832 (N_7832,N_4091,N_4980);
and U7833 (N_7833,N_4622,N_5184);
or U7834 (N_7834,N_4189,N_4375);
nor U7835 (N_7835,N_5250,N_4258);
nand U7836 (N_7836,N_4656,N_4030);
or U7837 (N_7837,N_4773,N_5375);
and U7838 (N_7838,N_4826,N_5733);
nand U7839 (N_7839,N_5998,N_4547);
nand U7840 (N_7840,N_5887,N_4484);
xnor U7841 (N_7841,N_4147,N_5655);
nand U7842 (N_7842,N_5124,N_5126);
and U7843 (N_7843,N_4702,N_4755);
nand U7844 (N_7844,N_5733,N_5064);
or U7845 (N_7845,N_5310,N_5847);
nand U7846 (N_7846,N_4949,N_4315);
or U7847 (N_7847,N_4279,N_5281);
and U7848 (N_7848,N_4134,N_4453);
and U7849 (N_7849,N_5986,N_4734);
and U7850 (N_7850,N_5759,N_5565);
nor U7851 (N_7851,N_5123,N_4185);
nor U7852 (N_7852,N_5989,N_5856);
xor U7853 (N_7853,N_4089,N_4001);
nand U7854 (N_7854,N_4393,N_5173);
xor U7855 (N_7855,N_4313,N_4758);
nand U7856 (N_7856,N_4646,N_5627);
xnor U7857 (N_7857,N_4756,N_4682);
and U7858 (N_7858,N_4932,N_4891);
nor U7859 (N_7859,N_5389,N_5847);
and U7860 (N_7860,N_5537,N_4870);
or U7861 (N_7861,N_5465,N_5536);
or U7862 (N_7862,N_5983,N_4070);
xor U7863 (N_7863,N_5670,N_4245);
nor U7864 (N_7864,N_4989,N_5957);
xor U7865 (N_7865,N_5990,N_4930);
nor U7866 (N_7866,N_4389,N_4948);
or U7867 (N_7867,N_4434,N_5648);
xnor U7868 (N_7868,N_5132,N_4364);
and U7869 (N_7869,N_5530,N_4301);
and U7870 (N_7870,N_5165,N_4372);
nor U7871 (N_7871,N_5752,N_4638);
xnor U7872 (N_7872,N_5647,N_4551);
nor U7873 (N_7873,N_4791,N_4022);
nor U7874 (N_7874,N_5995,N_4042);
and U7875 (N_7875,N_4125,N_4207);
nor U7876 (N_7876,N_4474,N_4933);
nand U7877 (N_7877,N_4811,N_4866);
and U7878 (N_7878,N_5740,N_5090);
nor U7879 (N_7879,N_5404,N_4228);
xor U7880 (N_7880,N_4105,N_4590);
xnor U7881 (N_7881,N_5443,N_5623);
nand U7882 (N_7882,N_5480,N_4236);
xor U7883 (N_7883,N_5544,N_4126);
nor U7884 (N_7884,N_4435,N_4371);
nor U7885 (N_7885,N_5963,N_5100);
and U7886 (N_7886,N_4303,N_4924);
and U7887 (N_7887,N_5282,N_4935);
and U7888 (N_7888,N_5943,N_5432);
or U7889 (N_7889,N_4338,N_4041);
nand U7890 (N_7890,N_5770,N_5790);
nor U7891 (N_7891,N_5238,N_5182);
nand U7892 (N_7892,N_5124,N_5633);
nor U7893 (N_7893,N_5685,N_4701);
or U7894 (N_7894,N_5737,N_5289);
and U7895 (N_7895,N_5740,N_5898);
or U7896 (N_7896,N_4362,N_5791);
or U7897 (N_7897,N_4833,N_5028);
or U7898 (N_7898,N_4149,N_5065);
xor U7899 (N_7899,N_4732,N_4807);
xor U7900 (N_7900,N_4403,N_4194);
or U7901 (N_7901,N_5940,N_5648);
or U7902 (N_7902,N_4439,N_5334);
xor U7903 (N_7903,N_5466,N_5878);
nor U7904 (N_7904,N_4499,N_4491);
xor U7905 (N_7905,N_4102,N_5863);
xnor U7906 (N_7906,N_5351,N_4525);
xnor U7907 (N_7907,N_4171,N_4859);
or U7908 (N_7908,N_4135,N_4663);
xor U7909 (N_7909,N_4738,N_4182);
or U7910 (N_7910,N_5174,N_4330);
xor U7911 (N_7911,N_5207,N_4469);
or U7912 (N_7912,N_5771,N_5704);
xor U7913 (N_7913,N_4790,N_5876);
or U7914 (N_7914,N_4329,N_5962);
and U7915 (N_7915,N_4387,N_4615);
and U7916 (N_7916,N_4362,N_4008);
xnor U7917 (N_7917,N_5159,N_4299);
nand U7918 (N_7918,N_4170,N_4702);
nor U7919 (N_7919,N_5042,N_5552);
nand U7920 (N_7920,N_4830,N_5438);
nor U7921 (N_7921,N_5856,N_5006);
xor U7922 (N_7922,N_4149,N_5555);
xor U7923 (N_7923,N_5438,N_4393);
and U7924 (N_7924,N_4599,N_4603);
and U7925 (N_7925,N_4968,N_5354);
or U7926 (N_7926,N_4210,N_4344);
or U7927 (N_7927,N_4085,N_4596);
and U7928 (N_7928,N_4343,N_4263);
nand U7929 (N_7929,N_5549,N_4017);
nor U7930 (N_7930,N_5063,N_4861);
or U7931 (N_7931,N_4926,N_4899);
xor U7932 (N_7932,N_4218,N_4048);
or U7933 (N_7933,N_4217,N_4673);
and U7934 (N_7934,N_5175,N_4251);
nand U7935 (N_7935,N_4635,N_4541);
and U7936 (N_7936,N_5255,N_4618);
and U7937 (N_7937,N_4712,N_4417);
and U7938 (N_7938,N_5135,N_4048);
nand U7939 (N_7939,N_5916,N_5851);
or U7940 (N_7940,N_5479,N_5481);
nand U7941 (N_7941,N_4249,N_4513);
or U7942 (N_7942,N_4221,N_4940);
nor U7943 (N_7943,N_5440,N_4419);
or U7944 (N_7944,N_4864,N_5497);
and U7945 (N_7945,N_4027,N_4052);
nand U7946 (N_7946,N_5620,N_5568);
or U7947 (N_7947,N_4727,N_5324);
xnor U7948 (N_7948,N_5053,N_4757);
or U7949 (N_7949,N_5078,N_5735);
and U7950 (N_7950,N_4510,N_4854);
and U7951 (N_7951,N_4355,N_4446);
and U7952 (N_7952,N_5753,N_5527);
xor U7953 (N_7953,N_4265,N_5396);
and U7954 (N_7954,N_4844,N_4727);
xnor U7955 (N_7955,N_4729,N_4983);
and U7956 (N_7956,N_5959,N_5004);
xor U7957 (N_7957,N_4285,N_5443);
and U7958 (N_7958,N_5293,N_5156);
nand U7959 (N_7959,N_5989,N_4642);
xnor U7960 (N_7960,N_4002,N_4973);
or U7961 (N_7961,N_4247,N_5118);
or U7962 (N_7962,N_5124,N_4420);
nand U7963 (N_7963,N_5492,N_5163);
nor U7964 (N_7964,N_5041,N_5936);
nor U7965 (N_7965,N_5173,N_4622);
and U7966 (N_7966,N_4300,N_5204);
or U7967 (N_7967,N_5271,N_4034);
nor U7968 (N_7968,N_4324,N_4837);
and U7969 (N_7969,N_4929,N_5952);
or U7970 (N_7970,N_4499,N_5793);
xor U7971 (N_7971,N_4111,N_5526);
nand U7972 (N_7972,N_4431,N_4705);
xnor U7973 (N_7973,N_5613,N_5532);
xnor U7974 (N_7974,N_5989,N_4629);
or U7975 (N_7975,N_5266,N_4188);
and U7976 (N_7976,N_5060,N_5040);
nand U7977 (N_7977,N_4244,N_4905);
nand U7978 (N_7978,N_4056,N_4184);
nand U7979 (N_7979,N_4614,N_5514);
xnor U7980 (N_7980,N_5229,N_4821);
nor U7981 (N_7981,N_5932,N_4085);
xnor U7982 (N_7982,N_5845,N_4582);
nand U7983 (N_7983,N_5461,N_5652);
nor U7984 (N_7984,N_4713,N_5989);
and U7985 (N_7985,N_4542,N_5531);
xnor U7986 (N_7986,N_5864,N_4568);
and U7987 (N_7987,N_5446,N_5944);
xnor U7988 (N_7988,N_4304,N_4853);
xnor U7989 (N_7989,N_5113,N_5576);
and U7990 (N_7990,N_4307,N_5087);
nor U7991 (N_7991,N_5025,N_4390);
xnor U7992 (N_7992,N_4998,N_4770);
xnor U7993 (N_7993,N_4861,N_5255);
and U7994 (N_7994,N_5897,N_4683);
xor U7995 (N_7995,N_5629,N_5099);
xor U7996 (N_7996,N_4878,N_5111);
nor U7997 (N_7997,N_5785,N_4389);
nand U7998 (N_7998,N_5943,N_5190);
nor U7999 (N_7999,N_5851,N_4209);
nor U8000 (N_8000,N_7295,N_7775);
or U8001 (N_8001,N_6930,N_6914);
and U8002 (N_8002,N_6271,N_7038);
nor U8003 (N_8003,N_7140,N_7312);
and U8004 (N_8004,N_6612,N_7734);
xor U8005 (N_8005,N_7618,N_7784);
nor U8006 (N_8006,N_6607,N_6753);
nor U8007 (N_8007,N_7078,N_6875);
nand U8008 (N_8008,N_7264,N_6281);
xor U8009 (N_8009,N_6379,N_6794);
nor U8010 (N_8010,N_7957,N_6334);
or U8011 (N_8011,N_6261,N_6879);
xnor U8012 (N_8012,N_7835,N_7811);
nor U8013 (N_8013,N_6815,N_7715);
or U8014 (N_8014,N_7699,N_6047);
nor U8015 (N_8015,N_6965,N_7073);
and U8016 (N_8016,N_7768,N_7194);
xor U8017 (N_8017,N_7976,N_7416);
xor U8018 (N_8018,N_7979,N_6501);
and U8019 (N_8019,N_7540,N_6128);
nor U8020 (N_8020,N_7920,N_6820);
nor U8021 (N_8021,N_6773,N_6731);
nand U8022 (N_8022,N_7372,N_7656);
xor U8023 (N_8023,N_7158,N_6113);
nand U8024 (N_8024,N_7070,N_7946);
xor U8025 (N_8025,N_6217,N_7686);
nor U8026 (N_8026,N_6955,N_7532);
xnor U8027 (N_8027,N_7858,N_7412);
or U8028 (N_8028,N_6092,N_6841);
or U8029 (N_8029,N_7752,N_6371);
nand U8030 (N_8030,N_7017,N_7812);
and U8031 (N_8031,N_7989,N_6249);
and U8032 (N_8032,N_6412,N_6748);
nand U8033 (N_8033,N_7243,N_7588);
nor U8034 (N_8034,N_6505,N_6272);
and U8035 (N_8035,N_6929,N_6206);
xnor U8036 (N_8036,N_7509,N_6585);
or U8037 (N_8037,N_6399,N_6054);
xnor U8038 (N_8038,N_7436,N_6978);
or U8039 (N_8039,N_6862,N_7596);
and U8040 (N_8040,N_7885,N_6961);
xnor U8041 (N_8041,N_6020,N_6735);
nand U8042 (N_8042,N_6609,N_7611);
nand U8043 (N_8043,N_7725,N_7007);
nand U8044 (N_8044,N_7395,N_6489);
or U8045 (N_8045,N_7987,N_7429);
or U8046 (N_8046,N_7467,N_6458);
or U8047 (N_8047,N_6297,N_6403);
xor U8048 (N_8048,N_6004,N_6477);
and U8049 (N_8049,N_6022,N_6284);
nor U8050 (N_8050,N_6590,N_6050);
and U8051 (N_8051,N_7761,N_6362);
xor U8052 (N_8052,N_7263,N_7622);
xnor U8053 (N_8053,N_6378,N_7266);
and U8054 (N_8054,N_6828,N_7777);
or U8055 (N_8055,N_7727,N_7164);
and U8056 (N_8056,N_7616,N_6035);
nand U8057 (N_8057,N_7703,N_7117);
and U8058 (N_8058,N_7672,N_6739);
and U8059 (N_8059,N_6594,N_6716);
or U8060 (N_8060,N_7292,N_7655);
xnor U8061 (N_8061,N_6204,N_6051);
nor U8062 (N_8062,N_6418,N_7685);
xor U8063 (N_8063,N_6960,N_6222);
xnor U8064 (N_8064,N_7548,N_7359);
xnor U8065 (N_8065,N_6627,N_7380);
nor U8066 (N_8066,N_7493,N_7492);
or U8067 (N_8067,N_6698,N_6394);
nor U8068 (N_8068,N_6372,N_7900);
or U8069 (N_8069,N_6808,N_6993);
nor U8070 (N_8070,N_6294,N_7658);
nor U8071 (N_8071,N_7317,N_6279);
nand U8072 (N_8072,N_7254,N_6523);
nand U8073 (N_8073,N_6009,N_7889);
nand U8074 (N_8074,N_7912,N_6405);
or U8075 (N_8075,N_6954,N_6974);
nor U8076 (N_8076,N_7260,N_6743);
nor U8077 (N_8077,N_6924,N_7082);
nand U8078 (N_8078,N_6327,N_7785);
nand U8079 (N_8079,N_6416,N_6262);
nand U8080 (N_8080,N_7817,N_6580);
nand U8081 (N_8081,N_6330,N_7119);
and U8082 (N_8082,N_7246,N_7178);
or U8083 (N_8083,N_7661,N_6397);
nand U8084 (N_8084,N_7864,N_7267);
and U8085 (N_8085,N_6560,N_7402);
and U8086 (N_8086,N_7696,N_7886);
or U8087 (N_8087,N_6830,N_7333);
nand U8088 (N_8088,N_7102,N_7430);
and U8089 (N_8089,N_6124,N_6832);
nand U8090 (N_8090,N_7407,N_6303);
or U8091 (N_8091,N_7508,N_7182);
and U8092 (N_8092,N_6650,N_7591);
xnor U8093 (N_8093,N_6717,N_7199);
nand U8094 (N_8094,N_7604,N_6805);
nand U8095 (N_8095,N_6931,N_6301);
or U8096 (N_8096,N_6525,N_6463);
nor U8097 (N_8097,N_7172,N_6094);
and U8098 (N_8098,N_6663,N_6583);
nand U8099 (N_8099,N_7838,N_6352);
nand U8100 (N_8100,N_7155,N_6364);
xor U8101 (N_8101,N_7062,N_7859);
xnor U8102 (N_8102,N_7855,N_6472);
nand U8103 (N_8103,N_7648,N_6771);
nand U8104 (N_8104,N_6316,N_7643);
and U8105 (N_8105,N_7918,N_6256);
xnor U8106 (N_8106,N_6162,N_7203);
nand U8107 (N_8107,N_6881,N_7634);
nand U8108 (N_8108,N_7684,N_6264);
xor U8109 (N_8109,N_7177,N_7413);
nor U8110 (N_8110,N_7081,N_6592);
nand U8111 (N_8111,N_6713,N_6780);
xor U8112 (N_8112,N_6269,N_7211);
nor U8113 (N_8113,N_7603,N_6604);
or U8114 (N_8114,N_6447,N_6427);
or U8115 (N_8115,N_7726,N_7871);
nand U8116 (N_8116,N_6431,N_6992);
and U8117 (N_8117,N_7356,N_6428);
nor U8118 (N_8118,N_7210,N_7428);
or U8119 (N_8119,N_7681,N_6564);
or U8120 (N_8120,N_7570,N_6761);
or U8121 (N_8121,N_6185,N_7612);
nand U8122 (N_8122,N_6918,N_7000);
nor U8123 (N_8123,N_7068,N_7579);
nand U8124 (N_8124,N_7016,N_7818);
nand U8125 (N_8125,N_6647,N_7472);
and U8126 (N_8126,N_7418,N_6161);
or U8127 (N_8127,N_6956,N_6917);
xor U8128 (N_8128,N_7444,N_7130);
nor U8129 (N_8129,N_7345,N_7251);
nor U8130 (N_8130,N_7795,N_6097);
nor U8131 (N_8131,N_7772,N_6706);
nor U8132 (N_8132,N_7015,N_6865);
nand U8133 (N_8133,N_7111,N_6621);
xnor U8134 (N_8134,N_7526,N_6677);
nand U8135 (N_8135,N_6312,N_6021);
xnor U8136 (N_8136,N_6145,N_7950);
nor U8137 (N_8137,N_7244,N_7660);
xnor U8138 (N_8138,N_7866,N_7257);
or U8139 (N_8139,N_6933,N_7948);
or U8140 (N_8140,N_6522,N_6894);
xor U8141 (N_8141,N_6365,N_7283);
nor U8142 (N_8142,N_6725,N_6878);
xnor U8143 (N_8143,N_6738,N_7956);
or U8144 (N_8144,N_6632,N_7298);
nand U8145 (N_8145,N_7272,N_7735);
xor U8146 (N_8146,N_7732,N_6423);
nand U8147 (N_8147,N_6223,N_7714);
or U8148 (N_8148,N_6969,N_6198);
or U8149 (N_8149,N_7488,N_6386);
nand U8150 (N_8150,N_6120,N_7473);
and U8151 (N_8151,N_7872,N_7138);
and U8152 (N_8152,N_6366,N_7455);
xor U8153 (N_8153,N_7037,N_6192);
and U8154 (N_8154,N_7797,N_6913);
nor U8155 (N_8155,N_7437,N_6532);
xor U8156 (N_8156,N_6376,N_6186);
xor U8157 (N_8157,N_6977,N_6860);
and U8158 (N_8158,N_7939,N_6578);
nor U8159 (N_8159,N_6190,N_7443);
xnor U8160 (N_8160,N_7340,N_6970);
nand U8161 (N_8161,N_6215,N_6488);
nand U8162 (N_8162,N_7644,N_6575);
and U8163 (N_8163,N_7439,N_7120);
xnor U8164 (N_8164,N_6963,N_6259);
and U8165 (N_8165,N_7708,N_7367);
nor U8166 (N_8166,N_7165,N_6498);
nand U8167 (N_8167,N_7227,N_7891);
xor U8168 (N_8168,N_6160,N_7927);
and U8169 (N_8169,N_7301,N_7999);
xnor U8170 (N_8170,N_7516,N_6343);
nand U8171 (N_8171,N_6644,N_7438);
nand U8172 (N_8172,N_6859,N_7212);
and U8173 (N_8173,N_6346,N_7464);
xnor U8174 (N_8174,N_6559,N_6539);
nand U8175 (N_8175,N_7013,N_7743);
or U8176 (N_8176,N_6165,N_7763);
xor U8177 (N_8177,N_6871,N_7836);
nor U8178 (N_8178,N_6642,N_6547);
nor U8179 (N_8179,N_7142,N_6686);
xnor U8180 (N_8180,N_7792,N_7309);
or U8181 (N_8181,N_7503,N_6587);
or U8182 (N_8182,N_6452,N_7929);
nor U8183 (N_8183,N_6229,N_7450);
nor U8184 (N_8184,N_6546,N_7654);
and U8185 (N_8185,N_7105,N_7274);
and U8186 (N_8186,N_6385,N_7711);
and U8187 (N_8187,N_7518,N_7973);
nand U8188 (N_8188,N_6854,N_7635);
xor U8189 (N_8189,N_7722,N_6473);
and U8190 (N_8190,N_6673,N_6430);
nor U8191 (N_8191,N_6197,N_6283);
xor U8192 (N_8192,N_6703,N_6638);
and U8193 (N_8193,N_7103,N_7747);
nor U8194 (N_8194,N_6895,N_7801);
nand U8195 (N_8195,N_7175,N_7159);
nand U8196 (N_8196,N_7149,N_7665);
or U8197 (N_8197,N_6628,N_7033);
or U8198 (N_8198,N_7147,N_7562);
nor U8199 (N_8199,N_6252,N_7977);
and U8200 (N_8200,N_7196,N_7083);
xnor U8201 (N_8201,N_7883,N_7851);
nor U8202 (N_8202,N_7168,N_6781);
and U8203 (N_8203,N_7750,N_6251);
nand U8204 (N_8204,N_6694,N_7406);
nand U8205 (N_8205,N_6643,N_6635);
xor U8206 (N_8206,N_7632,N_7335);
nor U8207 (N_8207,N_6085,N_6200);
or U8208 (N_8208,N_7066,N_6305);
nand U8209 (N_8209,N_7288,N_7151);
nand U8210 (N_8210,N_7781,N_6278);
xnor U8211 (N_8211,N_6136,N_7405);
xor U8212 (N_8212,N_7305,N_7967);
and U8213 (N_8213,N_6763,N_6103);
xor U8214 (N_8214,N_6112,N_6356);
and U8215 (N_8215,N_6337,N_6614);
nand U8216 (N_8216,N_6221,N_7993);
and U8217 (N_8217,N_6067,N_6119);
nor U8218 (N_8218,N_6086,N_7605);
nor U8219 (N_8219,N_7679,N_7360);
or U8220 (N_8220,N_7981,N_6013);
xor U8221 (N_8221,N_7024,N_6757);
or U8222 (N_8222,N_6806,N_7375);
nand U8223 (N_8223,N_6220,N_6766);
nor U8224 (N_8224,N_6089,N_6076);
or U8225 (N_8225,N_7381,N_7765);
nor U8226 (N_8226,N_7379,N_7982);
and U8227 (N_8227,N_7983,N_7124);
or U8228 (N_8228,N_7678,N_6581);
nor U8229 (N_8229,N_7718,N_6833);
nor U8230 (N_8230,N_6711,N_6979);
and U8231 (N_8231,N_7343,N_6801);
xnor U8232 (N_8232,N_7421,N_7086);
and U8233 (N_8233,N_7442,N_6110);
nand U8234 (N_8234,N_7700,N_7101);
nand U8235 (N_8235,N_7624,N_7563);
nand U8236 (N_8236,N_7557,N_6006);
nand U8237 (N_8237,N_7136,N_7809);
xnor U8238 (N_8238,N_6118,N_7284);
xor U8239 (N_8239,N_7206,N_6319);
nor U8240 (N_8240,N_7922,N_6056);
nand U8241 (N_8241,N_6670,N_6809);
xor U8242 (N_8242,N_6353,N_7840);
and U8243 (N_8243,N_6872,N_6922);
xor U8244 (N_8244,N_7424,N_6617);
nand U8245 (N_8245,N_6495,N_6726);
nand U8246 (N_8246,N_7352,N_7121);
xor U8247 (N_8247,N_6328,N_6823);
nor U8248 (N_8248,N_6422,N_6709);
xnor U8249 (N_8249,N_7691,N_6077);
xnor U8250 (N_8250,N_7319,N_7690);
nor U8251 (N_8251,N_6890,N_6361);
xor U8252 (N_8252,N_6905,N_7456);
or U8253 (N_8253,N_6537,N_6135);
and U8254 (N_8254,N_7067,N_7749);
or U8255 (N_8255,N_7890,N_6882);
xnor U8256 (N_8256,N_6964,N_6506);
xnor U8257 (N_8257,N_6762,N_6692);
nor U8258 (N_8258,N_7803,N_6286);
nand U8259 (N_8259,N_7565,N_6032);
and U8260 (N_8260,N_6363,N_7815);
nor U8261 (N_8261,N_7549,N_7020);
nor U8262 (N_8262,N_6904,N_6459);
nand U8263 (N_8263,N_6512,N_7054);
nand U8264 (N_8264,N_6742,N_7773);
or U8265 (N_8265,N_7645,N_7482);
and U8266 (N_8266,N_6658,N_6445);
or U8267 (N_8267,N_6849,N_6653);
xor U8268 (N_8268,N_6582,N_6008);
nor U8269 (N_8269,N_7693,N_6891);
nand U8270 (N_8270,N_7550,N_6513);
nand U8271 (N_8271,N_7213,N_7529);
or U8272 (N_8272,N_6595,N_7821);
or U8273 (N_8273,N_7329,N_6042);
xnor U8274 (N_8274,N_6333,N_6061);
nor U8275 (N_8275,N_6025,N_7807);
or U8276 (N_8276,N_7435,N_6856);
xor U8277 (N_8277,N_7357,N_7106);
xnor U8278 (N_8278,N_7831,N_7148);
xor U8279 (N_8279,N_7805,N_6325);
nand U8280 (N_8280,N_7875,N_7580);
xor U8281 (N_8281,N_6840,N_6851);
xor U8282 (N_8282,N_7525,N_7241);
xnor U8283 (N_8283,N_7842,N_6778);
and U8284 (N_8284,N_6637,N_7465);
nor U8285 (N_8285,N_7386,N_7731);
nand U8286 (N_8286,N_7631,N_7475);
and U8287 (N_8287,N_6615,N_7287);
nor U8288 (N_8288,N_6344,N_7951);
xnor U8289 (N_8289,N_7426,N_7417);
or U8290 (N_8290,N_7001,N_6681);
nand U8291 (N_8291,N_7867,N_6749);
nand U8292 (N_8292,N_6065,N_7209);
and U8293 (N_8293,N_6844,N_6669);
nor U8294 (N_8294,N_7262,N_6434);
xnor U8295 (N_8295,N_7471,N_6402);
nand U8296 (N_8296,N_7991,N_6026);
and U8297 (N_8297,N_6313,N_6737);
nor U8298 (N_8298,N_6940,N_6184);
xnor U8299 (N_8299,N_6419,N_6123);
nor U8300 (N_8300,N_7469,N_7245);
nor U8301 (N_8301,N_6375,N_7739);
and U8302 (N_8302,N_6521,N_7796);
nand U8303 (N_8303,N_7500,N_7152);
or U8304 (N_8304,N_7928,N_7915);
nor U8305 (N_8305,N_7810,N_6784);
and U8306 (N_8306,N_6242,N_6923);
xor U8307 (N_8307,N_6908,N_6996);
and U8308 (N_8308,N_7445,N_7729);
or U8309 (N_8309,N_7145,N_7895);
xor U8310 (N_8310,N_6699,N_6540);
nand U8311 (N_8311,N_6591,N_6927);
nor U8312 (N_8312,N_7330,N_7404);
nor U8313 (N_8313,N_6100,N_7326);
nand U8314 (N_8314,N_6314,N_7935);
nor U8315 (N_8315,N_7528,N_7804);
nor U8316 (N_8316,N_7598,N_6370);
nand U8317 (N_8317,N_6132,N_6465);
xor U8318 (N_8318,N_6819,N_7293);
or U8319 (N_8319,N_6600,N_6724);
xor U8320 (N_8320,N_7334,N_7794);
xnor U8321 (N_8321,N_6187,N_6906);
or U8322 (N_8322,N_6182,N_6705);
and U8323 (N_8323,N_6530,N_6439);
nor U8324 (N_8324,N_6255,N_6341);
or U8325 (N_8325,N_6526,N_6656);
xor U8326 (N_8326,N_6475,N_7051);
nand U8327 (N_8327,N_7962,N_7219);
or U8328 (N_8328,N_6693,N_7128);
nor U8329 (N_8329,N_7601,N_6049);
xor U8330 (N_8330,N_6792,N_6818);
or U8331 (N_8331,N_7474,N_6528);
nor U8332 (N_8332,N_7167,N_7931);
nor U8333 (N_8333,N_7852,N_7834);
nand U8334 (N_8334,N_6733,N_7131);
and U8335 (N_8335,N_6210,N_6280);
or U8336 (N_8336,N_7370,N_6115);
nand U8337 (N_8337,N_7391,N_6561);
and U8338 (N_8338,N_6935,N_6510);
or U8339 (N_8339,N_7127,N_6962);
nor U8340 (N_8340,N_7207,N_6276);
nand U8341 (N_8341,N_6406,N_6177);
and U8342 (N_8342,N_6641,N_6446);
and U8343 (N_8343,N_6899,N_7388);
xor U8344 (N_8344,N_6415,N_7936);
xor U8345 (N_8345,N_6852,N_6414);
nor U8346 (N_8346,N_7639,N_7778);
and U8347 (N_8347,N_6461,N_6413);
and U8348 (N_8348,N_7487,N_6554);
or U8349 (N_8349,N_7228,N_7239);
nand U8350 (N_8350,N_7599,N_7745);
nor U8351 (N_8351,N_6787,N_7191);
or U8352 (N_8352,N_6630,N_6104);
or U8353 (N_8353,N_7857,N_6777);
xor U8354 (N_8354,N_6588,N_6986);
xor U8355 (N_8355,N_7517,N_6323);
xor U8356 (N_8356,N_6816,N_7560);
and U8357 (N_8357,N_7533,N_6322);
nor U8358 (N_8358,N_7327,N_7965);
nand U8359 (N_8359,N_6728,N_6836);
and U8360 (N_8360,N_6626,N_6436);
or U8361 (N_8361,N_7916,N_6727);
nor U8362 (N_8362,N_6164,N_7315);
or U8363 (N_8363,N_6723,N_7606);
or U8364 (N_8364,N_7134,N_6072);
xnor U8365 (N_8365,N_7683,N_7316);
nand U8366 (N_8366,N_7337,N_7393);
nor U8367 (N_8367,N_7774,N_6892);
and U8368 (N_8368,N_6949,N_7233);
nand U8369 (N_8369,N_7448,N_7627);
nor U8370 (N_8370,N_6759,N_7197);
nand U8371 (N_8371,N_6338,N_6629);
nand U8372 (N_8372,N_6332,N_7411);
and U8373 (N_8373,N_6075,N_6624);
xnor U8374 (N_8374,N_7459,N_7363);
xnor U8375 (N_8375,N_6797,N_7776);
nor U8376 (N_8376,N_6106,N_7080);
and U8377 (N_8377,N_6141,N_6487);
xnor U8378 (N_8378,N_7535,N_6708);
nand U8379 (N_8379,N_6214,N_7921);
nor U8380 (N_8380,N_6570,N_6558);
and U8381 (N_8381,N_6139,N_6845);
nor U8382 (N_8382,N_6710,N_7730);
nand U8383 (N_8383,N_7940,N_6355);
nor U8384 (N_8384,N_7169,N_6449);
or U8385 (N_8385,N_7397,N_6007);
or U8386 (N_8386,N_6533,N_7760);
nor U8387 (N_8387,N_7365,N_6619);
or U8388 (N_8388,N_7355,N_6596);
xor U8389 (N_8389,N_7202,N_6888);
or U8390 (N_8390,N_7969,N_6391);
and U8391 (N_8391,N_7096,N_6444);
or U8392 (N_8392,N_6593,N_7275);
and U8393 (N_8393,N_7968,N_6146);
nor U8394 (N_8394,N_6968,N_7697);
nor U8395 (N_8395,N_6335,N_7414);
nand U8396 (N_8396,N_6055,N_6381);
or U8397 (N_8397,N_7385,N_7793);
and U8398 (N_8398,N_6660,N_7970);
or U8399 (N_8399,N_6339,N_7132);
and U8400 (N_8400,N_7139,N_7737);
nor U8401 (N_8401,N_6208,N_6997);
nor U8402 (N_8402,N_7187,N_6265);
or U8403 (N_8403,N_7499,N_7252);
or U8404 (N_8404,N_6864,N_6302);
and U8405 (N_8405,N_6307,N_7064);
or U8406 (N_8406,N_7942,N_7454);
and U8407 (N_8407,N_7741,N_6550);
nor U8408 (N_8408,N_6676,N_6896);
and U8409 (N_8409,N_7300,N_7278);
and U8410 (N_8410,N_7374,N_7582);
xnor U8411 (N_8411,N_7527,N_7341);
nand U8412 (N_8412,N_7253,N_7041);
nand U8413 (N_8413,N_7553,N_7907);
nand U8414 (N_8414,N_6180,N_6750);
and U8415 (N_8415,N_7476,N_7720);
nand U8416 (N_8416,N_7294,N_7285);
nor U8417 (N_8417,N_7512,N_7176);
and U8418 (N_8418,N_7118,N_7382);
nand U8419 (N_8419,N_6450,N_6245);
or U8420 (N_8420,N_7434,N_7577);
nor U8421 (N_8421,N_6340,N_6228);
and U8422 (N_8422,N_7546,N_7906);
and U8423 (N_8423,N_7350,N_7934);
nand U8424 (N_8424,N_7824,N_7462);
nand U8425 (N_8425,N_6382,N_7917);
and U8426 (N_8426,N_6044,N_6667);
or U8427 (N_8427,N_7109,N_6659);
nor U8428 (N_8428,N_6019,N_6838);
xnor U8429 (N_8429,N_7095,N_6770);
or U8430 (N_8430,N_7098,N_7047);
and U8431 (N_8431,N_6868,N_7384);
xnor U8432 (N_8432,N_6195,N_7566);
and U8433 (N_8433,N_7286,N_6620);
and U8434 (N_8434,N_7222,N_6001);
xnor U8435 (N_8435,N_6893,N_6573);
or U8436 (N_8436,N_6148,N_7161);
nor U8437 (N_8437,N_6524,N_6685);
nor U8438 (N_8438,N_7046,N_7994);
or U8439 (N_8439,N_7088,N_7280);
nor U8440 (N_8440,N_7063,N_7259);
xnor U8441 (N_8441,N_7432,N_6915);
nor U8442 (N_8442,N_6886,N_7229);
or U8443 (N_8443,N_7953,N_6606);
or U8444 (N_8444,N_7780,N_6129);
xnor U8445 (N_8445,N_6179,N_7310);
nand U8446 (N_8446,N_6577,N_6267);
or U8447 (N_8447,N_7256,N_6756);
or U8448 (N_8448,N_6945,N_7311);
or U8449 (N_8449,N_7997,N_6520);
or U8450 (N_8450,N_7195,N_6740);
or U8451 (N_8451,N_7820,N_6696);
nand U8452 (N_8452,N_7733,N_6441);
nor U8453 (N_8453,N_6985,N_6298);
nand U8454 (N_8454,N_7513,N_7036);
nor U8455 (N_8455,N_7537,N_7028);
and U8456 (N_8456,N_6701,N_7056);
xor U8457 (N_8457,N_7583,N_6719);
xor U8458 (N_8458,N_7494,N_6548);
nor U8459 (N_8459,N_6393,N_6912);
nand U8460 (N_8460,N_7273,N_6231);
and U8461 (N_8461,N_7180,N_6348);
or U8462 (N_8462,N_7626,N_7198);
and U8463 (N_8463,N_6074,N_7924);
or U8464 (N_8464,N_6508,N_7170);
xnor U8465 (N_8465,N_6690,N_6631);
nand U8466 (N_8466,N_6224,N_6318);
xnor U8467 (N_8467,N_7556,N_7153);
xnor U8468 (N_8468,N_7403,N_7141);
xnor U8469 (N_8469,N_7324,N_7304);
xor U8470 (N_8470,N_7415,N_7009);
nor U8471 (N_8471,N_7230,N_7204);
xnor U8472 (N_8472,N_7221,N_6936);
or U8473 (N_8473,N_6130,N_6274);
xor U8474 (N_8474,N_6213,N_7944);
nor U8475 (N_8475,N_6260,N_6804);
xor U8476 (N_8476,N_7572,N_6760);
and U8477 (N_8477,N_7966,N_7573);
nor U8478 (N_8478,N_7870,N_6466);
or U8479 (N_8479,N_6438,N_7061);
nor U8480 (N_8480,N_6932,N_7816);
or U8481 (N_8481,N_6939,N_6982);
nand U8482 (N_8482,N_6633,N_7477);
nor U8483 (N_8483,N_6679,N_6090);
xor U8484 (N_8484,N_6563,N_6201);
nor U8485 (N_8485,N_6033,N_7354);
xnor U8486 (N_8486,N_6857,N_7163);
or U8487 (N_8487,N_7313,N_7555);
xor U8488 (N_8488,N_6437,N_6266);
and U8489 (N_8489,N_6517,N_7574);
xor U8490 (N_8490,N_7584,N_6758);
nand U8491 (N_8491,N_7255,N_6697);
and U8492 (N_8492,N_6166,N_7261);
and U8493 (N_8493,N_6584,N_7276);
xor U8494 (N_8494,N_7092,N_6270);
or U8495 (N_8495,N_6108,N_6618);
or U8496 (N_8496,N_7349,N_7521);
or U8497 (N_8497,N_6174,N_7470);
and U8498 (N_8498,N_6167,N_6233);
nand U8499 (N_8499,N_6672,N_6030);
or U8500 (N_8500,N_6156,N_7463);
nor U8501 (N_8501,N_6435,N_6351);
xor U8502 (N_8502,N_7779,N_7709);
nand U8503 (N_8503,N_7530,N_7988);
nand U8504 (N_8504,N_7200,N_7964);
xor U8505 (N_8505,N_7721,N_7911);
xor U8506 (N_8506,N_7664,N_6451);
or U8507 (N_8507,N_6736,N_6105);
and U8508 (N_8508,N_7049,N_6623);
nand U8509 (N_8509,N_6774,N_6744);
and U8510 (N_8510,N_7216,N_6678);
or U8511 (N_8511,N_6388,N_6863);
xor U8512 (N_8512,N_6829,N_6947);
xor U8513 (N_8513,N_6668,N_6480);
and U8514 (N_8514,N_6490,N_6769);
and U8515 (N_8515,N_7394,N_6202);
xor U8516 (N_8516,N_7668,N_6036);
and U8517 (N_8517,N_7862,N_6919);
nand U8518 (N_8518,N_7748,N_6151);
or U8519 (N_8519,N_7150,N_6408);
and U8520 (N_8520,N_6636,N_7547);
and U8521 (N_8521,N_7505,N_6691);
and U8522 (N_8522,N_6052,N_7813);
and U8523 (N_8523,N_6188,N_7097);
and U8524 (N_8524,N_7523,N_6153);
nand U8525 (N_8525,N_7514,N_7542);
xor U8526 (N_8526,N_7069,N_6902);
nand U8527 (N_8527,N_7710,N_6099);
or U8528 (N_8528,N_6023,N_7461);
nand U8529 (N_8529,N_7554,N_6002);
xor U8530 (N_8530,N_6448,N_6825);
nor U8531 (N_8531,N_7787,N_7823);
or U8532 (N_8532,N_7232,N_6134);
nand U8533 (N_8533,N_7019,N_7223);
xnor U8534 (N_8534,N_6555,N_6661);
nor U8535 (N_8535,N_6576,N_6483);
nand U8536 (N_8536,N_7694,N_6814);
nand U8537 (N_8537,N_6295,N_6874);
xnor U8538 (N_8538,N_6682,N_6980);
nor U8539 (N_8539,N_6098,N_6846);
xnor U8540 (N_8540,N_6812,N_6114);
or U8541 (N_8541,N_6359,N_7390);
nand U8542 (N_8542,N_7717,N_7541);
nor U8543 (N_8543,N_6847,N_6746);
or U8544 (N_8544,N_7646,N_7568);
nand U8545 (N_8545,N_6455,N_7893);
or U8546 (N_8546,N_7832,N_7190);
nor U8547 (N_8547,N_7682,N_7874);
nor U8548 (N_8548,N_7348,N_7291);
or U8549 (N_8549,N_6154,N_6158);
xor U8550 (N_8550,N_7947,N_7186);
xor U8551 (N_8551,N_7090,N_7306);
xnor U8552 (N_8552,N_7201,N_7042);
nand U8553 (N_8553,N_7481,N_6039);
and U8554 (N_8554,N_7497,N_7713);
xor U8555 (N_8555,N_7123,N_6622);
or U8556 (N_8556,N_6903,N_6308);
and U8557 (N_8557,N_7843,N_6027);
or U8558 (N_8558,N_7849,N_6246);
or U8559 (N_8559,N_6171,N_6373);
xnor U8560 (N_8560,N_6951,N_6589);
and U8561 (N_8561,N_6579,N_6367);
or U8562 (N_8562,N_6831,N_7100);
nor U8563 (N_8563,N_6317,N_6810);
nor U8564 (N_8564,N_7453,N_6101);
nand U8565 (N_8565,N_6654,N_7844);
or U8566 (N_8566,N_7519,N_7837);
xor U8567 (N_8567,N_6973,N_6232);
nand U8568 (N_8568,N_6282,N_6257);
or U8569 (N_8569,N_6289,N_7044);
nand U8570 (N_8570,N_7850,N_7129);
and U8571 (N_8571,N_6684,N_6494);
nor U8572 (N_8572,N_7896,N_7235);
nor U8573 (N_8573,N_6789,N_7166);
nand U8574 (N_8574,N_7466,N_7218);
nand U8575 (N_8575,N_6291,N_6481);
nor U8576 (N_8576,N_6995,N_6544);
and U8577 (N_8577,N_6168,N_6107);
xor U8578 (N_8578,N_6640,N_7650);
and U8579 (N_8579,N_6028,N_6241);
or U8580 (N_8580,N_7502,N_7558);
or U8581 (N_8581,N_7035,N_6869);
or U8582 (N_8582,N_7071,N_7031);
nand U8583 (N_8583,N_7240,N_7822);
xor U8584 (N_8584,N_6861,N_6071);
or U8585 (N_8585,N_6529,N_6972);
or U8586 (N_8586,N_7496,N_7833);
nand U8587 (N_8587,N_6834,N_6655);
nor U8588 (N_8588,N_6803,N_7786);
and U8589 (N_8589,N_6835,N_6163);
or U8590 (N_8590,N_7561,N_7258);
nand U8591 (N_8591,N_7321,N_6380);
nand U8592 (N_8592,N_6254,N_7846);
and U8593 (N_8593,N_6880,N_7369);
xor U8594 (N_8594,N_6060,N_7022);
and U8595 (N_8595,N_6850,N_7888);
and U8596 (N_8596,N_7880,N_6527);
or U8597 (N_8597,N_7460,N_7783);
nand U8598 (N_8598,N_6247,N_6715);
and U8599 (N_8599,N_6943,N_7600);
nand U8600 (N_8600,N_6155,N_6843);
nand U8601 (N_8601,N_7137,N_7827);
nor U8602 (N_8602,N_7676,N_6981);
nor U8603 (N_8603,N_6253,N_7115);
xnor U8604 (N_8604,N_7173,N_6605);
nand U8605 (N_8605,N_7902,N_7825);
nor U8606 (N_8606,N_6898,N_7909);
nor U8607 (N_8607,N_6765,N_7894);
nand U8608 (N_8608,N_6574,N_6170);
nand U8609 (N_8609,N_6556,N_6425);
nor U8610 (N_8610,N_7531,N_7762);
nor U8611 (N_8611,N_6811,N_7806);
xor U8612 (N_8612,N_6116,N_7576);
and U8613 (N_8613,N_7491,N_7642);
nand U8614 (N_8614,N_6998,N_7226);
or U8615 (N_8615,N_6411,N_7480);
and U8616 (N_8616,N_7076,N_7279);
or U8617 (N_8617,N_6597,N_6602);
and U8618 (N_8618,N_7307,N_7026);
and U8619 (N_8619,N_6671,N_6783);
nand U8620 (N_8620,N_6387,N_7712);
nor U8621 (N_8621,N_6683,N_6193);
nor U8622 (N_8622,N_7706,N_7373);
or U8623 (N_8623,N_6384,N_7629);
and U8624 (N_8624,N_7234,N_6395);
xnor U8625 (N_8625,N_7620,N_6990);
nor U8626 (N_8626,N_7059,N_6354);
xor U8627 (N_8627,N_7913,N_7597);
nand U8628 (N_8628,N_6235,N_6976);
and U8629 (N_8629,N_6131,N_6230);
nand U8630 (N_8630,N_6514,N_7181);
xor U8631 (N_8631,N_6015,N_7602);
and U8632 (N_8632,N_6400,N_7625);
xor U8633 (N_8633,N_6538,N_7551);
or U8634 (N_8634,N_7670,N_6562);
or U8635 (N_8635,N_7425,N_6848);
nor U8636 (N_8636,N_7647,N_6429);
or U8637 (N_8637,N_6073,N_6536);
nor U8638 (N_8638,N_7881,N_6928);
nor U8639 (N_8639,N_7179,N_6453);
and U8640 (N_8640,N_7800,N_7972);
or U8641 (N_8641,N_7368,N_7651);
nor U8642 (N_8642,N_6542,N_6209);
xor U8643 (N_8643,N_6754,N_6290);
nand U8644 (N_8644,N_7157,N_6181);
nand U8645 (N_8645,N_7628,N_6024);
xor U8646 (N_8646,N_6485,N_6041);
xnor U8647 (N_8647,N_7027,N_6066);
nor U8648 (N_8648,N_6920,N_6610);
nor U8649 (N_8649,N_6712,N_6496);
xor U8650 (N_8650,N_7192,N_6639);
nor U8651 (N_8651,N_6948,N_6518);
nand U8652 (N_8652,N_7501,N_7652);
nand U8653 (N_8653,N_7869,N_7510);
xor U8654 (N_8654,N_6183,N_6285);
nor U8655 (N_8655,N_6788,N_6821);
xnor U8656 (N_8656,N_6407,N_7050);
nand U8657 (N_8657,N_6464,N_6479);
or U8658 (N_8658,N_7339,N_6941);
xnor U8659 (N_8659,N_6043,N_6031);
nor U8660 (N_8660,N_7039,N_6409);
xnor U8661 (N_8661,N_7879,N_6734);
nor U8662 (N_8662,N_6456,N_6250);
nor U8663 (N_8663,N_7828,N_7299);
or U8664 (N_8664,N_6907,N_7515);
or U8665 (N_8665,N_7231,N_6651);
xor U8666 (N_8666,N_6674,N_6142);
or U8667 (N_8667,N_7662,N_6499);
nor U8668 (N_8668,N_6046,N_6657);
xnor U8669 (N_8669,N_6011,N_7990);
nand U8670 (N_8670,N_7053,N_6509);
xor U8671 (N_8671,N_7108,N_6877);
nand U8672 (N_8672,N_6988,N_6999);
xnor U8673 (N_8673,N_6782,N_7451);
xnor U8674 (N_8674,N_7409,N_7766);
or U8675 (N_8675,N_6925,N_6331);
or U8676 (N_8676,N_6426,N_6987);
and U8677 (N_8677,N_7520,N_6243);
nand U8678 (N_8678,N_6557,N_7677);
xor U8679 (N_8679,N_7030,N_6133);
or U8680 (N_8680,N_7247,N_7376);
nand U8681 (N_8681,N_6944,N_6248);
nor U8682 (N_8682,N_7707,N_7978);
and U8683 (N_8683,N_6476,N_6772);
nand U8684 (N_8684,N_7564,N_7160);
nand U8685 (N_8685,N_6189,N_7091);
nand U8686 (N_8686,N_6689,N_6866);
nand U8687 (N_8687,N_7479,N_6421);
xor U8688 (N_8688,N_7992,N_6796);
xnor U8689 (N_8689,N_7673,N_7799);
nor U8690 (N_8690,N_6350,N_6883);
nand U8691 (N_8691,N_6608,N_7332);
and U8692 (N_8692,N_6152,N_7396);
nor U8693 (N_8693,N_7146,N_6296);
and U8694 (N_8694,N_7641,N_7539);
and U8695 (N_8695,N_7125,N_6634);
nand U8696 (N_8696,N_6837,N_7029);
and U8697 (N_8697,N_6326,N_6959);
xor U8698 (N_8698,N_7930,N_7790);
nor U8699 (N_8699,N_6345,N_7320);
and U8700 (N_8700,N_6300,N_6900);
xor U8701 (N_8701,N_7826,N_6320);
and U8702 (N_8702,N_6551,N_7208);
or U8703 (N_8703,N_7689,N_6360);
nor U8704 (N_8704,N_7344,N_6037);
xnor U8705 (N_8705,N_7308,N_7144);
nor U8706 (N_8706,N_7788,N_7468);
nand U8707 (N_8707,N_7014,N_6729);
or U8708 (N_8708,N_6793,N_7058);
xor U8709 (N_8709,N_6994,N_6611);
and U8710 (N_8710,N_6457,N_7789);
xnor U8711 (N_8711,N_6511,N_6396);
nand U8712 (N_8712,N_6079,N_7087);
xnor U8713 (N_8713,N_7698,N_6029);
nand U8714 (N_8714,N_7110,N_6680);
nand U8715 (N_8715,N_7882,N_7609);
and U8716 (N_8716,N_6212,N_6219);
and U8717 (N_8717,N_6942,N_6603);
nand U8718 (N_8718,N_6926,N_7006);
nor U8719 (N_8719,N_7093,N_7904);
and U8720 (N_8720,N_6975,N_7638);
nand U8721 (N_8721,N_6016,N_6953);
or U8722 (N_8722,N_7617,N_7094);
and U8723 (N_8723,N_6157,N_7543);
nand U8724 (N_8724,N_6791,N_7290);
nand U8725 (N_8725,N_6410,N_6675);
nand U8726 (N_8726,N_7238,N_6730);
nand U8727 (N_8727,N_6126,N_6827);
nand U8728 (N_8728,N_6652,N_6194);
nor U8729 (N_8729,N_6471,N_7236);
nand U8730 (N_8730,N_7571,N_6598);
xor U8731 (N_8731,N_7592,N_7587);
nand U8732 (N_8732,N_7084,N_7589);
and U8733 (N_8733,N_7423,N_6984);
xnor U8734 (N_8734,N_7008,N_7839);
and U8735 (N_8735,N_7829,N_6205);
xor U8736 (N_8736,N_7185,N_7072);
nand U8737 (N_8737,N_6800,N_6109);
nand U8738 (N_8738,N_7483,N_7325);
and U8739 (N_8739,N_7802,N_6482);
and U8740 (N_8740,N_7099,N_7452);
nor U8741 (N_8741,N_7695,N_7884);
nor U8742 (N_8742,N_7746,N_6034);
and U8743 (N_8743,N_6755,N_7897);
nor U8744 (N_8744,N_7559,N_7769);
xnor U8745 (N_8745,N_7408,N_7621);
or U8746 (N_8746,N_6064,N_7107);
or U8747 (N_8747,N_7898,N_6227);
nor U8748 (N_8748,N_7104,N_7389);
or U8749 (N_8749,N_7135,N_6858);
nand U8750 (N_8750,N_6432,N_7126);
nand U8751 (N_8751,N_7034,N_7538);
xor U8752 (N_8752,N_7861,N_7217);
xor U8753 (N_8753,N_6549,N_6971);
and U8754 (N_8754,N_7759,N_6275);
nor U8755 (N_8755,N_7331,N_6958);
nand U8756 (N_8756,N_6176,N_7723);
nand U8757 (N_8757,N_7753,N_7511);
xor U8758 (N_8758,N_6901,N_7669);
xnor U8759 (N_8759,N_7065,N_7581);
and U8760 (N_8760,N_7522,N_7590);
or U8761 (N_8761,N_6545,N_6911);
nand U8762 (N_8762,N_7675,N_6649);
or U8763 (N_8763,N_7985,N_6234);
nand U8764 (N_8764,N_6117,N_7277);
nand U8765 (N_8765,N_6442,N_6311);
or U8766 (N_8766,N_6143,N_7873);
xor U8767 (N_8767,N_7205,N_7003);
nor U8768 (N_8768,N_7923,N_7674);
or U8769 (N_8769,N_6172,N_7188);
nand U8770 (N_8770,N_6159,N_6443);
nor U8771 (N_8771,N_6855,N_6199);
or U8772 (N_8772,N_7498,N_7507);
nand U8773 (N_8773,N_7724,N_7899);
nor U8774 (N_8774,N_7841,N_7744);
and U8775 (N_8775,N_7392,N_6571);
and U8776 (N_8776,N_7608,N_7771);
xnor U8777 (N_8777,N_7045,N_6122);
xnor U8778 (N_8778,N_7666,N_7133);
nand U8779 (N_8779,N_7265,N_7012);
xor U8780 (N_8780,N_6102,N_6747);
nor U8781 (N_8781,N_7876,N_7892);
nand U8782 (N_8782,N_7653,N_6817);
or U8783 (N_8783,N_6802,N_7242);
or U8784 (N_8784,N_7719,N_6616);
nand U8785 (N_8785,N_6786,N_7986);
or U8786 (N_8786,N_6191,N_6078);
xor U8787 (N_8787,N_6569,N_6934);
xnor U8788 (N_8788,N_6454,N_6873);
and U8789 (N_8789,N_7984,N_6433);
or U8790 (N_8790,N_6909,N_7296);
xor U8791 (N_8791,N_6309,N_7594);
and U8792 (N_8792,N_6666,N_7010);
xor U8793 (N_8793,N_7701,N_7933);
or U8794 (N_8794,N_6383,N_6884);
and U8795 (N_8795,N_7819,N_6292);
nor U8796 (N_8796,N_6870,N_6287);
nor U8797 (N_8797,N_6096,N_7025);
xnor U8798 (N_8798,N_6404,N_6121);
and U8799 (N_8799,N_6702,N_7057);
xnor U8800 (N_8800,N_7268,N_6991);
and U8801 (N_8801,N_7457,N_6885);
or U8802 (N_8802,N_6059,N_7552);
and U8803 (N_8803,N_7756,N_7878);
or U8804 (N_8804,N_6484,N_6648);
or U8805 (N_8805,N_6776,N_7954);
and U8806 (N_8806,N_6824,N_6225);
xnor U8807 (N_8807,N_6504,N_7250);
nor U8808 (N_8808,N_6424,N_6460);
and U8809 (N_8809,N_7757,N_6081);
and U8810 (N_8810,N_7478,N_7323);
nor U8811 (N_8811,N_7544,N_6306);
or U8812 (N_8812,N_7925,N_6721);
or U8813 (N_8813,N_6795,N_7949);
nand U8814 (N_8814,N_7649,N_7422);
or U8815 (N_8815,N_6358,N_6087);
nand U8816 (N_8816,N_7995,N_6700);
nor U8817 (N_8817,N_7440,N_7830);
or U8818 (N_8818,N_6921,N_7495);
or U8819 (N_8819,N_7248,N_7449);
and U8820 (N_8820,N_7623,N_6258);
nand U8821 (N_8821,N_6417,N_7112);
nand U8822 (N_8822,N_6374,N_7156);
nor U8823 (N_8823,N_6502,N_7336);
or U8824 (N_8824,N_7433,N_6347);
or U8825 (N_8825,N_7998,N_7704);
and U8826 (N_8826,N_6625,N_7903);
xor U8827 (N_8827,N_7446,N_6138);
and U8828 (N_8828,N_6910,N_7963);
xnor U8829 (N_8829,N_6045,N_7863);
nor U8830 (N_8830,N_6552,N_6687);
nand U8831 (N_8831,N_6745,N_6057);
xor U8832 (N_8832,N_6127,N_7901);
nand U8833 (N_8833,N_7736,N_6752);
nor U8834 (N_8834,N_7399,N_6369);
nand U8835 (N_8835,N_6173,N_6012);
nand U8836 (N_8836,N_6534,N_7400);
xnor U8837 (N_8837,N_6175,N_6867);
xor U8838 (N_8838,N_7174,N_6741);
xor U8839 (N_8839,N_7791,N_7122);
nor U8840 (N_8840,N_6226,N_7116);
xor U8841 (N_8841,N_7613,N_7114);
xor U8842 (N_8842,N_7420,N_7941);
and U8843 (N_8843,N_6519,N_6646);
nor U8844 (N_8844,N_6541,N_6357);
or U8845 (N_8845,N_7458,N_7945);
or U8846 (N_8846,N_7524,N_7271);
nor U8847 (N_8847,N_7619,N_7595);
xnor U8848 (N_8848,N_7671,N_6807);
xor U8849 (N_8849,N_6665,N_7297);
nor U8850 (N_8850,N_6288,N_6613);
and U8851 (N_8851,N_7536,N_6040);
or U8852 (N_8852,N_7269,N_6989);
nand U8853 (N_8853,N_6293,N_7716);
xnor U8854 (N_8854,N_6144,N_6938);
nand U8855 (N_8855,N_7959,N_7705);
and U8856 (N_8856,N_6268,N_6420);
or U8857 (N_8857,N_7740,N_6053);
xnor U8858 (N_8858,N_7960,N_6273);
nor U8859 (N_8859,N_6467,N_6916);
nor U8860 (N_8860,N_6000,N_7079);
xnor U8861 (N_8861,N_7075,N_7361);
nor U8862 (N_8862,N_6785,N_7364);
and U8863 (N_8863,N_7636,N_6310);
or U8864 (N_8864,N_7506,N_6688);
nor U8865 (N_8865,N_6695,N_7004);
xor U8866 (N_8866,N_6014,N_7961);
nand U8867 (N_8867,N_6720,N_6779);
xnor U8868 (N_8868,N_6775,N_6091);
nand U8869 (N_8869,N_6342,N_6140);
xor U8870 (N_8870,N_6111,N_6398);
or U8871 (N_8871,N_7567,N_7758);
nor U8872 (N_8872,N_7958,N_7914);
or U8873 (N_8873,N_7754,N_7398);
or U8874 (N_8874,N_6062,N_6664);
nor U8875 (N_8875,N_7688,N_7887);
nand U8876 (N_8876,N_7214,N_6543);
and U8877 (N_8877,N_7362,N_7637);
nor U8878 (N_8878,N_7569,N_6083);
nand U8879 (N_8879,N_6790,N_6601);
and U8880 (N_8880,N_6068,N_6842);
nand U8881 (N_8881,N_6497,N_6218);
or U8882 (N_8882,N_6093,N_6565);
nand U8883 (N_8883,N_7782,N_6178);
nand U8884 (N_8884,N_7610,N_6718);
or U8885 (N_8885,N_7633,N_7322);
xor U8886 (N_8886,N_6440,N_7447);
xor U8887 (N_8887,N_6390,N_7657);
nand U8888 (N_8888,N_7937,N_6240);
xor U8889 (N_8889,N_7171,N_7347);
nor U8890 (N_8890,N_7032,N_6704);
and U8891 (N_8891,N_7659,N_6304);
and U8892 (N_8892,N_6377,N_7575);
and U8893 (N_8893,N_7853,N_7484);
xor U8894 (N_8894,N_6063,N_7184);
nand U8895 (N_8895,N_7346,N_7751);
nor U8896 (N_8896,N_6478,N_6389);
or U8897 (N_8897,N_6137,N_7085);
and U8898 (N_8898,N_7975,N_6500);
nand U8899 (N_8899,N_6503,N_7908);
and U8900 (N_8900,N_7578,N_7237);
nor U8901 (N_8901,N_7980,N_7302);
nor U8902 (N_8902,N_7074,N_7441);
and U8903 (N_8903,N_6568,N_7692);
xnor U8904 (N_8904,N_6799,N_7755);
or U8905 (N_8905,N_6277,N_6599);
nor U8906 (N_8906,N_7932,N_6567);
xor U8907 (N_8907,N_7905,N_7974);
nand U8908 (N_8908,N_7351,N_6826);
and U8909 (N_8909,N_6336,N_6535);
xor U8910 (N_8910,N_7630,N_6368);
and U8911 (N_8911,N_6084,N_6732);
or U8912 (N_8912,N_6764,N_6070);
xnor U8913 (N_8913,N_7378,N_7996);
or U8914 (N_8914,N_6018,N_6299);
nand U8915 (N_8915,N_6048,N_7281);
nand U8916 (N_8916,N_7154,N_7410);
and U8917 (N_8917,N_6003,N_7052);
and U8918 (N_8918,N_6469,N_7534);
nor U8919 (N_8919,N_6768,N_6349);
and U8920 (N_8920,N_7667,N_7431);
nand U8921 (N_8921,N_6515,N_6839);
xor U8922 (N_8922,N_7089,N_7486);
and U8923 (N_8923,N_7615,N_6507);
or U8924 (N_8924,N_6486,N_7303);
nand U8925 (N_8925,N_6751,N_7955);
or U8926 (N_8926,N_6216,N_6767);
xnor U8927 (N_8927,N_6401,N_6082);
and U8928 (N_8928,N_6010,N_7193);
or U8929 (N_8929,N_7358,N_7702);
xnor U8930 (N_8930,N_6967,N_7593);
and U8931 (N_8931,N_6069,N_7728);
xor U8932 (N_8932,N_7860,N_6889);
nand U8933 (N_8933,N_7011,N_7023);
nand U8934 (N_8934,N_6236,N_6263);
or U8935 (N_8935,N_6645,N_7814);
nand U8936 (N_8936,N_7318,N_6315);
or U8937 (N_8937,N_7282,N_7338);
nor U8938 (N_8938,N_6491,N_7162);
xor U8939 (N_8939,N_6722,N_7387);
nor U8940 (N_8940,N_6392,N_6662);
nor U8941 (N_8941,N_7952,N_6237);
and U8942 (N_8942,N_6321,N_6038);
and U8943 (N_8943,N_6017,N_6474);
xor U8944 (N_8944,N_6125,N_6005);
and U8945 (N_8945,N_7366,N_6058);
nor U8946 (N_8946,N_6707,N_7854);
and U8947 (N_8947,N_7738,N_6714);
nand U8948 (N_8948,N_7767,N_6493);
or U8949 (N_8949,N_6957,N_7607);
or U8950 (N_8950,N_7845,N_6211);
nand U8951 (N_8951,N_7371,N_7383);
nand U8952 (N_8952,N_6470,N_7005);
xnor U8953 (N_8953,N_7919,N_7225);
nor U8954 (N_8954,N_7848,N_7018);
nor U8955 (N_8955,N_6887,N_7798);
nand U8956 (N_8956,N_7490,N_6147);
or U8957 (N_8957,N_6876,N_7489);
nand U8958 (N_8958,N_7353,N_6207);
nand U8959 (N_8959,N_7856,N_7545);
nor U8960 (N_8960,N_7943,N_7377);
and U8961 (N_8961,N_6324,N_7401);
xor U8962 (N_8962,N_7938,N_6239);
and U8963 (N_8963,N_7687,N_7427);
nor U8964 (N_8964,N_6169,N_7770);
nand U8965 (N_8965,N_6203,N_7926);
and U8966 (N_8966,N_7680,N_7183);
xnor U8967 (N_8967,N_7189,N_6095);
nand U8968 (N_8968,N_6088,N_7289);
xnor U8969 (N_8969,N_6966,N_6572);
and U8970 (N_8970,N_7055,N_6492);
or U8971 (N_8971,N_6462,N_6952);
nand U8972 (N_8972,N_6329,N_6080);
or U8973 (N_8973,N_7314,N_7640);
xnor U8974 (N_8974,N_6531,N_6150);
xor U8975 (N_8975,N_7215,N_6586);
xnor U8976 (N_8976,N_6196,N_7971);
and U8977 (N_8977,N_6238,N_7868);
and U8978 (N_8978,N_7220,N_7040);
nand U8979 (N_8979,N_7910,N_7419);
xnor U8980 (N_8980,N_6813,N_7048);
or U8981 (N_8981,N_7504,N_7224);
nand U8982 (N_8982,N_7143,N_6897);
xnor U8983 (N_8983,N_6553,N_7614);
xor U8984 (N_8984,N_7043,N_7342);
xor U8985 (N_8985,N_7060,N_6937);
nor U8986 (N_8986,N_6853,N_7113);
or U8987 (N_8987,N_7877,N_7742);
nand U8988 (N_8988,N_7485,N_7077);
or U8989 (N_8989,N_6244,N_6822);
and U8990 (N_8990,N_6983,N_7021);
nor U8991 (N_8991,N_6950,N_7249);
nor U8992 (N_8992,N_6149,N_7328);
or U8993 (N_8993,N_7847,N_7764);
nand U8994 (N_8994,N_7002,N_6566);
and U8995 (N_8995,N_6516,N_7865);
nor U8996 (N_8996,N_7585,N_6798);
and U8997 (N_8997,N_7808,N_7663);
xnor U8998 (N_8998,N_6468,N_6946);
or U8999 (N_8999,N_7586,N_7270);
nand U9000 (N_9000,N_6326,N_7598);
or U9001 (N_9001,N_7579,N_6451);
nand U9002 (N_9002,N_7548,N_7804);
or U9003 (N_9003,N_7970,N_7856);
xor U9004 (N_9004,N_7934,N_7094);
nor U9005 (N_9005,N_6892,N_7984);
xnor U9006 (N_9006,N_6272,N_7347);
and U9007 (N_9007,N_6749,N_6854);
xnor U9008 (N_9008,N_6364,N_7261);
or U9009 (N_9009,N_6464,N_7886);
xnor U9010 (N_9010,N_7606,N_6678);
nand U9011 (N_9011,N_7127,N_7649);
and U9012 (N_9012,N_6100,N_6356);
nor U9013 (N_9013,N_6315,N_7952);
nand U9014 (N_9014,N_6006,N_6273);
nand U9015 (N_9015,N_6418,N_7935);
xor U9016 (N_9016,N_7001,N_6258);
or U9017 (N_9017,N_6817,N_6882);
nand U9018 (N_9018,N_6885,N_7911);
nor U9019 (N_9019,N_7665,N_6780);
and U9020 (N_9020,N_7966,N_7516);
nor U9021 (N_9021,N_6884,N_7382);
xor U9022 (N_9022,N_6135,N_7167);
xnor U9023 (N_9023,N_7120,N_6661);
xor U9024 (N_9024,N_6890,N_6846);
nand U9025 (N_9025,N_7552,N_6296);
and U9026 (N_9026,N_6740,N_6749);
and U9027 (N_9027,N_6894,N_7725);
xor U9028 (N_9028,N_7879,N_6353);
xnor U9029 (N_9029,N_6487,N_6296);
or U9030 (N_9030,N_7085,N_6043);
and U9031 (N_9031,N_7175,N_7525);
nor U9032 (N_9032,N_6367,N_6727);
nor U9033 (N_9033,N_6739,N_6279);
nand U9034 (N_9034,N_6400,N_6585);
xor U9035 (N_9035,N_6191,N_7647);
xor U9036 (N_9036,N_7281,N_7742);
or U9037 (N_9037,N_7912,N_7929);
and U9038 (N_9038,N_6529,N_7156);
and U9039 (N_9039,N_6537,N_7100);
and U9040 (N_9040,N_6119,N_6950);
and U9041 (N_9041,N_6857,N_7002);
and U9042 (N_9042,N_7215,N_7545);
nor U9043 (N_9043,N_6431,N_7293);
and U9044 (N_9044,N_6003,N_7637);
and U9045 (N_9045,N_6722,N_6020);
or U9046 (N_9046,N_6778,N_7165);
and U9047 (N_9047,N_6631,N_7315);
nor U9048 (N_9048,N_7515,N_6633);
nand U9049 (N_9049,N_6414,N_6601);
xnor U9050 (N_9050,N_6095,N_6300);
or U9051 (N_9051,N_7040,N_6908);
nand U9052 (N_9052,N_7932,N_7772);
or U9053 (N_9053,N_7407,N_7753);
and U9054 (N_9054,N_7467,N_7774);
nor U9055 (N_9055,N_7513,N_7866);
xnor U9056 (N_9056,N_6099,N_6450);
and U9057 (N_9057,N_7029,N_7890);
and U9058 (N_9058,N_7181,N_6687);
and U9059 (N_9059,N_7061,N_6171);
nor U9060 (N_9060,N_7086,N_6264);
and U9061 (N_9061,N_6578,N_6607);
nand U9062 (N_9062,N_7746,N_7409);
nand U9063 (N_9063,N_6129,N_6836);
nor U9064 (N_9064,N_6392,N_6846);
xnor U9065 (N_9065,N_7634,N_6637);
and U9066 (N_9066,N_6026,N_6507);
nand U9067 (N_9067,N_7879,N_6892);
xor U9068 (N_9068,N_6164,N_7526);
and U9069 (N_9069,N_6967,N_6267);
or U9070 (N_9070,N_6215,N_6005);
and U9071 (N_9071,N_7391,N_6458);
and U9072 (N_9072,N_6567,N_7775);
or U9073 (N_9073,N_6941,N_7568);
or U9074 (N_9074,N_6064,N_7787);
or U9075 (N_9075,N_6964,N_6806);
nor U9076 (N_9076,N_7265,N_7030);
nand U9077 (N_9077,N_6003,N_7350);
xor U9078 (N_9078,N_6402,N_6347);
nor U9079 (N_9079,N_7112,N_6326);
nand U9080 (N_9080,N_7333,N_6584);
xor U9081 (N_9081,N_6574,N_7761);
xor U9082 (N_9082,N_7274,N_6863);
nand U9083 (N_9083,N_7757,N_6007);
or U9084 (N_9084,N_6277,N_6136);
nor U9085 (N_9085,N_6005,N_7471);
xnor U9086 (N_9086,N_6519,N_7268);
nand U9087 (N_9087,N_7607,N_7081);
nor U9088 (N_9088,N_6306,N_7902);
and U9089 (N_9089,N_7891,N_6453);
nor U9090 (N_9090,N_7476,N_7934);
xor U9091 (N_9091,N_7420,N_7452);
and U9092 (N_9092,N_6222,N_7428);
nor U9093 (N_9093,N_6218,N_6523);
and U9094 (N_9094,N_7793,N_7294);
nor U9095 (N_9095,N_7462,N_6694);
nand U9096 (N_9096,N_7635,N_7040);
nand U9097 (N_9097,N_7327,N_7939);
nand U9098 (N_9098,N_7054,N_7254);
nand U9099 (N_9099,N_7348,N_7444);
nor U9100 (N_9100,N_6946,N_6449);
or U9101 (N_9101,N_6371,N_6416);
nor U9102 (N_9102,N_7121,N_6373);
nor U9103 (N_9103,N_6239,N_7249);
xnor U9104 (N_9104,N_6306,N_7330);
nand U9105 (N_9105,N_6793,N_6159);
nor U9106 (N_9106,N_7487,N_7969);
nand U9107 (N_9107,N_7276,N_6540);
xnor U9108 (N_9108,N_6109,N_6458);
nand U9109 (N_9109,N_7135,N_6622);
or U9110 (N_9110,N_7884,N_6400);
and U9111 (N_9111,N_6905,N_6017);
and U9112 (N_9112,N_6527,N_6474);
nor U9113 (N_9113,N_7837,N_7685);
nor U9114 (N_9114,N_7869,N_6326);
xnor U9115 (N_9115,N_7000,N_7463);
and U9116 (N_9116,N_7895,N_6397);
nor U9117 (N_9117,N_6714,N_7105);
or U9118 (N_9118,N_7149,N_6642);
nand U9119 (N_9119,N_6385,N_7981);
or U9120 (N_9120,N_6240,N_7814);
and U9121 (N_9121,N_6243,N_7096);
and U9122 (N_9122,N_6791,N_6920);
xor U9123 (N_9123,N_7987,N_6092);
and U9124 (N_9124,N_7898,N_7431);
xor U9125 (N_9125,N_7199,N_6996);
and U9126 (N_9126,N_7329,N_7099);
xor U9127 (N_9127,N_7444,N_6796);
nor U9128 (N_9128,N_7173,N_6049);
or U9129 (N_9129,N_7634,N_7087);
or U9130 (N_9130,N_7033,N_7355);
or U9131 (N_9131,N_6583,N_6188);
and U9132 (N_9132,N_6163,N_6201);
or U9133 (N_9133,N_6589,N_7475);
and U9134 (N_9134,N_6787,N_6224);
nand U9135 (N_9135,N_7489,N_6586);
nand U9136 (N_9136,N_7164,N_6154);
or U9137 (N_9137,N_7094,N_7674);
xor U9138 (N_9138,N_6186,N_7837);
and U9139 (N_9139,N_6658,N_7175);
nor U9140 (N_9140,N_6016,N_6705);
or U9141 (N_9141,N_6486,N_7672);
nor U9142 (N_9142,N_6576,N_6547);
or U9143 (N_9143,N_7930,N_6668);
and U9144 (N_9144,N_6281,N_6057);
or U9145 (N_9145,N_7462,N_6029);
or U9146 (N_9146,N_7791,N_7309);
xnor U9147 (N_9147,N_6423,N_7536);
or U9148 (N_9148,N_7021,N_6258);
nor U9149 (N_9149,N_6485,N_6741);
and U9150 (N_9150,N_6080,N_7616);
and U9151 (N_9151,N_6139,N_6178);
xor U9152 (N_9152,N_6276,N_7630);
nor U9153 (N_9153,N_6772,N_7460);
and U9154 (N_9154,N_6815,N_7384);
or U9155 (N_9155,N_7526,N_7512);
and U9156 (N_9156,N_7087,N_6678);
nand U9157 (N_9157,N_6097,N_6769);
xnor U9158 (N_9158,N_6345,N_7825);
nand U9159 (N_9159,N_6067,N_7527);
and U9160 (N_9160,N_7486,N_6736);
xnor U9161 (N_9161,N_7544,N_6966);
or U9162 (N_9162,N_6725,N_6322);
nand U9163 (N_9163,N_7764,N_6757);
nor U9164 (N_9164,N_6621,N_7578);
nand U9165 (N_9165,N_6584,N_7380);
and U9166 (N_9166,N_7306,N_7800);
or U9167 (N_9167,N_7339,N_7286);
and U9168 (N_9168,N_7707,N_7826);
nor U9169 (N_9169,N_6936,N_6717);
xor U9170 (N_9170,N_6324,N_6259);
or U9171 (N_9171,N_7325,N_7083);
nand U9172 (N_9172,N_6764,N_7898);
and U9173 (N_9173,N_7181,N_7364);
and U9174 (N_9174,N_7763,N_7232);
nand U9175 (N_9175,N_7280,N_6600);
or U9176 (N_9176,N_6924,N_6108);
or U9177 (N_9177,N_7888,N_7355);
xnor U9178 (N_9178,N_7734,N_6398);
or U9179 (N_9179,N_7141,N_7224);
or U9180 (N_9180,N_6423,N_6224);
and U9181 (N_9181,N_6173,N_7246);
and U9182 (N_9182,N_6882,N_7625);
nand U9183 (N_9183,N_7821,N_7338);
xnor U9184 (N_9184,N_6703,N_7696);
xnor U9185 (N_9185,N_7671,N_7646);
nand U9186 (N_9186,N_6539,N_7001);
nand U9187 (N_9187,N_6340,N_7528);
xor U9188 (N_9188,N_6182,N_7357);
or U9189 (N_9189,N_7866,N_6541);
or U9190 (N_9190,N_7730,N_7179);
or U9191 (N_9191,N_6861,N_7896);
or U9192 (N_9192,N_6661,N_6142);
nand U9193 (N_9193,N_7819,N_7002);
and U9194 (N_9194,N_6322,N_6437);
nor U9195 (N_9195,N_6664,N_7139);
nor U9196 (N_9196,N_6654,N_6528);
xnor U9197 (N_9197,N_7634,N_7374);
and U9198 (N_9198,N_7337,N_6995);
nor U9199 (N_9199,N_7324,N_6921);
nor U9200 (N_9200,N_6217,N_7003);
xnor U9201 (N_9201,N_6435,N_7615);
or U9202 (N_9202,N_7929,N_7530);
or U9203 (N_9203,N_6453,N_7169);
or U9204 (N_9204,N_6089,N_7483);
and U9205 (N_9205,N_7458,N_7597);
xnor U9206 (N_9206,N_6009,N_6270);
nand U9207 (N_9207,N_6625,N_6652);
nand U9208 (N_9208,N_7996,N_7505);
xor U9209 (N_9209,N_7226,N_7798);
nand U9210 (N_9210,N_6074,N_7863);
nor U9211 (N_9211,N_6921,N_7023);
and U9212 (N_9212,N_7966,N_6033);
nand U9213 (N_9213,N_7368,N_7237);
and U9214 (N_9214,N_7536,N_6201);
xnor U9215 (N_9215,N_7135,N_6638);
nand U9216 (N_9216,N_6257,N_6274);
nand U9217 (N_9217,N_6159,N_7793);
xnor U9218 (N_9218,N_7517,N_7590);
nor U9219 (N_9219,N_7166,N_6293);
xnor U9220 (N_9220,N_6106,N_6972);
and U9221 (N_9221,N_6666,N_7161);
nand U9222 (N_9222,N_7097,N_6407);
and U9223 (N_9223,N_7144,N_6656);
and U9224 (N_9224,N_6126,N_7082);
and U9225 (N_9225,N_6164,N_6971);
nor U9226 (N_9226,N_7392,N_7710);
nor U9227 (N_9227,N_6798,N_7799);
or U9228 (N_9228,N_6215,N_7864);
and U9229 (N_9229,N_7168,N_6865);
nand U9230 (N_9230,N_7345,N_6965);
and U9231 (N_9231,N_7209,N_7567);
nor U9232 (N_9232,N_7140,N_6516);
nor U9233 (N_9233,N_7475,N_6356);
nand U9234 (N_9234,N_7145,N_6569);
nand U9235 (N_9235,N_6683,N_7771);
and U9236 (N_9236,N_6600,N_7024);
nand U9237 (N_9237,N_7147,N_6355);
or U9238 (N_9238,N_6417,N_7078);
nor U9239 (N_9239,N_6635,N_7118);
nor U9240 (N_9240,N_6181,N_7236);
xnor U9241 (N_9241,N_7284,N_6695);
nor U9242 (N_9242,N_7952,N_6625);
or U9243 (N_9243,N_6004,N_7611);
or U9244 (N_9244,N_7242,N_6241);
and U9245 (N_9245,N_6917,N_7444);
nand U9246 (N_9246,N_7794,N_6991);
nand U9247 (N_9247,N_6778,N_6026);
and U9248 (N_9248,N_7840,N_6230);
nor U9249 (N_9249,N_7990,N_7723);
and U9250 (N_9250,N_7475,N_7628);
xor U9251 (N_9251,N_7046,N_6379);
xor U9252 (N_9252,N_7999,N_7393);
xor U9253 (N_9253,N_7285,N_6751);
nand U9254 (N_9254,N_7275,N_7500);
xnor U9255 (N_9255,N_7501,N_6098);
nor U9256 (N_9256,N_7121,N_7441);
or U9257 (N_9257,N_6034,N_6569);
or U9258 (N_9258,N_7099,N_6812);
or U9259 (N_9259,N_7269,N_7044);
nand U9260 (N_9260,N_7512,N_7153);
and U9261 (N_9261,N_7525,N_6413);
xnor U9262 (N_9262,N_7668,N_6403);
and U9263 (N_9263,N_6322,N_7654);
or U9264 (N_9264,N_6611,N_7538);
nand U9265 (N_9265,N_7011,N_7444);
nand U9266 (N_9266,N_6513,N_6366);
or U9267 (N_9267,N_7810,N_6793);
or U9268 (N_9268,N_7516,N_6011);
nand U9269 (N_9269,N_7788,N_6070);
xor U9270 (N_9270,N_7981,N_6491);
xor U9271 (N_9271,N_6331,N_7286);
nand U9272 (N_9272,N_7940,N_7103);
nor U9273 (N_9273,N_6302,N_7632);
nand U9274 (N_9274,N_7493,N_6653);
or U9275 (N_9275,N_6176,N_6339);
or U9276 (N_9276,N_7540,N_6089);
nor U9277 (N_9277,N_6265,N_6951);
and U9278 (N_9278,N_7909,N_6510);
xor U9279 (N_9279,N_6331,N_6965);
nor U9280 (N_9280,N_6379,N_7849);
xnor U9281 (N_9281,N_6806,N_7999);
nand U9282 (N_9282,N_7089,N_6088);
xnor U9283 (N_9283,N_6678,N_7958);
and U9284 (N_9284,N_7097,N_7502);
xor U9285 (N_9285,N_7017,N_6811);
or U9286 (N_9286,N_6818,N_7809);
and U9287 (N_9287,N_6626,N_6469);
xnor U9288 (N_9288,N_7184,N_7490);
or U9289 (N_9289,N_6776,N_6926);
and U9290 (N_9290,N_6543,N_7234);
nand U9291 (N_9291,N_6561,N_6707);
nor U9292 (N_9292,N_6536,N_6540);
or U9293 (N_9293,N_7176,N_7791);
nor U9294 (N_9294,N_7408,N_7215);
nor U9295 (N_9295,N_6961,N_7577);
or U9296 (N_9296,N_6424,N_7536);
or U9297 (N_9297,N_7641,N_6230);
nand U9298 (N_9298,N_7755,N_6665);
xnor U9299 (N_9299,N_7295,N_7694);
or U9300 (N_9300,N_7222,N_6561);
or U9301 (N_9301,N_7313,N_7796);
nand U9302 (N_9302,N_6469,N_6453);
nor U9303 (N_9303,N_6979,N_6166);
or U9304 (N_9304,N_7854,N_7532);
and U9305 (N_9305,N_6574,N_7762);
xnor U9306 (N_9306,N_6104,N_7042);
and U9307 (N_9307,N_6005,N_7771);
xor U9308 (N_9308,N_6352,N_7128);
xnor U9309 (N_9309,N_7160,N_7295);
nor U9310 (N_9310,N_6399,N_6583);
and U9311 (N_9311,N_6095,N_6102);
xnor U9312 (N_9312,N_6571,N_6320);
nor U9313 (N_9313,N_7569,N_6273);
or U9314 (N_9314,N_7835,N_6783);
nand U9315 (N_9315,N_7200,N_6484);
nand U9316 (N_9316,N_7940,N_7213);
and U9317 (N_9317,N_6965,N_7845);
nand U9318 (N_9318,N_7576,N_6312);
xor U9319 (N_9319,N_7404,N_6287);
nand U9320 (N_9320,N_7080,N_7876);
nand U9321 (N_9321,N_6461,N_6484);
xnor U9322 (N_9322,N_7780,N_6914);
xnor U9323 (N_9323,N_7374,N_6030);
or U9324 (N_9324,N_6967,N_7990);
or U9325 (N_9325,N_6307,N_6916);
nand U9326 (N_9326,N_7953,N_7722);
and U9327 (N_9327,N_7386,N_7739);
nand U9328 (N_9328,N_6531,N_7081);
nor U9329 (N_9329,N_7805,N_6117);
or U9330 (N_9330,N_7310,N_6534);
nand U9331 (N_9331,N_6902,N_6485);
nand U9332 (N_9332,N_6213,N_7926);
xnor U9333 (N_9333,N_7404,N_7460);
nor U9334 (N_9334,N_7297,N_7509);
or U9335 (N_9335,N_6952,N_6114);
or U9336 (N_9336,N_7184,N_6587);
or U9337 (N_9337,N_7214,N_7926);
nor U9338 (N_9338,N_6274,N_6599);
nor U9339 (N_9339,N_6715,N_6062);
or U9340 (N_9340,N_6019,N_6268);
nor U9341 (N_9341,N_7207,N_6193);
nand U9342 (N_9342,N_6264,N_6520);
nand U9343 (N_9343,N_7748,N_7960);
nand U9344 (N_9344,N_6361,N_6259);
nand U9345 (N_9345,N_6913,N_7479);
xor U9346 (N_9346,N_7756,N_7595);
and U9347 (N_9347,N_7146,N_7069);
nor U9348 (N_9348,N_6737,N_6604);
and U9349 (N_9349,N_7593,N_6110);
nor U9350 (N_9350,N_6234,N_6288);
nand U9351 (N_9351,N_7204,N_7018);
or U9352 (N_9352,N_7989,N_6030);
or U9353 (N_9353,N_6080,N_7541);
or U9354 (N_9354,N_6927,N_6609);
xnor U9355 (N_9355,N_6837,N_7642);
xor U9356 (N_9356,N_6241,N_6713);
nor U9357 (N_9357,N_7865,N_7170);
nand U9358 (N_9358,N_7609,N_7989);
nand U9359 (N_9359,N_6200,N_7028);
nor U9360 (N_9360,N_7128,N_6609);
and U9361 (N_9361,N_7477,N_7888);
and U9362 (N_9362,N_7129,N_7743);
xor U9363 (N_9363,N_6707,N_6119);
xor U9364 (N_9364,N_7687,N_7206);
or U9365 (N_9365,N_7600,N_6069);
or U9366 (N_9366,N_7849,N_6952);
and U9367 (N_9367,N_7259,N_6839);
nor U9368 (N_9368,N_6193,N_6752);
nor U9369 (N_9369,N_6320,N_7886);
or U9370 (N_9370,N_7101,N_7641);
or U9371 (N_9371,N_6135,N_7472);
or U9372 (N_9372,N_7026,N_6215);
or U9373 (N_9373,N_6193,N_7390);
nand U9374 (N_9374,N_6581,N_6806);
xnor U9375 (N_9375,N_7001,N_6604);
or U9376 (N_9376,N_7770,N_6723);
and U9377 (N_9377,N_7771,N_6163);
nand U9378 (N_9378,N_6835,N_7968);
or U9379 (N_9379,N_6033,N_6695);
xnor U9380 (N_9380,N_6685,N_6497);
or U9381 (N_9381,N_7720,N_6534);
or U9382 (N_9382,N_6658,N_6336);
nand U9383 (N_9383,N_7695,N_6838);
and U9384 (N_9384,N_6668,N_6236);
xnor U9385 (N_9385,N_6442,N_6103);
nand U9386 (N_9386,N_7694,N_6820);
xnor U9387 (N_9387,N_6519,N_7773);
and U9388 (N_9388,N_6053,N_6354);
or U9389 (N_9389,N_7781,N_6849);
nor U9390 (N_9390,N_7642,N_6318);
xor U9391 (N_9391,N_6890,N_7138);
or U9392 (N_9392,N_7009,N_6033);
xor U9393 (N_9393,N_6943,N_7782);
nor U9394 (N_9394,N_6701,N_7698);
and U9395 (N_9395,N_7497,N_6621);
nand U9396 (N_9396,N_7474,N_7935);
and U9397 (N_9397,N_6998,N_6041);
nor U9398 (N_9398,N_6727,N_7511);
xnor U9399 (N_9399,N_7754,N_7336);
nand U9400 (N_9400,N_7245,N_6141);
nor U9401 (N_9401,N_7568,N_7254);
and U9402 (N_9402,N_6743,N_6801);
xnor U9403 (N_9403,N_7721,N_7865);
and U9404 (N_9404,N_6507,N_6012);
and U9405 (N_9405,N_7641,N_7442);
xnor U9406 (N_9406,N_6785,N_7740);
xor U9407 (N_9407,N_6222,N_6802);
and U9408 (N_9408,N_7879,N_6092);
or U9409 (N_9409,N_6235,N_7407);
xnor U9410 (N_9410,N_6830,N_7883);
and U9411 (N_9411,N_7548,N_6434);
and U9412 (N_9412,N_6996,N_7566);
xor U9413 (N_9413,N_6624,N_7439);
nand U9414 (N_9414,N_7543,N_6589);
or U9415 (N_9415,N_6859,N_6629);
and U9416 (N_9416,N_6534,N_6905);
nor U9417 (N_9417,N_7452,N_6125);
nand U9418 (N_9418,N_7382,N_6124);
xor U9419 (N_9419,N_6939,N_7515);
xor U9420 (N_9420,N_6081,N_7428);
and U9421 (N_9421,N_7235,N_6238);
nand U9422 (N_9422,N_6510,N_7391);
and U9423 (N_9423,N_6153,N_6018);
and U9424 (N_9424,N_6530,N_6342);
or U9425 (N_9425,N_6819,N_6517);
and U9426 (N_9426,N_6765,N_6783);
xor U9427 (N_9427,N_7217,N_6062);
and U9428 (N_9428,N_6702,N_7900);
or U9429 (N_9429,N_7588,N_6293);
nor U9430 (N_9430,N_6401,N_6669);
or U9431 (N_9431,N_7784,N_6115);
or U9432 (N_9432,N_6967,N_7496);
or U9433 (N_9433,N_6172,N_7520);
xor U9434 (N_9434,N_7948,N_6389);
and U9435 (N_9435,N_7973,N_7955);
nor U9436 (N_9436,N_7764,N_7253);
nor U9437 (N_9437,N_7278,N_7944);
and U9438 (N_9438,N_7856,N_6956);
nand U9439 (N_9439,N_6787,N_6293);
or U9440 (N_9440,N_6941,N_6834);
nor U9441 (N_9441,N_7191,N_6027);
xnor U9442 (N_9442,N_6957,N_6127);
and U9443 (N_9443,N_7584,N_6582);
nand U9444 (N_9444,N_7263,N_6699);
nor U9445 (N_9445,N_6152,N_7569);
or U9446 (N_9446,N_7647,N_7420);
xnor U9447 (N_9447,N_6762,N_7635);
and U9448 (N_9448,N_6764,N_7360);
xnor U9449 (N_9449,N_6372,N_6544);
and U9450 (N_9450,N_6510,N_7653);
or U9451 (N_9451,N_7022,N_7892);
nor U9452 (N_9452,N_6845,N_6387);
xor U9453 (N_9453,N_7281,N_6158);
nand U9454 (N_9454,N_7148,N_6902);
nand U9455 (N_9455,N_6925,N_7332);
nor U9456 (N_9456,N_7319,N_7539);
or U9457 (N_9457,N_7491,N_7508);
and U9458 (N_9458,N_7743,N_7371);
nor U9459 (N_9459,N_6421,N_7606);
or U9460 (N_9460,N_6114,N_6247);
xnor U9461 (N_9461,N_6527,N_6883);
nand U9462 (N_9462,N_6363,N_7178);
or U9463 (N_9463,N_7843,N_7975);
or U9464 (N_9464,N_6723,N_6426);
and U9465 (N_9465,N_7934,N_6042);
or U9466 (N_9466,N_7440,N_7155);
nor U9467 (N_9467,N_6067,N_6326);
xnor U9468 (N_9468,N_6004,N_6055);
nor U9469 (N_9469,N_6201,N_7033);
and U9470 (N_9470,N_6886,N_6783);
xnor U9471 (N_9471,N_6556,N_6294);
nand U9472 (N_9472,N_6608,N_7722);
nand U9473 (N_9473,N_7155,N_7472);
and U9474 (N_9474,N_6136,N_6014);
and U9475 (N_9475,N_7538,N_7432);
nand U9476 (N_9476,N_6041,N_7659);
nand U9477 (N_9477,N_7231,N_6512);
or U9478 (N_9478,N_6289,N_6816);
or U9479 (N_9479,N_6575,N_6951);
and U9480 (N_9480,N_7070,N_6118);
nor U9481 (N_9481,N_6025,N_6919);
nor U9482 (N_9482,N_7114,N_6614);
xnor U9483 (N_9483,N_7668,N_7490);
nor U9484 (N_9484,N_7490,N_7604);
xnor U9485 (N_9485,N_7945,N_6238);
or U9486 (N_9486,N_6749,N_7230);
or U9487 (N_9487,N_6307,N_7959);
nor U9488 (N_9488,N_7207,N_6091);
and U9489 (N_9489,N_6708,N_6879);
and U9490 (N_9490,N_7655,N_6600);
and U9491 (N_9491,N_7458,N_7104);
nand U9492 (N_9492,N_6814,N_7895);
xnor U9493 (N_9493,N_7519,N_6120);
nor U9494 (N_9494,N_7483,N_7590);
nor U9495 (N_9495,N_7401,N_6239);
xnor U9496 (N_9496,N_7033,N_7571);
xor U9497 (N_9497,N_7255,N_7582);
xnor U9498 (N_9498,N_6789,N_6051);
and U9499 (N_9499,N_7625,N_7258);
nand U9500 (N_9500,N_7098,N_6616);
and U9501 (N_9501,N_7194,N_7542);
and U9502 (N_9502,N_6963,N_7055);
nor U9503 (N_9503,N_6515,N_7138);
xnor U9504 (N_9504,N_6888,N_7228);
nand U9505 (N_9505,N_7729,N_7789);
and U9506 (N_9506,N_7100,N_6671);
xnor U9507 (N_9507,N_6940,N_7049);
nor U9508 (N_9508,N_7228,N_6877);
or U9509 (N_9509,N_7940,N_7142);
or U9510 (N_9510,N_7568,N_7410);
or U9511 (N_9511,N_7353,N_6297);
or U9512 (N_9512,N_7764,N_7901);
xnor U9513 (N_9513,N_6916,N_7462);
nand U9514 (N_9514,N_7596,N_7063);
nor U9515 (N_9515,N_7364,N_7723);
nand U9516 (N_9516,N_7292,N_6229);
and U9517 (N_9517,N_6333,N_7681);
xor U9518 (N_9518,N_6619,N_7782);
nor U9519 (N_9519,N_6218,N_6801);
xnor U9520 (N_9520,N_7215,N_7497);
and U9521 (N_9521,N_7222,N_6289);
nor U9522 (N_9522,N_7735,N_7754);
nor U9523 (N_9523,N_7569,N_6631);
nand U9524 (N_9524,N_7794,N_6839);
and U9525 (N_9525,N_6200,N_6901);
and U9526 (N_9526,N_7401,N_6805);
xnor U9527 (N_9527,N_6677,N_7132);
xor U9528 (N_9528,N_6138,N_6906);
xnor U9529 (N_9529,N_7055,N_7858);
or U9530 (N_9530,N_6393,N_6655);
or U9531 (N_9531,N_6657,N_6904);
or U9532 (N_9532,N_7775,N_7928);
and U9533 (N_9533,N_6371,N_6992);
or U9534 (N_9534,N_7118,N_6780);
nor U9535 (N_9535,N_6068,N_6615);
or U9536 (N_9536,N_6033,N_6578);
and U9537 (N_9537,N_6519,N_7404);
xor U9538 (N_9538,N_6885,N_7628);
nand U9539 (N_9539,N_6465,N_7626);
nor U9540 (N_9540,N_7744,N_6082);
and U9541 (N_9541,N_7349,N_7357);
nor U9542 (N_9542,N_6709,N_6701);
xnor U9543 (N_9543,N_7214,N_7198);
nor U9544 (N_9544,N_7029,N_6035);
nor U9545 (N_9545,N_7512,N_6054);
nand U9546 (N_9546,N_6858,N_6974);
and U9547 (N_9547,N_7538,N_7009);
nor U9548 (N_9548,N_7573,N_7098);
or U9549 (N_9549,N_7191,N_6536);
and U9550 (N_9550,N_6217,N_6510);
nand U9551 (N_9551,N_6686,N_6402);
or U9552 (N_9552,N_6474,N_7264);
xor U9553 (N_9553,N_6354,N_6805);
xor U9554 (N_9554,N_7309,N_6862);
nor U9555 (N_9555,N_7240,N_7600);
nor U9556 (N_9556,N_7182,N_7742);
xor U9557 (N_9557,N_6620,N_7745);
nand U9558 (N_9558,N_6696,N_7951);
and U9559 (N_9559,N_7087,N_7418);
xnor U9560 (N_9560,N_7177,N_7037);
xnor U9561 (N_9561,N_6102,N_6916);
and U9562 (N_9562,N_7582,N_6561);
or U9563 (N_9563,N_7591,N_7764);
nor U9564 (N_9564,N_6536,N_6199);
xnor U9565 (N_9565,N_7680,N_6710);
and U9566 (N_9566,N_7336,N_7939);
nor U9567 (N_9567,N_7048,N_7398);
xor U9568 (N_9568,N_6611,N_7485);
nand U9569 (N_9569,N_6867,N_7824);
xor U9570 (N_9570,N_7893,N_6223);
nor U9571 (N_9571,N_7144,N_6163);
nor U9572 (N_9572,N_7482,N_7514);
xnor U9573 (N_9573,N_7275,N_6624);
and U9574 (N_9574,N_7139,N_6794);
nand U9575 (N_9575,N_7786,N_7115);
nor U9576 (N_9576,N_7440,N_7255);
nand U9577 (N_9577,N_7105,N_7805);
nand U9578 (N_9578,N_7256,N_7460);
and U9579 (N_9579,N_6058,N_6360);
or U9580 (N_9580,N_7516,N_6825);
and U9581 (N_9581,N_7229,N_6923);
xor U9582 (N_9582,N_6459,N_7754);
or U9583 (N_9583,N_7929,N_7979);
xor U9584 (N_9584,N_6773,N_7307);
nand U9585 (N_9585,N_6431,N_7742);
or U9586 (N_9586,N_7584,N_7529);
nand U9587 (N_9587,N_6987,N_7967);
nand U9588 (N_9588,N_6442,N_7177);
and U9589 (N_9589,N_7720,N_7180);
and U9590 (N_9590,N_6816,N_7098);
nand U9591 (N_9591,N_6006,N_6149);
nor U9592 (N_9592,N_6406,N_6445);
or U9593 (N_9593,N_7204,N_7899);
or U9594 (N_9594,N_6675,N_6807);
nor U9595 (N_9595,N_7189,N_6818);
xnor U9596 (N_9596,N_6512,N_6673);
nor U9597 (N_9597,N_6652,N_7989);
and U9598 (N_9598,N_6761,N_7619);
nor U9599 (N_9599,N_7493,N_7276);
and U9600 (N_9600,N_7137,N_7113);
nand U9601 (N_9601,N_7801,N_6090);
and U9602 (N_9602,N_6064,N_6548);
nand U9603 (N_9603,N_6425,N_6331);
nand U9604 (N_9604,N_7940,N_6301);
xor U9605 (N_9605,N_7478,N_7007);
xnor U9606 (N_9606,N_7686,N_6873);
and U9607 (N_9607,N_6283,N_6338);
xnor U9608 (N_9608,N_6748,N_7080);
xor U9609 (N_9609,N_6334,N_6221);
or U9610 (N_9610,N_6406,N_7753);
or U9611 (N_9611,N_7928,N_6858);
xnor U9612 (N_9612,N_7674,N_6898);
nand U9613 (N_9613,N_7502,N_7439);
or U9614 (N_9614,N_7570,N_7184);
xnor U9615 (N_9615,N_6290,N_7932);
and U9616 (N_9616,N_6536,N_6419);
and U9617 (N_9617,N_7678,N_6504);
xor U9618 (N_9618,N_7977,N_7301);
xor U9619 (N_9619,N_6588,N_7067);
or U9620 (N_9620,N_7303,N_6114);
nor U9621 (N_9621,N_7464,N_6162);
xor U9622 (N_9622,N_6180,N_6291);
or U9623 (N_9623,N_6511,N_7255);
and U9624 (N_9624,N_6777,N_6613);
or U9625 (N_9625,N_6850,N_6453);
and U9626 (N_9626,N_6247,N_6277);
nor U9627 (N_9627,N_6988,N_7884);
nand U9628 (N_9628,N_7583,N_7234);
or U9629 (N_9629,N_7431,N_6592);
nor U9630 (N_9630,N_6818,N_6289);
nand U9631 (N_9631,N_7864,N_6610);
xnor U9632 (N_9632,N_7251,N_6818);
nor U9633 (N_9633,N_7886,N_6566);
or U9634 (N_9634,N_7952,N_7217);
and U9635 (N_9635,N_6331,N_6601);
xnor U9636 (N_9636,N_7616,N_7677);
and U9637 (N_9637,N_6486,N_6349);
nand U9638 (N_9638,N_6321,N_7440);
or U9639 (N_9639,N_6079,N_6852);
xor U9640 (N_9640,N_7488,N_6223);
or U9641 (N_9641,N_6340,N_6436);
nand U9642 (N_9642,N_6600,N_6374);
xor U9643 (N_9643,N_7206,N_6866);
and U9644 (N_9644,N_6901,N_6071);
nand U9645 (N_9645,N_7246,N_6710);
or U9646 (N_9646,N_6970,N_6205);
nor U9647 (N_9647,N_7279,N_7453);
nand U9648 (N_9648,N_6816,N_7652);
xor U9649 (N_9649,N_7461,N_6525);
or U9650 (N_9650,N_7429,N_7300);
xor U9651 (N_9651,N_6879,N_6755);
nor U9652 (N_9652,N_7943,N_6162);
and U9653 (N_9653,N_7306,N_7330);
xnor U9654 (N_9654,N_7851,N_6728);
and U9655 (N_9655,N_7886,N_7407);
xnor U9656 (N_9656,N_7505,N_7001);
and U9657 (N_9657,N_6971,N_7490);
nor U9658 (N_9658,N_6207,N_6308);
or U9659 (N_9659,N_7573,N_7185);
xor U9660 (N_9660,N_6620,N_7446);
nand U9661 (N_9661,N_6605,N_7994);
or U9662 (N_9662,N_6561,N_6306);
nand U9663 (N_9663,N_6320,N_7832);
and U9664 (N_9664,N_7562,N_6315);
nand U9665 (N_9665,N_6026,N_7977);
nor U9666 (N_9666,N_7596,N_7317);
nand U9667 (N_9667,N_6050,N_6081);
xor U9668 (N_9668,N_6920,N_6473);
or U9669 (N_9669,N_6412,N_6534);
nand U9670 (N_9670,N_6690,N_6460);
xor U9671 (N_9671,N_6255,N_6115);
or U9672 (N_9672,N_7966,N_6682);
nor U9673 (N_9673,N_7216,N_7732);
nor U9674 (N_9674,N_7576,N_7571);
nor U9675 (N_9675,N_6721,N_6113);
nand U9676 (N_9676,N_6236,N_6636);
nand U9677 (N_9677,N_7866,N_7676);
xnor U9678 (N_9678,N_7435,N_7020);
or U9679 (N_9679,N_7544,N_6446);
and U9680 (N_9680,N_7492,N_6031);
nand U9681 (N_9681,N_6351,N_6710);
and U9682 (N_9682,N_6340,N_6932);
nand U9683 (N_9683,N_7262,N_7029);
or U9684 (N_9684,N_6008,N_6423);
nand U9685 (N_9685,N_7300,N_6618);
and U9686 (N_9686,N_6763,N_6703);
nor U9687 (N_9687,N_6683,N_7685);
nor U9688 (N_9688,N_6073,N_6961);
nand U9689 (N_9689,N_6189,N_6342);
nand U9690 (N_9690,N_6409,N_6434);
and U9691 (N_9691,N_6632,N_7811);
and U9692 (N_9692,N_6809,N_7171);
nor U9693 (N_9693,N_7354,N_6385);
nor U9694 (N_9694,N_6499,N_7306);
xnor U9695 (N_9695,N_7909,N_6177);
nor U9696 (N_9696,N_7264,N_7815);
and U9697 (N_9697,N_7312,N_7641);
nand U9698 (N_9698,N_7695,N_7205);
nor U9699 (N_9699,N_6922,N_6007);
nor U9700 (N_9700,N_6832,N_7409);
or U9701 (N_9701,N_6475,N_6164);
nand U9702 (N_9702,N_6522,N_7774);
or U9703 (N_9703,N_6355,N_6492);
nor U9704 (N_9704,N_6578,N_7647);
nand U9705 (N_9705,N_6777,N_7379);
or U9706 (N_9706,N_7993,N_6272);
nand U9707 (N_9707,N_7298,N_7538);
nand U9708 (N_9708,N_7972,N_6499);
xor U9709 (N_9709,N_7318,N_7299);
xnor U9710 (N_9710,N_6252,N_7061);
and U9711 (N_9711,N_7618,N_7839);
or U9712 (N_9712,N_7138,N_6067);
or U9713 (N_9713,N_7109,N_7600);
nand U9714 (N_9714,N_6838,N_6559);
or U9715 (N_9715,N_7544,N_6709);
nand U9716 (N_9716,N_7926,N_6582);
nand U9717 (N_9717,N_7787,N_6700);
nand U9718 (N_9718,N_6131,N_6150);
nand U9719 (N_9719,N_7435,N_7170);
xor U9720 (N_9720,N_7248,N_7029);
nor U9721 (N_9721,N_7731,N_6365);
and U9722 (N_9722,N_7302,N_6283);
nand U9723 (N_9723,N_7753,N_7548);
nor U9724 (N_9724,N_6805,N_7201);
nand U9725 (N_9725,N_7377,N_6928);
nand U9726 (N_9726,N_6381,N_7946);
and U9727 (N_9727,N_7372,N_6272);
nand U9728 (N_9728,N_6382,N_6697);
or U9729 (N_9729,N_6897,N_6098);
xor U9730 (N_9730,N_7291,N_7457);
xor U9731 (N_9731,N_6633,N_7001);
or U9732 (N_9732,N_6374,N_7926);
nor U9733 (N_9733,N_7434,N_7612);
nor U9734 (N_9734,N_6571,N_6052);
and U9735 (N_9735,N_6976,N_6124);
and U9736 (N_9736,N_6294,N_7875);
nor U9737 (N_9737,N_6016,N_7240);
xor U9738 (N_9738,N_6712,N_6324);
nand U9739 (N_9739,N_6501,N_6867);
nand U9740 (N_9740,N_6369,N_6378);
xor U9741 (N_9741,N_6639,N_7520);
or U9742 (N_9742,N_7236,N_6680);
or U9743 (N_9743,N_6636,N_7370);
and U9744 (N_9744,N_7687,N_7396);
or U9745 (N_9745,N_6814,N_7730);
xnor U9746 (N_9746,N_6217,N_6243);
nand U9747 (N_9747,N_7532,N_7756);
nor U9748 (N_9748,N_7626,N_6584);
nor U9749 (N_9749,N_7024,N_7998);
xnor U9750 (N_9750,N_6657,N_6155);
or U9751 (N_9751,N_6967,N_7627);
and U9752 (N_9752,N_7921,N_7678);
nor U9753 (N_9753,N_6874,N_7838);
nand U9754 (N_9754,N_7473,N_6697);
nand U9755 (N_9755,N_6607,N_7684);
nand U9756 (N_9756,N_6572,N_6009);
nand U9757 (N_9757,N_6881,N_7729);
xnor U9758 (N_9758,N_7748,N_7525);
nand U9759 (N_9759,N_6584,N_7099);
nor U9760 (N_9760,N_6853,N_7970);
nand U9761 (N_9761,N_7572,N_6238);
xor U9762 (N_9762,N_7444,N_7425);
nor U9763 (N_9763,N_7536,N_6281);
or U9764 (N_9764,N_7665,N_6070);
xnor U9765 (N_9765,N_6114,N_7486);
nand U9766 (N_9766,N_6716,N_6543);
and U9767 (N_9767,N_7652,N_7616);
xor U9768 (N_9768,N_7173,N_7483);
or U9769 (N_9769,N_6441,N_6350);
or U9770 (N_9770,N_6436,N_6613);
and U9771 (N_9771,N_6410,N_7520);
and U9772 (N_9772,N_7534,N_7536);
or U9773 (N_9773,N_6633,N_6101);
nand U9774 (N_9774,N_7684,N_7551);
nor U9775 (N_9775,N_7867,N_6360);
nand U9776 (N_9776,N_6194,N_7694);
nor U9777 (N_9777,N_7993,N_6654);
xor U9778 (N_9778,N_6146,N_7040);
nor U9779 (N_9779,N_7378,N_7736);
xnor U9780 (N_9780,N_7742,N_6475);
nor U9781 (N_9781,N_7047,N_6473);
nand U9782 (N_9782,N_7506,N_6017);
nor U9783 (N_9783,N_6881,N_7300);
nand U9784 (N_9784,N_7526,N_7329);
xor U9785 (N_9785,N_7101,N_7110);
or U9786 (N_9786,N_6149,N_6113);
xnor U9787 (N_9787,N_6917,N_6827);
xor U9788 (N_9788,N_7708,N_6834);
nor U9789 (N_9789,N_7481,N_7897);
or U9790 (N_9790,N_7646,N_7889);
and U9791 (N_9791,N_6770,N_6138);
nor U9792 (N_9792,N_6813,N_6141);
and U9793 (N_9793,N_6437,N_6384);
or U9794 (N_9794,N_6148,N_7506);
or U9795 (N_9795,N_6246,N_7416);
or U9796 (N_9796,N_6200,N_6261);
nand U9797 (N_9797,N_7805,N_6847);
xnor U9798 (N_9798,N_7135,N_6956);
or U9799 (N_9799,N_7055,N_7253);
xor U9800 (N_9800,N_6173,N_6237);
or U9801 (N_9801,N_6619,N_7552);
nor U9802 (N_9802,N_6970,N_7030);
and U9803 (N_9803,N_6178,N_6106);
nor U9804 (N_9804,N_7213,N_7452);
and U9805 (N_9805,N_6012,N_7552);
nor U9806 (N_9806,N_7418,N_7326);
xnor U9807 (N_9807,N_6285,N_6252);
or U9808 (N_9808,N_6310,N_7914);
and U9809 (N_9809,N_6622,N_7679);
xor U9810 (N_9810,N_7545,N_7308);
xnor U9811 (N_9811,N_7239,N_6094);
and U9812 (N_9812,N_7777,N_6716);
or U9813 (N_9813,N_6591,N_7616);
nor U9814 (N_9814,N_7076,N_6674);
nand U9815 (N_9815,N_7531,N_6190);
nand U9816 (N_9816,N_7338,N_7630);
nor U9817 (N_9817,N_7080,N_6413);
or U9818 (N_9818,N_6064,N_6401);
nor U9819 (N_9819,N_7863,N_6183);
and U9820 (N_9820,N_6207,N_6728);
and U9821 (N_9821,N_7326,N_6415);
nand U9822 (N_9822,N_7629,N_6652);
or U9823 (N_9823,N_6246,N_7625);
and U9824 (N_9824,N_7342,N_6397);
and U9825 (N_9825,N_6911,N_7131);
or U9826 (N_9826,N_6748,N_6392);
nand U9827 (N_9827,N_7144,N_6880);
nand U9828 (N_9828,N_6761,N_6215);
nand U9829 (N_9829,N_7532,N_6033);
nor U9830 (N_9830,N_7389,N_6899);
xnor U9831 (N_9831,N_7172,N_6470);
nor U9832 (N_9832,N_7108,N_6026);
xnor U9833 (N_9833,N_7840,N_7883);
nand U9834 (N_9834,N_7996,N_6102);
or U9835 (N_9835,N_7244,N_7348);
nand U9836 (N_9836,N_7605,N_6005);
nand U9837 (N_9837,N_6405,N_6378);
nor U9838 (N_9838,N_7129,N_6018);
xor U9839 (N_9839,N_6167,N_7694);
nor U9840 (N_9840,N_7325,N_6764);
nor U9841 (N_9841,N_7983,N_6765);
xor U9842 (N_9842,N_6313,N_6025);
or U9843 (N_9843,N_7657,N_7889);
nand U9844 (N_9844,N_7649,N_7543);
or U9845 (N_9845,N_7448,N_6525);
or U9846 (N_9846,N_7256,N_6516);
xor U9847 (N_9847,N_7543,N_6017);
or U9848 (N_9848,N_7326,N_6903);
and U9849 (N_9849,N_7083,N_7144);
xnor U9850 (N_9850,N_7062,N_7611);
and U9851 (N_9851,N_7985,N_6565);
xnor U9852 (N_9852,N_6679,N_7026);
nor U9853 (N_9853,N_6174,N_6341);
nand U9854 (N_9854,N_6243,N_6787);
and U9855 (N_9855,N_7551,N_7276);
nand U9856 (N_9856,N_6767,N_6099);
or U9857 (N_9857,N_6540,N_7685);
xor U9858 (N_9858,N_7969,N_6136);
xnor U9859 (N_9859,N_6471,N_7713);
or U9860 (N_9860,N_6004,N_6495);
xnor U9861 (N_9861,N_6238,N_6421);
nor U9862 (N_9862,N_7833,N_6402);
and U9863 (N_9863,N_6975,N_6749);
nand U9864 (N_9864,N_6454,N_7767);
xnor U9865 (N_9865,N_6529,N_7105);
nand U9866 (N_9866,N_6193,N_7988);
xnor U9867 (N_9867,N_6357,N_6397);
or U9868 (N_9868,N_7742,N_7779);
xor U9869 (N_9869,N_7608,N_6988);
and U9870 (N_9870,N_7878,N_6109);
or U9871 (N_9871,N_7568,N_7975);
and U9872 (N_9872,N_6129,N_6125);
and U9873 (N_9873,N_7359,N_7864);
nand U9874 (N_9874,N_6290,N_7338);
or U9875 (N_9875,N_7556,N_7908);
or U9876 (N_9876,N_6740,N_6861);
and U9877 (N_9877,N_6645,N_7799);
nor U9878 (N_9878,N_6153,N_6785);
xor U9879 (N_9879,N_6586,N_6949);
xnor U9880 (N_9880,N_6675,N_7903);
or U9881 (N_9881,N_7410,N_6988);
xnor U9882 (N_9882,N_6307,N_6414);
nand U9883 (N_9883,N_7047,N_7250);
or U9884 (N_9884,N_7857,N_6456);
and U9885 (N_9885,N_7357,N_6230);
nor U9886 (N_9886,N_6169,N_7877);
xnor U9887 (N_9887,N_6759,N_6173);
or U9888 (N_9888,N_7963,N_6678);
xnor U9889 (N_9889,N_6535,N_7333);
and U9890 (N_9890,N_6908,N_7739);
nor U9891 (N_9891,N_6209,N_6833);
and U9892 (N_9892,N_7142,N_6657);
xor U9893 (N_9893,N_6105,N_7758);
and U9894 (N_9894,N_6343,N_6590);
and U9895 (N_9895,N_6818,N_6177);
nand U9896 (N_9896,N_6315,N_6482);
and U9897 (N_9897,N_7450,N_6911);
nand U9898 (N_9898,N_7926,N_6742);
xnor U9899 (N_9899,N_7871,N_7964);
and U9900 (N_9900,N_7734,N_6702);
or U9901 (N_9901,N_6543,N_6547);
xnor U9902 (N_9902,N_6893,N_6607);
or U9903 (N_9903,N_7441,N_6973);
or U9904 (N_9904,N_7236,N_6851);
nor U9905 (N_9905,N_6312,N_6414);
xor U9906 (N_9906,N_6658,N_7416);
xnor U9907 (N_9907,N_6086,N_6221);
and U9908 (N_9908,N_6351,N_7427);
xor U9909 (N_9909,N_6389,N_7461);
xor U9910 (N_9910,N_6893,N_7894);
nand U9911 (N_9911,N_6038,N_6748);
nor U9912 (N_9912,N_7000,N_6365);
and U9913 (N_9913,N_7192,N_6701);
or U9914 (N_9914,N_7316,N_7426);
nor U9915 (N_9915,N_6348,N_7445);
nand U9916 (N_9916,N_7237,N_6129);
xnor U9917 (N_9917,N_6274,N_7085);
xor U9918 (N_9918,N_6527,N_6216);
nor U9919 (N_9919,N_7346,N_6656);
or U9920 (N_9920,N_6442,N_7362);
xnor U9921 (N_9921,N_6162,N_6073);
or U9922 (N_9922,N_7582,N_6660);
and U9923 (N_9923,N_7490,N_7442);
xor U9924 (N_9924,N_6147,N_7966);
xnor U9925 (N_9925,N_7402,N_7629);
xor U9926 (N_9926,N_7458,N_7264);
xnor U9927 (N_9927,N_6053,N_6246);
and U9928 (N_9928,N_7734,N_7603);
xnor U9929 (N_9929,N_6465,N_7257);
and U9930 (N_9930,N_6365,N_7892);
xor U9931 (N_9931,N_7426,N_7570);
or U9932 (N_9932,N_7489,N_7144);
and U9933 (N_9933,N_6928,N_7560);
nor U9934 (N_9934,N_6029,N_7432);
nor U9935 (N_9935,N_6127,N_6702);
nand U9936 (N_9936,N_7917,N_6350);
nand U9937 (N_9937,N_6569,N_6382);
nor U9938 (N_9938,N_6950,N_7549);
nor U9939 (N_9939,N_7136,N_6724);
and U9940 (N_9940,N_6321,N_7698);
or U9941 (N_9941,N_7563,N_7280);
or U9942 (N_9942,N_7779,N_6843);
and U9943 (N_9943,N_6938,N_6172);
or U9944 (N_9944,N_7351,N_6137);
xor U9945 (N_9945,N_6204,N_6411);
xor U9946 (N_9946,N_6631,N_6517);
and U9947 (N_9947,N_7579,N_7979);
nor U9948 (N_9948,N_7949,N_6903);
xnor U9949 (N_9949,N_6958,N_7011);
nand U9950 (N_9950,N_6202,N_6710);
nand U9951 (N_9951,N_6782,N_6732);
and U9952 (N_9952,N_7298,N_7025);
or U9953 (N_9953,N_7461,N_7269);
nor U9954 (N_9954,N_7490,N_6241);
nor U9955 (N_9955,N_6645,N_7510);
nand U9956 (N_9956,N_6358,N_7634);
nor U9957 (N_9957,N_7516,N_6902);
nor U9958 (N_9958,N_6420,N_7089);
xor U9959 (N_9959,N_7482,N_6038);
and U9960 (N_9960,N_7447,N_7085);
nand U9961 (N_9961,N_7226,N_6478);
nand U9962 (N_9962,N_7109,N_6295);
nor U9963 (N_9963,N_7239,N_6446);
and U9964 (N_9964,N_7746,N_7231);
and U9965 (N_9965,N_7481,N_6665);
nor U9966 (N_9966,N_7198,N_7220);
nand U9967 (N_9967,N_6090,N_6252);
or U9968 (N_9968,N_6897,N_7187);
and U9969 (N_9969,N_7997,N_6653);
nand U9970 (N_9970,N_6237,N_7959);
nand U9971 (N_9971,N_6923,N_6018);
nor U9972 (N_9972,N_6922,N_7108);
xnor U9973 (N_9973,N_6644,N_7878);
nor U9974 (N_9974,N_6679,N_7195);
or U9975 (N_9975,N_7963,N_6355);
xnor U9976 (N_9976,N_7415,N_6139);
nor U9977 (N_9977,N_6886,N_6758);
nor U9978 (N_9978,N_6292,N_7523);
xnor U9979 (N_9979,N_6081,N_6845);
nor U9980 (N_9980,N_7475,N_7305);
nor U9981 (N_9981,N_7930,N_6533);
or U9982 (N_9982,N_7177,N_6534);
or U9983 (N_9983,N_6753,N_6470);
nand U9984 (N_9984,N_7174,N_7646);
or U9985 (N_9985,N_7807,N_6337);
xnor U9986 (N_9986,N_7552,N_7478);
nand U9987 (N_9987,N_6112,N_6589);
and U9988 (N_9988,N_7400,N_7734);
xor U9989 (N_9989,N_6521,N_7492);
or U9990 (N_9990,N_6006,N_6316);
xor U9991 (N_9991,N_7715,N_7730);
or U9992 (N_9992,N_7150,N_6633);
nand U9993 (N_9993,N_7211,N_6418);
nor U9994 (N_9994,N_7993,N_6490);
or U9995 (N_9995,N_7876,N_7991);
nand U9996 (N_9996,N_6426,N_6278);
or U9997 (N_9997,N_6250,N_7300);
and U9998 (N_9998,N_6738,N_6595);
nor U9999 (N_9999,N_7031,N_6349);
and U10000 (N_10000,N_8192,N_9890);
or U10001 (N_10001,N_8255,N_9708);
and U10002 (N_10002,N_8605,N_9823);
and U10003 (N_10003,N_9574,N_9028);
xor U10004 (N_10004,N_9042,N_8771);
and U10005 (N_10005,N_9400,N_9460);
and U10006 (N_10006,N_9669,N_8082);
nor U10007 (N_10007,N_8707,N_9936);
or U10008 (N_10008,N_9044,N_9808);
or U10009 (N_10009,N_8327,N_8176);
xor U10010 (N_10010,N_8906,N_8646);
xnor U10011 (N_10011,N_8389,N_9921);
nand U10012 (N_10012,N_8154,N_8585);
and U10013 (N_10013,N_8766,N_8991);
nor U10014 (N_10014,N_8686,N_8347);
xnor U10015 (N_10015,N_9308,N_8713);
and U10016 (N_10016,N_8699,N_8424);
xor U10017 (N_10017,N_9862,N_9147);
or U10018 (N_10018,N_9564,N_8739);
or U10019 (N_10019,N_9242,N_9052);
or U10020 (N_10020,N_9321,N_8725);
nand U10021 (N_10021,N_8899,N_8979);
and U10022 (N_10022,N_9686,N_9264);
and U10023 (N_10023,N_9408,N_8383);
xnor U10024 (N_10024,N_8369,N_8554);
nor U10025 (N_10025,N_8795,N_8103);
or U10026 (N_10026,N_9067,N_8832);
or U10027 (N_10027,N_9123,N_8698);
nor U10028 (N_10028,N_9366,N_9703);
nand U10029 (N_10029,N_8622,N_8027);
or U10030 (N_10030,N_8547,N_9826);
xnor U10031 (N_10031,N_9002,N_8782);
xnor U10032 (N_10032,N_8432,N_8590);
nand U10033 (N_10033,N_8579,N_8271);
nor U10034 (N_10034,N_9150,N_8164);
xnor U10035 (N_10035,N_9309,N_8143);
nand U10036 (N_10036,N_8484,N_8737);
xnor U10037 (N_10037,N_8138,N_8134);
or U10038 (N_10038,N_9831,N_9461);
and U10039 (N_10039,N_8475,N_8244);
or U10040 (N_10040,N_8381,N_9134);
nor U10041 (N_10041,N_8038,N_9171);
or U10042 (N_10042,N_8153,N_8180);
xnor U10043 (N_10043,N_9156,N_9879);
nand U10044 (N_10044,N_9859,N_8118);
nand U10045 (N_10045,N_8478,N_8452);
or U10046 (N_10046,N_9733,N_9177);
or U10047 (N_10047,N_8351,N_8596);
and U10048 (N_10048,N_8530,N_8524);
xor U10049 (N_10049,N_8956,N_9565);
and U10050 (N_10050,N_8696,N_9911);
nor U10051 (N_10051,N_8288,N_9806);
nor U10052 (N_10052,N_8663,N_8802);
xor U10053 (N_10053,N_9160,N_8845);
nand U10054 (N_10054,N_9683,N_9277);
or U10055 (N_10055,N_9790,N_8498);
nor U10056 (N_10056,N_8607,N_8167);
nand U10057 (N_10057,N_8592,N_8717);
or U10058 (N_10058,N_8654,N_9718);
nor U10059 (N_10059,N_9927,N_8966);
and U10060 (N_10060,N_8961,N_9902);
or U10061 (N_10061,N_9809,N_8430);
xor U10062 (N_10062,N_9172,N_8673);
nand U10063 (N_10063,N_9724,N_8029);
xnor U10064 (N_10064,N_9009,N_8629);
nand U10065 (N_10065,N_8784,N_8923);
or U10066 (N_10066,N_9899,N_8088);
nand U10067 (N_10067,N_8871,N_9851);
xor U10068 (N_10068,N_9815,N_9057);
and U10069 (N_10069,N_8512,N_9228);
xor U10070 (N_10070,N_9431,N_9021);
nand U10071 (N_10071,N_8026,N_8815);
xor U10072 (N_10072,N_8689,N_8319);
or U10073 (N_10073,N_9688,N_9577);
nor U10074 (N_10074,N_8139,N_8587);
or U10075 (N_10075,N_8178,N_8773);
or U10076 (N_10076,N_9168,N_9896);
and U10077 (N_10077,N_9015,N_9447);
or U10078 (N_10078,N_9151,N_8515);
and U10079 (N_10079,N_8848,N_9612);
and U10080 (N_10080,N_9471,N_9212);
xnor U10081 (N_10081,N_9558,N_8057);
and U10082 (N_10082,N_8039,N_9934);
nor U10083 (N_10083,N_9483,N_9265);
and U10084 (N_10084,N_9738,N_8291);
and U10085 (N_10085,N_8031,N_9492);
xnor U10086 (N_10086,N_9882,N_9763);
and U10087 (N_10087,N_9105,N_8905);
xor U10088 (N_10088,N_9217,N_8047);
nand U10089 (N_10089,N_8804,N_9922);
or U10090 (N_10090,N_8929,N_9705);
or U10091 (N_10091,N_8419,N_8358);
nor U10092 (N_10092,N_9845,N_9040);
xor U10093 (N_10093,N_8313,N_8750);
xor U10094 (N_10094,N_9909,N_8538);
xor U10095 (N_10095,N_8551,N_8330);
or U10096 (N_10096,N_9698,N_8833);
and U10097 (N_10097,N_8416,N_8667);
or U10098 (N_10098,N_9116,N_8454);
xnor U10099 (N_10099,N_9645,N_8576);
nand U10100 (N_10100,N_8772,N_9777);
or U10101 (N_10101,N_8986,N_8356);
nor U10102 (N_10102,N_8578,N_8469);
or U10103 (N_10103,N_8857,N_8916);
or U10104 (N_10104,N_9534,N_8423);
xnor U10105 (N_10105,N_9096,N_8652);
xnor U10106 (N_10106,N_9668,N_9055);
nor U10107 (N_10107,N_8458,N_9155);
nand U10108 (N_10108,N_8907,N_9465);
nor U10109 (N_10109,N_9401,N_9399);
xor U10110 (N_10110,N_8035,N_8517);
nor U10111 (N_10111,N_8609,N_9275);
nor U10112 (N_10112,N_9749,N_9521);
nand U10113 (N_10113,N_8627,N_8449);
xor U10114 (N_10114,N_9499,N_8042);
nor U10115 (N_10115,N_8893,N_9538);
xnor U10116 (N_10116,N_8163,N_8457);
and U10117 (N_10117,N_9474,N_8075);
nand U10118 (N_10118,N_9083,N_8343);
nand U10119 (N_10119,N_8593,N_8106);
or U10120 (N_10120,N_8774,N_9557);
nor U10121 (N_10121,N_9712,N_8998);
xnor U10122 (N_10122,N_9775,N_9800);
nand U10123 (N_10123,N_9149,N_9878);
xor U10124 (N_10124,N_9258,N_8670);
nand U10125 (N_10125,N_9596,N_8162);
and U10126 (N_10126,N_9964,N_8051);
and U10127 (N_10127,N_8467,N_8009);
nor U10128 (N_10128,N_9306,N_8700);
or U10129 (N_10129,N_8544,N_8217);
xnor U10130 (N_10130,N_9629,N_9000);
nand U10131 (N_10131,N_9370,N_8441);
and U10132 (N_10132,N_9433,N_9758);
nor U10133 (N_10133,N_8561,N_9295);
or U10134 (N_10134,N_8438,N_9003);
xnor U10135 (N_10135,N_8535,N_9233);
nor U10136 (N_10136,N_8024,N_8294);
or U10137 (N_10137,N_9576,N_9850);
or U10138 (N_10138,N_9273,N_8716);
or U10139 (N_10139,N_9967,N_8166);
nor U10140 (N_10140,N_8948,N_9561);
nand U10141 (N_10141,N_9439,N_8333);
nand U10142 (N_10142,N_8341,N_9945);
or U10143 (N_10143,N_8641,N_9372);
or U10144 (N_10144,N_8494,N_8897);
xnor U10145 (N_10145,N_8382,N_9840);
or U10146 (N_10146,N_8232,N_8148);
and U10147 (N_10147,N_8496,N_8006);
nand U10148 (N_10148,N_9470,N_9545);
nor U10149 (N_10149,N_9428,N_9907);
nand U10150 (N_10150,N_9174,N_9307);
nand U10151 (N_10151,N_9239,N_8242);
xor U10152 (N_10152,N_9078,N_8140);
and U10153 (N_10153,N_8599,N_9200);
xor U10154 (N_10154,N_8245,N_9898);
nor U10155 (N_10155,N_8649,N_8884);
nand U10156 (N_10156,N_9631,N_8297);
and U10157 (N_10157,N_9848,N_8243);
nand U10158 (N_10158,N_9269,N_9988);
xnor U10159 (N_10159,N_9569,N_9737);
nor U10160 (N_10160,N_9720,N_8144);
nor U10161 (N_10161,N_8964,N_9989);
nor U10162 (N_10162,N_9572,N_8756);
and U10163 (N_10163,N_9259,N_9769);
nor U10164 (N_10164,N_9503,N_8455);
or U10165 (N_10165,N_8374,N_8055);
or U10166 (N_10166,N_8635,N_8115);
and U10167 (N_10167,N_8499,N_9732);
or U10168 (N_10168,N_9245,N_8236);
xnor U10169 (N_10169,N_9880,N_8439);
nor U10170 (N_10170,N_8212,N_8099);
nor U10171 (N_10171,N_9448,N_8968);
nor U10172 (N_10172,N_8885,N_9947);
or U10173 (N_10173,N_9327,N_9743);
or U10174 (N_10174,N_8807,N_9204);
or U10175 (N_10175,N_8844,N_8643);
nor U10176 (N_10176,N_8161,N_9736);
and U10177 (N_10177,N_9184,N_8872);
xnor U10178 (N_10178,N_9490,N_8056);
nor U10179 (N_10179,N_9349,N_8693);
and U10180 (N_10180,N_9871,N_8859);
nand U10181 (N_10181,N_9870,N_9373);
and U10182 (N_10182,N_8181,N_8738);
nand U10183 (N_10183,N_9525,N_8470);
xor U10184 (N_10184,N_9729,N_9451);
and U10185 (N_10185,N_9793,N_8918);
nor U10186 (N_10186,N_9092,N_8307);
or U10187 (N_10187,N_8710,N_8227);
or U10188 (N_10188,N_8728,N_8480);
nand U10189 (N_10189,N_9665,N_8486);
or U10190 (N_10190,N_8724,N_8669);
nor U10191 (N_10191,N_8894,N_9037);
nand U10192 (N_10192,N_9001,N_9908);
nor U10193 (N_10193,N_8363,N_9118);
and U10194 (N_10194,N_8919,N_8091);
and U10195 (N_10195,N_9225,N_9663);
and U10196 (N_10196,N_9106,N_9214);
or U10197 (N_10197,N_9832,N_9584);
nand U10198 (N_10198,N_9122,N_9056);
xnor U10199 (N_10199,N_9954,N_9328);
or U10200 (N_10200,N_9925,N_9025);
or U10201 (N_10201,N_9613,N_9262);
nand U10202 (N_10202,N_8934,N_8746);
xor U10203 (N_10203,N_9682,N_8437);
and U10204 (N_10204,N_9068,N_8822);
and U10205 (N_10205,N_8365,N_8546);
nor U10206 (N_10206,N_8472,N_9419);
xnor U10207 (N_10207,N_9075,N_8121);
nand U10208 (N_10208,N_9088,N_9514);
or U10209 (N_10209,N_9157,N_9772);
nor U10210 (N_10210,N_8062,N_8537);
or U10211 (N_10211,N_8235,N_9847);
nand U10212 (N_10212,N_8490,N_8838);
nand U10213 (N_10213,N_8981,N_8908);
and U10214 (N_10214,N_8639,N_8680);
nand U10215 (N_10215,N_9222,N_9335);
xnor U10216 (N_10216,N_8988,N_8401);
and U10217 (N_10217,N_8615,N_8044);
nor U10218 (N_10218,N_8214,N_8900);
nand U10219 (N_10219,N_8926,N_8955);
nand U10220 (N_10220,N_8241,N_8360);
nor U10221 (N_10221,N_9079,N_9783);
nand U10222 (N_10222,N_8136,N_8866);
and U10223 (N_10223,N_9413,N_8201);
or U10224 (N_10224,N_8002,N_9058);
nand U10225 (N_10225,N_9504,N_8065);
and U10226 (N_10226,N_8761,N_8760);
or U10227 (N_10227,N_8461,N_8915);
nor U10228 (N_10228,N_9607,N_9542);
nor U10229 (N_10229,N_8957,N_8765);
and U10230 (N_10230,N_9287,N_8616);
xnor U10231 (N_10231,N_9192,N_8558);
xnor U10232 (N_10232,N_9197,N_9585);
and U10233 (N_10233,N_9827,N_8265);
nor U10234 (N_10234,N_8415,N_9913);
nor U10235 (N_10235,N_9956,N_9263);
and U10236 (N_10236,N_9647,N_8312);
or U10237 (N_10237,N_8868,N_8559);
xor U10238 (N_10238,N_9027,N_9389);
nand U10239 (N_10239,N_8448,N_8944);
xnor U10240 (N_10240,N_9164,N_8058);
xnor U10241 (N_10241,N_9384,N_9364);
xnor U10242 (N_10242,N_8194,N_8744);
nand U10243 (N_10243,N_9700,N_8005);
and U10244 (N_10244,N_8174,N_8072);
xor U10245 (N_10245,N_9326,N_8016);
or U10246 (N_10246,N_9374,N_8837);
nand U10247 (N_10247,N_9017,N_9689);
xor U10248 (N_10248,N_9714,N_9511);
xnor U10249 (N_10249,N_9455,N_9325);
xnor U10250 (N_10250,N_9996,N_9959);
xnor U10251 (N_10251,N_8149,N_8690);
xor U10252 (N_10252,N_8618,N_9960);
and U10253 (N_10253,N_8577,N_9440);
xor U10254 (N_10254,N_9599,N_8963);
nor U10255 (N_10255,N_8462,N_9904);
nor U10256 (N_10256,N_9863,N_9424);
nor U10257 (N_10257,N_8340,N_9251);
nor U10258 (N_10258,N_8385,N_9169);
or U10259 (N_10259,N_8131,N_8507);
xor U10260 (N_10260,N_8390,N_9527);
and U10261 (N_10261,N_9608,N_9484);
nor U10262 (N_10262,N_8130,N_9208);
and U10263 (N_10263,N_9005,N_8160);
or U10264 (N_10264,N_8684,N_9442);
or U10265 (N_10265,N_8334,N_8092);
and U10266 (N_10266,N_9926,N_8946);
or U10267 (N_10267,N_9464,N_8878);
and U10268 (N_10268,N_9220,N_8060);
or U10269 (N_10269,N_9013,N_8623);
nor U10270 (N_10270,N_9953,N_8137);
nor U10271 (N_10271,N_9334,N_8425);
xnor U10272 (N_10272,N_9467,N_8671);
xnor U10273 (N_10273,N_8779,N_8196);
nand U10274 (N_10274,N_8621,N_8806);
xor U10275 (N_10275,N_8540,N_8568);
or U10276 (N_10276,N_8734,N_8190);
and U10277 (N_10277,N_8354,N_8011);
and U10278 (N_10278,N_9434,N_9201);
nor U10279 (N_10279,N_9430,N_8541);
or U10280 (N_10280,N_9114,N_8302);
nor U10281 (N_10281,N_8068,N_9477);
or U10282 (N_10282,N_8633,N_9961);
nor U10283 (N_10283,N_9978,N_8545);
or U10284 (N_10284,N_9980,N_8405);
or U10285 (N_10285,N_9004,N_9271);
xor U10286 (N_10286,N_9940,N_8662);
and U10287 (N_10287,N_8350,N_9556);
nand U10288 (N_10288,N_9674,N_9450);
or U10289 (N_10289,N_8071,N_9938);
or U10290 (N_10290,N_9779,N_8823);
xor U10291 (N_10291,N_9687,N_9801);
xor U10292 (N_10292,N_8266,N_8305);
and U10293 (N_10293,N_8995,N_8586);
and U10294 (N_10294,N_8109,N_9018);
or U10295 (N_10295,N_8422,N_8295);
and U10296 (N_10296,N_8598,N_8522);
xnor U10297 (N_10297,N_8270,N_9524);
xor U10298 (N_10298,N_9468,N_8818);
or U10299 (N_10299,N_9874,N_8536);
nor U10300 (N_10300,N_9316,N_9268);
nor U10301 (N_10301,N_9795,N_9643);
nand U10302 (N_10302,N_8159,N_8703);
and U10303 (N_10303,N_8993,N_9342);
nand U10304 (N_10304,N_8820,N_8485);
xnor U10305 (N_10305,N_8994,N_9411);
or U10306 (N_10306,N_8610,N_8589);
nor U10307 (N_10307,N_9968,N_8704);
nor U10308 (N_10308,N_8594,N_8040);
or U10309 (N_10309,N_8096,N_9093);
nand U10310 (N_10310,N_9802,N_8440);
and U10311 (N_10311,N_9064,N_8081);
nand U10312 (N_10312,N_8256,N_8008);
nand U10313 (N_10313,N_8322,N_8105);
xor U10314 (N_10314,N_8320,N_8850);
nor U10315 (N_10315,N_9741,N_8901);
and U10316 (N_10316,N_9713,N_8314);
and U10317 (N_10317,N_9590,N_8672);
nor U10318 (N_10318,N_9991,N_8695);
nand U10319 (N_10319,N_8752,N_9592);
nand U10320 (N_10320,N_8465,N_8098);
or U10321 (N_10321,N_8502,N_9866);
nor U10322 (N_10322,N_9523,N_8880);
nor U10323 (N_10323,N_8826,N_9670);
nor U10324 (N_10324,N_8418,N_9391);
and U10325 (N_10325,N_8157,N_8624);
and U10326 (N_10326,N_8357,N_8709);
nand U10327 (N_10327,N_9297,N_8151);
or U10328 (N_10328,N_9421,N_8973);
or U10329 (N_10329,N_8729,N_8574);
or U10330 (N_10330,N_8694,N_9165);
xnor U10331 (N_10331,N_8276,N_8625);
or U10332 (N_10332,N_8117,N_8797);
and U10333 (N_10333,N_9510,N_8539);
or U10334 (N_10334,N_8158,N_8488);
or U10335 (N_10335,N_9051,N_8917);
nor U10336 (N_10336,N_9528,N_9496);
xor U10337 (N_10337,N_9636,N_9338);
and U10338 (N_10338,N_9351,N_9887);
xor U10339 (N_10339,N_9628,N_8553);
xnor U10340 (N_10340,N_9332,N_9113);
nor U10341 (N_10341,N_9138,N_8751);
and U10342 (N_10342,N_8829,N_8384);
and U10343 (N_10343,N_9103,N_8264);
and U10344 (N_10344,N_9502,N_9548);
or U10345 (N_10345,N_8582,N_9546);
xnor U10346 (N_10346,N_9069,N_9918);
nor U10347 (N_10347,N_9662,N_9837);
nor U10348 (N_10348,N_9012,N_9161);
nor U10349 (N_10349,N_9322,N_9232);
xnor U10350 (N_10350,N_9255,N_9625);
nor U10351 (N_10351,N_8984,N_8887);
nor U10352 (N_10352,N_8768,N_8126);
xnor U10353 (N_10353,N_8775,N_8495);
nand U10354 (N_10354,N_9191,N_9770);
or U10355 (N_10355,N_9472,N_9133);
nor U10356 (N_10356,N_9285,N_9404);
nor U10357 (N_10357,N_9261,N_9563);
nand U10358 (N_10358,N_8013,N_8533);
and U10359 (N_10359,N_8501,N_9383);
nor U10360 (N_10360,N_9049,N_9623);
xnor U10361 (N_10361,N_8453,N_8825);
nor U10362 (N_10362,N_9167,N_8812);
xor U10363 (N_10363,N_8318,N_9661);
xnor U10364 (N_10364,N_8749,N_9942);
or U10365 (N_10365,N_8308,N_8810);
and U10366 (N_10366,N_8208,N_9573);
xnor U10367 (N_10367,N_9877,N_9031);
and U10368 (N_10368,N_9821,N_9966);
xnor U10369 (N_10369,N_9494,N_9281);
xor U10370 (N_10370,N_8003,N_8348);
and U10371 (N_10371,N_9835,N_9330);
nor U10372 (N_10372,N_8107,N_9868);
and U10373 (N_10373,N_8851,N_8464);
nand U10374 (N_10374,N_9520,N_9948);
xor U10375 (N_10375,N_9454,N_9579);
nand U10376 (N_10376,N_8007,N_8170);
or U10377 (N_10377,N_9047,N_8821);
or U10378 (N_10378,N_8834,N_9781);
or U10379 (N_10379,N_8043,N_8996);
and U10380 (N_10380,N_9681,N_9675);
nand U10381 (N_10381,N_8004,N_8104);
or U10382 (N_10382,N_8491,N_9253);
and U10383 (N_10383,N_8542,N_8875);
and U10384 (N_10384,N_8741,N_9331);
xor U10385 (N_10385,N_9535,N_9690);
or U10386 (N_10386,N_9867,N_8306);
nand U10387 (N_10387,N_8742,N_9469);
nor U10388 (N_10388,N_9302,N_8067);
or U10389 (N_10389,N_8402,N_9515);
xor U10390 (N_10390,N_8066,N_8952);
or U10391 (N_10391,N_9062,N_9032);
or U10392 (N_10392,N_9707,N_8846);
nor U10393 (N_10393,N_8400,N_8450);
nand U10394 (N_10394,N_9011,N_9594);
or U10395 (N_10395,N_9405,N_8967);
xnor U10396 (N_10396,N_9735,N_9933);
xnor U10397 (N_10397,N_9231,N_9227);
or U10398 (N_10398,N_8321,N_8510);
xnor U10399 (N_10399,N_8442,N_8714);
or U10400 (N_10400,N_8634,N_9347);
or U10401 (N_10401,N_9691,N_9230);
nand U10402 (N_10402,N_8113,N_9748);
and U10403 (N_10403,N_8188,N_8332);
nor U10404 (N_10404,N_9606,N_8959);
or U10405 (N_10405,N_9817,N_8904);
nand U10406 (N_10406,N_9089,N_9876);
nand U10407 (N_10407,N_9990,N_8511);
nor U10408 (N_10408,N_9102,N_8912);
nor U10409 (N_10409,N_8240,N_9799);
or U10410 (N_10410,N_8758,N_8165);
or U10411 (N_10411,N_8090,N_9822);
nand U10412 (N_10412,N_8776,N_8781);
or U10413 (N_10413,N_8869,N_8229);
and U10414 (N_10414,N_9109,N_9914);
xnor U10415 (N_10415,N_9701,N_8412);
or U10416 (N_10416,N_9975,N_8186);
nor U10417 (N_10417,N_9750,N_9892);
and U10418 (N_10418,N_9453,N_9935);
and U10419 (N_10419,N_9901,N_9048);
xnor U10420 (N_10420,N_8175,N_9583);
nor U10421 (N_10421,N_8602,N_8045);
nor U10422 (N_10422,N_8743,N_8969);
xnor U10423 (N_10423,N_8920,N_8520);
nand U10424 (N_10424,N_9387,N_8431);
nand U10425 (N_10425,N_8211,N_8015);
nor U10426 (N_10426,N_8444,N_8745);
or U10427 (N_10427,N_9386,N_8811);
nor U10428 (N_10428,N_9642,N_8388);
nor U10429 (N_10429,N_8664,N_9518);
xor U10430 (N_10430,N_8268,N_8556);
or U10431 (N_10431,N_9361,N_9213);
or U10432 (N_10432,N_9046,N_9180);
and U10433 (N_10433,N_9843,N_8199);
and U10434 (N_10434,N_9397,N_8142);
or U10435 (N_10435,N_8630,N_8614);
or U10436 (N_10436,N_9506,N_9183);
or U10437 (N_10437,N_8377,N_8410);
nand U10438 (N_10438,N_9081,N_8853);
or U10439 (N_10439,N_8277,N_9889);
and U10440 (N_10440,N_9226,N_8022);
and U10441 (N_10441,N_8626,N_8666);
xnor U10442 (N_10442,N_9323,N_9597);
nand U10443 (N_10443,N_9593,N_9098);
xnor U10444 (N_10444,N_9992,N_8376);
nand U10445 (N_10445,N_9693,N_9566);
or U10446 (N_10446,N_8847,N_9522);
or U10447 (N_10447,N_8977,N_8762);
or U10448 (N_10448,N_8702,N_9516);
nand U10449 (N_10449,N_9932,N_8064);
and U10450 (N_10450,N_9656,N_9620);
nand U10451 (N_10451,N_9358,N_8267);
nor U10452 (N_10452,N_9060,N_8862);
xnor U10453 (N_10453,N_9266,N_8179);
nand U10454 (N_10454,N_8945,N_9224);
nor U10455 (N_10455,N_8951,N_9751);
nor U10456 (N_10456,N_9756,N_9955);
nand U10457 (N_10457,N_9537,N_9381);
and U10458 (N_10458,N_9446,N_9324);
xnor U10459 (N_10459,N_8087,N_8651);
nand U10460 (N_10460,N_9478,N_8339);
nor U10461 (N_10461,N_9544,N_9969);
nand U10462 (N_10462,N_9854,N_9329);
or U10463 (N_10463,N_9252,N_8301);
and U10464 (N_10464,N_9452,N_8298);
nand U10465 (N_10465,N_9915,N_9313);
and U10466 (N_10466,N_9124,N_9965);
or U10467 (N_10467,N_9254,N_9211);
xnor U10468 (N_10468,N_9838,N_9276);
and U10469 (N_10469,N_9680,N_9580);
xnor U10470 (N_10470,N_8239,N_9747);
xnor U10471 (N_10471,N_8063,N_9059);
nor U10472 (N_10472,N_9717,N_8218);
xor U10473 (N_10473,N_8523,N_9298);
xor U10474 (N_10474,N_9355,N_9146);
xor U10475 (N_10475,N_9519,N_8938);
nand U10476 (N_10476,N_8791,N_8754);
nand U10477 (N_10477,N_8079,N_9137);
or U10478 (N_10478,N_9619,N_9834);
or U10479 (N_10479,N_8220,N_8195);
or U10480 (N_10480,N_8606,N_8407);
and U10481 (N_10481,N_8254,N_8466);
nand U10482 (N_10482,N_9210,N_9754);
xnor U10483 (N_10483,N_8017,N_8999);
nor U10484 (N_10484,N_8794,N_8344);
xnor U10485 (N_10485,N_8292,N_8805);
xor U10486 (N_10486,N_9664,N_9804);
and U10487 (N_10487,N_9292,N_9363);
or U10488 (N_10488,N_9536,N_9375);
xnor U10489 (N_10489,N_9020,N_8396);
xnor U10490 (N_10490,N_9897,N_9857);
nand U10491 (N_10491,N_9762,N_8931);
nand U10492 (N_10492,N_9820,N_9962);
nand U10493 (N_10493,N_8940,N_9110);
and U10494 (N_10494,N_8787,N_8580);
or U10495 (N_10495,N_9630,N_8283);
nand U10496 (N_10496,N_9666,N_8503);
nand U10497 (N_10497,N_8375,N_8359);
and U10498 (N_10498,N_8839,N_9090);
nand U10499 (N_10499,N_9154,N_9622);
nand U10500 (N_10500,N_9728,N_8398);
xnor U10501 (N_10501,N_8792,N_8513);
nand U10502 (N_10502,N_8910,N_8352);
nand U10503 (N_10503,N_8417,N_9949);
nor U10504 (N_10504,N_8085,N_8169);
and U10505 (N_10505,N_9198,N_9087);
nor U10506 (N_10506,N_8665,N_8653);
and U10507 (N_10507,N_8529,N_8675);
nand U10508 (N_10508,N_8572,N_9438);
or U10509 (N_10509,N_8840,N_9432);
xor U10510 (N_10510,N_8990,N_8207);
nand U10511 (N_10511,N_8721,N_8697);
and U10512 (N_10512,N_8852,N_8428);
xor U10513 (N_10513,N_8628,N_8659);
and U10514 (N_10514,N_8863,N_9441);
nand U10515 (N_10515,N_9120,N_8682);
or U10516 (N_10516,N_8206,N_9731);
nand U10517 (N_10517,N_8249,N_9970);
nor U10518 (N_10518,N_9603,N_9906);
and U10519 (N_10519,N_9186,N_9241);
xor U10520 (N_10520,N_9872,N_9173);
nor U10521 (N_10521,N_8282,N_9997);
and U10522 (N_10522,N_9716,N_9621);
nor U10523 (N_10523,N_9853,N_8858);
xnor U10524 (N_10524,N_9235,N_8095);
xnor U10525 (N_10525,N_8803,N_8619);
and U10526 (N_10526,N_8379,N_9345);
nand U10527 (N_10527,N_8150,N_8033);
xnor U10528 (N_10528,N_8645,N_8225);
and U10529 (N_10529,N_8168,N_8281);
or U10530 (N_10530,N_8769,N_9776);
nand U10531 (N_10531,N_9943,N_9318);
nor U10532 (N_10532,N_9637,N_8767);
xor U10533 (N_10533,N_8636,N_8234);
nor U10534 (N_10534,N_9797,N_9825);
nand U10535 (N_10535,N_9159,N_8565);
and U10536 (N_10536,N_9761,N_9082);
or U10537 (N_10537,N_9633,N_8835);
and U10538 (N_10538,N_9084,N_9053);
xor U10539 (N_10539,N_9951,N_8902);
or U10540 (N_10540,N_8303,N_9634);
or U10541 (N_10541,N_9500,N_8715);
or U10542 (N_10542,N_9508,N_9304);
xnor U10543 (N_10543,N_9554,N_9181);
nor U10544 (N_10544,N_8909,N_8816);
nor U10545 (N_10545,N_9884,N_9759);
nand U10546 (N_10546,N_9194,N_9648);
xnor U10547 (N_10547,N_9531,N_9881);
and U10548 (N_10548,N_8571,N_8928);
nor U10549 (N_10549,N_8155,N_9244);
and U10550 (N_10550,N_8290,N_9188);
xnor U10551 (N_10551,N_8247,N_9493);
and U10552 (N_10552,N_9115,N_9247);
and U10553 (N_10553,N_8278,N_8549);
xor U10554 (N_10554,N_9371,N_9380);
nand U10555 (N_10555,N_9812,N_9530);
or U10556 (N_10556,N_9144,N_9466);
xnor U10557 (N_10557,N_9730,N_8701);
and U10558 (N_10558,N_8911,N_8219);
xnor U10559 (N_10559,N_9903,N_9036);
nand U10560 (N_10560,N_9283,N_8061);
xor U10561 (N_10561,N_9141,N_8021);
nand U10562 (N_10562,N_8783,N_8189);
and U10563 (N_10563,N_8962,N_8032);
nand U10564 (N_10564,N_8950,N_9849);
or U10565 (N_10565,N_8202,N_9199);
or U10566 (N_10566,N_8285,N_8093);
nor U10567 (N_10567,N_8611,N_8146);
or U10568 (N_10568,N_9352,N_9396);
or U10569 (N_10569,N_9218,N_9547);
xor U10570 (N_10570,N_9998,N_8128);
xor U10571 (N_10571,N_9319,N_8329);
nand U10572 (N_10572,N_9498,N_9844);
nand U10573 (N_10573,N_9745,N_8975);
nor U10574 (N_10574,N_9301,N_8560);
xnor U10575 (N_10575,N_9333,N_8198);
nand U10576 (N_10576,N_8191,N_9362);
nand U10577 (N_10577,N_9641,N_8819);
xnor U10578 (N_10578,N_8780,N_9586);
nor U10579 (N_10579,N_8970,N_9415);
nand U10580 (N_10580,N_8112,N_9644);
nand U10581 (N_10581,N_8263,N_9394);
and U10582 (N_10582,N_8567,N_9559);
nor U10583 (N_10583,N_9312,N_9651);
and U10584 (N_10584,N_9274,N_9107);
xnor U10585 (N_10585,N_8740,N_9249);
xnor U10586 (N_10586,N_8555,N_9917);
xor U10587 (N_10587,N_9526,N_9063);
nor U10588 (N_10588,N_9829,N_8286);
or U10589 (N_10589,N_9019,N_9824);
or U10590 (N_10590,N_8193,N_9091);
or U10591 (N_10591,N_8748,N_8764);
or U10592 (N_10592,N_9869,N_8460);
xor U10593 (N_10593,N_8949,N_9650);
nand U10594 (N_10594,N_8446,N_9131);
nand U10595 (N_10595,N_8473,N_9207);
xor U10596 (N_10596,N_9679,N_8564);
and U10597 (N_10597,N_9614,N_9409);
and U10598 (N_10598,N_9189,N_8706);
xor U10599 (N_10599,N_9507,N_9976);
and U10600 (N_10600,N_8817,N_9350);
xor U10601 (N_10601,N_8604,N_8257);
nand U10602 (N_10602,N_9746,N_8489);
and U10603 (N_10603,N_9987,N_9395);
nor U10604 (N_10604,N_9982,N_9072);
xor U10605 (N_10605,N_9353,N_8289);
and U10606 (N_10606,N_9993,N_8346);
or U10607 (N_10607,N_9365,N_8246);
xor U10608 (N_10608,N_9382,N_9444);
nand U10609 (N_10609,N_8028,N_9320);
and U10610 (N_10610,N_8023,N_8296);
or U10611 (N_10611,N_9875,N_8936);
nor U10612 (N_10612,N_9550,N_9567);
nand U10613 (N_10613,N_9479,N_8924);
xor U10614 (N_10614,N_9828,N_9782);
or U10615 (N_10615,N_8250,N_9166);
nand U10616 (N_10616,N_9505,N_8620);
or U10617 (N_10617,N_9074,N_9203);
xnor U10618 (N_10618,N_9006,N_8637);
nand U10619 (N_10619,N_8830,N_8125);
or U10620 (N_10620,N_8925,N_8655);
or U10621 (N_10621,N_8371,N_8046);
nor U10622 (N_10622,N_9539,N_9425);
xor U10623 (N_10623,N_8504,N_8233);
or U10624 (N_10624,N_9420,N_9532);
or U10625 (N_10625,N_9485,N_8368);
and U10626 (N_10626,N_8932,N_9260);
xnor U10627 (N_10627,N_9459,N_8468);
nand U10628 (N_10628,N_9677,N_9445);
nor U10629 (N_10629,N_8674,N_9864);
and U10630 (N_10630,N_8974,N_8173);
nor U10631 (N_10631,N_8508,N_9340);
or U10632 (N_10632,N_9744,N_9449);
nor U10633 (N_10633,N_8342,N_9385);
xnor U10634 (N_10634,N_9930,N_9288);
xor U10635 (N_10635,N_9086,N_8736);
nand U10636 (N_10636,N_8237,N_9836);
nor U10637 (N_10637,N_9581,N_8617);
or U10638 (N_10638,N_9035,N_9604);
or U10639 (N_10639,N_9774,N_9673);
nor U10640 (N_10640,N_9126,N_8476);
or U10641 (N_10641,N_8287,N_8992);
nand U10642 (N_10642,N_8474,N_8753);
or U10643 (N_10643,N_8041,N_9671);
or U10644 (N_10644,N_8273,N_8323);
and U10645 (N_10645,N_8316,N_8111);
or U10646 (N_10646,N_9788,N_9080);
or U10647 (N_10647,N_8477,N_8077);
and U10648 (N_10648,N_8226,N_9398);
xnor U10649 (N_10649,N_9480,N_9418);
nand U10650 (N_10650,N_9711,N_9248);
nand U10651 (N_10651,N_8727,N_9294);
or U10652 (N_10652,N_9406,N_8683);
xnor U10653 (N_10653,N_9158,N_8747);
xor U10654 (N_10654,N_9653,N_8261);
or U10655 (N_10655,N_8274,N_8790);
and U10656 (N_10656,N_8987,N_9977);
xor U10657 (N_10657,N_9061,N_9299);
or U10658 (N_10658,N_8204,N_9609);
nor U10659 (N_10659,N_8353,N_9495);
nand U10660 (N_10660,N_9626,N_9885);
and U10661 (N_10661,N_9646,N_8933);
and U10662 (N_10662,N_9443,N_8935);
or U10663 (N_10663,N_9601,N_8972);
and U10664 (N_10664,N_9456,N_9475);
xnor U10665 (N_10665,N_9128,N_9284);
nand U10666 (N_10666,N_8326,N_8896);
nor U10667 (N_10667,N_8177,N_9457);
xor U10668 (N_10668,N_8757,N_9787);
nand U10669 (N_10669,N_9807,N_9894);
xor U10670 (N_10670,N_8566,N_9654);
nor U10671 (N_10671,N_8573,N_8613);
nand U10672 (N_10672,N_8723,N_9919);
nor U10673 (N_10673,N_8543,N_8965);
nor U10674 (N_10674,N_9344,N_9145);
or U10675 (N_10675,N_8279,N_8953);
nand U10676 (N_10676,N_9814,N_9236);
nor U10677 (N_10677,N_8552,N_9216);
or U10678 (N_10678,N_8678,N_9602);
and U10679 (N_10679,N_9811,N_9852);
nor U10680 (N_10680,N_8882,N_8814);
or U10681 (N_10681,N_9117,N_9767);
xnor U10682 (N_10682,N_8020,N_8799);
or U10683 (N_10683,N_9311,N_8718);
and U10684 (N_10684,N_9187,N_9639);
nand U10685 (N_10685,N_9752,N_9652);
xor U10686 (N_10686,N_8251,N_9710);
nand U10687 (N_10687,N_9196,N_9810);
or U10688 (N_10688,N_9981,N_9473);
xnor U10689 (N_10689,N_9286,N_9575);
nand U10690 (N_10690,N_8311,N_9562);
xor U10691 (N_10691,N_8650,N_8223);
nor U10692 (N_10692,N_9855,N_9010);
nor U10693 (N_10693,N_9692,N_8482);
and U10694 (N_10694,N_9549,N_8642);
nor U10695 (N_10695,N_8141,N_9765);
nand U10696 (N_10696,N_8569,N_9676);
xnor U10697 (N_10697,N_8248,N_9206);
or U10698 (N_10698,N_8711,N_9667);
and U10699 (N_10699,N_8200,N_8487);
nand U10700 (N_10700,N_9816,N_9234);
and U10701 (N_10701,N_8516,N_9813);
nor U10702 (N_10702,N_8941,N_9784);
or U10703 (N_10703,N_8788,N_8052);
and U10704 (N_10704,N_8433,N_9803);
nand U10705 (N_10705,N_9291,N_9140);
nor U10706 (N_10706,N_8238,N_9392);
xor U10707 (N_10707,N_9033,N_8514);
xor U10708 (N_10708,N_8132,N_8304);
xor U10709 (N_10709,N_8879,N_8881);
and U10710 (N_10710,N_8084,N_8392);
or U10711 (N_10711,N_9560,N_9112);
nor U10712 (N_10712,N_9412,N_9193);
xor U10713 (N_10713,N_9139,N_8101);
or U10714 (N_10714,N_9796,N_8755);
nor U10715 (N_10715,N_8397,N_9924);
nand U10716 (N_10716,N_9699,N_9073);
and U10717 (N_10717,N_9553,N_9219);
or U10718 (N_10718,N_8335,N_9846);
nand U10719 (N_10719,N_9640,N_8152);
or U10720 (N_10720,N_9238,N_8018);
or U10721 (N_10721,N_8980,N_8260);
xnor U10722 (N_10722,N_9367,N_9354);
or U10723 (N_10723,N_9706,N_9043);
and U10724 (N_10724,N_9791,N_9568);
and U10725 (N_10725,N_9153,N_8870);
xor U10726 (N_10726,N_8583,N_9931);
nand U10727 (N_10727,N_8921,N_8010);
or U10728 (N_10728,N_9709,N_9615);
nor U10729 (N_10729,N_9303,N_8861);
and U10730 (N_10730,N_8867,N_8349);
and U10731 (N_10731,N_9610,N_8681);
nor U10732 (N_10732,N_9999,N_9094);
xnor U10733 (N_10733,N_8386,N_9833);
nand U10734 (N_10734,N_8443,N_9026);
and U10735 (N_10735,N_9818,N_8836);
nand U10736 (N_10736,N_9368,N_9127);
xnor U10737 (N_10737,N_9272,N_8801);
or U10738 (N_10738,N_9039,N_8842);
nand U10739 (N_10739,N_8876,N_9481);
nor U10740 (N_10740,N_8284,N_8722);
nand U10741 (N_10741,N_9257,N_8903);
xnor U10742 (N_10742,N_9111,N_8414);
nand U10743 (N_10743,N_9916,N_9065);
xnor U10744 (N_10744,N_9760,N_8658);
and U10745 (N_10745,N_9587,N_9873);
nand U10746 (N_10746,N_9163,N_9798);
and U10747 (N_10747,N_8404,N_9223);
or U10748 (N_10748,N_8050,N_8854);
or U10749 (N_10749,N_8122,N_9423);
or U10750 (N_10750,N_9578,N_8661);
and U10751 (N_10751,N_8456,N_9403);
xnor U10752 (N_10752,N_8145,N_8989);
nand U10753 (N_10753,N_9888,N_8687);
or U10754 (N_10754,N_8299,N_9458);
or U10755 (N_10755,N_8083,N_9488);
nor U10756 (N_10756,N_8644,N_8692);
nor U10757 (N_10757,N_9509,N_8943);
and U10758 (N_10758,N_9179,N_9861);
or U10759 (N_10759,N_8372,N_8116);
nor U10760 (N_10760,N_9008,N_8786);
or U10761 (N_10761,N_9617,N_8985);
xor U10762 (N_10762,N_8364,N_9016);
xor U10763 (N_10763,N_9946,N_9958);
or U10764 (N_10764,N_9541,N_9910);
nand U10765 (N_10765,N_8129,N_8184);
and U10766 (N_10766,N_9489,N_8927);
or U10767 (N_10767,N_9221,N_8759);
and U10768 (N_10768,N_8197,N_9293);
or U10769 (N_10769,N_8463,N_9739);
xor U10770 (N_10770,N_9589,N_9119);
xor U10771 (N_10771,N_9178,N_8309);
xor U10772 (N_10772,N_9638,N_9858);
or U10773 (N_10773,N_9135,N_9972);
nand U10774 (N_10774,N_8688,N_8719);
or U10775 (N_10775,N_9721,N_8182);
and U10776 (N_10776,N_9130,N_9436);
nor U10777 (N_10777,N_8492,N_8548);
and U10778 (N_10778,N_9030,N_9132);
and U10779 (N_10779,N_9422,N_8300);
and U10780 (N_10780,N_9658,N_9512);
and U10781 (N_10781,N_9963,N_9805);
nor U10782 (N_10782,N_8459,N_9944);
nor U10783 (N_10783,N_9830,N_8726);
nor U10784 (N_10784,N_8070,N_9209);
nor U10785 (N_10785,N_8960,N_9176);
nand U10786 (N_10786,N_8831,N_8813);
or U10787 (N_10787,N_8720,N_8259);
xnor U10788 (N_10788,N_8841,N_9071);
or U10789 (N_10789,N_8434,N_8527);
or U10790 (N_10790,N_8147,N_8877);
xnor U10791 (N_10791,N_8100,N_9310);
nand U10792 (N_10792,N_9786,N_8493);
nand U10793 (N_10793,N_9856,N_9054);
nand U10794 (N_10794,N_8366,N_9794);
nand U10795 (N_10795,N_8976,N_9315);
xnor U10796 (N_10796,N_8230,N_9920);
or U10797 (N_10797,N_9552,N_9182);
xnor U10798 (N_10798,N_9376,N_9886);
nor U10799 (N_10799,N_9205,N_9346);
nor U10800 (N_10800,N_8049,N_8185);
or U10801 (N_10801,N_8954,N_8971);
xor U10802 (N_10802,N_9290,N_9250);
nand U10803 (N_10803,N_8873,N_9971);
xnor U10804 (N_10804,N_8001,N_9357);
nand U10805 (N_10805,N_9476,N_8519);
and U10806 (N_10806,N_9300,N_9202);
xnor U10807 (N_10807,N_8631,N_8019);
nand U10808 (N_10808,N_9390,N_8856);
and U10809 (N_10809,N_9267,N_8216);
nor U10810 (N_10810,N_9143,N_9595);
and U10811 (N_10811,N_9616,N_9725);
xor U10812 (N_10812,N_8676,N_8436);
and U10813 (N_10813,N_8373,N_9517);
and U10814 (N_10814,N_9034,N_8886);
or U10815 (N_10815,N_8293,N_9314);
nor U10816 (N_10816,N_8420,N_9279);
nand U10817 (N_10817,N_9792,N_9270);
or U10818 (N_10818,N_8657,N_8310);
nor U10819 (N_10819,N_9407,N_8429);
nand U10820 (N_10820,N_9170,N_9256);
xnor U10821 (N_10821,N_8958,N_9076);
nor U10822 (N_10822,N_9359,N_9136);
xor U10823 (N_10823,N_9378,N_9773);
nand U10824 (N_10824,N_9722,N_9839);
nand U10825 (N_10825,N_8883,N_8855);
and U10826 (N_10826,N_9571,N_8809);
nand U10827 (N_10827,N_9305,N_9819);
nor U10828 (N_10828,N_9695,N_8983);
or U10829 (N_10829,N_9923,N_8395);
xnor U10830 (N_10830,N_8123,N_9895);
and U10831 (N_10831,N_9605,N_8328);
nor U10832 (N_10832,N_9694,N_8172);
and U10833 (N_10833,N_9066,N_8210);
nand U10834 (N_10834,N_9995,N_9900);
and U10835 (N_10835,N_8156,N_8183);
and U10836 (N_10836,N_8660,N_9883);
xor U10837 (N_10837,N_9768,N_9766);
nor U10838 (N_10838,N_8471,N_8562);
and U10839 (N_10839,N_8733,N_9317);
nand U10840 (N_10840,N_9685,N_9727);
and U10841 (N_10841,N_9343,N_9427);
xnor U10842 (N_10842,N_9598,N_8114);
or U10843 (N_10843,N_8509,N_9237);
nand U10844 (N_10844,N_8526,N_9570);
and U10845 (N_10845,N_9435,N_9152);
nand U10846 (N_10846,N_9101,N_8435);
or U10847 (N_10847,N_9582,N_9753);
and U10848 (N_10848,N_9414,N_9771);
nor U10849 (N_10849,N_8012,N_8677);
and U10850 (N_10850,N_9591,N_9950);
nand U10851 (N_10851,N_9278,N_9697);
nand U10852 (N_10852,N_9734,N_9289);
nand U10853 (N_10853,N_8939,N_9282);
or U10854 (N_10854,N_8708,N_8324);
xor U10855 (N_10855,N_9437,N_8331);
or U10856 (N_10856,N_9195,N_8778);
nor U10857 (N_10857,N_9979,N_8231);
nand U10858 (N_10858,N_8367,N_8036);
or U10859 (N_10859,N_9660,N_8581);
xor U10860 (N_10860,N_9024,N_8253);
xor U10861 (N_10861,N_8393,N_9740);
xnor U10862 (N_10862,N_9416,N_8124);
nand U10863 (N_10863,N_8258,N_8843);
or U10864 (N_10864,N_8224,N_8864);
nand U10865 (N_10865,N_9983,N_9501);
nor U10866 (N_10866,N_9243,N_9757);
nor U10867 (N_10867,N_8849,N_8421);
nand U10868 (N_10868,N_9148,N_9865);
and U10869 (N_10869,N_9099,N_8073);
xor U10870 (N_10870,N_8550,N_8409);
or U10871 (N_10871,N_9905,N_8595);
and U10872 (N_10872,N_9939,N_8860);
xnor U10873 (N_10873,N_9125,N_9624);
nor U10874 (N_10874,N_8317,N_9543);
nand U10875 (N_10875,N_9215,N_9551);
xor U10876 (N_10876,N_9588,N_9402);
and U10877 (N_10877,N_9742,N_8575);
or U10878 (N_10878,N_9841,N_8213);
and U10879 (N_10879,N_9379,N_9029);
nand U10880 (N_10880,N_9041,N_8209);
and U10881 (N_10881,N_9696,N_9185);
and U10882 (N_10882,N_8048,N_8127);
nand U10883 (N_10883,N_8203,N_8532);
nor U10884 (N_10884,N_8770,N_9050);
and U10885 (N_10885,N_8603,N_8648);
or U10886 (N_10886,N_9860,N_9339);
and U10887 (N_10887,N_9097,N_9984);
nand U10888 (N_10888,N_8668,N_8025);
nand U10889 (N_10889,N_8447,N_8074);
and U10890 (N_10890,N_8557,N_8076);
or U10891 (N_10891,N_9336,N_9555);
xor U10892 (N_10892,N_8215,N_8171);
xor U10893 (N_10893,N_8262,N_9388);
or U10894 (N_10894,N_9985,N_8080);
nor U10895 (N_10895,N_8445,N_9463);
nand U10896 (N_10896,N_9045,N_9077);
and U10897 (N_10897,N_8525,N_8228);
nand U10898 (N_10898,N_8712,N_8483);
xor U10899 (N_10899,N_9377,N_9928);
and U10900 (N_10900,N_8097,N_8272);
and U10901 (N_10901,N_8656,N_9190);
nand U10902 (N_10902,N_8078,N_9929);
nor U10903 (N_10903,N_8891,N_8777);
xnor U10904 (N_10904,N_9974,N_8942);
or U10905 (N_10905,N_8205,N_8531);
or U10906 (N_10906,N_8089,N_9429);
nor U10907 (N_10907,N_8362,N_9014);
or U10908 (N_10908,N_8597,N_8037);
nand U10909 (N_10909,N_8110,N_9842);
nor U10910 (N_10910,N_9229,N_9497);
xor U10911 (N_10911,N_8355,N_8789);
nand U10912 (N_10912,N_8947,N_8785);
xnor U10913 (N_10913,N_8937,N_9618);
or U10914 (N_10914,N_8135,N_8391);
nand U10915 (N_10915,N_8588,N_8102);
nor U10916 (N_10916,N_8534,N_8796);
nand U10917 (N_10917,N_8888,N_8413);
nand U10918 (N_10918,N_9672,N_8735);
xnor U10919 (N_10919,N_8914,N_9240);
and U10920 (N_10920,N_9095,N_8763);
xor U10921 (N_10921,N_9280,N_8913);
xnor U10922 (N_10922,N_9635,N_8874);
xor U10923 (N_10923,N_8518,N_8647);
or U10924 (N_10924,N_9715,N_9393);
xor U10925 (N_10925,N_8034,N_9891);
nand U10926 (N_10926,N_8086,N_9684);
nand U10927 (N_10927,N_8133,N_9632);
nand U10928 (N_10928,N_8732,N_8982);
nand U10929 (N_10929,N_8481,N_8426);
xor U10930 (N_10930,N_8528,N_9426);
xor U10931 (N_10931,N_9723,N_9337);
nor U10932 (N_10932,N_8403,N_9600);
nand U10933 (N_10933,N_8380,N_9341);
nand U10934 (N_10934,N_8600,N_8187);
nand U10935 (N_10935,N_8275,N_8892);
nor U10936 (N_10936,N_8640,N_8632);
nand U10937 (N_10937,N_8479,N_8591);
nor U10938 (N_10938,N_8269,N_9410);
or U10939 (N_10939,N_8601,N_9678);
nor U10940 (N_10940,N_8922,N_9941);
and U10941 (N_10941,N_8793,N_8119);
xor U10942 (N_10942,N_9022,N_8679);
or U10943 (N_10943,N_9246,N_9649);
nand U10944 (N_10944,N_9704,N_9491);
or U10945 (N_10945,N_9486,N_8394);
or U10946 (N_10946,N_8427,N_8584);
xnor U10947 (N_10947,N_9627,N_8685);
or U10948 (N_10948,N_8505,N_9764);
xnor U10949 (N_10949,N_8054,N_9780);
nor U10950 (N_10950,N_8361,N_9023);
or U10951 (N_10951,N_8399,N_8612);
or U10952 (N_10952,N_8059,N_8000);
and U10953 (N_10953,N_8222,N_9360);
nor U10954 (N_10954,N_8053,N_8930);
and U10955 (N_10955,N_9789,N_8014);
and U10956 (N_10956,N_9038,N_8325);
or U10957 (N_10957,N_8638,N_9162);
xor U10958 (N_10958,N_9417,N_9129);
and U10959 (N_10959,N_9659,N_8094);
nand U10960 (N_10960,N_8730,N_9462);
nand U10961 (N_10961,N_9785,N_9296);
or U10962 (N_10962,N_8506,N_8800);
nor U10963 (N_10963,N_9957,N_8808);
nand U10964 (N_10964,N_9893,N_9937);
nand U10965 (N_10965,N_8798,N_9175);
nor U10966 (N_10966,N_9702,N_8705);
nor U10967 (N_10967,N_8406,N_9912);
nor U10968 (N_10968,N_9369,N_9540);
or U10969 (N_10969,N_9994,N_8898);
nor U10970 (N_10970,N_8315,N_9482);
nor U10971 (N_10971,N_8828,N_8824);
or U10972 (N_10972,N_9007,N_8345);
xor U10973 (N_10973,N_8978,N_8378);
nand U10974 (N_10974,N_8338,N_8731);
nand U10975 (N_10975,N_8221,N_8069);
xnor U10976 (N_10976,N_8563,N_8827);
and U10977 (N_10977,N_9356,N_8500);
and U10978 (N_10978,N_8336,N_9085);
nor U10979 (N_10979,N_9070,N_9348);
nor U10980 (N_10980,N_9986,N_8521);
nor U10981 (N_10981,N_8387,N_8895);
nor U10982 (N_10982,N_9513,N_8451);
nor U10983 (N_10983,N_8108,N_8890);
or U10984 (N_10984,N_8408,N_8865);
or U10985 (N_10985,N_9487,N_8120);
or U10986 (N_10986,N_9121,N_8280);
xnor U10987 (N_10987,N_9719,N_9100);
xor U10988 (N_10988,N_9142,N_9108);
and U10989 (N_10989,N_9973,N_9755);
or U10990 (N_10990,N_9726,N_8370);
nor U10991 (N_10991,N_8030,N_8997);
or U10992 (N_10992,N_8570,N_9657);
or U10993 (N_10993,N_9533,N_9104);
and U10994 (N_10994,N_9778,N_8497);
nor U10995 (N_10995,N_9611,N_9952);
nand U10996 (N_10996,N_8411,N_8608);
nand U10997 (N_10997,N_8337,N_9655);
and U10998 (N_10998,N_8252,N_8889);
nand U10999 (N_10999,N_8691,N_9529);
and U11000 (N_11000,N_9915,N_9017);
or U11001 (N_11001,N_9778,N_8058);
and U11002 (N_11002,N_9536,N_9974);
nand U11003 (N_11003,N_8673,N_8743);
nor U11004 (N_11004,N_9911,N_9118);
xnor U11005 (N_11005,N_9930,N_8544);
and U11006 (N_11006,N_8028,N_8314);
nand U11007 (N_11007,N_9111,N_9515);
or U11008 (N_11008,N_8424,N_8199);
or U11009 (N_11009,N_9323,N_9652);
nand U11010 (N_11010,N_9969,N_8731);
or U11011 (N_11011,N_8749,N_9106);
xor U11012 (N_11012,N_9126,N_9250);
xnor U11013 (N_11013,N_8431,N_8730);
or U11014 (N_11014,N_8616,N_8288);
or U11015 (N_11015,N_8492,N_9673);
nand U11016 (N_11016,N_8067,N_8101);
nand U11017 (N_11017,N_9726,N_8243);
nor U11018 (N_11018,N_8192,N_8039);
nand U11019 (N_11019,N_8885,N_9388);
and U11020 (N_11020,N_8641,N_8828);
nand U11021 (N_11021,N_9908,N_8496);
and U11022 (N_11022,N_8118,N_9570);
and U11023 (N_11023,N_8957,N_8364);
xnor U11024 (N_11024,N_9208,N_8618);
nor U11025 (N_11025,N_8717,N_9166);
nand U11026 (N_11026,N_8443,N_8484);
or U11027 (N_11027,N_9302,N_9327);
and U11028 (N_11028,N_9695,N_9188);
nor U11029 (N_11029,N_8848,N_9198);
xor U11030 (N_11030,N_8036,N_8694);
nand U11031 (N_11031,N_8505,N_9557);
nand U11032 (N_11032,N_9707,N_9025);
nand U11033 (N_11033,N_9734,N_8860);
and U11034 (N_11034,N_9021,N_9269);
nor U11035 (N_11035,N_9505,N_8235);
nor U11036 (N_11036,N_8287,N_8860);
xnor U11037 (N_11037,N_9130,N_9014);
nand U11038 (N_11038,N_8952,N_8670);
xor U11039 (N_11039,N_9377,N_8459);
nand U11040 (N_11040,N_9814,N_9284);
or U11041 (N_11041,N_8616,N_9985);
or U11042 (N_11042,N_8085,N_8010);
nor U11043 (N_11043,N_8301,N_8862);
xor U11044 (N_11044,N_9650,N_8968);
nand U11045 (N_11045,N_8650,N_9870);
xor U11046 (N_11046,N_8671,N_8278);
and U11047 (N_11047,N_8672,N_9667);
or U11048 (N_11048,N_9900,N_9348);
xnor U11049 (N_11049,N_8021,N_9228);
nor U11050 (N_11050,N_8223,N_9435);
and U11051 (N_11051,N_9019,N_9607);
and U11052 (N_11052,N_8017,N_8694);
xnor U11053 (N_11053,N_9321,N_8054);
or U11054 (N_11054,N_8359,N_8118);
xnor U11055 (N_11055,N_8081,N_9562);
nand U11056 (N_11056,N_9610,N_8365);
and U11057 (N_11057,N_8365,N_8990);
and U11058 (N_11058,N_9072,N_9706);
nor U11059 (N_11059,N_9267,N_8976);
nor U11060 (N_11060,N_8441,N_9221);
nand U11061 (N_11061,N_9510,N_8469);
or U11062 (N_11062,N_8013,N_8416);
or U11063 (N_11063,N_9221,N_9278);
nand U11064 (N_11064,N_9808,N_8081);
and U11065 (N_11065,N_8543,N_8430);
and U11066 (N_11066,N_8917,N_9942);
nand U11067 (N_11067,N_9331,N_9076);
and U11068 (N_11068,N_9993,N_9011);
and U11069 (N_11069,N_9360,N_9647);
and U11070 (N_11070,N_9176,N_8862);
and U11071 (N_11071,N_9144,N_8108);
xnor U11072 (N_11072,N_8844,N_9823);
xnor U11073 (N_11073,N_8579,N_9833);
and U11074 (N_11074,N_9100,N_8414);
nand U11075 (N_11075,N_8766,N_9470);
xor U11076 (N_11076,N_8963,N_9826);
xor U11077 (N_11077,N_8594,N_9991);
or U11078 (N_11078,N_9707,N_9748);
or U11079 (N_11079,N_8671,N_9814);
nor U11080 (N_11080,N_9792,N_8742);
nor U11081 (N_11081,N_8173,N_9247);
xor U11082 (N_11082,N_8782,N_9859);
nand U11083 (N_11083,N_8514,N_8053);
and U11084 (N_11084,N_8209,N_9546);
nand U11085 (N_11085,N_9793,N_8764);
nor U11086 (N_11086,N_8920,N_8740);
and U11087 (N_11087,N_9573,N_9500);
nand U11088 (N_11088,N_9161,N_8742);
or U11089 (N_11089,N_8888,N_9526);
and U11090 (N_11090,N_9858,N_8725);
and U11091 (N_11091,N_9971,N_8892);
nor U11092 (N_11092,N_8455,N_8821);
nand U11093 (N_11093,N_8841,N_9872);
and U11094 (N_11094,N_9055,N_9824);
nand U11095 (N_11095,N_9885,N_8155);
nand U11096 (N_11096,N_9575,N_8880);
nor U11097 (N_11097,N_8365,N_8082);
nand U11098 (N_11098,N_9677,N_8647);
nand U11099 (N_11099,N_8330,N_9829);
or U11100 (N_11100,N_9259,N_8148);
or U11101 (N_11101,N_8757,N_8697);
nor U11102 (N_11102,N_8310,N_9078);
or U11103 (N_11103,N_9780,N_8988);
nand U11104 (N_11104,N_9211,N_8731);
nand U11105 (N_11105,N_9566,N_9981);
nand U11106 (N_11106,N_8886,N_9115);
nand U11107 (N_11107,N_8397,N_9798);
or U11108 (N_11108,N_9063,N_8522);
nand U11109 (N_11109,N_8774,N_9657);
nand U11110 (N_11110,N_9234,N_9314);
nor U11111 (N_11111,N_9922,N_8113);
nand U11112 (N_11112,N_8196,N_9521);
or U11113 (N_11113,N_8979,N_8872);
nor U11114 (N_11114,N_9620,N_9293);
and U11115 (N_11115,N_8511,N_8392);
nor U11116 (N_11116,N_8798,N_8124);
nand U11117 (N_11117,N_8133,N_9012);
or U11118 (N_11118,N_9506,N_9416);
and U11119 (N_11119,N_9558,N_8617);
and U11120 (N_11120,N_9528,N_9404);
nor U11121 (N_11121,N_8540,N_8593);
and U11122 (N_11122,N_8217,N_8506);
and U11123 (N_11123,N_8039,N_8186);
nor U11124 (N_11124,N_9799,N_9901);
nand U11125 (N_11125,N_9193,N_9735);
nand U11126 (N_11126,N_8926,N_9071);
nand U11127 (N_11127,N_9380,N_8548);
nand U11128 (N_11128,N_8013,N_8805);
and U11129 (N_11129,N_8268,N_8242);
or U11130 (N_11130,N_9211,N_9943);
and U11131 (N_11131,N_8345,N_8409);
nand U11132 (N_11132,N_8203,N_9032);
and U11133 (N_11133,N_8495,N_8308);
or U11134 (N_11134,N_8276,N_8203);
or U11135 (N_11135,N_8375,N_9890);
or U11136 (N_11136,N_8200,N_8029);
nand U11137 (N_11137,N_9994,N_9211);
or U11138 (N_11138,N_9951,N_8930);
or U11139 (N_11139,N_9524,N_9226);
or U11140 (N_11140,N_9651,N_8311);
nor U11141 (N_11141,N_8950,N_9811);
xor U11142 (N_11142,N_9699,N_9588);
nor U11143 (N_11143,N_8673,N_9707);
nor U11144 (N_11144,N_8922,N_8639);
nand U11145 (N_11145,N_8016,N_9245);
nor U11146 (N_11146,N_8634,N_8628);
and U11147 (N_11147,N_9626,N_8134);
xor U11148 (N_11148,N_8647,N_9069);
or U11149 (N_11149,N_8317,N_8550);
nand U11150 (N_11150,N_8265,N_9095);
nand U11151 (N_11151,N_8619,N_9824);
nand U11152 (N_11152,N_9418,N_8371);
or U11153 (N_11153,N_9668,N_8927);
or U11154 (N_11154,N_9556,N_9685);
nor U11155 (N_11155,N_8433,N_8655);
xnor U11156 (N_11156,N_8254,N_8011);
nor U11157 (N_11157,N_8019,N_8480);
and U11158 (N_11158,N_9050,N_9902);
nor U11159 (N_11159,N_9784,N_9271);
nand U11160 (N_11160,N_8647,N_9046);
and U11161 (N_11161,N_8328,N_8940);
nor U11162 (N_11162,N_8628,N_9973);
and U11163 (N_11163,N_8178,N_9877);
or U11164 (N_11164,N_9762,N_8992);
nor U11165 (N_11165,N_9050,N_9383);
nor U11166 (N_11166,N_9016,N_9690);
xor U11167 (N_11167,N_8326,N_8179);
nand U11168 (N_11168,N_8219,N_9973);
nor U11169 (N_11169,N_8034,N_8383);
and U11170 (N_11170,N_8327,N_8393);
or U11171 (N_11171,N_8609,N_8031);
nand U11172 (N_11172,N_9183,N_8382);
or U11173 (N_11173,N_9685,N_9425);
xnor U11174 (N_11174,N_9905,N_8304);
nor U11175 (N_11175,N_8602,N_9732);
nand U11176 (N_11176,N_9653,N_8721);
or U11177 (N_11177,N_8605,N_9687);
nand U11178 (N_11178,N_8985,N_9022);
nand U11179 (N_11179,N_8270,N_8249);
nor U11180 (N_11180,N_9987,N_9363);
and U11181 (N_11181,N_9576,N_9427);
and U11182 (N_11182,N_8354,N_9877);
nand U11183 (N_11183,N_8329,N_9794);
xor U11184 (N_11184,N_9235,N_9773);
and U11185 (N_11185,N_9275,N_8727);
xnor U11186 (N_11186,N_9655,N_8949);
or U11187 (N_11187,N_8103,N_8369);
or U11188 (N_11188,N_8251,N_8954);
or U11189 (N_11189,N_9866,N_9675);
or U11190 (N_11190,N_9357,N_8110);
or U11191 (N_11191,N_9981,N_9901);
and U11192 (N_11192,N_8689,N_8034);
nor U11193 (N_11193,N_9524,N_9160);
xnor U11194 (N_11194,N_9116,N_9456);
nor U11195 (N_11195,N_8221,N_8134);
xnor U11196 (N_11196,N_9233,N_9131);
nand U11197 (N_11197,N_8617,N_8785);
nor U11198 (N_11198,N_9019,N_9681);
or U11199 (N_11199,N_9323,N_8046);
nor U11200 (N_11200,N_9826,N_8055);
nor U11201 (N_11201,N_9909,N_9591);
nor U11202 (N_11202,N_9591,N_8340);
xnor U11203 (N_11203,N_9682,N_9677);
nand U11204 (N_11204,N_9625,N_9404);
nor U11205 (N_11205,N_9884,N_9015);
xnor U11206 (N_11206,N_8112,N_8676);
or U11207 (N_11207,N_9140,N_9489);
nand U11208 (N_11208,N_9419,N_8394);
or U11209 (N_11209,N_9198,N_9886);
nand U11210 (N_11210,N_9869,N_8755);
or U11211 (N_11211,N_9866,N_9924);
nor U11212 (N_11212,N_8053,N_9113);
nand U11213 (N_11213,N_8131,N_9143);
xnor U11214 (N_11214,N_9193,N_9579);
or U11215 (N_11215,N_9512,N_9430);
or U11216 (N_11216,N_9308,N_8788);
nand U11217 (N_11217,N_9542,N_9488);
or U11218 (N_11218,N_8268,N_9121);
or U11219 (N_11219,N_8729,N_9669);
and U11220 (N_11220,N_9403,N_9516);
and U11221 (N_11221,N_8589,N_8897);
xnor U11222 (N_11222,N_9099,N_9469);
and U11223 (N_11223,N_9600,N_8621);
nor U11224 (N_11224,N_8995,N_8700);
nor U11225 (N_11225,N_8579,N_8512);
or U11226 (N_11226,N_9678,N_8892);
and U11227 (N_11227,N_9584,N_9261);
nor U11228 (N_11228,N_8058,N_9759);
and U11229 (N_11229,N_9517,N_8266);
xor U11230 (N_11230,N_8234,N_9514);
or U11231 (N_11231,N_8565,N_8377);
nor U11232 (N_11232,N_8270,N_9644);
nor U11233 (N_11233,N_9085,N_8967);
nand U11234 (N_11234,N_9650,N_8081);
nor U11235 (N_11235,N_8684,N_8607);
nor U11236 (N_11236,N_9244,N_9820);
and U11237 (N_11237,N_8401,N_9389);
nor U11238 (N_11238,N_8761,N_9416);
nor U11239 (N_11239,N_8702,N_8284);
nand U11240 (N_11240,N_8666,N_8609);
xor U11241 (N_11241,N_9342,N_9021);
or U11242 (N_11242,N_8359,N_9640);
xnor U11243 (N_11243,N_8061,N_9234);
nand U11244 (N_11244,N_9936,N_8581);
and U11245 (N_11245,N_9347,N_9941);
nand U11246 (N_11246,N_9663,N_8830);
or U11247 (N_11247,N_8961,N_8462);
and U11248 (N_11248,N_8051,N_9517);
nor U11249 (N_11249,N_8027,N_8629);
nand U11250 (N_11250,N_9256,N_9918);
or U11251 (N_11251,N_8610,N_8812);
xnor U11252 (N_11252,N_9021,N_8344);
nor U11253 (N_11253,N_9623,N_8425);
nor U11254 (N_11254,N_8306,N_8230);
and U11255 (N_11255,N_9780,N_8605);
nor U11256 (N_11256,N_9020,N_8926);
nand U11257 (N_11257,N_9896,N_9188);
or U11258 (N_11258,N_9165,N_8135);
nor U11259 (N_11259,N_8252,N_9134);
and U11260 (N_11260,N_9265,N_9940);
nor U11261 (N_11261,N_8271,N_9825);
or U11262 (N_11262,N_9404,N_8012);
nand U11263 (N_11263,N_9984,N_9211);
xor U11264 (N_11264,N_8911,N_9996);
or U11265 (N_11265,N_9803,N_8217);
nor U11266 (N_11266,N_9038,N_9404);
nor U11267 (N_11267,N_8375,N_9648);
and U11268 (N_11268,N_8265,N_9919);
xor U11269 (N_11269,N_8618,N_8374);
and U11270 (N_11270,N_9586,N_8274);
or U11271 (N_11271,N_8906,N_9346);
and U11272 (N_11272,N_9433,N_8168);
xor U11273 (N_11273,N_8645,N_8482);
xor U11274 (N_11274,N_9403,N_8959);
xor U11275 (N_11275,N_8259,N_9859);
or U11276 (N_11276,N_8622,N_8282);
or U11277 (N_11277,N_9986,N_9969);
or U11278 (N_11278,N_8552,N_8632);
nand U11279 (N_11279,N_8476,N_8313);
and U11280 (N_11280,N_8496,N_9205);
xnor U11281 (N_11281,N_9020,N_9222);
or U11282 (N_11282,N_8846,N_9849);
xnor U11283 (N_11283,N_9705,N_8442);
xor U11284 (N_11284,N_8955,N_9944);
nor U11285 (N_11285,N_8788,N_8476);
xnor U11286 (N_11286,N_8739,N_8806);
xor U11287 (N_11287,N_9935,N_8792);
or U11288 (N_11288,N_8083,N_9603);
or U11289 (N_11289,N_8866,N_8177);
xnor U11290 (N_11290,N_9935,N_9415);
nand U11291 (N_11291,N_9153,N_9544);
xnor U11292 (N_11292,N_9099,N_9204);
nor U11293 (N_11293,N_9881,N_9918);
and U11294 (N_11294,N_8363,N_9739);
nor U11295 (N_11295,N_8544,N_9433);
xnor U11296 (N_11296,N_8528,N_9425);
nor U11297 (N_11297,N_8697,N_9055);
nand U11298 (N_11298,N_8441,N_9264);
xor U11299 (N_11299,N_8706,N_9889);
or U11300 (N_11300,N_8282,N_8902);
and U11301 (N_11301,N_9358,N_9079);
and U11302 (N_11302,N_8059,N_9554);
or U11303 (N_11303,N_8399,N_8366);
xor U11304 (N_11304,N_9392,N_8673);
nand U11305 (N_11305,N_8361,N_8883);
nor U11306 (N_11306,N_8506,N_9845);
xnor U11307 (N_11307,N_9054,N_8229);
and U11308 (N_11308,N_9976,N_8605);
and U11309 (N_11309,N_8641,N_8350);
and U11310 (N_11310,N_9263,N_8953);
or U11311 (N_11311,N_9020,N_8399);
and U11312 (N_11312,N_8224,N_9114);
and U11313 (N_11313,N_8597,N_8756);
xor U11314 (N_11314,N_9799,N_9788);
nor U11315 (N_11315,N_8035,N_8686);
nand U11316 (N_11316,N_8701,N_9782);
nand U11317 (N_11317,N_8829,N_9553);
nor U11318 (N_11318,N_9803,N_9000);
nand U11319 (N_11319,N_9979,N_9329);
xor U11320 (N_11320,N_9455,N_8522);
nor U11321 (N_11321,N_8803,N_9280);
nor U11322 (N_11322,N_8429,N_8911);
nand U11323 (N_11323,N_8449,N_9566);
and U11324 (N_11324,N_9092,N_9745);
nand U11325 (N_11325,N_8899,N_8422);
and U11326 (N_11326,N_9404,N_9957);
or U11327 (N_11327,N_9498,N_8692);
nor U11328 (N_11328,N_9070,N_8244);
nor U11329 (N_11329,N_9392,N_8134);
and U11330 (N_11330,N_8870,N_9493);
nor U11331 (N_11331,N_9319,N_8332);
nor U11332 (N_11332,N_8482,N_8226);
nor U11333 (N_11333,N_8932,N_8769);
or U11334 (N_11334,N_8143,N_8011);
nand U11335 (N_11335,N_9983,N_8552);
nand U11336 (N_11336,N_9600,N_9546);
nand U11337 (N_11337,N_9190,N_8848);
or U11338 (N_11338,N_9213,N_8709);
xnor U11339 (N_11339,N_9528,N_8514);
and U11340 (N_11340,N_8707,N_8061);
nor U11341 (N_11341,N_8583,N_8287);
nor U11342 (N_11342,N_9897,N_8411);
and U11343 (N_11343,N_9448,N_9954);
xnor U11344 (N_11344,N_8609,N_9912);
nor U11345 (N_11345,N_8240,N_8572);
or U11346 (N_11346,N_9491,N_8297);
nor U11347 (N_11347,N_8688,N_8477);
or U11348 (N_11348,N_8885,N_8579);
nor U11349 (N_11349,N_9289,N_9243);
or U11350 (N_11350,N_8270,N_9421);
nor U11351 (N_11351,N_8054,N_9729);
and U11352 (N_11352,N_8482,N_9919);
and U11353 (N_11353,N_9543,N_8954);
nand U11354 (N_11354,N_8377,N_9094);
nor U11355 (N_11355,N_9446,N_9823);
or U11356 (N_11356,N_8617,N_8520);
and U11357 (N_11357,N_8083,N_8691);
or U11358 (N_11358,N_9275,N_8272);
xor U11359 (N_11359,N_8493,N_9043);
nor U11360 (N_11360,N_9991,N_8022);
and U11361 (N_11361,N_8513,N_9808);
nor U11362 (N_11362,N_9703,N_8869);
nand U11363 (N_11363,N_8758,N_8324);
and U11364 (N_11364,N_9349,N_8137);
nand U11365 (N_11365,N_9173,N_8172);
and U11366 (N_11366,N_9457,N_9269);
nand U11367 (N_11367,N_9365,N_9147);
or U11368 (N_11368,N_8193,N_9052);
xor U11369 (N_11369,N_9196,N_9310);
and U11370 (N_11370,N_9558,N_8839);
xor U11371 (N_11371,N_9921,N_8925);
xnor U11372 (N_11372,N_8419,N_8475);
nor U11373 (N_11373,N_8292,N_8533);
nor U11374 (N_11374,N_9254,N_8186);
nand U11375 (N_11375,N_9655,N_8304);
and U11376 (N_11376,N_8916,N_8996);
or U11377 (N_11377,N_8202,N_9988);
and U11378 (N_11378,N_9396,N_8198);
and U11379 (N_11379,N_9235,N_9579);
nor U11380 (N_11380,N_9234,N_9674);
nand U11381 (N_11381,N_8446,N_8630);
and U11382 (N_11382,N_8139,N_8740);
or U11383 (N_11383,N_9749,N_9060);
xor U11384 (N_11384,N_8813,N_8419);
or U11385 (N_11385,N_9943,N_8559);
nand U11386 (N_11386,N_9891,N_8170);
nand U11387 (N_11387,N_8511,N_9189);
xor U11388 (N_11388,N_8561,N_9631);
nor U11389 (N_11389,N_8967,N_8935);
nor U11390 (N_11390,N_8310,N_9624);
nand U11391 (N_11391,N_8011,N_8804);
nor U11392 (N_11392,N_8125,N_9915);
nand U11393 (N_11393,N_8702,N_9608);
or U11394 (N_11394,N_8180,N_8685);
and U11395 (N_11395,N_8447,N_8713);
nor U11396 (N_11396,N_8155,N_8420);
xnor U11397 (N_11397,N_8925,N_9559);
nor U11398 (N_11398,N_8321,N_8283);
or U11399 (N_11399,N_9522,N_8082);
nor U11400 (N_11400,N_9439,N_9097);
xor U11401 (N_11401,N_9394,N_8166);
xor U11402 (N_11402,N_9899,N_8379);
xor U11403 (N_11403,N_8138,N_9821);
and U11404 (N_11404,N_8566,N_8837);
nand U11405 (N_11405,N_9159,N_8698);
and U11406 (N_11406,N_9839,N_9083);
nand U11407 (N_11407,N_9463,N_9121);
or U11408 (N_11408,N_9980,N_9566);
nand U11409 (N_11409,N_8504,N_8249);
and U11410 (N_11410,N_8908,N_8433);
xor U11411 (N_11411,N_8427,N_8197);
xor U11412 (N_11412,N_9620,N_8883);
xnor U11413 (N_11413,N_9602,N_8817);
xnor U11414 (N_11414,N_8187,N_9759);
nand U11415 (N_11415,N_8577,N_8431);
nand U11416 (N_11416,N_9990,N_8570);
nor U11417 (N_11417,N_9183,N_8535);
nor U11418 (N_11418,N_9883,N_9624);
nand U11419 (N_11419,N_9700,N_9391);
xnor U11420 (N_11420,N_9275,N_8414);
or U11421 (N_11421,N_9404,N_8419);
xnor U11422 (N_11422,N_9600,N_8868);
and U11423 (N_11423,N_8602,N_9880);
nor U11424 (N_11424,N_8138,N_8063);
nor U11425 (N_11425,N_8595,N_8499);
and U11426 (N_11426,N_8190,N_9335);
xor U11427 (N_11427,N_8807,N_9360);
xnor U11428 (N_11428,N_9227,N_9598);
nand U11429 (N_11429,N_8261,N_8488);
nor U11430 (N_11430,N_9174,N_9160);
and U11431 (N_11431,N_9446,N_8746);
nor U11432 (N_11432,N_8921,N_8569);
or U11433 (N_11433,N_8941,N_9493);
nand U11434 (N_11434,N_9910,N_8638);
nor U11435 (N_11435,N_8969,N_8711);
or U11436 (N_11436,N_8037,N_9325);
nor U11437 (N_11437,N_9034,N_9286);
or U11438 (N_11438,N_9483,N_9204);
and U11439 (N_11439,N_8270,N_8945);
or U11440 (N_11440,N_9349,N_9287);
and U11441 (N_11441,N_8621,N_8273);
xor U11442 (N_11442,N_9711,N_8796);
and U11443 (N_11443,N_9252,N_9043);
or U11444 (N_11444,N_8340,N_9991);
xor U11445 (N_11445,N_9544,N_9028);
and U11446 (N_11446,N_8407,N_9577);
and U11447 (N_11447,N_9760,N_9569);
xnor U11448 (N_11448,N_9723,N_8869);
nor U11449 (N_11449,N_9773,N_9914);
nand U11450 (N_11450,N_9020,N_9649);
or U11451 (N_11451,N_8090,N_8139);
or U11452 (N_11452,N_8548,N_8458);
nor U11453 (N_11453,N_8689,N_8254);
nand U11454 (N_11454,N_9776,N_8614);
or U11455 (N_11455,N_9823,N_9121);
or U11456 (N_11456,N_8060,N_9983);
xnor U11457 (N_11457,N_9998,N_9962);
or U11458 (N_11458,N_9374,N_8540);
nand U11459 (N_11459,N_9902,N_9525);
nand U11460 (N_11460,N_9587,N_9423);
and U11461 (N_11461,N_8229,N_9532);
nor U11462 (N_11462,N_9731,N_9748);
or U11463 (N_11463,N_8496,N_9557);
or U11464 (N_11464,N_8608,N_8072);
and U11465 (N_11465,N_8606,N_8420);
and U11466 (N_11466,N_8036,N_9524);
nand U11467 (N_11467,N_9378,N_8593);
nand U11468 (N_11468,N_8474,N_9333);
xnor U11469 (N_11469,N_9382,N_8092);
or U11470 (N_11470,N_9098,N_9578);
xnor U11471 (N_11471,N_9926,N_8593);
xor U11472 (N_11472,N_9104,N_9929);
or U11473 (N_11473,N_8348,N_9938);
nand U11474 (N_11474,N_9070,N_9987);
xor U11475 (N_11475,N_8377,N_8350);
and U11476 (N_11476,N_9108,N_8674);
nand U11477 (N_11477,N_8795,N_8410);
nor U11478 (N_11478,N_8411,N_8927);
xor U11479 (N_11479,N_9079,N_9975);
or U11480 (N_11480,N_9956,N_8335);
nand U11481 (N_11481,N_8029,N_8900);
nand U11482 (N_11482,N_8909,N_9258);
or U11483 (N_11483,N_8409,N_8626);
nor U11484 (N_11484,N_8479,N_8810);
or U11485 (N_11485,N_9964,N_8140);
nor U11486 (N_11486,N_8135,N_9765);
xor U11487 (N_11487,N_8489,N_9732);
nor U11488 (N_11488,N_9476,N_9444);
and U11489 (N_11489,N_8016,N_8839);
xnor U11490 (N_11490,N_9652,N_8811);
or U11491 (N_11491,N_9325,N_8149);
nor U11492 (N_11492,N_9664,N_8287);
or U11493 (N_11493,N_9520,N_8038);
or U11494 (N_11494,N_8095,N_9977);
and U11495 (N_11495,N_8386,N_8855);
xnor U11496 (N_11496,N_9515,N_9909);
nand U11497 (N_11497,N_9016,N_8676);
nor U11498 (N_11498,N_9425,N_9090);
nand U11499 (N_11499,N_9456,N_9628);
nand U11500 (N_11500,N_9759,N_9819);
nor U11501 (N_11501,N_9724,N_9126);
xor U11502 (N_11502,N_9754,N_8478);
or U11503 (N_11503,N_9355,N_9519);
xor U11504 (N_11504,N_9961,N_8679);
nor U11505 (N_11505,N_9488,N_8713);
and U11506 (N_11506,N_9560,N_9973);
nand U11507 (N_11507,N_8945,N_9577);
nor U11508 (N_11508,N_8858,N_9031);
or U11509 (N_11509,N_9949,N_8815);
or U11510 (N_11510,N_9720,N_9848);
or U11511 (N_11511,N_9467,N_8892);
and U11512 (N_11512,N_9716,N_8537);
xor U11513 (N_11513,N_9656,N_9823);
and U11514 (N_11514,N_8919,N_8600);
or U11515 (N_11515,N_8520,N_9978);
and U11516 (N_11516,N_8642,N_9244);
xnor U11517 (N_11517,N_9974,N_8891);
xnor U11518 (N_11518,N_9902,N_9472);
and U11519 (N_11519,N_8238,N_8345);
and U11520 (N_11520,N_8212,N_8832);
or U11521 (N_11521,N_9720,N_9344);
or U11522 (N_11522,N_8276,N_8653);
and U11523 (N_11523,N_9952,N_9198);
nand U11524 (N_11524,N_8742,N_9595);
nand U11525 (N_11525,N_9253,N_8657);
xnor U11526 (N_11526,N_9077,N_9557);
or U11527 (N_11527,N_8902,N_9607);
nor U11528 (N_11528,N_9749,N_8495);
nand U11529 (N_11529,N_9523,N_8372);
nor U11530 (N_11530,N_8149,N_9937);
or U11531 (N_11531,N_9938,N_8414);
xnor U11532 (N_11532,N_9404,N_9215);
and U11533 (N_11533,N_8405,N_8354);
xnor U11534 (N_11534,N_9788,N_9846);
or U11535 (N_11535,N_8592,N_8582);
and U11536 (N_11536,N_8838,N_8060);
xnor U11537 (N_11537,N_9616,N_9560);
xnor U11538 (N_11538,N_9511,N_8522);
and U11539 (N_11539,N_8880,N_9193);
nand U11540 (N_11540,N_9218,N_8450);
nor U11541 (N_11541,N_8122,N_9630);
nor U11542 (N_11542,N_9625,N_9958);
xnor U11543 (N_11543,N_9917,N_9126);
or U11544 (N_11544,N_8054,N_9074);
and U11545 (N_11545,N_8160,N_8954);
xnor U11546 (N_11546,N_9436,N_9698);
xor U11547 (N_11547,N_9755,N_9047);
and U11548 (N_11548,N_8670,N_9685);
or U11549 (N_11549,N_8207,N_9133);
nand U11550 (N_11550,N_8516,N_9261);
or U11551 (N_11551,N_9969,N_8268);
or U11552 (N_11552,N_9539,N_8994);
or U11553 (N_11553,N_8425,N_8483);
nor U11554 (N_11554,N_9246,N_8808);
and U11555 (N_11555,N_8876,N_9179);
nand U11556 (N_11556,N_9000,N_9615);
and U11557 (N_11557,N_8679,N_8103);
or U11558 (N_11558,N_9472,N_9855);
or U11559 (N_11559,N_8064,N_9078);
and U11560 (N_11560,N_8583,N_8680);
or U11561 (N_11561,N_8238,N_9004);
and U11562 (N_11562,N_8721,N_8459);
nand U11563 (N_11563,N_9319,N_9834);
nor U11564 (N_11564,N_8168,N_9092);
xor U11565 (N_11565,N_9006,N_9864);
nand U11566 (N_11566,N_8285,N_8623);
and U11567 (N_11567,N_8651,N_9790);
xnor U11568 (N_11568,N_8244,N_8909);
nand U11569 (N_11569,N_8740,N_8487);
and U11570 (N_11570,N_9151,N_9972);
or U11571 (N_11571,N_8638,N_9938);
and U11572 (N_11572,N_9697,N_8944);
xor U11573 (N_11573,N_8243,N_9505);
xor U11574 (N_11574,N_9713,N_8003);
or U11575 (N_11575,N_8960,N_8955);
or U11576 (N_11576,N_9373,N_8313);
xor U11577 (N_11577,N_9170,N_9869);
or U11578 (N_11578,N_8737,N_9697);
and U11579 (N_11579,N_8465,N_9473);
xnor U11580 (N_11580,N_8674,N_9282);
or U11581 (N_11581,N_9739,N_8642);
or U11582 (N_11582,N_8234,N_8010);
xnor U11583 (N_11583,N_9201,N_8620);
and U11584 (N_11584,N_9178,N_8790);
or U11585 (N_11585,N_9443,N_8120);
or U11586 (N_11586,N_9992,N_9199);
nor U11587 (N_11587,N_8562,N_8953);
nor U11588 (N_11588,N_8509,N_9508);
and U11589 (N_11589,N_8629,N_8805);
or U11590 (N_11590,N_9067,N_9962);
nand U11591 (N_11591,N_9883,N_9220);
or U11592 (N_11592,N_8526,N_8218);
or U11593 (N_11593,N_8641,N_8144);
and U11594 (N_11594,N_8145,N_9564);
nand U11595 (N_11595,N_9419,N_8996);
nand U11596 (N_11596,N_8959,N_8983);
nor U11597 (N_11597,N_8389,N_9208);
or U11598 (N_11598,N_9272,N_9333);
or U11599 (N_11599,N_8624,N_9837);
nand U11600 (N_11600,N_9598,N_8292);
nor U11601 (N_11601,N_8713,N_8508);
xnor U11602 (N_11602,N_8883,N_8939);
or U11603 (N_11603,N_8589,N_9990);
nor U11604 (N_11604,N_9900,N_9138);
nor U11605 (N_11605,N_8642,N_9357);
nand U11606 (N_11606,N_8528,N_9113);
or U11607 (N_11607,N_8642,N_8389);
nor U11608 (N_11608,N_8389,N_9171);
xnor U11609 (N_11609,N_8608,N_8448);
and U11610 (N_11610,N_8333,N_8508);
nor U11611 (N_11611,N_8666,N_8579);
or U11612 (N_11612,N_8284,N_9353);
nor U11613 (N_11613,N_8813,N_8632);
nor U11614 (N_11614,N_8479,N_9834);
nand U11615 (N_11615,N_9304,N_9804);
nor U11616 (N_11616,N_9058,N_9354);
nor U11617 (N_11617,N_8966,N_8893);
nand U11618 (N_11618,N_9036,N_8049);
nor U11619 (N_11619,N_8196,N_9780);
and U11620 (N_11620,N_8294,N_9538);
and U11621 (N_11621,N_8387,N_8096);
and U11622 (N_11622,N_8542,N_8557);
nand U11623 (N_11623,N_9485,N_9319);
and U11624 (N_11624,N_9176,N_8744);
and U11625 (N_11625,N_9650,N_8901);
nand U11626 (N_11626,N_9018,N_8922);
xor U11627 (N_11627,N_8569,N_8142);
or U11628 (N_11628,N_8048,N_9475);
or U11629 (N_11629,N_9159,N_8749);
nand U11630 (N_11630,N_8732,N_9146);
nand U11631 (N_11631,N_8101,N_8470);
nand U11632 (N_11632,N_8203,N_9677);
nand U11633 (N_11633,N_8317,N_8413);
nand U11634 (N_11634,N_8175,N_8199);
xor U11635 (N_11635,N_8260,N_9780);
nand U11636 (N_11636,N_9075,N_9173);
xnor U11637 (N_11637,N_8133,N_9870);
xor U11638 (N_11638,N_9854,N_9010);
xor U11639 (N_11639,N_8911,N_8912);
or U11640 (N_11640,N_9365,N_8809);
nor U11641 (N_11641,N_8888,N_9041);
xnor U11642 (N_11642,N_9127,N_8824);
xnor U11643 (N_11643,N_8912,N_8897);
nand U11644 (N_11644,N_8578,N_9925);
nor U11645 (N_11645,N_9315,N_8037);
xor U11646 (N_11646,N_8935,N_8681);
and U11647 (N_11647,N_8757,N_8856);
nor U11648 (N_11648,N_9821,N_8420);
and U11649 (N_11649,N_8253,N_8446);
nand U11650 (N_11650,N_8928,N_9306);
nand U11651 (N_11651,N_8144,N_8663);
nor U11652 (N_11652,N_8017,N_8115);
and U11653 (N_11653,N_9932,N_9094);
nand U11654 (N_11654,N_8655,N_9396);
or U11655 (N_11655,N_8928,N_8407);
nor U11656 (N_11656,N_8661,N_9960);
and U11657 (N_11657,N_8275,N_8501);
or U11658 (N_11658,N_8901,N_8019);
and U11659 (N_11659,N_9085,N_9678);
or U11660 (N_11660,N_8893,N_8371);
and U11661 (N_11661,N_9765,N_8216);
and U11662 (N_11662,N_8560,N_9866);
and U11663 (N_11663,N_8118,N_9684);
and U11664 (N_11664,N_8428,N_9222);
and U11665 (N_11665,N_9961,N_9218);
or U11666 (N_11666,N_9144,N_9052);
or U11667 (N_11667,N_8408,N_9454);
and U11668 (N_11668,N_8905,N_8948);
and U11669 (N_11669,N_8839,N_8745);
and U11670 (N_11670,N_9930,N_8650);
or U11671 (N_11671,N_9760,N_8052);
nor U11672 (N_11672,N_8054,N_8081);
or U11673 (N_11673,N_8960,N_9228);
xnor U11674 (N_11674,N_8307,N_9975);
or U11675 (N_11675,N_9511,N_8206);
or U11676 (N_11676,N_8633,N_9438);
and U11677 (N_11677,N_9236,N_9700);
nor U11678 (N_11678,N_9878,N_9762);
xnor U11679 (N_11679,N_8427,N_9044);
or U11680 (N_11680,N_9222,N_8610);
xor U11681 (N_11681,N_9027,N_9620);
or U11682 (N_11682,N_8993,N_8775);
and U11683 (N_11683,N_9091,N_9544);
xor U11684 (N_11684,N_9352,N_8781);
and U11685 (N_11685,N_9308,N_8522);
xor U11686 (N_11686,N_8270,N_9373);
nand U11687 (N_11687,N_8932,N_9326);
xnor U11688 (N_11688,N_8594,N_8816);
or U11689 (N_11689,N_9651,N_9183);
nor U11690 (N_11690,N_8329,N_9612);
and U11691 (N_11691,N_8584,N_8646);
nor U11692 (N_11692,N_9640,N_8217);
or U11693 (N_11693,N_9448,N_9281);
xnor U11694 (N_11694,N_8612,N_9598);
nor U11695 (N_11695,N_8350,N_9077);
or U11696 (N_11696,N_9564,N_9740);
and U11697 (N_11697,N_9365,N_8333);
nor U11698 (N_11698,N_9408,N_9924);
nand U11699 (N_11699,N_8588,N_8683);
and U11700 (N_11700,N_8093,N_8092);
nor U11701 (N_11701,N_8283,N_9218);
xnor U11702 (N_11702,N_8059,N_9349);
nand U11703 (N_11703,N_8366,N_9221);
nand U11704 (N_11704,N_9907,N_9673);
nor U11705 (N_11705,N_8070,N_9410);
xnor U11706 (N_11706,N_8129,N_8915);
nor U11707 (N_11707,N_8147,N_8809);
nor U11708 (N_11708,N_9869,N_9187);
xnor U11709 (N_11709,N_9149,N_8934);
and U11710 (N_11710,N_8835,N_8272);
or U11711 (N_11711,N_8153,N_9690);
nand U11712 (N_11712,N_9181,N_9854);
nand U11713 (N_11713,N_9867,N_9289);
xor U11714 (N_11714,N_9950,N_9750);
xor U11715 (N_11715,N_8598,N_8993);
and U11716 (N_11716,N_9038,N_9748);
or U11717 (N_11717,N_9174,N_8610);
xor U11718 (N_11718,N_9530,N_9886);
nor U11719 (N_11719,N_9860,N_9550);
and U11720 (N_11720,N_8772,N_9215);
xor U11721 (N_11721,N_9157,N_8874);
and U11722 (N_11722,N_9573,N_9751);
or U11723 (N_11723,N_9872,N_9142);
and U11724 (N_11724,N_8443,N_9854);
nand U11725 (N_11725,N_9962,N_9161);
or U11726 (N_11726,N_9196,N_9735);
nand U11727 (N_11727,N_8943,N_9675);
or U11728 (N_11728,N_8422,N_9468);
and U11729 (N_11729,N_8834,N_8447);
nor U11730 (N_11730,N_8705,N_9813);
nor U11731 (N_11731,N_8823,N_8138);
or U11732 (N_11732,N_9360,N_8714);
and U11733 (N_11733,N_9735,N_8444);
or U11734 (N_11734,N_8344,N_8690);
nand U11735 (N_11735,N_8510,N_9289);
nor U11736 (N_11736,N_9249,N_8941);
xor U11737 (N_11737,N_9732,N_8431);
nand U11738 (N_11738,N_8556,N_8752);
or U11739 (N_11739,N_8059,N_9195);
nor U11740 (N_11740,N_8939,N_8916);
nand U11741 (N_11741,N_9965,N_9898);
and U11742 (N_11742,N_8350,N_8788);
xnor U11743 (N_11743,N_9798,N_9967);
or U11744 (N_11744,N_8979,N_8838);
nor U11745 (N_11745,N_8518,N_9563);
and U11746 (N_11746,N_9590,N_8454);
nand U11747 (N_11747,N_9612,N_8556);
xor U11748 (N_11748,N_9539,N_8757);
nor U11749 (N_11749,N_9162,N_8260);
nor U11750 (N_11750,N_9965,N_8488);
nor U11751 (N_11751,N_9573,N_9832);
and U11752 (N_11752,N_8680,N_9467);
and U11753 (N_11753,N_8666,N_9232);
nor U11754 (N_11754,N_8292,N_9633);
nand U11755 (N_11755,N_9033,N_8836);
and U11756 (N_11756,N_8362,N_8959);
and U11757 (N_11757,N_9267,N_9270);
nor U11758 (N_11758,N_8422,N_8640);
and U11759 (N_11759,N_9358,N_9883);
xor U11760 (N_11760,N_8850,N_9307);
nand U11761 (N_11761,N_8757,N_9948);
and U11762 (N_11762,N_9278,N_8889);
nor U11763 (N_11763,N_8287,N_8082);
or U11764 (N_11764,N_9645,N_8363);
xnor U11765 (N_11765,N_9570,N_9964);
or U11766 (N_11766,N_8425,N_9136);
nand U11767 (N_11767,N_9813,N_8925);
xor U11768 (N_11768,N_8601,N_9970);
nor U11769 (N_11769,N_9512,N_9501);
nand U11770 (N_11770,N_8323,N_8449);
nand U11771 (N_11771,N_9008,N_8035);
xnor U11772 (N_11772,N_9158,N_8606);
and U11773 (N_11773,N_9133,N_8236);
xor U11774 (N_11774,N_8625,N_9730);
and U11775 (N_11775,N_9881,N_8849);
xor U11776 (N_11776,N_9566,N_9836);
nand U11777 (N_11777,N_9196,N_8970);
and U11778 (N_11778,N_8586,N_8114);
and U11779 (N_11779,N_8033,N_9012);
and U11780 (N_11780,N_9239,N_9830);
nor U11781 (N_11781,N_8058,N_8236);
or U11782 (N_11782,N_8233,N_9450);
xnor U11783 (N_11783,N_9154,N_9930);
and U11784 (N_11784,N_8913,N_8853);
and U11785 (N_11785,N_8389,N_8743);
xor U11786 (N_11786,N_8791,N_9184);
xnor U11787 (N_11787,N_8699,N_9706);
xor U11788 (N_11788,N_8783,N_9279);
nand U11789 (N_11789,N_9179,N_9733);
and U11790 (N_11790,N_8006,N_8317);
nor U11791 (N_11791,N_8387,N_8459);
xnor U11792 (N_11792,N_8221,N_9371);
or U11793 (N_11793,N_8575,N_9308);
and U11794 (N_11794,N_9486,N_8910);
nor U11795 (N_11795,N_9107,N_8565);
nand U11796 (N_11796,N_8342,N_8246);
or U11797 (N_11797,N_8634,N_9180);
nor U11798 (N_11798,N_9147,N_9881);
xnor U11799 (N_11799,N_8064,N_9607);
xor U11800 (N_11800,N_9127,N_8869);
xor U11801 (N_11801,N_9635,N_9796);
nor U11802 (N_11802,N_8350,N_8145);
and U11803 (N_11803,N_8614,N_8873);
and U11804 (N_11804,N_9282,N_9661);
xnor U11805 (N_11805,N_8194,N_9983);
or U11806 (N_11806,N_9908,N_9667);
nor U11807 (N_11807,N_9026,N_9911);
or U11808 (N_11808,N_9896,N_8709);
and U11809 (N_11809,N_8256,N_8594);
nor U11810 (N_11810,N_8375,N_8990);
and U11811 (N_11811,N_9330,N_9514);
xor U11812 (N_11812,N_9092,N_9241);
and U11813 (N_11813,N_9382,N_9080);
nor U11814 (N_11814,N_8111,N_8599);
nor U11815 (N_11815,N_8190,N_8760);
and U11816 (N_11816,N_8664,N_9448);
xnor U11817 (N_11817,N_8355,N_8439);
or U11818 (N_11818,N_9027,N_8384);
and U11819 (N_11819,N_9407,N_9516);
xor U11820 (N_11820,N_8330,N_9409);
or U11821 (N_11821,N_8127,N_8182);
nor U11822 (N_11822,N_9079,N_9406);
nor U11823 (N_11823,N_8270,N_8502);
xor U11824 (N_11824,N_8033,N_9210);
or U11825 (N_11825,N_9769,N_8231);
xnor U11826 (N_11826,N_9106,N_8072);
xor U11827 (N_11827,N_8847,N_9614);
nand U11828 (N_11828,N_9417,N_9967);
xor U11829 (N_11829,N_8803,N_9891);
or U11830 (N_11830,N_9557,N_9922);
or U11831 (N_11831,N_9934,N_8669);
nand U11832 (N_11832,N_9044,N_9048);
and U11833 (N_11833,N_8085,N_8716);
and U11834 (N_11834,N_9131,N_9106);
xnor U11835 (N_11835,N_9395,N_8102);
and U11836 (N_11836,N_8834,N_9166);
or U11837 (N_11837,N_8896,N_9504);
nor U11838 (N_11838,N_8967,N_9239);
and U11839 (N_11839,N_9505,N_9879);
and U11840 (N_11840,N_8480,N_9537);
or U11841 (N_11841,N_8985,N_8408);
nand U11842 (N_11842,N_8945,N_9999);
nor U11843 (N_11843,N_8834,N_9159);
xor U11844 (N_11844,N_8922,N_8634);
nor U11845 (N_11845,N_8795,N_8677);
or U11846 (N_11846,N_8667,N_9014);
or U11847 (N_11847,N_8552,N_9809);
nor U11848 (N_11848,N_9243,N_8881);
xor U11849 (N_11849,N_9687,N_8504);
nand U11850 (N_11850,N_8657,N_8577);
xor U11851 (N_11851,N_8351,N_9019);
nand U11852 (N_11852,N_8137,N_8657);
nand U11853 (N_11853,N_9880,N_8801);
and U11854 (N_11854,N_9567,N_9268);
xor U11855 (N_11855,N_9619,N_9861);
nor U11856 (N_11856,N_8438,N_8219);
nor U11857 (N_11857,N_9919,N_9555);
xor U11858 (N_11858,N_8039,N_9436);
or U11859 (N_11859,N_9416,N_9356);
xnor U11860 (N_11860,N_9208,N_9188);
nor U11861 (N_11861,N_8304,N_8932);
nand U11862 (N_11862,N_9840,N_9105);
xnor U11863 (N_11863,N_9258,N_9084);
nand U11864 (N_11864,N_8146,N_9865);
nand U11865 (N_11865,N_9650,N_8925);
nor U11866 (N_11866,N_8085,N_8961);
and U11867 (N_11867,N_9912,N_8473);
nand U11868 (N_11868,N_9700,N_9131);
and U11869 (N_11869,N_8961,N_8542);
or U11870 (N_11870,N_9773,N_8463);
xor U11871 (N_11871,N_8342,N_9223);
and U11872 (N_11872,N_8113,N_8953);
xnor U11873 (N_11873,N_8859,N_9616);
xor U11874 (N_11874,N_9345,N_8608);
nand U11875 (N_11875,N_9485,N_9338);
xor U11876 (N_11876,N_8898,N_9477);
or U11877 (N_11877,N_9545,N_9312);
nand U11878 (N_11878,N_9358,N_8386);
and U11879 (N_11879,N_9606,N_8086);
nor U11880 (N_11880,N_8903,N_9818);
and U11881 (N_11881,N_9242,N_8204);
xor U11882 (N_11882,N_9918,N_8908);
or U11883 (N_11883,N_9026,N_9755);
and U11884 (N_11884,N_9645,N_8832);
and U11885 (N_11885,N_8884,N_9988);
nand U11886 (N_11886,N_9007,N_8065);
or U11887 (N_11887,N_8826,N_9902);
nor U11888 (N_11888,N_8937,N_9994);
nand U11889 (N_11889,N_9291,N_9779);
nor U11890 (N_11890,N_9184,N_9557);
nor U11891 (N_11891,N_9485,N_8578);
nand U11892 (N_11892,N_9936,N_9461);
or U11893 (N_11893,N_9152,N_8090);
xor U11894 (N_11894,N_9486,N_8694);
or U11895 (N_11895,N_8621,N_8175);
or U11896 (N_11896,N_8705,N_8984);
or U11897 (N_11897,N_9430,N_9486);
xor U11898 (N_11898,N_8989,N_8437);
nor U11899 (N_11899,N_8013,N_8433);
nor U11900 (N_11900,N_8550,N_9587);
nand U11901 (N_11901,N_8784,N_8887);
or U11902 (N_11902,N_9184,N_8423);
or U11903 (N_11903,N_8681,N_9178);
or U11904 (N_11904,N_8621,N_9840);
xnor U11905 (N_11905,N_9177,N_8175);
or U11906 (N_11906,N_9631,N_8290);
xor U11907 (N_11907,N_8740,N_8805);
or U11908 (N_11908,N_9111,N_9690);
xnor U11909 (N_11909,N_9396,N_9300);
nand U11910 (N_11910,N_8784,N_9144);
xnor U11911 (N_11911,N_8330,N_9928);
xor U11912 (N_11912,N_8148,N_8464);
nand U11913 (N_11913,N_9597,N_8469);
and U11914 (N_11914,N_8659,N_8888);
xor U11915 (N_11915,N_8405,N_9381);
and U11916 (N_11916,N_9837,N_8239);
xnor U11917 (N_11917,N_9858,N_8491);
nand U11918 (N_11918,N_8130,N_8108);
xnor U11919 (N_11919,N_8255,N_9992);
and U11920 (N_11920,N_9930,N_9885);
and U11921 (N_11921,N_8782,N_9042);
or U11922 (N_11922,N_9346,N_8258);
or U11923 (N_11923,N_8593,N_8439);
xor U11924 (N_11924,N_9192,N_8665);
or U11925 (N_11925,N_9346,N_8646);
or U11926 (N_11926,N_8818,N_9653);
nor U11927 (N_11927,N_8413,N_8488);
nor U11928 (N_11928,N_9571,N_8540);
nor U11929 (N_11929,N_9023,N_8651);
or U11930 (N_11930,N_8392,N_9220);
and U11931 (N_11931,N_8174,N_9363);
xnor U11932 (N_11932,N_9200,N_8070);
or U11933 (N_11933,N_8548,N_9326);
xor U11934 (N_11934,N_8717,N_8212);
and U11935 (N_11935,N_9954,N_9701);
and U11936 (N_11936,N_8457,N_8907);
or U11937 (N_11937,N_9718,N_8338);
xor U11938 (N_11938,N_8820,N_9151);
nor U11939 (N_11939,N_9576,N_8861);
nor U11940 (N_11940,N_8015,N_8344);
or U11941 (N_11941,N_8179,N_8690);
nand U11942 (N_11942,N_9357,N_9257);
xnor U11943 (N_11943,N_8807,N_8106);
and U11944 (N_11944,N_8887,N_9255);
and U11945 (N_11945,N_8177,N_9331);
nand U11946 (N_11946,N_9283,N_8377);
or U11947 (N_11947,N_9173,N_8402);
and U11948 (N_11948,N_9116,N_9252);
nor U11949 (N_11949,N_9563,N_9965);
or U11950 (N_11950,N_8880,N_8709);
or U11951 (N_11951,N_9821,N_8003);
or U11952 (N_11952,N_8030,N_9348);
nand U11953 (N_11953,N_8336,N_9730);
or U11954 (N_11954,N_9264,N_9439);
and U11955 (N_11955,N_9117,N_9359);
xnor U11956 (N_11956,N_8876,N_8303);
xnor U11957 (N_11957,N_9244,N_8131);
nor U11958 (N_11958,N_8363,N_8659);
nor U11959 (N_11959,N_9627,N_9722);
xnor U11960 (N_11960,N_9709,N_8009);
or U11961 (N_11961,N_8548,N_9900);
and U11962 (N_11962,N_8828,N_9214);
xor U11963 (N_11963,N_8724,N_9326);
and U11964 (N_11964,N_8017,N_9735);
xnor U11965 (N_11965,N_9943,N_8932);
nor U11966 (N_11966,N_8101,N_9389);
xnor U11967 (N_11967,N_8061,N_9678);
or U11968 (N_11968,N_8326,N_8966);
and U11969 (N_11969,N_8504,N_8225);
or U11970 (N_11970,N_8163,N_8463);
nor U11971 (N_11971,N_9587,N_8242);
nor U11972 (N_11972,N_9491,N_9999);
nor U11973 (N_11973,N_8047,N_8213);
nor U11974 (N_11974,N_8861,N_9906);
nand U11975 (N_11975,N_9350,N_8064);
or U11976 (N_11976,N_8108,N_8899);
nand U11977 (N_11977,N_9150,N_8153);
or U11978 (N_11978,N_8250,N_9168);
and U11979 (N_11979,N_9465,N_8493);
xor U11980 (N_11980,N_8817,N_8398);
and U11981 (N_11981,N_9212,N_8339);
xnor U11982 (N_11982,N_8890,N_8561);
nand U11983 (N_11983,N_8654,N_8212);
nor U11984 (N_11984,N_8469,N_8482);
and U11985 (N_11985,N_8745,N_9686);
nand U11986 (N_11986,N_8963,N_9007);
or U11987 (N_11987,N_9660,N_9598);
nor U11988 (N_11988,N_8524,N_8874);
nor U11989 (N_11989,N_8444,N_9542);
or U11990 (N_11990,N_8879,N_8291);
or U11991 (N_11991,N_9275,N_9125);
or U11992 (N_11992,N_9824,N_9688);
or U11993 (N_11993,N_8396,N_9843);
or U11994 (N_11994,N_9389,N_9580);
or U11995 (N_11995,N_8508,N_9146);
or U11996 (N_11996,N_9257,N_8706);
nor U11997 (N_11997,N_9457,N_8263);
nand U11998 (N_11998,N_9042,N_8570);
nor U11999 (N_11999,N_9236,N_9953);
nor U12000 (N_12000,N_10726,N_10631);
or U12001 (N_12001,N_11987,N_10196);
and U12002 (N_12002,N_11871,N_10009);
and U12003 (N_12003,N_10439,N_11506);
xor U12004 (N_12004,N_10594,N_11312);
and U12005 (N_12005,N_11501,N_11999);
and U12006 (N_12006,N_10056,N_11933);
or U12007 (N_12007,N_11235,N_11483);
xnor U12008 (N_12008,N_10936,N_10213);
nand U12009 (N_12009,N_10428,N_10808);
xnor U12010 (N_12010,N_11671,N_11746);
nor U12011 (N_12011,N_11587,N_11602);
nor U12012 (N_12012,N_11706,N_11583);
nand U12013 (N_12013,N_11254,N_11723);
nand U12014 (N_12014,N_11328,N_11337);
and U12015 (N_12015,N_10258,N_11864);
nand U12016 (N_12016,N_11000,N_10846);
nor U12017 (N_12017,N_11157,N_10335);
nand U12018 (N_12018,N_11414,N_10677);
xnor U12019 (N_12019,N_11816,N_10382);
or U12020 (N_12020,N_11975,N_11510);
and U12021 (N_12021,N_11817,N_11439);
nor U12022 (N_12022,N_11363,N_10577);
nand U12023 (N_12023,N_11520,N_10780);
nor U12024 (N_12024,N_11650,N_10195);
nor U12025 (N_12025,N_11278,N_10815);
xor U12026 (N_12026,N_10110,N_10272);
xnor U12027 (N_12027,N_11504,N_10167);
or U12028 (N_12028,N_11112,N_11799);
xnor U12029 (N_12029,N_10743,N_11589);
xnor U12030 (N_12030,N_11007,N_10522);
and U12031 (N_12031,N_11986,N_11804);
xor U12032 (N_12032,N_10850,N_10853);
nand U12033 (N_12033,N_10068,N_10061);
xor U12034 (N_12034,N_10896,N_10178);
or U12035 (N_12035,N_10361,N_10977);
xnor U12036 (N_12036,N_10429,N_10425);
or U12037 (N_12037,N_10779,N_11712);
xor U12038 (N_12038,N_10697,N_10922);
and U12039 (N_12039,N_11239,N_10705);
nand U12040 (N_12040,N_11862,N_11123);
xor U12041 (N_12041,N_10529,N_11751);
and U12042 (N_12042,N_11956,N_11702);
xnor U12043 (N_12043,N_11904,N_10290);
and U12044 (N_12044,N_10231,N_10042);
or U12045 (N_12045,N_11297,N_11279);
or U12046 (N_12046,N_10750,N_10444);
nand U12047 (N_12047,N_10207,N_11745);
nand U12048 (N_12048,N_10038,N_10398);
nor U12049 (N_12049,N_10812,N_10860);
xnor U12050 (N_12050,N_11866,N_11982);
nor U12051 (N_12051,N_11764,N_10700);
nand U12052 (N_12052,N_10232,N_10205);
xor U12053 (N_12053,N_10332,N_10895);
xor U12054 (N_12054,N_11051,N_10737);
or U12055 (N_12055,N_10498,N_11072);
and U12056 (N_12056,N_10451,N_11030);
nor U12057 (N_12057,N_10490,N_10802);
nand U12058 (N_12058,N_10010,N_10915);
nand U12059 (N_12059,N_11545,N_10740);
nor U12060 (N_12060,N_11559,N_10914);
and U12061 (N_12061,N_10655,N_11819);
nand U12062 (N_12062,N_10701,N_10172);
or U12063 (N_12063,N_11568,N_11089);
or U12064 (N_12064,N_11682,N_11640);
and U12065 (N_12065,N_11894,N_10098);
xor U12066 (N_12066,N_11515,N_10239);
nand U12067 (N_12067,N_10663,N_11042);
or U12068 (N_12068,N_11431,N_10659);
and U12069 (N_12069,N_10997,N_11073);
nor U12070 (N_12070,N_11884,N_10648);
and U12071 (N_12071,N_10596,N_11406);
or U12072 (N_12072,N_11162,N_10958);
xor U12073 (N_12073,N_11518,N_10461);
or U12074 (N_12074,N_10643,N_11181);
and U12075 (N_12075,N_10792,N_10400);
nor U12076 (N_12076,N_11202,N_10575);
nand U12077 (N_12077,N_11873,N_10970);
nand U12078 (N_12078,N_11018,N_11453);
nor U12079 (N_12079,N_11209,N_11293);
nand U12080 (N_12080,N_10557,N_11796);
or U12081 (N_12081,N_10587,N_11826);
nand U12082 (N_12082,N_11379,N_10026);
nand U12083 (N_12083,N_11789,N_11105);
xor U12084 (N_12084,N_10766,N_11582);
nand U12085 (N_12085,N_10025,N_11617);
and U12086 (N_12086,N_10560,N_10285);
xnor U12087 (N_12087,N_11497,N_11776);
and U12088 (N_12088,N_11377,N_10538);
xnor U12089 (N_12089,N_10670,N_10842);
and U12090 (N_12090,N_10475,N_11121);
nor U12091 (N_12091,N_10609,N_11075);
xnor U12092 (N_12092,N_10640,N_11410);
nor U12093 (N_12093,N_11253,N_10013);
nand U12094 (N_12094,N_11949,N_10411);
or U12095 (N_12095,N_11144,N_10122);
nor U12096 (N_12096,N_10987,N_11326);
or U12097 (N_12097,N_11918,N_11296);
nand U12098 (N_12098,N_11860,N_11141);
nand U12099 (N_12099,N_11781,N_11777);
or U12100 (N_12100,N_10313,N_10286);
nand U12101 (N_12101,N_10985,N_11644);
xnor U12102 (N_12102,N_10496,N_11450);
xnor U12103 (N_12103,N_10797,N_10480);
or U12104 (N_12104,N_10800,N_11138);
xnor U12105 (N_12105,N_11333,N_10765);
and U12106 (N_12106,N_11403,N_11736);
or U12107 (N_12107,N_10369,N_11445);
xor U12108 (N_12108,N_10913,N_11536);
xor U12109 (N_12109,N_11204,N_10569);
nor U12110 (N_12110,N_11772,N_10757);
nor U12111 (N_12111,N_10535,N_10464);
nor U12112 (N_12112,N_10789,N_11355);
xnor U12113 (N_12113,N_10069,N_11767);
or U12114 (N_12114,N_11897,N_11785);
or U12115 (N_12115,N_11045,N_10581);
nor U12116 (N_12116,N_10316,N_10455);
or U12117 (N_12117,N_10044,N_11649);
and U12118 (N_12118,N_10637,N_11662);
nor U12119 (N_12119,N_11538,N_11511);
and U12120 (N_12120,N_10248,N_11359);
or U12121 (N_12121,N_10152,N_11747);
and U12122 (N_12122,N_10889,N_10019);
xnor U12123 (N_12123,N_10409,N_11319);
or U12124 (N_12124,N_10988,N_10549);
or U12125 (N_12125,N_10857,N_10747);
or U12126 (N_12126,N_10270,N_10015);
and U12127 (N_12127,N_11820,N_10040);
xnor U12128 (N_12128,N_10518,N_11651);
and U12129 (N_12129,N_10228,N_11216);
nand U12130 (N_12130,N_10884,N_11464);
or U12131 (N_12131,N_10082,N_11783);
nor U12132 (N_12132,N_10991,N_10874);
or U12133 (N_12133,N_11093,N_11201);
or U12134 (N_12134,N_11806,N_11726);
nand U12135 (N_12135,N_10407,N_11482);
nor U12136 (N_12136,N_11957,N_11594);
xnor U12137 (N_12137,N_11125,N_11686);
and U12138 (N_12138,N_10442,N_10841);
or U12139 (N_12139,N_10224,N_10667);
or U12140 (N_12140,N_11461,N_10719);
nand U12141 (N_12141,N_11366,N_11596);
nor U12142 (N_12142,N_10163,N_10410);
and U12143 (N_12143,N_10683,N_11985);
or U12144 (N_12144,N_11234,N_10030);
nand U12145 (N_12145,N_10756,N_10331);
nand U12146 (N_12146,N_10337,N_11930);
or U12147 (N_12147,N_10097,N_11610);
and U12148 (N_12148,N_11291,N_10778);
and U12149 (N_12149,N_11586,N_11529);
xnor U12150 (N_12150,N_10347,N_11967);
and U12151 (N_12151,N_10665,N_11766);
or U12152 (N_12152,N_10927,N_10062);
nor U12153 (N_12153,N_10008,N_10482);
xnor U12154 (N_12154,N_11564,N_10657);
nand U12155 (N_12155,N_11437,N_10277);
nor U12156 (N_12156,N_10311,N_10000);
xnor U12157 (N_12157,N_11939,N_11146);
and U12158 (N_12158,N_10317,N_11019);
and U12159 (N_12159,N_11094,N_11169);
xor U12160 (N_12160,N_10767,N_11067);
xnor U12161 (N_12161,N_11350,N_11740);
nand U12162 (N_12162,N_10489,N_11922);
nand U12163 (N_12163,N_10553,N_10809);
and U12164 (N_12164,N_10295,N_11632);
nor U12165 (N_12165,N_11412,N_10945);
nand U12166 (N_12166,N_11033,N_10516);
xor U12167 (N_12167,N_10982,N_10505);
nor U12168 (N_12168,N_11593,N_11393);
nand U12169 (N_12169,N_10832,N_10269);
xnor U12170 (N_12170,N_10894,N_10605);
and U12171 (N_12171,N_10626,N_10865);
nand U12172 (N_12172,N_11352,N_11277);
nor U12173 (N_12173,N_10817,N_10979);
nor U12174 (N_12174,N_11635,N_10261);
nor U12175 (N_12175,N_11074,N_11679);
or U12176 (N_12176,N_11211,N_10103);
nand U12177 (N_12177,N_10628,N_10322);
or U12178 (N_12178,N_10969,N_10137);
or U12179 (N_12179,N_11775,N_10380);
nor U12180 (N_12180,N_11696,N_10194);
and U12181 (N_12181,N_11032,N_11264);
or U12182 (N_12182,N_11378,N_11976);
or U12183 (N_12183,N_11875,N_10078);
xnor U12184 (N_12184,N_11150,N_10129);
nor U12185 (N_12185,N_10217,N_11595);
or U12186 (N_12186,N_11334,N_11080);
nand U12187 (N_12187,N_11056,N_10084);
xnor U12188 (N_12188,N_11044,N_11699);
nand U12189 (N_12189,N_10028,N_11100);
xor U12190 (N_12190,N_10158,N_10859);
or U12191 (N_12191,N_10179,N_10054);
nand U12192 (N_12192,N_11579,N_10171);
nor U12193 (N_12193,N_11308,N_10121);
nand U12194 (N_12194,N_11707,N_10828);
nand U12195 (N_12195,N_10704,N_10996);
or U12196 (N_12196,N_10572,N_11238);
and U12197 (N_12197,N_10067,N_11843);
nor U12198 (N_12198,N_10707,N_11441);
or U12199 (N_12199,N_11742,N_11294);
xor U12200 (N_12200,N_11349,N_10983);
or U12201 (N_12201,N_11143,N_11332);
or U12202 (N_12202,N_10055,N_11286);
xnor U12203 (N_12203,N_11171,N_10512);
xor U12204 (N_12204,N_11274,N_10112);
or U12205 (N_12205,N_11857,N_10826);
nor U12206 (N_12206,N_10452,N_11365);
xnor U12207 (N_12207,N_11315,N_10764);
and U12208 (N_12208,N_10250,N_11313);
or U12209 (N_12209,N_11547,N_10672);
and U12210 (N_12210,N_10928,N_10556);
or U12211 (N_12211,N_10708,N_11495);
and U12212 (N_12212,N_10245,N_11174);
xnor U12213 (N_12213,N_11267,N_11229);
xor U12214 (N_12214,N_11544,N_10241);
nand U12215 (N_12215,N_11280,N_10159);
nor U12216 (N_12216,N_10187,N_10762);
or U12217 (N_12217,N_11401,N_10488);
nor U12218 (N_12218,N_11903,N_10905);
and U12219 (N_12219,N_11036,N_10681);
and U12220 (N_12220,N_11654,N_10036);
nor U12221 (N_12221,N_11320,N_11060);
xnor U12222 (N_12222,N_11118,N_10118);
and U12223 (N_12223,N_10106,N_10325);
and U12224 (N_12224,N_11295,N_10579);
xnor U12225 (N_12225,N_10304,N_11448);
nor U12226 (N_12226,N_11103,N_11489);
or U12227 (N_12227,N_11537,N_10023);
nand U12228 (N_12228,N_10554,N_10869);
xnor U12229 (N_12229,N_11344,N_11847);
nor U12230 (N_12230,N_10301,N_11387);
nor U12231 (N_12231,N_11020,N_11895);
xnor U12232 (N_12232,N_11752,N_11227);
nand U12233 (N_12233,N_11400,N_10260);
nor U12234 (N_12234,N_11762,N_11372);
xnor U12235 (N_12235,N_11805,N_10746);
nor U12236 (N_12236,N_11442,N_11630);
or U12237 (N_12237,N_10547,N_11941);
and U12238 (N_12238,N_10170,N_10733);
nand U12239 (N_12239,N_11914,N_10882);
nor U12240 (N_12240,N_11021,N_10117);
xnor U12241 (N_12241,N_11733,N_11323);
nor U12242 (N_12242,N_11912,N_10578);
or U12243 (N_12243,N_10471,N_10059);
nand U12244 (N_12244,N_11732,N_10555);
or U12245 (N_12245,N_11688,N_11833);
nand U12246 (N_12246,N_11505,N_11485);
nor U12247 (N_12247,N_10775,N_11135);
nand U12248 (N_12248,N_10240,N_11656);
xnor U12249 (N_12249,N_11932,N_11503);
nor U12250 (N_12250,N_11576,N_10323);
or U12251 (N_12251,N_11142,N_10660);
nor U12252 (N_12252,N_10266,N_10508);
nor U12253 (N_12253,N_11413,N_10495);
or U12254 (N_12254,N_11787,N_10289);
nand U12255 (N_12255,N_11164,N_11402);
or U12256 (N_12256,N_11797,N_11698);
or U12257 (N_12257,N_10956,N_10976);
xor U12258 (N_12258,N_10012,N_10709);
or U12259 (N_12259,N_11486,N_10145);
xor U12260 (N_12260,N_10847,N_10748);
xor U12261 (N_12261,N_11149,N_10345);
nand U12262 (N_12262,N_11172,N_11853);
and U12263 (N_12263,N_11512,N_10702);
and U12264 (N_12264,N_10005,N_11147);
nand U12265 (N_12265,N_10146,N_10920);
nor U12266 (N_12266,N_10220,N_11900);
or U12267 (N_12267,N_11447,N_10706);
and U12268 (N_12268,N_11024,N_11066);
nand U12269 (N_12269,N_10080,N_10811);
or U12270 (N_12270,N_10203,N_11327);
and U12271 (N_12271,N_10181,N_11906);
and U12272 (N_12272,N_10161,N_10511);
and U12273 (N_12273,N_11331,N_11119);
or U12274 (N_12274,N_11513,N_10014);
xor U12275 (N_12275,N_10230,N_10823);
xnor U12276 (N_12276,N_10052,N_11492);
nand U12277 (N_12277,N_11523,N_10673);
nand U12278 (N_12278,N_11658,N_10786);
nand U12279 (N_12279,N_11068,N_10132);
nor U12280 (N_12280,N_11339,N_10598);
xnor U12281 (N_12281,N_10046,N_10177);
or U12282 (N_12282,N_10543,N_10022);
nand U12283 (N_12283,N_10388,N_10507);
nor U12284 (N_12284,N_10074,N_10263);
or U12285 (N_12285,N_11354,N_11309);
nand U12286 (N_12286,N_11531,N_10453);
nand U12287 (N_12287,N_11759,N_11034);
xor U12288 (N_12288,N_11116,N_10405);
and U12289 (N_12289,N_11476,N_11233);
or U12290 (N_12290,N_10227,N_10933);
xnor U12291 (N_12291,N_10190,N_10592);
nor U12292 (N_12292,N_10477,N_11053);
and U12293 (N_12293,N_11770,N_11876);
or U12294 (N_12294,N_11472,N_10472);
and U12295 (N_12295,N_10342,N_11009);
and U12296 (N_12296,N_10136,N_10206);
and U12297 (N_12297,N_10492,N_11952);
or U12298 (N_12298,N_10049,N_11756);
xor U12299 (N_12299,N_11604,N_10680);
or U12300 (N_12300,N_10413,N_10381);
nand U12301 (N_12301,N_11769,N_11385);
xnor U12302 (N_12302,N_11728,N_11316);
or U12303 (N_12303,N_11257,N_11054);
and U12304 (N_12304,N_10794,N_11913);
and U12305 (N_12305,N_11383,N_10688);
nor U12306 (N_12306,N_10840,N_10037);
nand U12307 (N_12307,N_11660,N_11029);
or U12308 (N_12308,N_11388,N_10386);
xor U12309 (N_12309,N_11394,N_11236);
xnor U12310 (N_12310,N_11446,N_10645);
nor U12311 (N_12311,N_10478,N_11189);
nand U12312 (N_12312,N_11893,N_11697);
or U12313 (N_12313,N_10109,N_11182);
nor U12314 (N_12314,N_11028,N_10276);
and U12315 (N_12315,N_10283,N_11719);
xnor U12316 (N_12316,N_10018,N_10359);
and U12317 (N_12317,N_11006,N_11151);
nand U12318 (N_12318,N_11621,N_10613);
nor U12319 (N_12319,N_11376,N_11082);
and U12320 (N_12320,N_10917,N_10404);
nand U12321 (N_12321,N_10449,N_10868);
nor U12322 (N_12322,N_11969,N_11451);
nor U12323 (N_12323,N_11546,N_10566);
nor U12324 (N_12324,N_10684,N_11065);
or U12325 (N_12325,N_10935,N_10744);
xnor U12326 (N_12326,N_11578,N_10218);
nor U12327 (N_12327,N_10534,N_10952);
nand U12328 (N_12328,N_10938,N_11270);
or U12329 (N_12329,N_10338,N_11902);
nor U12330 (N_12330,N_10070,N_10873);
xor U12331 (N_12331,N_10953,N_10561);
xor U12332 (N_12332,N_10918,N_11916);
nand U12333 (N_12333,N_11481,N_10612);
nor U12334 (N_12334,N_11432,N_10047);
or U12335 (N_12335,N_10354,N_11812);
nand U12336 (N_12336,N_11101,N_11842);
xnor U12337 (N_12337,N_10924,N_10769);
and U12338 (N_12338,N_11543,N_11207);
xnor U12339 (N_12339,N_10259,N_11592);
or U12340 (N_12340,N_10622,N_10607);
nand U12341 (N_12341,N_11829,N_10777);
or U12342 (N_12342,N_10813,N_10830);
nor U12343 (N_12343,N_11725,N_11888);
nand U12344 (N_12344,N_10265,N_11892);
and U12345 (N_12345,N_11250,N_10154);
xor U12346 (N_12346,N_10793,N_10751);
or U12347 (N_12347,N_11200,N_10362);
nor U12348 (N_12348,N_11087,N_11477);
nand U12349 (N_12349,N_10827,N_10545);
xor U12350 (N_12350,N_11490,N_10950);
nand U12351 (N_12351,N_11920,N_10457);
xnor U12352 (N_12352,N_10002,N_11611);
nand U12353 (N_12353,N_11645,N_11273);
nor U12354 (N_12354,N_10053,N_11416);
and U12355 (N_12355,N_10866,N_10336);
xnor U12356 (N_12356,N_11824,N_11516);
nand U12357 (N_12357,N_10698,N_10906);
nand U12358 (N_12358,N_10685,N_11931);
and U12359 (N_12359,N_11836,N_10877);
and U12360 (N_12360,N_11247,N_10377);
and U12361 (N_12361,N_10458,N_11569);
or U12362 (N_12362,N_11591,N_11924);
xnor U12363 (N_12363,N_10091,N_10975);
nor U12364 (N_12364,N_10763,N_11553);
nand U12365 (N_12365,N_10741,N_11782);
nor U12366 (N_12366,N_11950,N_11026);
xnor U12367 (N_12367,N_10804,N_10689);
and U12368 (N_12368,N_11220,N_10774);
or U12369 (N_12369,N_11438,N_11452);
and U12370 (N_12370,N_10288,N_11960);
or U12371 (N_12371,N_10192,N_11744);
nor U12372 (N_12372,N_10200,N_11137);
nand U12373 (N_12373,N_10424,N_11471);
nor U12374 (N_12374,N_11071,N_10222);
nor U12375 (N_12375,N_11289,N_11565);
nand U12376 (N_12376,N_10450,N_10414);
nor U12377 (N_12377,N_11727,N_10324);
nor U12378 (N_12378,N_11830,N_11374);
xnor U12379 (N_12379,N_11768,N_11222);
nor U12380 (N_12380,N_11680,N_10155);
nand U12381 (N_12381,N_11132,N_11643);
nor U12382 (N_12382,N_10327,N_10406);
nor U12383 (N_12383,N_10372,N_11556);
and U12384 (N_12384,N_11117,N_11714);
nand U12385 (N_12385,N_10831,N_10422);
and U12386 (N_12386,N_10093,N_10050);
xnor U12387 (N_12387,N_10135,N_10807);
xor U12388 (N_12388,N_10166,N_10676);
xnor U12389 (N_12389,N_11700,N_11231);
and U12390 (N_12390,N_11599,N_11979);
and U12391 (N_12391,N_11195,N_10147);
xor U12392 (N_12392,N_10908,N_10293);
nor U12393 (N_12393,N_10716,N_10770);
nand U12394 (N_12394,N_10493,N_11272);
or U12395 (N_12395,N_10686,N_11667);
or U12396 (N_12396,N_11124,N_10870);
nor U12397 (N_12397,N_10368,N_10510);
nor U12398 (N_12398,N_10588,N_10041);
and U12399 (N_12399,N_11059,N_10108);
nor U12400 (N_12400,N_10140,N_11104);
xor U12401 (N_12401,N_10102,N_11574);
and U12402 (N_12402,N_10394,N_11618);
or U12403 (N_12403,N_10189,N_10524);
and U12404 (N_12404,N_10517,N_10034);
nand U12405 (N_12405,N_11223,N_11647);
or U12406 (N_12406,N_10848,N_10113);
nand U12407 (N_12407,N_10968,N_10732);
xnor U12408 (N_12408,N_11739,N_10459);
or U12409 (N_12409,N_11384,N_10635);
or U12410 (N_12410,N_10173,N_11981);
or U12411 (N_12411,N_10986,N_10086);
nand U12412 (N_12412,N_10902,N_11525);
xnor U12413 (N_12413,N_10421,N_11380);
xor U12414 (N_12414,N_10574,N_11735);
nand U12415 (N_12415,N_10785,N_11226);
or U12416 (N_12416,N_11984,N_10937);
xor U12417 (N_12417,N_10485,N_10799);
and U12418 (N_12418,N_10964,N_10654);
xnor U12419 (N_12419,N_10717,N_11259);
nor U12420 (N_12420,N_11214,N_11502);
xnor U12421 (N_12421,N_11798,N_11815);
xnor U12422 (N_12422,N_11346,N_10509);
or U12423 (N_12423,N_11269,N_11340);
or U12424 (N_12424,N_10237,N_11803);
or U12425 (N_12425,N_11887,N_10514);
nand U12426 (N_12426,N_10900,N_11710);
xnor U12427 (N_12427,N_10946,N_11668);
and U12428 (N_12428,N_11039,N_11153);
nor U12429 (N_12429,N_10352,N_11832);
or U12430 (N_12430,N_10749,N_10564);
xor U12431 (N_12431,N_10923,N_11616);
nand U12432 (N_12432,N_11549,N_11301);
nor U12433 (N_12433,N_11625,N_10142);
xnor U12434 (N_12434,N_10223,N_11780);
xor U12435 (N_12435,N_10298,N_11290);
nor U12436 (N_12436,N_11844,N_10710);
nand U12437 (N_12437,N_10065,N_11426);
or U12438 (N_12438,N_10585,N_10888);
nand U12439 (N_12439,N_11588,N_10085);
nor U12440 (N_12440,N_10818,N_10590);
nand U12441 (N_12441,N_10836,N_10638);
xnor U12442 (N_12442,N_10233,N_11534);
nor U12443 (N_12443,N_10878,N_10990);
nand U12444 (N_12444,N_10433,N_10552);
nor U12445 (N_12445,N_10835,N_10718);
or U12446 (N_12446,N_10910,N_11687);
and U12447 (N_12447,N_11191,N_11993);
nand U12448 (N_12448,N_11889,N_11178);
xnor U12449 (N_12449,N_11911,N_10519);
nor U12450 (N_12450,N_10466,N_11262);
or U12451 (N_12451,N_11694,N_11014);
nand U12452 (N_12452,N_10401,N_11934);
or U12453 (N_12453,N_11827,N_10760);
or U12454 (N_12454,N_11314,N_11825);
xnor U12455 (N_12455,N_10297,N_10119);
nand U12456 (N_12456,N_11851,N_11002);
or U12457 (N_12457,N_10963,N_11003);
nor U12458 (N_12458,N_11695,N_11245);
nor U12459 (N_12459,N_11869,N_11557);
or U12460 (N_12460,N_11653,N_10803);
or U12461 (N_12461,N_11937,N_11677);
nand U12462 (N_12462,N_11821,N_11057);
nor U12463 (N_12463,N_10175,N_11743);
xor U12464 (N_12464,N_10758,N_11282);
or U12465 (N_12465,N_11637,N_10476);
nand U12466 (N_12466,N_10530,N_11997);
xnor U12467 (N_12467,N_11584,N_11901);
xnor U12468 (N_12468,N_11040,N_10833);
nand U12469 (N_12469,N_11008,N_11753);
nand U12470 (N_12470,N_10378,N_11995);
xor U12471 (N_12471,N_10864,N_11642);
nand U12472 (N_12472,N_11013,N_10045);
nor U12473 (N_12473,N_10951,N_11715);
xnor U12474 (N_12474,N_10202,N_11165);
xnor U12475 (N_12475,N_10282,N_10788);
or U12476 (N_12476,N_10491,N_10576);
or U12477 (N_12477,N_11685,N_11167);
nand U12478 (N_12478,N_11455,N_11962);
xor U12479 (N_12479,N_11404,N_11943);
nand U12480 (N_12480,N_10736,N_10912);
or U12481 (N_12481,N_11088,N_11846);
or U12482 (N_12482,N_11307,N_11923);
and U12483 (N_12483,N_10973,N_11266);
xnor U12484 (N_12484,N_11411,N_10387);
nand U12485 (N_12485,N_11136,N_11938);
nor U12486 (N_12486,N_11133,N_11325);
xor U12487 (N_12487,N_11241,N_10739);
xnor U12488 (N_12488,N_10210,N_10426);
nand U12489 (N_12489,N_11757,N_11217);
or U12490 (N_12490,N_11140,N_11620);
nand U12491 (N_12491,N_11940,N_11083);
nand U12492 (N_12492,N_11417,N_10995);
xnor U12493 (N_12493,N_10043,N_11122);
nand U12494 (N_12494,N_11397,N_10370);
or U12495 (N_12495,N_11945,N_11703);
nand U12496 (N_12496,N_11213,N_11391);
xnor U12497 (N_12497,N_11590,N_10271);
xor U12498 (N_12498,N_10017,N_10076);
or U12499 (N_12499,N_11347,N_10253);
or U12500 (N_12500,N_11638,N_11128);
xnor U12501 (N_12501,N_10723,N_10584);
nor U12502 (N_12502,N_11530,N_10903);
xnor U12503 (N_12503,N_10416,N_10721);
xor U12504 (N_12504,N_11351,N_10989);
or U12505 (N_12505,N_11305,N_10219);
or U12506 (N_12506,N_10214,N_11225);
or U12507 (N_12507,N_10801,N_11935);
xor U12508 (N_12508,N_11158,N_10443);
xnor U12509 (N_12509,N_10427,N_10363);
nor U12510 (N_12510,N_10057,N_10226);
and U12511 (N_12511,N_10696,N_11463);
or U12512 (N_12512,N_11669,N_11598);
or U12513 (N_12513,N_11808,N_11023);
nand U12514 (N_12514,N_11362,N_11716);
and U12515 (N_12515,N_11251,N_10264);
xnor U12516 (N_12516,N_11246,N_10312);
nand U12517 (N_12517,N_10412,N_11929);
and U12518 (N_12518,N_11069,N_11988);
or U12519 (N_12519,N_10160,N_10174);
nor U12520 (N_12520,N_10502,N_10198);
xor U12521 (N_12521,N_10887,N_10360);
and U12522 (N_12522,N_11771,N_11629);
and U12523 (N_12523,N_11859,N_11341);
or U12524 (N_12524,N_11120,N_11398);
and U12525 (N_12525,N_10423,N_10334);
nand U12526 (N_12526,N_11881,N_10096);
xor U12527 (N_12527,N_11288,N_11657);
xnor U12528 (N_12528,N_11449,N_11130);
nor U12529 (N_12529,N_10504,N_11792);
or U12530 (N_12530,N_11183,N_11734);
nand U12531 (N_12531,N_11459,N_11898);
and U12532 (N_12532,N_10348,N_10081);
xor U12533 (N_12533,N_10911,N_10176);
xnor U12534 (N_12534,N_11196,N_11562);
nand U12535 (N_12535,N_10820,N_10366);
nor U12536 (N_12536,N_11188,N_11001);
nor U12537 (N_12537,N_11357,N_10357);
or U12538 (N_12538,N_11854,N_11237);
or U12539 (N_12539,N_11612,N_10284);
nor U12540 (N_12540,N_10941,N_10861);
and U12541 (N_12541,N_11551,N_11795);
nor U12542 (N_12542,N_10599,N_11509);
nand U12543 (N_12543,N_11615,N_10291);
and U12544 (N_12544,N_11641,N_10690);
nand U12545 (N_12545,N_11358,N_10186);
or U12546 (N_12546,N_11255,N_11905);
xnor U12547 (N_12547,N_10351,N_10650);
or U12548 (N_12548,N_11878,N_10460);
and U12549 (N_12549,N_11963,N_11050);
xnor U12550 (N_12550,N_11228,N_11025);
and U12551 (N_12551,N_10305,N_11915);
nand U12552 (N_12552,N_11457,N_11998);
xnor U12553 (N_12553,N_11692,N_11947);
and U12554 (N_12554,N_11194,N_11203);
nand U12555 (N_12555,N_10713,N_11891);
or U12556 (N_12556,N_10791,N_10185);
and U12557 (N_12557,N_10618,N_11396);
nor U12558 (N_12558,N_11978,N_11467);
and U12559 (N_12559,N_10441,N_11478);
and U12560 (N_12560,N_10408,N_10116);
nand U12561 (N_12561,N_10246,N_10940);
xnor U12562 (N_12562,N_10879,N_11925);
nand U12563 (N_12563,N_11711,N_11343);
or U12564 (N_12564,N_10183,N_10326);
nand U12565 (N_12565,N_10497,N_11936);
and U12566 (N_12566,N_11532,N_11198);
nor U12567 (N_12567,N_10101,N_11336);
xnor U12568 (N_12568,N_10075,N_10897);
or U12569 (N_12569,N_11555,N_11159);
or U12570 (N_12570,N_11199,N_10852);
xnor U12571 (N_12571,N_11306,N_11192);
nand U12572 (N_12572,N_11390,N_10314);
nor U12573 (N_12573,N_11542,N_11919);
xor U12574 (N_12574,N_11874,N_10615);
nand U12575 (N_12575,N_10204,N_11841);
or U12576 (N_12576,N_10463,N_11983);
nand U12577 (N_12577,N_10063,N_11990);
nand U12578 (N_12578,N_11422,N_10738);
and U12579 (N_12579,N_10420,N_11970);
nand U12580 (N_12580,N_11802,N_10402);
or U12581 (N_12581,N_10541,N_11521);
nand U12582 (N_12582,N_10930,N_10620);
or U12583 (N_12583,N_11047,N_11959);
xor U12584 (N_12584,N_10854,N_10356);
nor U12585 (N_12585,N_10715,N_11670);
or U12586 (N_12586,N_10006,N_11623);
nand U12587 (N_12587,N_11152,N_11335);
xor U12588 (N_12588,N_10845,N_10473);
nand U12589 (N_12589,N_11330,N_10446);
or U12590 (N_12590,N_11717,N_10099);
nand U12591 (N_12591,N_11527,N_11953);
nand U12592 (N_12592,N_11389,N_11041);
or U12593 (N_12593,N_11899,N_11129);
xor U12594 (N_12594,N_10862,N_11965);
and U12595 (N_12595,N_11908,N_10087);
xnor U12596 (N_12596,N_10971,N_10114);
nand U12597 (N_12597,N_11790,N_10647);
or U12598 (N_12598,N_10340,N_11705);
nor U12599 (N_12599,N_10071,N_11382);
and U12600 (N_12600,N_10838,N_11721);
xor U12601 (N_12601,N_11664,N_11016);
or U12602 (N_12602,N_10687,N_10771);
and U12603 (N_12603,N_10944,N_11224);
or U12604 (N_12604,N_11822,N_10652);
or U12605 (N_12605,N_11148,N_11737);
and U12606 (N_12606,N_11974,N_11600);
or U12607 (N_12607,N_10755,N_10661);
or U12608 (N_12608,N_10965,N_10153);
xnor U12609 (N_12609,N_11855,N_10383);
xnor U12610 (N_12610,N_11880,N_10024);
nor U12611 (N_12611,N_11896,N_11786);
nand U12612 (N_12612,N_11535,N_11801);
nor U12613 (N_12613,N_10948,N_10095);
and U12614 (N_12614,N_10191,N_10397);
nor U12615 (N_12615,N_10610,N_11111);
or U12616 (N_12616,N_10090,N_10583);
nand U12617 (N_12617,N_11865,N_11460);
nand U12618 (N_12618,N_10391,N_10532);
nor U12619 (N_12619,N_10287,N_10787);
nor U12620 (N_12620,N_10100,N_10904);
and U12621 (N_12621,N_10837,N_10515);
or U12622 (N_12622,N_11917,N_11749);
nor U12623 (N_12623,N_10967,N_11012);
xnor U12624 (N_12624,N_10379,N_11479);
xnor U12625 (N_12625,N_10440,N_10693);
xnor U12626 (N_12626,N_10367,N_10039);
nor U12627 (N_12627,N_11964,N_10959);
or U12628 (N_12628,N_11090,N_11672);
and U12629 (N_12629,N_10089,N_11318);
and U12630 (N_12630,N_11064,N_10481);
or U12631 (N_12631,N_11260,N_11704);
nor U12632 (N_12632,N_11176,N_11367);
or U12633 (N_12633,N_10188,N_10525);
nand U12634 (N_12634,N_11927,N_10724);
or U12635 (N_12635,N_11193,N_11818);
nand U12636 (N_12636,N_10201,N_10921);
and U12637 (N_12637,N_11170,N_10849);
xor U12638 (N_12638,N_10392,N_11469);
nand U12639 (N_12639,N_10582,N_11420);
nand U12640 (N_12640,N_10695,N_10734);
and U12641 (N_12641,N_11788,N_10972);
and U12642 (N_12642,N_10725,N_11581);
nand U12643 (N_12643,N_10768,N_10679);
and U12644 (N_12644,N_11256,N_10621);
nand U12645 (N_12645,N_10669,N_10344);
xor U12646 (N_12646,N_11639,N_11877);
and U12647 (N_12647,N_10759,N_10267);
nor U12648 (N_12648,N_10321,N_10784);
nor U12649 (N_12649,N_10567,N_11879);
and U12650 (N_12650,N_11971,N_10867);
xnor U12651 (N_12651,N_10292,N_10728);
xnor U12652 (N_12652,N_11070,N_10925);
nor U12653 (N_12653,N_11849,N_10550);
nor U12654 (N_12654,N_10916,N_11955);
xnor U12655 (N_12655,N_11648,N_10761);
xor U12656 (N_12656,N_11977,N_10373);
xnor U12657 (N_12657,N_11863,N_11741);
nor U12658 (N_12658,N_11989,N_11038);
and U12659 (N_12659,N_11415,N_10072);
or U12660 (N_12660,N_11175,N_11310);
nor U12661 (N_12661,N_10134,N_10124);
and U12662 (N_12662,N_11748,N_10961);
or U12663 (N_12663,N_10932,N_10694);
nand U12664 (N_12664,N_10559,N_11106);
nor U12665 (N_12665,N_10664,N_11996);
or U12666 (N_12666,N_11603,N_10551);
nand U12667 (N_12667,N_11261,N_11265);
and U12668 (N_12668,N_11561,N_10467);
nor U12669 (N_12669,N_10262,N_11046);
xnor U12670 (N_12670,N_11252,N_11760);
or U12671 (N_12671,N_10671,N_10130);
and U12672 (N_12672,N_11381,N_11329);
or U12673 (N_12673,N_10563,N_10625);
nor U12674 (N_12674,N_11673,N_11548);
nand U12675 (N_12675,N_11373,N_10462);
or U12676 (N_12676,N_10353,N_11454);
nor U12677 (N_12677,N_10573,N_10528);
or U12678 (N_12678,N_11284,N_11552);
nand U12679 (N_12679,N_11765,N_10494);
nor U12680 (N_12680,N_10315,N_10539);
nand U12681 (N_12681,N_10329,N_10162);
and U12682 (N_12682,N_10235,N_10814);
or U12683 (N_12683,N_10795,N_10893);
or U12684 (N_12684,N_10001,N_11814);
xor U12685 (N_12685,N_10568,N_10376);
xnor U12686 (N_12686,N_10330,N_10675);
xor U12687 (N_12687,N_10855,N_11550);
xor U12688 (N_12688,N_11809,N_11838);
nor U12689 (N_12689,N_11807,N_11300);
and U12690 (N_12690,N_11800,N_10431);
or U12691 (N_12691,N_10714,N_11356);
or U12692 (N_12692,N_11440,N_10127);
or U12693 (N_12693,N_10520,N_10623);
nor U12694 (N_12694,N_11585,N_10144);
xor U12695 (N_12695,N_11709,N_10506);
and U12696 (N_12696,N_10180,N_10674);
nand U12697 (N_12697,N_11205,N_11473);
nor U12698 (N_12698,N_10033,N_10521);
xnor U12699 (N_12699,N_11168,N_10339);
xnor U12700 (N_12700,N_11951,N_10021);
nor U12701 (N_12701,N_11249,N_11361);
nor U12702 (N_12702,N_10993,N_10875);
xor U12703 (N_12703,N_10562,N_11627);
and U12704 (N_12704,N_11468,N_10542);
or U12705 (N_12705,N_11156,N_10608);
or U12706 (N_12706,N_10602,N_10960);
or U12707 (N_12707,N_11661,N_10088);
nor U12708 (N_12708,N_10133,N_11944);
nand U12709 (N_12709,N_11628,N_11622);
or U12710 (N_12710,N_10051,N_11980);
xor U12711 (N_12711,N_10302,N_10216);
nand U12712 (N_12712,N_10310,N_10624);
nand U12713 (N_12713,N_10796,N_10333);
and U12714 (N_12714,N_10111,N_10934);
xor U12715 (N_12715,N_11519,N_11353);
nor U12716 (N_12716,N_10468,N_11921);
nand U12717 (N_12717,N_11499,N_11210);
xnor U12718 (N_12718,N_10527,N_11858);
nand U12719 (N_12719,N_11856,N_10469);
nand U12720 (N_12720,N_11948,N_10242);
and U12721 (N_12721,N_10128,N_10540);
or U12722 (N_12722,N_11185,N_10143);
and U12723 (N_12723,N_10595,N_10126);
xor U12724 (N_12724,N_10066,N_11834);
nand U12725 (N_12725,N_11077,N_11861);
nand U12726 (N_12726,N_11689,N_11099);
xor U12727 (N_12727,N_11973,N_11368);
nor U12728 (N_12728,N_10123,N_11160);
and U12729 (N_12729,N_11010,N_11244);
nand U12730 (N_12730,N_10994,N_10668);
nand U12731 (N_12731,N_10891,N_10341);
xnor U12732 (N_12732,N_10772,N_10212);
and U12733 (N_12733,N_11738,N_11281);
or U12734 (N_12734,N_10629,N_10589);
nand U12735 (N_12735,N_10844,N_10678);
xor U12736 (N_12736,N_10448,N_11731);
nand U12737 (N_12737,N_10531,N_11419);
or U12738 (N_12738,N_10798,N_10003);
nor U12739 (N_12739,N_10805,N_11232);
xnor U12740 (N_12740,N_10978,N_10225);
nand U12741 (N_12741,N_10454,N_11145);
nand U12742 (N_12742,N_11161,N_10658);
nand U12743 (N_12743,N_10546,N_11095);
nand U12744 (N_12744,N_10364,N_11774);
nor U12745 (N_12745,N_11540,N_10931);
xor U12746 (N_12746,N_10148,N_10954);
nand U12747 (N_12747,N_11794,N_10007);
or U12748 (N_12748,N_10107,N_11166);
nor U12749 (N_12749,N_10255,N_10955);
nor U12750 (N_12750,N_10822,N_10419);
xnor U12751 (N_12751,N_10371,N_10909);
or U12752 (N_12752,N_11248,N_10399);
and U12753 (N_12753,N_10943,N_10606);
xnor U12754 (N_12754,N_10503,N_11342);
nor U12755 (N_12755,N_10880,N_11126);
xnor U12756 (N_12756,N_11215,N_11408);
nor U12757 (N_12757,N_11605,N_11304);
nand U12758 (N_12758,N_11601,N_10415);
and U12759 (N_12759,N_11197,N_11691);
nand U12760 (N_12760,N_10790,N_10565);
xnor U12761 (N_12761,N_11392,N_10465);
and U12762 (N_12762,N_10632,N_11480);
or U12763 (N_12763,N_10249,N_10011);
and U12764 (N_12764,N_10389,N_11275);
xnor U12765 (N_12765,N_10244,N_11423);
and U12766 (N_12766,N_10892,N_10487);
nor U12767 (N_12767,N_10974,N_10484);
and U12768 (N_12768,N_10499,N_11498);
nor U12769 (N_12769,N_11494,N_10278);
nand U12770 (N_12770,N_11405,N_10843);
xnor U12771 (N_12771,N_10435,N_10169);
nand U12772 (N_12772,N_10729,N_11675);
or U12773 (N_12773,N_10571,N_11035);
or U12774 (N_12774,N_10004,N_10300);
nand U12775 (N_12775,N_10526,N_11263);
nand U12776 (N_12776,N_11434,N_10328);
nand U12777 (N_12777,N_10604,N_11429);
xor U12778 (N_12778,N_11163,N_11631);
and U12779 (N_12779,N_10825,N_10193);
nor U12780 (N_12780,N_11613,N_10156);
and U12781 (N_12781,N_10699,N_11507);
or U12782 (N_12782,N_11575,N_11154);
and U12783 (N_12783,N_11242,N_10883);
or U12784 (N_12784,N_11187,N_10149);
xnor U12785 (N_12785,N_11681,N_10251);
xnor U12786 (N_12786,N_10600,N_11085);
xor U12787 (N_12787,N_11835,N_10395);
nand U12788 (N_12788,N_11043,N_10720);
or U12789 (N_12789,N_11676,N_10580);
or U12790 (N_12790,N_10558,N_10586);
nor U12791 (N_12791,N_11155,N_10619);
or U12792 (N_12792,N_10168,N_10350);
and U12793 (N_12793,N_11666,N_11190);
nor U12794 (N_12794,N_11465,N_10703);
and U12795 (N_12795,N_10275,N_11011);
nor U12796 (N_12796,N_10656,N_10773);
nor U12797 (N_12797,N_11539,N_10630);
nor U12798 (N_12798,N_10999,N_11646);
nor U12799 (N_12799,N_10810,N_10470);
nand U12800 (N_12800,N_10474,N_11427);
and U12801 (N_12801,N_10273,N_11399);
nor U12802 (N_12802,N_10616,N_11219);
xor U12803 (N_12803,N_11127,N_10027);
xor U12804 (N_12804,N_11597,N_11614);
xor U12805 (N_12805,N_11338,N_11386);
nand U12806 (N_12806,N_10486,N_10984);
and U12807 (N_12807,N_11991,N_10209);
or U12808 (N_12808,N_10603,N_11496);
and U12809 (N_12809,N_10886,N_10479);
nand U12810 (N_12810,N_11724,N_10032);
nand U12811 (N_12811,N_11514,N_11867);
xnor U12812 (N_12812,N_10863,N_10064);
and U12813 (N_12813,N_10048,N_11180);
and U12814 (N_12814,N_11364,N_10384);
nor U12815 (N_12815,N_11607,N_10644);
and U12816 (N_12816,N_11567,N_11558);
nand U12817 (N_12817,N_11317,N_11755);
xnor U12818 (N_12818,N_11287,N_11369);
xnor U12819 (N_12819,N_11580,N_11533);
and U12820 (N_12820,N_11395,N_11475);
or U12821 (N_12821,N_11212,N_11324);
nand U12822 (N_12822,N_10642,N_11092);
nand U12823 (N_12823,N_11528,N_11221);
nand U12824 (N_12824,N_11890,N_10731);
nand U12825 (N_12825,N_11872,N_10150);
nand U12826 (N_12826,N_10634,N_10268);
xor U12827 (N_12827,N_10501,N_10651);
or U12828 (N_12828,N_10839,N_11131);
nand U12829 (N_12829,N_10141,N_10318);
nand U12830 (N_12830,N_10980,N_10020);
nor U12831 (N_12831,N_10856,N_10742);
xor U12832 (N_12832,N_10164,N_11321);
nor U12833 (N_12833,N_11793,N_11754);
nand U12834 (N_12834,N_11823,N_10299);
nor U12835 (N_12835,N_11954,N_11828);
nor U12836 (N_12836,N_11779,N_10138);
nand U12837 (N_12837,N_10735,N_10730);
or U12838 (N_12838,N_11831,N_11665);
and U12839 (N_12839,N_10430,N_11690);
nand U12840 (N_12840,N_10094,N_10711);
xnor U12841 (N_12841,N_11466,N_11678);
or U12842 (N_12842,N_11571,N_11017);
xnor U12843 (N_12843,N_10029,N_11609);
nor U12844 (N_12844,N_10346,N_11102);
or U12845 (N_12845,N_11554,N_11443);
nand U12846 (N_12846,N_11348,N_10593);
nor U12847 (N_12847,N_10753,N_11701);
nor U12848 (N_12848,N_10806,N_11619);
or U12849 (N_12849,N_11958,N_11061);
or U12850 (N_12850,N_11302,N_10816);
xnor U12851 (N_12851,N_10396,N_11684);
nand U12852 (N_12852,N_10682,N_10434);
and U12853 (N_12853,N_11840,N_11285);
and U12854 (N_12854,N_11560,N_11436);
and U12855 (N_12855,N_11375,N_11062);
nor U12856 (N_12856,N_10403,N_10998);
nand U12857 (N_12857,N_11186,N_10834);
xor U12858 (N_12858,N_11430,N_11139);
or U12859 (N_12859,N_10436,N_11109);
nand U12860 (N_12860,N_10929,N_10890);
xnor U12861 (N_12861,N_10851,N_10208);
or U12862 (N_12862,N_11076,N_11462);
xnor U12863 (N_12863,N_11663,N_11885);
nor U12864 (N_12864,N_11522,N_11882);
nor U12865 (N_12865,N_10858,N_10781);
and U12866 (N_12866,N_11474,N_10390);
nand U12867 (N_12867,N_10919,N_11813);
nand U12868 (N_12868,N_11720,N_10418);
nor U12869 (N_12869,N_11811,N_10876);
or U12870 (N_12870,N_11444,N_10881);
xor U12871 (N_12871,N_11243,N_10907);
nor U12872 (N_12872,N_10365,N_10274);
nand U12873 (N_12873,N_10754,N_10303);
and U12874 (N_12874,N_10752,N_10992);
and U12875 (N_12875,N_11433,N_11946);
and U12876 (N_12876,N_11837,N_10627);
nand U12877 (N_12877,N_10949,N_10872);
and U12878 (N_12878,N_10374,N_11458);
nor U12879 (N_12879,N_10727,N_11791);
nand U12880 (N_12880,N_10438,N_10898);
xnor U12881 (N_12881,N_10597,N_10281);
nor U12882 (N_12882,N_11208,N_11299);
and U12883 (N_12883,N_10236,N_11470);
or U12884 (N_12884,N_11425,N_10035);
and U12885 (N_12885,N_10355,N_11992);
and U12886 (N_12886,N_10611,N_10139);
nand U12887 (N_12887,N_10280,N_10199);
nor U12888 (N_12888,N_11079,N_10483);
and U12889 (N_12889,N_10662,N_11435);
or U12890 (N_12890,N_11566,N_11230);
nor U12891 (N_12891,N_11910,N_10016);
nand U12892 (N_12892,N_11345,N_11418);
and U12893 (N_12893,N_11636,N_10885);
nand U12894 (N_12894,N_10456,N_10309);
or U12895 (N_12895,N_10060,N_10646);
nand U12896 (N_12896,N_10077,N_11500);
and U12897 (N_12897,N_11852,N_11966);
or U12898 (N_12898,N_11022,N_10417);
nand U12899 (N_12899,N_11276,N_10614);
and U12900 (N_12900,N_11303,N_11493);
xor U12901 (N_12901,N_10358,N_10824);
nor U12902 (N_12902,N_10537,N_10819);
or U12903 (N_12903,N_11078,N_11541);
nand U12904 (N_12904,N_11524,N_10296);
and U12905 (N_12905,N_11773,N_11968);
nand U12906 (N_12906,N_11110,N_11730);
or U12907 (N_12907,N_11371,N_10432);
or U12908 (N_12908,N_11722,N_10247);
nor U12909 (N_12909,N_10513,N_10073);
and U12910 (N_12910,N_11693,N_10197);
and U12911 (N_12911,N_10393,N_10092);
or U12912 (N_12912,N_10165,N_10385);
xor U12913 (N_12913,N_11298,N_11761);
or U12914 (N_12914,N_11049,N_11037);
xnor U12915 (N_12915,N_10079,N_11570);
nand U12916 (N_12916,N_10229,N_11926);
nand U12917 (N_12917,N_10131,N_11240);
nor U12918 (N_12918,N_11407,N_11108);
or U12919 (N_12919,N_10157,N_11907);
xnor U12920 (N_12920,N_11683,N_10899);
and U12921 (N_12921,N_11114,N_11218);
xor U12922 (N_12922,N_11508,N_10031);
nand U12923 (N_12923,N_11961,N_11886);
nand U12924 (N_12924,N_10692,N_11086);
nand U12925 (N_12925,N_10782,N_10544);
and U12926 (N_12926,N_11928,N_10105);
xor U12927 (N_12927,N_11179,N_11370);
or U12928 (N_12928,N_11942,N_11173);
nor U12929 (N_12929,N_10722,N_11004);
nor U12930 (N_12930,N_10234,N_11052);
nand U12931 (N_12931,N_11883,N_10548);
and U12932 (N_12932,N_10829,N_11870);
or U12933 (N_12933,N_11098,N_11268);
xnor U12934 (N_12934,N_10120,N_10447);
nor U12935 (N_12935,N_11311,N_10343);
and U12936 (N_12936,N_11091,N_11634);
nor U12937 (N_12937,N_11484,N_11031);
and U12938 (N_12938,N_11633,N_11563);
or U12939 (N_12939,N_10939,N_11517);
xnor U12940 (N_12940,N_10349,N_11360);
or U12941 (N_12941,N_11909,N_10437);
nand U12942 (N_12942,N_10256,N_10294);
nor U12943 (N_12943,N_10279,N_10666);
xnor U12944 (N_12944,N_11994,N_10871);
nor U12945 (N_12945,N_10901,N_11107);
or U12946 (N_12946,N_10617,N_11729);
nand U12947 (N_12947,N_10058,N_10243);
or U12948 (N_12948,N_10570,N_11713);
nor U12949 (N_12949,N_11322,N_11258);
or U12950 (N_12950,N_10712,N_10307);
nand U12951 (N_12951,N_11134,N_11015);
xnor U12952 (N_12952,N_11573,N_11058);
or U12953 (N_12953,N_11177,N_11624);
or U12954 (N_12954,N_11097,N_10783);
nand U12955 (N_12955,N_11084,N_11839);
and U12956 (N_12956,N_11850,N_11708);
xor U12957 (N_12957,N_11081,N_10215);
and U12958 (N_12958,N_10776,N_11784);
nand U12959 (N_12959,N_10966,N_10252);
nor U12960 (N_12960,N_10115,N_11491);
nand U12961 (N_12961,N_10633,N_11868);
or U12962 (N_12962,N_11428,N_10221);
or U12963 (N_12963,N_10254,N_10184);
and U12964 (N_12964,N_11271,N_11424);
xnor U12965 (N_12965,N_11778,N_10308);
nor U12966 (N_12966,N_10238,N_10151);
nor U12967 (N_12967,N_11763,N_11655);
nor U12968 (N_12968,N_10306,N_10649);
xor U12969 (N_12969,N_11027,N_11409);
nand U12970 (N_12970,N_11096,N_10523);
nor U12971 (N_12971,N_11487,N_11572);
and U12972 (N_12972,N_10942,N_10636);
or U12973 (N_12973,N_10926,N_11113);
nor U12974 (N_12974,N_11577,N_10319);
or U12975 (N_12975,N_11292,N_10104);
nand U12976 (N_12976,N_11115,N_10962);
and U12977 (N_12977,N_11421,N_11810);
nand U12978 (N_12978,N_11626,N_10981);
nand U12979 (N_12979,N_11456,N_11283);
or U12980 (N_12980,N_10533,N_11206);
or U12981 (N_12981,N_10639,N_11055);
xor U12982 (N_12982,N_11184,N_10445);
nand U12983 (N_12983,N_11848,N_11750);
xor U12984 (N_12984,N_11674,N_10375);
xnor U12985 (N_12985,N_10653,N_11608);
nand U12986 (N_12986,N_10745,N_10591);
xnor U12987 (N_12987,N_10957,N_11063);
xnor U12988 (N_12988,N_11048,N_11659);
nand U12989 (N_12989,N_10821,N_10083);
or U12990 (N_12990,N_10947,N_10257);
xor U12991 (N_12991,N_10211,N_10182);
or U12992 (N_12992,N_10691,N_11758);
or U12993 (N_12993,N_10641,N_11488);
or U12994 (N_12994,N_10601,N_11972);
and U12995 (N_12995,N_10320,N_11652);
nor U12996 (N_12996,N_11718,N_11526);
nor U12997 (N_12997,N_10125,N_10536);
nand U12998 (N_12998,N_11845,N_11606);
xor U12999 (N_12999,N_11005,N_10500);
xor U13000 (N_13000,N_10002,N_11227);
nand U13001 (N_13001,N_10916,N_10013);
xnor U13002 (N_13002,N_10807,N_11680);
or U13003 (N_13003,N_11765,N_11368);
nor U13004 (N_13004,N_10922,N_10594);
or U13005 (N_13005,N_10355,N_10026);
and U13006 (N_13006,N_11931,N_11174);
and U13007 (N_13007,N_10833,N_11086);
and U13008 (N_13008,N_11552,N_11008);
and U13009 (N_13009,N_11496,N_10763);
nand U13010 (N_13010,N_11028,N_10008);
and U13011 (N_13011,N_11701,N_11115);
and U13012 (N_13012,N_11396,N_11407);
nand U13013 (N_13013,N_10891,N_11831);
and U13014 (N_13014,N_11537,N_10614);
or U13015 (N_13015,N_10249,N_10635);
xor U13016 (N_13016,N_11808,N_11095);
or U13017 (N_13017,N_10813,N_10975);
and U13018 (N_13018,N_10030,N_10997);
nand U13019 (N_13019,N_11222,N_11923);
nor U13020 (N_13020,N_11031,N_11506);
nand U13021 (N_13021,N_11322,N_11306);
nor U13022 (N_13022,N_11611,N_11863);
or U13023 (N_13023,N_10575,N_10053);
nor U13024 (N_13024,N_10471,N_11345);
xnor U13025 (N_13025,N_11721,N_11614);
and U13026 (N_13026,N_10449,N_11313);
xor U13027 (N_13027,N_11522,N_10190);
nor U13028 (N_13028,N_10811,N_10212);
xor U13029 (N_13029,N_11281,N_11439);
nand U13030 (N_13030,N_10037,N_10201);
xor U13031 (N_13031,N_11358,N_11398);
xor U13032 (N_13032,N_11603,N_10790);
nor U13033 (N_13033,N_10256,N_10715);
and U13034 (N_13034,N_10324,N_11028);
and U13035 (N_13035,N_11326,N_10517);
nor U13036 (N_13036,N_10346,N_11816);
and U13037 (N_13037,N_11351,N_10485);
nor U13038 (N_13038,N_11899,N_10245);
nand U13039 (N_13039,N_11049,N_11406);
xor U13040 (N_13040,N_11799,N_11712);
nand U13041 (N_13041,N_10375,N_10581);
or U13042 (N_13042,N_11396,N_11793);
nor U13043 (N_13043,N_11499,N_11087);
xnor U13044 (N_13044,N_11259,N_10579);
nand U13045 (N_13045,N_11497,N_10383);
nand U13046 (N_13046,N_11431,N_10712);
and U13047 (N_13047,N_11257,N_11445);
and U13048 (N_13048,N_11239,N_11561);
nand U13049 (N_13049,N_11284,N_11146);
nor U13050 (N_13050,N_10535,N_10252);
or U13051 (N_13051,N_11178,N_11490);
nor U13052 (N_13052,N_10046,N_11955);
or U13053 (N_13053,N_11914,N_11797);
and U13054 (N_13054,N_11366,N_11455);
or U13055 (N_13055,N_11742,N_11489);
nor U13056 (N_13056,N_11788,N_10030);
or U13057 (N_13057,N_11160,N_11347);
xnor U13058 (N_13058,N_11901,N_11947);
and U13059 (N_13059,N_11761,N_11252);
nor U13060 (N_13060,N_10812,N_11186);
nand U13061 (N_13061,N_10995,N_11962);
xnor U13062 (N_13062,N_10659,N_11025);
nand U13063 (N_13063,N_10985,N_10848);
and U13064 (N_13064,N_11894,N_10336);
nand U13065 (N_13065,N_11014,N_11359);
xnor U13066 (N_13066,N_11725,N_10787);
nand U13067 (N_13067,N_11624,N_11022);
nand U13068 (N_13068,N_10154,N_10349);
or U13069 (N_13069,N_11638,N_11192);
nor U13070 (N_13070,N_11974,N_10888);
nor U13071 (N_13071,N_10518,N_11760);
and U13072 (N_13072,N_10283,N_11304);
nor U13073 (N_13073,N_11973,N_11858);
nand U13074 (N_13074,N_10620,N_11395);
or U13075 (N_13075,N_10162,N_10297);
nor U13076 (N_13076,N_10485,N_11215);
nand U13077 (N_13077,N_11766,N_11457);
xnor U13078 (N_13078,N_11536,N_10507);
xor U13079 (N_13079,N_11168,N_11321);
nand U13080 (N_13080,N_11233,N_11172);
or U13081 (N_13081,N_11043,N_11197);
xor U13082 (N_13082,N_11293,N_11623);
nand U13083 (N_13083,N_11731,N_10818);
nor U13084 (N_13084,N_11417,N_11753);
and U13085 (N_13085,N_11126,N_10705);
nand U13086 (N_13086,N_11305,N_10748);
nand U13087 (N_13087,N_10017,N_10205);
xnor U13088 (N_13088,N_10220,N_11921);
nor U13089 (N_13089,N_10394,N_11722);
nor U13090 (N_13090,N_10644,N_11896);
xor U13091 (N_13091,N_11797,N_10378);
or U13092 (N_13092,N_10366,N_11470);
xor U13093 (N_13093,N_11374,N_10442);
and U13094 (N_13094,N_10329,N_10279);
nand U13095 (N_13095,N_10389,N_10793);
nor U13096 (N_13096,N_10243,N_11775);
and U13097 (N_13097,N_10219,N_11752);
xnor U13098 (N_13098,N_11377,N_11854);
xnor U13099 (N_13099,N_11368,N_11873);
or U13100 (N_13100,N_10312,N_10977);
and U13101 (N_13101,N_10166,N_10765);
xnor U13102 (N_13102,N_11711,N_11463);
and U13103 (N_13103,N_11920,N_11295);
nor U13104 (N_13104,N_11052,N_11102);
and U13105 (N_13105,N_10515,N_10766);
and U13106 (N_13106,N_10935,N_10234);
xnor U13107 (N_13107,N_11775,N_10086);
and U13108 (N_13108,N_10427,N_10518);
and U13109 (N_13109,N_11202,N_10099);
and U13110 (N_13110,N_10670,N_11742);
and U13111 (N_13111,N_10370,N_11370);
or U13112 (N_13112,N_11475,N_11520);
or U13113 (N_13113,N_11795,N_10127);
or U13114 (N_13114,N_10959,N_11070);
nor U13115 (N_13115,N_10143,N_10225);
nand U13116 (N_13116,N_10004,N_11836);
or U13117 (N_13117,N_10984,N_11212);
nand U13118 (N_13118,N_10575,N_11741);
nand U13119 (N_13119,N_11987,N_10292);
or U13120 (N_13120,N_10165,N_11155);
nand U13121 (N_13121,N_10398,N_11864);
and U13122 (N_13122,N_10556,N_10766);
nand U13123 (N_13123,N_11764,N_11655);
or U13124 (N_13124,N_10651,N_10569);
nand U13125 (N_13125,N_10634,N_10109);
nand U13126 (N_13126,N_10053,N_11672);
or U13127 (N_13127,N_11687,N_11639);
and U13128 (N_13128,N_11297,N_11839);
and U13129 (N_13129,N_11967,N_11488);
or U13130 (N_13130,N_11096,N_10530);
xor U13131 (N_13131,N_10357,N_10397);
nor U13132 (N_13132,N_11943,N_11258);
or U13133 (N_13133,N_10273,N_11388);
xor U13134 (N_13134,N_11994,N_10064);
or U13135 (N_13135,N_11796,N_10954);
nand U13136 (N_13136,N_10530,N_10811);
xnor U13137 (N_13137,N_10642,N_10363);
and U13138 (N_13138,N_10494,N_11119);
and U13139 (N_13139,N_11352,N_11628);
nor U13140 (N_13140,N_11480,N_11870);
and U13141 (N_13141,N_10001,N_11798);
and U13142 (N_13142,N_11468,N_11338);
nor U13143 (N_13143,N_11902,N_10922);
xnor U13144 (N_13144,N_10956,N_11191);
nor U13145 (N_13145,N_11909,N_10463);
nand U13146 (N_13146,N_11913,N_10507);
and U13147 (N_13147,N_11594,N_10247);
nor U13148 (N_13148,N_11665,N_11599);
or U13149 (N_13149,N_11972,N_10557);
and U13150 (N_13150,N_11214,N_10661);
or U13151 (N_13151,N_11027,N_11587);
and U13152 (N_13152,N_10917,N_10533);
and U13153 (N_13153,N_11602,N_11759);
or U13154 (N_13154,N_10274,N_11862);
xor U13155 (N_13155,N_11811,N_11788);
and U13156 (N_13156,N_10753,N_11850);
nand U13157 (N_13157,N_11237,N_10174);
and U13158 (N_13158,N_10926,N_10762);
or U13159 (N_13159,N_10061,N_11120);
or U13160 (N_13160,N_11458,N_11422);
nor U13161 (N_13161,N_11128,N_11849);
nor U13162 (N_13162,N_11667,N_11105);
and U13163 (N_13163,N_10164,N_11742);
nand U13164 (N_13164,N_10251,N_11074);
nand U13165 (N_13165,N_11152,N_11457);
nor U13166 (N_13166,N_11919,N_10624);
nor U13167 (N_13167,N_10706,N_10876);
and U13168 (N_13168,N_11822,N_11943);
nand U13169 (N_13169,N_11959,N_11614);
and U13170 (N_13170,N_10729,N_10626);
and U13171 (N_13171,N_10570,N_11733);
or U13172 (N_13172,N_10227,N_11700);
nand U13173 (N_13173,N_11220,N_11789);
or U13174 (N_13174,N_11945,N_10008);
and U13175 (N_13175,N_11595,N_10195);
or U13176 (N_13176,N_11999,N_11272);
nand U13177 (N_13177,N_10927,N_11733);
nor U13178 (N_13178,N_11661,N_11020);
and U13179 (N_13179,N_10364,N_11095);
nand U13180 (N_13180,N_11578,N_10026);
nor U13181 (N_13181,N_10912,N_11621);
and U13182 (N_13182,N_11572,N_11319);
nand U13183 (N_13183,N_10577,N_11657);
and U13184 (N_13184,N_10529,N_11960);
and U13185 (N_13185,N_10810,N_10953);
xnor U13186 (N_13186,N_10118,N_10132);
nand U13187 (N_13187,N_11089,N_11711);
nor U13188 (N_13188,N_10134,N_11922);
or U13189 (N_13189,N_11501,N_10000);
xnor U13190 (N_13190,N_10065,N_11986);
nor U13191 (N_13191,N_10356,N_10949);
nand U13192 (N_13192,N_10382,N_11645);
or U13193 (N_13193,N_10362,N_10109);
xnor U13194 (N_13194,N_11510,N_10069);
nand U13195 (N_13195,N_11003,N_10324);
nand U13196 (N_13196,N_10665,N_11276);
and U13197 (N_13197,N_11446,N_11492);
or U13198 (N_13198,N_11310,N_11762);
xnor U13199 (N_13199,N_10464,N_11979);
nor U13200 (N_13200,N_11090,N_10719);
nand U13201 (N_13201,N_11911,N_11280);
and U13202 (N_13202,N_11285,N_10388);
and U13203 (N_13203,N_10875,N_10834);
nand U13204 (N_13204,N_11866,N_10980);
nand U13205 (N_13205,N_11028,N_11801);
nor U13206 (N_13206,N_11867,N_10876);
nor U13207 (N_13207,N_10464,N_10713);
xor U13208 (N_13208,N_10425,N_10986);
and U13209 (N_13209,N_11927,N_10610);
and U13210 (N_13210,N_11495,N_10406);
or U13211 (N_13211,N_10566,N_10030);
nand U13212 (N_13212,N_11255,N_11613);
nand U13213 (N_13213,N_11331,N_10849);
nor U13214 (N_13214,N_10291,N_10451);
nand U13215 (N_13215,N_11230,N_10028);
nor U13216 (N_13216,N_10658,N_11421);
xnor U13217 (N_13217,N_10108,N_10823);
nor U13218 (N_13218,N_11676,N_11866);
or U13219 (N_13219,N_11291,N_11434);
nor U13220 (N_13220,N_11713,N_11368);
or U13221 (N_13221,N_10402,N_10410);
xor U13222 (N_13222,N_11490,N_11160);
xnor U13223 (N_13223,N_10932,N_11064);
nand U13224 (N_13224,N_10721,N_10078);
xnor U13225 (N_13225,N_11667,N_11687);
and U13226 (N_13226,N_11731,N_10516);
xnor U13227 (N_13227,N_11195,N_10330);
and U13228 (N_13228,N_10867,N_11533);
xor U13229 (N_13229,N_10508,N_11552);
nand U13230 (N_13230,N_11222,N_11375);
and U13231 (N_13231,N_11195,N_10410);
or U13232 (N_13232,N_10680,N_10382);
or U13233 (N_13233,N_11683,N_11415);
nor U13234 (N_13234,N_11941,N_11549);
nand U13235 (N_13235,N_10157,N_11546);
or U13236 (N_13236,N_10867,N_11445);
xor U13237 (N_13237,N_10671,N_11337);
and U13238 (N_13238,N_10349,N_10781);
xor U13239 (N_13239,N_11484,N_11333);
and U13240 (N_13240,N_11239,N_10563);
nor U13241 (N_13241,N_11374,N_10816);
xnor U13242 (N_13242,N_10742,N_11399);
nor U13243 (N_13243,N_11596,N_10679);
or U13244 (N_13244,N_11585,N_10849);
or U13245 (N_13245,N_10578,N_11823);
nor U13246 (N_13246,N_10292,N_11290);
or U13247 (N_13247,N_11081,N_10170);
and U13248 (N_13248,N_11683,N_10697);
or U13249 (N_13249,N_11161,N_10834);
and U13250 (N_13250,N_11610,N_11665);
or U13251 (N_13251,N_11451,N_10907);
or U13252 (N_13252,N_10048,N_10328);
xor U13253 (N_13253,N_11907,N_10033);
nor U13254 (N_13254,N_10530,N_10764);
nor U13255 (N_13255,N_11189,N_11092);
nand U13256 (N_13256,N_10039,N_10091);
xor U13257 (N_13257,N_11697,N_10912);
xor U13258 (N_13258,N_11783,N_11431);
or U13259 (N_13259,N_10762,N_10180);
and U13260 (N_13260,N_11220,N_10734);
and U13261 (N_13261,N_11581,N_10866);
and U13262 (N_13262,N_11781,N_10866);
and U13263 (N_13263,N_11950,N_11561);
and U13264 (N_13264,N_11854,N_11807);
xor U13265 (N_13265,N_10518,N_10302);
or U13266 (N_13266,N_10600,N_10489);
nand U13267 (N_13267,N_10230,N_11259);
nand U13268 (N_13268,N_11802,N_10574);
nand U13269 (N_13269,N_11329,N_11845);
nand U13270 (N_13270,N_11190,N_10341);
or U13271 (N_13271,N_10378,N_10281);
nor U13272 (N_13272,N_10507,N_11063);
nor U13273 (N_13273,N_10060,N_10369);
or U13274 (N_13274,N_10902,N_10842);
and U13275 (N_13275,N_11703,N_10943);
xnor U13276 (N_13276,N_11831,N_10777);
and U13277 (N_13277,N_11582,N_10059);
and U13278 (N_13278,N_11871,N_10301);
nand U13279 (N_13279,N_10616,N_11028);
xor U13280 (N_13280,N_11481,N_10381);
and U13281 (N_13281,N_11667,N_10324);
and U13282 (N_13282,N_11843,N_11960);
or U13283 (N_13283,N_11586,N_10280);
or U13284 (N_13284,N_10489,N_11368);
or U13285 (N_13285,N_11327,N_10226);
and U13286 (N_13286,N_11223,N_10236);
or U13287 (N_13287,N_10243,N_11178);
xnor U13288 (N_13288,N_11373,N_11357);
nor U13289 (N_13289,N_10794,N_10247);
xor U13290 (N_13290,N_11261,N_10921);
and U13291 (N_13291,N_10511,N_11866);
and U13292 (N_13292,N_11914,N_11268);
nor U13293 (N_13293,N_10561,N_10548);
and U13294 (N_13294,N_11736,N_10530);
xor U13295 (N_13295,N_10372,N_10111);
xor U13296 (N_13296,N_10529,N_11607);
xor U13297 (N_13297,N_10888,N_11708);
nand U13298 (N_13298,N_10446,N_10168);
and U13299 (N_13299,N_11919,N_10288);
nor U13300 (N_13300,N_10339,N_11303);
and U13301 (N_13301,N_10159,N_11989);
or U13302 (N_13302,N_10647,N_10107);
or U13303 (N_13303,N_10171,N_11208);
nor U13304 (N_13304,N_11644,N_10542);
or U13305 (N_13305,N_11586,N_11526);
and U13306 (N_13306,N_10780,N_11944);
and U13307 (N_13307,N_10105,N_11146);
xor U13308 (N_13308,N_10499,N_11154);
xnor U13309 (N_13309,N_11966,N_10381);
and U13310 (N_13310,N_10114,N_11213);
and U13311 (N_13311,N_10983,N_11387);
nor U13312 (N_13312,N_11628,N_11821);
xor U13313 (N_13313,N_10732,N_11349);
nor U13314 (N_13314,N_10209,N_11145);
nor U13315 (N_13315,N_11810,N_10117);
xnor U13316 (N_13316,N_10548,N_11421);
xor U13317 (N_13317,N_10560,N_10266);
or U13318 (N_13318,N_10827,N_10507);
xor U13319 (N_13319,N_10629,N_11558);
and U13320 (N_13320,N_10600,N_10625);
or U13321 (N_13321,N_11841,N_11437);
nor U13322 (N_13322,N_10082,N_11955);
and U13323 (N_13323,N_10026,N_11845);
nor U13324 (N_13324,N_11632,N_11948);
and U13325 (N_13325,N_10813,N_11816);
nor U13326 (N_13326,N_10851,N_11175);
nor U13327 (N_13327,N_10685,N_10708);
and U13328 (N_13328,N_10743,N_11939);
nor U13329 (N_13329,N_11255,N_10176);
xor U13330 (N_13330,N_11204,N_11655);
or U13331 (N_13331,N_10104,N_10432);
nor U13332 (N_13332,N_11044,N_11136);
nor U13333 (N_13333,N_10811,N_11807);
or U13334 (N_13334,N_10710,N_11423);
and U13335 (N_13335,N_11233,N_10545);
xnor U13336 (N_13336,N_11926,N_10942);
nand U13337 (N_13337,N_11332,N_11466);
nand U13338 (N_13338,N_11267,N_10021);
and U13339 (N_13339,N_11315,N_10596);
xor U13340 (N_13340,N_10117,N_11340);
nor U13341 (N_13341,N_11664,N_11338);
and U13342 (N_13342,N_11975,N_11199);
or U13343 (N_13343,N_11937,N_11717);
nand U13344 (N_13344,N_10765,N_11445);
nor U13345 (N_13345,N_10018,N_11553);
nor U13346 (N_13346,N_10137,N_10896);
xnor U13347 (N_13347,N_11330,N_10044);
nand U13348 (N_13348,N_11860,N_10378);
or U13349 (N_13349,N_10577,N_10906);
nor U13350 (N_13350,N_11339,N_11513);
nor U13351 (N_13351,N_10909,N_11897);
or U13352 (N_13352,N_10155,N_11875);
xor U13353 (N_13353,N_10323,N_11779);
xnor U13354 (N_13354,N_10088,N_11313);
xor U13355 (N_13355,N_10963,N_11851);
xnor U13356 (N_13356,N_11548,N_11267);
xnor U13357 (N_13357,N_10595,N_10949);
xnor U13358 (N_13358,N_10115,N_11627);
nand U13359 (N_13359,N_10240,N_10576);
or U13360 (N_13360,N_10021,N_11726);
xnor U13361 (N_13361,N_11936,N_11687);
and U13362 (N_13362,N_11288,N_10772);
nand U13363 (N_13363,N_10766,N_11546);
xor U13364 (N_13364,N_11654,N_11123);
xor U13365 (N_13365,N_10535,N_10194);
nand U13366 (N_13366,N_11490,N_10722);
nor U13367 (N_13367,N_10571,N_11810);
nand U13368 (N_13368,N_10021,N_10910);
xor U13369 (N_13369,N_11632,N_11646);
and U13370 (N_13370,N_11385,N_11167);
nor U13371 (N_13371,N_11010,N_11508);
xor U13372 (N_13372,N_11320,N_11775);
or U13373 (N_13373,N_10906,N_10575);
and U13374 (N_13374,N_10499,N_11442);
xnor U13375 (N_13375,N_10695,N_10745);
and U13376 (N_13376,N_11910,N_10715);
nand U13377 (N_13377,N_10023,N_11598);
xor U13378 (N_13378,N_11389,N_11506);
and U13379 (N_13379,N_11977,N_11129);
nor U13380 (N_13380,N_11648,N_10277);
and U13381 (N_13381,N_11719,N_11698);
and U13382 (N_13382,N_11760,N_10319);
nor U13383 (N_13383,N_11896,N_11981);
or U13384 (N_13384,N_10139,N_10159);
nand U13385 (N_13385,N_10141,N_11257);
or U13386 (N_13386,N_10363,N_11539);
and U13387 (N_13387,N_11102,N_10014);
xnor U13388 (N_13388,N_10381,N_10650);
nand U13389 (N_13389,N_10240,N_10982);
xnor U13390 (N_13390,N_11841,N_10424);
xnor U13391 (N_13391,N_11888,N_11471);
or U13392 (N_13392,N_11349,N_10234);
and U13393 (N_13393,N_10961,N_10989);
nand U13394 (N_13394,N_10152,N_11582);
nor U13395 (N_13395,N_11404,N_10050);
or U13396 (N_13396,N_11681,N_10768);
or U13397 (N_13397,N_10825,N_10406);
nand U13398 (N_13398,N_10328,N_10596);
xnor U13399 (N_13399,N_10626,N_11408);
and U13400 (N_13400,N_10640,N_11120);
and U13401 (N_13401,N_10643,N_10891);
or U13402 (N_13402,N_10288,N_10530);
nand U13403 (N_13403,N_10019,N_10500);
nor U13404 (N_13404,N_11019,N_10173);
and U13405 (N_13405,N_11746,N_11198);
and U13406 (N_13406,N_10237,N_11233);
nor U13407 (N_13407,N_10439,N_10676);
or U13408 (N_13408,N_10290,N_10930);
nand U13409 (N_13409,N_10300,N_11407);
xnor U13410 (N_13410,N_10582,N_11248);
or U13411 (N_13411,N_10198,N_11862);
nand U13412 (N_13412,N_10149,N_10232);
nand U13413 (N_13413,N_11426,N_11822);
or U13414 (N_13414,N_11520,N_11789);
nor U13415 (N_13415,N_10125,N_11911);
nor U13416 (N_13416,N_10906,N_10361);
or U13417 (N_13417,N_11677,N_10790);
nand U13418 (N_13418,N_11244,N_10357);
nor U13419 (N_13419,N_11468,N_10093);
or U13420 (N_13420,N_11353,N_11344);
xnor U13421 (N_13421,N_11721,N_11324);
and U13422 (N_13422,N_10997,N_11801);
xor U13423 (N_13423,N_11338,N_10349);
nand U13424 (N_13424,N_11864,N_11059);
or U13425 (N_13425,N_11993,N_11121);
xnor U13426 (N_13426,N_10354,N_11618);
xor U13427 (N_13427,N_11865,N_11238);
xor U13428 (N_13428,N_11823,N_11043);
and U13429 (N_13429,N_11357,N_11075);
nand U13430 (N_13430,N_11308,N_11371);
or U13431 (N_13431,N_10467,N_11516);
xnor U13432 (N_13432,N_10222,N_10545);
and U13433 (N_13433,N_10235,N_10422);
nand U13434 (N_13434,N_11163,N_11592);
nor U13435 (N_13435,N_10386,N_10822);
nor U13436 (N_13436,N_10702,N_10532);
xnor U13437 (N_13437,N_10911,N_11168);
nand U13438 (N_13438,N_10085,N_11002);
xnor U13439 (N_13439,N_10963,N_10870);
and U13440 (N_13440,N_11557,N_11884);
and U13441 (N_13441,N_11101,N_10567);
and U13442 (N_13442,N_10770,N_11609);
and U13443 (N_13443,N_11384,N_10871);
xor U13444 (N_13444,N_11032,N_10328);
and U13445 (N_13445,N_10341,N_11215);
nand U13446 (N_13446,N_11789,N_10071);
or U13447 (N_13447,N_11768,N_10047);
and U13448 (N_13448,N_11221,N_11004);
or U13449 (N_13449,N_10191,N_10401);
or U13450 (N_13450,N_11711,N_11827);
nor U13451 (N_13451,N_11982,N_10075);
nor U13452 (N_13452,N_11315,N_10494);
and U13453 (N_13453,N_11548,N_11554);
and U13454 (N_13454,N_11304,N_11323);
or U13455 (N_13455,N_11007,N_11404);
nor U13456 (N_13456,N_11599,N_11141);
and U13457 (N_13457,N_10025,N_10538);
xnor U13458 (N_13458,N_10353,N_10745);
xnor U13459 (N_13459,N_10373,N_10899);
and U13460 (N_13460,N_10018,N_11238);
nor U13461 (N_13461,N_10154,N_10453);
xor U13462 (N_13462,N_11225,N_11199);
nor U13463 (N_13463,N_10048,N_10827);
or U13464 (N_13464,N_11747,N_11215);
xnor U13465 (N_13465,N_11777,N_10362);
and U13466 (N_13466,N_10762,N_11993);
and U13467 (N_13467,N_10038,N_10640);
nor U13468 (N_13468,N_10729,N_11732);
and U13469 (N_13469,N_11348,N_11954);
nor U13470 (N_13470,N_10863,N_11789);
and U13471 (N_13471,N_11982,N_10245);
nand U13472 (N_13472,N_11780,N_10121);
nand U13473 (N_13473,N_10404,N_10074);
xor U13474 (N_13474,N_10128,N_11685);
nand U13475 (N_13475,N_10122,N_11836);
and U13476 (N_13476,N_10404,N_10948);
nor U13477 (N_13477,N_10712,N_10928);
and U13478 (N_13478,N_11595,N_10600);
nor U13479 (N_13479,N_10567,N_10794);
and U13480 (N_13480,N_11949,N_10947);
nand U13481 (N_13481,N_10896,N_10701);
xor U13482 (N_13482,N_10375,N_10047);
nor U13483 (N_13483,N_11873,N_10111);
nand U13484 (N_13484,N_11457,N_10919);
xor U13485 (N_13485,N_10949,N_11747);
xor U13486 (N_13486,N_11674,N_10484);
xnor U13487 (N_13487,N_11409,N_10080);
or U13488 (N_13488,N_10064,N_11804);
nor U13489 (N_13489,N_10809,N_11995);
nand U13490 (N_13490,N_11944,N_11020);
and U13491 (N_13491,N_11465,N_11448);
xor U13492 (N_13492,N_11265,N_11590);
and U13493 (N_13493,N_10519,N_11687);
xnor U13494 (N_13494,N_11325,N_11052);
xnor U13495 (N_13495,N_11181,N_10548);
nor U13496 (N_13496,N_10395,N_11449);
nor U13497 (N_13497,N_11454,N_11489);
and U13498 (N_13498,N_10728,N_10071);
xnor U13499 (N_13499,N_10812,N_10344);
nor U13500 (N_13500,N_11596,N_10157);
nand U13501 (N_13501,N_11066,N_10407);
xor U13502 (N_13502,N_10467,N_10398);
xor U13503 (N_13503,N_10713,N_10265);
xor U13504 (N_13504,N_11995,N_11568);
xnor U13505 (N_13505,N_11107,N_11684);
xnor U13506 (N_13506,N_11881,N_11636);
xnor U13507 (N_13507,N_10151,N_10196);
xnor U13508 (N_13508,N_11335,N_10606);
xor U13509 (N_13509,N_11373,N_10729);
nand U13510 (N_13510,N_11520,N_11900);
and U13511 (N_13511,N_11892,N_10237);
and U13512 (N_13512,N_11416,N_11014);
xor U13513 (N_13513,N_10961,N_10388);
and U13514 (N_13514,N_10636,N_10107);
nor U13515 (N_13515,N_11749,N_11190);
nor U13516 (N_13516,N_10686,N_10672);
or U13517 (N_13517,N_10877,N_10378);
nand U13518 (N_13518,N_10753,N_10169);
or U13519 (N_13519,N_10240,N_10926);
or U13520 (N_13520,N_10494,N_11000);
and U13521 (N_13521,N_11191,N_10064);
xor U13522 (N_13522,N_10855,N_11272);
nand U13523 (N_13523,N_11607,N_11641);
nor U13524 (N_13524,N_10735,N_11706);
nand U13525 (N_13525,N_10232,N_10529);
nor U13526 (N_13526,N_11813,N_10291);
and U13527 (N_13527,N_11068,N_10529);
nor U13528 (N_13528,N_10520,N_10118);
nor U13529 (N_13529,N_11310,N_10474);
nand U13530 (N_13530,N_10965,N_10938);
xor U13531 (N_13531,N_10214,N_10952);
xnor U13532 (N_13532,N_11919,N_11190);
nand U13533 (N_13533,N_10935,N_10088);
xor U13534 (N_13534,N_11065,N_11664);
or U13535 (N_13535,N_10069,N_10897);
or U13536 (N_13536,N_10198,N_11587);
and U13537 (N_13537,N_11184,N_11721);
or U13538 (N_13538,N_10933,N_10682);
or U13539 (N_13539,N_11152,N_11255);
and U13540 (N_13540,N_10294,N_10738);
nor U13541 (N_13541,N_11665,N_10244);
xnor U13542 (N_13542,N_11918,N_11716);
nand U13543 (N_13543,N_11235,N_10750);
or U13544 (N_13544,N_11524,N_10129);
or U13545 (N_13545,N_11378,N_11308);
and U13546 (N_13546,N_10703,N_11809);
nor U13547 (N_13547,N_11311,N_11523);
xnor U13548 (N_13548,N_11764,N_11816);
nand U13549 (N_13549,N_11734,N_11292);
and U13550 (N_13550,N_10773,N_11007);
or U13551 (N_13551,N_10487,N_10836);
nor U13552 (N_13552,N_11300,N_10039);
xnor U13553 (N_13553,N_10875,N_11874);
nor U13554 (N_13554,N_11337,N_11716);
or U13555 (N_13555,N_11944,N_10703);
xor U13556 (N_13556,N_10322,N_11456);
nand U13557 (N_13557,N_11490,N_11423);
xor U13558 (N_13558,N_11466,N_11740);
nor U13559 (N_13559,N_11388,N_10361);
xnor U13560 (N_13560,N_11463,N_10898);
or U13561 (N_13561,N_10020,N_10703);
nand U13562 (N_13562,N_10774,N_11912);
and U13563 (N_13563,N_10757,N_10903);
and U13564 (N_13564,N_11159,N_10015);
or U13565 (N_13565,N_10378,N_10444);
nor U13566 (N_13566,N_10151,N_11896);
and U13567 (N_13567,N_10830,N_11604);
or U13568 (N_13568,N_10084,N_11072);
nor U13569 (N_13569,N_11146,N_11169);
nor U13570 (N_13570,N_10563,N_11922);
nand U13571 (N_13571,N_10630,N_11126);
nor U13572 (N_13572,N_10282,N_11603);
or U13573 (N_13573,N_11535,N_10528);
and U13574 (N_13574,N_11743,N_11878);
xnor U13575 (N_13575,N_11842,N_10558);
or U13576 (N_13576,N_10887,N_11395);
or U13577 (N_13577,N_11046,N_11829);
nand U13578 (N_13578,N_10218,N_11183);
nor U13579 (N_13579,N_11710,N_11979);
nor U13580 (N_13580,N_10483,N_10330);
nand U13581 (N_13581,N_11467,N_11646);
and U13582 (N_13582,N_10032,N_10409);
nor U13583 (N_13583,N_10969,N_10373);
or U13584 (N_13584,N_11673,N_10354);
or U13585 (N_13585,N_10966,N_11568);
nor U13586 (N_13586,N_10849,N_10751);
nor U13587 (N_13587,N_10973,N_11986);
xor U13588 (N_13588,N_11926,N_11383);
xor U13589 (N_13589,N_11234,N_10029);
and U13590 (N_13590,N_10762,N_11273);
xor U13591 (N_13591,N_11535,N_11699);
or U13592 (N_13592,N_10863,N_11781);
nand U13593 (N_13593,N_11921,N_10179);
nor U13594 (N_13594,N_10535,N_10349);
nand U13595 (N_13595,N_11184,N_10401);
or U13596 (N_13596,N_11511,N_11043);
or U13597 (N_13597,N_11676,N_10874);
and U13598 (N_13598,N_10650,N_11964);
xor U13599 (N_13599,N_10625,N_10149);
nor U13600 (N_13600,N_10180,N_11452);
and U13601 (N_13601,N_10230,N_10221);
xor U13602 (N_13602,N_10160,N_11658);
nand U13603 (N_13603,N_10573,N_10445);
nor U13604 (N_13604,N_11072,N_10390);
and U13605 (N_13605,N_10100,N_11337);
xor U13606 (N_13606,N_11265,N_11134);
nor U13607 (N_13607,N_10415,N_11939);
nor U13608 (N_13608,N_10361,N_10234);
and U13609 (N_13609,N_11422,N_10698);
and U13610 (N_13610,N_11456,N_11979);
and U13611 (N_13611,N_11086,N_10592);
nor U13612 (N_13612,N_11799,N_10092);
nand U13613 (N_13613,N_10298,N_10397);
nand U13614 (N_13614,N_11957,N_10620);
nand U13615 (N_13615,N_11615,N_10545);
nand U13616 (N_13616,N_11754,N_10087);
and U13617 (N_13617,N_10618,N_10450);
or U13618 (N_13618,N_10056,N_10877);
nor U13619 (N_13619,N_11554,N_11956);
or U13620 (N_13620,N_11944,N_10953);
nor U13621 (N_13621,N_10651,N_11628);
nor U13622 (N_13622,N_11405,N_11857);
or U13623 (N_13623,N_10302,N_11893);
and U13624 (N_13624,N_11241,N_10189);
xnor U13625 (N_13625,N_10586,N_11778);
and U13626 (N_13626,N_11576,N_10359);
nor U13627 (N_13627,N_11924,N_10255);
nor U13628 (N_13628,N_11139,N_10562);
nor U13629 (N_13629,N_11322,N_10369);
xnor U13630 (N_13630,N_10650,N_10494);
nor U13631 (N_13631,N_11037,N_10280);
nand U13632 (N_13632,N_11754,N_10955);
and U13633 (N_13633,N_11481,N_10087);
xnor U13634 (N_13634,N_10092,N_11352);
and U13635 (N_13635,N_10180,N_11045);
nand U13636 (N_13636,N_10920,N_11833);
nor U13637 (N_13637,N_11629,N_11012);
or U13638 (N_13638,N_10442,N_10235);
and U13639 (N_13639,N_10403,N_10503);
xnor U13640 (N_13640,N_10936,N_10016);
nand U13641 (N_13641,N_11274,N_10439);
or U13642 (N_13642,N_11448,N_10858);
nor U13643 (N_13643,N_11559,N_11163);
nor U13644 (N_13644,N_11200,N_11065);
xnor U13645 (N_13645,N_10727,N_10562);
nand U13646 (N_13646,N_10671,N_11383);
nand U13647 (N_13647,N_10580,N_11158);
nand U13648 (N_13648,N_11604,N_11731);
nand U13649 (N_13649,N_10450,N_10675);
and U13650 (N_13650,N_11559,N_10467);
or U13651 (N_13651,N_10973,N_11132);
and U13652 (N_13652,N_11382,N_11838);
and U13653 (N_13653,N_11149,N_11612);
nor U13654 (N_13654,N_10735,N_10393);
nand U13655 (N_13655,N_10166,N_10817);
and U13656 (N_13656,N_11034,N_10524);
nand U13657 (N_13657,N_11549,N_10030);
or U13658 (N_13658,N_11807,N_10294);
nor U13659 (N_13659,N_11773,N_11761);
nand U13660 (N_13660,N_10022,N_10403);
nand U13661 (N_13661,N_10658,N_11401);
nand U13662 (N_13662,N_11621,N_10661);
or U13663 (N_13663,N_11068,N_10724);
or U13664 (N_13664,N_11167,N_11831);
and U13665 (N_13665,N_11568,N_10009);
and U13666 (N_13666,N_10149,N_11679);
or U13667 (N_13667,N_11140,N_10889);
nor U13668 (N_13668,N_10530,N_10302);
or U13669 (N_13669,N_11480,N_10112);
nand U13670 (N_13670,N_11999,N_11994);
nand U13671 (N_13671,N_11796,N_10045);
and U13672 (N_13672,N_10899,N_10491);
or U13673 (N_13673,N_11538,N_10658);
nand U13674 (N_13674,N_10715,N_10981);
or U13675 (N_13675,N_11473,N_11358);
xnor U13676 (N_13676,N_11731,N_10419);
and U13677 (N_13677,N_11360,N_10434);
xnor U13678 (N_13678,N_11287,N_10493);
nand U13679 (N_13679,N_10979,N_10051);
and U13680 (N_13680,N_11502,N_11447);
nor U13681 (N_13681,N_10263,N_10485);
or U13682 (N_13682,N_10701,N_11716);
or U13683 (N_13683,N_10654,N_11280);
nand U13684 (N_13684,N_10399,N_11650);
nor U13685 (N_13685,N_10129,N_10482);
xor U13686 (N_13686,N_11143,N_10215);
or U13687 (N_13687,N_10546,N_10402);
nor U13688 (N_13688,N_10098,N_10656);
xnor U13689 (N_13689,N_10875,N_11600);
xnor U13690 (N_13690,N_11737,N_11175);
nand U13691 (N_13691,N_10695,N_10469);
nor U13692 (N_13692,N_10619,N_11834);
nor U13693 (N_13693,N_11754,N_11735);
or U13694 (N_13694,N_11055,N_10579);
xor U13695 (N_13695,N_10284,N_10463);
nand U13696 (N_13696,N_10014,N_10725);
xor U13697 (N_13697,N_10547,N_10266);
and U13698 (N_13698,N_11045,N_11683);
nor U13699 (N_13699,N_11736,N_11772);
nor U13700 (N_13700,N_11689,N_10703);
xor U13701 (N_13701,N_11917,N_11872);
nand U13702 (N_13702,N_11188,N_11169);
or U13703 (N_13703,N_11067,N_10848);
and U13704 (N_13704,N_11664,N_11790);
nor U13705 (N_13705,N_10451,N_11119);
xor U13706 (N_13706,N_10298,N_11884);
nor U13707 (N_13707,N_10578,N_11058);
xor U13708 (N_13708,N_10789,N_11312);
xnor U13709 (N_13709,N_10164,N_11686);
nor U13710 (N_13710,N_10506,N_11801);
nor U13711 (N_13711,N_10443,N_11704);
nand U13712 (N_13712,N_11946,N_10189);
xnor U13713 (N_13713,N_10830,N_10471);
nand U13714 (N_13714,N_10689,N_10251);
and U13715 (N_13715,N_10939,N_10978);
nor U13716 (N_13716,N_11758,N_10580);
and U13717 (N_13717,N_10788,N_10018);
or U13718 (N_13718,N_10449,N_11990);
nand U13719 (N_13719,N_11313,N_11781);
nand U13720 (N_13720,N_11468,N_11795);
and U13721 (N_13721,N_11666,N_11836);
nand U13722 (N_13722,N_10920,N_10450);
nand U13723 (N_13723,N_10249,N_10053);
and U13724 (N_13724,N_10106,N_11093);
nand U13725 (N_13725,N_11991,N_10593);
and U13726 (N_13726,N_10184,N_10566);
xnor U13727 (N_13727,N_11951,N_10494);
and U13728 (N_13728,N_11915,N_11447);
or U13729 (N_13729,N_11171,N_10813);
and U13730 (N_13730,N_11990,N_10429);
nand U13731 (N_13731,N_10506,N_10200);
xor U13732 (N_13732,N_10331,N_10376);
or U13733 (N_13733,N_11603,N_10822);
nor U13734 (N_13734,N_11028,N_10120);
or U13735 (N_13735,N_10092,N_10064);
nand U13736 (N_13736,N_10931,N_11003);
xnor U13737 (N_13737,N_11542,N_11174);
or U13738 (N_13738,N_11202,N_11433);
nor U13739 (N_13739,N_10022,N_11148);
and U13740 (N_13740,N_11954,N_10430);
and U13741 (N_13741,N_11988,N_11786);
nor U13742 (N_13742,N_11913,N_10526);
xor U13743 (N_13743,N_11538,N_10308);
xor U13744 (N_13744,N_11739,N_10504);
or U13745 (N_13745,N_11993,N_11648);
or U13746 (N_13746,N_11375,N_11057);
or U13747 (N_13747,N_11398,N_11362);
and U13748 (N_13748,N_10223,N_11225);
nand U13749 (N_13749,N_10512,N_10019);
xnor U13750 (N_13750,N_10363,N_11443);
and U13751 (N_13751,N_11899,N_11397);
nand U13752 (N_13752,N_11696,N_11796);
and U13753 (N_13753,N_10692,N_11390);
nor U13754 (N_13754,N_11863,N_11186);
nand U13755 (N_13755,N_11653,N_10518);
nand U13756 (N_13756,N_11277,N_10846);
and U13757 (N_13757,N_10644,N_11818);
or U13758 (N_13758,N_10962,N_10193);
or U13759 (N_13759,N_10398,N_10206);
or U13760 (N_13760,N_10218,N_11495);
xnor U13761 (N_13761,N_11484,N_11892);
xor U13762 (N_13762,N_10588,N_11375);
or U13763 (N_13763,N_11503,N_11523);
and U13764 (N_13764,N_11249,N_10910);
or U13765 (N_13765,N_10119,N_10029);
and U13766 (N_13766,N_10273,N_10794);
nor U13767 (N_13767,N_11515,N_10949);
nand U13768 (N_13768,N_10628,N_10440);
nand U13769 (N_13769,N_10333,N_11314);
xnor U13770 (N_13770,N_11185,N_10382);
xnor U13771 (N_13771,N_10319,N_10013);
xnor U13772 (N_13772,N_10286,N_10912);
xnor U13773 (N_13773,N_10534,N_10038);
or U13774 (N_13774,N_11216,N_11210);
or U13775 (N_13775,N_11843,N_11805);
and U13776 (N_13776,N_10961,N_11902);
or U13777 (N_13777,N_10304,N_11364);
xnor U13778 (N_13778,N_11899,N_11344);
or U13779 (N_13779,N_10871,N_10821);
nand U13780 (N_13780,N_10091,N_10201);
nand U13781 (N_13781,N_10867,N_10431);
nor U13782 (N_13782,N_10937,N_10764);
or U13783 (N_13783,N_11687,N_11868);
nand U13784 (N_13784,N_10449,N_11342);
or U13785 (N_13785,N_11388,N_11832);
xor U13786 (N_13786,N_11894,N_11260);
xnor U13787 (N_13787,N_11285,N_11538);
or U13788 (N_13788,N_10230,N_11675);
or U13789 (N_13789,N_11110,N_11206);
nor U13790 (N_13790,N_10241,N_11858);
and U13791 (N_13791,N_11855,N_10157);
xnor U13792 (N_13792,N_10627,N_11129);
nor U13793 (N_13793,N_10951,N_10933);
and U13794 (N_13794,N_10209,N_11903);
nand U13795 (N_13795,N_10038,N_10247);
nand U13796 (N_13796,N_11582,N_10696);
nand U13797 (N_13797,N_10835,N_10140);
and U13798 (N_13798,N_10014,N_10475);
nand U13799 (N_13799,N_10157,N_11605);
or U13800 (N_13800,N_10341,N_10880);
nand U13801 (N_13801,N_11794,N_11790);
or U13802 (N_13802,N_11524,N_10720);
and U13803 (N_13803,N_11924,N_11339);
xnor U13804 (N_13804,N_10339,N_11201);
xor U13805 (N_13805,N_11198,N_10776);
xnor U13806 (N_13806,N_10082,N_11058);
or U13807 (N_13807,N_10957,N_11128);
xor U13808 (N_13808,N_11034,N_11732);
nand U13809 (N_13809,N_11948,N_11704);
and U13810 (N_13810,N_11425,N_11012);
or U13811 (N_13811,N_10124,N_11914);
nor U13812 (N_13812,N_10004,N_10240);
xnor U13813 (N_13813,N_11007,N_10633);
xor U13814 (N_13814,N_11829,N_10380);
or U13815 (N_13815,N_10601,N_10518);
or U13816 (N_13816,N_11764,N_11315);
xnor U13817 (N_13817,N_10017,N_10999);
or U13818 (N_13818,N_10843,N_10612);
nor U13819 (N_13819,N_10498,N_10137);
nor U13820 (N_13820,N_11584,N_11697);
or U13821 (N_13821,N_10695,N_10621);
and U13822 (N_13822,N_11365,N_11576);
or U13823 (N_13823,N_10531,N_11823);
or U13824 (N_13824,N_11353,N_11178);
or U13825 (N_13825,N_10008,N_10387);
nor U13826 (N_13826,N_10396,N_10937);
nor U13827 (N_13827,N_10462,N_11749);
and U13828 (N_13828,N_11417,N_11247);
nor U13829 (N_13829,N_11479,N_11169);
nand U13830 (N_13830,N_11493,N_10316);
xor U13831 (N_13831,N_11646,N_10011);
xnor U13832 (N_13832,N_11097,N_10722);
and U13833 (N_13833,N_11310,N_11096);
xnor U13834 (N_13834,N_11600,N_11876);
nor U13835 (N_13835,N_10414,N_10508);
xor U13836 (N_13836,N_10547,N_11505);
and U13837 (N_13837,N_10602,N_11852);
xor U13838 (N_13838,N_10552,N_10158);
and U13839 (N_13839,N_10551,N_11206);
nand U13840 (N_13840,N_10578,N_11862);
or U13841 (N_13841,N_10195,N_11900);
nand U13842 (N_13842,N_11528,N_11157);
xor U13843 (N_13843,N_10735,N_11466);
nand U13844 (N_13844,N_11770,N_10873);
nor U13845 (N_13845,N_10441,N_10974);
xor U13846 (N_13846,N_10593,N_10801);
and U13847 (N_13847,N_11855,N_11667);
nand U13848 (N_13848,N_10062,N_10310);
or U13849 (N_13849,N_10992,N_10610);
xnor U13850 (N_13850,N_11866,N_11416);
nor U13851 (N_13851,N_10079,N_10310);
or U13852 (N_13852,N_11682,N_10823);
xnor U13853 (N_13853,N_10474,N_11375);
nand U13854 (N_13854,N_10141,N_11468);
or U13855 (N_13855,N_11312,N_10552);
or U13856 (N_13856,N_10075,N_10969);
xor U13857 (N_13857,N_10403,N_10311);
or U13858 (N_13858,N_10831,N_10733);
or U13859 (N_13859,N_11560,N_11026);
or U13860 (N_13860,N_10288,N_11805);
and U13861 (N_13861,N_11370,N_11265);
nor U13862 (N_13862,N_10142,N_11750);
and U13863 (N_13863,N_11238,N_11942);
and U13864 (N_13864,N_10217,N_10262);
or U13865 (N_13865,N_11767,N_11508);
nand U13866 (N_13866,N_11575,N_10612);
or U13867 (N_13867,N_11736,N_10837);
or U13868 (N_13868,N_11757,N_11719);
nand U13869 (N_13869,N_10172,N_10627);
nor U13870 (N_13870,N_10118,N_10587);
or U13871 (N_13871,N_11449,N_11286);
and U13872 (N_13872,N_11799,N_10258);
nor U13873 (N_13873,N_11156,N_10949);
xnor U13874 (N_13874,N_11431,N_11530);
or U13875 (N_13875,N_11551,N_11280);
or U13876 (N_13876,N_11643,N_10871);
or U13877 (N_13877,N_10149,N_11788);
or U13878 (N_13878,N_11758,N_10212);
and U13879 (N_13879,N_10909,N_10666);
nand U13880 (N_13880,N_11800,N_10791);
nand U13881 (N_13881,N_11813,N_11684);
nor U13882 (N_13882,N_11832,N_10760);
nor U13883 (N_13883,N_11583,N_10035);
xnor U13884 (N_13884,N_11026,N_10280);
nor U13885 (N_13885,N_11257,N_10684);
or U13886 (N_13886,N_11982,N_10449);
and U13887 (N_13887,N_10693,N_11522);
nor U13888 (N_13888,N_11695,N_11580);
or U13889 (N_13889,N_11006,N_11745);
nor U13890 (N_13890,N_10290,N_10508);
nor U13891 (N_13891,N_10240,N_11186);
and U13892 (N_13892,N_10476,N_10678);
or U13893 (N_13893,N_10430,N_10315);
nand U13894 (N_13894,N_10142,N_11715);
xor U13895 (N_13895,N_11568,N_11329);
and U13896 (N_13896,N_11072,N_10566);
or U13897 (N_13897,N_11612,N_10372);
xor U13898 (N_13898,N_11685,N_11221);
xor U13899 (N_13899,N_11778,N_10589);
and U13900 (N_13900,N_11172,N_10112);
or U13901 (N_13901,N_11160,N_11248);
xnor U13902 (N_13902,N_11800,N_10135);
xnor U13903 (N_13903,N_10878,N_10222);
and U13904 (N_13904,N_11712,N_11156);
or U13905 (N_13905,N_10773,N_10976);
xor U13906 (N_13906,N_11216,N_11342);
nand U13907 (N_13907,N_10433,N_10852);
and U13908 (N_13908,N_10692,N_10214);
nor U13909 (N_13909,N_11251,N_10675);
nor U13910 (N_13910,N_11452,N_10220);
and U13911 (N_13911,N_10086,N_11160);
nor U13912 (N_13912,N_11719,N_10754);
nand U13913 (N_13913,N_10764,N_10097);
and U13914 (N_13914,N_11354,N_11400);
nor U13915 (N_13915,N_10676,N_11049);
nor U13916 (N_13916,N_11301,N_11916);
xnor U13917 (N_13917,N_10745,N_11810);
xor U13918 (N_13918,N_11339,N_10539);
and U13919 (N_13919,N_11375,N_10275);
nand U13920 (N_13920,N_11132,N_11125);
xor U13921 (N_13921,N_10025,N_11150);
nor U13922 (N_13922,N_10497,N_11538);
xnor U13923 (N_13923,N_10514,N_10547);
xnor U13924 (N_13924,N_11566,N_11223);
nand U13925 (N_13925,N_11338,N_10184);
xor U13926 (N_13926,N_10709,N_11776);
nor U13927 (N_13927,N_10941,N_10799);
or U13928 (N_13928,N_10215,N_10589);
nand U13929 (N_13929,N_11234,N_10700);
nand U13930 (N_13930,N_10094,N_11977);
or U13931 (N_13931,N_11621,N_10277);
or U13932 (N_13932,N_11830,N_11668);
and U13933 (N_13933,N_11955,N_10724);
xor U13934 (N_13934,N_10773,N_11510);
xnor U13935 (N_13935,N_11002,N_11106);
nand U13936 (N_13936,N_11277,N_10470);
nor U13937 (N_13937,N_10509,N_10135);
xor U13938 (N_13938,N_10878,N_11304);
and U13939 (N_13939,N_11523,N_11406);
or U13940 (N_13940,N_11226,N_10828);
nand U13941 (N_13941,N_10638,N_11018);
nand U13942 (N_13942,N_10919,N_11393);
and U13943 (N_13943,N_10084,N_11112);
nor U13944 (N_13944,N_11703,N_11490);
and U13945 (N_13945,N_11605,N_10328);
xnor U13946 (N_13946,N_11880,N_10667);
xor U13947 (N_13947,N_10530,N_10320);
nand U13948 (N_13948,N_11552,N_11686);
and U13949 (N_13949,N_11751,N_10633);
or U13950 (N_13950,N_10687,N_11677);
or U13951 (N_13951,N_10288,N_10259);
xnor U13952 (N_13952,N_11555,N_10132);
nor U13953 (N_13953,N_10781,N_10820);
and U13954 (N_13954,N_11360,N_11509);
nand U13955 (N_13955,N_10945,N_10188);
nor U13956 (N_13956,N_11743,N_11048);
nand U13957 (N_13957,N_10698,N_11770);
or U13958 (N_13958,N_10748,N_11911);
or U13959 (N_13959,N_10642,N_11606);
or U13960 (N_13960,N_11499,N_11804);
nor U13961 (N_13961,N_10552,N_10631);
and U13962 (N_13962,N_10761,N_11694);
or U13963 (N_13963,N_10698,N_11038);
nand U13964 (N_13964,N_11468,N_11767);
nor U13965 (N_13965,N_10605,N_10956);
nor U13966 (N_13966,N_10504,N_10362);
xor U13967 (N_13967,N_11703,N_10353);
nor U13968 (N_13968,N_10956,N_10780);
or U13969 (N_13969,N_10999,N_11922);
or U13970 (N_13970,N_10789,N_11218);
nor U13971 (N_13971,N_10886,N_10455);
and U13972 (N_13972,N_10890,N_11406);
nor U13973 (N_13973,N_10064,N_10682);
nor U13974 (N_13974,N_11562,N_10588);
nor U13975 (N_13975,N_10680,N_10960);
nand U13976 (N_13976,N_10765,N_11409);
and U13977 (N_13977,N_10250,N_11058);
xnor U13978 (N_13978,N_10443,N_11008);
nor U13979 (N_13979,N_10427,N_10346);
nor U13980 (N_13980,N_10549,N_11533);
or U13981 (N_13981,N_11777,N_10688);
xor U13982 (N_13982,N_11414,N_11115);
xnor U13983 (N_13983,N_11124,N_10098);
nand U13984 (N_13984,N_11429,N_10990);
xor U13985 (N_13985,N_11144,N_11795);
nand U13986 (N_13986,N_11506,N_10147);
or U13987 (N_13987,N_10057,N_10642);
and U13988 (N_13988,N_10379,N_11005);
and U13989 (N_13989,N_10481,N_11710);
xor U13990 (N_13990,N_11520,N_10440);
and U13991 (N_13991,N_11843,N_11176);
nor U13992 (N_13992,N_10773,N_11560);
nand U13993 (N_13993,N_11566,N_11581);
and U13994 (N_13994,N_11942,N_10523);
or U13995 (N_13995,N_11097,N_11954);
nand U13996 (N_13996,N_11854,N_11988);
or U13997 (N_13997,N_10890,N_10753);
nand U13998 (N_13998,N_10173,N_10889);
or U13999 (N_13999,N_10589,N_11302);
or U14000 (N_14000,N_13955,N_13368);
xnor U14001 (N_14001,N_12557,N_12194);
nand U14002 (N_14002,N_12016,N_12404);
nor U14003 (N_14003,N_13631,N_12343);
nor U14004 (N_14004,N_12221,N_12268);
and U14005 (N_14005,N_12551,N_13171);
or U14006 (N_14006,N_13464,N_12337);
nor U14007 (N_14007,N_12466,N_12601);
and U14008 (N_14008,N_13770,N_13522);
nand U14009 (N_14009,N_13506,N_12274);
or U14010 (N_14010,N_12552,N_12403);
and U14011 (N_14011,N_13192,N_13622);
or U14012 (N_14012,N_12570,N_13503);
nor U14013 (N_14013,N_13287,N_12596);
nand U14014 (N_14014,N_13474,N_12257);
and U14015 (N_14015,N_12514,N_13206);
nor U14016 (N_14016,N_12294,N_13352);
nor U14017 (N_14017,N_13065,N_12774);
xor U14018 (N_14018,N_12058,N_12757);
and U14019 (N_14019,N_13175,N_12032);
and U14020 (N_14020,N_13919,N_12939);
or U14021 (N_14021,N_13433,N_12112);
or U14022 (N_14022,N_13607,N_13008);
nand U14023 (N_14023,N_13187,N_13725);
xnor U14024 (N_14024,N_13609,N_13434);
nand U14025 (N_14025,N_13222,N_13145);
and U14026 (N_14026,N_12180,N_13494);
xor U14027 (N_14027,N_12270,N_12346);
nand U14028 (N_14028,N_12906,N_13298);
or U14029 (N_14029,N_13032,N_13533);
and U14030 (N_14030,N_12796,N_13826);
or U14031 (N_14031,N_13965,N_12679);
xnor U14032 (N_14032,N_13193,N_12487);
xnor U14033 (N_14033,N_13665,N_13751);
and U14034 (N_14034,N_13651,N_13015);
or U14035 (N_14035,N_13742,N_13849);
nand U14036 (N_14036,N_13407,N_12742);
and U14037 (N_14037,N_12879,N_13325);
nor U14038 (N_14038,N_12749,N_13313);
xor U14039 (N_14039,N_12756,N_13796);
or U14040 (N_14040,N_13322,N_12431);
xor U14041 (N_14041,N_12946,N_12116);
or U14042 (N_14042,N_12159,N_12623);
nor U14043 (N_14043,N_12761,N_12536);
xor U14044 (N_14044,N_13667,N_12741);
xnor U14045 (N_14045,N_13271,N_12452);
or U14046 (N_14046,N_12818,N_12957);
or U14047 (N_14047,N_13677,N_12951);
or U14048 (N_14048,N_12018,N_13197);
xor U14049 (N_14049,N_13726,N_12884);
nor U14050 (N_14050,N_13366,N_13549);
and U14051 (N_14051,N_13381,N_13260);
xnor U14052 (N_14052,N_12923,N_12590);
xor U14053 (N_14053,N_12657,N_13165);
xor U14054 (N_14054,N_13164,N_13396);
xor U14055 (N_14055,N_13010,N_12232);
xnor U14056 (N_14056,N_13315,N_13447);
xnor U14057 (N_14057,N_12656,N_12333);
nand U14058 (N_14058,N_12920,N_13612);
xor U14059 (N_14059,N_12791,N_12300);
nand U14060 (N_14060,N_13033,N_12760);
nand U14061 (N_14061,N_13388,N_12430);
xnor U14062 (N_14062,N_13227,N_12241);
xor U14063 (N_14063,N_12661,N_13401);
and U14064 (N_14064,N_13129,N_12190);
or U14065 (N_14065,N_13217,N_13611);
xnor U14066 (N_14066,N_12125,N_13473);
nor U14067 (N_14067,N_13740,N_13870);
and U14068 (N_14068,N_12812,N_12823);
or U14069 (N_14069,N_13654,N_13804);
and U14070 (N_14070,N_12305,N_12523);
or U14071 (N_14071,N_12535,N_12031);
and U14072 (N_14072,N_13463,N_13701);
and U14073 (N_14073,N_13021,N_13053);
or U14074 (N_14074,N_13096,N_12696);
xnor U14075 (N_14075,N_12807,N_12490);
xnor U14076 (N_14076,N_12599,N_13989);
nor U14077 (N_14077,N_13783,N_13162);
nor U14078 (N_14078,N_12352,N_13294);
xnor U14079 (N_14079,N_12720,N_13143);
or U14080 (N_14080,N_12071,N_13185);
and U14081 (N_14081,N_13582,N_13597);
nand U14082 (N_14082,N_12531,N_13158);
and U14083 (N_14083,N_13242,N_12777);
and U14084 (N_14084,N_13137,N_13682);
xnor U14085 (N_14085,N_12817,N_12783);
xnor U14086 (N_14086,N_13801,N_12788);
or U14087 (N_14087,N_12867,N_13468);
and U14088 (N_14088,N_12893,N_12267);
xnor U14089 (N_14089,N_12646,N_13105);
xnor U14090 (N_14090,N_12694,N_12455);
xnor U14091 (N_14091,N_12967,N_13018);
nor U14092 (N_14092,N_13556,N_12844);
or U14093 (N_14093,N_12559,N_13709);
nor U14094 (N_14094,N_13952,N_13089);
xnor U14095 (N_14095,N_12735,N_12958);
and U14096 (N_14096,N_12500,N_12424);
or U14097 (N_14097,N_13357,N_12949);
nor U14098 (N_14098,N_12406,N_12326);
nor U14099 (N_14099,N_12912,N_13283);
nand U14100 (N_14100,N_13146,N_13417);
nor U14101 (N_14101,N_13174,N_13780);
xnor U14102 (N_14102,N_13775,N_12631);
or U14103 (N_14103,N_13684,N_12437);
or U14104 (N_14104,N_12496,N_13560);
nand U14105 (N_14105,N_13948,N_13517);
xnor U14106 (N_14106,N_12229,N_13029);
and U14107 (N_14107,N_13946,N_12492);
nor U14108 (N_14108,N_13276,N_13718);
and U14109 (N_14109,N_13099,N_13215);
nor U14110 (N_14110,N_13571,N_12688);
nor U14111 (N_14111,N_12915,N_13765);
nand U14112 (N_14112,N_13661,N_12191);
nand U14113 (N_14113,N_12815,N_13305);
or U14114 (N_14114,N_13112,N_12594);
nor U14115 (N_14115,N_12717,N_13973);
nor U14116 (N_14116,N_12718,N_12769);
or U14117 (N_14117,N_13257,N_13178);
xnor U14118 (N_14118,N_12779,N_13431);
or U14119 (N_14119,N_13152,N_12520);
or U14120 (N_14120,N_13170,N_12182);
xnor U14121 (N_14121,N_12789,N_13871);
or U14122 (N_14122,N_13130,N_13216);
xor U14123 (N_14123,N_13861,N_13834);
or U14124 (N_14124,N_12135,N_13499);
nand U14125 (N_14125,N_12830,N_12703);
nand U14126 (N_14126,N_12310,N_13452);
xor U14127 (N_14127,N_13251,N_13927);
and U14128 (N_14128,N_13716,N_13127);
nor U14129 (N_14129,N_13617,N_13856);
nand U14130 (N_14130,N_13538,N_12507);
nand U14131 (N_14131,N_12185,N_12321);
nand U14132 (N_14132,N_12090,N_13580);
nand U14133 (N_14133,N_13954,N_12209);
and U14134 (N_14134,N_13062,N_13457);
nand U14135 (N_14135,N_13606,N_13619);
nand U14136 (N_14136,N_12519,N_12651);
or U14137 (N_14137,N_12637,N_13991);
nor U14138 (N_14138,N_12253,N_12615);
and U14139 (N_14139,N_12555,N_13996);
xor U14140 (N_14140,N_12260,N_13759);
nand U14141 (N_14141,N_13031,N_12060);
and U14142 (N_14142,N_13299,N_12499);
nand U14143 (N_14143,N_13256,N_12649);
and U14144 (N_14144,N_13199,N_12065);
nand U14145 (N_14145,N_13916,N_13578);
xor U14146 (N_14146,N_13928,N_12130);
xnor U14147 (N_14147,N_12620,N_13771);
and U14148 (N_14148,N_12087,N_12778);
or U14149 (N_14149,N_13840,N_13832);
xnor U14150 (N_14150,N_12330,N_12117);
or U14151 (N_14151,N_12868,N_13600);
xor U14152 (N_14152,N_12744,N_12020);
xnor U14153 (N_14153,N_12612,N_12436);
nor U14154 (N_14154,N_13354,N_12276);
and U14155 (N_14155,N_13076,N_13043);
xor U14156 (N_14156,N_12273,N_12362);
nor U14157 (N_14157,N_13167,N_12292);
nand U14158 (N_14158,N_13022,N_13639);
xor U14159 (N_14159,N_13882,N_13425);
nand U14160 (N_14160,N_12814,N_12173);
nor U14161 (N_14161,N_12243,N_12894);
xor U14162 (N_14162,N_13747,N_13679);
or U14163 (N_14163,N_13423,N_13243);
and U14164 (N_14164,N_13420,N_13234);
nand U14165 (N_14165,N_12377,N_12279);
xnor U14166 (N_14166,N_12347,N_12317);
and U14167 (N_14167,N_13318,N_12228);
xnor U14168 (N_14168,N_12467,N_13618);
and U14169 (N_14169,N_12149,N_13229);
and U14170 (N_14170,N_13254,N_13488);
nor U14171 (N_14171,N_12632,N_13702);
and U14172 (N_14172,N_12785,N_13527);
and U14173 (N_14173,N_13439,N_12219);
nand U14174 (N_14174,N_12953,N_12203);
nor U14175 (N_14175,N_13255,N_13923);
or U14176 (N_14176,N_13492,N_13157);
nand U14177 (N_14177,N_13109,N_12409);
and U14178 (N_14178,N_13110,N_13190);
nor U14179 (N_14179,N_12441,N_12699);
nor U14180 (N_14180,N_13534,N_13012);
nand U14181 (N_14181,N_13947,N_13083);
or U14182 (N_14182,N_12883,N_12107);
nor U14183 (N_14183,N_12160,N_13913);
nor U14184 (N_14184,N_12944,N_12043);
and U14185 (N_14185,N_12148,N_12617);
or U14186 (N_14186,N_12996,N_12704);
and U14187 (N_14187,N_12419,N_13487);
xor U14188 (N_14188,N_12375,N_12240);
and U14189 (N_14189,N_13876,N_12766);
xor U14190 (N_14190,N_13833,N_12764);
nand U14191 (N_14191,N_13296,N_13554);
or U14192 (N_14192,N_12554,N_13521);
nor U14193 (N_14193,N_13126,N_12534);
xor U14194 (N_14194,N_12813,N_12937);
nand U14195 (N_14195,N_12443,N_13176);
and U14196 (N_14196,N_12484,N_12605);
nand U14197 (N_14197,N_12984,N_13280);
nor U14198 (N_14198,N_13992,N_12763);
or U14199 (N_14199,N_12172,N_12410);
nor U14200 (N_14200,N_12841,N_13017);
nor U14201 (N_14201,N_13787,N_13392);
or U14202 (N_14202,N_13981,N_12610);
xnor U14203 (N_14203,N_12349,N_12449);
nor U14204 (N_14204,N_12296,N_13529);
or U14205 (N_14205,N_13847,N_12085);
nor U14206 (N_14206,N_12390,N_13699);
and U14207 (N_14207,N_12320,N_13743);
or U14208 (N_14208,N_12361,N_13259);
xor U14209 (N_14209,N_13093,N_13986);
or U14210 (N_14210,N_12181,N_13752);
and U14211 (N_14211,N_13685,N_12691);
xor U14212 (N_14212,N_12075,N_12663);
or U14213 (N_14213,N_12524,N_13630);
and U14214 (N_14214,N_13144,N_12510);
or U14215 (N_14215,N_12716,N_13598);
or U14216 (N_14216,N_12607,N_12597);
or U14217 (N_14217,N_13098,N_12099);
nor U14218 (N_14218,N_13442,N_13807);
xnor U14219 (N_14219,N_13041,N_12943);
or U14220 (N_14220,N_12411,N_12952);
and U14221 (N_14221,N_13561,N_12142);
nand U14222 (N_14222,N_13049,N_12629);
nor U14223 (N_14223,N_12114,N_13118);
xnor U14224 (N_14224,N_13084,N_12652);
nand U14225 (N_14225,N_12684,N_12239);
or U14226 (N_14226,N_12722,N_13769);
nand U14227 (N_14227,N_12680,N_12158);
nand U14228 (N_14228,N_13250,N_13841);
and U14229 (N_14229,N_13704,N_12550);
nor U14230 (N_14230,N_12336,N_12976);
xnor U14231 (N_14231,N_13498,N_12754);
and U14232 (N_14232,N_12877,N_12916);
xnor U14233 (N_14233,N_12565,N_12798);
nor U14234 (N_14234,N_13738,N_13642);
or U14235 (N_14235,N_13868,N_12029);
or U14236 (N_14236,N_12972,N_12281);
xor U14237 (N_14237,N_13230,N_12329);
nor U14238 (N_14238,N_12801,N_12236);
xor U14239 (N_14239,N_13774,N_12383);
and U14240 (N_14240,N_13412,N_13646);
nand U14241 (N_14241,N_13269,N_13390);
nand U14242 (N_14242,N_13025,N_12875);
or U14243 (N_14243,N_13450,N_13975);
nor U14244 (N_14244,N_13415,N_12187);
xnor U14245 (N_14245,N_12682,N_13444);
nor U14246 (N_14246,N_12457,N_13231);
and U14247 (N_14247,N_12451,N_13858);
xnor U14248 (N_14248,N_13080,N_12512);
xor U14249 (N_14249,N_12285,N_13339);
xnor U14250 (N_14250,N_13154,N_12829);
xor U14251 (N_14251,N_13111,N_12360);
nand U14252 (N_14252,N_13963,N_13720);
or U14253 (N_14253,N_12028,N_12479);
or U14254 (N_14254,N_13912,N_13785);
or U14255 (N_14255,N_12643,N_13791);
xnor U14256 (N_14256,N_12302,N_12433);
xor U14257 (N_14257,N_12693,N_13343);
nand U14258 (N_14258,N_13375,N_12325);
xor U14259 (N_14259,N_12364,N_12206);
nor U14260 (N_14260,N_12563,N_13161);
nor U14261 (N_14261,N_12578,N_13194);
and U14262 (N_14262,N_13878,N_12393);
or U14263 (N_14263,N_13418,N_13413);
xnor U14264 (N_14264,N_13275,N_12730);
nand U14265 (N_14265,N_13133,N_12262);
nand U14266 (N_14266,N_13956,N_13263);
xnor U14267 (N_14267,N_13356,N_12344);
nand U14268 (N_14268,N_12571,N_12880);
xnor U14269 (N_14269,N_12111,N_12444);
nor U14270 (N_14270,N_12865,N_12928);
nand U14271 (N_14271,N_13393,N_13942);
and U14272 (N_14272,N_12725,N_12978);
xnor U14273 (N_14273,N_12126,N_13933);
and U14274 (N_14274,N_12908,N_13848);
nand U14275 (N_14275,N_13384,N_12439);
nor U14276 (N_14276,N_13301,N_13887);
or U14277 (N_14277,N_13835,N_12989);
nor U14278 (N_14278,N_13753,N_12064);
nor U14279 (N_14279,N_13957,N_13536);
or U14280 (N_14280,N_13812,N_12573);
or U14281 (N_14281,N_13827,N_12385);
xor U14282 (N_14282,N_12583,N_12269);
or U14283 (N_14283,N_13813,N_12354);
and U14284 (N_14284,N_13419,N_12743);
or U14285 (N_14285,N_13967,N_13553);
nor U14286 (N_14286,N_13931,N_12073);
nand U14287 (N_14287,N_13943,N_13545);
nor U14288 (N_14288,N_13671,N_12088);
nor U14289 (N_14289,N_12752,N_12711);
nand U14290 (N_14290,N_12840,N_12141);
xor U14291 (N_14291,N_12794,N_12047);
and U14292 (N_14292,N_13577,N_12380);
or U14293 (N_14293,N_12174,N_12247);
and U14294 (N_14294,N_12220,N_12278);
nand U14295 (N_14295,N_12799,N_13805);
or U14296 (N_14296,N_12904,N_12950);
xor U14297 (N_14297,N_12539,N_13088);
or U14298 (N_14298,N_13344,N_13662);
or U14299 (N_14299,N_12460,N_13095);
nor U14300 (N_14300,N_12113,N_13237);
nor U14301 (N_14301,N_12399,N_12965);
xnor U14302 (N_14302,N_12707,N_13641);
nand U14303 (N_14303,N_13497,N_13938);
or U14304 (N_14304,N_12066,N_12889);
nor U14305 (N_14305,N_13623,N_12739);
or U14306 (N_14306,N_13857,N_13042);
nor U14307 (N_14307,N_13377,N_13903);
nor U14308 (N_14308,N_13106,N_13908);
xor U14309 (N_14309,N_12506,N_12721);
xor U14310 (N_14310,N_12205,N_13458);
and U14311 (N_14311,N_12314,N_12413);
or U14312 (N_14312,N_13048,N_13186);
nor U14313 (N_14313,N_13451,N_13820);
or U14314 (N_14314,N_12245,N_13472);
nor U14315 (N_14315,N_12898,N_13274);
nand U14316 (N_14316,N_12049,N_13934);
nand U14317 (N_14317,N_13372,N_12835);
or U14318 (N_14318,N_13311,N_12922);
xnor U14319 (N_14319,N_13781,N_13120);
and U14320 (N_14320,N_13729,N_12969);
or U14321 (N_14321,N_13940,N_12034);
xnor U14322 (N_14322,N_12025,N_12831);
nand U14323 (N_14323,N_12356,N_13976);
and U14324 (N_14324,N_13360,N_13914);
and U14325 (N_14325,N_12521,N_12471);
nand U14326 (N_14326,N_13614,N_12223);
xor U14327 (N_14327,N_12522,N_12706);
xnor U14328 (N_14328,N_12474,N_12195);
or U14329 (N_14329,N_12529,N_13530);
or U14330 (N_14330,N_12613,N_13002);
xor U14331 (N_14331,N_13063,N_13794);
nor U14332 (N_14332,N_13125,N_13666);
nand U14333 (N_14333,N_13670,N_12138);
nor U14334 (N_14334,N_13309,N_12304);
xnor U14335 (N_14335,N_13636,N_13683);
nor U14336 (N_14336,N_12104,N_13897);
xnor U14337 (N_14337,N_13920,N_13790);
or U14338 (N_14338,N_12638,N_12295);
xor U14339 (N_14339,N_13789,N_13475);
and U14340 (N_14340,N_12945,N_13700);
nand U14341 (N_14341,N_12671,N_12669);
xnor U14342 (N_14342,N_13141,N_12040);
and U14343 (N_14343,N_13226,N_13650);
nor U14344 (N_14344,N_12157,N_12863);
and U14345 (N_14345,N_12048,N_12415);
nor U14346 (N_14346,N_12103,N_12980);
nor U14347 (N_14347,N_13353,N_13427);
nor U14348 (N_14348,N_12005,N_13978);
and U14349 (N_14349,N_13091,N_13964);
xnor U14350 (N_14350,N_13477,N_12780);
and U14351 (N_14351,N_12155,N_13852);
xor U14352 (N_14352,N_12100,N_13588);
or U14353 (N_14353,N_12402,N_12664);
nand U14354 (N_14354,N_13621,N_13410);
nand U14355 (N_14355,N_12373,N_12350);
xor U14356 (N_14356,N_13072,N_12662);
xor U14357 (N_14357,N_12482,N_12477);
nand U14358 (N_14358,N_13668,N_12131);
xnor U14359 (N_14359,N_13816,N_13800);
nor U14360 (N_14360,N_13349,N_12940);
nand U14361 (N_14361,N_13551,N_12151);
or U14362 (N_14362,N_12021,N_13373);
xnor U14363 (N_14363,N_12962,N_12518);
or U14364 (N_14364,N_12227,N_13632);
nor U14365 (N_14365,N_12556,N_12254);
and U14366 (N_14366,N_12004,N_13590);
nand U14367 (N_14367,N_13592,N_12564);
and U14368 (N_14368,N_13486,N_13830);
or U14369 (N_14369,N_12290,N_12608);
nand U14370 (N_14370,N_13505,N_12727);
and U14371 (N_14371,N_12398,N_12003);
nand U14372 (N_14372,N_13335,N_13949);
and U14373 (N_14373,N_13241,N_13262);
or U14374 (N_14374,N_13198,N_13603);
and U14375 (N_14375,N_12332,N_13620);
or U14376 (N_14376,N_12516,N_13988);
xnor U14377 (N_14377,N_13179,N_13050);
and U14378 (N_14378,N_12081,N_12913);
nand U14379 (N_14379,N_12611,N_12987);
and U14380 (N_14380,N_13809,N_12082);
or U14381 (N_14381,N_12307,N_12587);
or U14382 (N_14382,N_13645,N_13404);
nor U14383 (N_14383,N_12309,N_12074);
or U14384 (N_14384,N_13471,N_12386);
xor U14385 (N_14385,N_12572,N_13584);
xor U14386 (N_14386,N_12926,N_13212);
nor U14387 (N_14387,N_12494,N_13663);
or U14388 (N_14388,N_13220,N_12231);
nor U14389 (N_14389,N_12022,N_13994);
nor U14390 (N_14390,N_13524,N_13548);
xor U14391 (N_14391,N_12803,N_13173);
nor U14392 (N_14392,N_13838,N_12050);
xor U14393 (N_14393,N_13839,N_13290);
nand U14394 (N_14394,N_12357,N_13574);
nand U14395 (N_14395,N_13026,N_12491);
or U14396 (N_14396,N_12737,N_12395);
nand U14397 (N_14397,N_12850,N_13634);
nor U14398 (N_14398,N_13884,N_12574);
nor U14399 (N_14399,N_12869,N_13749);
or U14400 (N_14400,N_12878,N_12569);
nand U14401 (N_14401,N_12767,N_12225);
or U14402 (N_14402,N_13310,N_13961);
and U14403 (N_14403,N_13984,N_12170);
nor U14404 (N_14404,N_13828,N_12026);
nor U14405 (N_14405,N_12848,N_12624);
xnor U14406 (N_14406,N_12027,N_12224);
and U14407 (N_14407,N_12150,N_13625);
xnor U14408 (N_14408,N_12019,N_12351);
and U14409 (N_14409,N_13862,N_12024);
and U14410 (N_14410,N_13273,N_12006);
and U14411 (N_14411,N_13055,N_12660);
nor U14412 (N_14412,N_13077,N_12199);
xnor U14413 (N_14413,N_12000,N_12566);
xnor U14414 (N_14414,N_12171,N_12122);
xor U14415 (N_14415,N_13660,N_13124);
nand U14416 (N_14416,N_13900,N_12339);
nor U14417 (N_14417,N_13378,N_13030);
xnor U14418 (N_14418,N_13877,N_13128);
nand U14419 (N_14419,N_12200,N_13090);
xnor U14420 (N_14420,N_12188,N_12975);
or U14421 (N_14421,N_13006,N_12655);
nand U14422 (N_14422,N_13092,N_12715);
xnor U14423 (N_14423,N_13177,N_12348);
or U14424 (N_14424,N_12907,N_12983);
or U14425 (N_14425,N_12667,N_12775);
xnor U14426 (N_14426,N_13071,N_13104);
nor U14427 (N_14427,N_13509,N_12825);
nand U14428 (N_14428,N_12526,N_13402);
nor U14429 (N_14429,N_12327,N_12483);
nor U14430 (N_14430,N_12540,N_12425);
nand U14431 (N_14431,N_12995,N_13842);
or U14432 (N_14432,N_12234,N_13939);
or U14433 (N_14433,N_12502,N_13583);
and U14434 (N_14434,N_12838,N_12265);
nor U14435 (N_14435,N_12054,N_12713);
nand U14436 (N_14436,N_12886,N_13019);
nor U14437 (N_14437,N_12288,N_13034);
nand U14438 (N_14438,N_12790,N_12532);
xor U14439 (N_14439,N_12233,N_12145);
or U14440 (N_14440,N_13168,N_13901);
nand U14441 (N_14441,N_13435,N_12129);
or U14442 (N_14442,N_12137,N_13586);
xor U14443 (N_14443,N_13697,N_12810);
or U14444 (N_14444,N_12947,N_12593);
or U14445 (N_14445,N_12673,N_12579);
or U14446 (N_14446,N_12837,N_12924);
xnor U14447 (N_14447,N_13428,N_13508);
xnor U14448 (N_14448,N_13389,N_12833);
and U14449 (N_14449,N_12396,N_13564);
nor U14450 (N_14450,N_12193,N_12910);
and U14451 (N_14451,N_12475,N_13778);
xnor U14452 (N_14452,N_12297,N_12407);
xnor U14453 (N_14453,N_12678,N_12648);
nand U14454 (N_14454,N_13085,N_13565);
and U14455 (N_14455,N_13204,N_12561);
xnor U14456 (N_14456,N_12497,N_13895);
or U14457 (N_14457,N_12039,N_12079);
or U14458 (N_14458,N_12435,N_13020);
nand U14459 (N_14459,N_13116,N_13723);
or U14460 (N_14460,N_12740,N_13902);
nor U14461 (N_14461,N_12509,N_13532);
nand U14462 (N_14462,N_12977,N_13993);
nand U14463 (N_14463,N_13108,N_13672);
nor U14464 (N_14464,N_13731,N_12069);
nand U14465 (N_14465,N_13664,N_13866);
xor U14466 (N_14466,N_13223,N_13758);
nor U14467 (N_14467,N_12993,N_13694);
nand U14468 (N_14468,N_13755,N_13119);
nor U14469 (N_14469,N_12063,N_12991);
nand U14470 (N_14470,N_12576,N_13734);
nor U14471 (N_14471,N_12672,N_12515);
nand U14472 (N_14472,N_13891,N_12315);
and U14473 (N_14473,N_13485,N_12363);
nor U14474 (N_14474,N_13448,N_13968);
and U14475 (N_14475,N_13886,N_13345);
and U14476 (N_14476,N_12668,N_12609);
nand U14477 (N_14477,N_13653,N_13982);
nor U14478 (N_14478,N_13113,N_12675);
xnor U14479 (N_14479,N_12930,N_13079);
and U14480 (N_14480,N_12936,N_12909);
and U14481 (N_14481,N_13889,N_12824);
xnor U14482 (N_14482,N_13114,N_13024);
nor U14483 (N_14483,N_12714,N_13382);
nor U14484 (N_14484,N_12603,N_13371);
xnor U14485 (N_14485,N_13546,N_12773);
nand U14486 (N_14486,N_12712,N_12885);
and U14487 (N_14487,N_12123,N_13151);
xnor U14488 (N_14488,N_13674,N_13482);
nor U14489 (N_14489,N_13219,N_13297);
or U14490 (N_14490,N_12870,N_13138);
or U14491 (N_14491,N_13935,N_12513);
xnor U14492 (N_14492,N_13558,N_12284);
xnor U14493 (N_14493,N_12486,N_12072);
nand U14494 (N_14494,N_12674,N_12465);
nor U14495 (N_14495,N_13907,N_12676);
and U14496 (N_14496,N_12175,N_12851);
and U14497 (N_14497,N_12218,N_12447);
and U14498 (N_14498,N_12371,N_12263);
nand U14499 (N_14499,N_12731,N_13456);
nand U14500 (N_14500,N_12919,N_13860);
nand U14501 (N_14501,N_13288,N_12708);
xnor U14502 (N_14502,N_13792,N_12979);
nand U14503 (N_14503,N_12323,N_13971);
or U14504 (N_14504,N_13046,N_12164);
nand U14505 (N_14505,N_12345,N_12115);
and U14506 (N_14506,N_12046,N_12316);
nor U14507 (N_14507,N_12689,N_12765);
and U14508 (N_14508,N_12666,N_13330);
nor U14509 (N_14509,N_13515,N_13676);
nand U14510 (N_14510,N_12547,N_13040);
and U14511 (N_14511,N_13693,N_13817);
xor U14512 (N_14512,N_13806,N_13652);
nor U14513 (N_14513,N_13896,N_12313);
or U14514 (N_14514,N_13921,N_13380);
or U14515 (N_14515,N_13459,N_12728);
nand U14516 (N_14516,N_12960,N_13863);
xor U14517 (N_14517,N_12729,N_12165);
or U14518 (N_14518,N_12598,N_13510);
nand U14519 (N_14519,N_13075,N_12562);
and U14520 (N_14520,N_13972,N_13385);
nor U14521 (N_14521,N_13054,N_12461);
nand U14522 (N_14522,N_12068,N_12308);
and U14523 (N_14523,N_13869,N_13047);
or U14524 (N_14524,N_12770,N_13710);
xnor U14525 (N_14525,N_12982,N_12143);
nand U14526 (N_14526,N_12681,N_13678);
nand U14527 (N_14527,N_12719,N_13240);
nor U14528 (N_14528,N_12319,N_13189);
nor U14529 (N_14529,N_13235,N_13541);
nand U14530 (N_14530,N_13784,N_13762);
nand U14531 (N_14531,N_12035,N_13763);
or U14532 (N_14532,N_12198,N_13730);
or U14533 (N_14533,N_13979,N_13926);
or U14534 (N_14534,N_12834,N_13067);
xnor U14535 (N_14535,N_13818,N_13005);
nor U14536 (N_14536,N_12002,N_12934);
nand U14537 (N_14537,N_12935,N_13815);
nor U14538 (N_14538,N_12341,N_13566);
nor U14539 (N_14539,N_12378,N_12146);
nor U14540 (N_14540,N_13074,N_13713);
nand U14541 (N_14541,N_12110,N_13793);
or U14542 (N_14542,N_13898,N_12804);
or U14543 (N_14543,N_12811,N_13542);
or U14544 (N_14544,N_13628,N_12768);
nand U14545 (N_14545,N_13593,N_13248);
nand U14546 (N_14546,N_13070,N_12528);
xnor U14547 (N_14547,N_13616,N_12981);
nand U14548 (N_14548,N_13911,N_13312);
xnor U14549 (N_14549,N_12762,N_13058);
nand U14550 (N_14550,N_13405,N_12809);
nor U14551 (N_14551,N_12543,N_12136);
and U14552 (N_14552,N_12581,N_13708);
nand U14553 (N_14553,N_12903,N_12828);
xor U14554 (N_14554,N_13478,N_13873);
or U14555 (N_14555,N_13421,N_13342);
nor U14556 (N_14556,N_13557,N_13350);
and U14557 (N_14557,N_12955,N_13233);
nand U14558 (N_14558,N_12845,N_13656);
and U14559 (N_14559,N_13881,N_13408);
nand U14560 (N_14560,N_12686,N_12537);
or U14561 (N_14561,N_13319,N_12010);
or U14562 (N_14562,N_13727,N_12214);
or U14563 (N_14563,N_12335,N_12095);
and U14564 (N_14564,N_12097,N_12450);
and U14565 (N_14565,N_13056,N_13461);
xnor U14566 (N_14566,N_12902,N_12871);
nor U14567 (N_14567,N_12261,N_13998);
nor U14568 (N_14568,N_12128,N_12405);
nand U14569 (N_14569,N_13003,N_13314);
nand U14570 (N_14570,N_12856,N_13648);
and U14571 (N_14571,N_13466,N_13136);
nand U14572 (N_14572,N_12849,N_12575);
nand U14573 (N_14573,N_12213,N_12445);
xor U14574 (N_14574,N_12478,N_12489);
nand U14575 (N_14575,N_13153,N_12698);
xor U14576 (N_14576,N_13027,N_13224);
xor U14577 (N_14577,N_13277,N_13864);
nor U14578 (N_14578,N_12446,N_13329);
nand U14579 (N_14579,N_12772,N_12179);
xnor U14580 (N_14580,N_13822,N_13414);
xor U14581 (N_14581,N_12751,N_13121);
and U14582 (N_14582,N_13983,N_12710);
and U14583 (N_14583,N_12517,N_13493);
nand U14584 (N_14584,N_12334,N_12299);
and U14585 (N_14585,N_12560,N_12106);
or U14586 (N_14586,N_13200,N_13845);
xor U14587 (N_14587,N_12985,N_13962);
xnor U14588 (N_14588,N_13507,N_12259);
and U14589 (N_14589,N_12086,N_12248);
xnor U14590 (N_14590,N_13232,N_12968);
or U14591 (N_14591,N_12897,N_12282);
and U14592 (N_14592,N_12062,N_12933);
nand U14593 (N_14593,N_13358,N_13712);
or U14594 (N_14594,N_12009,N_12567);
or U14595 (N_14595,N_12634,N_13953);
and U14596 (N_14596,N_12258,N_12359);
nand U14597 (N_14597,N_12498,N_12367);
and U14598 (N_14598,N_13985,N_13245);
xnor U14599 (N_14599,N_12291,N_12639);
or U14600 (N_14600,N_12255,N_13406);
xnor U14601 (N_14601,N_13196,N_13591);
nand U14602 (N_14602,N_13722,N_13865);
or U14603 (N_14603,N_12015,N_12644);
and U14604 (N_14604,N_13773,N_13181);
or U14605 (N_14605,N_12230,N_13811);
xor U14606 (N_14606,N_12287,N_13159);
and U14607 (N_14607,N_13516,N_13374);
nor U14608 (N_14608,N_13995,N_13244);
and U14609 (N_14609,N_13585,N_13550);
nand U14610 (N_14610,N_12216,N_13706);
nand U14611 (N_14611,N_12217,N_13221);
xor U14612 (N_14612,N_12932,N_12827);
nor U14613 (N_14613,N_12853,N_12453);
nand U14614 (N_14614,N_12108,N_12249);
xor U14615 (N_14615,N_12215,N_13009);
and U14616 (N_14616,N_12917,N_13635);
and U14617 (N_14617,N_13843,N_12585);
xnor U14618 (N_14618,N_12670,N_12508);
and U14619 (N_14619,N_13037,N_13737);
xnor U14620 (N_14620,N_12476,N_12012);
and U14621 (N_14621,N_12311,N_13205);
nor U14622 (N_14622,N_12961,N_13540);
nand U14623 (N_14623,N_12745,N_13253);
or U14624 (N_14624,N_12931,N_12876);
nand U14625 (N_14625,N_13432,N_13411);
or U14626 (N_14626,N_12429,N_12376);
nand U14627 (N_14627,N_12368,N_12918);
nand U14628 (N_14628,N_13086,N_13362);
or U14629 (N_14629,N_13629,N_12527);
xor U14630 (N_14630,N_13559,N_13370);
and U14631 (N_14631,N_13707,N_13552);
nand U14632 (N_14632,N_12511,N_13361);
xnor U14633 (N_14633,N_12914,N_12842);
nor U14634 (N_14634,N_12872,N_12041);
or U14635 (N_14635,N_12732,N_13531);
or U14636 (N_14636,N_12102,N_12238);
xnor U14637 (N_14637,N_13915,N_12473);
and U14638 (N_14638,N_12161,N_13686);
xnor U14639 (N_14639,N_12692,N_12588);
xnor U14640 (N_14640,N_13579,N_13337);
and U14641 (N_14641,N_13930,N_12816);
or U14642 (N_14642,N_13799,N_12503);
nor U14643 (N_14643,N_12797,N_13182);
or U14644 (N_14644,N_13123,N_13465);
or U14645 (N_14645,N_12784,N_12895);
nor U14646 (N_14646,N_12901,N_13397);
and U14647 (N_14647,N_12469,N_12966);
or U14648 (N_14648,N_12548,N_13844);
nand U14649 (N_14649,N_13334,N_12887);
and U14650 (N_14650,N_12423,N_12013);
xnor U14651 (N_14651,N_12211,N_12250);
and U14652 (N_14652,N_13140,N_13107);
nor U14653 (N_14653,N_12454,N_12726);
or U14654 (N_14654,N_13733,N_13596);
or U14655 (N_14655,N_12162,N_12382);
xor U14656 (N_14656,N_13673,N_13469);
or U14657 (N_14657,N_13581,N_12630);
and U14658 (N_14658,N_13798,N_13036);
nor U14659 (N_14659,N_12891,N_13454);
or U14660 (N_14660,N_12558,N_13750);
nor U14661 (N_14661,N_12379,N_12747);
or U14662 (N_14662,N_12992,N_12485);
nand U14663 (N_14663,N_13480,N_13746);
or U14664 (N_14664,N_12998,N_13476);
or U14665 (N_14665,N_13172,N_13724);
xor U14666 (N_14666,N_12802,N_13195);
xor U14667 (N_14667,N_12192,N_13906);
or U14668 (N_14668,N_12076,N_12324);
nand U14669 (N_14669,N_13101,N_13997);
nand U14670 (N_14670,N_12963,N_12459);
or U14671 (N_14671,N_13208,N_12625);
or U14672 (N_14672,N_13655,N_13855);
nor U14673 (N_14673,N_12045,N_12826);
and U14674 (N_14674,N_13004,N_13819);
nor U14675 (N_14675,N_13249,N_13265);
xnor U14676 (N_14676,N_13624,N_12470);
xor U14677 (N_14677,N_12189,N_12549);
xnor U14678 (N_14678,N_12890,N_13387);
nand U14679 (N_14679,N_13644,N_13073);
xor U14680 (N_14680,N_12252,N_12272);
or U14681 (N_14681,N_12408,N_12251);
xor U14682 (N_14682,N_12458,N_12283);
xor U14683 (N_14683,N_13867,N_12821);
and U14684 (N_14684,N_13929,N_13258);
or U14685 (N_14685,N_13284,N_13155);
or U14686 (N_14686,N_13403,N_13761);
nor U14687 (N_14687,N_12805,N_12036);
or U14688 (N_14688,N_12568,N_12776);
xor U14689 (N_14689,N_13810,N_13803);
and U14690 (N_14690,N_13608,N_12621);
and U14691 (N_14691,N_12759,N_12892);
xor U14692 (N_14692,N_13543,N_12734);
or U14693 (N_14693,N_13714,N_12077);
and U14694 (N_14694,N_13537,N_13264);
nand U14695 (N_14695,N_13735,N_13400);
nand U14696 (N_14696,N_13490,N_13148);
xor U14697 (N_14697,N_13376,N_12636);
or U14698 (N_14698,N_12888,N_12653);
nand U14699 (N_14699,N_13449,N_13149);
and U14700 (N_14700,N_12859,N_13150);
and U14701 (N_14701,N_12700,N_13122);
nand U14702 (N_14702,N_13484,N_13739);
and U14703 (N_14703,N_13899,N_12633);
nand U14704 (N_14704,N_12822,N_13637);
or U14705 (N_14705,N_12580,N_12806);
xor U14706 (N_14706,N_12008,N_13306);
and U14707 (N_14707,N_12748,N_12096);
and U14708 (N_14708,N_13980,N_12365);
or U14709 (N_14709,N_13332,N_12169);
xnor U14710 (N_14710,N_12542,N_12011);
xor U14711 (N_14711,N_12723,N_13535);
nand U14712 (N_14712,N_12153,N_12861);
nand U14713 (N_14713,N_12685,N_13757);
nor U14714 (N_14714,N_12586,N_12140);
nor U14715 (N_14715,N_12353,N_12246);
and U14716 (N_14716,N_13333,N_13568);
or U14717 (N_14717,N_13977,N_13501);
nand U14718 (N_14718,N_13691,N_13268);
xnor U14719 (N_14719,N_13604,N_13688);
nor U14720 (N_14720,N_13051,N_12954);
and U14721 (N_14721,N_13489,N_13643);
xnor U14722 (N_14722,N_13990,N_12462);
and U14723 (N_14723,N_12001,N_12858);
and U14724 (N_14724,N_12614,N_12124);
and U14725 (N_14725,N_13057,N_13282);
and U14726 (N_14726,N_13359,N_13772);
nor U14727 (N_14727,N_12440,N_13028);
nor U14728 (N_14728,N_12226,N_12427);
and U14729 (N_14729,N_13348,N_12340);
nor U14730 (N_14730,N_13379,N_13436);
xor U14731 (N_14731,N_13768,N_13117);
and U14732 (N_14732,N_12204,N_13894);
xor U14733 (N_14733,N_13872,N_13504);
nand U14734 (N_14734,N_12592,N_12659);
or U14735 (N_14735,N_12481,N_12546);
and U14736 (N_14736,N_13572,N_13821);
xnor U14737 (N_14737,N_13575,N_12168);
or U14738 (N_14738,N_13347,N_13690);
or U14739 (N_14739,N_13917,N_12293);
nand U14740 (N_14740,N_12280,N_13695);
nand U14741 (N_14741,N_12618,N_12121);
nor U14742 (N_14742,N_12650,N_13880);
nand U14743 (N_14743,N_13853,N_13328);
nand U14744 (N_14744,N_13038,N_13627);
or U14745 (N_14745,N_12070,N_12120);
nor U14746 (N_14746,N_13814,N_13308);
nand U14747 (N_14747,N_13918,N_13307);
nor U14748 (N_14748,N_13286,N_13295);
nand U14749 (N_14749,N_13369,N_12970);
and U14750 (N_14750,N_13941,N_12038);
xnor U14751 (N_14751,N_12078,N_12622);
or U14752 (N_14752,N_13570,N_13767);
nand U14753 (N_14753,N_12464,N_13681);
xnor U14754 (N_14754,N_12755,N_12298);
nand U14755 (N_14755,N_13859,N_12438);
nand U14756 (N_14756,N_13601,N_13569);
xor U14757 (N_14757,N_12683,N_12210);
or U14758 (N_14758,N_12388,N_13649);
nand U14759 (N_14759,N_13786,N_12852);
nand U14760 (N_14760,N_13239,N_12616);
and U14761 (N_14761,N_12595,N_13539);
or U14762 (N_14762,N_12358,N_13825);
xnor U14763 (N_14763,N_12400,N_12758);
nor U14764 (N_14764,N_12056,N_12619);
nand U14765 (N_14765,N_13659,N_12178);
or U14766 (N_14766,N_12750,N_13610);
nand U14767 (N_14767,N_13013,N_13395);
and U14768 (N_14768,N_13455,N_13958);
or U14769 (N_14769,N_13851,N_13443);
or U14770 (N_14770,N_12468,N_13365);
or U14771 (N_14771,N_13936,N_13555);
and U14772 (N_14772,N_13831,N_12640);
or U14773 (N_14773,N_13698,N_13278);
and U14774 (N_14774,N_13201,N_13850);
nand U14775 (N_14775,N_12974,N_13987);
and U14776 (N_14776,N_13715,N_12421);
and U14777 (N_14777,N_12053,N_12927);
nor U14778 (N_14778,N_12084,N_12956);
and U14779 (N_14779,N_12196,N_13512);
or U14780 (N_14780,N_12235,N_13669);
xnor U14781 (N_14781,N_12873,N_13745);
nand U14782 (N_14782,N_13760,N_12422);
nor U14783 (N_14783,N_12301,N_13836);
nor U14784 (N_14784,N_12836,N_13061);
nor U14785 (N_14785,N_12338,N_13909);
and U14786 (N_14786,N_12808,N_13777);
or U14787 (N_14787,N_12051,N_13523);
or U14788 (N_14788,N_12899,N_13399);
or U14789 (N_14789,N_12677,N_12426);
xnor U14790 (N_14790,N_12387,N_13802);
xor U14791 (N_14791,N_13326,N_13426);
or U14792 (N_14792,N_12820,N_13910);
nor U14793 (N_14793,N_13782,N_13082);
nor U14794 (N_14794,N_12533,N_13429);
and U14795 (N_14795,N_13445,N_12911);
nand U14796 (N_14796,N_13479,N_13689);
nand U14797 (N_14797,N_13135,N_12746);
nor U14798 (N_14798,N_13594,N_12819);
nor U14799 (N_14799,N_12237,N_13272);
xor U14800 (N_14800,N_13068,N_12442);
or U14801 (N_14801,N_12042,N_12017);
xnor U14802 (N_14802,N_12553,N_12303);
or U14803 (N_14803,N_13317,N_12266);
xnor U14804 (N_14804,N_13658,N_12434);
and U14805 (N_14805,N_13925,N_12654);
or U14806 (N_14806,N_12342,N_12971);
nand U14807 (N_14807,N_13892,N_12089);
or U14808 (N_14808,N_13211,N_12154);
and U14809 (N_14809,N_12709,N_13721);
nand U14810 (N_14810,N_13779,N_12584);
and U14811 (N_14811,N_13795,N_13131);
nand U14812 (N_14812,N_13970,N_12147);
nor U14813 (N_14813,N_12736,N_13969);
nand U14814 (N_14814,N_12782,N_12033);
nand U14815 (N_14815,N_12900,N_12418);
or U14816 (N_14816,N_12994,N_13302);
xnor U14817 (N_14817,N_12530,N_13705);
xnor U14818 (N_14818,N_13097,N_12545);
or U14819 (N_14819,N_13924,N_12176);
and U14820 (N_14820,N_13383,N_13363);
nand U14821 (N_14821,N_13711,N_13441);
xor U14822 (N_14822,N_12793,N_12312);
or U14823 (N_14823,N_13209,N_13132);
nor U14824 (N_14824,N_13576,N_12105);
and U14825 (N_14825,N_12589,N_12052);
nand U14826 (N_14826,N_12416,N_12602);
xnor U14827 (N_14827,N_13094,N_12420);
nor U14828 (N_14828,N_13776,N_12412);
or U14829 (N_14829,N_12094,N_13696);
or U14830 (N_14830,N_12697,N_13511);
and U14831 (N_14831,N_13069,N_13267);
nand U14832 (N_14832,N_13142,N_13470);
xnor U14833 (N_14833,N_13160,N_13950);
nand U14834 (N_14834,N_13945,N_13687);
nand U14835 (N_14835,N_13453,N_12059);
and U14836 (N_14836,N_12397,N_12092);
nand U14837 (N_14837,N_13460,N_13797);
and U14838 (N_14838,N_13589,N_13246);
nor U14839 (N_14839,N_13331,N_13045);
and U14840 (N_14840,N_12183,N_12771);
xor U14841 (N_14841,N_13854,N_13039);
and U14842 (N_14842,N_13270,N_13188);
nor U14843 (N_14843,N_13437,N_12480);
nor U14844 (N_14844,N_12463,N_12392);
and U14845 (N_14845,N_12695,N_13102);
and U14846 (N_14846,N_12591,N_12244);
nor U14847 (N_14847,N_12495,N_13398);
xnor U14848 (N_14848,N_12472,N_13210);
and U14849 (N_14849,N_13218,N_13766);
xnor U14850 (N_14850,N_13595,N_12306);
nor U14851 (N_14851,N_12134,N_12389);
and U14852 (N_14852,N_12642,N_12862);
nor U14853 (N_14853,N_12525,N_13520);
nand U14854 (N_14854,N_13180,N_13893);
and U14855 (N_14855,N_13846,N_13207);
nor U14856 (N_14856,N_13213,N_13281);
nor U14857 (N_14857,N_13587,N_13647);
or U14858 (N_14858,N_13156,N_12055);
and U14859 (N_14859,N_13885,N_13340);
and U14860 (N_14860,N_13544,N_13922);
nand U14861 (N_14861,N_12448,N_13657);
or U14862 (N_14862,N_13424,N_12197);
nand U14863 (N_14863,N_12504,N_12786);
or U14864 (N_14864,N_13719,N_13748);
nor U14865 (N_14865,N_13321,N_12119);
or U14866 (N_14866,N_13364,N_13338);
or U14867 (N_14867,N_12456,N_13367);
and U14868 (N_14868,N_13823,N_13147);
nand U14869 (N_14869,N_13717,N_12690);
xnor U14870 (N_14870,N_12037,N_12921);
nor U14871 (N_14871,N_13500,N_12057);
nand U14872 (N_14872,N_13764,N_12384);
and U14873 (N_14873,N_12792,N_13134);
xor U14874 (N_14874,N_13440,N_12641);
xnor U14875 (N_14875,N_13346,N_13905);
nand U14876 (N_14876,N_13615,N_12874);
xor U14877 (N_14877,N_13052,N_12144);
xnor U14878 (N_14878,N_13951,N_12401);
nor U14879 (N_14879,N_13890,N_12847);
nor U14880 (N_14880,N_12030,N_12372);
and U14881 (N_14881,N_12860,N_13491);
xnor U14882 (N_14882,N_12800,N_13513);
nand U14883 (N_14883,N_13808,N_12882);
xnor U14884 (N_14884,N_12414,N_13303);
nor U14885 (N_14885,N_13023,N_13238);
nor U14886 (N_14886,N_12538,N_13279);
and U14887 (N_14887,N_13044,N_12381);
xor U14888 (N_14888,N_13496,N_13202);
nand U14889 (N_14889,N_13300,N_13519);
or U14890 (N_14890,N_13087,N_12275);
xor U14891 (N_14891,N_13289,N_13115);
or U14892 (N_14892,N_12541,N_13355);
xnor U14893 (N_14893,N_13100,N_12929);
and U14894 (N_14894,N_13732,N_13324);
xnor U14895 (N_14895,N_12207,N_12881);
and U14896 (N_14896,N_12369,N_12864);
xnor U14897 (N_14897,N_12289,N_12101);
xor U14898 (N_14898,N_13495,N_13183);
xnor U14899 (N_14899,N_13547,N_12355);
nand U14900 (N_14900,N_12156,N_12091);
and U14901 (N_14901,N_12986,N_13514);
or U14902 (N_14902,N_12839,N_13394);
nor U14903 (N_14903,N_13829,N_12264);
or U14904 (N_14904,N_13974,N_12132);
or U14905 (N_14905,N_13875,N_12118);
nand U14906 (N_14906,N_12705,N_12394);
xor U14907 (N_14907,N_13203,N_13035);
nor U14908 (N_14908,N_13386,N_13736);
and U14909 (N_14909,N_12999,N_13103);
or U14910 (N_14910,N_13320,N_13247);
and U14911 (N_14911,N_13351,N_13788);
or U14912 (N_14912,N_13059,N_13261);
nand U14913 (N_14913,N_12061,N_12328);
nor U14914 (N_14914,N_12493,N_12753);
or U14915 (N_14915,N_13562,N_13567);
xor U14916 (N_14916,N_12186,N_12152);
or U14917 (N_14917,N_12577,N_12687);
nand U14918 (N_14918,N_12604,N_12832);
nor U14919 (N_14919,N_13169,N_12488);
nor U14920 (N_14920,N_12014,N_12212);
xor U14921 (N_14921,N_12787,N_12391);
nor U14922 (N_14922,N_12582,N_13573);
nand U14923 (N_14923,N_12896,N_12139);
nor U14924 (N_14924,N_13703,N_12428);
or U14925 (N_14925,N_13446,N_13191);
nor U14926 (N_14926,N_12432,N_13741);
xor U14927 (N_14927,N_13754,N_13166);
and U14928 (N_14928,N_13064,N_13430);
nand U14929 (N_14929,N_12166,N_13563);
and U14930 (N_14930,N_13692,N_12866);
or U14931 (N_14931,N_12080,N_12322);
xor U14932 (N_14932,N_13291,N_12959);
xnor U14933 (N_14933,N_12208,N_12271);
nand U14934 (N_14934,N_12948,N_13824);
and U14935 (N_14935,N_13837,N_13640);
or U14936 (N_14936,N_13323,N_13081);
or U14937 (N_14937,N_12318,N_13066);
nor U14938 (N_14938,N_13888,N_13225);
or U14939 (N_14939,N_13883,N_12997);
or U14940 (N_14940,N_13944,N_12702);
or U14941 (N_14941,N_13001,N_12202);
and U14942 (N_14942,N_13744,N_13728);
xnor U14943 (N_14943,N_12505,N_13438);
and U14944 (N_14944,N_12857,N_12942);
nand U14945 (N_14945,N_13602,N_13675);
nor U14946 (N_14946,N_13462,N_12647);
or U14947 (N_14947,N_13904,N_13007);
nor U14948 (N_14948,N_12701,N_12658);
xor U14949 (N_14949,N_13626,N_12854);
and U14950 (N_14950,N_13638,N_12738);
nor U14951 (N_14951,N_13422,N_13932);
and U14952 (N_14952,N_13292,N_13000);
xor U14953 (N_14953,N_12627,N_12133);
nor U14954 (N_14954,N_12370,N_13014);
xor U14955 (N_14955,N_12795,N_12044);
nand U14956 (N_14956,N_13481,N_12184);
nor U14957 (N_14957,N_12083,N_13316);
xor U14958 (N_14958,N_12626,N_12938);
nand U14959 (N_14959,N_12964,N_13016);
and U14960 (N_14960,N_13266,N_13228);
nand U14961 (N_14961,N_12606,N_13304);
nand U14962 (N_14962,N_12023,N_12628);
and U14963 (N_14963,N_13341,N_13966);
and U14964 (N_14964,N_12925,N_12331);
nor U14965 (N_14965,N_13613,N_13060);
or U14966 (N_14966,N_13252,N_12098);
nor U14967 (N_14967,N_13518,N_12665);
or U14968 (N_14968,N_12222,N_13528);
and U14969 (N_14969,N_13525,N_12109);
and U14970 (N_14970,N_13680,N_13336);
or U14971 (N_14971,N_12277,N_12366);
nand U14972 (N_14972,N_12733,N_12544);
xor U14973 (N_14973,N_13467,N_13139);
or U14974 (N_14974,N_12781,N_12990);
nor U14975 (N_14975,N_12007,N_12256);
nand U14976 (N_14976,N_12724,N_12973);
nand U14977 (N_14977,N_12067,N_12127);
nor U14978 (N_14978,N_13163,N_13960);
nand U14979 (N_14979,N_13285,N_12846);
or U14980 (N_14980,N_13502,N_13959);
xor U14981 (N_14981,N_12843,N_12635);
and U14982 (N_14982,N_12177,N_13184);
nor U14983 (N_14983,N_12242,N_12093);
xor U14984 (N_14984,N_13874,N_13999);
nor U14985 (N_14985,N_12374,N_13214);
xnor U14986 (N_14986,N_13327,N_12645);
xnor U14987 (N_14987,N_12201,N_13011);
and U14988 (N_14988,N_13391,N_13599);
xnor U14989 (N_14989,N_13409,N_13483);
or U14990 (N_14990,N_12600,N_12855);
xor U14991 (N_14991,N_12905,N_13879);
nand U14992 (N_14992,N_13526,N_12988);
xnor U14993 (N_14993,N_12167,N_12163);
xor U14994 (N_14994,N_12417,N_12941);
or U14995 (N_14995,N_13937,N_13236);
and U14996 (N_14996,N_13078,N_13293);
nor U14997 (N_14997,N_13633,N_12286);
nor U14998 (N_14998,N_13605,N_13416);
nor U14999 (N_14999,N_12501,N_13756);
nor U15000 (N_15000,N_13873,N_12698);
nand U15001 (N_15001,N_13696,N_12901);
xnor U15002 (N_15002,N_13931,N_12588);
or U15003 (N_15003,N_12571,N_13771);
or U15004 (N_15004,N_12677,N_13886);
or U15005 (N_15005,N_12424,N_12847);
nor U15006 (N_15006,N_13244,N_13087);
and U15007 (N_15007,N_13374,N_13409);
xor U15008 (N_15008,N_13037,N_12080);
nand U15009 (N_15009,N_13508,N_12135);
nor U15010 (N_15010,N_12943,N_12444);
xnor U15011 (N_15011,N_12792,N_12819);
xnor U15012 (N_15012,N_12473,N_13960);
and U15013 (N_15013,N_13159,N_12190);
nor U15014 (N_15014,N_13214,N_13662);
or U15015 (N_15015,N_13411,N_13616);
and U15016 (N_15016,N_12889,N_13957);
nand U15017 (N_15017,N_13041,N_13479);
or U15018 (N_15018,N_12739,N_13962);
and U15019 (N_15019,N_13109,N_12412);
or U15020 (N_15020,N_12650,N_12843);
or U15021 (N_15021,N_13839,N_12604);
nor U15022 (N_15022,N_12694,N_13483);
or U15023 (N_15023,N_12809,N_12228);
xnor U15024 (N_15024,N_12300,N_12120);
nor U15025 (N_15025,N_12959,N_12845);
nand U15026 (N_15026,N_12746,N_12529);
nand U15027 (N_15027,N_12452,N_13145);
and U15028 (N_15028,N_13610,N_12211);
nand U15029 (N_15029,N_12161,N_12801);
nor U15030 (N_15030,N_13966,N_13096);
or U15031 (N_15031,N_12217,N_12506);
or U15032 (N_15032,N_13737,N_13465);
xor U15033 (N_15033,N_12741,N_13646);
and U15034 (N_15034,N_13186,N_13236);
xor U15035 (N_15035,N_12461,N_12428);
xor U15036 (N_15036,N_13333,N_12495);
or U15037 (N_15037,N_13269,N_12716);
nor U15038 (N_15038,N_13741,N_13190);
nor U15039 (N_15039,N_12900,N_13176);
nor U15040 (N_15040,N_13993,N_13644);
nand U15041 (N_15041,N_12091,N_13996);
or U15042 (N_15042,N_12125,N_13582);
and U15043 (N_15043,N_12245,N_12042);
or U15044 (N_15044,N_13434,N_12626);
nand U15045 (N_15045,N_13564,N_13917);
nand U15046 (N_15046,N_13589,N_12671);
xor U15047 (N_15047,N_13294,N_13707);
xnor U15048 (N_15048,N_13667,N_13374);
nand U15049 (N_15049,N_12985,N_12265);
and U15050 (N_15050,N_12091,N_12351);
xnor U15051 (N_15051,N_12677,N_13180);
or U15052 (N_15052,N_12774,N_13827);
and U15053 (N_15053,N_12818,N_13460);
and U15054 (N_15054,N_12324,N_13774);
xnor U15055 (N_15055,N_13259,N_13330);
xnor U15056 (N_15056,N_13350,N_12115);
and U15057 (N_15057,N_12190,N_13469);
xor U15058 (N_15058,N_12402,N_13499);
or U15059 (N_15059,N_12767,N_13487);
nand U15060 (N_15060,N_12852,N_12748);
nand U15061 (N_15061,N_13808,N_13685);
xnor U15062 (N_15062,N_13443,N_12882);
or U15063 (N_15063,N_12972,N_13145);
nand U15064 (N_15064,N_12631,N_13489);
and U15065 (N_15065,N_12816,N_13325);
xor U15066 (N_15066,N_12374,N_12572);
nor U15067 (N_15067,N_13680,N_12262);
nand U15068 (N_15068,N_13463,N_12025);
nor U15069 (N_15069,N_13669,N_12720);
nor U15070 (N_15070,N_13032,N_13211);
and U15071 (N_15071,N_12006,N_12713);
nor U15072 (N_15072,N_12378,N_13667);
nand U15073 (N_15073,N_13756,N_12532);
and U15074 (N_15074,N_13500,N_12848);
and U15075 (N_15075,N_12869,N_12903);
xnor U15076 (N_15076,N_12859,N_12051);
or U15077 (N_15077,N_12610,N_13825);
xor U15078 (N_15078,N_13264,N_13011);
or U15079 (N_15079,N_13238,N_13909);
nor U15080 (N_15080,N_13646,N_12598);
or U15081 (N_15081,N_13187,N_12194);
nand U15082 (N_15082,N_13325,N_12897);
or U15083 (N_15083,N_13716,N_13859);
and U15084 (N_15084,N_13300,N_13582);
nand U15085 (N_15085,N_13199,N_12937);
and U15086 (N_15086,N_12663,N_12593);
nor U15087 (N_15087,N_12189,N_13629);
and U15088 (N_15088,N_12749,N_13870);
nor U15089 (N_15089,N_13570,N_12290);
xnor U15090 (N_15090,N_12023,N_12678);
xor U15091 (N_15091,N_13457,N_13413);
xor U15092 (N_15092,N_12193,N_12376);
nand U15093 (N_15093,N_12586,N_12728);
and U15094 (N_15094,N_13479,N_12596);
xnor U15095 (N_15095,N_12855,N_13970);
and U15096 (N_15096,N_12958,N_13154);
nand U15097 (N_15097,N_12189,N_13571);
or U15098 (N_15098,N_12901,N_13770);
nor U15099 (N_15099,N_13065,N_13594);
nor U15100 (N_15100,N_13467,N_12636);
or U15101 (N_15101,N_13351,N_12811);
nor U15102 (N_15102,N_12929,N_13507);
and U15103 (N_15103,N_13636,N_12712);
xnor U15104 (N_15104,N_13177,N_12279);
or U15105 (N_15105,N_13396,N_13174);
nor U15106 (N_15106,N_13606,N_12880);
and U15107 (N_15107,N_13843,N_12285);
or U15108 (N_15108,N_12462,N_13543);
xnor U15109 (N_15109,N_12961,N_13282);
and U15110 (N_15110,N_12281,N_13965);
nor U15111 (N_15111,N_13428,N_13163);
nor U15112 (N_15112,N_12075,N_13534);
xnor U15113 (N_15113,N_12243,N_13993);
nor U15114 (N_15114,N_13280,N_13480);
nor U15115 (N_15115,N_12033,N_13663);
or U15116 (N_15116,N_13754,N_12918);
or U15117 (N_15117,N_13553,N_12106);
nor U15118 (N_15118,N_12859,N_12578);
and U15119 (N_15119,N_12257,N_13413);
and U15120 (N_15120,N_13405,N_12090);
or U15121 (N_15121,N_12778,N_12668);
nand U15122 (N_15122,N_13652,N_13765);
xor U15123 (N_15123,N_12291,N_12960);
nor U15124 (N_15124,N_12044,N_12733);
and U15125 (N_15125,N_13210,N_12830);
and U15126 (N_15126,N_12032,N_13738);
nand U15127 (N_15127,N_12797,N_13695);
and U15128 (N_15128,N_13567,N_13085);
nand U15129 (N_15129,N_12977,N_13339);
nand U15130 (N_15130,N_12653,N_13579);
and U15131 (N_15131,N_13582,N_12236);
nor U15132 (N_15132,N_12271,N_12861);
nand U15133 (N_15133,N_12528,N_13023);
or U15134 (N_15134,N_13477,N_12232);
nor U15135 (N_15135,N_13754,N_13327);
nor U15136 (N_15136,N_12226,N_13842);
nand U15137 (N_15137,N_13715,N_12506);
nor U15138 (N_15138,N_12790,N_12353);
xor U15139 (N_15139,N_12623,N_13241);
or U15140 (N_15140,N_13727,N_13989);
xnor U15141 (N_15141,N_12272,N_12005);
nand U15142 (N_15142,N_12360,N_12854);
or U15143 (N_15143,N_12874,N_12791);
or U15144 (N_15144,N_13299,N_12224);
xor U15145 (N_15145,N_13756,N_13517);
or U15146 (N_15146,N_13474,N_12136);
nor U15147 (N_15147,N_13153,N_13667);
or U15148 (N_15148,N_13692,N_13790);
xor U15149 (N_15149,N_12103,N_12659);
xor U15150 (N_15150,N_13383,N_13812);
nor U15151 (N_15151,N_13304,N_13265);
and U15152 (N_15152,N_13284,N_13087);
nor U15153 (N_15153,N_13692,N_12433);
xor U15154 (N_15154,N_12346,N_12144);
nand U15155 (N_15155,N_12035,N_12865);
nand U15156 (N_15156,N_13471,N_12514);
nor U15157 (N_15157,N_12908,N_12710);
xor U15158 (N_15158,N_12479,N_12717);
xnor U15159 (N_15159,N_12226,N_12969);
nand U15160 (N_15160,N_13417,N_12232);
nand U15161 (N_15161,N_12785,N_12427);
and U15162 (N_15162,N_12203,N_13362);
xor U15163 (N_15163,N_13677,N_12949);
and U15164 (N_15164,N_12179,N_12982);
xnor U15165 (N_15165,N_12813,N_12182);
nand U15166 (N_15166,N_12116,N_13755);
or U15167 (N_15167,N_12443,N_13809);
nand U15168 (N_15168,N_13982,N_12027);
nor U15169 (N_15169,N_13505,N_12309);
and U15170 (N_15170,N_13022,N_13121);
xnor U15171 (N_15171,N_13786,N_12783);
and U15172 (N_15172,N_12852,N_12902);
or U15173 (N_15173,N_13730,N_12794);
and U15174 (N_15174,N_12367,N_12988);
or U15175 (N_15175,N_12376,N_12289);
xor U15176 (N_15176,N_12962,N_13452);
xnor U15177 (N_15177,N_13491,N_12822);
xor U15178 (N_15178,N_13678,N_12861);
xor U15179 (N_15179,N_12327,N_12653);
xnor U15180 (N_15180,N_13802,N_13061);
nor U15181 (N_15181,N_12464,N_13817);
nor U15182 (N_15182,N_13469,N_13921);
nor U15183 (N_15183,N_12056,N_13789);
or U15184 (N_15184,N_13142,N_13662);
or U15185 (N_15185,N_12078,N_13918);
nor U15186 (N_15186,N_12273,N_13091);
nor U15187 (N_15187,N_12731,N_13383);
nand U15188 (N_15188,N_12405,N_12828);
or U15189 (N_15189,N_13394,N_13650);
xnor U15190 (N_15190,N_12354,N_12753);
nand U15191 (N_15191,N_13336,N_13562);
xor U15192 (N_15192,N_12032,N_13753);
or U15193 (N_15193,N_12625,N_12624);
and U15194 (N_15194,N_12663,N_13233);
or U15195 (N_15195,N_13773,N_13688);
xor U15196 (N_15196,N_12901,N_12876);
and U15197 (N_15197,N_12532,N_12291);
and U15198 (N_15198,N_12909,N_13148);
and U15199 (N_15199,N_12641,N_13740);
and U15200 (N_15200,N_12119,N_12382);
and U15201 (N_15201,N_13308,N_13619);
and U15202 (N_15202,N_13505,N_13131);
or U15203 (N_15203,N_13770,N_12621);
and U15204 (N_15204,N_13587,N_13055);
nand U15205 (N_15205,N_13156,N_12083);
or U15206 (N_15206,N_12096,N_13078);
and U15207 (N_15207,N_13613,N_13317);
nand U15208 (N_15208,N_13248,N_13974);
or U15209 (N_15209,N_12933,N_13519);
and U15210 (N_15210,N_12274,N_13700);
and U15211 (N_15211,N_12474,N_13174);
nand U15212 (N_15212,N_12172,N_13845);
xnor U15213 (N_15213,N_12681,N_13554);
xnor U15214 (N_15214,N_12748,N_12514);
xnor U15215 (N_15215,N_12639,N_13203);
and U15216 (N_15216,N_12917,N_13278);
nand U15217 (N_15217,N_13925,N_12817);
or U15218 (N_15218,N_12834,N_12102);
or U15219 (N_15219,N_12061,N_13906);
nor U15220 (N_15220,N_13389,N_13683);
or U15221 (N_15221,N_13138,N_12869);
or U15222 (N_15222,N_13047,N_13503);
nand U15223 (N_15223,N_12898,N_13954);
xnor U15224 (N_15224,N_12457,N_13215);
and U15225 (N_15225,N_13981,N_13379);
nor U15226 (N_15226,N_12999,N_13436);
nor U15227 (N_15227,N_13307,N_12822);
nand U15228 (N_15228,N_12136,N_13747);
xor U15229 (N_15229,N_12679,N_12099);
nor U15230 (N_15230,N_12797,N_12009);
or U15231 (N_15231,N_13379,N_12530);
nand U15232 (N_15232,N_13651,N_13409);
xor U15233 (N_15233,N_13333,N_13967);
nand U15234 (N_15234,N_12551,N_12154);
and U15235 (N_15235,N_13525,N_13520);
and U15236 (N_15236,N_13033,N_13926);
and U15237 (N_15237,N_13504,N_13562);
nand U15238 (N_15238,N_12788,N_13421);
or U15239 (N_15239,N_13392,N_12320);
or U15240 (N_15240,N_12608,N_12578);
and U15241 (N_15241,N_12420,N_13256);
and U15242 (N_15242,N_13697,N_12673);
xnor U15243 (N_15243,N_12602,N_12316);
xor U15244 (N_15244,N_12607,N_12218);
xor U15245 (N_15245,N_12090,N_12149);
or U15246 (N_15246,N_13159,N_13988);
nand U15247 (N_15247,N_12916,N_13382);
xor U15248 (N_15248,N_13518,N_13807);
or U15249 (N_15249,N_12613,N_12223);
xnor U15250 (N_15250,N_13471,N_12737);
nor U15251 (N_15251,N_13470,N_12419);
and U15252 (N_15252,N_13404,N_13467);
xnor U15253 (N_15253,N_12962,N_13870);
nor U15254 (N_15254,N_13388,N_12078);
nor U15255 (N_15255,N_12457,N_12831);
or U15256 (N_15256,N_13805,N_13244);
or U15257 (N_15257,N_12104,N_12548);
nor U15258 (N_15258,N_13710,N_13504);
and U15259 (N_15259,N_13878,N_13105);
xnor U15260 (N_15260,N_13230,N_12680);
xor U15261 (N_15261,N_13481,N_13566);
nand U15262 (N_15262,N_12762,N_13018);
and U15263 (N_15263,N_12973,N_12398);
and U15264 (N_15264,N_12833,N_12222);
xor U15265 (N_15265,N_13419,N_13575);
xnor U15266 (N_15266,N_12147,N_13059);
nor U15267 (N_15267,N_12468,N_12121);
xor U15268 (N_15268,N_13458,N_13761);
xor U15269 (N_15269,N_13509,N_12331);
xnor U15270 (N_15270,N_13346,N_13249);
nand U15271 (N_15271,N_13432,N_13399);
xor U15272 (N_15272,N_12010,N_12991);
xor U15273 (N_15273,N_13914,N_12165);
and U15274 (N_15274,N_12866,N_12719);
nor U15275 (N_15275,N_13568,N_12119);
xor U15276 (N_15276,N_12841,N_12213);
nor U15277 (N_15277,N_13694,N_12983);
xnor U15278 (N_15278,N_13413,N_12287);
nand U15279 (N_15279,N_12871,N_13762);
nand U15280 (N_15280,N_12463,N_13948);
xnor U15281 (N_15281,N_12640,N_13539);
nor U15282 (N_15282,N_12549,N_13642);
or U15283 (N_15283,N_13144,N_13468);
xnor U15284 (N_15284,N_13998,N_13760);
and U15285 (N_15285,N_12773,N_12134);
xnor U15286 (N_15286,N_13348,N_13471);
nor U15287 (N_15287,N_13856,N_12057);
xor U15288 (N_15288,N_12522,N_13699);
nor U15289 (N_15289,N_12588,N_12078);
nand U15290 (N_15290,N_13098,N_13690);
nand U15291 (N_15291,N_12825,N_12572);
and U15292 (N_15292,N_13017,N_12675);
nand U15293 (N_15293,N_12335,N_13184);
or U15294 (N_15294,N_13288,N_13965);
and U15295 (N_15295,N_12106,N_13722);
or U15296 (N_15296,N_13009,N_12610);
nor U15297 (N_15297,N_13032,N_13777);
and U15298 (N_15298,N_13682,N_12290);
xor U15299 (N_15299,N_12616,N_12112);
nor U15300 (N_15300,N_13250,N_12724);
nand U15301 (N_15301,N_13261,N_12071);
and U15302 (N_15302,N_13382,N_13782);
and U15303 (N_15303,N_12735,N_12449);
nor U15304 (N_15304,N_12135,N_12509);
xor U15305 (N_15305,N_13489,N_13768);
and U15306 (N_15306,N_12956,N_13978);
nand U15307 (N_15307,N_12744,N_12364);
nor U15308 (N_15308,N_13494,N_13291);
nand U15309 (N_15309,N_13499,N_12162);
xor U15310 (N_15310,N_12257,N_12450);
nand U15311 (N_15311,N_13787,N_13999);
or U15312 (N_15312,N_13351,N_13015);
nand U15313 (N_15313,N_12746,N_12174);
and U15314 (N_15314,N_13682,N_12937);
and U15315 (N_15315,N_12667,N_13613);
and U15316 (N_15316,N_12172,N_13710);
nand U15317 (N_15317,N_13121,N_13094);
nand U15318 (N_15318,N_12614,N_12205);
nor U15319 (N_15319,N_12263,N_12219);
xnor U15320 (N_15320,N_12061,N_12508);
nand U15321 (N_15321,N_13562,N_13003);
xnor U15322 (N_15322,N_13957,N_13004);
or U15323 (N_15323,N_13710,N_13387);
or U15324 (N_15324,N_12290,N_13365);
nand U15325 (N_15325,N_13830,N_12194);
or U15326 (N_15326,N_12139,N_12122);
and U15327 (N_15327,N_13395,N_13001);
and U15328 (N_15328,N_12470,N_13585);
nand U15329 (N_15329,N_12475,N_13174);
or U15330 (N_15330,N_13348,N_12713);
and U15331 (N_15331,N_13982,N_13299);
nand U15332 (N_15332,N_13598,N_12053);
nor U15333 (N_15333,N_12215,N_13929);
nor U15334 (N_15334,N_12651,N_12293);
nor U15335 (N_15335,N_13714,N_13809);
xor U15336 (N_15336,N_13396,N_13686);
nor U15337 (N_15337,N_12537,N_12190);
nand U15338 (N_15338,N_12815,N_12391);
nand U15339 (N_15339,N_13995,N_12297);
or U15340 (N_15340,N_12072,N_12502);
nand U15341 (N_15341,N_12905,N_13814);
nor U15342 (N_15342,N_13255,N_12165);
or U15343 (N_15343,N_13212,N_13026);
and U15344 (N_15344,N_12323,N_13348);
xor U15345 (N_15345,N_13908,N_13201);
nor U15346 (N_15346,N_12315,N_13847);
nand U15347 (N_15347,N_13477,N_13864);
xnor U15348 (N_15348,N_13162,N_12111);
nor U15349 (N_15349,N_13008,N_12182);
and U15350 (N_15350,N_12165,N_12032);
or U15351 (N_15351,N_12358,N_13807);
nor U15352 (N_15352,N_13013,N_13523);
or U15353 (N_15353,N_13876,N_12675);
nand U15354 (N_15354,N_13390,N_13033);
nand U15355 (N_15355,N_12682,N_13546);
or U15356 (N_15356,N_12630,N_12280);
xnor U15357 (N_15357,N_12190,N_12111);
nor U15358 (N_15358,N_12583,N_12769);
nand U15359 (N_15359,N_13271,N_13510);
xor U15360 (N_15360,N_13361,N_13119);
or U15361 (N_15361,N_13562,N_12651);
nand U15362 (N_15362,N_13685,N_12806);
nand U15363 (N_15363,N_13968,N_12197);
nor U15364 (N_15364,N_13058,N_12740);
and U15365 (N_15365,N_12493,N_12527);
nand U15366 (N_15366,N_13805,N_13775);
or U15367 (N_15367,N_12552,N_12571);
nor U15368 (N_15368,N_13060,N_13337);
nor U15369 (N_15369,N_12635,N_13693);
nor U15370 (N_15370,N_13246,N_13295);
nor U15371 (N_15371,N_13323,N_12059);
and U15372 (N_15372,N_12932,N_13203);
nand U15373 (N_15373,N_12416,N_13384);
nor U15374 (N_15374,N_13694,N_13181);
and U15375 (N_15375,N_13736,N_12377);
nand U15376 (N_15376,N_12231,N_13234);
nor U15377 (N_15377,N_12876,N_13604);
or U15378 (N_15378,N_12807,N_12858);
and U15379 (N_15379,N_13443,N_12726);
and U15380 (N_15380,N_12575,N_12399);
or U15381 (N_15381,N_13814,N_13888);
and U15382 (N_15382,N_13891,N_12121);
nor U15383 (N_15383,N_12780,N_13928);
or U15384 (N_15384,N_13694,N_12067);
or U15385 (N_15385,N_13325,N_12570);
or U15386 (N_15386,N_12024,N_13176);
and U15387 (N_15387,N_13965,N_12644);
and U15388 (N_15388,N_13738,N_13452);
nand U15389 (N_15389,N_12128,N_13138);
xnor U15390 (N_15390,N_12023,N_12592);
and U15391 (N_15391,N_12335,N_12905);
and U15392 (N_15392,N_12735,N_13416);
and U15393 (N_15393,N_13810,N_13619);
and U15394 (N_15394,N_12384,N_12397);
nor U15395 (N_15395,N_12880,N_12081);
and U15396 (N_15396,N_12691,N_13086);
xnor U15397 (N_15397,N_12726,N_12589);
nand U15398 (N_15398,N_12754,N_13284);
nor U15399 (N_15399,N_13891,N_13462);
nor U15400 (N_15400,N_12168,N_12786);
xnor U15401 (N_15401,N_12926,N_13738);
or U15402 (N_15402,N_12794,N_13066);
and U15403 (N_15403,N_13928,N_12544);
and U15404 (N_15404,N_13723,N_12248);
nor U15405 (N_15405,N_12415,N_13305);
nor U15406 (N_15406,N_12952,N_12822);
nand U15407 (N_15407,N_12768,N_13601);
xnor U15408 (N_15408,N_12066,N_12036);
and U15409 (N_15409,N_12628,N_12780);
nor U15410 (N_15410,N_13909,N_13303);
or U15411 (N_15411,N_13009,N_12928);
nor U15412 (N_15412,N_12137,N_13529);
and U15413 (N_15413,N_13218,N_13648);
or U15414 (N_15414,N_12269,N_12319);
and U15415 (N_15415,N_13546,N_13879);
or U15416 (N_15416,N_13989,N_12514);
nor U15417 (N_15417,N_12464,N_12951);
and U15418 (N_15418,N_12151,N_12355);
and U15419 (N_15419,N_13763,N_12229);
nor U15420 (N_15420,N_12602,N_13925);
nor U15421 (N_15421,N_13150,N_13411);
xor U15422 (N_15422,N_13604,N_13731);
or U15423 (N_15423,N_13185,N_13840);
or U15424 (N_15424,N_12432,N_13197);
nor U15425 (N_15425,N_13856,N_12711);
or U15426 (N_15426,N_13970,N_12979);
nand U15427 (N_15427,N_13288,N_13876);
nand U15428 (N_15428,N_13464,N_13430);
or U15429 (N_15429,N_13885,N_12325);
nor U15430 (N_15430,N_12767,N_13481);
and U15431 (N_15431,N_12513,N_13644);
or U15432 (N_15432,N_13582,N_12404);
and U15433 (N_15433,N_12582,N_12923);
nand U15434 (N_15434,N_13751,N_12828);
or U15435 (N_15435,N_12230,N_12876);
or U15436 (N_15436,N_12156,N_12417);
nor U15437 (N_15437,N_12401,N_13788);
nand U15438 (N_15438,N_13663,N_13561);
or U15439 (N_15439,N_12682,N_13753);
xor U15440 (N_15440,N_12098,N_13513);
nor U15441 (N_15441,N_12250,N_12946);
and U15442 (N_15442,N_13845,N_12005);
nand U15443 (N_15443,N_12132,N_12875);
nor U15444 (N_15444,N_13708,N_12963);
and U15445 (N_15445,N_13869,N_13106);
or U15446 (N_15446,N_13251,N_12442);
nand U15447 (N_15447,N_12482,N_12465);
or U15448 (N_15448,N_12928,N_13904);
xor U15449 (N_15449,N_12579,N_13343);
or U15450 (N_15450,N_12655,N_13628);
nand U15451 (N_15451,N_13713,N_12125);
or U15452 (N_15452,N_13402,N_13515);
xor U15453 (N_15453,N_12182,N_12539);
or U15454 (N_15454,N_12285,N_13690);
nor U15455 (N_15455,N_13321,N_13357);
nand U15456 (N_15456,N_13703,N_13364);
xnor U15457 (N_15457,N_13600,N_13742);
xor U15458 (N_15458,N_13183,N_12747);
xor U15459 (N_15459,N_13606,N_12213);
nand U15460 (N_15460,N_12357,N_12705);
xor U15461 (N_15461,N_12468,N_13724);
xor U15462 (N_15462,N_12271,N_13067);
nand U15463 (N_15463,N_12804,N_13458);
nand U15464 (N_15464,N_13721,N_12396);
xor U15465 (N_15465,N_12083,N_12847);
nand U15466 (N_15466,N_12896,N_12503);
nor U15467 (N_15467,N_13961,N_12709);
and U15468 (N_15468,N_13246,N_12011);
nand U15469 (N_15469,N_13009,N_12606);
or U15470 (N_15470,N_13766,N_12445);
xnor U15471 (N_15471,N_12853,N_13288);
and U15472 (N_15472,N_13747,N_13082);
nand U15473 (N_15473,N_12978,N_12991);
nand U15474 (N_15474,N_12069,N_12515);
nand U15475 (N_15475,N_13009,N_13066);
nand U15476 (N_15476,N_12601,N_13212);
xnor U15477 (N_15477,N_12283,N_12516);
nor U15478 (N_15478,N_13661,N_13503);
xor U15479 (N_15479,N_13873,N_12808);
nand U15480 (N_15480,N_13418,N_13097);
xnor U15481 (N_15481,N_13401,N_12399);
xnor U15482 (N_15482,N_12309,N_13991);
or U15483 (N_15483,N_12901,N_12085);
xnor U15484 (N_15484,N_12819,N_12492);
or U15485 (N_15485,N_13120,N_12106);
nand U15486 (N_15486,N_13835,N_13828);
xnor U15487 (N_15487,N_13068,N_13679);
xor U15488 (N_15488,N_13668,N_12878);
xnor U15489 (N_15489,N_13660,N_12089);
nor U15490 (N_15490,N_13132,N_12666);
or U15491 (N_15491,N_13144,N_12413);
nand U15492 (N_15492,N_12683,N_12030);
nand U15493 (N_15493,N_12486,N_12813);
or U15494 (N_15494,N_12662,N_12980);
nand U15495 (N_15495,N_12240,N_13335);
nor U15496 (N_15496,N_13359,N_12379);
nand U15497 (N_15497,N_13368,N_12240);
or U15498 (N_15498,N_12140,N_13056);
and U15499 (N_15499,N_12640,N_13247);
xor U15500 (N_15500,N_12370,N_12263);
xnor U15501 (N_15501,N_13587,N_12505);
or U15502 (N_15502,N_13426,N_13399);
or U15503 (N_15503,N_12903,N_12732);
nor U15504 (N_15504,N_12864,N_12117);
xor U15505 (N_15505,N_12111,N_12965);
xnor U15506 (N_15506,N_12607,N_12426);
nor U15507 (N_15507,N_12514,N_13153);
or U15508 (N_15508,N_13083,N_12885);
and U15509 (N_15509,N_12077,N_13383);
xor U15510 (N_15510,N_12945,N_13164);
xnor U15511 (N_15511,N_13442,N_12471);
or U15512 (N_15512,N_13513,N_13888);
nand U15513 (N_15513,N_12503,N_12980);
nand U15514 (N_15514,N_13228,N_13261);
or U15515 (N_15515,N_13016,N_12934);
xnor U15516 (N_15516,N_12858,N_13308);
xor U15517 (N_15517,N_12494,N_12633);
and U15518 (N_15518,N_13007,N_13998);
xor U15519 (N_15519,N_13307,N_13790);
or U15520 (N_15520,N_13976,N_12937);
and U15521 (N_15521,N_12341,N_12793);
nor U15522 (N_15522,N_13332,N_13401);
or U15523 (N_15523,N_12555,N_13727);
nor U15524 (N_15524,N_12458,N_13866);
or U15525 (N_15525,N_12928,N_13243);
nor U15526 (N_15526,N_13637,N_12824);
and U15527 (N_15527,N_12644,N_12158);
or U15528 (N_15528,N_13144,N_12307);
and U15529 (N_15529,N_13854,N_13843);
xnor U15530 (N_15530,N_13311,N_13432);
nor U15531 (N_15531,N_13084,N_13379);
nor U15532 (N_15532,N_13447,N_12679);
and U15533 (N_15533,N_12150,N_12499);
xnor U15534 (N_15534,N_13721,N_12179);
or U15535 (N_15535,N_12102,N_13864);
nor U15536 (N_15536,N_13936,N_13443);
and U15537 (N_15537,N_12837,N_12455);
and U15538 (N_15538,N_12051,N_12225);
nand U15539 (N_15539,N_12686,N_13534);
or U15540 (N_15540,N_13719,N_12036);
nand U15541 (N_15541,N_13268,N_13906);
or U15542 (N_15542,N_12015,N_13795);
xnor U15543 (N_15543,N_12236,N_12050);
xor U15544 (N_15544,N_13100,N_13810);
nor U15545 (N_15545,N_13640,N_13570);
or U15546 (N_15546,N_13718,N_13974);
xor U15547 (N_15547,N_13657,N_13852);
nor U15548 (N_15548,N_12728,N_12145);
xnor U15549 (N_15549,N_13688,N_13795);
nor U15550 (N_15550,N_12129,N_13181);
or U15551 (N_15551,N_12536,N_13963);
or U15552 (N_15552,N_12473,N_13987);
nand U15553 (N_15553,N_12404,N_12536);
and U15554 (N_15554,N_13901,N_13765);
and U15555 (N_15555,N_12288,N_12788);
or U15556 (N_15556,N_12025,N_12668);
and U15557 (N_15557,N_12241,N_12909);
or U15558 (N_15558,N_12584,N_13750);
nand U15559 (N_15559,N_13187,N_13470);
or U15560 (N_15560,N_13567,N_12281);
nor U15561 (N_15561,N_13058,N_12353);
nor U15562 (N_15562,N_13189,N_12657);
nand U15563 (N_15563,N_13123,N_12971);
nor U15564 (N_15564,N_13118,N_12977);
or U15565 (N_15565,N_13303,N_13328);
and U15566 (N_15566,N_12673,N_13350);
nor U15567 (N_15567,N_12124,N_12333);
nor U15568 (N_15568,N_13363,N_12441);
xnor U15569 (N_15569,N_13936,N_13563);
nor U15570 (N_15570,N_13113,N_12737);
xnor U15571 (N_15571,N_13085,N_12353);
or U15572 (N_15572,N_12138,N_13263);
nand U15573 (N_15573,N_12171,N_12466);
or U15574 (N_15574,N_12710,N_13310);
and U15575 (N_15575,N_12797,N_12771);
or U15576 (N_15576,N_13023,N_13530);
or U15577 (N_15577,N_13011,N_12255);
and U15578 (N_15578,N_13185,N_13564);
xnor U15579 (N_15579,N_12988,N_12537);
xor U15580 (N_15580,N_12605,N_12451);
nor U15581 (N_15581,N_13417,N_12727);
and U15582 (N_15582,N_12846,N_12860);
xor U15583 (N_15583,N_12646,N_12163);
nor U15584 (N_15584,N_13040,N_13375);
xor U15585 (N_15585,N_13398,N_12417);
nand U15586 (N_15586,N_12786,N_13658);
or U15587 (N_15587,N_12820,N_13737);
or U15588 (N_15588,N_13250,N_13452);
nor U15589 (N_15589,N_12880,N_12005);
nor U15590 (N_15590,N_13183,N_13492);
xnor U15591 (N_15591,N_13852,N_12031);
xor U15592 (N_15592,N_13848,N_13852);
xor U15593 (N_15593,N_13916,N_12873);
nor U15594 (N_15594,N_13699,N_12070);
nor U15595 (N_15595,N_12954,N_13141);
nand U15596 (N_15596,N_13263,N_13861);
or U15597 (N_15597,N_13774,N_12829);
and U15598 (N_15598,N_12860,N_12424);
and U15599 (N_15599,N_12926,N_12703);
or U15600 (N_15600,N_12139,N_13076);
nor U15601 (N_15601,N_12414,N_13810);
and U15602 (N_15602,N_12116,N_13823);
nand U15603 (N_15603,N_13780,N_12994);
nor U15604 (N_15604,N_13514,N_13099);
and U15605 (N_15605,N_12833,N_12868);
nor U15606 (N_15606,N_13602,N_13235);
xor U15607 (N_15607,N_13464,N_12988);
nor U15608 (N_15608,N_13000,N_12773);
or U15609 (N_15609,N_13760,N_13280);
nand U15610 (N_15610,N_12462,N_12710);
and U15611 (N_15611,N_13580,N_12944);
and U15612 (N_15612,N_12583,N_12121);
nor U15613 (N_15613,N_13891,N_13550);
and U15614 (N_15614,N_13084,N_13225);
nand U15615 (N_15615,N_12352,N_12178);
or U15616 (N_15616,N_12062,N_13710);
or U15617 (N_15617,N_12312,N_13235);
or U15618 (N_15618,N_12136,N_12739);
xnor U15619 (N_15619,N_12718,N_12075);
or U15620 (N_15620,N_13242,N_12273);
and U15621 (N_15621,N_12485,N_13607);
xor U15622 (N_15622,N_13680,N_12770);
or U15623 (N_15623,N_13001,N_13393);
nor U15624 (N_15624,N_13633,N_13701);
nor U15625 (N_15625,N_12576,N_12966);
nor U15626 (N_15626,N_13672,N_13298);
nor U15627 (N_15627,N_13669,N_12735);
or U15628 (N_15628,N_13297,N_13067);
or U15629 (N_15629,N_12703,N_13062);
xor U15630 (N_15630,N_13091,N_12758);
nor U15631 (N_15631,N_12323,N_12481);
xor U15632 (N_15632,N_13140,N_13384);
nor U15633 (N_15633,N_13859,N_12850);
xnor U15634 (N_15634,N_12429,N_13795);
or U15635 (N_15635,N_12302,N_13697);
or U15636 (N_15636,N_12377,N_13107);
or U15637 (N_15637,N_12440,N_12173);
nand U15638 (N_15638,N_13553,N_12530);
nor U15639 (N_15639,N_13617,N_13007);
or U15640 (N_15640,N_12281,N_13837);
nor U15641 (N_15641,N_12542,N_12932);
and U15642 (N_15642,N_12826,N_13180);
and U15643 (N_15643,N_13322,N_13416);
nand U15644 (N_15644,N_13133,N_12278);
nand U15645 (N_15645,N_13895,N_12398);
xnor U15646 (N_15646,N_12141,N_12907);
xnor U15647 (N_15647,N_13247,N_12598);
nand U15648 (N_15648,N_12450,N_13041);
or U15649 (N_15649,N_13346,N_12347);
or U15650 (N_15650,N_12398,N_13908);
xor U15651 (N_15651,N_13099,N_12567);
nor U15652 (N_15652,N_13129,N_12113);
or U15653 (N_15653,N_12125,N_13812);
and U15654 (N_15654,N_12891,N_12237);
and U15655 (N_15655,N_13579,N_13608);
and U15656 (N_15656,N_13615,N_13773);
or U15657 (N_15657,N_12912,N_12456);
and U15658 (N_15658,N_13920,N_13324);
nor U15659 (N_15659,N_12551,N_12228);
nand U15660 (N_15660,N_12102,N_13625);
or U15661 (N_15661,N_13445,N_12755);
nor U15662 (N_15662,N_13602,N_12526);
nand U15663 (N_15663,N_13808,N_13423);
nor U15664 (N_15664,N_13057,N_13508);
nand U15665 (N_15665,N_12774,N_13707);
and U15666 (N_15666,N_13873,N_12926);
xor U15667 (N_15667,N_13559,N_13043);
nor U15668 (N_15668,N_13192,N_13684);
and U15669 (N_15669,N_12777,N_13896);
and U15670 (N_15670,N_13872,N_13668);
nor U15671 (N_15671,N_12169,N_13134);
and U15672 (N_15672,N_13130,N_12659);
nand U15673 (N_15673,N_12305,N_13464);
or U15674 (N_15674,N_13043,N_13124);
nand U15675 (N_15675,N_12148,N_13329);
nor U15676 (N_15676,N_12884,N_13343);
and U15677 (N_15677,N_13647,N_12481);
xnor U15678 (N_15678,N_13979,N_13486);
and U15679 (N_15679,N_12467,N_12205);
or U15680 (N_15680,N_13134,N_12494);
nand U15681 (N_15681,N_12142,N_12223);
nand U15682 (N_15682,N_12282,N_12901);
nand U15683 (N_15683,N_13542,N_13549);
or U15684 (N_15684,N_12809,N_12526);
nand U15685 (N_15685,N_13003,N_12737);
nor U15686 (N_15686,N_13285,N_13229);
and U15687 (N_15687,N_12673,N_12316);
xnor U15688 (N_15688,N_13351,N_12189);
nor U15689 (N_15689,N_12743,N_13566);
or U15690 (N_15690,N_12293,N_12565);
nand U15691 (N_15691,N_13193,N_12102);
nand U15692 (N_15692,N_13808,N_12674);
or U15693 (N_15693,N_13241,N_13126);
or U15694 (N_15694,N_12669,N_12501);
xor U15695 (N_15695,N_13093,N_13257);
or U15696 (N_15696,N_13623,N_13725);
nand U15697 (N_15697,N_12819,N_12301);
nor U15698 (N_15698,N_12367,N_13774);
nor U15699 (N_15699,N_13958,N_13656);
xnor U15700 (N_15700,N_12132,N_13074);
or U15701 (N_15701,N_13027,N_13221);
and U15702 (N_15702,N_13684,N_12575);
xnor U15703 (N_15703,N_13495,N_12199);
and U15704 (N_15704,N_13231,N_13269);
nor U15705 (N_15705,N_12971,N_13269);
nand U15706 (N_15706,N_13967,N_12579);
or U15707 (N_15707,N_12476,N_13159);
or U15708 (N_15708,N_13779,N_13353);
nor U15709 (N_15709,N_12476,N_13887);
or U15710 (N_15710,N_13943,N_13293);
xnor U15711 (N_15711,N_12575,N_13939);
nand U15712 (N_15712,N_12424,N_12813);
nand U15713 (N_15713,N_12077,N_13923);
and U15714 (N_15714,N_13904,N_13760);
nor U15715 (N_15715,N_12686,N_13997);
nand U15716 (N_15716,N_13102,N_12324);
nor U15717 (N_15717,N_12289,N_13764);
nor U15718 (N_15718,N_13384,N_12966);
and U15719 (N_15719,N_12234,N_13393);
or U15720 (N_15720,N_12589,N_12526);
xnor U15721 (N_15721,N_12380,N_12261);
and U15722 (N_15722,N_12366,N_12421);
nor U15723 (N_15723,N_13887,N_13982);
xor U15724 (N_15724,N_12090,N_12977);
or U15725 (N_15725,N_13650,N_12840);
nor U15726 (N_15726,N_12874,N_13846);
nand U15727 (N_15727,N_12581,N_12449);
and U15728 (N_15728,N_13864,N_13829);
or U15729 (N_15729,N_13345,N_13475);
or U15730 (N_15730,N_12871,N_13506);
nor U15731 (N_15731,N_12465,N_12521);
or U15732 (N_15732,N_12687,N_13474);
xor U15733 (N_15733,N_12507,N_12526);
and U15734 (N_15734,N_13709,N_12476);
and U15735 (N_15735,N_12379,N_13435);
xnor U15736 (N_15736,N_12415,N_13050);
nand U15737 (N_15737,N_13487,N_12962);
and U15738 (N_15738,N_13633,N_12008);
nor U15739 (N_15739,N_13134,N_13689);
nor U15740 (N_15740,N_12116,N_12231);
and U15741 (N_15741,N_12439,N_13708);
nor U15742 (N_15742,N_12471,N_12284);
nor U15743 (N_15743,N_12199,N_13836);
nor U15744 (N_15744,N_13798,N_12519);
xnor U15745 (N_15745,N_12962,N_13124);
nand U15746 (N_15746,N_13672,N_12577);
xor U15747 (N_15747,N_12452,N_13025);
nor U15748 (N_15748,N_13147,N_12737);
or U15749 (N_15749,N_13645,N_12939);
nor U15750 (N_15750,N_12031,N_13587);
or U15751 (N_15751,N_12017,N_12931);
nor U15752 (N_15752,N_13239,N_12628);
and U15753 (N_15753,N_13375,N_13058);
nor U15754 (N_15754,N_12234,N_12011);
nand U15755 (N_15755,N_13943,N_12212);
or U15756 (N_15756,N_12478,N_13261);
xnor U15757 (N_15757,N_13858,N_13155);
or U15758 (N_15758,N_13007,N_13911);
xnor U15759 (N_15759,N_13621,N_13603);
nand U15760 (N_15760,N_12391,N_13377);
nand U15761 (N_15761,N_13857,N_13549);
and U15762 (N_15762,N_13613,N_13856);
or U15763 (N_15763,N_12854,N_13791);
and U15764 (N_15764,N_13306,N_13022);
nor U15765 (N_15765,N_12161,N_13261);
xor U15766 (N_15766,N_12934,N_12833);
xnor U15767 (N_15767,N_12867,N_13483);
and U15768 (N_15768,N_13629,N_12100);
or U15769 (N_15769,N_12069,N_12345);
xnor U15770 (N_15770,N_12379,N_12511);
nand U15771 (N_15771,N_12911,N_13734);
nand U15772 (N_15772,N_13556,N_12739);
or U15773 (N_15773,N_13247,N_12207);
xor U15774 (N_15774,N_13037,N_13424);
or U15775 (N_15775,N_13861,N_13835);
and U15776 (N_15776,N_12049,N_13897);
or U15777 (N_15777,N_12535,N_12737);
and U15778 (N_15778,N_13866,N_13531);
and U15779 (N_15779,N_12983,N_12898);
nor U15780 (N_15780,N_13418,N_13006);
nand U15781 (N_15781,N_13706,N_13118);
or U15782 (N_15782,N_13201,N_12497);
xnor U15783 (N_15783,N_12833,N_13775);
nor U15784 (N_15784,N_13022,N_12330);
nand U15785 (N_15785,N_12797,N_13227);
xor U15786 (N_15786,N_13977,N_13523);
and U15787 (N_15787,N_13335,N_13593);
nand U15788 (N_15788,N_12722,N_13052);
and U15789 (N_15789,N_12086,N_12661);
xor U15790 (N_15790,N_12141,N_12778);
or U15791 (N_15791,N_12123,N_12819);
xnor U15792 (N_15792,N_13732,N_13125);
xor U15793 (N_15793,N_12561,N_13492);
or U15794 (N_15794,N_13639,N_12578);
or U15795 (N_15795,N_12963,N_13864);
xor U15796 (N_15796,N_12879,N_12624);
xor U15797 (N_15797,N_12550,N_13417);
nand U15798 (N_15798,N_13128,N_13747);
nand U15799 (N_15799,N_13238,N_12195);
nor U15800 (N_15800,N_12489,N_13589);
or U15801 (N_15801,N_12419,N_13922);
nor U15802 (N_15802,N_12921,N_12556);
and U15803 (N_15803,N_12754,N_12773);
or U15804 (N_15804,N_12013,N_13245);
nor U15805 (N_15805,N_12548,N_13888);
nor U15806 (N_15806,N_12517,N_12693);
nand U15807 (N_15807,N_13901,N_13550);
nor U15808 (N_15808,N_12830,N_13721);
nor U15809 (N_15809,N_13538,N_12194);
and U15810 (N_15810,N_13109,N_13791);
and U15811 (N_15811,N_13382,N_12927);
nor U15812 (N_15812,N_12756,N_13744);
nor U15813 (N_15813,N_12713,N_13480);
nor U15814 (N_15814,N_12985,N_13646);
and U15815 (N_15815,N_12983,N_13970);
or U15816 (N_15816,N_12841,N_13410);
and U15817 (N_15817,N_13356,N_13186);
nand U15818 (N_15818,N_13638,N_12718);
xnor U15819 (N_15819,N_13676,N_13972);
nor U15820 (N_15820,N_13700,N_12064);
and U15821 (N_15821,N_12593,N_12346);
nand U15822 (N_15822,N_13383,N_12321);
nand U15823 (N_15823,N_12930,N_13126);
nor U15824 (N_15824,N_13846,N_13251);
xnor U15825 (N_15825,N_12329,N_13177);
nand U15826 (N_15826,N_13385,N_13221);
nor U15827 (N_15827,N_12419,N_13098);
nand U15828 (N_15828,N_13922,N_12832);
xnor U15829 (N_15829,N_13166,N_13081);
xnor U15830 (N_15830,N_13788,N_12589);
nand U15831 (N_15831,N_13405,N_12411);
and U15832 (N_15832,N_12056,N_13105);
nor U15833 (N_15833,N_13941,N_13581);
or U15834 (N_15834,N_12699,N_13380);
xor U15835 (N_15835,N_13587,N_12368);
xor U15836 (N_15836,N_13640,N_12780);
nand U15837 (N_15837,N_12402,N_13220);
nor U15838 (N_15838,N_12803,N_12258);
nand U15839 (N_15839,N_12643,N_13325);
and U15840 (N_15840,N_13357,N_13584);
xor U15841 (N_15841,N_12866,N_12663);
nand U15842 (N_15842,N_13140,N_12972);
nor U15843 (N_15843,N_12903,N_12193);
and U15844 (N_15844,N_13217,N_12522);
xnor U15845 (N_15845,N_12588,N_12001);
xnor U15846 (N_15846,N_12444,N_12648);
nand U15847 (N_15847,N_12148,N_12283);
and U15848 (N_15848,N_13893,N_13384);
nor U15849 (N_15849,N_12948,N_13339);
xor U15850 (N_15850,N_13112,N_12625);
or U15851 (N_15851,N_12407,N_12212);
nor U15852 (N_15852,N_12073,N_12980);
nand U15853 (N_15853,N_12486,N_12146);
xor U15854 (N_15854,N_13110,N_12095);
nand U15855 (N_15855,N_13082,N_13406);
xnor U15856 (N_15856,N_12577,N_13991);
or U15857 (N_15857,N_12907,N_12414);
xor U15858 (N_15858,N_13111,N_13260);
nand U15859 (N_15859,N_13149,N_13719);
nor U15860 (N_15860,N_12592,N_13148);
and U15861 (N_15861,N_12454,N_12953);
xor U15862 (N_15862,N_12805,N_13473);
or U15863 (N_15863,N_13221,N_13629);
nor U15864 (N_15864,N_13339,N_13317);
or U15865 (N_15865,N_13902,N_12837);
and U15866 (N_15866,N_12176,N_12056);
nand U15867 (N_15867,N_13625,N_12851);
or U15868 (N_15868,N_12209,N_13412);
xor U15869 (N_15869,N_12872,N_12619);
or U15870 (N_15870,N_12225,N_12096);
and U15871 (N_15871,N_13417,N_12043);
nand U15872 (N_15872,N_13333,N_13878);
and U15873 (N_15873,N_13185,N_13761);
nand U15874 (N_15874,N_12917,N_13663);
and U15875 (N_15875,N_12725,N_13294);
nand U15876 (N_15876,N_12221,N_13591);
xnor U15877 (N_15877,N_12623,N_13134);
xnor U15878 (N_15878,N_13762,N_12656);
and U15879 (N_15879,N_12867,N_12124);
nor U15880 (N_15880,N_13161,N_12889);
or U15881 (N_15881,N_13471,N_13067);
nand U15882 (N_15882,N_12586,N_13837);
nor U15883 (N_15883,N_13322,N_13427);
and U15884 (N_15884,N_13227,N_12222);
or U15885 (N_15885,N_12132,N_13727);
nand U15886 (N_15886,N_12016,N_13252);
nand U15887 (N_15887,N_12734,N_13398);
and U15888 (N_15888,N_13236,N_12439);
nor U15889 (N_15889,N_12377,N_12790);
and U15890 (N_15890,N_12729,N_13663);
or U15891 (N_15891,N_13994,N_13451);
and U15892 (N_15892,N_13318,N_13948);
or U15893 (N_15893,N_12949,N_13502);
xnor U15894 (N_15894,N_12270,N_13366);
nand U15895 (N_15895,N_12666,N_13259);
and U15896 (N_15896,N_12674,N_12393);
xnor U15897 (N_15897,N_12588,N_12343);
nor U15898 (N_15898,N_12514,N_13431);
nor U15899 (N_15899,N_13248,N_12854);
xnor U15900 (N_15900,N_12600,N_13028);
nor U15901 (N_15901,N_13598,N_13982);
nor U15902 (N_15902,N_12898,N_13705);
and U15903 (N_15903,N_13613,N_13768);
xnor U15904 (N_15904,N_12467,N_12834);
and U15905 (N_15905,N_12450,N_13347);
or U15906 (N_15906,N_12028,N_12691);
nand U15907 (N_15907,N_12617,N_13050);
nand U15908 (N_15908,N_13453,N_12672);
nor U15909 (N_15909,N_13502,N_12432);
nor U15910 (N_15910,N_13846,N_12540);
or U15911 (N_15911,N_12058,N_13287);
and U15912 (N_15912,N_12807,N_13992);
or U15913 (N_15913,N_13935,N_13950);
nor U15914 (N_15914,N_13745,N_12347);
xnor U15915 (N_15915,N_13541,N_12239);
or U15916 (N_15916,N_13344,N_12321);
and U15917 (N_15917,N_13027,N_12790);
and U15918 (N_15918,N_13863,N_13185);
or U15919 (N_15919,N_12321,N_12138);
xor U15920 (N_15920,N_13824,N_12180);
or U15921 (N_15921,N_12935,N_12691);
xor U15922 (N_15922,N_12746,N_12095);
xor U15923 (N_15923,N_13995,N_12213);
nor U15924 (N_15924,N_12498,N_12978);
xor U15925 (N_15925,N_12381,N_13196);
and U15926 (N_15926,N_12046,N_12821);
or U15927 (N_15927,N_13170,N_13415);
nand U15928 (N_15928,N_13564,N_12482);
and U15929 (N_15929,N_12095,N_12591);
and U15930 (N_15930,N_12789,N_12442);
or U15931 (N_15931,N_12860,N_13362);
nand U15932 (N_15932,N_12193,N_12250);
nor U15933 (N_15933,N_12387,N_13590);
xor U15934 (N_15934,N_12073,N_13894);
xor U15935 (N_15935,N_13950,N_12200);
or U15936 (N_15936,N_13902,N_13516);
xnor U15937 (N_15937,N_12375,N_13254);
xnor U15938 (N_15938,N_13930,N_12769);
nor U15939 (N_15939,N_13655,N_12068);
nand U15940 (N_15940,N_12855,N_12496);
and U15941 (N_15941,N_12346,N_12330);
and U15942 (N_15942,N_13320,N_12673);
and U15943 (N_15943,N_13741,N_12458);
and U15944 (N_15944,N_13937,N_12408);
xnor U15945 (N_15945,N_12503,N_12426);
xnor U15946 (N_15946,N_13257,N_13084);
nand U15947 (N_15947,N_13294,N_13743);
nand U15948 (N_15948,N_12659,N_12274);
nor U15949 (N_15949,N_13048,N_13796);
nand U15950 (N_15950,N_13352,N_13908);
xor U15951 (N_15951,N_13282,N_12024);
and U15952 (N_15952,N_12480,N_13214);
and U15953 (N_15953,N_13954,N_13629);
or U15954 (N_15954,N_13542,N_12118);
or U15955 (N_15955,N_13927,N_13204);
and U15956 (N_15956,N_13282,N_13893);
nand U15957 (N_15957,N_12874,N_13965);
xnor U15958 (N_15958,N_12236,N_12277);
or U15959 (N_15959,N_12295,N_13959);
and U15960 (N_15960,N_13686,N_12127);
nor U15961 (N_15961,N_13045,N_12228);
and U15962 (N_15962,N_12454,N_12312);
xnor U15963 (N_15963,N_13341,N_12193);
nor U15964 (N_15964,N_12496,N_13982);
xnor U15965 (N_15965,N_13066,N_12353);
and U15966 (N_15966,N_13774,N_12960);
xnor U15967 (N_15967,N_12008,N_12976);
or U15968 (N_15968,N_12711,N_12137);
and U15969 (N_15969,N_12038,N_13201);
nor U15970 (N_15970,N_13000,N_12779);
nor U15971 (N_15971,N_13108,N_13791);
nor U15972 (N_15972,N_12007,N_12164);
nor U15973 (N_15973,N_13385,N_13329);
nand U15974 (N_15974,N_12756,N_12831);
and U15975 (N_15975,N_12132,N_13292);
or U15976 (N_15976,N_12840,N_13974);
and U15977 (N_15977,N_13635,N_13860);
xnor U15978 (N_15978,N_13590,N_13937);
nand U15979 (N_15979,N_13386,N_12699);
nor U15980 (N_15980,N_13948,N_12419);
nor U15981 (N_15981,N_13374,N_13704);
nand U15982 (N_15982,N_12060,N_12609);
xnor U15983 (N_15983,N_12600,N_12335);
nor U15984 (N_15984,N_12346,N_13991);
and U15985 (N_15985,N_13782,N_13330);
xor U15986 (N_15986,N_13121,N_12068);
nand U15987 (N_15987,N_13107,N_12446);
nand U15988 (N_15988,N_12951,N_12056);
nand U15989 (N_15989,N_13152,N_13983);
nand U15990 (N_15990,N_12594,N_13470);
nand U15991 (N_15991,N_13935,N_12535);
and U15992 (N_15992,N_13989,N_13438);
or U15993 (N_15993,N_12288,N_13431);
nor U15994 (N_15994,N_13895,N_12983);
nand U15995 (N_15995,N_13203,N_13760);
and U15996 (N_15996,N_13705,N_13559);
and U15997 (N_15997,N_13434,N_12093);
xnor U15998 (N_15998,N_12080,N_13264);
nand U15999 (N_15999,N_12833,N_13766);
xnor U16000 (N_16000,N_15647,N_15557);
or U16001 (N_16001,N_15899,N_15372);
or U16002 (N_16002,N_15287,N_15247);
or U16003 (N_16003,N_14236,N_15397);
nor U16004 (N_16004,N_14345,N_14352);
nand U16005 (N_16005,N_14517,N_15875);
nand U16006 (N_16006,N_15742,N_15982);
xor U16007 (N_16007,N_14976,N_15399);
nand U16008 (N_16008,N_14753,N_15869);
or U16009 (N_16009,N_14578,N_14566);
and U16010 (N_16010,N_15333,N_14619);
or U16011 (N_16011,N_15022,N_15893);
nand U16012 (N_16012,N_15963,N_14128);
or U16013 (N_16013,N_14932,N_14375);
and U16014 (N_16014,N_15428,N_15579);
and U16015 (N_16015,N_15745,N_14823);
nor U16016 (N_16016,N_14110,N_14290);
or U16017 (N_16017,N_15817,N_14704);
nor U16018 (N_16018,N_15794,N_15880);
xor U16019 (N_16019,N_14489,N_14938);
nand U16020 (N_16020,N_15774,N_15970);
nor U16021 (N_16021,N_15635,N_14648);
and U16022 (N_16022,N_15180,N_14701);
nand U16023 (N_16023,N_14802,N_15531);
nand U16024 (N_16024,N_14668,N_15525);
nor U16025 (N_16025,N_14356,N_14847);
nor U16026 (N_16026,N_15427,N_15024);
xnor U16027 (N_16027,N_14913,N_14385);
nor U16028 (N_16028,N_14059,N_14123);
and U16029 (N_16029,N_14867,N_15274);
or U16030 (N_16030,N_14732,N_14239);
nand U16031 (N_16031,N_15425,N_14889);
nor U16032 (N_16032,N_14731,N_15409);
or U16033 (N_16033,N_15757,N_14049);
nand U16034 (N_16034,N_15270,N_14971);
xor U16035 (N_16035,N_14167,N_14705);
nor U16036 (N_16036,N_14429,N_15596);
nor U16037 (N_16037,N_15373,N_14979);
xor U16038 (N_16038,N_14945,N_14189);
nor U16039 (N_16039,N_14198,N_15710);
xor U16040 (N_16040,N_15407,N_15637);
or U16041 (N_16041,N_15888,N_14816);
nor U16042 (N_16042,N_15789,N_15153);
or U16043 (N_16043,N_15870,N_15175);
and U16044 (N_16044,N_14699,N_15844);
and U16045 (N_16045,N_15071,N_15630);
or U16046 (N_16046,N_14591,N_14496);
nor U16047 (N_16047,N_14240,N_14102);
and U16048 (N_16048,N_15897,N_14069);
xor U16049 (N_16049,N_14113,N_15898);
and U16050 (N_16050,N_15191,N_14819);
xnor U16051 (N_16051,N_14691,N_14320);
or U16052 (N_16052,N_14514,N_15879);
and U16053 (N_16053,N_15594,N_15959);
nand U16054 (N_16054,N_15536,N_15743);
or U16055 (N_16055,N_14106,N_15940);
xnor U16056 (N_16056,N_14277,N_14894);
nor U16057 (N_16057,N_15656,N_15593);
nor U16058 (N_16058,N_14808,N_14287);
and U16059 (N_16059,N_14525,N_14444);
or U16060 (N_16060,N_14233,N_14117);
nor U16061 (N_16061,N_15118,N_14792);
and U16062 (N_16062,N_14549,N_14223);
and U16063 (N_16063,N_14683,N_14048);
nor U16064 (N_16064,N_14494,N_14582);
nand U16065 (N_16065,N_15735,N_15986);
and U16066 (N_16066,N_14775,N_15586);
xnor U16067 (N_16067,N_15734,N_15384);
and U16068 (N_16068,N_14219,N_15008);
and U16069 (N_16069,N_14641,N_15129);
nor U16070 (N_16070,N_14773,N_14101);
or U16071 (N_16071,N_14221,N_14646);
or U16072 (N_16072,N_15361,N_14642);
or U16073 (N_16073,N_15324,N_14053);
or U16074 (N_16074,N_14120,N_14937);
xnor U16075 (N_16075,N_14562,N_15808);
xnor U16076 (N_16076,N_15674,N_15758);
or U16077 (N_16077,N_14697,N_15631);
nand U16078 (N_16078,N_15646,N_14666);
nor U16079 (N_16079,N_15605,N_15379);
xor U16080 (N_16080,N_15436,N_14321);
nor U16081 (N_16081,N_15755,N_15194);
nor U16082 (N_16082,N_14232,N_14686);
and U16083 (N_16083,N_15339,N_15500);
xnor U16084 (N_16084,N_15983,N_14528);
or U16085 (N_16085,N_14421,N_15860);
nor U16086 (N_16086,N_15106,N_15414);
or U16087 (N_16087,N_14279,N_14625);
and U16088 (N_16088,N_15469,N_14095);
xor U16089 (N_16089,N_15042,N_15989);
nand U16090 (N_16090,N_15169,N_15447);
xor U16091 (N_16091,N_15606,N_15292);
nor U16092 (N_16092,N_14785,N_14185);
nand U16093 (N_16093,N_15771,N_15878);
or U16094 (N_16094,N_15722,N_14361);
or U16095 (N_16095,N_15341,N_15289);
and U16096 (N_16096,N_15137,N_14651);
or U16097 (N_16097,N_14903,N_14464);
xor U16098 (N_16098,N_15634,N_15435);
xnor U16099 (N_16099,N_14853,N_15249);
xor U16100 (N_16100,N_15306,N_15505);
xnor U16101 (N_16101,N_15615,N_15573);
nor U16102 (N_16102,N_15255,N_14963);
nor U16103 (N_16103,N_14466,N_14615);
xor U16104 (N_16104,N_14427,N_14249);
nand U16105 (N_16105,N_14974,N_14492);
nor U16106 (N_16106,N_14687,N_15592);
nand U16107 (N_16107,N_15296,N_15811);
nor U16108 (N_16108,N_15651,N_15585);
xnor U16109 (N_16109,N_14506,N_14431);
or U16110 (N_16110,N_14784,N_14138);
or U16111 (N_16111,N_14447,N_14378);
and U16112 (N_16112,N_14599,N_14748);
nor U16113 (N_16113,N_15784,N_15250);
nand U16114 (N_16114,N_15465,N_15291);
and U16115 (N_16115,N_14843,N_15495);
or U16116 (N_16116,N_15739,N_14084);
nand U16117 (N_16117,N_14146,N_14220);
or U16118 (N_16118,N_14706,N_14303);
nand U16119 (N_16119,N_14688,N_15666);
or U16120 (N_16120,N_14374,N_15038);
xor U16121 (N_16121,N_14746,N_15028);
xor U16122 (N_16122,N_15921,N_14139);
or U16123 (N_16123,N_15183,N_15261);
and U16124 (N_16124,N_14271,N_14398);
xor U16125 (N_16125,N_15491,N_15891);
and U16126 (N_16126,N_15763,N_15812);
xnor U16127 (N_16127,N_14793,N_15377);
nor U16128 (N_16128,N_14907,N_15124);
and U16129 (N_16129,N_14891,N_15972);
xor U16130 (N_16130,N_15081,N_14174);
xnor U16131 (N_16131,N_15325,N_14594);
xnor U16132 (N_16132,N_14597,N_14912);
nor U16133 (N_16133,N_14344,N_14803);
xor U16134 (N_16134,N_14608,N_14264);
xor U16135 (N_16135,N_14631,N_15098);
nand U16136 (N_16136,N_14719,N_15564);
and U16137 (N_16137,N_14136,N_15257);
or U16138 (N_16138,N_15696,N_14436);
and U16139 (N_16139,N_15093,N_15562);
nor U16140 (N_16140,N_14116,N_15913);
and U16141 (N_16141,N_15003,N_14424);
and U16142 (N_16142,N_14411,N_14788);
and U16143 (N_16143,N_15352,N_14024);
nor U16144 (N_16144,N_15541,N_14399);
xnor U16145 (N_16145,N_14484,N_14851);
and U16146 (N_16146,N_14040,N_14939);
nor U16147 (N_16147,N_14677,N_14030);
or U16148 (N_16148,N_14010,N_14448);
xor U16149 (N_16149,N_15321,N_14868);
or U16150 (N_16150,N_14195,N_15707);
and U16151 (N_16151,N_14289,N_15062);
or U16152 (N_16152,N_14629,N_15991);
nor U16153 (N_16153,N_15344,N_15569);
nand U16154 (N_16154,N_14414,N_15506);
xor U16155 (N_16155,N_14897,N_14884);
xnor U16156 (N_16156,N_14125,N_15697);
nor U16157 (N_16157,N_15919,N_15240);
nor U16158 (N_16158,N_14310,N_14451);
and U16159 (N_16159,N_14710,N_14592);
nand U16160 (N_16160,N_14127,N_14355);
nor U16161 (N_16161,N_15480,N_14986);
nand U16162 (N_16162,N_14111,N_15149);
and U16163 (N_16163,N_14933,N_15957);
nor U16164 (N_16164,N_15104,N_14047);
or U16165 (N_16165,N_14767,N_15351);
xnor U16166 (N_16166,N_15978,N_14627);
nor U16167 (N_16167,N_14899,N_15589);
nor U16168 (N_16168,N_14953,N_14993);
xor U16169 (N_16169,N_15984,N_15790);
nand U16170 (N_16170,N_14812,N_15552);
nand U16171 (N_16171,N_15601,N_14459);
nand U16172 (N_16172,N_15501,N_15026);
nand U16173 (N_16173,N_14299,N_14927);
or U16174 (N_16174,N_15155,N_15803);
nand U16175 (N_16175,N_14760,N_14322);
or U16176 (N_16176,N_14527,N_14995);
nand U16177 (N_16177,N_15456,N_15723);
and U16178 (N_16178,N_15229,N_14382);
nand U16179 (N_16179,N_14610,N_15969);
and U16180 (N_16180,N_14863,N_15788);
nor U16181 (N_16181,N_14243,N_15752);
nor U16182 (N_16182,N_15086,N_14401);
and U16183 (N_16183,N_14441,N_14028);
nor U16184 (N_16184,N_14650,N_14634);
or U16185 (N_16185,N_14073,N_15199);
xnor U16186 (N_16186,N_14476,N_15727);
and U16187 (N_16187,N_14256,N_15020);
nor U16188 (N_16188,N_15826,N_14300);
or U16189 (N_16189,N_15222,N_15680);
nor U16190 (N_16190,N_15205,N_14392);
and U16191 (N_16191,N_14777,N_15850);
nor U16192 (N_16192,N_14914,N_14538);
or U16193 (N_16193,N_15203,N_14319);
nor U16194 (N_16194,N_15614,N_15968);
nor U16195 (N_16195,N_14600,N_14042);
nor U16196 (N_16196,N_15625,N_14328);
nand U16197 (N_16197,N_15286,N_14413);
nand U16198 (N_16198,N_14131,N_14789);
and U16199 (N_16199,N_15034,N_14855);
or U16200 (N_16200,N_14928,N_14032);
xor U16201 (N_16201,N_14261,N_14992);
nor U16202 (N_16202,N_15507,N_14662);
xnor U16203 (N_16203,N_15396,N_14561);
xnor U16204 (N_16204,N_14272,N_14568);
and U16205 (N_16205,N_14104,N_14961);
nand U16206 (N_16206,N_14021,N_15871);
nor U16207 (N_16207,N_15157,N_15740);
nand U16208 (N_16208,N_14917,N_15493);
nand U16209 (N_16209,N_14529,N_14554);
and U16210 (N_16210,N_14013,N_14726);
xor U16211 (N_16211,N_14770,N_14759);
nand U16212 (N_16212,N_15942,N_15559);
nor U16213 (N_16213,N_15017,N_15931);
or U16214 (N_16214,N_14334,N_14340);
or U16215 (N_16215,N_15027,N_14880);
nand U16216 (N_16216,N_15954,N_15235);
and U16217 (N_16217,N_14100,N_14052);
and U16218 (N_16218,N_15336,N_15934);
and U16219 (N_16219,N_14029,N_15643);
and U16220 (N_16220,N_14479,N_14061);
nand U16221 (N_16221,N_14665,N_15295);
xnor U16222 (N_16222,N_14311,N_15300);
and U16223 (N_16223,N_15702,N_14780);
xnor U16224 (N_16224,N_14535,N_14983);
xnor U16225 (N_16225,N_14285,N_14577);
xnor U16226 (N_16226,N_15809,N_15842);
xnor U16227 (N_16227,N_15574,N_14446);
and U16228 (N_16228,N_15294,N_15489);
nor U16229 (N_16229,N_15563,N_14596);
nor U16230 (N_16230,N_14434,N_15956);
nand U16231 (N_16231,N_15170,N_14990);
nand U16232 (N_16232,N_14004,N_14003);
and U16233 (N_16233,N_14703,N_15187);
nand U16234 (N_16234,N_14199,N_15549);
nor U16235 (N_16235,N_15004,N_14327);
and U16236 (N_16236,N_14016,N_14358);
and U16237 (N_16237,N_14604,N_15577);
nand U16238 (N_16238,N_14893,N_15089);
nor U16239 (N_16239,N_14071,N_15304);
nor U16240 (N_16240,N_15896,N_15141);
and U16241 (N_16241,N_15000,N_14055);
nand U16242 (N_16242,N_14291,N_15314);
or U16243 (N_16243,N_15219,N_15620);
and U16244 (N_16244,N_15402,N_14150);
or U16245 (N_16245,N_14583,N_14294);
nor U16246 (N_16246,N_15953,N_14196);
nand U16247 (N_16247,N_14950,N_14350);
or U16248 (N_16248,N_15009,N_15484);
nand U16249 (N_16249,N_15091,N_14715);
nor U16250 (N_16250,N_15193,N_15964);
or U16251 (N_16251,N_15163,N_15225);
or U16252 (N_16252,N_15168,N_14957);
and U16253 (N_16253,N_14533,N_15952);
xor U16254 (N_16254,N_14367,N_15439);
nor U16255 (N_16255,N_14716,N_15400);
nand U16256 (N_16256,N_15437,N_15772);
nand U16257 (N_16257,N_14837,N_14829);
nand U16258 (N_16258,N_14524,N_14832);
and U16259 (N_16259,N_14409,N_15522);
or U16260 (N_16260,N_15068,N_15328);
or U16261 (N_16261,N_15025,N_14712);
and U16262 (N_16262,N_15543,N_14519);
nor U16263 (N_16263,N_14203,N_15512);
nand U16264 (N_16264,N_14143,N_15472);
or U16265 (N_16265,N_14944,N_15408);
nand U16266 (N_16266,N_15410,N_14909);
and U16267 (N_16267,N_15482,N_15041);
nand U16268 (N_16268,N_14833,N_15116);
nand U16269 (N_16269,N_15530,N_14551);
nor U16270 (N_16270,N_14564,N_15110);
nor U16271 (N_16271,N_14313,N_14363);
xor U16272 (N_16272,N_15502,N_15603);
or U16273 (N_16273,N_14204,N_14681);
nand U16274 (N_16274,N_15099,N_15622);
xnor U16275 (N_16275,N_15079,N_15002);
or U16276 (N_16276,N_15652,N_15883);
nor U16277 (N_16277,N_14735,N_14806);
nand U16278 (N_16278,N_14273,N_15477);
xor U16279 (N_16279,N_14636,N_14491);
and U16280 (N_16280,N_15908,N_15650);
and U16281 (N_16281,N_14137,N_14509);
nor U16282 (N_16282,N_14338,N_14145);
nor U16283 (N_16283,N_15115,N_14543);
nand U16284 (N_16284,N_14086,N_14941);
or U16285 (N_16285,N_15539,N_15417);
xor U16286 (N_16286,N_14002,N_14418);
nand U16287 (N_16287,N_14407,N_14623);
nor U16288 (N_16288,N_14864,N_14000);
and U16289 (N_16289,N_15738,N_14486);
xnor U16290 (N_16290,N_15545,N_14559);
nor U16291 (N_16291,N_15253,N_14955);
xor U16292 (N_16292,N_14384,N_14756);
xor U16293 (N_16293,N_14191,N_15192);
nand U16294 (N_16294,N_14018,N_14540);
xor U16295 (N_16295,N_15648,N_14121);
or U16296 (N_16296,N_14711,N_15362);
or U16297 (N_16297,N_15876,N_15103);
or U16298 (N_16298,N_14947,N_15985);
nor U16299 (N_16299,N_15977,N_15101);
nand U16300 (N_16300,N_15962,N_15468);
nand U16301 (N_16301,N_15462,N_14695);
nor U16302 (N_16302,N_14870,N_14357);
or U16303 (N_16303,N_15754,N_14848);
or U16304 (N_16304,N_15945,N_14815);
and U16305 (N_16305,N_15320,N_15102);
nor U16306 (N_16306,N_15166,N_14742);
or U16307 (N_16307,N_14675,N_14613);
or U16308 (N_16308,N_15750,N_14058);
nand U16309 (N_16309,N_15729,N_15698);
or U16310 (N_16310,N_14333,N_14275);
and U16311 (N_16311,N_15737,N_15457);
nor U16312 (N_16312,N_15242,N_14569);
and U16313 (N_16313,N_14638,N_14881);
xor U16314 (N_16314,N_14019,N_14173);
xnor U16315 (N_16315,N_14325,N_15466);
or U16316 (N_16316,N_14585,N_15829);
and U16317 (N_16317,N_15381,N_14680);
and U16318 (N_16318,N_15209,N_15868);
or U16319 (N_16319,N_15073,N_14453);
nand U16320 (N_16320,N_14406,N_15282);
nor U16321 (N_16321,N_15496,N_15127);
nor U16322 (N_16322,N_15867,N_15759);
or U16323 (N_16323,N_15332,N_15052);
and U16324 (N_16324,N_15451,N_15418);
xor U16325 (N_16325,N_14498,N_14589);
nand U16326 (N_16326,N_15459,N_15591);
nand U16327 (N_16327,N_15901,N_14471);
xor U16328 (N_16328,N_14210,N_15715);
or U16329 (N_16329,N_15455,N_14088);
nand U16330 (N_16330,N_15335,N_15849);
xor U16331 (N_16331,N_14133,N_15690);
nor U16332 (N_16332,N_15950,N_14495);
nor U16333 (N_16333,N_14628,N_14532);
nor U16334 (N_16334,N_14520,N_15830);
and U16335 (N_16335,N_14822,N_14366);
nor U16336 (N_16336,N_15914,N_15602);
or U16337 (N_16337,N_15354,N_14440);
xor U16338 (N_16338,N_15910,N_14056);
xor U16339 (N_16339,N_14946,N_15391);
and U16340 (N_16340,N_14126,N_15616);
or U16341 (N_16341,N_14316,N_15857);
nor U16342 (N_16342,N_14461,N_15224);
nand U16343 (N_16343,N_15277,N_15252);
nand U16344 (N_16344,N_15481,N_15043);
xnor U16345 (N_16345,N_14373,N_15509);
or U16346 (N_16346,N_14033,N_14419);
xor U16347 (N_16347,N_15265,N_14685);
and U16348 (N_16348,N_14852,N_14635);
or U16349 (N_16349,N_14159,N_14389);
or U16350 (N_16350,N_14750,N_14330);
xnor U16351 (N_16351,N_14902,N_15177);
nand U16352 (N_16352,N_14188,N_14149);
nand U16353 (N_16353,N_14764,N_14670);
nor U16354 (N_16354,N_14781,N_14339);
nor U16355 (N_16355,N_15799,N_15773);
nand U16356 (N_16356,N_15302,N_14626);
nor U16357 (N_16357,N_15390,N_14215);
xnor U16358 (N_16358,N_15267,N_15313);
xnor U16359 (N_16359,N_15864,N_15995);
xnor U16360 (N_16360,N_15892,N_15230);
and U16361 (N_16361,N_14603,N_14107);
or U16362 (N_16362,N_14964,N_14014);
and U16363 (N_16363,N_15162,N_15076);
and U16364 (N_16364,N_15094,N_15831);
xnor U16365 (N_16365,N_14151,N_15244);
nand U16366 (N_16366,N_14276,N_14546);
nand U16367 (N_16367,N_14644,N_15279);
nor U16368 (N_16368,N_15519,N_14765);
xor U16369 (N_16369,N_14882,N_14283);
xnor U16370 (N_16370,N_14904,N_15285);
xor U16371 (N_16371,N_14214,N_15444);
nand U16372 (N_16372,N_15546,N_15654);
xor U16373 (N_16373,N_15273,N_14423);
and U16374 (N_16374,N_14175,N_14072);
and U16375 (N_16375,N_14972,N_14521);
nand U16376 (N_16376,N_14224,N_15672);
and U16377 (N_16377,N_14534,N_15973);
nand U16378 (N_16378,N_14335,N_15420);
nor U16379 (N_16379,N_15884,N_14544);
nand U16380 (N_16380,N_15392,N_15143);
nand U16381 (N_16381,N_15121,N_14207);
or U16382 (N_16382,N_15526,N_14255);
nand U16383 (N_16383,N_15037,N_15951);
nor U16384 (N_16384,N_14797,N_14557);
nor U16385 (N_16385,N_15975,N_15718);
nor U16386 (N_16386,N_14011,N_14877);
or U16387 (N_16387,N_14751,N_15571);
nor U16388 (N_16388,N_15236,N_15368);
nand U16389 (N_16389,N_14836,N_14402);
nand U16390 (N_16390,N_14553,N_15657);
nand U16391 (N_16391,N_15767,N_15612);
nand U16392 (N_16392,N_15107,N_14241);
or U16393 (N_16393,N_15846,N_14380);
and U16394 (N_16394,N_15558,N_14508);
or U16395 (N_16395,N_14462,N_14831);
and U16396 (N_16396,N_14845,N_14722);
nor U16397 (N_16397,N_14152,N_14298);
xor U16398 (N_16398,N_15889,N_14799);
and U16399 (N_16399,N_15663,N_14351);
or U16400 (N_16400,N_15785,N_14244);
and U16401 (N_16401,N_14229,N_14844);
xnor U16402 (N_16402,N_14027,N_15713);
nand U16403 (N_16403,N_14682,N_14284);
xor U16404 (N_16404,N_14170,N_14739);
xor U16405 (N_16405,N_15597,N_14396);
and U16406 (N_16406,N_14200,N_14342);
nand U16407 (N_16407,N_15958,N_14645);
nor U16408 (N_16408,N_15080,N_14570);
xnor U16409 (N_16409,N_15665,N_15238);
nand U16410 (N_16410,N_14160,N_15717);
nand U16411 (N_16411,N_14359,N_15258);
nor U16412 (N_16412,N_15376,N_14977);
and U16413 (N_16413,N_15035,N_14050);
or U16414 (N_16414,N_14692,N_14856);
xnor U16415 (N_16415,N_14371,N_15303);
and U16416 (N_16416,N_14892,N_15355);
nor U16417 (N_16417,N_14573,N_15403);
or U16418 (N_16418,N_14001,N_15479);
nor U16419 (N_16419,N_14772,N_14368);
nor U16420 (N_16420,N_14346,N_15007);
nor U16421 (N_16421,N_15529,N_15448);
and U16422 (N_16422,N_15036,N_14839);
or U16423 (N_16423,N_15269,N_15033);
xnor U16424 (N_16424,N_15185,N_15587);
nor U16425 (N_16425,N_14761,N_15382);
and U16426 (N_16426,N_14728,N_15318);
or U16427 (N_16427,N_15572,N_15393);
or U16428 (N_16428,N_15768,N_14251);
xor U16429 (N_16429,N_15019,N_15746);
or U16430 (N_16430,N_14262,N_15761);
nor U16431 (N_16431,N_14168,N_15640);
nor U16432 (N_16432,N_15014,N_15056);
or U16433 (N_16433,N_14846,N_15415);
nand U16434 (N_16434,N_15173,N_14581);
or U16435 (N_16435,N_15912,N_15450);
or U16436 (N_16436,N_15171,N_15161);
nand U16437 (N_16437,N_14245,N_14022);
nand U16438 (N_16438,N_14743,N_15204);
xnor U16439 (N_16439,N_14266,N_15720);
or U16440 (N_16440,N_14208,N_15751);
nand U16441 (N_16441,N_14179,N_15781);
or U16442 (N_16442,N_14091,N_14511);
xor U16443 (N_16443,N_14593,N_14394);
nand U16444 (N_16444,N_15851,N_15946);
nor U16445 (N_16445,N_14135,N_15406);
or U16446 (N_16446,N_14388,N_15366);
nand U16447 (N_16447,N_14672,N_14984);
nand U16448 (N_16448,N_15638,N_15966);
xnor U16449 (N_16449,N_14607,N_14075);
nand U16450 (N_16450,N_15618,N_14166);
xnor U16451 (N_16451,N_15461,N_15974);
xor U16452 (N_16452,N_15695,N_14659);
or U16453 (N_16453,N_14456,N_15057);
xor U16454 (N_16454,N_14369,N_15109);
nor U16455 (N_16455,N_15580,N_15590);
or U16456 (N_16456,N_14194,N_14305);
xor U16457 (N_16457,N_14959,N_15686);
nand U16458 (N_16458,N_15624,N_14099);
nand U16459 (N_16459,N_15350,N_15067);
nor U16460 (N_16460,N_15814,N_14437);
nor U16461 (N_16461,N_15677,N_15097);
or U16462 (N_16462,N_15824,N_14575);
and U16463 (N_16463,N_15327,N_15547);
nor U16464 (N_16464,N_14488,N_14940);
or U16465 (N_16465,N_14618,N_14910);
nand U16466 (N_16466,N_15906,N_14779);
nor U16467 (N_16467,N_14124,N_15488);
nor U16468 (N_16468,N_14841,N_15449);
nor U16469 (N_16469,N_14978,N_14744);
xor U16470 (N_16470,N_15948,N_15716);
xor U16471 (N_16471,N_15342,N_14526);
nand U16472 (N_16472,N_14624,N_15981);
or U16473 (N_16473,N_14336,N_15426);
nor U16474 (N_16474,N_15044,N_15976);
nand U16475 (N_16475,N_14376,N_14433);
or U16476 (N_16476,N_15440,N_15566);
xor U16477 (N_16477,N_15841,N_15711);
and U16478 (N_16478,N_14263,N_14747);
or U16479 (N_16479,N_14301,N_14714);
or U16480 (N_16480,N_15066,N_15923);
and U16481 (N_16481,N_15232,N_14122);
nor U16482 (N_16482,N_15049,N_15176);
or U16483 (N_16483,N_15941,N_15074);
nand U16484 (N_16484,N_14038,N_14827);
nor U16485 (N_16485,N_14838,N_14031);
or U16486 (N_16486,N_14994,N_15018);
nor U16487 (N_16487,N_15012,N_15508);
or U16488 (N_16488,N_14502,N_15560);
or U16489 (N_16489,N_15343,N_14490);
nand U16490 (N_16490,N_15221,N_14507);
and U16491 (N_16491,N_15241,N_14804);
xor U16492 (N_16492,N_15031,N_15706);
or U16493 (N_16493,N_15917,N_14567);
nand U16494 (N_16494,N_14468,N_15213);
and U16495 (N_16495,N_14609,N_15905);
or U16496 (N_16496,N_14309,N_15932);
xor U16497 (N_16497,N_14674,N_14397);
and U16498 (N_16498,N_14998,N_15992);
or U16499 (N_16499,N_14193,N_15865);
xor U16500 (N_16500,N_14684,N_15309);
xnor U16501 (N_16501,N_14826,N_15828);
xnor U16502 (N_16502,N_14046,N_14026);
or U16503 (N_16503,N_14782,N_14663);
xor U16504 (N_16504,N_15023,N_14721);
and U16505 (N_16505,N_14885,N_14671);
nor U16506 (N_16506,N_14850,N_15297);
and U16507 (N_16507,N_15126,N_15920);
nor U16508 (N_16508,N_15822,N_15565);
and U16509 (N_16509,N_14501,N_15212);
nand U16510 (N_16510,N_14017,N_15345);
nand U16511 (N_16511,N_15144,N_15548);
nand U16512 (N_16512,N_14201,N_14878);
xnor U16513 (N_16513,N_14970,N_15001);
nand U16514 (N_16514,N_14536,N_15394);
and U16515 (N_16515,N_15655,N_14405);
or U16516 (N_16516,N_14738,N_15206);
nor U16517 (N_16517,N_15900,N_14842);
or U16518 (N_16518,N_15188,N_14304);
and U16519 (N_16519,N_14144,N_15159);
xor U16520 (N_16520,N_14070,N_15764);
and U16521 (N_16521,N_15470,N_15979);
nand U16522 (N_16522,N_15272,N_14025);
and U16523 (N_16523,N_15211,N_15125);
or U16524 (N_16524,N_15401,N_14469);
nand U16525 (N_16525,N_14951,N_15112);
nor U16526 (N_16526,N_14515,N_14281);
nor U16527 (N_16527,N_14148,N_15123);
nand U16528 (N_16528,N_15217,N_15105);
nand U16529 (N_16529,N_14445,N_14840);
xor U16530 (N_16530,N_15092,N_14545);
nor U16531 (N_16531,N_14632,N_15725);
nor U16532 (N_16532,N_15485,N_15416);
or U16533 (N_16533,N_14326,N_15233);
and U16534 (N_16534,N_14176,N_14463);
or U16535 (N_16535,N_14481,N_15748);
nor U16536 (N_16536,N_14871,N_14595);
nand U16537 (N_16537,N_15980,N_14089);
and U16538 (N_16538,N_15852,N_14859);
xnor U16539 (N_16539,N_14916,N_15013);
or U16540 (N_16540,N_14778,N_15021);
or U16541 (N_16541,N_15190,N_14432);
and U16542 (N_16542,N_15237,N_15518);
nand U16543 (N_16543,N_14817,N_14769);
and U16544 (N_16544,N_14293,N_14548);
nand U16545 (N_16545,N_15524,N_14036);
nor U16546 (N_16546,N_15692,N_14087);
nand U16547 (N_16547,N_15227,N_14694);
xor U16548 (N_16548,N_14531,N_15645);
nor U16549 (N_16549,N_14713,N_15783);
nor U16550 (N_16550,N_15818,N_15108);
and U16551 (N_16551,N_14134,N_15681);
nor U16552 (N_16552,N_14297,N_14552);
xnor U16553 (N_16553,N_15312,N_15911);
nor U16554 (N_16554,N_15264,N_15122);
or U16555 (N_16555,N_15460,N_15786);
or U16556 (N_16556,N_15669,N_14158);
and U16557 (N_16557,N_15554,N_14365);
nand U16558 (N_16558,N_14857,N_15070);
nor U16559 (N_16559,N_15429,N_14154);
xnor U16560 (N_16560,N_15644,N_14470);
and U16561 (N_16561,N_15796,N_14639);
xnor U16562 (N_16562,N_15388,N_14354);
nor U16563 (N_16563,N_15639,N_15039);
or U16564 (N_16564,N_15072,N_15578);
and U16565 (N_16565,N_15576,N_14982);
and U16566 (N_16566,N_14206,N_15584);
xor U16567 (N_16567,N_15924,N_15172);
nor U16568 (N_16568,N_14317,N_15128);
nand U16569 (N_16569,N_15453,N_14873);
nand U16570 (N_16570,N_14966,N_15276);
nor U16571 (N_16571,N_14776,N_15676);
nor U16572 (N_16572,N_14094,N_15517);
and U16573 (N_16573,N_15197,N_14637);
nand U16574 (N_16574,N_15872,N_14347);
nand U16575 (N_16575,N_15156,N_15165);
and U16576 (N_16576,N_15938,N_14678);
xnor U16577 (N_16577,N_15138,N_15278);
and U16578 (N_16578,N_14090,N_14006);
or U16579 (N_16579,N_14924,N_15281);
nand U16580 (N_16580,N_14112,N_15550);
or U16581 (N_16581,N_15700,N_14888);
and U16582 (N_16582,N_15778,N_14455);
xor U16583 (N_16583,N_14919,N_15780);
xnor U16584 (N_16584,N_14343,N_14268);
or U16585 (N_16585,N_14755,N_15766);
nand U16586 (N_16586,N_14798,N_15854);
nor U16587 (N_16587,N_14835,N_15095);
xnor U16588 (N_16588,N_15894,N_15527);
or U16589 (N_16589,N_14679,N_14901);
nand U16590 (N_16590,N_15357,N_15551);
or U16591 (N_16591,N_15490,N_14667);
and U16592 (N_16592,N_14362,N_15999);
and U16593 (N_16593,N_15201,N_15553);
or U16594 (N_16594,N_15949,N_15843);
nand U16595 (N_16595,N_15475,N_14661);
nor U16596 (N_16596,N_14250,N_14428);
xor U16597 (N_16597,N_15486,N_15805);
xnor U16598 (N_16598,N_14169,N_15863);
nand U16599 (N_16599,N_15016,N_14943);
or U16600 (N_16600,N_14898,N_14766);
nand U16601 (N_16601,N_14230,N_14598);
and U16602 (N_16602,N_14956,N_14825);
nand U16603 (N_16603,N_14216,N_15895);
nand U16604 (N_16604,N_15685,N_15083);
or U16605 (N_16605,N_14274,N_14736);
nor U16606 (N_16606,N_14922,N_15542);
or U16607 (N_16607,N_15452,N_15256);
nand U16608 (N_16608,N_15806,N_14969);
or U16609 (N_16609,N_14190,N_15629);
nor U16610 (N_16610,N_15463,N_15434);
or U16611 (N_16611,N_14257,N_15521);
xor U16612 (N_16612,N_15323,N_15322);
nand U16613 (N_16613,N_14620,N_15378);
or U16614 (N_16614,N_15111,N_15326);
and U16615 (N_16615,N_14296,N_15389);
or U16616 (N_16616,N_14601,N_15065);
nand U16617 (N_16617,N_15096,N_14571);
or U16618 (N_16618,N_15186,N_15714);
and U16619 (N_16619,N_15356,N_14795);
or U16620 (N_16620,N_15833,N_15858);
and U16621 (N_16621,N_14973,N_15364);
and U16622 (N_16622,N_15928,N_14085);
nor U16623 (N_16623,N_14153,N_15661);
or U16624 (N_16624,N_15816,N_15015);
and U16625 (N_16625,N_14370,N_14114);
nor U16626 (N_16626,N_15499,N_14612);
nor U16627 (N_16627,N_15497,N_14260);
or U16628 (N_16628,N_15664,N_14062);
and U16629 (N_16629,N_14295,N_15228);
nand U16630 (N_16630,N_15855,N_14530);
and U16631 (N_16631,N_14602,N_14809);
nand U16632 (N_16632,N_15859,N_14866);
xor U16633 (N_16633,N_15215,N_15998);
and U16634 (N_16634,N_14246,N_15231);
and U16635 (N_16635,N_15653,N_15131);
nor U16636 (N_16636,N_15691,N_14875);
xnor U16637 (N_16637,N_14588,N_14876);
nor U16638 (N_16638,N_14348,N_14796);
and U16639 (N_16639,N_14403,N_15011);
nand U16640 (N_16640,N_15347,N_15063);
or U16641 (N_16641,N_15467,N_15904);
nor U16642 (N_16642,N_14824,N_15513);
nor U16643 (N_16643,N_14830,N_15607);
and U16644 (N_16644,N_14081,N_14222);
xor U16645 (N_16645,N_14905,N_14129);
and U16646 (N_16646,N_15311,N_15632);
and U16647 (N_16647,N_14872,N_14556);
or U16648 (N_16648,N_14109,N_14745);
nor U16649 (N_16649,N_15922,N_14740);
nand U16650 (N_16650,N_14079,N_14162);
nand U16651 (N_16651,N_15595,N_14555);
or U16652 (N_16652,N_15515,N_14814);
xnor U16653 (N_16653,N_14051,N_15747);
nand U16654 (N_16654,N_15433,N_14306);
nor U16655 (N_16655,N_14439,N_15712);
nand U16656 (N_16656,N_15365,N_14563);
or U16657 (N_16657,N_15413,N_15262);
nor U16658 (N_16658,N_15902,N_15610);
nor U16659 (N_16659,N_15167,N_14505);
or U16660 (N_16660,N_15259,N_14991);
or U16661 (N_16661,N_14252,N_14768);
nor U16662 (N_16662,N_14155,N_15280);
nor U16663 (N_16663,N_15682,N_15360);
xnor U16664 (N_16664,N_14586,N_14171);
nor U16665 (N_16665,N_15907,N_14954);
or U16666 (N_16666,N_15363,N_14387);
and U16667 (N_16667,N_15100,N_15120);
and U16668 (N_16668,N_15937,N_15588);
or U16669 (N_16669,N_15133,N_14660);
xnor U16670 (N_16670,N_15346,N_14630);
or U16671 (N_16671,N_15349,N_15623);
nand U16672 (N_16672,N_15198,N_14443);
xnor U16673 (N_16673,N_14377,N_14936);
and U16674 (N_16674,N_15820,N_14009);
or U16675 (N_16675,N_15756,N_15528);
nor U16676 (N_16676,N_15483,N_15117);
nor U16677 (N_16677,N_15135,N_14008);
nand U16678 (N_16678,N_14353,N_14513);
nand U16679 (N_16679,N_15329,N_15776);
nor U16680 (N_16680,N_14066,N_14654);
nor U16681 (N_16681,N_15848,N_14700);
or U16682 (N_16682,N_14805,N_14472);
nand U16683 (N_16683,N_15078,N_15662);
nand U16684 (N_16684,N_15423,N_15441);
and U16685 (N_16685,N_15837,N_15220);
and U16686 (N_16686,N_14288,N_14142);
or U16687 (N_16687,N_14865,N_14364);
or U16688 (N_16688,N_15840,N_15158);
xnor U16689 (N_16689,N_14989,N_14269);
or U16690 (N_16690,N_14247,N_14093);
xnor U16691 (N_16691,N_14887,N_15770);
nand U16692 (N_16692,N_14935,N_15040);
or U16693 (N_16693,N_14709,N_15568);
nand U16694 (N_16694,N_14308,N_15214);
nor U16695 (N_16695,N_15053,N_14331);
or U16696 (N_16696,N_15069,N_14165);
xor U16697 (N_16697,N_15926,N_14329);
xor U16698 (N_16698,N_15189,N_15825);
and U16699 (N_16699,N_14242,N_15334);
nand U16700 (N_16700,N_14516,N_15877);
xnor U16701 (N_16701,N_15744,N_15385);
xor U16702 (N_16702,N_14132,N_14043);
and U16703 (N_16703,N_14923,N_14952);
nand U16704 (N_16704,N_14708,N_15792);
or U16705 (N_16705,N_14975,N_15659);
and U16706 (N_16706,N_15422,N_14460);
or U16707 (N_16707,N_14115,N_15088);
nand U16708 (N_16708,N_14547,N_14020);
and U16709 (N_16709,N_15010,N_15454);
xor U16710 (N_16710,N_14828,N_15380);
or U16711 (N_16711,N_15555,N_14622);
nand U16712 (N_16712,N_14438,N_15246);
xnor U16713 (N_16713,N_15432,N_14140);
nor U16714 (N_16714,N_15055,N_14186);
or U16715 (N_16715,N_14482,N_15800);
and U16716 (N_16716,N_14161,N_15866);
xor U16717 (N_16717,N_15310,N_14874);
nor U16718 (N_16718,N_15741,N_15719);
or U16719 (N_16719,N_15791,N_14475);
nor U16720 (N_16720,N_14253,N_15678);
xnor U16721 (N_16721,N_14395,N_15927);
or U16722 (N_16722,N_14834,N_15795);
nor U16723 (N_16723,N_15930,N_14758);
and U16724 (N_16724,N_14633,N_14119);
xnor U16725 (N_16725,N_15688,N_15150);
nand U16726 (N_16726,N_14467,N_15369);
and U16727 (N_16727,N_15248,N_14425);
xnor U16728 (N_16728,N_14314,N_15782);
nor U16729 (N_16729,N_15284,N_15836);
and U16730 (N_16730,N_14417,N_15819);
xnor U16731 (N_16731,N_15510,N_14900);
or U16732 (N_16732,N_15315,N_15728);
and U16733 (N_16733,N_15987,N_15045);
xnor U16734 (N_16734,N_14225,N_15704);
nand U16735 (N_16735,N_15260,N_15216);
nand U16736 (N_16736,N_14211,N_14435);
nand U16737 (N_16737,N_14757,N_15990);
or U16738 (N_16738,N_14512,N_14854);
xnor U16739 (N_16739,N_15046,N_14942);
and U16740 (N_16740,N_14458,N_14248);
and U16741 (N_16741,N_15487,N_15404);
nor U16742 (N_16742,N_15473,N_15140);
nor U16743 (N_16743,N_14915,N_14673);
and U16744 (N_16744,N_15006,N_14226);
nor U16745 (N_16745,N_14762,N_15749);
or U16746 (N_16746,N_15374,N_15827);
nor U16747 (N_16747,N_14749,N_14821);
nor U16748 (N_16748,N_14318,N_15210);
or U16749 (N_16749,N_15769,N_15054);
nand U16750 (N_16750,N_14861,N_14987);
and U16751 (N_16751,N_15540,N_14172);
nand U16752 (N_16752,N_14076,N_15705);
or U16753 (N_16753,N_15916,N_15395);
xnor U16754 (N_16754,N_15458,N_14258);
or U16755 (N_16755,N_14164,N_15600);
xor U16756 (N_16756,N_15724,N_15887);
and U16757 (N_16757,N_14267,N_14410);
and U16758 (N_16758,N_14282,N_15777);
or U16759 (N_16759,N_15668,N_15613);
nand U16760 (N_16760,N_14985,N_15136);
nor U16761 (N_16761,N_15730,N_14752);
nand U16762 (N_16762,N_14080,N_14181);
nand U16763 (N_16763,N_15317,N_14118);
nand U16764 (N_16764,N_15130,N_14858);
and U16765 (N_16765,N_14896,N_14477);
or U16766 (N_16766,N_15853,N_15628);
xnor U16767 (N_16767,N_14156,N_14408);
xnor U16768 (N_16768,N_15234,N_15835);
nor U16769 (N_16769,N_15925,N_15299);
and U16770 (N_16770,N_15514,N_15762);
nor U16771 (N_16771,N_15847,N_14576);
xor U16772 (N_16772,N_14689,N_15290);
xor U16773 (N_16773,N_14412,N_15059);
nand U16774 (N_16774,N_15340,N_14254);
nand U16775 (N_16775,N_14217,N_14931);
nand U16776 (N_16776,N_15492,N_14584);
and U16777 (N_16777,N_15051,N_14063);
nand U16778 (N_16778,N_14231,N_14652);
or U16779 (N_16779,N_14183,N_14930);
nand U16780 (N_16780,N_15047,N_14730);
or U16781 (N_16781,N_15331,N_14209);
nor U16782 (N_16782,N_14035,N_15032);
nor U16783 (N_16783,N_14478,N_14404);
and U16784 (N_16784,N_15997,N_14064);
or U16785 (N_16785,N_14860,N_15832);
nor U16786 (N_16786,N_14442,N_14141);
nor U16787 (N_16787,N_15298,N_14182);
nor U16788 (N_16788,N_15061,N_14718);
xnor U16789 (N_16789,N_15503,N_15708);
and U16790 (N_16790,N_14202,N_14383);
xor U16791 (N_16791,N_15348,N_15533);
and U16792 (N_16792,N_14259,N_15520);
or U16793 (N_16793,N_15882,N_14324);
and U16794 (N_16794,N_15226,N_15683);
nor U16795 (N_16795,N_15405,N_15839);
xnor U16796 (N_16796,N_14302,N_15544);
and U16797 (N_16797,N_14067,N_14737);
nor U16798 (N_16798,N_14669,N_15005);
or U16799 (N_16799,N_14197,N_15733);
or U16800 (N_16800,N_14658,N_14542);
nor U16801 (N_16801,N_15760,N_15251);
xnor U16802 (N_16802,N_14499,N_15804);
xnor U16803 (N_16803,N_14649,N_14657);
xnor U16804 (N_16804,N_15617,N_15821);
nand U16805 (N_16805,N_14541,N_15075);
and U16806 (N_16806,N_15085,N_14474);
nand U16807 (N_16807,N_14337,N_15765);
nand U16808 (N_16808,N_15050,N_14422);
nand U16809 (N_16809,N_14693,N_15687);
nor U16810 (N_16810,N_15633,N_14518);
or U16811 (N_16811,N_15516,N_14925);
nor U16812 (N_16812,N_14640,N_15801);
xnor U16813 (N_16813,N_14381,N_14082);
and U16814 (N_16814,N_15787,N_14655);
and U16815 (N_16815,N_14886,N_15575);
or U16816 (N_16816,N_15430,N_14921);
nor U16817 (N_16817,N_14237,N_14729);
and U16818 (N_16818,N_14265,N_15431);
nor U16819 (N_16819,N_15375,N_14849);
or U16820 (N_16820,N_14934,N_15200);
and U16821 (N_16821,N_14180,N_14015);
nor U16822 (N_16822,N_14587,N_15845);
nand U16823 (N_16823,N_15996,N_14393);
and U16824 (N_16824,N_15307,N_14926);
and U16825 (N_16825,N_14487,N_15598);
nor U16826 (N_16826,N_14341,N_14372);
nor U16827 (N_16827,N_14522,N_14783);
nand U16828 (N_16828,N_15599,N_15721);
xor U16829 (N_16829,N_14698,N_15703);
xnor U16830 (N_16830,N_15556,N_14270);
nor U16831 (N_16831,N_15498,N_14130);
nand U16832 (N_16832,N_14480,N_14493);
xor U16833 (N_16833,N_15476,N_14965);
and U16834 (N_16834,N_14212,N_15890);
or U16835 (N_16835,N_15443,N_14801);
xor U16836 (N_16836,N_15504,N_15838);
xnor U16837 (N_16837,N_14537,N_14147);
xnor U16838 (N_16838,N_14426,N_14483);
and U16839 (N_16839,N_14996,N_14163);
nand U16840 (N_16840,N_15960,N_15604);
nand U16841 (N_16841,N_14213,N_14981);
and U16842 (N_16842,N_15029,N_15268);
nand U16843 (N_16843,N_14187,N_15641);
xnor U16844 (N_16844,N_14192,N_14560);
xnor U16845 (N_16845,N_14790,N_14077);
or U16846 (N_16846,N_15660,N_15933);
nor U16847 (N_16847,N_14550,N_15305);
nand U16848 (N_16848,N_15132,N_14643);
and U16849 (N_16849,N_15207,N_15967);
xor U16850 (N_16850,N_15386,N_15196);
xor U16851 (N_16851,N_15699,N_15810);
or U16852 (N_16852,N_15077,N_15807);
nor U16853 (N_16853,N_14510,N_15208);
nor U16854 (N_16854,N_15421,N_15626);
and U16855 (N_16855,N_14948,N_14890);
or U16856 (N_16856,N_14616,N_15670);
xor U16857 (N_16857,N_14664,N_15178);
nor U16858 (N_16858,N_14012,N_14920);
nor U16859 (N_16859,N_14676,N_15358);
or U16860 (N_16860,N_15271,N_15667);
nor U16861 (N_16861,N_14332,N_15561);
and U16862 (N_16862,N_14280,N_14041);
and U16863 (N_16863,N_15523,N_15064);
or U16864 (N_16864,N_15684,N_15943);
xnor U16865 (N_16865,N_15873,N_15793);
or U16866 (N_16866,N_14074,N_14096);
and U16867 (N_16867,N_15570,N_15709);
xor U16868 (N_16868,N_15288,N_15619);
nor U16869 (N_16869,N_14960,N_15689);
and U16870 (N_16870,N_15048,N_14818);
or U16871 (N_16871,N_15511,N_14774);
nor U16872 (N_16872,N_14105,N_14906);
and U16873 (N_16873,N_15301,N_15856);
and U16874 (N_16874,N_14278,N_15151);
nand U16875 (N_16875,N_15971,N_15147);
nand U16876 (N_16876,N_15862,N_15030);
nor U16877 (N_16877,N_14720,N_15731);
or U16878 (N_16878,N_14184,N_15182);
xnor U16879 (N_16879,N_14473,N_15367);
nand U16880 (N_16880,N_14386,N_15438);
and U16881 (N_16881,N_14724,N_15642);
and U16882 (N_16882,N_14177,N_14690);
or U16883 (N_16883,N_14023,N_14416);
or U16884 (N_16884,N_14929,N_14108);
xnor U16885 (N_16885,N_15732,N_15445);
and U16886 (N_16886,N_15918,N_15779);
xor U16887 (N_16887,N_15202,N_14590);
and U16888 (N_16888,N_15160,N_15223);
nand U16889 (N_16889,N_15353,N_15993);
and U16890 (N_16890,N_14323,N_15442);
nand U16891 (N_16891,N_14103,N_15145);
and U16892 (N_16892,N_14068,N_15266);
xnor U16893 (N_16893,N_15798,N_14235);
nor U16894 (N_16894,N_14820,N_15947);
nand U16895 (N_16895,N_14485,N_14786);
or U16896 (N_16896,N_14879,N_15815);
and U16897 (N_16897,N_15412,N_15535);
nor U16898 (N_16898,N_14379,N_15609);
and U16899 (N_16899,N_15474,N_15239);
nor U16900 (N_16900,N_14653,N_15939);
nand U16901 (N_16901,N_14218,N_14450);
or U16902 (N_16902,N_14503,N_14178);
nand U16903 (N_16903,N_14238,N_14968);
xnor U16904 (N_16904,N_14656,N_15994);
nor U16905 (N_16905,N_14312,N_14454);
nand U16906 (N_16906,N_14606,N_15988);
and U16907 (N_16907,N_15398,N_14400);
or U16908 (N_16908,N_15446,N_14558);
and U16909 (N_16909,N_14572,N_15611);
or U16910 (N_16910,N_15679,N_14999);
nor U16911 (N_16911,N_15701,N_14717);
nor U16912 (N_16912,N_14605,N_14862);
xor U16913 (N_16913,N_14360,N_14078);
nor U16914 (N_16914,N_15861,N_15058);
nand U16915 (N_16915,N_15694,N_14523);
xnor U16916 (N_16916,N_15179,N_15243);
and U16917 (N_16917,N_14065,N_14349);
or U16918 (N_16918,N_14092,N_15621);
nand U16919 (N_16919,N_14723,N_14980);
and U16920 (N_16920,N_14228,N_15195);
nand U16921 (N_16921,N_15753,N_14918);
xor U16922 (N_16922,N_14097,N_15961);
and U16923 (N_16923,N_15308,N_15148);
or U16924 (N_16924,N_14292,N_14005);
nor U16925 (N_16925,N_14734,N_15338);
nand U16926 (N_16926,N_15134,N_15881);
or U16927 (N_16927,N_15909,N_14647);
nand U16928 (N_16928,N_15371,N_15154);
xnor U16929 (N_16929,N_15538,N_15283);
nor U16930 (N_16930,N_15658,N_14997);
xor U16931 (N_16931,N_15582,N_14614);
xor U16932 (N_16932,N_15944,N_14962);
xnor U16933 (N_16933,N_14791,N_14967);
and U16934 (N_16934,N_14390,N_15263);
and U16935 (N_16935,N_15319,N_14449);
nor U16936 (N_16936,N_15090,N_15797);
nor U16937 (N_16937,N_15218,N_14574);
nand U16938 (N_16938,N_14045,N_15316);
and U16939 (N_16939,N_14949,N_15675);
or U16940 (N_16940,N_15537,N_15387);
or U16941 (N_16941,N_14811,N_15802);
and U16942 (N_16942,N_15478,N_15164);
or U16943 (N_16943,N_15726,N_14098);
nor U16944 (N_16944,N_15370,N_15936);
or U16945 (N_16945,N_15627,N_15965);
nor U16946 (N_16946,N_14391,N_15671);
nand U16947 (N_16947,N_14452,N_15113);
and U16948 (N_16948,N_15114,N_14054);
nor U16949 (N_16949,N_15885,N_14741);
and U16950 (N_16950,N_14807,N_15060);
or U16951 (N_16951,N_14813,N_14794);
xor U16952 (N_16952,N_14286,N_14039);
or U16953 (N_16953,N_14430,N_15649);
xnor U16954 (N_16954,N_15886,N_14580);
xor U16955 (N_16955,N_15532,N_15775);
and U16956 (N_16956,N_15152,N_15184);
xnor U16957 (N_16957,N_15583,N_15359);
and U16958 (N_16958,N_14234,N_14707);
nor U16959 (N_16959,N_14315,N_15494);
nor U16960 (N_16960,N_14227,N_15464);
xnor U16961 (N_16961,N_15608,N_15693);
nand U16962 (N_16962,N_15254,N_15330);
nand U16963 (N_16963,N_14611,N_14205);
xnor U16964 (N_16964,N_15084,N_15903);
nand U16965 (N_16965,N_14911,N_14465);
nor U16966 (N_16966,N_14500,N_15181);
nand U16967 (N_16967,N_15146,N_15174);
xnor U16968 (N_16968,N_14579,N_14908);
or U16969 (N_16969,N_14988,N_15673);
xnor U16970 (N_16970,N_15082,N_15534);
nor U16971 (N_16971,N_15337,N_14415);
and U16972 (N_16972,N_14763,N_14621);
or U16973 (N_16973,N_15142,N_14060);
xor U16974 (N_16974,N_15915,N_15834);
xor U16975 (N_16975,N_15119,N_14771);
or U16976 (N_16976,N_14083,N_15929);
nand U16977 (N_16977,N_14504,N_14037);
and U16978 (N_16978,N_15424,N_14420);
xor U16979 (N_16979,N_14007,N_14044);
nand U16980 (N_16980,N_14725,N_14787);
or U16981 (N_16981,N_15935,N_15275);
and U16982 (N_16982,N_15581,N_14895);
and U16983 (N_16983,N_15955,N_14727);
nand U16984 (N_16984,N_14702,N_15567);
and U16985 (N_16985,N_15087,N_14869);
or U16986 (N_16986,N_14733,N_14565);
or U16987 (N_16987,N_14307,N_14539);
xnor U16988 (N_16988,N_15874,N_15736);
and U16989 (N_16989,N_15419,N_15383);
and U16990 (N_16990,N_15823,N_14034);
nand U16991 (N_16991,N_15636,N_14497);
nor U16992 (N_16992,N_14810,N_14057);
nand U16993 (N_16993,N_15245,N_14157);
nor U16994 (N_16994,N_14883,N_15471);
nand U16995 (N_16995,N_15293,N_14754);
or U16996 (N_16996,N_14457,N_14617);
or U16997 (N_16997,N_14696,N_14800);
xor U16998 (N_16998,N_15139,N_15813);
and U16999 (N_16999,N_15411,N_14958);
nor U17000 (N_17000,N_14706,N_14666);
xor U17001 (N_17001,N_14331,N_14193);
or U17002 (N_17002,N_14292,N_14356);
xnor U17003 (N_17003,N_14378,N_15591);
xor U17004 (N_17004,N_14440,N_14441);
xnor U17005 (N_17005,N_14932,N_15541);
xor U17006 (N_17006,N_15688,N_14158);
and U17007 (N_17007,N_14917,N_14316);
nor U17008 (N_17008,N_14384,N_15961);
or U17009 (N_17009,N_14054,N_15127);
and U17010 (N_17010,N_14080,N_15328);
and U17011 (N_17011,N_15599,N_15173);
xnor U17012 (N_17012,N_15078,N_15774);
or U17013 (N_17013,N_15064,N_14394);
and U17014 (N_17014,N_14999,N_14245);
xor U17015 (N_17015,N_14299,N_14337);
and U17016 (N_17016,N_15133,N_15653);
nor U17017 (N_17017,N_14522,N_15570);
xor U17018 (N_17018,N_14759,N_14875);
or U17019 (N_17019,N_14869,N_14525);
and U17020 (N_17020,N_15769,N_15196);
and U17021 (N_17021,N_14560,N_15493);
nand U17022 (N_17022,N_14782,N_15096);
or U17023 (N_17023,N_15015,N_14586);
and U17024 (N_17024,N_14967,N_15361);
and U17025 (N_17025,N_14092,N_14806);
nand U17026 (N_17026,N_15960,N_14029);
or U17027 (N_17027,N_15944,N_15735);
nand U17028 (N_17028,N_15383,N_14357);
and U17029 (N_17029,N_15024,N_14780);
xnor U17030 (N_17030,N_15611,N_15031);
and U17031 (N_17031,N_14080,N_15837);
xnor U17032 (N_17032,N_15862,N_14983);
xnor U17033 (N_17033,N_15365,N_14595);
and U17034 (N_17034,N_15817,N_15212);
or U17035 (N_17035,N_15168,N_15989);
nor U17036 (N_17036,N_15569,N_14620);
nand U17037 (N_17037,N_15874,N_14214);
xnor U17038 (N_17038,N_15370,N_15978);
or U17039 (N_17039,N_14750,N_14910);
nand U17040 (N_17040,N_15323,N_15027);
and U17041 (N_17041,N_15896,N_14947);
and U17042 (N_17042,N_14953,N_14709);
nand U17043 (N_17043,N_14780,N_14609);
or U17044 (N_17044,N_15007,N_15795);
xor U17045 (N_17045,N_15214,N_14094);
nand U17046 (N_17046,N_14518,N_15454);
nor U17047 (N_17047,N_14938,N_15779);
nor U17048 (N_17048,N_14525,N_15614);
and U17049 (N_17049,N_14356,N_15005);
nand U17050 (N_17050,N_14210,N_14178);
and U17051 (N_17051,N_14207,N_14457);
nand U17052 (N_17052,N_15785,N_15385);
xnor U17053 (N_17053,N_14315,N_14133);
xnor U17054 (N_17054,N_14940,N_15701);
and U17055 (N_17055,N_14834,N_15806);
and U17056 (N_17056,N_14275,N_14546);
and U17057 (N_17057,N_14435,N_15129);
nor U17058 (N_17058,N_15604,N_15526);
xor U17059 (N_17059,N_14388,N_14791);
xor U17060 (N_17060,N_15697,N_15786);
nand U17061 (N_17061,N_15144,N_14282);
or U17062 (N_17062,N_14670,N_14103);
and U17063 (N_17063,N_15776,N_15061);
and U17064 (N_17064,N_15513,N_15490);
or U17065 (N_17065,N_14324,N_14463);
and U17066 (N_17066,N_15262,N_15912);
xor U17067 (N_17067,N_15897,N_14474);
or U17068 (N_17068,N_14158,N_14949);
and U17069 (N_17069,N_14948,N_14074);
xnor U17070 (N_17070,N_15881,N_14125);
nand U17071 (N_17071,N_15925,N_15491);
or U17072 (N_17072,N_14622,N_15166);
or U17073 (N_17073,N_15902,N_14995);
nor U17074 (N_17074,N_14267,N_15577);
nand U17075 (N_17075,N_14829,N_14108);
nand U17076 (N_17076,N_14487,N_15059);
or U17077 (N_17077,N_15109,N_15055);
nand U17078 (N_17078,N_14259,N_14146);
nor U17079 (N_17079,N_14240,N_15582);
xnor U17080 (N_17080,N_14234,N_15014);
and U17081 (N_17081,N_14572,N_15905);
and U17082 (N_17082,N_15192,N_14392);
and U17083 (N_17083,N_14621,N_15358);
nand U17084 (N_17084,N_15135,N_15466);
nand U17085 (N_17085,N_15175,N_15987);
xnor U17086 (N_17086,N_14520,N_15645);
xnor U17087 (N_17087,N_14877,N_15792);
or U17088 (N_17088,N_15487,N_14203);
or U17089 (N_17089,N_14917,N_15999);
or U17090 (N_17090,N_15398,N_14138);
and U17091 (N_17091,N_15707,N_15426);
xnor U17092 (N_17092,N_15565,N_15640);
xor U17093 (N_17093,N_14368,N_14744);
nor U17094 (N_17094,N_15589,N_15797);
xor U17095 (N_17095,N_15333,N_15012);
or U17096 (N_17096,N_14155,N_15372);
xnor U17097 (N_17097,N_14640,N_15260);
nand U17098 (N_17098,N_14331,N_15886);
nand U17099 (N_17099,N_14927,N_15732);
and U17100 (N_17100,N_15157,N_14198);
and U17101 (N_17101,N_15237,N_15325);
nor U17102 (N_17102,N_14024,N_15666);
or U17103 (N_17103,N_14952,N_15861);
nor U17104 (N_17104,N_14203,N_15231);
xor U17105 (N_17105,N_14531,N_14316);
nand U17106 (N_17106,N_15667,N_14970);
nand U17107 (N_17107,N_14253,N_14485);
nor U17108 (N_17108,N_15930,N_14026);
nor U17109 (N_17109,N_15807,N_15850);
nor U17110 (N_17110,N_14693,N_14947);
or U17111 (N_17111,N_15394,N_14616);
nand U17112 (N_17112,N_14756,N_14845);
or U17113 (N_17113,N_14373,N_14383);
xnor U17114 (N_17114,N_14226,N_14779);
nor U17115 (N_17115,N_15696,N_14862);
and U17116 (N_17116,N_15804,N_15186);
or U17117 (N_17117,N_15140,N_15978);
xnor U17118 (N_17118,N_14416,N_14626);
and U17119 (N_17119,N_14940,N_15777);
and U17120 (N_17120,N_15880,N_14389);
nand U17121 (N_17121,N_15134,N_15389);
xnor U17122 (N_17122,N_15173,N_15844);
and U17123 (N_17123,N_15336,N_14063);
nand U17124 (N_17124,N_14928,N_15046);
and U17125 (N_17125,N_15320,N_15612);
or U17126 (N_17126,N_15431,N_15347);
nor U17127 (N_17127,N_14767,N_15863);
nor U17128 (N_17128,N_14118,N_15924);
nor U17129 (N_17129,N_15020,N_15687);
nor U17130 (N_17130,N_14896,N_15845);
and U17131 (N_17131,N_15729,N_15016);
xnor U17132 (N_17132,N_14133,N_15305);
and U17133 (N_17133,N_14463,N_15148);
and U17134 (N_17134,N_14710,N_14022);
nor U17135 (N_17135,N_15230,N_15193);
nand U17136 (N_17136,N_14175,N_14540);
nor U17137 (N_17137,N_14974,N_14763);
and U17138 (N_17138,N_14903,N_14965);
and U17139 (N_17139,N_15349,N_14863);
xnor U17140 (N_17140,N_14571,N_14212);
xor U17141 (N_17141,N_15953,N_14549);
or U17142 (N_17142,N_15378,N_14834);
nand U17143 (N_17143,N_14888,N_14661);
or U17144 (N_17144,N_15835,N_14466);
xnor U17145 (N_17145,N_15995,N_15246);
xor U17146 (N_17146,N_14111,N_15393);
xnor U17147 (N_17147,N_15405,N_15824);
xnor U17148 (N_17148,N_15532,N_15618);
and U17149 (N_17149,N_15411,N_14174);
nand U17150 (N_17150,N_15410,N_15650);
xnor U17151 (N_17151,N_14790,N_14949);
and U17152 (N_17152,N_14147,N_15859);
and U17153 (N_17153,N_14501,N_14405);
and U17154 (N_17154,N_15347,N_15393);
or U17155 (N_17155,N_14049,N_14192);
xor U17156 (N_17156,N_14386,N_15947);
and U17157 (N_17157,N_15187,N_14727);
xnor U17158 (N_17158,N_15908,N_14189);
and U17159 (N_17159,N_15414,N_15907);
and U17160 (N_17160,N_14742,N_15114);
or U17161 (N_17161,N_14083,N_15707);
nand U17162 (N_17162,N_14587,N_15033);
nand U17163 (N_17163,N_15550,N_14811);
and U17164 (N_17164,N_15296,N_15275);
and U17165 (N_17165,N_14788,N_14013);
and U17166 (N_17166,N_15531,N_14670);
or U17167 (N_17167,N_14269,N_15340);
or U17168 (N_17168,N_15366,N_15939);
or U17169 (N_17169,N_15523,N_15011);
nand U17170 (N_17170,N_14212,N_15628);
and U17171 (N_17171,N_14008,N_15562);
nor U17172 (N_17172,N_14499,N_14939);
or U17173 (N_17173,N_14432,N_14781);
xnor U17174 (N_17174,N_14389,N_15901);
and U17175 (N_17175,N_14344,N_15469);
and U17176 (N_17176,N_15711,N_15999);
xnor U17177 (N_17177,N_15257,N_14690);
nand U17178 (N_17178,N_15138,N_15903);
xnor U17179 (N_17179,N_15923,N_15884);
xor U17180 (N_17180,N_15665,N_15318);
nand U17181 (N_17181,N_14986,N_15194);
and U17182 (N_17182,N_15135,N_14020);
and U17183 (N_17183,N_15106,N_14349);
or U17184 (N_17184,N_14974,N_15998);
nor U17185 (N_17185,N_15840,N_15251);
xnor U17186 (N_17186,N_15200,N_15769);
nor U17187 (N_17187,N_14204,N_15601);
and U17188 (N_17188,N_14607,N_14541);
xnor U17189 (N_17189,N_14914,N_15987);
or U17190 (N_17190,N_14487,N_15912);
or U17191 (N_17191,N_15209,N_14740);
or U17192 (N_17192,N_15786,N_14687);
nand U17193 (N_17193,N_14766,N_15288);
and U17194 (N_17194,N_14162,N_14138);
and U17195 (N_17195,N_14436,N_14312);
nand U17196 (N_17196,N_14903,N_14435);
or U17197 (N_17197,N_14554,N_14129);
and U17198 (N_17198,N_14688,N_14886);
nand U17199 (N_17199,N_14599,N_15807);
nand U17200 (N_17200,N_14591,N_14338);
nor U17201 (N_17201,N_15930,N_15264);
and U17202 (N_17202,N_14917,N_14382);
nand U17203 (N_17203,N_15044,N_14203);
nand U17204 (N_17204,N_15811,N_15283);
xnor U17205 (N_17205,N_15201,N_15345);
nand U17206 (N_17206,N_14776,N_15528);
and U17207 (N_17207,N_15424,N_14270);
nand U17208 (N_17208,N_15621,N_15782);
nand U17209 (N_17209,N_15038,N_15629);
and U17210 (N_17210,N_14183,N_15611);
and U17211 (N_17211,N_15813,N_14014);
and U17212 (N_17212,N_15560,N_15929);
nor U17213 (N_17213,N_15670,N_15302);
and U17214 (N_17214,N_15995,N_15844);
xor U17215 (N_17215,N_15227,N_14587);
nand U17216 (N_17216,N_14469,N_15218);
nand U17217 (N_17217,N_15105,N_14517);
or U17218 (N_17218,N_15373,N_14408);
or U17219 (N_17219,N_14735,N_15916);
nor U17220 (N_17220,N_14282,N_15378);
xnor U17221 (N_17221,N_15834,N_14848);
and U17222 (N_17222,N_15079,N_15048);
nor U17223 (N_17223,N_15125,N_15054);
nand U17224 (N_17224,N_15516,N_14689);
nand U17225 (N_17225,N_15687,N_14641);
nand U17226 (N_17226,N_14728,N_15513);
nor U17227 (N_17227,N_15063,N_14111);
or U17228 (N_17228,N_15755,N_14148);
and U17229 (N_17229,N_15677,N_15588);
nand U17230 (N_17230,N_15468,N_14471);
nand U17231 (N_17231,N_14684,N_14139);
nor U17232 (N_17232,N_15649,N_14014);
nor U17233 (N_17233,N_14053,N_14040);
or U17234 (N_17234,N_15025,N_15951);
and U17235 (N_17235,N_15578,N_15859);
and U17236 (N_17236,N_15669,N_15876);
and U17237 (N_17237,N_15217,N_15997);
xnor U17238 (N_17238,N_14066,N_15296);
nand U17239 (N_17239,N_15356,N_15273);
and U17240 (N_17240,N_15642,N_15137);
nor U17241 (N_17241,N_14829,N_15649);
or U17242 (N_17242,N_15009,N_14628);
or U17243 (N_17243,N_15354,N_14711);
xnor U17244 (N_17244,N_14018,N_14407);
or U17245 (N_17245,N_15948,N_14493);
or U17246 (N_17246,N_15864,N_15127);
nand U17247 (N_17247,N_14331,N_14837);
nand U17248 (N_17248,N_14219,N_14287);
or U17249 (N_17249,N_15807,N_15558);
xnor U17250 (N_17250,N_15914,N_14852);
xnor U17251 (N_17251,N_14192,N_15963);
xor U17252 (N_17252,N_14667,N_15819);
and U17253 (N_17253,N_14643,N_15842);
or U17254 (N_17254,N_14434,N_15106);
nand U17255 (N_17255,N_14206,N_15262);
nor U17256 (N_17256,N_14691,N_15610);
or U17257 (N_17257,N_14996,N_14528);
xor U17258 (N_17258,N_15996,N_15506);
or U17259 (N_17259,N_14873,N_14804);
xnor U17260 (N_17260,N_15110,N_15694);
nand U17261 (N_17261,N_15606,N_14437);
or U17262 (N_17262,N_15213,N_14125);
or U17263 (N_17263,N_15733,N_15336);
or U17264 (N_17264,N_14301,N_14078);
xnor U17265 (N_17265,N_15326,N_14995);
nand U17266 (N_17266,N_15881,N_14304);
xnor U17267 (N_17267,N_15575,N_14313);
xor U17268 (N_17268,N_14750,N_14635);
or U17269 (N_17269,N_15998,N_15669);
xor U17270 (N_17270,N_14334,N_14225);
nand U17271 (N_17271,N_14030,N_15645);
xor U17272 (N_17272,N_14609,N_14579);
and U17273 (N_17273,N_14314,N_15090);
nor U17274 (N_17274,N_14360,N_14813);
nor U17275 (N_17275,N_15647,N_14910);
and U17276 (N_17276,N_15496,N_15528);
or U17277 (N_17277,N_14430,N_14509);
and U17278 (N_17278,N_14892,N_15880);
nand U17279 (N_17279,N_14463,N_15533);
nand U17280 (N_17280,N_15905,N_15885);
nor U17281 (N_17281,N_15088,N_15184);
and U17282 (N_17282,N_14095,N_14701);
xnor U17283 (N_17283,N_14560,N_14317);
xor U17284 (N_17284,N_15709,N_15035);
and U17285 (N_17285,N_15794,N_14378);
nand U17286 (N_17286,N_14382,N_14393);
xnor U17287 (N_17287,N_15852,N_15065);
nand U17288 (N_17288,N_15327,N_15453);
and U17289 (N_17289,N_15802,N_15883);
or U17290 (N_17290,N_15972,N_15174);
nor U17291 (N_17291,N_14977,N_15180);
nand U17292 (N_17292,N_15866,N_14298);
xnor U17293 (N_17293,N_14079,N_14075);
nand U17294 (N_17294,N_15623,N_14516);
xor U17295 (N_17295,N_15445,N_15398);
nand U17296 (N_17296,N_14950,N_15697);
and U17297 (N_17297,N_14320,N_15046);
and U17298 (N_17298,N_15494,N_15749);
or U17299 (N_17299,N_15582,N_14700);
and U17300 (N_17300,N_14869,N_14634);
or U17301 (N_17301,N_14382,N_15863);
nor U17302 (N_17302,N_14701,N_15386);
nor U17303 (N_17303,N_14789,N_14206);
nand U17304 (N_17304,N_14267,N_15144);
and U17305 (N_17305,N_15214,N_15866);
nand U17306 (N_17306,N_15649,N_15564);
or U17307 (N_17307,N_14670,N_15255);
and U17308 (N_17308,N_14440,N_14331);
nand U17309 (N_17309,N_15374,N_14280);
nor U17310 (N_17310,N_14275,N_15279);
nor U17311 (N_17311,N_14931,N_14301);
xor U17312 (N_17312,N_14480,N_14380);
nand U17313 (N_17313,N_15039,N_15352);
and U17314 (N_17314,N_14715,N_15757);
xnor U17315 (N_17315,N_15444,N_14489);
or U17316 (N_17316,N_14271,N_14293);
or U17317 (N_17317,N_14656,N_14621);
xor U17318 (N_17318,N_15646,N_14994);
and U17319 (N_17319,N_15244,N_15383);
or U17320 (N_17320,N_14247,N_15333);
and U17321 (N_17321,N_15959,N_14919);
xor U17322 (N_17322,N_15781,N_14207);
or U17323 (N_17323,N_14333,N_15838);
or U17324 (N_17324,N_15181,N_15484);
xor U17325 (N_17325,N_15211,N_14715);
xor U17326 (N_17326,N_15556,N_14188);
and U17327 (N_17327,N_15311,N_14293);
or U17328 (N_17328,N_15878,N_15643);
and U17329 (N_17329,N_15710,N_15900);
and U17330 (N_17330,N_14669,N_14274);
nand U17331 (N_17331,N_15838,N_14592);
xnor U17332 (N_17332,N_15171,N_15268);
nand U17333 (N_17333,N_15091,N_14291);
or U17334 (N_17334,N_15238,N_15630);
nor U17335 (N_17335,N_14534,N_15304);
or U17336 (N_17336,N_15853,N_14035);
or U17337 (N_17337,N_15356,N_15155);
xnor U17338 (N_17338,N_14636,N_15378);
and U17339 (N_17339,N_15804,N_14192);
nand U17340 (N_17340,N_14157,N_15595);
nor U17341 (N_17341,N_14828,N_14730);
xnor U17342 (N_17342,N_14116,N_15570);
nor U17343 (N_17343,N_14917,N_14558);
nor U17344 (N_17344,N_14524,N_14435);
xor U17345 (N_17345,N_14456,N_15734);
xor U17346 (N_17346,N_15095,N_14660);
xnor U17347 (N_17347,N_14505,N_15499);
or U17348 (N_17348,N_14029,N_14856);
or U17349 (N_17349,N_15848,N_14963);
xor U17350 (N_17350,N_14357,N_15625);
or U17351 (N_17351,N_14446,N_14626);
xor U17352 (N_17352,N_15964,N_15745);
or U17353 (N_17353,N_15837,N_15467);
nand U17354 (N_17354,N_15604,N_15088);
xnor U17355 (N_17355,N_14276,N_14114);
or U17356 (N_17356,N_15067,N_14523);
nor U17357 (N_17357,N_15746,N_14310);
nor U17358 (N_17358,N_15376,N_14094);
and U17359 (N_17359,N_15312,N_14807);
nor U17360 (N_17360,N_15250,N_15307);
nand U17361 (N_17361,N_15706,N_14340);
xnor U17362 (N_17362,N_14467,N_14138);
and U17363 (N_17363,N_14681,N_14218);
nand U17364 (N_17364,N_15829,N_14426);
xor U17365 (N_17365,N_14080,N_15067);
nor U17366 (N_17366,N_15735,N_14861);
and U17367 (N_17367,N_14477,N_14472);
or U17368 (N_17368,N_15873,N_15913);
and U17369 (N_17369,N_14985,N_15889);
nor U17370 (N_17370,N_15478,N_14748);
xnor U17371 (N_17371,N_15764,N_14173);
or U17372 (N_17372,N_14153,N_15207);
nand U17373 (N_17373,N_14501,N_15476);
and U17374 (N_17374,N_14887,N_15619);
and U17375 (N_17375,N_14398,N_14083);
or U17376 (N_17376,N_15337,N_14314);
or U17377 (N_17377,N_15726,N_14436);
and U17378 (N_17378,N_14883,N_14773);
nor U17379 (N_17379,N_15917,N_15294);
xnor U17380 (N_17380,N_15436,N_15693);
or U17381 (N_17381,N_15019,N_14077);
and U17382 (N_17382,N_15885,N_14470);
or U17383 (N_17383,N_14645,N_14393);
nor U17384 (N_17384,N_14069,N_14869);
nor U17385 (N_17385,N_15276,N_15979);
and U17386 (N_17386,N_14870,N_15105);
xor U17387 (N_17387,N_15610,N_15991);
or U17388 (N_17388,N_15754,N_14027);
or U17389 (N_17389,N_14682,N_14268);
or U17390 (N_17390,N_14201,N_15110);
nand U17391 (N_17391,N_15787,N_14593);
xnor U17392 (N_17392,N_14710,N_15582);
nor U17393 (N_17393,N_15233,N_15099);
and U17394 (N_17394,N_14761,N_14973);
or U17395 (N_17395,N_14903,N_14262);
or U17396 (N_17396,N_15711,N_15785);
nand U17397 (N_17397,N_14414,N_15367);
xnor U17398 (N_17398,N_15484,N_15720);
and U17399 (N_17399,N_15157,N_14216);
nor U17400 (N_17400,N_14559,N_14810);
nand U17401 (N_17401,N_14987,N_15171);
xnor U17402 (N_17402,N_14675,N_15932);
nand U17403 (N_17403,N_14092,N_15096);
or U17404 (N_17404,N_15227,N_15404);
or U17405 (N_17405,N_14657,N_14584);
nand U17406 (N_17406,N_15670,N_14677);
nand U17407 (N_17407,N_15528,N_14572);
nor U17408 (N_17408,N_14880,N_15200);
xnor U17409 (N_17409,N_14396,N_15271);
and U17410 (N_17410,N_15012,N_14503);
and U17411 (N_17411,N_14550,N_14658);
nand U17412 (N_17412,N_14643,N_15537);
nand U17413 (N_17413,N_15127,N_15498);
nor U17414 (N_17414,N_15853,N_15827);
nor U17415 (N_17415,N_15683,N_14691);
nor U17416 (N_17416,N_14075,N_14209);
xnor U17417 (N_17417,N_14847,N_15330);
nand U17418 (N_17418,N_14855,N_14922);
or U17419 (N_17419,N_15014,N_15503);
and U17420 (N_17420,N_14306,N_15231);
nor U17421 (N_17421,N_14364,N_14159);
nand U17422 (N_17422,N_14265,N_14478);
xnor U17423 (N_17423,N_15637,N_15919);
nand U17424 (N_17424,N_15157,N_15959);
nand U17425 (N_17425,N_14643,N_15854);
xor U17426 (N_17426,N_15162,N_15361);
xnor U17427 (N_17427,N_14913,N_15426);
xor U17428 (N_17428,N_14620,N_14760);
xor U17429 (N_17429,N_14921,N_15305);
or U17430 (N_17430,N_14694,N_15203);
and U17431 (N_17431,N_14277,N_15900);
nor U17432 (N_17432,N_14695,N_14468);
nor U17433 (N_17433,N_14705,N_14159);
xor U17434 (N_17434,N_14789,N_15056);
nand U17435 (N_17435,N_14582,N_15038);
xnor U17436 (N_17436,N_14139,N_15509);
and U17437 (N_17437,N_15549,N_14207);
or U17438 (N_17438,N_14044,N_14119);
or U17439 (N_17439,N_15802,N_14324);
nand U17440 (N_17440,N_15402,N_14404);
xor U17441 (N_17441,N_14474,N_14311);
xor U17442 (N_17442,N_15437,N_15530);
nand U17443 (N_17443,N_14139,N_14177);
nor U17444 (N_17444,N_14681,N_14588);
nand U17445 (N_17445,N_14872,N_15043);
nand U17446 (N_17446,N_15465,N_15550);
or U17447 (N_17447,N_14393,N_15724);
nand U17448 (N_17448,N_14645,N_15226);
and U17449 (N_17449,N_14462,N_15702);
nand U17450 (N_17450,N_15122,N_15259);
or U17451 (N_17451,N_14133,N_15565);
or U17452 (N_17452,N_15249,N_14453);
xnor U17453 (N_17453,N_15053,N_15551);
nor U17454 (N_17454,N_15118,N_14265);
nor U17455 (N_17455,N_14799,N_15500);
nor U17456 (N_17456,N_15416,N_14612);
and U17457 (N_17457,N_14625,N_14120);
xor U17458 (N_17458,N_14420,N_14219);
nor U17459 (N_17459,N_15596,N_15221);
and U17460 (N_17460,N_14005,N_15052);
or U17461 (N_17461,N_14194,N_14509);
nor U17462 (N_17462,N_14194,N_15198);
xnor U17463 (N_17463,N_15738,N_14834);
xor U17464 (N_17464,N_14586,N_14229);
or U17465 (N_17465,N_15898,N_14588);
and U17466 (N_17466,N_15322,N_14050);
xor U17467 (N_17467,N_15845,N_14912);
nand U17468 (N_17468,N_15905,N_15446);
nand U17469 (N_17469,N_14717,N_14803);
or U17470 (N_17470,N_15716,N_15262);
and U17471 (N_17471,N_15599,N_14865);
xnor U17472 (N_17472,N_15946,N_15716);
nor U17473 (N_17473,N_14389,N_14941);
or U17474 (N_17474,N_14413,N_15278);
or U17475 (N_17475,N_15242,N_14000);
or U17476 (N_17476,N_15828,N_15695);
or U17477 (N_17477,N_15819,N_15462);
or U17478 (N_17478,N_15435,N_15352);
or U17479 (N_17479,N_15334,N_15204);
xnor U17480 (N_17480,N_15903,N_15104);
nor U17481 (N_17481,N_14984,N_15541);
or U17482 (N_17482,N_15680,N_14904);
xnor U17483 (N_17483,N_15561,N_14310);
or U17484 (N_17484,N_15164,N_15071);
xor U17485 (N_17485,N_14444,N_15059);
xnor U17486 (N_17486,N_14766,N_15443);
and U17487 (N_17487,N_15298,N_15707);
xor U17488 (N_17488,N_15501,N_15625);
nand U17489 (N_17489,N_14800,N_15073);
and U17490 (N_17490,N_15031,N_15927);
and U17491 (N_17491,N_14344,N_15215);
xor U17492 (N_17492,N_14092,N_15774);
nor U17493 (N_17493,N_15237,N_14735);
nor U17494 (N_17494,N_14927,N_15035);
nand U17495 (N_17495,N_15772,N_15860);
nand U17496 (N_17496,N_15135,N_15602);
and U17497 (N_17497,N_14754,N_14459);
nand U17498 (N_17498,N_14984,N_14526);
or U17499 (N_17499,N_15242,N_14697);
and U17500 (N_17500,N_14328,N_14578);
and U17501 (N_17501,N_15603,N_14902);
or U17502 (N_17502,N_14969,N_15105);
xnor U17503 (N_17503,N_14289,N_15831);
and U17504 (N_17504,N_14975,N_15661);
or U17505 (N_17505,N_14083,N_14476);
nand U17506 (N_17506,N_14715,N_15094);
xnor U17507 (N_17507,N_14981,N_14503);
xnor U17508 (N_17508,N_15993,N_15878);
or U17509 (N_17509,N_14634,N_14940);
and U17510 (N_17510,N_15134,N_14507);
or U17511 (N_17511,N_15910,N_15947);
nand U17512 (N_17512,N_15685,N_14549);
xor U17513 (N_17513,N_14806,N_14807);
nor U17514 (N_17514,N_14128,N_14665);
nor U17515 (N_17515,N_15205,N_15570);
and U17516 (N_17516,N_14436,N_14075);
nand U17517 (N_17517,N_15487,N_15477);
nand U17518 (N_17518,N_15270,N_15728);
and U17519 (N_17519,N_14222,N_15714);
nand U17520 (N_17520,N_14761,N_14448);
or U17521 (N_17521,N_15438,N_14639);
xor U17522 (N_17522,N_15384,N_15979);
nor U17523 (N_17523,N_15077,N_14945);
and U17524 (N_17524,N_15317,N_14011);
and U17525 (N_17525,N_15323,N_14591);
xnor U17526 (N_17526,N_15967,N_15128);
and U17527 (N_17527,N_14350,N_14477);
nor U17528 (N_17528,N_14549,N_15296);
and U17529 (N_17529,N_15855,N_14416);
nand U17530 (N_17530,N_14910,N_15092);
nor U17531 (N_17531,N_14460,N_15521);
or U17532 (N_17532,N_14304,N_14515);
and U17533 (N_17533,N_15098,N_14598);
and U17534 (N_17534,N_14624,N_14715);
or U17535 (N_17535,N_14620,N_14845);
nor U17536 (N_17536,N_14447,N_15183);
xnor U17537 (N_17537,N_14777,N_14736);
nor U17538 (N_17538,N_15270,N_14700);
and U17539 (N_17539,N_14769,N_15868);
nand U17540 (N_17540,N_14368,N_15740);
nor U17541 (N_17541,N_14027,N_15344);
nand U17542 (N_17542,N_14103,N_14198);
nor U17543 (N_17543,N_14282,N_14039);
xnor U17544 (N_17544,N_15808,N_14482);
nor U17545 (N_17545,N_14421,N_14471);
and U17546 (N_17546,N_14332,N_15864);
and U17547 (N_17547,N_14567,N_15657);
xor U17548 (N_17548,N_14963,N_14996);
nor U17549 (N_17549,N_15105,N_14705);
nor U17550 (N_17550,N_14852,N_15878);
xnor U17551 (N_17551,N_15387,N_15973);
nand U17552 (N_17552,N_14433,N_14410);
xor U17553 (N_17553,N_14977,N_14051);
nor U17554 (N_17554,N_14811,N_14689);
and U17555 (N_17555,N_14910,N_15643);
or U17556 (N_17556,N_14274,N_14754);
or U17557 (N_17557,N_15413,N_15319);
xnor U17558 (N_17558,N_15019,N_14605);
and U17559 (N_17559,N_14812,N_14568);
nor U17560 (N_17560,N_15377,N_14584);
or U17561 (N_17561,N_14766,N_14077);
xor U17562 (N_17562,N_15747,N_15922);
xor U17563 (N_17563,N_15944,N_14984);
xor U17564 (N_17564,N_15737,N_15111);
nor U17565 (N_17565,N_14345,N_14187);
and U17566 (N_17566,N_15897,N_15288);
nor U17567 (N_17567,N_15992,N_14646);
nand U17568 (N_17568,N_15076,N_15919);
xor U17569 (N_17569,N_15390,N_15623);
xnor U17570 (N_17570,N_15794,N_14593);
and U17571 (N_17571,N_15474,N_15199);
nand U17572 (N_17572,N_15896,N_14049);
nor U17573 (N_17573,N_14748,N_14249);
or U17574 (N_17574,N_15979,N_14134);
and U17575 (N_17575,N_14155,N_14471);
or U17576 (N_17576,N_15489,N_14865);
and U17577 (N_17577,N_15470,N_15713);
xnor U17578 (N_17578,N_15168,N_14195);
nand U17579 (N_17579,N_14908,N_15614);
nor U17580 (N_17580,N_14550,N_15841);
and U17581 (N_17581,N_15488,N_15481);
nand U17582 (N_17582,N_14087,N_15212);
nand U17583 (N_17583,N_15994,N_14226);
nand U17584 (N_17584,N_15026,N_14889);
xnor U17585 (N_17585,N_15902,N_14531);
nor U17586 (N_17586,N_14333,N_15038);
or U17587 (N_17587,N_14221,N_15741);
xor U17588 (N_17588,N_15409,N_14196);
or U17589 (N_17589,N_15426,N_14930);
nor U17590 (N_17590,N_15493,N_15176);
or U17591 (N_17591,N_15156,N_15136);
nor U17592 (N_17592,N_15657,N_15712);
xnor U17593 (N_17593,N_14703,N_14979);
nand U17594 (N_17594,N_15499,N_14575);
nand U17595 (N_17595,N_14198,N_14098);
nand U17596 (N_17596,N_14854,N_15357);
and U17597 (N_17597,N_15340,N_14076);
xnor U17598 (N_17598,N_14948,N_15972);
xor U17599 (N_17599,N_15884,N_14758);
xnor U17600 (N_17600,N_15781,N_14680);
nor U17601 (N_17601,N_15486,N_14943);
nand U17602 (N_17602,N_15651,N_15382);
and U17603 (N_17603,N_14830,N_15525);
or U17604 (N_17604,N_15203,N_14432);
xnor U17605 (N_17605,N_15469,N_14126);
nor U17606 (N_17606,N_15268,N_15674);
nor U17607 (N_17607,N_15474,N_14566);
xnor U17608 (N_17608,N_15813,N_14685);
nand U17609 (N_17609,N_15980,N_14173);
nor U17610 (N_17610,N_15079,N_15496);
nand U17611 (N_17611,N_14473,N_15727);
xnor U17612 (N_17612,N_15976,N_15131);
nand U17613 (N_17613,N_15493,N_15623);
xor U17614 (N_17614,N_14324,N_15790);
and U17615 (N_17615,N_14513,N_14548);
and U17616 (N_17616,N_15782,N_14860);
nand U17617 (N_17617,N_14116,N_15265);
or U17618 (N_17618,N_15901,N_15656);
nor U17619 (N_17619,N_15741,N_15314);
nor U17620 (N_17620,N_15390,N_14598);
or U17621 (N_17621,N_15899,N_15599);
xnor U17622 (N_17622,N_15483,N_14949);
or U17623 (N_17623,N_14917,N_15410);
or U17624 (N_17624,N_14021,N_15809);
or U17625 (N_17625,N_15484,N_14696);
nand U17626 (N_17626,N_14603,N_14032);
nand U17627 (N_17627,N_14514,N_14202);
nand U17628 (N_17628,N_14808,N_14655);
and U17629 (N_17629,N_15356,N_15347);
nand U17630 (N_17630,N_15907,N_15203);
xnor U17631 (N_17631,N_14956,N_15434);
nor U17632 (N_17632,N_14396,N_15282);
nor U17633 (N_17633,N_14602,N_14651);
xnor U17634 (N_17634,N_14642,N_15232);
or U17635 (N_17635,N_15232,N_15654);
and U17636 (N_17636,N_15008,N_14921);
xnor U17637 (N_17637,N_14985,N_15488);
nand U17638 (N_17638,N_15105,N_15300);
xor U17639 (N_17639,N_15786,N_15828);
nand U17640 (N_17640,N_14435,N_14443);
nor U17641 (N_17641,N_14046,N_15875);
nor U17642 (N_17642,N_14618,N_15597);
xnor U17643 (N_17643,N_15234,N_14992);
nand U17644 (N_17644,N_14388,N_14925);
or U17645 (N_17645,N_15785,N_15703);
nand U17646 (N_17646,N_14419,N_14502);
and U17647 (N_17647,N_15227,N_14363);
nor U17648 (N_17648,N_15436,N_14916);
nor U17649 (N_17649,N_14769,N_14411);
nor U17650 (N_17650,N_14788,N_15098);
or U17651 (N_17651,N_14813,N_15233);
nand U17652 (N_17652,N_14536,N_14818);
and U17653 (N_17653,N_15588,N_15218);
xnor U17654 (N_17654,N_14437,N_15496);
or U17655 (N_17655,N_14483,N_15434);
nor U17656 (N_17656,N_15151,N_15670);
and U17657 (N_17657,N_15534,N_14274);
nand U17658 (N_17658,N_15592,N_14989);
nor U17659 (N_17659,N_14525,N_14587);
or U17660 (N_17660,N_15948,N_15616);
nand U17661 (N_17661,N_15499,N_15491);
and U17662 (N_17662,N_15918,N_15968);
xnor U17663 (N_17663,N_14219,N_15550);
xnor U17664 (N_17664,N_14966,N_15407);
nor U17665 (N_17665,N_15868,N_15954);
and U17666 (N_17666,N_14576,N_15342);
nand U17667 (N_17667,N_15833,N_14602);
and U17668 (N_17668,N_15439,N_15706);
or U17669 (N_17669,N_15367,N_15066);
and U17670 (N_17670,N_14147,N_15447);
and U17671 (N_17671,N_14038,N_15900);
nand U17672 (N_17672,N_14777,N_14743);
or U17673 (N_17673,N_14072,N_15130);
or U17674 (N_17674,N_14245,N_14317);
xnor U17675 (N_17675,N_14115,N_15390);
nand U17676 (N_17676,N_14805,N_14429);
nor U17677 (N_17677,N_14098,N_14869);
and U17678 (N_17678,N_15919,N_14426);
xor U17679 (N_17679,N_15485,N_15799);
xor U17680 (N_17680,N_14535,N_14686);
nor U17681 (N_17681,N_14723,N_15957);
and U17682 (N_17682,N_14506,N_14378);
xor U17683 (N_17683,N_15876,N_14889);
xor U17684 (N_17684,N_15925,N_14668);
or U17685 (N_17685,N_15781,N_15039);
xor U17686 (N_17686,N_15713,N_14281);
nor U17687 (N_17687,N_14234,N_15812);
xor U17688 (N_17688,N_14463,N_15423);
or U17689 (N_17689,N_15733,N_14561);
nand U17690 (N_17690,N_15118,N_14569);
xnor U17691 (N_17691,N_14243,N_15664);
nand U17692 (N_17692,N_15085,N_14047);
nor U17693 (N_17693,N_14271,N_15746);
xor U17694 (N_17694,N_14195,N_15773);
nor U17695 (N_17695,N_14373,N_15338);
nand U17696 (N_17696,N_15664,N_14647);
or U17697 (N_17697,N_15524,N_14502);
or U17698 (N_17698,N_14839,N_14100);
nand U17699 (N_17699,N_15740,N_15571);
and U17700 (N_17700,N_14520,N_15841);
nor U17701 (N_17701,N_15705,N_15508);
nand U17702 (N_17702,N_14822,N_15403);
nand U17703 (N_17703,N_14931,N_14713);
or U17704 (N_17704,N_15425,N_15094);
or U17705 (N_17705,N_14853,N_14328);
nand U17706 (N_17706,N_14999,N_15276);
or U17707 (N_17707,N_14891,N_15097);
or U17708 (N_17708,N_15763,N_14554);
xnor U17709 (N_17709,N_14209,N_14585);
nand U17710 (N_17710,N_14090,N_14067);
or U17711 (N_17711,N_14116,N_15193);
nand U17712 (N_17712,N_15961,N_14885);
nor U17713 (N_17713,N_14521,N_15694);
xnor U17714 (N_17714,N_14993,N_15960);
xor U17715 (N_17715,N_15369,N_14497);
nand U17716 (N_17716,N_14493,N_15310);
nand U17717 (N_17717,N_14591,N_14984);
nand U17718 (N_17718,N_15325,N_14921);
or U17719 (N_17719,N_15447,N_14654);
nor U17720 (N_17720,N_14944,N_15948);
and U17721 (N_17721,N_15096,N_14845);
xor U17722 (N_17722,N_15018,N_15053);
nand U17723 (N_17723,N_15199,N_14346);
and U17724 (N_17724,N_15431,N_15195);
and U17725 (N_17725,N_15613,N_15169);
xnor U17726 (N_17726,N_14328,N_15265);
or U17727 (N_17727,N_14812,N_14417);
or U17728 (N_17728,N_15336,N_14473);
nand U17729 (N_17729,N_15034,N_14398);
nand U17730 (N_17730,N_14095,N_14112);
or U17731 (N_17731,N_15795,N_14773);
and U17732 (N_17732,N_14967,N_15193);
nand U17733 (N_17733,N_14173,N_14177);
xor U17734 (N_17734,N_14315,N_14786);
nand U17735 (N_17735,N_15426,N_14028);
and U17736 (N_17736,N_14242,N_15174);
xnor U17737 (N_17737,N_15865,N_15824);
xor U17738 (N_17738,N_14739,N_14346);
and U17739 (N_17739,N_15162,N_15063);
nor U17740 (N_17740,N_15121,N_14490);
xor U17741 (N_17741,N_15974,N_14225);
and U17742 (N_17742,N_14633,N_14970);
or U17743 (N_17743,N_15944,N_15388);
and U17744 (N_17744,N_15642,N_14046);
xnor U17745 (N_17745,N_15078,N_15711);
xor U17746 (N_17746,N_14127,N_14290);
or U17747 (N_17747,N_15790,N_15168);
nor U17748 (N_17748,N_15482,N_14864);
or U17749 (N_17749,N_15445,N_14155);
and U17750 (N_17750,N_14356,N_14611);
or U17751 (N_17751,N_14742,N_14251);
and U17752 (N_17752,N_15001,N_15173);
xnor U17753 (N_17753,N_15551,N_15279);
nor U17754 (N_17754,N_14755,N_14017);
xnor U17755 (N_17755,N_15308,N_14257);
nor U17756 (N_17756,N_15872,N_14855);
nand U17757 (N_17757,N_14330,N_15141);
nand U17758 (N_17758,N_15609,N_15222);
nand U17759 (N_17759,N_15288,N_15051);
or U17760 (N_17760,N_14632,N_15752);
or U17761 (N_17761,N_15211,N_14944);
nor U17762 (N_17762,N_15476,N_14066);
or U17763 (N_17763,N_14773,N_14373);
and U17764 (N_17764,N_15880,N_15136);
nand U17765 (N_17765,N_15156,N_14763);
xnor U17766 (N_17766,N_15689,N_15265);
xnor U17767 (N_17767,N_15758,N_14386);
nor U17768 (N_17768,N_15428,N_14925);
nand U17769 (N_17769,N_15662,N_14056);
nor U17770 (N_17770,N_15746,N_15403);
nor U17771 (N_17771,N_14179,N_15618);
or U17772 (N_17772,N_15054,N_15536);
xor U17773 (N_17773,N_14126,N_14903);
nand U17774 (N_17774,N_15766,N_14314);
xnor U17775 (N_17775,N_14613,N_15380);
or U17776 (N_17776,N_14093,N_14880);
or U17777 (N_17777,N_15464,N_14018);
nor U17778 (N_17778,N_15659,N_15855);
xnor U17779 (N_17779,N_15192,N_15961);
nor U17780 (N_17780,N_15718,N_15407);
and U17781 (N_17781,N_14692,N_14037);
or U17782 (N_17782,N_14319,N_14953);
nand U17783 (N_17783,N_15469,N_15705);
nand U17784 (N_17784,N_14369,N_15329);
xnor U17785 (N_17785,N_14895,N_14673);
nor U17786 (N_17786,N_14997,N_15625);
nor U17787 (N_17787,N_14287,N_14532);
nand U17788 (N_17788,N_15607,N_15515);
xor U17789 (N_17789,N_15318,N_15854);
xnor U17790 (N_17790,N_14996,N_14675);
and U17791 (N_17791,N_15839,N_15477);
and U17792 (N_17792,N_15042,N_14339);
xor U17793 (N_17793,N_15802,N_15038);
or U17794 (N_17794,N_15124,N_14614);
nor U17795 (N_17795,N_15521,N_15553);
nand U17796 (N_17796,N_15798,N_14100);
or U17797 (N_17797,N_14422,N_15734);
nand U17798 (N_17798,N_14323,N_15929);
nor U17799 (N_17799,N_15512,N_14442);
xor U17800 (N_17800,N_15547,N_15711);
nor U17801 (N_17801,N_15876,N_14295);
xnor U17802 (N_17802,N_15045,N_14935);
nand U17803 (N_17803,N_14048,N_15286);
and U17804 (N_17804,N_15905,N_14402);
nand U17805 (N_17805,N_15135,N_15843);
and U17806 (N_17806,N_14160,N_15733);
and U17807 (N_17807,N_14273,N_14057);
and U17808 (N_17808,N_15686,N_14084);
nand U17809 (N_17809,N_15259,N_15102);
and U17810 (N_17810,N_15354,N_15720);
and U17811 (N_17811,N_14338,N_14228);
nor U17812 (N_17812,N_14249,N_14217);
xnor U17813 (N_17813,N_14231,N_15417);
xor U17814 (N_17814,N_15216,N_15513);
nor U17815 (N_17815,N_14399,N_15438);
or U17816 (N_17816,N_15513,N_15880);
and U17817 (N_17817,N_15043,N_15619);
and U17818 (N_17818,N_15695,N_14094);
xnor U17819 (N_17819,N_15714,N_14336);
xnor U17820 (N_17820,N_15484,N_15246);
nor U17821 (N_17821,N_14282,N_15092);
nand U17822 (N_17822,N_15376,N_14659);
nand U17823 (N_17823,N_14696,N_14543);
nand U17824 (N_17824,N_14082,N_15131);
nor U17825 (N_17825,N_15388,N_15178);
xnor U17826 (N_17826,N_14791,N_15239);
and U17827 (N_17827,N_14618,N_15194);
and U17828 (N_17828,N_14623,N_15937);
xor U17829 (N_17829,N_14546,N_14079);
and U17830 (N_17830,N_14327,N_15906);
and U17831 (N_17831,N_15829,N_15048);
xnor U17832 (N_17832,N_14489,N_15380);
nor U17833 (N_17833,N_15842,N_15708);
nor U17834 (N_17834,N_15419,N_15451);
nand U17835 (N_17835,N_15461,N_14149);
xnor U17836 (N_17836,N_15116,N_14675);
nand U17837 (N_17837,N_15834,N_15445);
or U17838 (N_17838,N_15653,N_14127);
or U17839 (N_17839,N_15239,N_14548);
xor U17840 (N_17840,N_14096,N_15459);
nand U17841 (N_17841,N_14789,N_14734);
xnor U17842 (N_17842,N_14472,N_15230);
nor U17843 (N_17843,N_15037,N_14308);
and U17844 (N_17844,N_14486,N_15320);
nor U17845 (N_17845,N_14933,N_15846);
xnor U17846 (N_17846,N_15855,N_15089);
nor U17847 (N_17847,N_15649,N_14772);
or U17848 (N_17848,N_15674,N_14120);
nor U17849 (N_17849,N_14074,N_15046);
or U17850 (N_17850,N_15299,N_14586);
nand U17851 (N_17851,N_15126,N_14573);
nor U17852 (N_17852,N_14221,N_14028);
nand U17853 (N_17853,N_15712,N_15614);
or U17854 (N_17854,N_14066,N_15243);
or U17855 (N_17855,N_14760,N_15372);
xor U17856 (N_17856,N_14364,N_15716);
and U17857 (N_17857,N_15204,N_14317);
nor U17858 (N_17858,N_15066,N_15751);
or U17859 (N_17859,N_14629,N_14077);
or U17860 (N_17860,N_15871,N_14741);
or U17861 (N_17861,N_14283,N_15232);
xor U17862 (N_17862,N_14098,N_14834);
nand U17863 (N_17863,N_14469,N_14415);
and U17864 (N_17864,N_14764,N_15941);
xnor U17865 (N_17865,N_15331,N_14686);
nand U17866 (N_17866,N_15178,N_15962);
nor U17867 (N_17867,N_15505,N_15780);
nand U17868 (N_17868,N_15701,N_15546);
and U17869 (N_17869,N_14456,N_15433);
xnor U17870 (N_17870,N_15254,N_14166);
nor U17871 (N_17871,N_14007,N_15146);
and U17872 (N_17872,N_14101,N_14918);
or U17873 (N_17873,N_15058,N_14532);
and U17874 (N_17874,N_15769,N_15663);
nand U17875 (N_17875,N_15210,N_15049);
nor U17876 (N_17876,N_15748,N_15043);
xor U17877 (N_17877,N_15335,N_15423);
nand U17878 (N_17878,N_15527,N_15950);
and U17879 (N_17879,N_15220,N_15006);
nor U17880 (N_17880,N_14566,N_14399);
and U17881 (N_17881,N_14388,N_14428);
xor U17882 (N_17882,N_14990,N_15865);
and U17883 (N_17883,N_14888,N_14153);
nor U17884 (N_17884,N_14573,N_15135);
and U17885 (N_17885,N_14508,N_14074);
or U17886 (N_17886,N_15423,N_14535);
nor U17887 (N_17887,N_14410,N_15005);
nor U17888 (N_17888,N_14494,N_15532);
nand U17889 (N_17889,N_15659,N_15834);
xor U17890 (N_17890,N_14833,N_14058);
xor U17891 (N_17891,N_14126,N_15330);
xnor U17892 (N_17892,N_14034,N_15925);
xnor U17893 (N_17893,N_15770,N_15622);
xor U17894 (N_17894,N_15405,N_14597);
or U17895 (N_17895,N_15673,N_14481);
nand U17896 (N_17896,N_15430,N_14272);
and U17897 (N_17897,N_14771,N_15956);
xnor U17898 (N_17898,N_15104,N_14419);
or U17899 (N_17899,N_15794,N_15321);
and U17900 (N_17900,N_15597,N_15180);
and U17901 (N_17901,N_15883,N_14358);
nor U17902 (N_17902,N_15574,N_15865);
and U17903 (N_17903,N_15429,N_14484);
nand U17904 (N_17904,N_15913,N_14156);
nand U17905 (N_17905,N_14825,N_14472);
xnor U17906 (N_17906,N_14632,N_15453);
xor U17907 (N_17907,N_14434,N_15590);
or U17908 (N_17908,N_15340,N_14136);
nor U17909 (N_17909,N_14089,N_15669);
or U17910 (N_17910,N_14724,N_14742);
or U17911 (N_17911,N_14266,N_15893);
and U17912 (N_17912,N_14229,N_14507);
and U17913 (N_17913,N_14199,N_14328);
xor U17914 (N_17914,N_14537,N_14579);
or U17915 (N_17915,N_14092,N_14829);
nor U17916 (N_17916,N_15918,N_15769);
nor U17917 (N_17917,N_15600,N_15372);
xnor U17918 (N_17918,N_14445,N_14151);
or U17919 (N_17919,N_15959,N_14580);
nand U17920 (N_17920,N_15389,N_14195);
and U17921 (N_17921,N_15869,N_15418);
and U17922 (N_17922,N_15328,N_15719);
and U17923 (N_17923,N_15080,N_15114);
nand U17924 (N_17924,N_15101,N_14156);
or U17925 (N_17925,N_14186,N_14281);
nor U17926 (N_17926,N_14168,N_15951);
nand U17927 (N_17927,N_14731,N_15670);
and U17928 (N_17928,N_15500,N_14175);
xnor U17929 (N_17929,N_14648,N_14978);
xor U17930 (N_17930,N_14010,N_15128);
or U17931 (N_17931,N_15071,N_14480);
or U17932 (N_17932,N_15186,N_15082);
nand U17933 (N_17933,N_14669,N_15853);
and U17934 (N_17934,N_15282,N_14327);
and U17935 (N_17935,N_15565,N_14701);
xnor U17936 (N_17936,N_14547,N_14319);
nand U17937 (N_17937,N_14745,N_15947);
xor U17938 (N_17938,N_15340,N_14852);
xor U17939 (N_17939,N_14545,N_15078);
and U17940 (N_17940,N_14886,N_15999);
or U17941 (N_17941,N_15445,N_14689);
and U17942 (N_17942,N_15726,N_14566);
xor U17943 (N_17943,N_14093,N_15186);
nor U17944 (N_17944,N_14408,N_15238);
or U17945 (N_17945,N_14812,N_15787);
or U17946 (N_17946,N_14841,N_15383);
nor U17947 (N_17947,N_14019,N_15753);
nand U17948 (N_17948,N_14320,N_14545);
xor U17949 (N_17949,N_15533,N_14803);
xor U17950 (N_17950,N_15011,N_15216);
and U17951 (N_17951,N_14331,N_15214);
xnor U17952 (N_17952,N_15259,N_14092);
and U17953 (N_17953,N_15513,N_14710);
and U17954 (N_17954,N_15673,N_15945);
xor U17955 (N_17955,N_15215,N_15670);
and U17956 (N_17956,N_14146,N_14249);
and U17957 (N_17957,N_15066,N_14918);
and U17958 (N_17958,N_15872,N_14078);
and U17959 (N_17959,N_14894,N_15220);
nor U17960 (N_17960,N_14830,N_15647);
nand U17961 (N_17961,N_15815,N_15223);
nor U17962 (N_17962,N_14527,N_14178);
xor U17963 (N_17963,N_14543,N_14422);
or U17964 (N_17964,N_14041,N_15934);
nor U17965 (N_17965,N_15512,N_14592);
nor U17966 (N_17966,N_14674,N_14150);
xor U17967 (N_17967,N_14995,N_15967);
xnor U17968 (N_17968,N_14992,N_15702);
nor U17969 (N_17969,N_15925,N_14469);
or U17970 (N_17970,N_15192,N_14784);
xor U17971 (N_17971,N_14590,N_14441);
nor U17972 (N_17972,N_15437,N_14900);
xor U17973 (N_17973,N_15499,N_14642);
or U17974 (N_17974,N_15963,N_15295);
nand U17975 (N_17975,N_15472,N_14804);
nor U17976 (N_17976,N_15936,N_15654);
or U17977 (N_17977,N_15281,N_15138);
or U17978 (N_17978,N_15708,N_15630);
nor U17979 (N_17979,N_14664,N_15207);
and U17980 (N_17980,N_14623,N_14319);
xnor U17981 (N_17981,N_15104,N_15651);
and U17982 (N_17982,N_15799,N_15883);
nor U17983 (N_17983,N_14386,N_14875);
xor U17984 (N_17984,N_15963,N_14339);
or U17985 (N_17985,N_15495,N_15718);
nand U17986 (N_17986,N_14319,N_15166);
nor U17987 (N_17987,N_15813,N_15223);
xor U17988 (N_17988,N_15496,N_15697);
and U17989 (N_17989,N_15721,N_14324);
nor U17990 (N_17990,N_15974,N_15386);
xnor U17991 (N_17991,N_14840,N_14421);
nor U17992 (N_17992,N_15250,N_15032);
and U17993 (N_17993,N_15968,N_15046);
nor U17994 (N_17994,N_14809,N_15601);
nor U17995 (N_17995,N_14736,N_14171);
nor U17996 (N_17996,N_15326,N_14452);
or U17997 (N_17997,N_14186,N_14464);
nand U17998 (N_17998,N_15510,N_15067);
xnor U17999 (N_17999,N_15122,N_15604);
nand U18000 (N_18000,N_16801,N_16909);
or U18001 (N_18001,N_17930,N_16800);
nand U18002 (N_18002,N_16564,N_16168);
xor U18003 (N_18003,N_17941,N_16252);
nor U18004 (N_18004,N_16085,N_16795);
nand U18005 (N_18005,N_17756,N_16754);
xor U18006 (N_18006,N_17480,N_17044);
nand U18007 (N_18007,N_17345,N_17051);
xnor U18008 (N_18008,N_16844,N_17934);
nand U18009 (N_18009,N_16456,N_16724);
nand U18010 (N_18010,N_16601,N_17655);
xor U18011 (N_18011,N_16481,N_16420);
and U18012 (N_18012,N_16772,N_17737);
nor U18013 (N_18013,N_17547,N_16256);
and U18014 (N_18014,N_17382,N_17230);
nor U18015 (N_18015,N_16857,N_16770);
xnor U18016 (N_18016,N_17103,N_17939);
nand U18017 (N_18017,N_17404,N_17327);
xnor U18018 (N_18018,N_17238,N_17426);
and U18019 (N_18019,N_17138,N_17469);
or U18020 (N_18020,N_17159,N_17007);
nand U18021 (N_18021,N_16209,N_16120);
nor U18022 (N_18022,N_17068,N_16982);
and U18023 (N_18023,N_17920,N_16683);
or U18024 (N_18024,N_16340,N_17525);
and U18025 (N_18025,N_16359,N_17052);
xnor U18026 (N_18026,N_17267,N_17447);
nand U18027 (N_18027,N_16297,N_16031);
nor U18028 (N_18028,N_16884,N_16693);
xnor U18029 (N_18029,N_16314,N_17643);
and U18030 (N_18030,N_16437,N_16415);
xor U18031 (N_18031,N_16237,N_17681);
nor U18032 (N_18032,N_17035,N_16161);
nor U18033 (N_18033,N_17039,N_16759);
xor U18034 (N_18034,N_16956,N_16465);
nor U18035 (N_18035,N_16814,N_17465);
nand U18036 (N_18036,N_16307,N_17748);
nand U18037 (N_18037,N_17272,N_16740);
xor U18038 (N_18038,N_17227,N_17126);
nand U18039 (N_18039,N_16331,N_17593);
or U18040 (N_18040,N_17600,N_17064);
or U18041 (N_18041,N_16952,N_17651);
or U18042 (N_18042,N_17770,N_16017);
nand U18043 (N_18043,N_17030,N_17178);
nor U18044 (N_18044,N_17149,N_16788);
nand U18045 (N_18045,N_16624,N_17925);
nor U18046 (N_18046,N_17164,N_17478);
xnor U18047 (N_18047,N_16293,N_16024);
and U18048 (N_18048,N_17792,N_17229);
xor U18049 (N_18049,N_16885,N_17496);
and U18050 (N_18050,N_17191,N_16512);
nand U18051 (N_18051,N_17485,N_16353);
or U18052 (N_18052,N_16692,N_17019);
and U18053 (N_18053,N_16295,N_16774);
nor U18054 (N_18054,N_17320,N_17251);
xor U18055 (N_18055,N_17658,N_16935);
or U18056 (N_18056,N_17607,N_17602);
nand U18057 (N_18057,N_16375,N_16521);
or U18058 (N_18058,N_17468,N_16078);
nor U18059 (N_18059,N_17460,N_17568);
and U18060 (N_18060,N_17606,N_16912);
nand U18061 (N_18061,N_16527,N_16253);
or U18062 (N_18062,N_17546,N_16696);
xnor U18063 (N_18063,N_17734,N_17528);
or U18064 (N_18064,N_16918,N_17249);
and U18065 (N_18065,N_17803,N_16779);
nand U18066 (N_18066,N_16294,N_17586);
nand U18067 (N_18067,N_16183,N_17882);
and U18068 (N_18068,N_17569,N_16407);
nor U18069 (N_18069,N_17660,N_16445);
and U18070 (N_18070,N_17384,N_16530);
and U18071 (N_18071,N_16549,N_16942);
and U18072 (N_18072,N_17054,N_16271);
or U18073 (N_18073,N_16852,N_16171);
nor U18074 (N_18074,N_16069,N_17332);
xor U18075 (N_18075,N_16762,N_16081);
nor U18076 (N_18076,N_17685,N_17859);
and U18077 (N_18077,N_16062,N_17334);
xnor U18078 (N_18078,N_16002,N_16948);
nand U18079 (N_18079,N_16750,N_17245);
or U18080 (N_18080,N_17890,N_16144);
xor U18081 (N_18081,N_16215,N_16094);
and U18082 (N_18082,N_16400,N_17183);
or U18083 (N_18083,N_16634,N_16323);
xor U18084 (N_18084,N_17169,N_17193);
xnor U18085 (N_18085,N_16810,N_17599);
nor U18086 (N_18086,N_17806,N_17142);
and U18087 (N_18087,N_17550,N_17309);
xor U18088 (N_18088,N_17872,N_17432);
and U18089 (N_18089,N_17451,N_16391);
nand U18090 (N_18090,N_17242,N_16711);
and U18091 (N_18091,N_17621,N_17036);
nor U18092 (N_18092,N_16819,N_17697);
nor U18093 (N_18093,N_16931,N_16495);
nor U18094 (N_18094,N_16454,N_16686);
nand U18095 (N_18095,N_16257,N_17832);
nor U18096 (N_18096,N_16090,N_17058);
or U18097 (N_18097,N_16838,N_16480);
and U18098 (N_18098,N_17491,N_16304);
or U18099 (N_18099,N_16139,N_16694);
nor U18100 (N_18100,N_17099,N_17217);
nand U18101 (N_18101,N_16608,N_17665);
xor U18102 (N_18102,N_16042,N_17758);
or U18103 (N_18103,N_17693,N_17707);
and U18104 (N_18104,N_17118,N_17701);
nand U18105 (N_18105,N_16650,N_16537);
and U18106 (N_18106,N_16211,N_16269);
and U18107 (N_18107,N_16673,N_16292);
xnor U18108 (N_18108,N_17290,N_16141);
nand U18109 (N_18109,N_16685,N_16467);
nor U18110 (N_18110,N_16337,N_17834);
xor U18111 (N_18111,N_17911,N_16434);
xor U18112 (N_18112,N_17298,N_16346);
or U18113 (N_18113,N_17801,N_16343);
or U18114 (N_18114,N_16172,N_17107);
or U18115 (N_18115,N_16700,N_16140);
nand U18116 (N_18116,N_17296,N_17316);
xor U18117 (N_18117,N_17605,N_17596);
nand U18118 (N_18118,N_16725,N_17458);
or U18119 (N_18119,N_17151,N_17720);
nand U18120 (N_18120,N_16843,N_16023);
xnor U18121 (N_18121,N_17495,N_17132);
nand U18122 (N_18122,N_17883,N_16846);
nand U18123 (N_18123,N_16996,N_16344);
nand U18124 (N_18124,N_17955,N_16243);
nor U18125 (N_18125,N_17056,N_16071);
nand U18126 (N_18126,N_16833,N_16433);
or U18127 (N_18127,N_16203,N_17603);
nand U18128 (N_18128,N_17899,N_16980);
nand U18129 (N_18129,N_17153,N_16084);
nor U18130 (N_18130,N_17269,N_16937);
nand U18131 (N_18131,N_17161,N_16338);
and U18132 (N_18132,N_17264,N_17223);
nor U18133 (N_18133,N_17993,N_17457);
nand U18134 (N_18134,N_17117,N_17340);
or U18135 (N_18135,N_17990,N_17235);
nand U18136 (N_18136,N_16721,N_16515);
and U18137 (N_18137,N_17255,N_16995);
xnor U18138 (N_18138,N_17415,N_16543);
nor U18139 (N_18139,N_16922,N_17696);
nor U18140 (N_18140,N_17517,N_17979);
nor U18141 (N_18141,N_17575,N_16888);
nor U18142 (N_18142,N_16164,N_17555);
and U18143 (N_18143,N_17816,N_16599);
xnor U18144 (N_18144,N_16580,N_16399);
xor U18145 (N_18145,N_16967,N_16339);
xor U18146 (N_18146,N_16881,N_17175);
or U18147 (N_18147,N_16315,N_16504);
xnor U18148 (N_18148,N_17545,N_17841);
nor U18149 (N_18149,N_17166,N_16904);
or U18150 (N_18150,N_17112,N_16986);
nand U18151 (N_18151,N_16575,N_17083);
xor U18152 (N_18152,N_17954,N_16545);
nand U18153 (N_18153,N_17704,N_17644);
and U18154 (N_18154,N_17474,N_17718);
and U18155 (N_18155,N_17472,N_16831);
nand U18156 (N_18156,N_16773,N_17139);
xnor U18157 (N_18157,N_16757,N_17127);
and U18158 (N_18158,N_17425,N_17443);
and U18159 (N_18159,N_16742,N_17160);
xor U18160 (N_18160,N_16127,N_17810);
xor U18161 (N_18161,N_17656,N_16901);
and U18162 (N_18162,N_17745,N_17817);
or U18163 (N_18163,N_17140,N_16476);
or U18164 (N_18164,N_16370,N_17520);
xor U18165 (N_18165,N_16897,N_16224);
xnor U18166 (N_18166,N_17900,N_17736);
nand U18167 (N_18167,N_16104,N_17595);
nand U18168 (N_18168,N_17738,N_17487);
xnor U18169 (N_18169,N_16500,N_16697);
nand U18170 (N_18170,N_16286,N_16201);
nor U18171 (N_18171,N_17612,N_17145);
or U18172 (N_18172,N_17972,N_17304);
xor U18173 (N_18173,N_17262,N_16733);
xor U18174 (N_18174,N_16109,N_16382);
and U18175 (N_18175,N_17870,N_17403);
nor U18176 (N_18176,N_16786,N_16197);
and U18177 (N_18177,N_17395,N_17985);
xnor U18178 (N_18178,N_17998,N_16080);
or U18179 (N_18179,N_16014,N_17312);
xor U18180 (N_18180,N_17089,N_17186);
nor U18181 (N_18181,N_17221,N_16933);
and U18182 (N_18182,N_16186,N_16616);
nand U18183 (N_18183,N_16923,N_17020);
or U18184 (N_18184,N_16726,N_17683);
nor U18185 (N_18185,N_17016,N_16064);
nand U18186 (N_18186,N_16548,N_16646);
or U18187 (N_18187,N_17833,N_16620);
nand U18188 (N_18188,N_17779,N_17638);
nand U18189 (N_18189,N_17809,N_17530);
or U18190 (N_18190,N_16479,N_16440);
nor U18191 (N_18191,N_17562,N_17503);
and U18192 (N_18192,N_17589,N_17659);
nor U18193 (N_18193,N_16503,N_16414);
and U18194 (N_18194,N_17009,N_17928);
nand U18195 (N_18195,N_16832,N_17452);
nor U18196 (N_18196,N_16571,N_17034);
nand U18197 (N_18197,N_16525,N_16588);
nor U18198 (N_18198,N_17579,N_16924);
xnor U18199 (N_18199,N_17845,N_17764);
xnor U18200 (N_18200,N_17887,N_16143);
nor U18201 (N_18201,N_17322,N_16491);
nor U18202 (N_18202,N_16988,N_17829);
or U18203 (N_18203,N_17971,N_17960);
and U18204 (N_18204,N_17556,N_17772);
and U18205 (N_18205,N_17592,N_17408);
or U18206 (N_18206,N_16609,N_17398);
or U18207 (N_18207,N_17891,N_16026);
nand U18208 (N_18208,N_17771,N_16475);
and U18209 (N_18209,N_17668,N_16802);
and U18210 (N_18210,N_16817,N_16121);
nand U18211 (N_18211,N_17086,N_16054);
or U18212 (N_18212,N_16863,N_16134);
and U18213 (N_18213,N_17385,N_17308);
nor U18214 (N_18214,N_16413,N_17987);
nor U18215 (N_18215,N_17753,N_17130);
and U18216 (N_18216,N_16283,N_16342);
or U18217 (N_18217,N_16122,N_16446);
nand U18218 (N_18218,N_16805,N_16883);
nor U18219 (N_18219,N_16984,N_16036);
and U18220 (N_18220,N_17553,N_17512);
and U18221 (N_18221,N_17288,N_17361);
nor U18222 (N_18222,N_16493,N_16579);
nand U18223 (N_18223,N_16751,N_16153);
xor U18224 (N_18224,N_16688,N_16979);
nand U18225 (N_18225,N_17261,N_16566);
or U18226 (N_18226,N_17096,N_17949);
xnor U18227 (N_18227,N_17195,N_17807);
nand U18228 (N_18228,N_17860,N_16507);
nor U18229 (N_18229,N_17134,N_16428);
or U18230 (N_18230,N_16214,N_17893);
nand U18231 (N_18231,N_17709,N_16514);
nand U18232 (N_18232,N_16739,N_16990);
nand U18233 (N_18233,N_16011,N_16418);
or U18234 (N_18234,N_16939,N_16510);
nor U18235 (N_18235,N_16859,N_17319);
and U18236 (N_18236,N_17077,N_16066);
or U18237 (N_18237,N_17078,N_17079);
xnor U18238 (N_18238,N_16112,N_17348);
nor U18239 (N_18239,N_16334,N_16189);
nor U18240 (N_18240,N_16424,N_17690);
or U18241 (N_18241,N_16657,N_17208);
nor U18242 (N_18242,N_16185,N_16596);
or U18243 (N_18243,N_17097,N_16861);
or U18244 (N_18244,N_16871,N_16508);
and U18245 (N_18245,N_16971,N_16992);
nand U18246 (N_18246,N_17511,N_17179);
or U18247 (N_18247,N_17411,N_17610);
xnor U18248 (N_18248,N_17435,N_16749);
nor U18249 (N_18249,N_17703,N_16964);
and U18250 (N_18250,N_17866,N_16691);
xor U18251 (N_18251,N_17198,N_16277);
xnor U18252 (N_18252,N_16787,N_16652);
nor U18253 (N_18253,N_17090,N_16132);
nor U18254 (N_18254,N_17847,N_17396);
and U18255 (N_18255,N_16572,N_17342);
nand U18256 (N_18256,N_17513,N_16238);
or U18257 (N_18257,N_16917,N_16597);
nand U18258 (N_18258,N_17826,N_17677);
xnor U18259 (N_18259,N_17494,N_16276);
and U18260 (N_18260,N_16517,N_17306);
nor U18261 (N_18261,N_16086,N_16825);
nor U18262 (N_18262,N_17909,N_16605);
or U18263 (N_18263,N_16060,N_17409);
xnor U18264 (N_18264,N_16803,N_17420);
or U18265 (N_18265,N_16676,N_16371);
nand U18266 (N_18266,N_17314,N_17733);
nor U18267 (N_18267,N_16151,N_16460);
nand U18268 (N_18268,N_17601,N_17956);
nand U18269 (N_18269,N_16973,N_16160);
or U18270 (N_18270,N_17258,N_17002);
or U18271 (N_18271,N_16578,N_17021);
or U18272 (N_18272,N_16645,N_17046);
nand U18273 (N_18273,N_16505,N_17578);
and U18274 (N_18274,N_17618,N_17490);
or U18275 (N_18275,N_16077,N_16560);
and U18276 (N_18276,N_16226,N_16748);
or U18277 (N_18277,N_16305,N_16797);
xnor U18278 (N_18278,N_16858,N_17973);
and U18279 (N_18279,N_17347,N_17184);
and U18280 (N_18280,N_17984,N_16099);
and U18281 (N_18281,N_16722,N_17011);
nand U18282 (N_18282,N_16533,N_16870);
xnor U18283 (N_18283,N_16589,N_17522);
xor U18284 (N_18284,N_17781,N_17699);
or U18285 (N_18285,N_16875,N_16594);
or U18286 (N_18286,N_16181,N_17880);
nor U18287 (N_18287,N_16894,N_16671);
xnor U18288 (N_18288,N_17504,N_16007);
nor U18289 (N_18289,N_17042,N_17957);
nand U18290 (N_18290,N_16585,N_17561);
xnor U18291 (N_18291,N_16532,N_17529);
xnor U18292 (N_18292,N_16959,N_16674);
nor U18293 (N_18293,N_17004,N_17028);
and U18294 (N_18294,N_16473,N_16963);
and U18295 (N_18295,N_17233,N_16115);
xnor U18296 (N_18296,N_16372,N_16022);
and U18297 (N_18297,N_17231,N_16010);
nor U18298 (N_18298,N_17855,N_16622);
and U18299 (N_18299,N_16734,N_17263);
nand U18300 (N_18300,N_16053,N_16651);
nor U18301 (N_18301,N_17811,N_16577);
and U18302 (N_18302,N_16272,N_17199);
and U18303 (N_18303,N_17067,N_16553);
and U18304 (N_18304,N_16488,N_17102);
xnor U18305 (N_18305,N_17317,N_17326);
nand U18306 (N_18306,N_16267,N_17624);
or U18307 (N_18307,N_17869,N_17678);
and U18308 (N_18308,N_17167,N_17481);
nand U18309 (N_18309,N_16777,N_16983);
nor U18310 (N_18310,N_16157,N_16463);
or U18311 (N_18311,N_17148,N_17910);
nor U18312 (N_18312,N_16771,N_17172);
xor U18313 (N_18313,N_16329,N_16619);
or U18314 (N_18314,N_16710,N_17266);
xnor U18315 (N_18315,N_16953,N_16233);
nand U18316 (N_18316,N_17563,N_17414);
nor U18317 (N_18317,N_17275,N_17006);
xor U18318 (N_18318,N_16856,N_16173);
or U18319 (N_18319,N_16001,N_16117);
xor U18320 (N_18320,N_17749,N_16430);
xnor U18321 (N_18321,N_16868,N_17774);
xor U18322 (N_18322,N_16075,N_17615);
and U18323 (N_18323,N_16326,N_17544);
nor U18324 (N_18324,N_17372,N_16860);
nand U18325 (N_18325,N_16705,N_16393);
xor U18326 (N_18326,N_16116,N_17280);
nand U18327 (N_18327,N_17588,N_16535);
nand U18328 (N_18328,N_17785,N_17370);
and U18329 (N_18329,N_16902,N_16177);
or U18330 (N_18330,N_17669,N_16898);
or U18331 (N_18331,N_17551,N_16494);
nor U18332 (N_18332,N_16730,N_16887);
xnor U18333 (N_18333,N_17081,N_16546);
or U18334 (N_18334,N_16039,N_17968);
and U18335 (N_18335,N_17210,N_17339);
nor U18336 (N_18336,N_16999,N_17767);
nand U18337 (N_18337,N_17093,N_17234);
nand U18338 (N_18338,N_17514,N_16110);
nor U18339 (N_18339,N_16526,N_16679);
or U18340 (N_18340,N_17057,N_16408);
nand U18341 (N_18341,N_17988,N_16487);
nor U18342 (N_18342,N_16641,N_17804);
or U18343 (N_18343,N_16431,N_17903);
nand U18344 (N_18344,N_17824,N_17356);
nor U18345 (N_18345,N_16354,N_16236);
nor U18346 (N_18346,N_16732,N_17653);
nor U18347 (N_18347,N_16669,N_17115);
nor U18348 (N_18348,N_16621,N_16643);
or U18349 (N_18349,N_17947,N_16944);
nor U18350 (N_18350,N_17325,N_16205);
xor U18351 (N_18351,N_16389,N_17508);
and U18352 (N_18352,N_16135,N_16222);
nor U18353 (N_18353,N_17815,N_17446);
and U18354 (N_18354,N_16497,N_16125);
and U18355 (N_18355,N_16264,N_16296);
or U18356 (N_18356,N_16013,N_17688);
or U18357 (N_18357,N_17477,N_17228);
and U18358 (N_18358,N_16174,N_16442);
nor U18359 (N_18359,N_16715,N_17085);
nor U18360 (N_18360,N_17843,N_17591);
nand U18361 (N_18361,N_17784,N_17800);
and U18362 (N_18362,N_16511,N_16103);
xnor U18363 (N_18363,N_17453,N_16028);
xnor U18364 (N_18364,N_17691,N_17302);
nand U18365 (N_18365,N_17566,N_16718);
and U18366 (N_18366,N_16321,N_16630);
nand U18367 (N_18367,N_17486,N_16111);
nor U18368 (N_18368,N_16358,N_16877);
nand U18369 (N_18369,N_16325,N_17884);
nor U18370 (N_18370,N_17360,N_17715);
nor U18371 (N_18371,N_16486,N_16204);
nor U18372 (N_18372,N_16438,N_16290);
or U18373 (N_18373,N_17397,N_17462);
nand U18374 (N_18374,N_16170,N_16416);
or U18375 (N_18375,N_16347,N_17676);
nor U18376 (N_18376,N_17023,N_16386);
and U18377 (N_18377,N_17141,N_17277);
nor U18378 (N_18378,N_17997,N_16466);
xor U18379 (N_18379,N_17136,N_16761);
nor U18380 (N_18380,N_16941,N_16012);
nand U18381 (N_18381,N_17428,N_17466);
or U18382 (N_18382,N_16083,N_17790);
and U18383 (N_18383,N_16576,N_16464);
nand U18384 (N_18384,N_17844,N_16152);
and U18385 (N_18385,N_17521,N_16513);
nor U18386 (N_18386,N_17782,N_16441);
xor U18387 (N_18387,N_16969,N_16449);
nor U18388 (N_18388,N_17284,N_16108);
nand U18389 (N_18389,N_16426,N_16743);
nor U18390 (N_18390,N_16310,N_17448);
xor U18391 (N_18391,N_16425,N_16113);
nor U18392 (N_18392,N_17388,N_16301);
and U18393 (N_18393,N_17819,N_17323);
xnor U18394 (N_18394,N_17366,N_16583);
or U18395 (N_18395,N_17597,N_16397);
nand U18396 (N_18396,N_17357,N_16394);
or U18397 (N_18397,N_16736,N_16854);
or U18398 (N_18398,N_17524,N_16390);
and U18399 (N_18399,N_16586,N_17560);
nor U18400 (N_18400,N_17055,N_16167);
or U18401 (N_18401,N_17037,N_17976);
or U18402 (N_18402,N_17461,N_16395);
nor U18403 (N_18403,N_16096,N_17125);
or U18404 (N_18404,N_16220,N_17212);
and U18405 (N_18405,N_17265,N_17247);
xnor U18406 (N_18406,N_17885,N_16383);
nor U18407 (N_18407,N_17814,N_16960);
or U18408 (N_18408,N_16044,N_17611);
nor U18409 (N_18409,N_16385,N_17013);
xor U18410 (N_18410,N_17392,N_16444);
or U18411 (N_18411,N_17619,N_16462);
and U18412 (N_18412,N_16194,N_17661);
nand U18413 (N_18413,N_17454,N_17837);
nor U18414 (N_18414,N_16058,N_17029);
nor U18415 (N_18415,N_16753,N_16516);
or U18416 (N_18416,N_17307,N_17857);
or U18417 (N_18417,N_17202,N_17427);
xor U18418 (N_18418,N_16274,N_17338);
and U18419 (N_18419,N_16855,N_16794);
nand U18420 (N_18420,N_16632,N_16542);
nand U18421 (N_18421,N_17390,N_17436);
xnor U18422 (N_18422,N_16807,N_16138);
or U18423 (N_18423,N_16929,N_16250);
nor U18424 (N_18424,N_16541,N_16617);
and U18425 (N_18425,N_16539,N_16218);
xnor U18426 (N_18426,N_16925,N_16792);
and U18427 (N_18427,N_17080,N_16328);
or U18428 (N_18428,N_16492,N_16148);
nor U18429 (N_18429,N_17673,N_16768);
nor U18430 (N_18430,N_16972,N_16489);
and U18431 (N_18431,N_16166,N_17587);
or U18432 (N_18432,N_16945,N_17027);
nor U18433 (N_18433,N_16633,N_17576);
and U18434 (N_18434,N_16207,N_16478);
nand U18435 (N_18435,N_16208,N_17146);
xor U18436 (N_18436,N_16610,N_16196);
or U18437 (N_18437,N_17672,N_16363);
and U18438 (N_18438,N_17399,N_16200);
xor U18439 (N_18439,N_16997,N_16065);
or U18440 (N_18440,N_16581,N_17573);
or U18441 (N_18441,N_16627,N_16607);
nand U18442 (N_18442,N_16092,N_17725);
xnor U18443 (N_18443,N_16752,N_17268);
nand U18444 (N_18444,N_17680,N_17209);
or U18445 (N_18445,N_17516,N_17482);
nor U18446 (N_18446,N_17331,N_17025);
nand U18447 (N_18447,N_16049,N_16662);
nor U18448 (N_18448,N_16745,N_17059);
and U18449 (N_18449,N_17789,N_16509);
nand U18450 (N_18450,N_16019,N_17548);
nor U18451 (N_18451,N_17813,N_16558);
nand U18452 (N_18452,N_16260,N_16443);
xor U18453 (N_18453,N_17113,N_17510);
nand U18454 (N_18454,N_16074,N_17625);
or U18455 (N_18455,N_17200,N_17959);
and U18456 (N_18456,N_17005,N_17978);
xnor U18457 (N_18457,N_17786,N_17286);
nand U18458 (N_18458,N_17996,N_17507);
nand U18459 (N_18459,N_17867,N_16038);
and U18460 (N_18460,N_17418,N_16682);
nand U18461 (N_18461,N_16618,N_16198);
nand U18462 (N_18462,N_16760,N_17483);
or U18463 (N_18463,N_17122,N_16896);
nand U18464 (N_18464,N_16298,N_16848);
nor U18465 (N_18465,N_17726,N_16247);
nand U18466 (N_18466,N_16406,N_17747);
nand U18467 (N_18467,N_17250,N_16658);
nor U18468 (N_18468,N_17048,N_17620);
nand U18469 (N_18469,N_16087,N_16920);
or U18470 (N_18470,N_16958,N_16384);
and U18471 (N_18471,N_16365,N_17675);
nand U18472 (N_18472,N_16806,N_17763);
and U18473 (N_18473,N_16891,N_16584);
and U18474 (N_18474,N_17654,N_17123);
nor U18475 (N_18475,N_16239,N_17635);
nor U18476 (N_18476,N_17329,N_16879);
xnor U18477 (N_18477,N_16769,N_17904);
xor U18478 (N_18478,N_16661,N_17073);
and U18479 (N_18479,N_17594,N_16699);
xnor U18480 (N_18480,N_17907,N_17886);
xnor U18481 (N_18481,N_16573,N_16570);
nand U18482 (N_18482,N_16206,N_17818);
nor U18483 (N_18483,N_16317,N_17951);
nor U18484 (N_18484,N_17087,N_17564);
nor U18485 (N_18485,N_16279,N_17211);
nor U18486 (N_18486,N_17889,N_16823);
nor U18487 (N_18487,N_16427,N_16072);
nand U18488 (N_18488,N_17853,N_16993);
xnor U18489 (N_18489,N_17359,N_16341);
nor U18490 (N_18490,N_17389,N_16974);
or U18491 (N_18491,N_17684,N_17032);
and U18492 (N_18492,N_16635,N_16114);
and U18493 (N_18493,N_17358,N_17922);
nand U18494 (N_18494,N_16333,N_16303);
and U18495 (N_18495,N_16865,N_16849);
and U18496 (N_18496,N_17430,N_17858);
or U18497 (N_18497,N_17194,N_16559);
or U18498 (N_18498,N_17613,N_16035);
nand U18499 (N_18499,N_17670,N_17614);
or U18500 (N_18500,N_17986,N_17901);
and U18501 (N_18501,N_17927,N_16677);
xor U18502 (N_18502,N_16193,N_16006);
or U18503 (N_18503,N_17964,N_17791);
or U18504 (N_18504,N_17967,N_17040);
xor U18505 (N_18505,N_16895,N_17041);
and U18506 (N_18506,N_17567,N_16182);
xor U18507 (N_18507,N_16815,N_17671);
or U18508 (N_18508,N_17850,N_17963);
nand U18509 (N_18509,N_16082,N_16936);
or U18510 (N_18510,N_17994,N_16978);
xor U18511 (N_18511,N_16401,N_17154);
xor U18512 (N_18512,N_16351,N_17554);
xor U18513 (N_18513,N_16380,N_17049);
nand U18514 (N_18514,N_17727,N_16563);
nor U18515 (N_18515,N_17535,N_17240);
or U18516 (N_18516,N_17173,N_16240);
xnor U18517 (N_18517,N_17352,N_17515);
nand U18518 (N_18518,N_16519,N_16899);
and U18519 (N_18519,N_17995,N_17641);
or U18520 (N_18520,N_16921,N_16192);
or U18521 (N_18521,N_16951,N_17918);
nand U18522 (N_18522,N_17757,N_16088);
or U18523 (N_18523,N_16411,N_16100);
nand U18524 (N_18524,N_16606,N_17463);
nor U18525 (N_18525,N_16142,N_17735);
and U18526 (N_18526,N_17645,N_17741);
nor U18527 (N_18527,N_16499,N_16528);
and U18528 (N_18528,N_17527,N_16020);
and U18529 (N_18529,N_17022,N_16009);
xnor U18530 (N_18530,N_17038,N_17788);
and U18531 (N_18531,N_17892,N_16033);
xnor U18532 (N_18532,N_17623,N_16587);
and U18533 (N_18533,N_17768,N_16714);
nand U18534 (N_18534,N_16919,N_17616);
and U18535 (N_18535,N_16522,N_16723);
xor U18536 (N_18536,N_17794,N_16713);
and U18537 (N_18537,N_16309,N_17337);
nand U18538 (N_18538,N_16158,N_16763);
and U18539 (N_18539,N_17689,N_17371);
nor U18540 (N_18540,N_17752,N_17121);
xnor U18541 (N_18541,N_17831,N_17874);
or U18542 (N_18542,N_16938,N_17248);
nand U18543 (N_18543,N_16005,N_16977);
and U18544 (N_18544,N_17537,N_17271);
xor U18545 (N_18545,N_17559,N_16934);
or U18546 (N_18546,N_16822,N_16629);
and U18547 (N_18547,N_16133,N_16502);
or U18548 (N_18548,N_16808,N_17921);
xor U18549 (N_18549,N_16387,N_16813);
nand U18550 (N_18550,N_16318,N_16656);
and U18551 (N_18551,N_17050,N_16241);
or U18552 (N_18552,N_16107,N_17254);
and U18553 (N_18553,N_17923,N_16423);
nand U18554 (N_18554,N_16095,N_16379);
nor U18555 (N_18555,N_16003,N_16287);
xor U18556 (N_18556,N_16335,N_17953);
xnor U18557 (N_18557,N_17877,N_17863);
or U18558 (N_18558,N_17917,N_17297);
xor U18559 (N_18559,N_17662,N_17642);
nand U18560 (N_18560,N_16275,N_17473);
and U18561 (N_18561,N_16778,N_17000);
nand U18562 (N_18562,N_16320,N_16202);
nand U18563 (N_18563,N_16962,N_17285);
nand U18564 (N_18564,N_16940,N_17731);
xor U18565 (N_18565,N_16998,N_16811);
nor U18566 (N_18566,N_16916,N_17449);
nor U18567 (N_18567,N_17256,N_16348);
or U18568 (N_18568,N_17876,N_17378);
nor U18569 (N_18569,N_16712,N_16506);
and U18570 (N_18570,N_17075,N_17765);
or U18571 (N_18571,N_17065,N_17224);
nor U18572 (N_18572,N_16332,N_16524);
nand U18573 (N_18573,N_16738,N_17293);
nand U18574 (N_18574,N_16242,N_17730);
or U18575 (N_18575,N_17188,N_17295);
or U18576 (N_18576,N_16637,N_16690);
or U18577 (N_18577,N_17137,N_17830);
nor U18578 (N_18578,N_17180,N_16366);
and U18579 (N_18579,N_17270,N_16518);
or U18580 (N_18580,N_17700,N_17970);
or U18581 (N_18581,N_16367,N_17201);
xor U18582 (N_18582,N_16653,N_17419);
and U18583 (N_18583,N_16647,N_17156);
nor U18584 (N_18584,N_16052,N_17565);
nor U18585 (N_18585,N_16642,N_16364);
nand U18586 (N_18586,N_16655,N_17629);
and U18587 (N_18587,N_16150,N_17335);
or U18588 (N_18588,N_17407,N_16450);
nor U18589 (N_18589,N_17539,N_17914);
nand U18590 (N_18590,N_16876,N_16649);
and U18591 (N_18591,N_16258,N_16396);
nor U18592 (N_18592,N_17375,N_16728);
nand U18593 (N_18593,N_16403,N_16529);
nor U18594 (N_18594,N_16105,N_16664);
and U18595 (N_18595,N_17861,N_16316);
xnor U18596 (N_18596,N_17871,N_16229);
nor U18597 (N_18597,N_17740,N_16284);
and U18598 (N_18598,N_16034,N_16567);
and U18599 (N_18599,N_16191,N_17341);
nor U18600 (N_18600,N_16322,N_17413);
xnor U18601 (N_18601,N_16015,N_16793);
and U18602 (N_18602,N_17572,N_17958);
nor U18603 (N_18603,N_16994,N_16392);
nor U18604 (N_18604,N_17732,N_16886);
nor U18605 (N_18605,N_16631,N_17098);
and U18606 (N_18606,N_16246,N_16612);
and U18607 (N_18607,N_17253,N_17484);
nand U18608 (N_18608,N_17364,N_17260);
nor U18609 (N_18609,N_17835,N_17849);
xnor U18610 (N_18610,N_16747,N_16903);
nor U18611 (N_18611,N_17232,N_17031);
nand U18612 (N_18612,N_16136,N_16225);
or U18613 (N_18613,N_16966,N_16663);
or U18614 (N_18614,N_16744,N_17823);
and U18615 (N_18615,N_16289,N_17218);
and U18616 (N_18616,N_17674,N_17429);
and U18617 (N_18617,N_17303,N_17437);
nand U18618 (N_18618,N_16217,N_17590);
xnor U18619 (N_18619,N_17424,N_17150);
xor U18620 (N_18620,N_16531,N_17336);
xor U18621 (N_18621,N_16369,N_17147);
nand U18622 (N_18622,N_17760,N_17383);
nand U18623 (N_18623,N_17394,N_16862);
and U18624 (N_18624,N_16534,N_16595);
nor U18625 (N_18625,N_16299,N_16569);
and U18626 (N_18626,N_16212,N_17365);
nand U18627 (N_18627,N_16949,N_17283);
xor U18628 (N_18628,N_16930,N_16568);
nand U18629 (N_18629,N_17489,N_16781);
xnor U18630 (N_18630,N_17281,N_16668);
xor U18631 (N_18631,N_17192,N_16356);
xor U18632 (N_18632,N_16536,N_17328);
xor U18633 (N_18633,N_17533,N_17205);
xor U18634 (N_18634,N_16667,N_16636);
or U18635 (N_18635,N_17091,N_16523);
or U18636 (N_18636,N_17915,N_17724);
and U18637 (N_18637,N_17444,N_16552);
or U18638 (N_18638,N_16041,N_16417);
nand U18639 (N_18639,N_16538,N_16459);
nor U18640 (N_18640,N_16602,N_16412);
and U18641 (N_18641,N_17505,N_17467);
and U18642 (N_18642,N_16175,N_17558);
and U18643 (N_18643,N_16735,N_16235);
xnor U18644 (N_18644,N_17931,N_16291);
and U18645 (N_18645,N_16251,N_17557);
nor U18646 (N_18646,N_17543,N_17750);
or U18647 (N_18647,N_17082,N_16357);
or U18648 (N_18648,N_17464,N_17220);
or U18649 (N_18649,N_16300,N_16821);
and U18650 (N_18650,N_17313,N_16056);
nand U18651 (N_18651,N_16613,N_17300);
or U18652 (N_18652,N_17416,N_16180);
or U18653 (N_18653,N_17157,N_16050);
xor U18654 (N_18654,N_16681,N_17024);
nand U18655 (N_18655,N_17840,N_16470);
or U18656 (N_18656,N_17761,N_17330);
xor U18657 (N_18657,N_17744,N_16227);
xnor U18658 (N_18658,N_17708,N_17652);
xor U18659 (N_18659,N_16282,N_17318);
or U18660 (N_18660,N_16263,N_16927);
or U18661 (N_18661,N_17913,N_16178);
nor U18662 (N_18662,N_17932,N_16872);
and U18663 (N_18663,N_17694,N_17476);
and U18664 (N_18664,N_17060,N_16043);
xor U18665 (N_18665,N_16791,N_16840);
xnor U18666 (N_18666,N_16890,N_17942);
nor U18667 (N_18667,N_17924,N_17321);
nand U18668 (N_18668,N_17310,N_16708);
and U18669 (N_18669,N_16265,N_17001);
nand U18670 (N_18670,N_16234,N_16302);
xor U18671 (N_18671,N_16675,N_16782);
and U18672 (N_18672,N_17975,N_17155);
nand U18673 (N_18673,N_16270,N_16368);
nor U18674 (N_18674,N_16232,N_17983);
and U18675 (N_18675,N_17053,N_16068);
xnor U18676 (N_18676,N_16447,N_17120);
and U18677 (N_18677,N_16654,N_17581);
or U18678 (N_18678,N_16405,N_17204);
nor U18679 (N_18679,N_17379,N_16824);
and U18680 (N_18680,N_17391,N_16163);
nand U18681 (N_18681,N_17937,N_16716);
xor U18682 (N_18682,N_16402,N_16016);
nor U18683 (N_18683,N_17165,N_16565);
nand U18684 (N_18684,N_16623,N_17189);
nor U18685 (N_18685,N_16847,N_16021);
nor U18686 (N_18686,N_17519,N_17999);
nor U18687 (N_18687,N_17351,N_17965);
xor U18688 (N_18688,N_17584,N_17292);
and U18689 (N_18689,N_17762,N_16834);
xnor U18690 (N_18690,N_17061,N_17992);
nor U18691 (N_18691,N_16336,N_17438);
or U18692 (N_18692,N_16169,N_16288);
or U18693 (N_18693,N_17908,N_17881);
and U18694 (N_18694,N_17825,N_16561);
nor U18695 (N_18695,N_17174,N_17634);
and U18696 (N_18696,N_17518,N_16550);
or U18697 (N_18697,N_17094,N_16955);
and U18698 (N_18698,N_17627,N_17241);
nor U18699 (N_18699,N_16970,N_17109);
xor U18700 (N_18700,N_17666,N_17943);
nor U18701 (N_18701,N_16432,N_17380);
or U18702 (N_18702,N_17856,N_17962);
xor U18703 (N_18703,N_17777,N_16882);
or U18704 (N_18704,N_17033,N_17354);
nand U18705 (N_18705,N_17092,N_17754);
nor U18706 (N_18706,N_16910,N_16866);
nor U18707 (N_18707,N_16907,N_17244);
nand U18708 (N_18708,N_16162,N_17609);
and U18709 (N_18709,N_17207,N_16231);
nand U18710 (N_18710,N_17775,N_17349);
nor U18711 (N_18711,N_16555,N_16737);
nor U18712 (N_18712,N_16373,N_16900);
nor U18713 (N_18713,N_16377,N_16210);
and U18714 (N_18714,N_17152,N_17664);
xnor U18715 (N_18715,N_17176,N_17226);
nand U18716 (N_18716,N_16626,N_16954);
and U18717 (N_18717,N_16471,N_17177);
nor U18718 (N_18718,N_16767,N_16461);
and U18719 (N_18719,N_16027,N_16482);
and U18720 (N_18720,N_17129,N_17100);
or U18721 (N_18721,N_16051,N_17362);
nand U18722 (N_18722,N_17470,N_16458);
or U18723 (N_18723,N_17222,N_17273);
nand U18724 (N_18724,N_17868,N_16439);
and U18725 (N_18725,N_17509,N_17713);
and U18726 (N_18726,N_16118,N_17440);
nor U18727 (N_18727,N_17206,N_16073);
or U18728 (N_18728,N_17014,N_17095);
and U18729 (N_18729,N_17812,N_17439);
nand U18730 (N_18730,N_16689,N_17719);
xnor U18731 (N_18731,N_16764,N_17864);
nand U18732 (N_18732,N_16851,N_16436);
xor U18733 (N_18733,N_16985,N_16991);
or U18734 (N_18734,N_17219,N_17343);
nor U18735 (N_18735,N_16574,N_16809);
xnor U18736 (N_18736,N_16130,N_16409);
and U18737 (N_18737,N_17898,N_16741);
nor U18738 (N_18738,N_17433,N_17353);
and U18739 (N_18739,N_16047,N_16032);
or U18740 (N_18740,N_17633,N_17896);
nand U18741 (N_18741,N_17854,N_17369);
and U18742 (N_18742,N_16199,N_16829);
nand U18743 (N_18743,N_17906,N_17196);
nor U18744 (N_18744,N_17015,N_17948);
xor U18745 (N_18745,N_16244,N_17894);
nor U18746 (N_18746,N_17531,N_16603);
or U18747 (N_18747,N_16796,N_16483);
and U18748 (N_18748,N_16349,N_16614);
xor U18749 (N_18749,N_17702,N_16248);
nor U18750 (N_18750,N_16404,N_16477);
or U18751 (N_18751,N_16154,N_16453);
and U18752 (N_18752,N_16701,N_17929);
nand U18753 (N_18753,N_16746,N_16262);
nor U18754 (N_18754,N_17974,N_16145);
nand U18755 (N_18755,N_17966,N_16448);
nor U18756 (N_18756,N_17492,N_17344);
nor U18757 (N_18757,N_17821,N_16398);
xor U18758 (N_18758,N_17066,N_16867);
or U18759 (N_18759,N_16281,N_17632);
and U18760 (N_18760,N_17766,N_17101);
or U18761 (N_18761,N_16421,N_17950);
nand U18762 (N_18762,N_17311,N_16000);
xnor U18763 (N_18763,N_16451,N_16947);
and U18764 (N_18764,N_16091,N_17170);
nor U18765 (N_18765,N_16485,N_17969);
and U18766 (N_18766,N_16784,N_16278);
nand U18767 (N_18767,N_17536,N_17523);
or U18768 (N_18768,N_17582,N_17778);
nor U18769 (N_18769,N_17946,N_17549);
nor U18770 (N_18770,N_17069,N_16932);
or U18771 (N_18771,N_17798,N_17422);
nor U18772 (N_18772,N_16914,N_17162);
nor U18773 (N_18773,N_17583,N_16376);
nor U18774 (N_18774,N_17018,N_16223);
xnor U18775 (N_18775,N_16119,N_16709);
and U18776 (N_18776,N_16704,N_17787);
nand U18777 (N_18777,N_16702,N_17695);
xnor U18778 (N_18778,N_16950,N_16845);
nand U18779 (N_18779,N_17500,N_17729);
and U18780 (N_18780,N_16419,N_16915);
xor U18781 (N_18781,N_17679,N_16975);
or U18782 (N_18782,N_17291,N_16837);
or U18783 (N_18783,N_16600,N_17008);
nand U18784 (N_18784,N_17236,N_16057);
xnor U18785 (N_18785,N_16249,N_16592);
nand U18786 (N_18786,N_16640,N_17526);
nand U18787 (N_18787,N_17074,N_16374);
nor U18788 (N_18788,N_16018,N_16987);
or U18789 (N_18789,N_17216,N_16255);
nor U18790 (N_18790,N_16037,N_16869);
and U18791 (N_18791,N_16123,N_17128);
and U18792 (N_18792,N_16828,N_17497);
xnor U18793 (N_18793,N_16147,N_16961);
nand U18794 (N_18794,N_17839,N_16812);
xor U18795 (N_18795,N_17755,N_16228);
and U18796 (N_18796,N_16818,N_16727);
nand U18797 (N_18797,N_16455,N_17628);
nor U18798 (N_18798,N_17421,N_16625);
or U18799 (N_18799,N_16665,N_16490);
nor U18800 (N_18800,N_17105,N_16965);
xnor U18801 (N_18801,N_17940,N_17862);
nand U18802 (N_18802,N_16706,N_16680);
nor U18803 (N_18803,N_16659,N_17299);
and U18804 (N_18804,N_16864,N_17278);
nor U18805 (N_18805,N_17982,N_17190);
nand U18806 (N_18806,N_17650,N_17187);
and U18807 (N_18807,N_16765,N_16946);
xnor U18808 (N_18808,N_17181,N_16273);
nor U18809 (N_18809,N_17919,N_17751);
and U18810 (N_18810,N_17406,N_17716);
nor U18811 (N_18811,N_17088,N_16678);
nor U18812 (N_18812,N_17977,N_16155);
and U18813 (N_18813,N_17598,N_17493);
nand U18814 (N_18814,N_16219,N_17423);
xor U18815 (N_18815,N_16190,N_17728);
xnor U18816 (N_18816,N_17852,N_17043);
xnor U18817 (N_18817,N_17315,N_17604);
nand U18818 (N_18818,N_17114,N_17711);
xor U18819 (N_18819,N_16230,N_17836);
or U18820 (N_18820,N_16245,N_16008);
xnor U18821 (N_18821,N_16804,N_17279);
nor U18822 (N_18822,N_16707,N_17355);
nor U18823 (N_18823,N_17062,N_16591);
nor U18824 (N_18824,N_17552,N_16195);
nand U18825 (N_18825,N_16319,N_16055);
xor U18826 (N_18826,N_16775,N_16261);
and U18827 (N_18827,N_17802,N_16540);
nor U18828 (N_18828,N_17215,N_16660);
nand U18829 (N_18829,N_16590,N_17991);
nor U18830 (N_18830,N_17879,N_17450);
nand U18831 (N_18831,N_17571,N_17626);
xor U18832 (N_18832,N_17412,N_17289);
nand U18833 (N_18833,N_16128,N_16976);
and U18834 (N_18834,N_17705,N_16345);
nand U18835 (N_18835,N_17131,N_16089);
nor U18836 (N_18836,N_17257,N_17637);
and U18837 (N_18837,N_17796,N_17808);
and U18838 (N_18838,N_16179,N_16981);
nor U18839 (N_18839,N_16030,N_16165);
or U18840 (N_18840,N_17350,N_16452);
and U18841 (N_18841,N_17471,N_17459);
or U18842 (N_18842,N_17116,N_16029);
or U18843 (N_18843,N_16381,N_17646);
nor U18844 (N_18844,N_16638,N_17010);
xor U18845 (N_18845,N_17305,N_17622);
or U18846 (N_18846,N_17541,N_16308);
nand U18847 (N_18847,N_16124,N_16004);
xnor U18848 (N_18848,N_16280,N_16457);
nor U18849 (N_18849,N_16352,N_17063);
and U18850 (N_18850,N_17739,N_17805);
nand U18851 (N_18851,N_17442,N_17003);
nand U18852 (N_18852,N_16378,N_17045);
and U18853 (N_18853,N_17608,N_17902);
nor U18854 (N_18854,N_16703,N_16176);
nor U18855 (N_18855,N_16048,N_17698);
and U18856 (N_18856,N_17499,N_17933);
or U18857 (N_18857,N_17225,N_17124);
nand U18858 (N_18858,N_17276,N_17538);
and U18859 (N_18859,N_17070,N_17301);
or U18860 (N_18860,N_17405,N_17506);
and U18861 (N_18861,N_16097,N_16820);
nand U18862 (N_18862,N_16698,N_16429);
nor U18863 (N_18863,N_17916,N_16213);
or U18864 (N_18864,N_17071,N_17441);
xnor U18865 (N_18865,N_17410,N_17431);
nand U18866 (N_18866,N_17848,N_16360);
or U18867 (N_18867,N_16905,N_16484);
nand U18868 (N_18868,N_16880,N_17981);
nand U18869 (N_18869,N_17722,N_16149);
xnor U18870 (N_18870,N_17989,N_17944);
and U18871 (N_18871,N_17926,N_16785);
nor U18872 (N_18872,N_17773,N_16776);
or U18873 (N_18873,N_17498,N_16731);
nand U18874 (N_18874,N_16025,N_17714);
nor U18875 (N_18875,N_17912,N_17780);
nor U18876 (N_18876,N_17259,N_16350);
nand U18877 (N_18877,N_17822,N_16388);
or U18878 (N_18878,N_17282,N_16926);
and U18879 (N_18879,N_17373,N_17742);
nor U18880 (N_18880,N_16059,N_16327);
nand U18881 (N_18881,N_16551,N_17776);
xor U18882 (N_18882,N_16593,N_17851);
nand U18883 (N_18883,N_16557,N_17865);
xnor U18884 (N_18884,N_17197,N_17386);
nand U18885 (N_18885,N_17542,N_16268);
and U18886 (N_18886,N_17746,N_16547);
nand U18887 (N_18887,N_17938,N_17213);
nand U18888 (N_18888,N_17630,N_16498);
nor U18889 (N_18889,N_16496,N_17363);
xnor U18890 (N_18890,N_16968,N_16719);
nand U18891 (N_18891,N_16410,N_16835);
nor U18892 (N_18892,N_16131,N_17108);
and U18893 (N_18893,N_17717,N_17455);
or U18894 (N_18894,N_17047,N_16729);
nor U18895 (N_18895,N_17402,N_17888);
and U18896 (N_18896,N_17182,N_17712);
nor U18897 (N_18897,N_16628,N_16093);
nor U18898 (N_18898,N_16259,N_16106);
nand U18899 (N_18899,N_16188,N_17663);
nand U18900 (N_18900,N_17710,N_16046);
or U18901 (N_18901,N_16783,N_17110);
and U18902 (N_18902,N_16766,N_16853);
xnor U18903 (N_18903,N_17119,N_17936);
nor U18904 (N_18904,N_17842,N_16598);
nor U18905 (N_18905,N_17617,N_17106);
xor U18906 (N_18906,N_16913,N_17488);
nand U18907 (N_18907,N_16362,N_16216);
nand U18908 (N_18908,N_17076,N_16639);
nor U18909 (N_18909,N_16893,N_16873);
nor U18910 (N_18910,N_16313,N_16717);
nand U18911 (N_18911,N_17274,N_17895);
xnor U18912 (N_18912,N_17647,N_16129);
xor U18913 (N_18913,N_16556,N_16422);
xor U18914 (N_18914,N_16474,N_17686);
nand U18915 (N_18915,N_16644,N_17577);
nand U18916 (N_18916,N_17368,N_17163);
or U18917 (N_18917,N_17143,N_17952);
or U18918 (N_18918,N_17203,N_17243);
nand U18919 (N_18919,N_17873,N_17401);
and U18920 (N_18920,N_16756,N_17783);
nor U18921 (N_18921,N_16070,N_16061);
xor U18922 (N_18922,N_16311,N_16544);
xnor U18923 (N_18923,N_16361,N_16928);
xnor U18924 (N_18924,N_16780,N_17502);
and U18925 (N_18925,N_17961,N_16469);
nor U18926 (N_18926,N_17878,N_17017);
or U18927 (N_18927,N_16648,N_16067);
and U18928 (N_18928,N_17387,N_17104);
or U18929 (N_18929,N_16908,N_17585);
xor U18930 (N_18930,N_16790,N_16874);
xnor U18931 (N_18931,N_16957,N_16285);
and U18932 (N_18932,N_16137,N_16684);
and U18933 (N_18933,N_17367,N_16146);
or U18934 (N_18934,N_16827,N_17158);
and U18935 (N_18935,N_17111,N_17434);
or U18936 (N_18936,N_16501,N_17648);
or U18937 (N_18937,N_17376,N_17721);
or U18938 (N_18938,N_17692,N_17026);
nand U18939 (N_18939,N_17400,N_16306);
nand U18940 (N_18940,N_16045,N_17682);
and U18941 (N_18941,N_17501,N_17769);
nand U18942 (N_18942,N_16943,N_17640);
or U18943 (N_18943,N_17540,N_17294);
xor U18944 (N_18944,N_17846,N_16989);
nand U18945 (N_18945,N_16159,N_16850);
nor U18946 (N_18946,N_16611,N_16816);
xor U18947 (N_18947,N_16687,N_17377);
and U18948 (N_18948,N_16695,N_16842);
and U18949 (N_18949,N_16098,N_17374);
nor U18950 (N_18950,N_17475,N_17667);
or U18951 (N_18951,N_17252,N_17144);
xnor U18952 (N_18952,N_16472,N_16906);
and U18953 (N_18953,N_17168,N_17239);
and U18954 (N_18954,N_17479,N_16187);
xor U18955 (N_18955,N_17246,N_16720);
nand U18956 (N_18956,N_17935,N_17214);
nor U18957 (N_18957,N_16554,N_17324);
nor U18958 (N_18958,N_16221,N_16841);
or U18959 (N_18959,N_16312,N_17534);
nor U18960 (N_18960,N_16520,N_17417);
and U18961 (N_18961,N_16562,N_17346);
nor U18962 (N_18962,N_16079,N_16063);
or U18963 (N_18963,N_17580,N_17574);
xnor U18964 (N_18964,N_16892,N_17706);
xor U18965 (N_18965,N_17084,N_16672);
or U18966 (N_18966,N_17657,N_16156);
xor U18967 (N_18967,N_17631,N_16789);
or U18968 (N_18968,N_17135,N_17759);
xor U18969 (N_18969,N_17133,N_17799);
or U18970 (N_18970,N_17237,N_16666);
nor U18971 (N_18971,N_17381,N_16126);
or U18972 (N_18972,N_16468,N_17897);
or U18973 (N_18973,N_16889,N_17171);
xnor U18974 (N_18974,N_17797,N_17820);
nor U18975 (N_18975,N_16102,N_16254);
xor U18976 (N_18976,N_17743,N_17649);
nor U18977 (N_18977,N_16435,N_17636);
nand U18978 (N_18978,N_16755,N_16040);
nor U18979 (N_18979,N_16604,N_17945);
nand U18980 (N_18980,N_17333,N_17456);
nand U18981 (N_18981,N_16911,N_17795);
nand U18982 (N_18982,N_16830,N_17445);
nor U18983 (N_18983,N_17393,N_17532);
nor U18984 (N_18984,N_16670,N_16798);
xnor U18985 (N_18985,N_17827,N_17828);
xor U18986 (N_18986,N_16101,N_17723);
and U18987 (N_18987,N_17687,N_17185);
nor U18988 (N_18988,N_17012,N_16836);
or U18989 (N_18989,N_17570,N_16076);
xnor U18990 (N_18990,N_17639,N_16355);
xor U18991 (N_18991,N_16184,N_16799);
nand U18992 (N_18992,N_17287,N_16582);
nor U18993 (N_18993,N_17875,N_17980);
xor U18994 (N_18994,N_17838,N_17905);
nor U18995 (N_18995,N_16839,N_16615);
and U18996 (N_18996,N_16758,N_16324);
or U18997 (N_18997,N_16266,N_17793);
nor U18998 (N_18998,N_16826,N_16878);
and U18999 (N_18999,N_17072,N_16330);
and U19000 (N_19000,N_16287,N_16877);
xnor U19001 (N_19001,N_16106,N_17560);
nor U19002 (N_19002,N_17626,N_16699);
and U19003 (N_19003,N_16337,N_17810);
nor U19004 (N_19004,N_16538,N_17241);
and U19005 (N_19005,N_17820,N_17091);
xnor U19006 (N_19006,N_16134,N_17852);
and U19007 (N_19007,N_16144,N_16424);
and U19008 (N_19008,N_17026,N_17162);
or U19009 (N_19009,N_17948,N_16024);
xor U19010 (N_19010,N_16386,N_17764);
nor U19011 (N_19011,N_16740,N_16389);
xor U19012 (N_19012,N_16288,N_16184);
or U19013 (N_19013,N_16254,N_17920);
nor U19014 (N_19014,N_17934,N_16274);
nand U19015 (N_19015,N_17205,N_16615);
and U19016 (N_19016,N_16655,N_17048);
and U19017 (N_19017,N_16466,N_16391);
or U19018 (N_19018,N_16594,N_17500);
nand U19019 (N_19019,N_16914,N_17744);
nand U19020 (N_19020,N_16344,N_16259);
and U19021 (N_19021,N_17019,N_16028);
nor U19022 (N_19022,N_16514,N_17792);
nor U19023 (N_19023,N_17986,N_16570);
and U19024 (N_19024,N_16413,N_16907);
nand U19025 (N_19025,N_17022,N_17614);
and U19026 (N_19026,N_17353,N_16885);
nand U19027 (N_19027,N_17825,N_17255);
or U19028 (N_19028,N_17617,N_16156);
or U19029 (N_19029,N_17134,N_17698);
xor U19030 (N_19030,N_17685,N_16050);
and U19031 (N_19031,N_16479,N_17784);
and U19032 (N_19032,N_17251,N_17847);
or U19033 (N_19033,N_17418,N_16805);
nand U19034 (N_19034,N_16016,N_17910);
or U19035 (N_19035,N_17402,N_17175);
or U19036 (N_19036,N_16771,N_16190);
nor U19037 (N_19037,N_17707,N_17559);
nor U19038 (N_19038,N_16401,N_17739);
and U19039 (N_19039,N_17004,N_16598);
and U19040 (N_19040,N_17625,N_16180);
xnor U19041 (N_19041,N_17537,N_16909);
nor U19042 (N_19042,N_16779,N_16814);
or U19043 (N_19043,N_17113,N_17236);
xnor U19044 (N_19044,N_16303,N_17141);
nand U19045 (N_19045,N_17198,N_17368);
nor U19046 (N_19046,N_17456,N_17316);
and U19047 (N_19047,N_17038,N_16491);
nand U19048 (N_19048,N_17111,N_17733);
or U19049 (N_19049,N_16093,N_16031);
xnor U19050 (N_19050,N_16189,N_16946);
nand U19051 (N_19051,N_16597,N_16718);
or U19052 (N_19052,N_16962,N_17163);
or U19053 (N_19053,N_17466,N_17454);
and U19054 (N_19054,N_17394,N_17096);
or U19055 (N_19055,N_17030,N_17477);
nor U19056 (N_19056,N_16216,N_16693);
nor U19057 (N_19057,N_17510,N_17307);
nor U19058 (N_19058,N_17585,N_16800);
or U19059 (N_19059,N_16008,N_17434);
nor U19060 (N_19060,N_16021,N_17894);
xor U19061 (N_19061,N_17928,N_17673);
nor U19062 (N_19062,N_17993,N_17083);
or U19063 (N_19063,N_16549,N_16222);
and U19064 (N_19064,N_17557,N_16250);
and U19065 (N_19065,N_17079,N_16203);
and U19066 (N_19066,N_17111,N_16202);
and U19067 (N_19067,N_17699,N_17021);
or U19068 (N_19068,N_17308,N_16129);
nor U19069 (N_19069,N_17196,N_16223);
or U19070 (N_19070,N_16805,N_16564);
and U19071 (N_19071,N_16146,N_17178);
xor U19072 (N_19072,N_17715,N_16484);
and U19073 (N_19073,N_16652,N_16856);
and U19074 (N_19074,N_16236,N_16231);
or U19075 (N_19075,N_16158,N_17930);
and U19076 (N_19076,N_17159,N_16454);
or U19077 (N_19077,N_16078,N_16899);
or U19078 (N_19078,N_17668,N_16493);
and U19079 (N_19079,N_16167,N_17134);
and U19080 (N_19080,N_16183,N_16514);
xor U19081 (N_19081,N_16410,N_16328);
or U19082 (N_19082,N_16408,N_17056);
nor U19083 (N_19083,N_16909,N_16605);
nor U19084 (N_19084,N_17141,N_17355);
or U19085 (N_19085,N_16513,N_16925);
and U19086 (N_19086,N_16149,N_16983);
xnor U19087 (N_19087,N_16602,N_16425);
or U19088 (N_19088,N_16396,N_16944);
or U19089 (N_19089,N_16080,N_16321);
nor U19090 (N_19090,N_17228,N_17766);
nor U19091 (N_19091,N_16877,N_17686);
and U19092 (N_19092,N_16618,N_16016);
nor U19093 (N_19093,N_16621,N_16733);
and U19094 (N_19094,N_17921,N_16627);
xor U19095 (N_19095,N_17575,N_17352);
xor U19096 (N_19096,N_16639,N_16097);
nor U19097 (N_19097,N_16735,N_17392);
or U19098 (N_19098,N_16139,N_17777);
nand U19099 (N_19099,N_16792,N_17095);
nand U19100 (N_19100,N_17426,N_16670);
nor U19101 (N_19101,N_17884,N_16556);
nor U19102 (N_19102,N_16421,N_17394);
nor U19103 (N_19103,N_17236,N_16181);
or U19104 (N_19104,N_16628,N_17802);
or U19105 (N_19105,N_16857,N_16482);
xor U19106 (N_19106,N_17429,N_17298);
xor U19107 (N_19107,N_17896,N_17862);
nand U19108 (N_19108,N_17580,N_16498);
or U19109 (N_19109,N_17567,N_17878);
xor U19110 (N_19110,N_17128,N_17164);
or U19111 (N_19111,N_16725,N_17918);
nor U19112 (N_19112,N_16526,N_16692);
xor U19113 (N_19113,N_17984,N_17387);
and U19114 (N_19114,N_17473,N_17458);
nand U19115 (N_19115,N_16312,N_17426);
nand U19116 (N_19116,N_16833,N_17845);
and U19117 (N_19117,N_16829,N_17204);
and U19118 (N_19118,N_16181,N_16183);
or U19119 (N_19119,N_16749,N_17731);
nor U19120 (N_19120,N_17547,N_17358);
nor U19121 (N_19121,N_16566,N_16364);
or U19122 (N_19122,N_16941,N_17214);
or U19123 (N_19123,N_16153,N_17525);
nand U19124 (N_19124,N_17994,N_16674);
and U19125 (N_19125,N_17127,N_16952);
nor U19126 (N_19126,N_17361,N_16824);
or U19127 (N_19127,N_17536,N_17159);
nor U19128 (N_19128,N_17347,N_17939);
xor U19129 (N_19129,N_16019,N_17116);
and U19130 (N_19130,N_16671,N_16646);
xor U19131 (N_19131,N_16433,N_16459);
nand U19132 (N_19132,N_16414,N_16672);
nor U19133 (N_19133,N_17014,N_16479);
nor U19134 (N_19134,N_16213,N_16144);
or U19135 (N_19135,N_16724,N_17622);
nor U19136 (N_19136,N_16084,N_16316);
nor U19137 (N_19137,N_16834,N_16215);
xor U19138 (N_19138,N_16788,N_16118);
and U19139 (N_19139,N_16989,N_16373);
or U19140 (N_19140,N_17581,N_17694);
xnor U19141 (N_19141,N_17847,N_16053);
xor U19142 (N_19142,N_17665,N_17404);
and U19143 (N_19143,N_17750,N_16474);
xor U19144 (N_19144,N_16557,N_17785);
and U19145 (N_19145,N_17923,N_17468);
xnor U19146 (N_19146,N_16807,N_17166);
and U19147 (N_19147,N_17731,N_16862);
and U19148 (N_19148,N_17702,N_16445);
nor U19149 (N_19149,N_16441,N_16972);
xnor U19150 (N_19150,N_17592,N_17713);
nor U19151 (N_19151,N_16742,N_17499);
xor U19152 (N_19152,N_17673,N_16003);
and U19153 (N_19153,N_17775,N_16290);
nor U19154 (N_19154,N_16865,N_17318);
and U19155 (N_19155,N_16582,N_17584);
nor U19156 (N_19156,N_16499,N_16988);
and U19157 (N_19157,N_17086,N_17581);
xnor U19158 (N_19158,N_16279,N_16118);
or U19159 (N_19159,N_16334,N_17934);
and U19160 (N_19160,N_16654,N_16177);
nor U19161 (N_19161,N_16836,N_17431);
nand U19162 (N_19162,N_17838,N_17729);
and U19163 (N_19163,N_17631,N_16276);
nand U19164 (N_19164,N_16239,N_16429);
xor U19165 (N_19165,N_17780,N_17595);
or U19166 (N_19166,N_17483,N_17676);
or U19167 (N_19167,N_17420,N_16438);
nand U19168 (N_19168,N_17213,N_16158);
and U19169 (N_19169,N_17348,N_17316);
and U19170 (N_19170,N_16256,N_17708);
and U19171 (N_19171,N_16505,N_17682);
or U19172 (N_19172,N_17788,N_17780);
nand U19173 (N_19173,N_16462,N_17322);
and U19174 (N_19174,N_16964,N_17209);
nor U19175 (N_19175,N_16411,N_16192);
and U19176 (N_19176,N_16071,N_16301);
or U19177 (N_19177,N_16233,N_17328);
nor U19178 (N_19178,N_17457,N_17468);
nand U19179 (N_19179,N_17993,N_16099);
nor U19180 (N_19180,N_17969,N_16274);
nor U19181 (N_19181,N_17077,N_17920);
nor U19182 (N_19182,N_16669,N_17516);
or U19183 (N_19183,N_17956,N_16449);
or U19184 (N_19184,N_16524,N_17713);
and U19185 (N_19185,N_16445,N_16724);
and U19186 (N_19186,N_17145,N_17225);
nor U19187 (N_19187,N_16620,N_17846);
xnor U19188 (N_19188,N_16841,N_17833);
and U19189 (N_19189,N_16682,N_17403);
nand U19190 (N_19190,N_17315,N_16783);
nor U19191 (N_19191,N_17154,N_16118);
nor U19192 (N_19192,N_17919,N_17806);
xnor U19193 (N_19193,N_16542,N_16405);
nor U19194 (N_19194,N_16320,N_17488);
or U19195 (N_19195,N_16693,N_17635);
and U19196 (N_19196,N_16292,N_17767);
xor U19197 (N_19197,N_16113,N_17134);
nand U19198 (N_19198,N_17648,N_17440);
nand U19199 (N_19199,N_17930,N_16551);
xnor U19200 (N_19200,N_16413,N_17799);
or U19201 (N_19201,N_16745,N_17559);
and U19202 (N_19202,N_16643,N_16095);
or U19203 (N_19203,N_16873,N_17321);
or U19204 (N_19204,N_17006,N_17900);
nand U19205 (N_19205,N_17087,N_17457);
nand U19206 (N_19206,N_17328,N_17965);
nand U19207 (N_19207,N_16950,N_17013);
nand U19208 (N_19208,N_16941,N_16334);
nor U19209 (N_19209,N_17712,N_16634);
nor U19210 (N_19210,N_17711,N_17513);
nor U19211 (N_19211,N_17086,N_17534);
nand U19212 (N_19212,N_16281,N_16484);
or U19213 (N_19213,N_16662,N_16131);
nor U19214 (N_19214,N_17411,N_16303);
nand U19215 (N_19215,N_17863,N_16811);
and U19216 (N_19216,N_17434,N_17341);
and U19217 (N_19217,N_17129,N_17428);
or U19218 (N_19218,N_16333,N_16681);
nor U19219 (N_19219,N_16870,N_16672);
or U19220 (N_19220,N_16848,N_17928);
xnor U19221 (N_19221,N_16586,N_17538);
and U19222 (N_19222,N_17081,N_16170);
and U19223 (N_19223,N_16317,N_16564);
nand U19224 (N_19224,N_16427,N_16304);
nand U19225 (N_19225,N_17912,N_17201);
nand U19226 (N_19226,N_17994,N_17349);
and U19227 (N_19227,N_16193,N_17816);
and U19228 (N_19228,N_16574,N_16078);
nand U19229 (N_19229,N_16134,N_17844);
or U19230 (N_19230,N_17688,N_16331);
and U19231 (N_19231,N_16510,N_17448);
or U19232 (N_19232,N_16951,N_16725);
nor U19233 (N_19233,N_17211,N_17529);
xor U19234 (N_19234,N_17994,N_16739);
xnor U19235 (N_19235,N_17591,N_16357);
and U19236 (N_19236,N_17764,N_17212);
xor U19237 (N_19237,N_16738,N_16469);
or U19238 (N_19238,N_16838,N_16490);
or U19239 (N_19239,N_16297,N_17332);
xnor U19240 (N_19240,N_17027,N_17282);
nand U19241 (N_19241,N_17993,N_16308);
or U19242 (N_19242,N_16829,N_16046);
and U19243 (N_19243,N_17589,N_17770);
xnor U19244 (N_19244,N_17567,N_17459);
and U19245 (N_19245,N_17453,N_16775);
nor U19246 (N_19246,N_16069,N_17173);
xor U19247 (N_19247,N_17976,N_16664);
nor U19248 (N_19248,N_17269,N_16236);
xnor U19249 (N_19249,N_17753,N_17747);
or U19250 (N_19250,N_16479,N_16079);
nor U19251 (N_19251,N_17220,N_16009);
xnor U19252 (N_19252,N_17571,N_17635);
nand U19253 (N_19253,N_16437,N_16605);
nand U19254 (N_19254,N_16852,N_16454);
and U19255 (N_19255,N_17491,N_16409);
nand U19256 (N_19256,N_17721,N_16493);
xnor U19257 (N_19257,N_16967,N_16079);
nand U19258 (N_19258,N_17240,N_17792);
and U19259 (N_19259,N_17618,N_16059);
xor U19260 (N_19260,N_16955,N_17016);
or U19261 (N_19261,N_17194,N_17948);
nor U19262 (N_19262,N_17531,N_16669);
nand U19263 (N_19263,N_17711,N_17305);
or U19264 (N_19264,N_17481,N_17765);
or U19265 (N_19265,N_17384,N_17937);
or U19266 (N_19266,N_16987,N_17589);
and U19267 (N_19267,N_17760,N_16722);
or U19268 (N_19268,N_16540,N_16375);
and U19269 (N_19269,N_17463,N_17687);
and U19270 (N_19270,N_16215,N_16907);
xor U19271 (N_19271,N_17502,N_17943);
xnor U19272 (N_19272,N_17610,N_17671);
or U19273 (N_19273,N_16871,N_16928);
nor U19274 (N_19274,N_17921,N_16124);
nor U19275 (N_19275,N_17207,N_16877);
nand U19276 (N_19276,N_17264,N_16648);
xnor U19277 (N_19277,N_17363,N_17158);
and U19278 (N_19278,N_17633,N_17711);
xnor U19279 (N_19279,N_16334,N_17146);
nor U19280 (N_19280,N_17994,N_16767);
and U19281 (N_19281,N_16915,N_17820);
or U19282 (N_19282,N_16465,N_17902);
xor U19283 (N_19283,N_16511,N_16426);
nand U19284 (N_19284,N_17404,N_16571);
xor U19285 (N_19285,N_17829,N_17483);
or U19286 (N_19286,N_16218,N_17333);
nand U19287 (N_19287,N_17199,N_16287);
or U19288 (N_19288,N_16650,N_16200);
nor U19289 (N_19289,N_17796,N_17464);
and U19290 (N_19290,N_17438,N_17228);
nand U19291 (N_19291,N_17204,N_17869);
nor U19292 (N_19292,N_16043,N_17571);
and U19293 (N_19293,N_17745,N_16623);
xor U19294 (N_19294,N_17763,N_17699);
nor U19295 (N_19295,N_17688,N_16701);
and U19296 (N_19296,N_16475,N_17611);
or U19297 (N_19297,N_16044,N_16482);
nor U19298 (N_19298,N_17711,N_17470);
and U19299 (N_19299,N_17735,N_16841);
xnor U19300 (N_19300,N_17043,N_16664);
or U19301 (N_19301,N_16077,N_17889);
or U19302 (N_19302,N_17322,N_17418);
or U19303 (N_19303,N_16864,N_16187);
xor U19304 (N_19304,N_17078,N_16209);
or U19305 (N_19305,N_16505,N_16503);
nand U19306 (N_19306,N_17154,N_16497);
or U19307 (N_19307,N_17234,N_16499);
nor U19308 (N_19308,N_16903,N_17307);
nand U19309 (N_19309,N_16982,N_16734);
or U19310 (N_19310,N_16598,N_16117);
nor U19311 (N_19311,N_17292,N_17374);
or U19312 (N_19312,N_16879,N_17342);
and U19313 (N_19313,N_16120,N_17899);
xnor U19314 (N_19314,N_17546,N_16213);
nor U19315 (N_19315,N_16945,N_17537);
nand U19316 (N_19316,N_17202,N_16796);
xor U19317 (N_19317,N_16840,N_17978);
xor U19318 (N_19318,N_16432,N_16285);
or U19319 (N_19319,N_17875,N_16467);
xnor U19320 (N_19320,N_17863,N_16779);
nor U19321 (N_19321,N_17311,N_16871);
nor U19322 (N_19322,N_16786,N_16716);
nand U19323 (N_19323,N_16648,N_17837);
nor U19324 (N_19324,N_17224,N_16900);
xnor U19325 (N_19325,N_16829,N_16355);
nor U19326 (N_19326,N_17613,N_16854);
nor U19327 (N_19327,N_16850,N_17063);
or U19328 (N_19328,N_17264,N_17332);
nand U19329 (N_19329,N_17023,N_17758);
and U19330 (N_19330,N_17087,N_17244);
nand U19331 (N_19331,N_17945,N_17873);
or U19332 (N_19332,N_16740,N_16441);
or U19333 (N_19333,N_17870,N_16452);
and U19334 (N_19334,N_17377,N_17433);
and U19335 (N_19335,N_16465,N_17856);
and U19336 (N_19336,N_16992,N_17390);
xor U19337 (N_19337,N_16793,N_16138);
nand U19338 (N_19338,N_16031,N_17052);
or U19339 (N_19339,N_17631,N_16768);
xor U19340 (N_19340,N_16532,N_16911);
nor U19341 (N_19341,N_17911,N_16660);
or U19342 (N_19342,N_16295,N_16277);
or U19343 (N_19343,N_17408,N_16275);
nand U19344 (N_19344,N_16689,N_17182);
and U19345 (N_19345,N_17980,N_16853);
nand U19346 (N_19346,N_16607,N_17110);
nor U19347 (N_19347,N_16988,N_17674);
nand U19348 (N_19348,N_17011,N_16624);
nor U19349 (N_19349,N_16874,N_17478);
nor U19350 (N_19350,N_16875,N_16153);
and U19351 (N_19351,N_16343,N_17104);
nand U19352 (N_19352,N_16588,N_16960);
and U19353 (N_19353,N_16157,N_17783);
and U19354 (N_19354,N_17008,N_16648);
xnor U19355 (N_19355,N_17149,N_16434);
nand U19356 (N_19356,N_17278,N_17988);
nor U19357 (N_19357,N_17244,N_16715);
nand U19358 (N_19358,N_16636,N_17693);
nor U19359 (N_19359,N_17994,N_17005);
xnor U19360 (N_19360,N_17752,N_17692);
and U19361 (N_19361,N_16025,N_16318);
or U19362 (N_19362,N_16652,N_17837);
xor U19363 (N_19363,N_17582,N_17449);
and U19364 (N_19364,N_16132,N_16762);
nor U19365 (N_19365,N_17094,N_17389);
xnor U19366 (N_19366,N_17697,N_16934);
nand U19367 (N_19367,N_17773,N_16762);
nand U19368 (N_19368,N_16336,N_17906);
nand U19369 (N_19369,N_16549,N_17168);
and U19370 (N_19370,N_17356,N_16386);
xnor U19371 (N_19371,N_17967,N_17794);
xor U19372 (N_19372,N_17797,N_16798);
nand U19373 (N_19373,N_17306,N_16381);
nand U19374 (N_19374,N_17200,N_16464);
or U19375 (N_19375,N_16385,N_17916);
xnor U19376 (N_19376,N_17000,N_17388);
xnor U19377 (N_19377,N_16484,N_16374);
xnor U19378 (N_19378,N_16109,N_16725);
or U19379 (N_19379,N_17012,N_16693);
and U19380 (N_19380,N_16514,N_16203);
xor U19381 (N_19381,N_17422,N_16956);
xor U19382 (N_19382,N_16684,N_17803);
xnor U19383 (N_19383,N_17382,N_16986);
xnor U19384 (N_19384,N_16679,N_16064);
nor U19385 (N_19385,N_17586,N_17144);
xnor U19386 (N_19386,N_17073,N_17087);
nand U19387 (N_19387,N_16543,N_16284);
and U19388 (N_19388,N_17157,N_17489);
and U19389 (N_19389,N_17541,N_17068);
xnor U19390 (N_19390,N_17731,N_17915);
xor U19391 (N_19391,N_16665,N_17477);
and U19392 (N_19392,N_17461,N_17839);
and U19393 (N_19393,N_16336,N_16182);
or U19394 (N_19394,N_17101,N_16436);
xor U19395 (N_19395,N_17861,N_17790);
nand U19396 (N_19396,N_17023,N_17335);
or U19397 (N_19397,N_17857,N_16399);
nor U19398 (N_19398,N_16694,N_17159);
xnor U19399 (N_19399,N_17473,N_16966);
nand U19400 (N_19400,N_17068,N_17920);
nor U19401 (N_19401,N_17957,N_17444);
nor U19402 (N_19402,N_16996,N_16584);
nand U19403 (N_19403,N_16619,N_17355);
xor U19404 (N_19404,N_16260,N_16228);
and U19405 (N_19405,N_16144,N_17460);
nand U19406 (N_19406,N_17405,N_16678);
and U19407 (N_19407,N_17852,N_16065);
nor U19408 (N_19408,N_16510,N_17462);
nand U19409 (N_19409,N_17678,N_16184);
and U19410 (N_19410,N_16075,N_16496);
and U19411 (N_19411,N_17540,N_17853);
nand U19412 (N_19412,N_17484,N_17622);
nor U19413 (N_19413,N_16464,N_16687);
and U19414 (N_19414,N_17225,N_17311);
nor U19415 (N_19415,N_17532,N_16661);
nor U19416 (N_19416,N_17826,N_17969);
xor U19417 (N_19417,N_17894,N_17923);
xnor U19418 (N_19418,N_16794,N_17469);
or U19419 (N_19419,N_17864,N_17085);
nand U19420 (N_19420,N_16022,N_16510);
xnor U19421 (N_19421,N_16037,N_17560);
and U19422 (N_19422,N_16405,N_17155);
and U19423 (N_19423,N_17295,N_17305);
xor U19424 (N_19424,N_17701,N_17770);
and U19425 (N_19425,N_17117,N_16211);
xnor U19426 (N_19426,N_17096,N_16340);
xor U19427 (N_19427,N_17201,N_16009);
or U19428 (N_19428,N_16215,N_17314);
or U19429 (N_19429,N_17366,N_17746);
or U19430 (N_19430,N_16737,N_17795);
nor U19431 (N_19431,N_17133,N_16226);
xor U19432 (N_19432,N_16245,N_16895);
nand U19433 (N_19433,N_16435,N_17051);
and U19434 (N_19434,N_16663,N_17709);
nand U19435 (N_19435,N_17762,N_17489);
nand U19436 (N_19436,N_17386,N_16841);
or U19437 (N_19437,N_16474,N_17407);
and U19438 (N_19438,N_17372,N_16219);
nand U19439 (N_19439,N_17631,N_16227);
and U19440 (N_19440,N_17133,N_17955);
nand U19441 (N_19441,N_16512,N_16596);
xnor U19442 (N_19442,N_17731,N_17657);
xnor U19443 (N_19443,N_17121,N_17226);
or U19444 (N_19444,N_17319,N_17998);
and U19445 (N_19445,N_16782,N_16993);
and U19446 (N_19446,N_17093,N_17764);
nor U19447 (N_19447,N_16246,N_17689);
nand U19448 (N_19448,N_16091,N_17910);
xor U19449 (N_19449,N_17996,N_17429);
nand U19450 (N_19450,N_17437,N_16730);
xor U19451 (N_19451,N_16607,N_16878);
or U19452 (N_19452,N_16199,N_17905);
nand U19453 (N_19453,N_16004,N_17721);
and U19454 (N_19454,N_17982,N_17165);
and U19455 (N_19455,N_16051,N_16747);
or U19456 (N_19456,N_17159,N_17145);
nand U19457 (N_19457,N_16265,N_17950);
or U19458 (N_19458,N_17194,N_17499);
and U19459 (N_19459,N_17013,N_16668);
xnor U19460 (N_19460,N_17797,N_16454);
nor U19461 (N_19461,N_17901,N_17207);
xnor U19462 (N_19462,N_17618,N_16757);
xnor U19463 (N_19463,N_17216,N_17780);
nand U19464 (N_19464,N_17210,N_17827);
nor U19465 (N_19465,N_17638,N_17496);
xor U19466 (N_19466,N_17793,N_16469);
xnor U19467 (N_19467,N_16360,N_17551);
xnor U19468 (N_19468,N_17853,N_16445);
and U19469 (N_19469,N_16336,N_17223);
xnor U19470 (N_19470,N_17110,N_16818);
nand U19471 (N_19471,N_17764,N_16884);
nand U19472 (N_19472,N_17776,N_16418);
or U19473 (N_19473,N_17677,N_17157);
nand U19474 (N_19474,N_17316,N_17713);
or U19475 (N_19475,N_16448,N_17244);
xnor U19476 (N_19476,N_16859,N_16535);
or U19477 (N_19477,N_17312,N_17919);
and U19478 (N_19478,N_17431,N_17842);
nor U19479 (N_19479,N_17917,N_17816);
nor U19480 (N_19480,N_16312,N_17767);
or U19481 (N_19481,N_16084,N_17699);
nand U19482 (N_19482,N_16124,N_17467);
or U19483 (N_19483,N_17718,N_16601);
or U19484 (N_19484,N_17733,N_16613);
nand U19485 (N_19485,N_16661,N_16742);
nand U19486 (N_19486,N_16583,N_16202);
nand U19487 (N_19487,N_16614,N_16601);
nor U19488 (N_19488,N_16573,N_17706);
and U19489 (N_19489,N_16967,N_16398);
or U19490 (N_19490,N_16713,N_16890);
or U19491 (N_19491,N_17264,N_17719);
and U19492 (N_19492,N_17657,N_17221);
xnor U19493 (N_19493,N_17006,N_17296);
or U19494 (N_19494,N_17811,N_16835);
or U19495 (N_19495,N_17305,N_16115);
nor U19496 (N_19496,N_16857,N_16794);
and U19497 (N_19497,N_17076,N_16836);
nand U19498 (N_19498,N_17691,N_17163);
nand U19499 (N_19499,N_16631,N_16010);
nand U19500 (N_19500,N_17820,N_17808);
or U19501 (N_19501,N_17770,N_16335);
nand U19502 (N_19502,N_17913,N_16451);
and U19503 (N_19503,N_17747,N_16645);
and U19504 (N_19504,N_16279,N_17406);
xor U19505 (N_19505,N_16630,N_17783);
nor U19506 (N_19506,N_16787,N_16305);
or U19507 (N_19507,N_16662,N_17159);
xor U19508 (N_19508,N_16641,N_16860);
and U19509 (N_19509,N_17455,N_16560);
or U19510 (N_19510,N_16233,N_17704);
or U19511 (N_19511,N_16871,N_17796);
or U19512 (N_19512,N_16581,N_17944);
xor U19513 (N_19513,N_17738,N_17422);
and U19514 (N_19514,N_17852,N_16727);
xnor U19515 (N_19515,N_17608,N_17518);
nor U19516 (N_19516,N_17913,N_16267);
nand U19517 (N_19517,N_16634,N_17883);
nand U19518 (N_19518,N_16491,N_17481);
nor U19519 (N_19519,N_16040,N_17495);
or U19520 (N_19520,N_17744,N_17116);
and U19521 (N_19521,N_16289,N_16593);
nand U19522 (N_19522,N_16060,N_16284);
xor U19523 (N_19523,N_16010,N_17375);
xor U19524 (N_19524,N_17851,N_17596);
nor U19525 (N_19525,N_16184,N_17600);
nor U19526 (N_19526,N_16380,N_17614);
nand U19527 (N_19527,N_17835,N_17879);
or U19528 (N_19528,N_16844,N_16139);
nand U19529 (N_19529,N_17765,N_17444);
nand U19530 (N_19530,N_17508,N_17380);
and U19531 (N_19531,N_16753,N_17903);
or U19532 (N_19532,N_17466,N_16553);
nand U19533 (N_19533,N_16858,N_17282);
nand U19534 (N_19534,N_17509,N_16571);
nor U19535 (N_19535,N_16637,N_17370);
xnor U19536 (N_19536,N_16291,N_16089);
nand U19537 (N_19537,N_16836,N_17436);
xnor U19538 (N_19538,N_17964,N_16791);
nor U19539 (N_19539,N_16504,N_16905);
or U19540 (N_19540,N_17989,N_17156);
and U19541 (N_19541,N_17802,N_17102);
xor U19542 (N_19542,N_16395,N_16612);
and U19543 (N_19543,N_17309,N_17020);
nor U19544 (N_19544,N_17653,N_16684);
and U19545 (N_19545,N_16930,N_16911);
and U19546 (N_19546,N_17976,N_17995);
and U19547 (N_19547,N_16758,N_17904);
xnor U19548 (N_19548,N_16760,N_16996);
or U19549 (N_19549,N_16275,N_16059);
or U19550 (N_19550,N_17342,N_17758);
or U19551 (N_19551,N_16096,N_17250);
and U19552 (N_19552,N_16895,N_16278);
or U19553 (N_19553,N_17697,N_16176);
or U19554 (N_19554,N_16189,N_16778);
nand U19555 (N_19555,N_17084,N_16440);
xnor U19556 (N_19556,N_17486,N_17078);
nand U19557 (N_19557,N_17354,N_17538);
and U19558 (N_19558,N_16110,N_17680);
nor U19559 (N_19559,N_17682,N_16935);
nor U19560 (N_19560,N_17040,N_16389);
nand U19561 (N_19561,N_17547,N_16753);
and U19562 (N_19562,N_17932,N_17812);
or U19563 (N_19563,N_17259,N_17201);
xnor U19564 (N_19564,N_16276,N_16656);
or U19565 (N_19565,N_17192,N_16496);
nor U19566 (N_19566,N_16713,N_16593);
or U19567 (N_19567,N_17780,N_17929);
or U19568 (N_19568,N_16277,N_16207);
xnor U19569 (N_19569,N_16602,N_16178);
nand U19570 (N_19570,N_16766,N_16654);
or U19571 (N_19571,N_17537,N_17881);
or U19572 (N_19572,N_16731,N_17509);
nand U19573 (N_19573,N_17432,N_17759);
or U19574 (N_19574,N_16190,N_17302);
or U19575 (N_19575,N_17439,N_17257);
and U19576 (N_19576,N_17972,N_17400);
and U19577 (N_19577,N_16201,N_16640);
and U19578 (N_19578,N_17991,N_16661);
nor U19579 (N_19579,N_17464,N_17553);
nand U19580 (N_19580,N_16408,N_16417);
nor U19581 (N_19581,N_17688,N_17368);
xor U19582 (N_19582,N_17186,N_16941);
and U19583 (N_19583,N_17194,N_16804);
or U19584 (N_19584,N_17251,N_16603);
xnor U19585 (N_19585,N_16052,N_16042);
nor U19586 (N_19586,N_16285,N_16294);
nand U19587 (N_19587,N_17664,N_17250);
or U19588 (N_19588,N_16601,N_17752);
xnor U19589 (N_19589,N_17132,N_17321);
or U19590 (N_19590,N_16232,N_17855);
or U19591 (N_19591,N_17683,N_16059);
xor U19592 (N_19592,N_16800,N_17940);
xor U19593 (N_19593,N_17759,N_17587);
nor U19594 (N_19594,N_17625,N_16654);
nand U19595 (N_19595,N_17523,N_16140);
nand U19596 (N_19596,N_17994,N_16098);
nor U19597 (N_19597,N_16611,N_16971);
xnor U19598 (N_19598,N_16438,N_16303);
nand U19599 (N_19599,N_16083,N_17762);
xor U19600 (N_19600,N_17109,N_16497);
xor U19601 (N_19601,N_16636,N_17193);
xor U19602 (N_19602,N_17356,N_17947);
nor U19603 (N_19603,N_17338,N_16948);
and U19604 (N_19604,N_16182,N_16826);
and U19605 (N_19605,N_17412,N_16197);
or U19606 (N_19606,N_16137,N_16389);
xor U19607 (N_19607,N_16761,N_17043);
nand U19608 (N_19608,N_17601,N_16011);
nor U19609 (N_19609,N_16073,N_17595);
and U19610 (N_19610,N_17105,N_16816);
nor U19611 (N_19611,N_16714,N_17437);
nor U19612 (N_19612,N_16920,N_16043);
xor U19613 (N_19613,N_17562,N_16705);
and U19614 (N_19614,N_17323,N_16351);
xnor U19615 (N_19615,N_16703,N_17949);
xnor U19616 (N_19616,N_17150,N_17265);
nor U19617 (N_19617,N_17891,N_17550);
and U19618 (N_19618,N_16268,N_16143);
or U19619 (N_19619,N_17502,N_16808);
or U19620 (N_19620,N_17873,N_16534);
or U19621 (N_19621,N_17950,N_16224);
nand U19622 (N_19622,N_16531,N_16901);
nor U19623 (N_19623,N_16688,N_16842);
xnor U19624 (N_19624,N_17603,N_16542);
nor U19625 (N_19625,N_17155,N_16233);
or U19626 (N_19626,N_17235,N_17234);
nand U19627 (N_19627,N_16072,N_16243);
or U19628 (N_19628,N_16684,N_17377);
nand U19629 (N_19629,N_17881,N_16384);
xor U19630 (N_19630,N_16962,N_16475);
nor U19631 (N_19631,N_17786,N_17805);
nand U19632 (N_19632,N_16124,N_16895);
and U19633 (N_19633,N_16955,N_16972);
nand U19634 (N_19634,N_17203,N_16924);
or U19635 (N_19635,N_16580,N_17171);
xnor U19636 (N_19636,N_16997,N_16191);
nor U19637 (N_19637,N_17088,N_16418);
nand U19638 (N_19638,N_16570,N_16602);
xnor U19639 (N_19639,N_17446,N_17407);
xnor U19640 (N_19640,N_16882,N_17872);
nor U19641 (N_19641,N_17912,N_16412);
or U19642 (N_19642,N_17526,N_16057);
nand U19643 (N_19643,N_16272,N_16457);
nand U19644 (N_19644,N_16057,N_17746);
or U19645 (N_19645,N_16390,N_16594);
or U19646 (N_19646,N_16163,N_17384);
nor U19647 (N_19647,N_16158,N_17172);
nand U19648 (N_19648,N_17994,N_17703);
nor U19649 (N_19649,N_17469,N_16997);
xor U19650 (N_19650,N_17350,N_17039);
xnor U19651 (N_19651,N_17751,N_16691);
and U19652 (N_19652,N_16711,N_16972);
nand U19653 (N_19653,N_17889,N_17509);
and U19654 (N_19654,N_17501,N_17033);
nor U19655 (N_19655,N_16138,N_17085);
nor U19656 (N_19656,N_17201,N_17268);
and U19657 (N_19657,N_17841,N_17271);
nand U19658 (N_19658,N_16570,N_17216);
nand U19659 (N_19659,N_16215,N_16860);
or U19660 (N_19660,N_16678,N_16759);
and U19661 (N_19661,N_17765,N_16237);
xnor U19662 (N_19662,N_16921,N_17639);
or U19663 (N_19663,N_17755,N_16595);
nand U19664 (N_19664,N_17353,N_17416);
xnor U19665 (N_19665,N_16033,N_17116);
nand U19666 (N_19666,N_16941,N_17542);
and U19667 (N_19667,N_17155,N_16018);
nand U19668 (N_19668,N_16907,N_17125);
or U19669 (N_19669,N_17542,N_16924);
nand U19670 (N_19670,N_17096,N_17355);
or U19671 (N_19671,N_17834,N_16978);
and U19672 (N_19672,N_16117,N_17900);
nand U19673 (N_19673,N_16270,N_16440);
nand U19674 (N_19674,N_17887,N_16469);
or U19675 (N_19675,N_17304,N_16111);
nor U19676 (N_19676,N_16174,N_16993);
or U19677 (N_19677,N_17876,N_17151);
or U19678 (N_19678,N_16835,N_16195);
nor U19679 (N_19679,N_17492,N_17059);
xor U19680 (N_19680,N_17073,N_16655);
nor U19681 (N_19681,N_16316,N_16909);
nand U19682 (N_19682,N_16238,N_17801);
xor U19683 (N_19683,N_16390,N_16455);
and U19684 (N_19684,N_17275,N_17763);
and U19685 (N_19685,N_17198,N_16070);
and U19686 (N_19686,N_17655,N_17599);
or U19687 (N_19687,N_16903,N_16297);
nor U19688 (N_19688,N_16635,N_17487);
and U19689 (N_19689,N_17563,N_17485);
or U19690 (N_19690,N_17076,N_16886);
and U19691 (N_19691,N_17322,N_17119);
and U19692 (N_19692,N_17487,N_16349);
and U19693 (N_19693,N_16243,N_17992);
and U19694 (N_19694,N_17501,N_16809);
and U19695 (N_19695,N_17490,N_16080);
nand U19696 (N_19696,N_17210,N_16687);
and U19697 (N_19697,N_17789,N_16225);
and U19698 (N_19698,N_16254,N_16688);
or U19699 (N_19699,N_17689,N_17588);
nand U19700 (N_19700,N_17965,N_16072);
and U19701 (N_19701,N_16378,N_17858);
nor U19702 (N_19702,N_17019,N_16129);
or U19703 (N_19703,N_16145,N_16507);
nand U19704 (N_19704,N_17384,N_17842);
nand U19705 (N_19705,N_17107,N_17839);
or U19706 (N_19706,N_17592,N_16345);
or U19707 (N_19707,N_17623,N_16379);
nor U19708 (N_19708,N_17048,N_16116);
or U19709 (N_19709,N_17539,N_17738);
and U19710 (N_19710,N_17603,N_16858);
nor U19711 (N_19711,N_16422,N_17289);
or U19712 (N_19712,N_16827,N_17999);
nor U19713 (N_19713,N_17270,N_16043);
xor U19714 (N_19714,N_16918,N_16916);
nand U19715 (N_19715,N_16909,N_17825);
nand U19716 (N_19716,N_16545,N_17381);
xor U19717 (N_19717,N_17763,N_16127);
xnor U19718 (N_19718,N_16205,N_17856);
nor U19719 (N_19719,N_17612,N_16937);
xnor U19720 (N_19720,N_16569,N_16321);
nand U19721 (N_19721,N_17295,N_17567);
nor U19722 (N_19722,N_17831,N_17592);
xnor U19723 (N_19723,N_16758,N_17499);
nor U19724 (N_19724,N_17468,N_17427);
nand U19725 (N_19725,N_16968,N_16035);
and U19726 (N_19726,N_16418,N_16275);
and U19727 (N_19727,N_16231,N_16967);
nand U19728 (N_19728,N_16787,N_16532);
and U19729 (N_19729,N_17658,N_16543);
nor U19730 (N_19730,N_17099,N_16197);
and U19731 (N_19731,N_16830,N_17286);
xor U19732 (N_19732,N_17479,N_17524);
or U19733 (N_19733,N_17308,N_16752);
xnor U19734 (N_19734,N_17704,N_16945);
xor U19735 (N_19735,N_17294,N_16951);
or U19736 (N_19736,N_16928,N_16015);
xor U19737 (N_19737,N_16315,N_16680);
xor U19738 (N_19738,N_16183,N_16939);
nand U19739 (N_19739,N_16473,N_16971);
and U19740 (N_19740,N_16016,N_17864);
or U19741 (N_19741,N_17280,N_16373);
nor U19742 (N_19742,N_16455,N_17257);
and U19743 (N_19743,N_16713,N_16461);
and U19744 (N_19744,N_17307,N_17605);
and U19745 (N_19745,N_17754,N_16605);
nand U19746 (N_19746,N_17099,N_16198);
or U19747 (N_19747,N_16548,N_17007);
xnor U19748 (N_19748,N_16405,N_16241);
xnor U19749 (N_19749,N_17461,N_17558);
xor U19750 (N_19750,N_17019,N_16719);
nor U19751 (N_19751,N_17112,N_16866);
nor U19752 (N_19752,N_17025,N_16808);
xnor U19753 (N_19753,N_17201,N_16438);
xor U19754 (N_19754,N_16800,N_16583);
and U19755 (N_19755,N_17831,N_17501);
xnor U19756 (N_19756,N_17156,N_16315);
and U19757 (N_19757,N_16102,N_17868);
and U19758 (N_19758,N_16748,N_16687);
or U19759 (N_19759,N_16688,N_16848);
or U19760 (N_19760,N_17041,N_17019);
xor U19761 (N_19761,N_17966,N_16590);
nand U19762 (N_19762,N_17479,N_17188);
or U19763 (N_19763,N_16733,N_17436);
xnor U19764 (N_19764,N_17763,N_17429);
nor U19765 (N_19765,N_17031,N_17630);
nand U19766 (N_19766,N_16986,N_16940);
xor U19767 (N_19767,N_16562,N_16441);
nor U19768 (N_19768,N_16523,N_16339);
nor U19769 (N_19769,N_17864,N_17475);
xor U19770 (N_19770,N_16040,N_17579);
or U19771 (N_19771,N_17917,N_17653);
and U19772 (N_19772,N_16816,N_17938);
or U19773 (N_19773,N_17190,N_17842);
nor U19774 (N_19774,N_16196,N_17760);
and U19775 (N_19775,N_17869,N_17298);
or U19776 (N_19776,N_17525,N_17531);
nand U19777 (N_19777,N_17354,N_16793);
and U19778 (N_19778,N_17775,N_16663);
or U19779 (N_19779,N_16297,N_16536);
or U19780 (N_19780,N_16356,N_17442);
nor U19781 (N_19781,N_17888,N_16392);
nand U19782 (N_19782,N_17947,N_17251);
and U19783 (N_19783,N_16512,N_16966);
nand U19784 (N_19784,N_17122,N_17045);
nand U19785 (N_19785,N_16310,N_16452);
and U19786 (N_19786,N_16590,N_16186);
xor U19787 (N_19787,N_17721,N_16487);
nand U19788 (N_19788,N_17508,N_16019);
and U19789 (N_19789,N_16000,N_17085);
nand U19790 (N_19790,N_17199,N_17132);
and U19791 (N_19791,N_16230,N_17028);
nor U19792 (N_19792,N_16890,N_16555);
nor U19793 (N_19793,N_16437,N_17131);
nand U19794 (N_19794,N_17861,N_17691);
nor U19795 (N_19795,N_17330,N_16769);
nor U19796 (N_19796,N_17166,N_16056);
and U19797 (N_19797,N_17808,N_17077);
and U19798 (N_19798,N_17598,N_17987);
or U19799 (N_19799,N_17363,N_16641);
and U19800 (N_19800,N_16828,N_17009);
nand U19801 (N_19801,N_17222,N_17180);
nor U19802 (N_19802,N_17744,N_17280);
nand U19803 (N_19803,N_16722,N_17106);
and U19804 (N_19804,N_17202,N_16828);
and U19805 (N_19805,N_17232,N_17679);
nand U19806 (N_19806,N_16100,N_16393);
nor U19807 (N_19807,N_16306,N_16995);
or U19808 (N_19808,N_17884,N_16224);
nand U19809 (N_19809,N_16631,N_16820);
or U19810 (N_19810,N_16613,N_16754);
xnor U19811 (N_19811,N_17252,N_17303);
xor U19812 (N_19812,N_17637,N_16213);
and U19813 (N_19813,N_16267,N_17470);
nand U19814 (N_19814,N_17070,N_16140);
or U19815 (N_19815,N_17944,N_17595);
xor U19816 (N_19816,N_16970,N_17653);
nor U19817 (N_19817,N_17192,N_16041);
nor U19818 (N_19818,N_17557,N_16733);
and U19819 (N_19819,N_17125,N_16200);
xnor U19820 (N_19820,N_16760,N_16293);
and U19821 (N_19821,N_16908,N_16429);
xor U19822 (N_19822,N_17098,N_16591);
xnor U19823 (N_19823,N_16468,N_17863);
xnor U19824 (N_19824,N_17460,N_16827);
nand U19825 (N_19825,N_16188,N_17430);
nand U19826 (N_19826,N_17440,N_16110);
nand U19827 (N_19827,N_16809,N_17527);
xor U19828 (N_19828,N_17014,N_16049);
xnor U19829 (N_19829,N_16085,N_16112);
and U19830 (N_19830,N_16298,N_16460);
xor U19831 (N_19831,N_16947,N_17725);
xor U19832 (N_19832,N_17082,N_17654);
nand U19833 (N_19833,N_17616,N_16952);
nor U19834 (N_19834,N_17203,N_17883);
nand U19835 (N_19835,N_16132,N_17752);
xnor U19836 (N_19836,N_16708,N_17195);
xnor U19837 (N_19837,N_17136,N_17963);
nor U19838 (N_19838,N_17522,N_17162);
or U19839 (N_19839,N_16856,N_17352);
nor U19840 (N_19840,N_16042,N_17733);
nand U19841 (N_19841,N_17173,N_17732);
and U19842 (N_19842,N_16232,N_16047);
nor U19843 (N_19843,N_17917,N_17275);
nand U19844 (N_19844,N_16798,N_17018);
nor U19845 (N_19845,N_16980,N_17907);
xnor U19846 (N_19846,N_16580,N_16759);
or U19847 (N_19847,N_17744,N_17940);
nor U19848 (N_19848,N_17721,N_17437);
nand U19849 (N_19849,N_17525,N_16841);
and U19850 (N_19850,N_16027,N_16769);
xnor U19851 (N_19851,N_17116,N_17691);
nor U19852 (N_19852,N_17182,N_17725);
and U19853 (N_19853,N_16588,N_17812);
or U19854 (N_19854,N_17419,N_16660);
or U19855 (N_19855,N_16464,N_17546);
and U19856 (N_19856,N_16835,N_16883);
xnor U19857 (N_19857,N_16950,N_16175);
or U19858 (N_19858,N_16105,N_16799);
and U19859 (N_19859,N_16317,N_16536);
nand U19860 (N_19860,N_17681,N_17160);
xor U19861 (N_19861,N_16913,N_16426);
xor U19862 (N_19862,N_16937,N_17818);
nor U19863 (N_19863,N_17711,N_17186);
xor U19864 (N_19864,N_17871,N_16283);
xor U19865 (N_19865,N_17808,N_17973);
xor U19866 (N_19866,N_17409,N_17827);
nor U19867 (N_19867,N_17282,N_16209);
nand U19868 (N_19868,N_17054,N_16719);
or U19869 (N_19869,N_16066,N_16972);
or U19870 (N_19870,N_17876,N_17966);
nor U19871 (N_19871,N_17951,N_16139);
xnor U19872 (N_19872,N_16309,N_16056);
nor U19873 (N_19873,N_16166,N_17466);
nand U19874 (N_19874,N_16987,N_17490);
nand U19875 (N_19875,N_16860,N_17839);
nand U19876 (N_19876,N_17622,N_16133);
xor U19877 (N_19877,N_16001,N_16358);
xnor U19878 (N_19878,N_16236,N_17064);
nand U19879 (N_19879,N_17835,N_17344);
xor U19880 (N_19880,N_17418,N_16003);
and U19881 (N_19881,N_17758,N_16642);
nand U19882 (N_19882,N_17118,N_17539);
or U19883 (N_19883,N_16088,N_17917);
nor U19884 (N_19884,N_16017,N_16551);
xnor U19885 (N_19885,N_16503,N_16804);
nand U19886 (N_19886,N_17365,N_16104);
and U19887 (N_19887,N_16374,N_17084);
and U19888 (N_19888,N_17514,N_16727);
nor U19889 (N_19889,N_17888,N_16503);
or U19890 (N_19890,N_16066,N_17616);
or U19891 (N_19891,N_17544,N_16541);
or U19892 (N_19892,N_17123,N_16932);
and U19893 (N_19893,N_16006,N_16869);
and U19894 (N_19894,N_16458,N_16659);
or U19895 (N_19895,N_17995,N_16187);
xor U19896 (N_19896,N_17842,N_16533);
and U19897 (N_19897,N_17771,N_16969);
nor U19898 (N_19898,N_17822,N_16360);
nand U19899 (N_19899,N_16984,N_17890);
nand U19900 (N_19900,N_17045,N_17418);
and U19901 (N_19901,N_16759,N_16526);
and U19902 (N_19902,N_17215,N_17937);
or U19903 (N_19903,N_16309,N_16341);
and U19904 (N_19904,N_16383,N_16484);
nand U19905 (N_19905,N_16904,N_16432);
nand U19906 (N_19906,N_17519,N_16211);
nor U19907 (N_19907,N_16891,N_16191);
nand U19908 (N_19908,N_16359,N_16604);
xnor U19909 (N_19909,N_16846,N_17599);
nor U19910 (N_19910,N_16164,N_17662);
nor U19911 (N_19911,N_16309,N_16242);
xor U19912 (N_19912,N_17124,N_17715);
xnor U19913 (N_19913,N_16282,N_17715);
nand U19914 (N_19914,N_16434,N_16303);
and U19915 (N_19915,N_17964,N_17631);
or U19916 (N_19916,N_16770,N_17826);
xnor U19917 (N_19917,N_16147,N_17098);
nor U19918 (N_19918,N_16230,N_17835);
xnor U19919 (N_19919,N_16641,N_16527);
xnor U19920 (N_19920,N_17410,N_16302);
nor U19921 (N_19921,N_16031,N_17259);
xor U19922 (N_19922,N_16987,N_16539);
and U19923 (N_19923,N_16576,N_16588);
nand U19924 (N_19924,N_16969,N_17294);
nand U19925 (N_19925,N_16583,N_16899);
nor U19926 (N_19926,N_16427,N_16011);
or U19927 (N_19927,N_17389,N_16853);
nor U19928 (N_19928,N_17413,N_16247);
xor U19929 (N_19929,N_17694,N_16227);
nor U19930 (N_19930,N_16390,N_16690);
or U19931 (N_19931,N_17294,N_17188);
xnor U19932 (N_19932,N_17284,N_17492);
or U19933 (N_19933,N_17579,N_16502);
nor U19934 (N_19934,N_16008,N_16884);
and U19935 (N_19935,N_16983,N_16546);
xnor U19936 (N_19936,N_17036,N_16143);
nand U19937 (N_19937,N_17470,N_16905);
nand U19938 (N_19938,N_17855,N_16547);
nand U19939 (N_19939,N_16834,N_16842);
and U19940 (N_19940,N_16300,N_17178);
nand U19941 (N_19941,N_16298,N_16589);
and U19942 (N_19942,N_17358,N_17177);
nand U19943 (N_19943,N_17890,N_16328);
xnor U19944 (N_19944,N_16369,N_17471);
or U19945 (N_19945,N_17385,N_17255);
and U19946 (N_19946,N_17838,N_17889);
nor U19947 (N_19947,N_16563,N_17123);
nor U19948 (N_19948,N_17685,N_17805);
and U19949 (N_19949,N_16556,N_16608);
nor U19950 (N_19950,N_16556,N_16973);
nor U19951 (N_19951,N_16883,N_17721);
nand U19952 (N_19952,N_17645,N_17966);
nand U19953 (N_19953,N_16277,N_16272);
or U19954 (N_19954,N_16312,N_16521);
xor U19955 (N_19955,N_17837,N_17224);
or U19956 (N_19956,N_16244,N_17836);
nand U19957 (N_19957,N_16433,N_16037);
nor U19958 (N_19958,N_16159,N_16710);
and U19959 (N_19959,N_17994,N_16328);
or U19960 (N_19960,N_16838,N_16173);
or U19961 (N_19961,N_17884,N_17178);
and U19962 (N_19962,N_16820,N_16456);
or U19963 (N_19963,N_17968,N_17764);
nand U19964 (N_19964,N_17717,N_17329);
or U19965 (N_19965,N_16258,N_17781);
xor U19966 (N_19966,N_17811,N_17207);
and U19967 (N_19967,N_17561,N_16463);
and U19968 (N_19968,N_17108,N_17825);
nand U19969 (N_19969,N_17745,N_17794);
xnor U19970 (N_19970,N_16427,N_16057);
nand U19971 (N_19971,N_16465,N_16981);
or U19972 (N_19972,N_16953,N_16811);
xnor U19973 (N_19973,N_16712,N_17881);
nand U19974 (N_19974,N_16943,N_17365);
or U19975 (N_19975,N_17787,N_17589);
nand U19976 (N_19976,N_16684,N_17419);
nor U19977 (N_19977,N_16818,N_16272);
or U19978 (N_19978,N_16380,N_16560);
or U19979 (N_19979,N_17889,N_17081);
and U19980 (N_19980,N_16943,N_16148);
xor U19981 (N_19981,N_16792,N_17397);
nor U19982 (N_19982,N_17806,N_16494);
nand U19983 (N_19983,N_17443,N_16399);
and U19984 (N_19984,N_16676,N_16439);
xor U19985 (N_19985,N_17729,N_16474);
xor U19986 (N_19986,N_16390,N_16192);
or U19987 (N_19987,N_17086,N_16075);
and U19988 (N_19988,N_17049,N_16833);
and U19989 (N_19989,N_17207,N_16180);
nand U19990 (N_19990,N_16361,N_16074);
xor U19991 (N_19991,N_16716,N_17836);
or U19992 (N_19992,N_17200,N_17976);
nor U19993 (N_19993,N_16929,N_16664);
nand U19994 (N_19994,N_17492,N_16097);
and U19995 (N_19995,N_16174,N_16636);
nor U19996 (N_19996,N_17620,N_17518);
xor U19997 (N_19997,N_16818,N_17661);
and U19998 (N_19998,N_17168,N_17435);
or U19999 (N_19999,N_17134,N_17397);
nand U20000 (N_20000,N_18181,N_18276);
and U20001 (N_20001,N_18344,N_19818);
xor U20002 (N_20002,N_18949,N_18453);
or U20003 (N_20003,N_18214,N_18783);
or U20004 (N_20004,N_18103,N_18871);
nand U20005 (N_20005,N_19394,N_18139);
and U20006 (N_20006,N_19119,N_19343);
nor U20007 (N_20007,N_18784,N_19959);
and U20008 (N_20008,N_19782,N_18705);
and U20009 (N_20009,N_19479,N_19191);
or U20010 (N_20010,N_18252,N_19141);
nand U20011 (N_20011,N_19897,N_19703);
xnor U20012 (N_20012,N_19049,N_19433);
nor U20013 (N_20013,N_18492,N_18065);
nand U20014 (N_20014,N_18433,N_18408);
or U20015 (N_20015,N_19991,N_18971);
or U20016 (N_20016,N_19279,N_19184);
nand U20017 (N_20017,N_19659,N_18685);
and U20018 (N_20018,N_19307,N_18747);
nor U20019 (N_20019,N_18017,N_18954);
xnor U20020 (N_20020,N_18004,N_18948);
or U20021 (N_20021,N_18363,N_18273);
and U20022 (N_20022,N_18209,N_19319);
and U20023 (N_20023,N_19549,N_18441);
or U20024 (N_20024,N_19737,N_19910);
or U20025 (N_20025,N_19366,N_19166);
xor U20026 (N_20026,N_18397,N_19682);
nand U20027 (N_20027,N_19605,N_18880);
or U20028 (N_20028,N_18764,N_19930);
or U20029 (N_20029,N_19144,N_19137);
xor U20030 (N_20030,N_18179,N_18084);
nand U20031 (N_20031,N_19265,N_19778);
and U20032 (N_20032,N_19106,N_19270);
xnor U20033 (N_20033,N_19811,N_18835);
nand U20034 (N_20034,N_19837,N_18845);
or U20035 (N_20035,N_19362,N_18798);
xnor U20036 (N_20036,N_19743,N_18289);
and U20037 (N_20037,N_18975,N_18268);
nor U20038 (N_20038,N_18015,N_18074);
xnor U20039 (N_20039,N_18391,N_18269);
nand U20040 (N_20040,N_19722,N_19906);
or U20041 (N_20041,N_19926,N_19392);
nand U20042 (N_20042,N_18559,N_18473);
xor U20043 (N_20043,N_19446,N_18140);
xnor U20044 (N_20044,N_19601,N_18354);
xor U20045 (N_20045,N_19805,N_18929);
nand U20046 (N_20046,N_19048,N_19323);
nor U20047 (N_20047,N_19123,N_19611);
nor U20048 (N_20048,N_19208,N_19125);
nor U20049 (N_20049,N_19476,N_19620);
and U20050 (N_20050,N_19529,N_19354);
nand U20051 (N_20051,N_18699,N_18120);
nor U20052 (N_20052,N_19239,N_18598);
nand U20053 (N_20053,N_18762,N_18827);
nand U20054 (N_20054,N_19760,N_18199);
and U20055 (N_20055,N_19165,N_19967);
xor U20056 (N_20056,N_18687,N_18914);
and U20057 (N_20057,N_18321,N_19316);
nor U20058 (N_20058,N_18424,N_19506);
nor U20059 (N_20059,N_19448,N_18236);
nand U20060 (N_20060,N_19757,N_18907);
nor U20061 (N_20061,N_19415,N_19627);
nand U20062 (N_20062,N_18070,N_18516);
or U20063 (N_20063,N_18230,N_19105);
xor U20064 (N_20064,N_19101,N_19092);
nor U20065 (N_20065,N_18356,N_19041);
nor U20066 (N_20066,N_19477,N_19538);
nor U20067 (N_20067,N_18045,N_18901);
nor U20068 (N_20068,N_18471,N_18044);
nor U20069 (N_20069,N_19421,N_19725);
xor U20070 (N_20070,N_18723,N_18384);
nor U20071 (N_20071,N_18201,N_18920);
nor U20072 (N_20072,N_19864,N_18107);
or U20073 (N_20073,N_19245,N_19413);
and U20074 (N_20074,N_18266,N_19016);
xor U20075 (N_20075,N_19320,N_19197);
and U20076 (N_20076,N_19887,N_19423);
or U20077 (N_20077,N_19940,N_19247);
and U20078 (N_20078,N_19790,N_18922);
and U20079 (N_20079,N_19430,N_18930);
nor U20080 (N_20080,N_19034,N_18876);
xor U20081 (N_20081,N_19707,N_19751);
nand U20082 (N_20082,N_18742,N_18618);
and U20083 (N_20083,N_18437,N_19764);
nand U20084 (N_20084,N_19796,N_18115);
nor U20085 (N_20085,N_19591,N_18781);
or U20086 (N_20086,N_18864,N_18246);
or U20087 (N_20087,N_19965,N_19717);
and U20088 (N_20088,N_19237,N_19327);
nand U20089 (N_20089,N_18719,N_19289);
or U20090 (N_20090,N_18089,N_18648);
and U20091 (N_20091,N_18466,N_19345);
and U20092 (N_20092,N_19336,N_19787);
xor U20093 (N_20093,N_18805,N_19128);
and U20094 (N_20094,N_19422,N_18357);
nor U20095 (N_20095,N_19256,N_19290);
and U20096 (N_20096,N_19585,N_19693);
xnor U20097 (N_20097,N_19885,N_18106);
xnor U20098 (N_20098,N_19076,N_18241);
nor U20099 (N_20099,N_18317,N_18899);
and U20100 (N_20100,N_18995,N_18878);
and U20101 (N_20101,N_19522,N_19524);
and U20102 (N_20102,N_19969,N_18096);
nand U20103 (N_20103,N_19443,N_19589);
nand U20104 (N_20104,N_18814,N_18231);
nand U20105 (N_20105,N_18955,N_19839);
nor U20106 (N_20106,N_18405,N_18690);
nor U20107 (N_20107,N_19026,N_18756);
and U20108 (N_20108,N_19395,N_19326);
or U20109 (N_20109,N_19139,N_18389);
nor U20110 (N_20110,N_18879,N_18564);
nand U20111 (N_20111,N_18005,N_19153);
nand U20112 (N_20112,N_18320,N_18615);
or U20113 (N_20113,N_18688,N_18720);
nor U20114 (N_20114,N_19892,N_18788);
xor U20115 (N_20115,N_19633,N_18030);
xor U20116 (N_20116,N_18658,N_18640);
nor U20117 (N_20117,N_19329,N_18581);
nand U20118 (N_20118,N_19713,N_19062);
xor U20119 (N_20119,N_19770,N_18154);
nand U20120 (N_20120,N_19911,N_19008);
nand U20121 (N_20121,N_18331,N_19573);
or U20122 (N_20122,N_18675,N_18050);
nand U20123 (N_20123,N_19745,N_19739);
nand U20124 (N_20124,N_19110,N_18663);
nand U20125 (N_20125,N_18137,N_19877);
or U20126 (N_20126,N_19907,N_19124);
nor U20127 (N_20127,N_19070,N_19848);
or U20128 (N_20128,N_18020,N_18039);
nand U20129 (N_20129,N_19259,N_18122);
nor U20130 (N_20130,N_19003,N_19575);
xnor U20131 (N_20131,N_19656,N_19578);
or U20132 (N_20132,N_19935,N_19814);
and U20133 (N_20133,N_19939,N_18082);
nor U20134 (N_20134,N_19450,N_18457);
or U20135 (N_20135,N_19428,N_19813);
or U20136 (N_20136,N_19618,N_18462);
nand U20137 (N_20137,N_18821,N_19871);
xnor U20138 (N_20138,N_18852,N_18296);
and U20139 (N_20139,N_19867,N_18961);
and U20140 (N_20140,N_18114,N_18570);
xor U20141 (N_20141,N_18001,N_19138);
nand U20142 (N_20142,N_18434,N_19229);
or U20143 (N_20143,N_18672,N_19673);
or U20144 (N_20144,N_18253,N_19634);
xnor U20145 (N_20145,N_19521,N_19983);
nor U20146 (N_20146,N_18942,N_19810);
nor U20147 (N_20147,N_18813,N_19360);
xnor U20148 (N_20148,N_18249,N_19334);
and U20149 (N_20149,N_19590,N_18659);
or U20150 (N_20150,N_18505,N_19338);
or U20151 (N_20151,N_19396,N_19361);
nand U20152 (N_20152,N_18562,N_18048);
nor U20153 (N_20153,N_19744,N_18300);
nand U20154 (N_20154,N_19681,N_18409);
nor U20155 (N_20155,N_18332,N_19143);
or U20156 (N_20156,N_19410,N_18586);
xor U20157 (N_20157,N_19039,N_18576);
xor U20158 (N_20158,N_18873,N_19022);
or U20159 (N_20159,N_18449,N_19071);
or U20160 (N_20160,N_19439,N_19834);
and U20161 (N_20161,N_19363,N_19257);
or U20162 (N_20162,N_19655,N_18069);
or U20163 (N_20163,N_19777,N_18972);
xor U20164 (N_20164,N_18067,N_19017);
nor U20165 (N_20165,N_18085,N_19884);
or U20166 (N_20166,N_19631,N_18578);
and U20167 (N_20167,N_18442,N_18816);
or U20168 (N_20168,N_18713,N_18446);
nand U20169 (N_20169,N_18410,N_18667);
xnor U20170 (N_20170,N_18224,N_18313);
nand U20171 (N_20171,N_19828,N_19407);
xnor U20172 (N_20172,N_18771,N_18116);
nand U20173 (N_20173,N_18868,N_18587);
xnor U20174 (N_20174,N_18923,N_18965);
nand U20175 (N_20175,N_19238,N_18744);
and U20176 (N_20176,N_19977,N_19669);
xnor U20177 (N_20177,N_18303,N_18202);
and U20178 (N_20178,N_18606,N_18888);
nor U20179 (N_20179,N_18588,N_19023);
xnor U20180 (N_20180,N_18078,N_18959);
xnor U20181 (N_20181,N_19175,N_19670);
nor U20182 (N_20182,N_18143,N_19132);
and U20183 (N_20183,N_19024,N_19331);
nand U20184 (N_20184,N_18401,N_19306);
nor U20185 (N_20185,N_19462,N_18609);
and U20186 (N_20186,N_19369,N_18537);
nor U20187 (N_20187,N_18019,N_18655);
nor U20188 (N_20188,N_18622,N_19136);
xor U20189 (N_20189,N_18943,N_18770);
xnor U20190 (N_20190,N_19018,N_19944);
xnor U20191 (N_20191,N_19762,N_18536);
and U20192 (N_20192,N_18498,N_19261);
nor U20193 (N_20193,N_18306,N_18823);
nor U20194 (N_20194,N_18799,N_18820);
or U20195 (N_20195,N_18350,N_19516);
or U20196 (N_20196,N_19518,N_19164);
xor U20197 (N_20197,N_19950,N_19704);
nand U20198 (N_20198,N_18228,N_18619);
xnor U20199 (N_20199,N_19458,N_18169);
nand U20200 (N_20200,N_19021,N_18708);
nor U20201 (N_20201,N_18785,N_19142);
nand U20202 (N_20202,N_18242,N_18299);
or U20203 (N_20203,N_18937,N_18524);
xnor U20204 (N_20204,N_18240,N_18502);
or U20205 (N_20205,N_19901,N_19242);
and U20206 (N_20206,N_18522,N_18247);
and U20207 (N_20207,N_19929,N_18915);
nor U20208 (N_20208,N_19927,N_18220);
xnor U20209 (N_20209,N_18765,N_18365);
nand U20210 (N_20210,N_19636,N_19758);
and U20211 (N_20211,N_18308,N_19335);
nor U20212 (N_20212,N_18414,N_19474);
nor U20213 (N_20213,N_18337,N_18964);
nor U20214 (N_20214,N_19356,N_18867);
nand U20215 (N_20215,N_19157,N_18599);
xnor U20216 (N_20216,N_18985,N_18432);
and U20217 (N_20217,N_18523,N_19598);
nor U20218 (N_20218,N_19614,N_18271);
or U20219 (N_20219,N_19667,N_19577);
and U20220 (N_20220,N_19974,N_18893);
nor U20221 (N_20221,N_18396,N_19403);
and U20222 (N_20222,N_19613,N_19696);
xor U20223 (N_20223,N_19683,N_18007);
nor U20224 (N_20224,N_19154,N_18189);
and U20225 (N_20225,N_18525,N_18259);
or U20226 (N_20226,N_19699,N_18894);
nor U20227 (N_20227,N_18786,N_19461);
and U20228 (N_20228,N_18324,N_18666);
xor U20229 (N_20229,N_18552,N_18861);
nand U20230 (N_20230,N_18539,N_19639);
nand U20231 (N_20231,N_19485,N_18286);
or U20232 (N_20232,N_19612,N_18472);
nand U20233 (N_20233,N_18135,N_19738);
nand U20234 (N_20234,N_18183,N_19583);
nand U20235 (N_20235,N_19582,N_18425);
nor U20236 (N_20236,N_19908,N_19066);
xnor U20237 (N_20237,N_19653,N_19187);
nand U20238 (N_20238,N_18913,N_19408);
xor U20239 (N_20239,N_18800,N_18073);
nand U20240 (N_20240,N_18438,N_19315);
and U20241 (N_20241,N_19000,N_18841);
or U20242 (N_20242,N_18594,N_18497);
xor U20243 (N_20243,N_18338,N_19419);
or U20244 (N_20244,N_19204,N_18532);
and U20245 (N_20245,N_18314,N_19209);
nor U20246 (N_20246,N_18194,N_18822);
nand U20247 (N_20247,N_18156,N_19542);
xnor U20248 (N_20248,N_18651,N_18883);
nand U20249 (N_20249,N_18585,N_19176);
nor U20250 (N_20250,N_19380,N_18787);
or U20251 (N_20251,N_19833,N_19030);
and U20252 (N_20252,N_19749,N_18026);
nand U20253 (N_20253,N_18239,N_18460);
nor U20254 (N_20254,N_19444,N_19754);
nand U20255 (N_20255,N_18254,N_18219);
and U20256 (N_20256,N_18161,N_19720);
nor U20257 (N_20257,N_19127,N_18766);
or U20258 (N_20258,N_19414,N_19074);
or U20259 (N_20259,N_18468,N_18611);
and U20260 (N_20260,N_18171,N_18571);
nor U20261 (N_20261,N_18364,N_19708);
nor U20262 (N_20262,N_18167,N_18099);
nand U20263 (N_20263,N_18909,N_18533);
and U20264 (N_20264,N_19296,N_18164);
and U20265 (N_20265,N_19604,N_18682);
or U20266 (N_20266,N_18309,N_19317);
xnor U20267 (N_20267,N_18953,N_19843);
xor U20268 (N_20268,N_19140,N_19009);
or U20269 (N_20269,N_19437,N_19891);
nor U20270 (N_20270,N_19946,N_18866);
xor U20271 (N_20271,N_18634,N_18646);
and U20272 (N_20272,N_19719,N_18939);
nor U20273 (N_20273,N_18126,N_18162);
or U20274 (N_20274,N_19999,N_18006);
nor U20275 (N_20275,N_19268,N_18003);
nand U20276 (N_20276,N_18779,N_19469);
or U20277 (N_20277,N_18060,N_19688);
nor U20278 (N_20278,N_18451,N_18582);
nand U20279 (N_20279,N_18417,N_18612);
nor U20280 (N_20280,N_18144,N_19304);
and U20281 (N_20281,N_18027,N_18825);
or U20282 (N_20282,N_19292,N_18395);
or U20283 (N_20283,N_19120,N_19227);
and U20284 (N_20284,N_19498,N_18383);
and U20285 (N_20285,N_18080,N_19919);
nand U20286 (N_20286,N_19200,N_18245);
nor U20287 (N_20287,N_19493,N_19133);
or U20288 (N_20288,N_19701,N_18349);
nor U20289 (N_20289,N_18166,N_19145);
nand U20290 (N_20290,N_19957,N_19453);
nand U20291 (N_20291,N_19425,N_19882);
nor U20292 (N_20292,N_18511,N_18243);
xnor U20293 (N_20293,N_18662,N_19569);
nand U20294 (N_20294,N_18294,N_18643);
nor U20295 (N_20295,N_19888,N_19266);
nor U20296 (N_20296,N_19951,N_18898);
nand U20297 (N_20297,N_19500,N_19883);
or U20298 (N_20298,N_18858,N_19530);
nand U20299 (N_20299,N_18420,N_19515);
nand U20300 (N_20300,N_19122,N_18288);
and U20301 (N_20301,N_19340,N_19815);
xor U20302 (N_20302,N_19355,N_18633);
nand U20303 (N_20303,N_18413,N_19378);
and U20304 (N_20304,N_18741,N_18547);
nor U20305 (N_20305,N_19973,N_18627);
nor U20306 (N_20306,N_18887,N_18530);
nor U20307 (N_20307,N_19564,N_19217);
and U20308 (N_20308,N_19172,N_19889);
or U20309 (N_20309,N_19960,N_18217);
xor U20310 (N_20310,N_19218,N_19994);
xor U20311 (N_20311,N_18870,N_19607);
xnor U20312 (N_20312,N_18057,N_18427);
and U20313 (N_20313,N_19922,N_18444);
and U20314 (N_20314,N_19287,N_19121);
nand U20315 (N_20315,N_19010,N_19517);
nor U20316 (N_20316,N_18695,N_18091);
or U20317 (N_20317,N_19002,N_18047);
and U20318 (N_20318,N_18376,N_18318);
xor U20319 (N_20319,N_19630,N_18951);
nor U20320 (N_20320,N_19251,N_18275);
or U20321 (N_20321,N_18347,N_19112);
or U20322 (N_20322,N_18066,N_19832);
nor U20323 (N_20323,N_19635,N_18649);
nand U20324 (N_20324,N_18155,N_18422);
xnor U20325 (N_20325,N_18684,N_18173);
and U20326 (N_20326,N_19663,N_18234);
or U20327 (N_20327,N_18558,N_18042);
nand U20328 (N_20328,N_18706,N_18223);
nor U20329 (N_20329,N_18508,N_19748);
nand U20330 (N_20330,N_19183,N_18653);
or U20331 (N_20331,N_19324,N_18808);
nand U20332 (N_20332,N_18660,N_18863);
nand U20333 (N_20333,N_18669,N_19253);
and U20334 (N_20334,N_19563,N_19997);
and U20335 (N_20335,N_18411,N_19987);
xor U20336 (N_20336,N_18076,N_19936);
xnor U20337 (N_20337,N_18573,N_18373);
xnor U20338 (N_20338,N_18415,N_19706);
and U20339 (N_20339,N_18426,N_19916);
nand U20340 (N_20340,N_19075,N_19241);
and U20341 (N_20341,N_18304,N_18416);
nor U20342 (N_20342,N_18812,N_19761);
and U20343 (N_20343,N_18121,N_19866);
nor U20344 (N_20344,N_18734,N_19056);
nand U20345 (N_20345,N_19733,N_18575);
or U20346 (N_20346,N_19118,N_18727);
xnor U20347 (N_20347,N_19225,N_18108);
and U20348 (N_20348,N_18485,N_19181);
or U20349 (N_20349,N_18418,N_19841);
nor U20350 (N_20350,N_18488,N_19258);
or U20351 (N_20351,N_19823,N_19321);
nand U20352 (N_20352,N_19189,N_19234);
and U20353 (N_20353,N_18302,N_19005);
or U20354 (N_20354,N_18345,N_19586);
nand U20355 (N_20355,N_19020,N_19060);
or U20356 (N_20356,N_19351,N_18833);
nand U20357 (N_20357,N_19617,N_18804);
nor U20358 (N_20358,N_19525,N_19505);
xnor U20359 (N_20359,N_19385,N_18777);
xnor U20360 (N_20360,N_18512,N_19250);
xor U20361 (N_20361,N_19742,N_18210);
xor U20362 (N_20362,N_19186,N_19384);
nand U20363 (N_20363,N_19107,N_19382);
xor U20364 (N_20364,N_18518,N_19735);
and U20365 (N_20365,N_18514,N_19192);
xor U20366 (N_20366,N_19089,N_19771);
xnor U20367 (N_20367,N_18890,N_19019);
or U20368 (N_20368,N_18305,N_19857);
and U20369 (N_20369,N_19429,N_18200);
xnor U20370 (N_20370,N_18791,N_18875);
nand U20371 (N_20371,N_18281,N_18423);
nand U20372 (N_20372,N_19054,N_19223);
xnor U20373 (N_20373,N_19551,N_19700);
nand U20374 (N_20374,N_18185,N_18105);
xnor U20375 (N_20375,N_18645,N_19836);
and U20376 (N_20376,N_18597,N_18479);
or U20377 (N_20377,N_19114,N_18267);
nor U20378 (N_20378,N_18257,N_19497);
or U20379 (N_20379,N_19540,N_18014);
nor U20380 (N_20380,N_19817,N_19104);
nor U20381 (N_20381,N_18732,N_18342);
or U20382 (N_20382,N_18436,N_19531);
and U20383 (N_20383,N_19822,N_18538);
or U20384 (N_20384,N_19342,N_18726);
xnor U20385 (N_20385,N_19792,N_18233);
or U20386 (N_20386,N_18693,N_19464);
and U20387 (N_20387,N_18819,N_19081);
and U20388 (N_20388,N_18385,N_18795);
nand U20389 (N_20389,N_19799,N_18832);
nand U20390 (N_20390,N_19216,N_18421);
nor U20391 (N_20391,N_19073,N_19890);
nor U20392 (N_20392,N_18464,N_18158);
and U20393 (N_20393,N_18095,N_18644);
nor U20394 (N_20394,N_18381,N_19894);
nand U20395 (N_20395,N_18931,N_18407);
nand U20396 (N_20396,N_18509,N_19028);
and U20397 (N_20397,N_19674,N_19202);
or U20398 (N_20398,N_19678,N_19077);
xor U20399 (N_20399,N_19093,N_19246);
or U20400 (N_20400,N_19135,N_18661);
xor U20401 (N_20401,N_19219,N_18149);
or U20402 (N_20402,N_19685,N_19278);
nand U20403 (N_20403,N_19948,N_18962);
and U20404 (N_20404,N_19849,N_18119);
nand U20405 (N_20405,N_19687,N_18987);
nand U20406 (N_20406,N_18463,N_19621);
or U20407 (N_20407,N_19511,N_19170);
xor U20408 (N_20408,N_19178,N_19155);
nand U20409 (N_20409,N_18041,N_18531);
and U20410 (N_20410,N_19083,N_18307);
xor U20411 (N_20411,N_18796,N_18043);
xor U20412 (N_20412,N_18974,N_19100);
xor U20413 (N_20413,N_18809,N_18452);
xnor U20414 (N_20414,N_19824,N_18704);
and U20415 (N_20415,N_19859,N_19405);
nand U20416 (N_20416,N_19881,N_18340);
xnor U20417 (N_20417,N_18256,N_18709);
xor U20418 (N_20418,N_19486,N_19193);
and U20419 (N_20419,N_18624,N_18343);
nand U20420 (N_20420,N_19001,N_18163);
and U20421 (N_20421,N_18996,N_19691);
and U20422 (N_20422,N_19766,N_19947);
xor U20423 (N_20423,N_19094,N_19252);
or U20424 (N_20424,N_18792,N_19496);
xnor U20425 (N_20425,N_18717,N_18842);
or U20426 (N_20426,N_19554,N_19150);
and U20427 (N_20427,N_19404,N_19492);
nand U20428 (N_20428,N_18759,N_19567);
xnor U20429 (N_20429,N_19190,N_18950);
or U20430 (N_20430,N_18725,N_19214);
nor U20431 (N_20431,N_19007,N_18550);
nand U20432 (N_20432,N_18270,N_18297);
nor U20433 (N_20433,N_19014,N_18903);
or U20434 (N_20434,N_18580,N_19169);
and U20435 (N_20435,N_18021,N_19199);
nand U20436 (N_20436,N_18977,N_18094);
or U20437 (N_20437,N_18638,N_18853);
xor U20438 (N_20438,N_18574,N_19924);
nor U20439 (N_20439,N_18419,N_19043);
and U20440 (N_20440,N_19116,N_18993);
and U20441 (N_20441,N_19765,N_19029);
and U20442 (N_20442,N_18767,N_19643);
xor U20443 (N_20443,N_19364,N_19286);
xnor U20444 (N_20444,N_18123,N_19949);
nor U20445 (N_20445,N_18834,N_19330);
nand U20446 (N_20446,N_18483,N_19807);
and U20447 (N_20447,N_19724,N_18815);
or U20448 (N_20448,N_18075,N_18063);
nand U20449 (N_20449,N_18211,N_19844);
and U20450 (N_20450,N_19510,N_18641);
or U20451 (N_20451,N_18008,N_19979);
nor U20452 (N_20452,N_18431,N_19872);
or U20453 (N_20453,N_18399,N_19236);
nor U20454 (N_20454,N_18495,N_18282);
or U20455 (N_20455,N_19282,N_18592);
xor U20456 (N_20456,N_19456,N_18885);
nand U20457 (N_20457,N_18430,N_19090);
xor U20458 (N_20458,N_19357,N_18983);
xnor U20459 (N_20459,N_18774,N_18404);
or U20460 (N_20460,N_18896,N_19543);
or U20461 (N_20461,N_19096,N_18712);
or U20462 (N_20462,N_18250,N_18098);
or U20463 (N_20463,N_19665,N_18847);
xor U20464 (N_20464,N_18900,N_18077);
xor U20465 (N_20465,N_18049,N_18142);
nor U20466 (N_20466,N_19318,N_18928);
nor U20467 (N_20467,N_19953,N_18711);
and U20468 (N_20468,N_19809,N_18761);
nand U20469 (N_20469,N_19523,N_18617);
nand U20470 (N_20470,N_18680,N_18738);
and U20471 (N_20471,N_19767,N_19716);
nand U20472 (N_20472,N_18130,N_18190);
nand U20473 (N_20473,N_19163,N_18100);
and U20474 (N_20474,N_19185,N_18177);
or U20475 (N_20475,N_19705,N_18292);
or U20476 (N_20476,N_18892,N_19103);
xnor U20477 (N_20477,N_18590,N_18941);
xor U20478 (N_20478,N_19873,N_18938);
or U20479 (N_20479,N_19281,N_18172);
nand U20480 (N_20480,N_19562,N_18068);
nand U20481 (N_20481,N_18461,N_19381);
xnor U20482 (N_20482,N_19855,N_18776);
nor U20483 (N_20483,N_18970,N_18475);
and U20484 (N_20484,N_19267,N_18593);
or U20485 (N_20485,N_18957,N_18639);
nand U20486 (N_20486,N_19438,N_18544);
nor U20487 (N_20487,N_19417,N_19393);
xor U20488 (N_20488,N_19455,N_18117);
nor U20489 (N_20489,N_19058,N_18353);
nor U20490 (N_20490,N_18601,N_19442);
nand U20491 (N_20491,N_18636,N_18513);
or U20492 (N_20492,N_18002,N_18600);
nand U20493 (N_20493,N_19791,N_19055);
or U20494 (N_20494,N_19078,N_19389);
and U20495 (N_20495,N_19398,N_19721);
nor U20496 (N_20496,N_19695,N_19248);
and U20497 (N_20497,N_19769,N_19314);
xnor U20498 (N_20498,N_18118,N_18101);
nor U20499 (N_20499,N_19156,N_18377);
xor U20500 (N_20500,N_19006,N_19552);
and U20501 (N_20501,N_19339,N_18104);
nor U20502 (N_20502,N_18386,N_19915);
nor U20503 (N_20503,N_19220,N_19905);
and U20504 (N_20504,N_19491,N_18577);
nor U20505 (N_20505,N_19276,N_19179);
nand U20506 (N_20506,N_19283,N_19938);
or U20507 (N_20507,N_18032,N_18872);
or U20508 (N_20508,N_19499,N_18195);
xnor U20509 (N_20509,N_19602,N_18133);
nor U20510 (N_20510,N_19232,N_19876);
and U20511 (N_20511,N_18840,N_19303);
or U20512 (N_20512,N_18009,N_18197);
and U20513 (N_20513,N_19033,N_18794);
or U20514 (N_20514,N_19657,N_19037);
xnor U20515 (N_20515,N_19599,N_19875);
nand U20516 (N_20516,N_19298,N_19986);
and U20517 (N_20517,N_19870,N_18310);
nor U20518 (N_20518,N_19117,N_19955);
nand U20519 (N_20519,N_18691,N_19988);
or U20520 (N_20520,N_19862,N_19806);
or U20521 (N_20521,N_19013,N_18689);
nand U20522 (N_20522,N_19235,N_18566);
xor U20523 (N_20523,N_19920,N_19160);
or U20524 (N_20524,N_19053,N_19652);
xor U20525 (N_20525,N_18626,N_18569);
or U20526 (N_20526,N_19819,N_18454);
and U20527 (N_20527,N_19012,N_19694);
and U20528 (N_20528,N_19383,N_19418);
nor U20529 (N_20529,N_18010,N_19064);
nor U20530 (N_20530,N_18710,N_19654);
or U20531 (N_20531,N_18191,N_19971);
xnor U20532 (N_20532,N_18750,N_19904);
or U20533 (N_20533,N_19463,N_18311);
or U20534 (N_20534,N_18735,N_19374);
nand U20535 (N_20535,N_18677,N_19457);
xor U20536 (N_20536,N_18981,N_18013);
or U20537 (N_20537,N_19271,N_19619);
and U20538 (N_20538,N_18359,N_18697);
or U20539 (N_20539,N_18838,N_18718);
and U20540 (N_20540,N_18824,N_18527);
nand U20541 (N_20541,N_18647,N_18628);
or U20542 (N_20542,N_19785,N_18037);
nand U20543 (N_20543,N_19294,N_18775);
and U20544 (N_20544,N_18222,N_18174);
nor U20545 (N_20545,N_19108,N_19545);
nand U20546 (N_20546,N_18956,N_18428);
xnor U20547 (N_20547,N_18402,N_19854);
or U20548 (N_20548,N_18132,N_18613);
and U20549 (N_20549,N_19194,N_19489);
or U20550 (N_20550,N_19390,N_19780);
xnor U20551 (N_20551,N_19626,N_18459);
and U20552 (N_20552,N_19560,N_19397);
and U20553 (N_20553,N_19734,N_19391);
xor U20554 (N_20554,N_19865,N_18072);
and U20555 (N_20555,N_18328,N_19526);
or U20556 (N_20556,N_18440,N_18702);
xnor U20557 (N_20557,N_18301,N_19963);
or U20558 (N_20558,N_18455,N_18874);
or U20559 (N_20559,N_19921,N_18496);
and U20560 (N_20560,N_19454,N_19660);
or U20561 (N_20561,N_19297,N_19786);
nand U20562 (N_20562,N_18035,N_18607);
nor U20563 (N_20563,N_18011,N_18721);
and U20564 (N_20564,N_19804,N_19547);
or U20565 (N_20565,N_19750,N_19050);
xnor U20566 (N_20566,N_18567,N_18470);
nor U20567 (N_20567,N_18031,N_18782);
or U20568 (N_20568,N_18940,N_18754);
or U20569 (N_20569,N_18274,N_18160);
nor U20570 (N_20570,N_19481,N_18052);
nand U20571 (N_20571,N_18925,N_18212);
xor U20572 (N_20572,N_19344,N_18982);
and U20573 (N_20573,N_18351,N_18227);
and U20574 (N_20574,N_19623,N_19795);
or U20575 (N_20575,N_19295,N_19918);
xnor U20576 (N_20576,N_19507,N_18012);
xnor U20577 (N_20577,N_19856,N_18087);
nor U20578 (N_20578,N_19273,N_19113);
nand U20579 (N_20579,N_18146,N_19495);
or U20580 (N_20580,N_19874,N_18589);
or U20581 (N_20581,N_19640,N_19553);
xor U20582 (N_20582,N_18447,N_18186);
or U20583 (N_20583,N_18188,N_18650);
or U20584 (N_20584,N_19992,N_18261);
nor U20585 (N_20585,N_18621,N_19942);
nand U20586 (N_20586,N_18665,N_18596);
and U20587 (N_20587,N_18542,N_18676);
or U20588 (N_20588,N_19188,N_18400);
nand U20589 (N_20589,N_18504,N_18990);
xnor U20590 (N_20590,N_19431,N_19566);
or U20591 (N_20591,N_19679,N_18207);
and U20592 (N_20592,N_18284,N_19411);
or U20593 (N_20593,N_18232,N_19661);
nor U20594 (N_20594,N_18758,N_18855);
nand U20595 (N_20595,N_19680,N_19820);
or U20596 (N_20596,N_19755,N_18369);
and U20597 (N_20597,N_18683,N_19311);
nand U20598 (N_20598,N_18595,N_18062);
nand U20599 (N_20599,N_19972,N_19976);
nand U20600 (N_20600,N_19789,N_18806);
or U20601 (N_20601,N_19923,N_18968);
nand U20602 (N_20602,N_19313,N_19206);
or U20603 (N_20603,N_18773,N_19468);
and U20604 (N_20604,N_18360,N_19490);
or U20605 (N_20605,N_19173,N_18204);
and U20606 (N_20606,N_19561,N_18326);
nand U20607 (N_20607,N_19645,N_18797);
and U20608 (N_20608,N_19580,N_19349);
nor U20609 (N_20609,N_19471,N_18448);
and U20610 (N_20610,N_18869,N_18258);
nand U20611 (N_20611,N_18579,N_19460);
xnor U20612 (N_20612,N_19753,N_18817);
nand U20613 (N_20613,N_19426,N_19328);
or U20614 (N_20614,N_18467,N_19291);
and U20615 (N_20615,N_18752,N_19851);
xor U20616 (N_20616,N_19584,N_18387);
nand U20617 (N_20617,N_18745,N_19594);
and U20618 (N_20618,N_19098,N_19201);
nor U20619 (N_20619,N_18477,N_19858);
nand U20620 (N_20620,N_19260,N_18443);
nand U20621 (N_20621,N_18673,N_18213);
xor U20622 (N_20622,N_19945,N_18912);
nand U20623 (N_20623,N_18406,N_18291);
xnor U20624 (N_20624,N_19781,N_18642);
nor U20625 (N_20625,N_19729,N_18681);
and U20626 (N_20626,N_18584,N_19367);
nor U20627 (N_20627,N_18656,N_18203);
xor U20628 (N_20628,N_19962,N_18674);
and U20629 (N_20629,N_19537,N_19459);
xnor U20630 (N_20630,N_19980,N_18670);
and U20631 (N_20631,N_18637,N_19608);
or U20632 (N_20632,N_18147,N_18362);
and U20633 (N_20633,N_18802,N_19210);
xor U20634 (N_20634,N_18946,N_19830);
and U20635 (N_20635,N_19084,N_18958);
and U20636 (N_20636,N_18724,N_18679);
or U20637 (N_20637,N_18986,N_18857);
and U20638 (N_20638,N_18079,N_18548);
and U20639 (N_20639,N_18358,N_19662);
and U20640 (N_20640,N_18760,N_19368);
or U20641 (N_20641,N_18022,N_18378);
and U20642 (N_20642,N_18908,N_18093);
or U20643 (N_20643,N_18563,N_19099);
or U20644 (N_20644,N_19111,N_18215);
or U20645 (N_20645,N_19535,N_19115);
nor U20646 (N_20646,N_18412,N_19896);
nor U20647 (N_20647,N_19177,N_18846);
and U20648 (N_20648,N_19167,N_19982);
nor U20649 (N_20649,N_18629,N_19467);
or U20650 (N_20650,N_18054,N_19726);
or U20651 (N_20651,N_19269,N_18469);
or U20652 (N_20652,N_19686,N_18476);
xnor U20653 (N_20653,N_19231,N_18265);
nand U20654 (N_20654,N_19195,N_19480);
nand U20655 (N_20655,N_18616,N_19300);
or U20656 (N_20656,N_18346,N_19434);
and U20657 (N_20657,N_18316,N_19379);
xnor U20658 (N_20658,N_19913,N_18790);
nand U20659 (N_20659,N_18945,N_19341);
nand U20660 (N_20660,N_19226,N_18934);
nor U20661 (N_20661,N_19513,N_19718);
nand U20662 (N_20662,N_19148,N_19574);
xnor U20663 (N_20663,N_19171,N_18083);
or U20664 (N_20664,N_18753,N_18728);
nor U20665 (N_20665,N_19072,N_19386);
nand U20666 (N_20666,N_18620,N_18748);
nor U20667 (N_20667,N_19642,N_19998);
xor U20668 (N_20668,N_19277,N_18714);
nor U20669 (N_20669,N_18591,N_19768);
nor U20670 (N_20670,N_19353,N_19420);
and U20671 (N_20671,N_18722,N_18390);
xnor U20672 (N_20672,N_19559,N_19348);
and U20673 (N_20673,N_19063,N_19162);
or U20674 (N_20674,N_19581,N_18947);
or U20675 (N_20675,N_19903,N_19676);
or U20676 (N_20676,N_19447,N_18631);
nor U20677 (N_20677,N_19091,N_19221);
xor U20678 (N_20678,N_19821,N_18394);
nand U20679 (N_20679,N_19322,N_18371);
and U20680 (N_20680,N_18671,N_18484);
nor U20681 (N_20681,N_19233,N_19416);
nand U20682 (N_20682,N_19829,N_19488);
or U20683 (N_20683,N_18549,N_19714);
nand U20684 (N_20684,N_18465,N_18124);
xor U20685 (N_20685,N_19376,N_18884);
and U20686 (N_20686,N_18102,N_19047);
nand U20687 (N_20687,N_19067,N_19377);
or U20688 (N_20688,N_19052,N_19736);
nand U20689 (N_20689,N_19784,N_18327);
and U20690 (N_20690,N_19365,N_18664);
nor U20691 (N_20691,N_18339,N_18976);
and U20692 (N_20692,N_18244,N_18280);
xnor U20693 (N_20693,N_19032,N_18517);
nor U20694 (N_20694,N_19779,N_19989);
nor U20695 (N_20695,N_19995,N_19182);
xor U20696 (N_20696,N_18482,N_18831);
or U20697 (N_20697,N_18507,N_18789);
xnor U20698 (N_20698,N_19035,N_19375);
or U20699 (N_20699,N_19595,N_18998);
xor U20700 (N_20700,N_18319,N_18604);
nand U20701 (N_20701,N_19800,N_18715);
or U20702 (N_20702,N_18323,N_19044);
nor U20703 (N_20703,N_18138,N_19697);
or U20704 (N_20704,N_19042,N_18262);
nand U20705 (N_20705,N_19978,N_19933);
xor U20706 (N_20706,N_18778,N_19061);
or U20707 (N_20707,N_18113,N_19299);
xnor U20708 (N_20708,N_18810,N_19637);
and U20709 (N_20709,N_19671,N_18150);
or U20710 (N_20710,N_18180,N_18733);
xnor U20711 (N_20711,N_18780,N_19352);
xnor U20712 (N_20712,N_19472,N_18370);
and U20713 (N_20713,N_19808,N_18141);
nand U20714 (N_20714,N_18251,N_18828);
nor U20715 (N_20715,N_19644,N_18023);
or U20716 (N_20716,N_19672,N_19051);
and U20717 (N_20717,N_18196,N_19198);
and U20718 (N_20718,N_18630,N_19534);
nand U20719 (N_20719,N_18551,N_18368);
and U20720 (N_20720,N_18086,N_19224);
xor U20721 (N_20721,N_19544,N_19424);
xor U20722 (N_20722,N_19159,N_18487);
or U20723 (N_20723,N_19309,N_19548);
nand U20724 (N_20724,N_19036,N_18895);
xor U20725 (N_20725,N_18330,N_18392);
xor U20726 (N_20726,N_19388,N_18029);
xor U20727 (N_20727,N_18145,N_19880);
and U20728 (N_20728,N_18263,N_19827);
nor U20729 (N_20729,N_18526,N_19558);
or U20730 (N_20730,N_19168,N_19180);
xor U20731 (N_20731,N_19372,N_19196);
xnor U20732 (N_20732,N_18829,N_19943);
or U20733 (N_20733,N_18919,N_19503);
xor U20734 (N_20734,N_18285,N_18290);
or U20735 (N_20735,N_18111,N_18372);
nand U20736 (N_20736,N_18602,N_19350);
nor U20737 (N_20737,N_19895,N_18016);
and U20738 (N_20738,N_18134,N_19088);
or U20739 (N_20739,N_19147,N_19284);
nand U20740 (N_20740,N_19015,N_19993);
or U20741 (N_20741,N_19387,N_18746);
nand U20742 (N_20742,N_19520,N_19031);
and U20743 (N_20743,N_18889,N_19146);
nor U20744 (N_20744,N_19305,N_18904);
nor U20745 (N_20745,N_18737,N_18749);
and U20746 (N_20746,N_19592,N_18152);
xor U20747 (N_20747,N_19941,N_18902);
and U20748 (N_20748,N_18374,N_18226);
and U20749 (N_20749,N_18603,N_18905);
nor U20750 (N_20750,N_18515,N_18112);
and U20751 (N_20751,N_19373,N_18393);
xor U20752 (N_20752,N_18917,N_18848);
nor U20753 (N_20753,N_18877,N_18891);
and U20754 (N_20754,N_19912,N_19514);
and U20755 (N_20755,N_19850,N_19293);
nand U20756 (N_20756,N_18260,N_19346);
nor U20757 (N_20757,N_19648,N_18994);
nor U20758 (N_20758,N_19325,N_18860);
nand U20759 (N_20759,N_18493,N_19732);
or U20760 (N_20760,N_19675,N_19937);
or U20761 (N_20761,N_18071,N_19763);
nor U20762 (N_20762,N_18897,N_19600);
nand U20763 (N_20763,N_18528,N_18333);
xor U20764 (N_20764,N_18125,N_18736);
and U20765 (N_20765,N_18850,N_18109);
nor U20766 (N_20766,N_18836,N_19069);
nand U20767 (N_20767,N_19371,N_18543);
nand U20768 (N_20768,N_18382,N_19205);
and U20769 (N_20769,N_19952,N_18984);
nor U20770 (N_20770,N_19557,N_19715);
or U20771 (N_20771,N_19255,N_19095);
xor U20772 (N_20772,N_19451,N_18916);
nand U20773 (N_20773,N_19087,N_18973);
or U20774 (N_20774,N_19658,N_18610);
nor U20775 (N_20775,N_18491,N_19126);
xnor U20776 (N_20776,N_18605,N_19158);
nand U20777 (N_20777,N_19853,N_19861);
and U20778 (N_20778,N_18131,N_18334);
nor U20779 (N_20779,N_19909,N_19046);
or U20780 (N_20780,N_18398,N_19596);
or U20781 (N_20781,N_19783,N_18729);
xnor U20782 (N_20782,N_19027,N_18148);
nand U20783 (N_20783,N_19961,N_19449);
nor U20784 (N_20784,N_18283,N_19649);
nand U20785 (N_20785,N_19134,N_18963);
xnor U20786 (N_20786,N_19302,N_18168);
nor U20787 (N_20787,N_19692,N_18678);
or U20788 (N_20788,N_19587,N_19222);
and U20789 (N_20789,N_19109,N_18136);
nand U20790 (N_20790,N_18992,N_19203);
nand U20791 (N_20791,N_18967,N_19478);
nor U20792 (N_20792,N_19568,N_19402);
and U20793 (N_20793,N_18264,N_18489);
nand U20794 (N_20794,N_19151,N_19332);
nand U20795 (N_20795,N_19958,N_18859);
and U20796 (N_20796,N_18960,N_19964);
xor U20797 (N_20797,N_18206,N_19536);
nor U20798 (N_20798,N_18743,N_19576);
or U20799 (N_20799,N_18429,N_18830);
xor U20800 (N_20800,N_19501,N_18336);
nand U20801 (N_20801,N_18403,N_18456);
nand U20802 (N_20802,N_19508,N_19632);
nor U20803 (N_20803,N_19565,N_18906);
and U20804 (N_20804,N_18763,N_18352);
xnor U20805 (N_20805,N_19555,N_19690);
xnor U20806 (N_20806,N_18807,N_19914);
nand U20807 (N_20807,N_18935,N_19684);
nor U20808 (N_20808,N_19798,N_19057);
xnor U20809 (N_20809,N_18040,N_18170);
nor U20810 (N_20810,N_18038,N_19931);
or U20811 (N_20811,N_19406,N_19512);
xor U20812 (N_20812,N_18450,N_19504);
nor U20813 (N_20813,N_18478,N_19731);
and U20814 (N_20814,N_19131,N_19572);
nor U20815 (N_20815,N_18110,N_18519);
and U20816 (N_20816,N_19709,N_18028);
xor U20817 (N_20817,N_18686,N_19102);
or U20818 (N_20818,N_19606,N_18999);
and U20819 (N_20819,N_18851,N_19243);
and U20820 (N_20820,N_19466,N_19934);
nand U20821 (N_20821,N_18716,N_19759);
nor U20822 (N_20822,N_19710,N_18237);
nor U20823 (N_20823,N_19615,N_18024);
nor U20824 (N_20824,N_18731,N_19863);
nor U20825 (N_20825,N_19747,N_18295);
xnor U20826 (N_20826,N_19370,N_19174);
or U20827 (N_20827,N_18036,N_18635);
xor U20828 (N_20828,N_19746,N_19597);
or U20829 (N_20829,N_18772,N_18059);
and U20830 (N_20830,N_18856,N_18361);
xor U20831 (N_20831,N_18157,N_19541);
and U20832 (N_20832,N_18033,N_19080);
nor U20833 (N_20833,N_19925,N_19228);
or U20834 (N_20834,N_19794,N_19465);
and U20835 (N_20835,N_19869,N_18312);
xnor U20836 (N_20836,N_18988,N_18886);
nor U20837 (N_20837,N_19550,N_19059);
nand U20838 (N_20838,N_18952,N_19625);
nand U20839 (N_20839,N_18127,N_18924);
nand U20840 (N_20840,N_19264,N_18439);
xor U20841 (N_20841,N_18911,N_19040);
nor U20842 (N_20842,N_19129,N_18844);
nor U20843 (N_20843,N_19668,N_19244);
xor U20844 (N_20844,N_19068,N_19275);
and U20845 (N_20845,N_18555,N_18692);
nor U20846 (N_20846,N_18698,N_19975);
xnor U20847 (N_20847,N_18090,N_19097);
nand U20848 (N_20848,N_19624,N_19740);
nor U20849 (N_20849,N_19985,N_19571);
nor U20850 (N_20850,N_18989,N_19845);
xor U20851 (N_20851,N_19533,N_18769);
xnor U20852 (N_20852,N_18811,N_18921);
xnor U20853 (N_20853,N_19641,N_19698);
nand U20854 (N_20854,N_18272,N_18221);
nor U20855 (N_20855,N_18445,N_19773);
or U20856 (N_20856,N_19482,N_19262);
or U20857 (N_20857,N_19527,N_18793);
or U20858 (N_20858,N_18153,N_19435);
nor U20859 (N_20859,N_19902,N_18235);
nor U20860 (N_20860,N_18218,N_18388);
nand U20861 (N_20861,N_18572,N_18053);
nand U20862 (N_20862,N_19445,N_19149);
or U20863 (N_20863,N_18503,N_18435);
nand U20864 (N_20864,N_18051,N_19556);
and U20865 (N_20865,N_18055,N_19730);
xor U20866 (N_20866,N_19473,N_18700);
or U20867 (N_20867,N_18927,N_18966);
and U20868 (N_20868,N_19215,N_18521);
nor U20869 (N_20869,N_18315,N_18751);
nand U20870 (N_20870,N_19878,N_18865);
nand U20871 (N_20871,N_18707,N_19990);
and U20872 (N_20872,N_18740,N_18703);
nor U20873 (N_20873,N_18545,N_18335);
nand U20874 (N_20874,N_18696,N_19025);
and U20875 (N_20875,N_18128,N_19825);
nor U20876 (N_20876,N_19310,N_19475);
nand U20877 (N_20877,N_18064,N_18129);
or U20878 (N_20878,N_18554,N_18208);
and U20879 (N_20879,N_18474,N_18614);
nand U20880 (N_20880,N_19045,N_18380);
nor U20881 (N_20881,N_19886,N_19285);
or U20882 (N_20882,N_19852,N_19546);
xnor U20883 (N_20883,N_19230,N_18632);
nand U20884 (N_20884,N_19966,N_19711);
nand U20885 (N_20885,N_19358,N_19793);
nand U20886 (N_20886,N_19756,N_18494);
nor U20887 (N_20887,N_19802,N_18481);
and U20888 (N_20888,N_19570,N_18216);
xor U20889 (N_20889,N_19629,N_19752);
xnor U20890 (N_20890,N_18480,N_19288);
xnor U20891 (N_20891,N_18755,N_18991);
xor U20892 (N_20892,N_19409,N_19666);
xnor U20893 (N_20893,N_19399,N_19337);
nand U20894 (N_20894,N_19956,N_19212);
nor U20895 (N_20895,N_18944,N_19954);
nand U20896 (N_20896,N_19484,N_18701);
nand U20897 (N_20897,N_18854,N_18837);
and U20898 (N_20898,N_18056,N_19441);
or U20899 (N_20899,N_19401,N_19440);
xor U20900 (N_20900,N_18768,N_18205);
and U20901 (N_20901,N_19772,N_19400);
nor U20902 (N_20902,N_19011,N_19898);
nand U20903 (N_20903,N_18801,N_18936);
nor U20904 (N_20904,N_19741,N_18348);
nand U20905 (N_20905,N_18255,N_18978);
nand U20906 (N_20906,N_19579,N_19664);
nand U20907 (N_20907,N_18979,N_19085);
or U20908 (N_20908,N_18034,N_18694);
nand U20909 (N_20909,N_19532,N_19152);
or U20910 (N_20910,N_19130,N_18458);
or U20911 (N_20911,N_18862,N_18623);
and U20912 (N_20912,N_19797,N_18910);
nand U20913 (N_20913,N_19213,N_19588);
nor U20914 (N_20914,N_19254,N_19727);
xnor U20915 (N_20915,N_18843,N_19628);
xor U20916 (N_20916,N_19263,N_19427);
xor U20917 (N_20917,N_18159,N_19436);
xor U20918 (N_20918,N_18583,N_18818);
and U20919 (N_20919,N_18325,N_18025);
and U20920 (N_20920,N_19968,N_18165);
nor U20921 (N_20921,N_19470,N_18061);
nor U20922 (N_20922,N_19487,N_18248);
nand U20923 (N_20923,N_19803,N_18541);
nand U20924 (N_20924,N_18486,N_18329);
xor U20925 (N_20925,N_18657,N_19838);
nand U20926 (N_20926,N_19312,N_18561);
and U20927 (N_20927,N_19646,N_18277);
xnor U20928 (N_20928,N_18546,N_19868);
xor U20929 (N_20929,N_19677,N_18187);
nor U20930 (N_20930,N_18826,N_19846);
nor U20931 (N_20931,N_18757,N_18933);
or U20932 (N_20932,N_19812,N_18081);
and U20933 (N_20933,N_19775,N_19432);
or U20934 (N_20934,N_19728,N_18176);
nand U20935 (N_20935,N_18535,N_18500);
and U20936 (N_20936,N_19842,N_19509);
nand U20937 (N_20937,N_19996,N_19847);
or U20938 (N_20938,N_19840,N_18490);
or U20939 (N_20939,N_19928,N_18980);
nand U20940 (N_20940,N_19651,N_18560);
and U20941 (N_20941,N_19240,N_18668);
or U20942 (N_20942,N_18341,N_18184);
and U20943 (N_20943,N_19788,N_19528);
nand U20944 (N_20944,N_19774,N_18225);
or U20945 (N_20945,N_18556,N_18565);
or U20946 (N_20946,N_19650,N_19702);
nand U20947 (N_20947,N_18151,N_19333);
and U20948 (N_20948,N_18608,N_18182);
nand U20949 (N_20949,N_19917,N_19689);
nor U20950 (N_20950,N_19816,N_19274);
nor U20951 (N_20951,N_18175,N_18926);
and U20952 (N_20952,N_18018,N_18278);
xnor U20953 (N_20953,N_19801,N_18193);
nor U20954 (N_20954,N_19622,N_19082);
or U20955 (N_20955,N_19519,N_18520);
nand U20956 (N_20956,N_18557,N_19086);
and U20957 (N_20957,N_18997,N_19712);
xnor U20958 (N_20958,N_19616,N_18501);
nand U20959 (N_20959,N_18529,N_19301);
nand U20960 (N_20960,N_19603,N_19638);
or U20961 (N_20961,N_18510,N_19647);
nor U20962 (N_20962,N_19826,N_19308);
nand U20963 (N_20963,N_18293,N_19359);
nor U20964 (N_20964,N_18882,N_19483);
xnor U20965 (N_20965,N_19412,N_19981);
or U20966 (N_20966,N_19900,N_19835);
nand U20967 (N_20967,N_18092,N_19079);
nand U20968 (N_20968,N_19004,N_19347);
or U20969 (N_20969,N_19723,N_19539);
nor U20970 (N_20970,N_19984,N_19038);
nor U20971 (N_20971,N_19776,N_18238);
and U20972 (N_20972,N_18534,N_18046);
xor U20973 (N_20973,N_18499,N_19280);
and U20974 (N_20974,N_18379,N_19207);
nand U20975 (N_20975,N_19452,N_18625);
nand U20976 (N_20976,N_18652,N_18839);
and U20977 (N_20977,N_18803,N_19272);
or U20978 (N_20978,N_19161,N_18730);
and U20979 (N_20979,N_19899,N_18918);
xor U20980 (N_20980,N_18198,N_19860);
and U20981 (N_20981,N_19494,N_18553);
nand U20982 (N_20982,N_18568,N_19249);
nor U20983 (N_20983,N_19593,N_18279);
xnor U20984 (N_20984,N_19502,N_18000);
or U20985 (N_20985,N_19609,N_18367);
and U20986 (N_20986,N_18881,N_19211);
or U20987 (N_20987,N_18849,N_18355);
nand U20988 (N_20988,N_18506,N_18298);
nand U20989 (N_20989,N_18932,N_19932);
and U20990 (N_20990,N_18097,N_18192);
nor U20991 (N_20991,N_18366,N_18375);
or U20992 (N_20992,N_18058,N_18322);
nand U20993 (N_20993,N_18654,N_19610);
and U20994 (N_20994,N_18287,N_18229);
or U20995 (N_20995,N_18178,N_19893);
or U20996 (N_20996,N_19065,N_18088);
or U20997 (N_20997,N_18969,N_18739);
nor U20998 (N_20998,N_19831,N_18540);
and U20999 (N_20999,N_19970,N_19879);
or U21000 (N_21000,N_19234,N_19155);
xor U21001 (N_21001,N_18150,N_19660);
and U21002 (N_21002,N_18283,N_19770);
xor U21003 (N_21003,N_18011,N_19263);
nor U21004 (N_21004,N_19981,N_18981);
or U21005 (N_21005,N_18616,N_18405);
nand U21006 (N_21006,N_19002,N_19882);
and U21007 (N_21007,N_19773,N_19737);
nand U21008 (N_21008,N_18816,N_19627);
nand U21009 (N_21009,N_19095,N_19737);
nor U21010 (N_21010,N_19155,N_19826);
nor U21011 (N_21011,N_19457,N_19562);
xor U21012 (N_21012,N_19749,N_18880);
and U21013 (N_21013,N_18163,N_19277);
and U21014 (N_21014,N_18514,N_19061);
and U21015 (N_21015,N_18907,N_18131);
and U21016 (N_21016,N_18130,N_19292);
nor U21017 (N_21017,N_18994,N_18960);
nand U21018 (N_21018,N_18542,N_18641);
nor U21019 (N_21019,N_19440,N_18772);
and U21020 (N_21020,N_18794,N_18672);
or U21021 (N_21021,N_19992,N_18171);
nor U21022 (N_21022,N_18496,N_18691);
or U21023 (N_21023,N_19306,N_18092);
nand U21024 (N_21024,N_19817,N_18626);
nand U21025 (N_21025,N_19684,N_19669);
or U21026 (N_21026,N_19379,N_18483);
nand U21027 (N_21027,N_19146,N_18038);
and U21028 (N_21028,N_19406,N_19794);
nand U21029 (N_21029,N_18452,N_19432);
xor U21030 (N_21030,N_19276,N_18749);
or U21031 (N_21031,N_18431,N_19707);
nand U21032 (N_21032,N_18716,N_18667);
or U21033 (N_21033,N_18339,N_19312);
nand U21034 (N_21034,N_18325,N_19482);
nand U21035 (N_21035,N_19564,N_19969);
or U21036 (N_21036,N_18977,N_19346);
or U21037 (N_21037,N_19578,N_19131);
nor U21038 (N_21038,N_18051,N_18746);
nor U21039 (N_21039,N_19279,N_19059);
or U21040 (N_21040,N_19659,N_19937);
or U21041 (N_21041,N_19349,N_19844);
nand U21042 (N_21042,N_18643,N_19495);
nor U21043 (N_21043,N_19866,N_19443);
nand U21044 (N_21044,N_19303,N_19658);
or U21045 (N_21045,N_19041,N_18448);
nand U21046 (N_21046,N_19157,N_19474);
nand U21047 (N_21047,N_18404,N_19427);
nand U21048 (N_21048,N_18540,N_18557);
nor U21049 (N_21049,N_18318,N_19584);
nor U21050 (N_21050,N_19682,N_18244);
nand U21051 (N_21051,N_19544,N_19977);
nor U21052 (N_21052,N_19850,N_18930);
nor U21053 (N_21053,N_18790,N_18662);
nand U21054 (N_21054,N_18815,N_18518);
xor U21055 (N_21055,N_18542,N_18138);
xor U21056 (N_21056,N_18580,N_18900);
or U21057 (N_21057,N_18490,N_18292);
xnor U21058 (N_21058,N_19691,N_18995);
nor U21059 (N_21059,N_19631,N_18696);
xnor U21060 (N_21060,N_18665,N_19860);
xor U21061 (N_21061,N_18722,N_18529);
nor U21062 (N_21062,N_18780,N_18996);
xor U21063 (N_21063,N_18937,N_19233);
nor U21064 (N_21064,N_19178,N_19408);
nor U21065 (N_21065,N_19084,N_19552);
and U21066 (N_21066,N_19121,N_19618);
xor U21067 (N_21067,N_19547,N_19352);
nor U21068 (N_21068,N_18680,N_18262);
nor U21069 (N_21069,N_18784,N_19891);
or U21070 (N_21070,N_19949,N_19615);
xor U21071 (N_21071,N_18418,N_19096);
xor U21072 (N_21072,N_19879,N_18326);
and U21073 (N_21073,N_19657,N_19662);
or U21074 (N_21074,N_19247,N_19101);
xnor U21075 (N_21075,N_18405,N_18350);
nor U21076 (N_21076,N_18147,N_19454);
xor U21077 (N_21077,N_19637,N_19440);
xor U21078 (N_21078,N_18080,N_19749);
and U21079 (N_21079,N_18545,N_19791);
or U21080 (N_21080,N_18400,N_19921);
nor U21081 (N_21081,N_19928,N_18863);
nor U21082 (N_21082,N_18695,N_19834);
xnor U21083 (N_21083,N_19515,N_18572);
nor U21084 (N_21084,N_19311,N_19514);
xor U21085 (N_21085,N_18614,N_18018);
nor U21086 (N_21086,N_19498,N_18946);
xnor U21087 (N_21087,N_19155,N_19250);
nor U21088 (N_21088,N_18329,N_18771);
nand U21089 (N_21089,N_18839,N_19907);
or U21090 (N_21090,N_19169,N_19415);
nand U21091 (N_21091,N_18034,N_19421);
nand U21092 (N_21092,N_18092,N_18719);
nor U21093 (N_21093,N_19291,N_18085);
xnor U21094 (N_21094,N_18314,N_18562);
nand U21095 (N_21095,N_19090,N_19076);
or U21096 (N_21096,N_19515,N_18887);
nor U21097 (N_21097,N_19506,N_18187);
nor U21098 (N_21098,N_19090,N_19069);
and U21099 (N_21099,N_18124,N_18963);
and U21100 (N_21100,N_19576,N_19480);
nand U21101 (N_21101,N_18763,N_18273);
or U21102 (N_21102,N_18531,N_19402);
and U21103 (N_21103,N_19311,N_18825);
or U21104 (N_21104,N_19781,N_18327);
and U21105 (N_21105,N_19834,N_18589);
nand U21106 (N_21106,N_18002,N_18631);
and U21107 (N_21107,N_18333,N_19674);
and U21108 (N_21108,N_19915,N_18701);
nor U21109 (N_21109,N_19056,N_19382);
or U21110 (N_21110,N_19632,N_19898);
nor U21111 (N_21111,N_18602,N_19426);
xnor U21112 (N_21112,N_19883,N_19525);
nor U21113 (N_21113,N_18597,N_19185);
nand U21114 (N_21114,N_19274,N_18759);
nand U21115 (N_21115,N_18014,N_19910);
or U21116 (N_21116,N_18824,N_18743);
xnor U21117 (N_21117,N_19212,N_18469);
nor U21118 (N_21118,N_18076,N_19870);
nor U21119 (N_21119,N_19555,N_18056);
xor U21120 (N_21120,N_18239,N_19272);
or U21121 (N_21121,N_18734,N_18282);
or U21122 (N_21122,N_19691,N_19988);
and U21123 (N_21123,N_19939,N_19208);
xnor U21124 (N_21124,N_18518,N_18980);
xnor U21125 (N_21125,N_18607,N_19041);
nand U21126 (N_21126,N_18607,N_18585);
xor U21127 (N_21127,N_18210,N_19180);
or U21128 (N_21128,N_19351,N_18983);
and U21129 (N_21129,N_18948,N_19683);
nand U21130 (N_21130,N_19907,N_18819);
and U21131 (N_21131,N_18919,N_18773);
xnor U21132 (N_21132,N_18762,N_18057);
xor U21133 (N_21133,N_18577,N_18806);
and U21134 (N_21134,N_19245,N_19667);
or U21135 (N_21135,N_18389,N_18246);
nand U21136 (N_21136,N_18271,N_19352);
and U21137 (N_21137,N_18566,N_19406);
xnor U21138 (N_21138,N_18251,N_18117);
or U21139 (N_21139,N_18638,N_18901);
nor U21140 (N_21140,N_19418,N_18226);
xor U21141 (N_21141,N_18025,N_19628);
nand U21142 (N_21142,N_18224,N_18890);
xnor U21143 (N_21143,N_18335,N_19013);
nand U21144 (N_21144,N_19454,N_18814);
nand U21145 (N_21145,N_19611,N_19600);
and U21146 (N_21146,N_18486,N_19967);
xor U21147 (N_21147,N_19445,N_18116);
nand U21148 (N_21148,N_19500,N_18376);
or U21149 (N_21149,N_19757,N_18355);
or U21150 (N_21150,N_18338,N_18606);
xor U21151 (N_21151,N_19609,N_19451);
and U21152 (N_21152,N_19324,N_19638);
or U21153 (N_21153,N_18422,N_18789);
xnor U21154 (N_21154,N_18094,N_19443);
and U21155 (N_21155,N_19735,N_19527);
or U21156 (N_21156,N_18890,N_19217);
xnor U21157 (N_21157,N_19816,N_18631);
xor U21158 (N_21158,N_19221,N_19189);
nand U21159 (N_21159,N_19061,N_18286);
nor U21160 (N_21160,N_19828,N_18590);
or U21161 (N_21161,N_19250,N_19333);
nand U21162 (N_21162,N_19486,N_18002);
or U21163 (N_21163,N_18821,N_18685);
nand U21164 (N_21164,N_19988,N_18694);
or U21165 (N_21165,N_18423,N_19379);
nor U21166 (N_21166,N_18649,N_19976);
nor U21167 (N_21167,N_18282,N_18125);
nand U21168 (N_21168,N_19793,N_19756);
nand U21169 (N_21169,N_19882,N_19962);
xor U21170 (N_21170,N_18962,N_18111);
xnor U21171 (N_21171,N_19063,N_19179);
nand U21172 (N_21172,N_18192,N_18782);
or U21173 (N_21173,N_18807,N_19805);
nor U21174 (N_21174,N_19822,N_19433);
nor U21175 (N_21175,N_19536,N_19613);
nor U21176 (N_21176,N_18112,N_18438);
nor U21177 (N_21177,N_18465,N_18610);
and U21178 (N_21178,N_19248,N_19947);
xor U21179 (N_21179,N_19658,N_19848);
nand U21180 (N_21180,N_19858,N_19314);
or U21181 (N_21181,N_19194,N_18377);
or U21182 (N_21182,N_19224,N_18586);
nand U21183 (N_21183,N_19523,N_19327);
and U21184 (N_21184,N_19641,N_19109);
or U21185 (N_21185,N_19127,N_18244);
or U21186 (N_21186,N_19514,N_18414);
and U21187 (N_21187,N_19191,N_18012);
or U21188 (N_21188,N_18377,N_18412);
and U21189 (N_21189,N_18751,N_18940);
and U21190 (N_21190,N_18450,N_19659);
and U21191 (N_21191,N_19691,N_18982);
and U21192 (N_21192,N_19752,N_19212);
and U21193 (N_21193,N_19930,N_19563);
or U21194 (N_21194,N_19383,N_19962);
nand U21195 (N_21195,N_18127,N_19720);
and U21196 (N_21196,N_18669,N_18228);
nor U21197 (N_21197,N_19471,N_19745);
or U21198 (N_21198,N_18921,N_19388);
xnor U21199 (N_21199,N_19274,N_18591);
and U21200 (N_21200,N_19637,N_19192);
xnor U21201 (N_21201,N_19458,N_19044);
or U21202 (N_21202,N_19504,N_18536);
or U21203 (N_21203,N_19388,N_18588);
or U21204 (N_21204,N_19272,N_19143);
or U21205 (N_21205,N_18883,N_19410);
nand U21206 (N_21206,N_19364,N_18219);
or U21207 (N_21207,N_18642,N_19792);
nor U21208 (N_21208,N_18737,N_19410);
nor U21209 (N_21209,N_18151,N_18032);
nor U21210 (N_21210,N_19050,N_18885);
nor U21211 (N_21211,N_18268,N_18972);
nor U21212 (N_21212,N_19800,N_18802);
xnor U21213 (N_21213,N_19972,N_18255);
nand U21214 (N_21214,N_18263,N_19054);
or U21215 (N_21215,N_19476,N_19522);
nand U21216 (N_21216,N_19498,N_19283);
nand U21217 (N_21217,N_19786,N_18232);
nor U21218 (N_21218,N_18245,N_18929);
xnor U21219 (N_21219,N_18553,N_18674);
and U21220 (N_21220,N_19426,N_18109);
nand U21221 (N_21221,N_19828,N_19938);
and U21222 (N_21222,N_19521,N_19979);
nor U21223 (N_21223,N_19380,N_19078);
or U21224 (N_21224,N_19993,N_18203);
nor U21225 (N_21225,N_19687,N_18461);
nand U21226 (N_21226,N_18714,N_19615);
nand U21227 (N_21227,N_18870,N_19072);
and U21228 (N_21228,N_18570,N_18121);
and U21229 (N_21229,N_18276,N_19846);
nand U21230 (N_21230,N_19058,N_18818);
nor U21231 (N_21231,N_18510,N_18178);
and U21232 (N_21232,N_18490,N_19751);
xnor U21233 (N_21233,N_18766,N_18247);
nor U21234 (N_21234,N_19827,N_19846);
xor U21235 (N_21235,N_18101,N_18882);
nor U21236 (N_21236,N_19056,N_19100);
nor U21237 (N_21237,N_19248,N_19253);
nand U21238 (N_21238,N_19296,N_18179);
nand U21239 (N_21239,N_18150,N_19765);
or U21240 (N_21240,N_18046,N_18715);
nand U21241 (N_21241,N_18568,N_19895);
nand U21242 (N_21242,N_18840,N_18015);
or U21243 (N_21243,N_19621,N_18772);
or U21244 (N_21244,N_19529,N_18568);
nor U21245 (N_21245,N_19863,N_19664);
nand U21246 (N_21246,N_18069,N_19832);
xnor U21247 (N_21247,N_19723,N_18403);
nand U21248 (N_21248,N_18091,N_19448);
nand U21249 (N_21249,N_18328,N_18097);
or U21250 (N_21250,N_18586,N_18543);
nor U21251 (N_21251,N_18889,N_18019);
or U21252 (N_21252,N_18282,N_18848);
or U21253 (N_21253,N_19320,N_18898);
or U21254 (N_21254,N_19604,N_18387);
nand U21255 (N_21255,N_18804,N_18604);
xnor U21256 (N_21256,N_18241,N_19572);
and U21257 (N_21257,N_19838,N_19111);
nand U21258 (N_21258,N_19995,N_18750);
nor U21259 (N_21259,N_18360,N_19758);
nor U21260 (N_21260,N_18743,N_18554);
xor U21261 (N_21261,N_18156,N_18210);
and U21262 (N_21262,N_18507,N_19184);
and U21263 (N_21263,N_18828,N_19362);
nand U21264 (N_21264,N_19740,N_18039);
nor U21265 (N_21265,N_18822,N_19334);
or U21266 (N_21266,N_18940,N_19409);
and U21267 (N_21267,N_18523,N_19726);
nand U21268 (N_21268,N_18875,N_18540);
or U21269 (N_21269,N_18312,N_19176);
nor U21270 (N_21270,N_19906,N_19764);
nor U21271 (N_21271,N_19106,N_18289);
nor U21272 (N_21272,N_18969,N_19812);
nor U21273 (N_21273,N_19434,N_18991);
and U21274 (N_21274,N_19132,N_19419);
nor U21275 (N_21275,N_19078,N_19420);
and U21276 (N_21276,N_19378,N_18210);
and U21277 (N_21277,N_18839,N_18515);
and U21278 (N_21278,N_19129,N_18792);
nand U21279 (N_21279,N_18778,N_19473);
nand U21280 (N_21280,N_18023,N_18482);
xor U21281 (N_21281,N_18903,N_19791);
nor U21282 (N_21282,N_19757,N_18710);
nand U21283 (N_21283,N_18807,N_19723);
and U21284 (N_21284,N_19793,N_18290);
or U21285 (N_21285,N_18847,N_19410);
and U21286 (N_21286,N_19186,N_19827);
or U21287 (N_21287,N_19763,N_19044);
xor U21288 (N_21288,N_19143,N_18686);
nor U21289 (N_21289,N_18457,N_18991);
and U21290 (N_21290,N_18177,N_18613);
nor U21291 (N_21291,N_19163,N_19395);
or U21292 (N_21292,N_19752,N_19278);
or U21293 (N_21293,N_19365,N_18993);
xor U21294 (N_21294,N_18428,N_19536);
xor U21295 (N_21295,N_19477,N_18254);
xor U21296 (N_21296,N_18354,N_19293);
and U21297 (N_21297,N_18289,N_18785);
and U21298 (N_21298,N_19796,N_18371);
nor U21299 (N_21299,N_18507,N_18882);
and U21300 (N_21300,N_18999,N_18089);
nor U21301 (N_21301,N_18830,N_18679);
xor U21302 (N_21302,N_18794,N_19308);
and U21303 (N_21303,N_18537,N_19146);
and U21304 (N_21304,N_19017,N_19810);
xnor U21305 (N_21305,N_18836,N_19425);
and U21306 (N_21306,N_19680,N_19219);
or U21307 (N_21307,N_19280,N_18319);
and U21308 (N_21308,N_19431,N_19891);
nand U21309 (N_21309,N_18400,N_19815);
xor U21310 (N_21310,N_19513,N_19279);
and U21311 (N_21311,N_18798,N_19022);
xnor U21312 (N_21312,N_18300,N_18218);
xnor U21313 (N_21313,N_18399,N_19434);
or U21314 (N_21314,N_18165,N_18329);
nor U21315 (N_21315,N_18647,N_18755);
nand U21316 (N_21316,N_19470,N_18181);
and U21317 (N_21317,N_19668,N_18791);
nand U21318 (N_21318,N_18176,N_18437);
nor U21319 (N_21319,N_19439,N_19739);
or U21320 (N_21320,N_19845,N_18099);
or U21321 (N_21321,N_18576,N_18824);
nand U21322 (N_21322,N_18887,N_18637);
nand U21323 (N_21323,N_19228,N_18389);
or U21324 (N_21324,N_19396,N_19855);
and U21325 (N_21325,N_18097,N_18748);
or U21326 (N_21326,N_18896,N_19489);
and U21327 (N_21327,N_19167,N_18277);
and U21328 (N_21328,N_19323,N_18566);
xor U21329 (N_21329,N_18610,N_18239);
nand U21330 (N_21330,N_19221,N_18480);
xor U21331 (N_21331,N_18538,N_19609);
or U21332 (N_21332,N_19984,N_19192);
nor U21333 (N_21333,N_19029,N_19217);
and U21334 (N_21334,N_19388,N_18500);
nand U21335 (N_21335,N_19498,N_19513);
and U21336 (N_21336,N_18074,N_18580);
nand U21337 (N_21337,N_18928,N_18656);
xnor U21338 (N_21338,N_19376,N_18503);
or U21339 (N_21339,N_19270,N_18228);
nand U21340 (N_21340,N_19796,N_18679);
or U21341 (N_21341,N_19196,N_19805);
nand U21342 (N_21342,N_18265,N_18332);
and U21343 (N_21343,N_19508,N_18849);
nor U21344 (N_21344,N_19817,N_18379);
nand U21345 (N_21345,N_19430,N_19262);
nand U21346 (N_21346,N_18760,N_18973);
and U21347 (N_21347,N_18393,N_19602);
or U21348 (N_21348,N_19020,N_18076);
nand U21349 (N_21349,N_18469,N_19646);
xor U21350 (N_21350,N_19600,N_19630);
or U21351 (N_21351,N_19245,N_18435);
or U21352 (N_21352,N_18826,N_19941);
xor U21353 (N_21353,N_18756,N_18714);
xnor U21354 (N_21354,N_18416,N_18435);
nor U21355 (N_21355,N_19242,N_19804);
xor U21356 (N_21356,N_18818,N_19462);
and U21357 (N_21357,N_18094,N_19504);
and U21358 (N_21358,N_19063,N_18834);
or U21359 (N_21359,N_19376,N_18458);
xnor U21360 (N_21360,N_19150,N_18971);
and U21361 (N_21361,N_18719,N_18123);
nor U21362 (N_21362,N_19108,N_19640);
nand U21363 (N_21363,N_18836,N_19024);
xor U21364 (N_21364,N_19768,N_19038);
and U21365 (N_21365,N_18722,N_19922);
or U21366 (N_21366,N_19424,N_18117);
xnor U21367 (N_21367,N_18871,N_19184);
and U21368 (N_21368,N_19192,N_19767);
nor U21369 (N_21369,N_18931,N_19479);
nand U21370 (N_21370,N_19400,N_19399);
nor U21371 (N_21371,N_19334,N_19327);
nor U21372 (N_21372,N_19509,N_19143);
nor U21373 (N_21373,N_19633,N_18239);
and U21374 (N_21374,N_19721,N_18596);
and U21375 (N_21375,N_18478,N_19232);
nor U21376 (N_21376,N_19294,N_18198);
or U21377 (N_21377,N_19413,N_19237);
and U21378 (N_21378,N_19763,N_19007);
and U21379 (N_21379,N_18287,N_18601);
or U21380 (N_21380,N_18052,N_19200);
and U21381 (N_21381,N_18093,N_18935);
or U21382 (N_21382,N_19711,N_19270);
and U21383 (N_21383,N_19008,N_19579);
or U21384 (N_21384,N_18123,N_19659);
and U21385 (N_21385,N_18157,N_19608);
or U21386 (N_21386,N_18933,N_18704);
nand U21387 (N_21387,N_19323,N_19690);
xnor U21388 (N_21388,N_18690,N_18669);
nand U21389 (N_21389,N_19602,N_19258);
nand U21390 (N_21390,N_19517,N_18038);
and U21391 (N_21391,N_18269,N_19417);
and U21392 (N_21392,N_19158,N_18077);
nor U21393 (N_21393,N_18404,N_19696);
nand U21394 (N_21394,N_18493,N_19293);
xnor U21395 (N_21395,N_19499,N_19734);
nor U21396 (N_21396,N_18097,N_18899);
nand U21397 (N_21397,N_19641,N_19895);
nand U21398 (N_21398,N_19124,N_18917);
and U21399 (N_21399,N_18038,N_18054);
or U21400 (N_21400,N_19921,N_19013);
or U21401 (N_21401,N_19542,N_18377);
nor U21402 (N_21402,N_19957,N_19363);
xnor U21403 (N_21403,N_19028,N_18372);
nor U21404 (N_21404,N_18829,N_18853);
xnor U21405 (N_21405,N_19251,N_18166);
or U21406 (N_21406,N_19806,N_19753);
nor U21407 (N_21407,N_19752,N_19949);
nor U21408 (N_21408,N_18926,N_18345);
and U21409 (N_21409,N_18323,N_18241);
and U21410 (N_21410,N_19883,N_18939);
and U21411 (N_21411,N_18016,N_19296);
xor U21412 (N_21412,N_18242,N_19360);
xor U21413 (N_21413,N_18007,N_19826);
or U21414 (N_21414,N_18971,N_18391);
and U21415 (N_21415,N_18868,N_18904);
xor U21416 (N_21416,N_18367,N_18981);
nor U21417 (N_21417,N_19040,N_18146);
xnor U21418 (N_21418,N_18960,N_19965);
nand U21419 (N_21419,N_18923,N_19901);
nor U21420 (N_21420,N_19629,N_19623);
or U21421 (N_21421,N_18454,N_19416);
nand U21422 (N_21422,N_19595,N_18551);
nor U21423 (N_21423,N_18712,N_18340);
or U21424 (N_21424,N_19825,N_19504);
nor U21425 (N_21425,N_19902,N_19989);
xnor U21426 (N_21426,N_18493,N_19645);
or U21427 (N_21427,N_19189,N_18770);
nor U21428 (N_21428,N_18648,N_19494);
or U21429 (N_21429,N_18170,N_19943);
nand U21430 (N_21430,N_19471,N_19578);
nand U21431 (N_21431,N_19140,N_18862);
and U21432 (N_21432,N_18037,N_19502);
nor U21433 (N_21433,N_19423,N_19996);
nand U21434 (N_21434,N_18875,N_19460);
xnor U21435 (N_21435,N_19498,N_18579);
or U21436 (N_21436,N_19937,N_19657);
xnor U21437 (N_21437,N_19320,N_18793);
or U21438 (N_21438,N_18757,N_18516);
and U21439 (N_21439,N_19554,N_19790);
nor U21440 (N_21440,N_19661,N_19253);
or U21441 (N_21441,N_19147,N_18827);
and U21442 (N_21442,N_19694,N_19875);
xor U21443 (N_21443,N_19023,N_19485);
or U21444 (N_21444,N_19807,N_19406);
nand U21445 (N_21445,N_18101,N_19542);
xnor U21446 (N_21446,N_19657,N_19552);
nand U21447 (N_21447,N_19723,N_19739);
xor U21448 (N_21448,N_18708,N_19999);
nor U21449 (N_21449,N_18843,N_19560);
nand U21450 (N_21450,N_19534,N_19253);
nor U21451 (N_21451,N_19798,N_19272);
or U21452 (N_21452,N_18804,N_19818);
or U21453 (N_21453,N_19115,N_19208);
nand U21454 (N_21454,N_18305,N_19606);
nand U21455 (N_21455,N_18187,N_19053);
nor U21456 (N_21456,N_18171,N_19777);
or U21457 (N_21457,N_18041,N_19966);
and U21458 (N_21458,N_18666,N_19924);
nand U21459 (N_21459,N_18095,N_18459);
nor U21460 (N_21460,N_18363,N_18800);
nor U21461 (N_21461,N_18512,N_18309);
nand U21462 (N_21462,N_18758,N_18262);
nand U21463 (N_21463,N_18228,N_19849);
nor U21464 (N_21464,N_19935,N_18338);
nor U21465 (N_21465,N_19951,N_18023);
xor U21466 (N_21466,N_18722,N_19852);
or U21467 (N_21467,N_18794,N_18598);
nand U21468 (N_21468,N_19057,N_18650);
xnor U21469 (N_21469,N_18754,N_19534);
xnor U21470 (N_21470,N_19194,N_19995);
nor U21471 (N_21471,N_18995,N_19478);
nand U21472 (N_21472,N_19352,N_19398);
or U21473 (N_21473,N_18580,N_18739);
and U21474 (N_21474,N_18454,N_18191);
and U21475 (N_21475,N_18027,N_18846);
or U21476 (N_21476,N_19950,N_18582);
nor U21477 (N_21477,N_19649,N_19820);
nor U21478 (N_21478,N_19975,N_19102);
and U21479 (N_21479,N_19242,N_19960);
and U21480 (N_21480,N_19687,N_18457);
xor U21481 (N_21481,N_19047,N_19481);
xnor U21482 (N_21482,N_19468,N_19612);
nor U21483 (N_21483,N_18162,N_18506);
nor U21484 (N_21484,N_19911,N_19313);
nand U21485 (N_21485,N_18527,N_18404);
xor U21486 (N_21486,N_19951,N_19168);
and U21487 (N_21487,N_19316,N_19662);
or U21488 (N_21488,N_19858,N_19562);
and U21489 (N_21489,N_18497,N_18466);
nor U21490 (N_21490,N_18173,N_18635);
and U21491 (N_21491,N_19750,N_18727);
nand U21492 (N_21492,N_19281,N_18477);
nor U21493 (N_21493,N_18686,N_19527);
nand U21494 (N_21494,N_19023,N_19639);
and U21495 (N_21495,N_18217,N_18324);
or U21496 (N_21496,N_19256,N_19409);
nor U21497 (N_21497,N_18191,N_18331);
or U21498 (N_21498,N_19743,N_18397);
or U21499 (N_21499,N_18379,N_19460);
and U21500 (N_21500,N_18117,N_19629);
nand U21501 (N_21501,N_19338,N_19459);
nor U21502 (N_21502,N_18932,N_19163);
or U21503 (N_21503,N_19310,N_18660);
nand U21504 (N_21504,N_18564,N_18982);
nor U21505 (N_21505,N_18002,N_19463);
xor U21506 (N_21506,N_19289,N_18977);
xnor U21507 (N_21507,N_19651,N_19707);
nand U21508 (N_21508,N_19918,N_18399);
or U21509 (N_21509,N_19619,N_19941);
nor U21510 (N_21510,N_19510,N_19317);
nand U21511 (N_21511,N_19358,N_18444);
and U21512 (N_21512,N_19923,N_18148);
xnor U21513 (N_21513,N_19103,N_18825);
nor U21514 (N_21514,N_19119,N_18254);
or U21515 (N_21515,N_18877,N_19801);
or U21516 (N_21516,N_18494,N_18624);
xor U21517 (N_21517,N_19164,N_19432);
xor U21518 (N_21518,N_18707,N_18236);
nand U21519 (N_21519,N_18393,N_18906);
nand U21520 (N_21520,N_18983,N_18463);
and U21521 (N_21521,N_19404,N_18072);
nand U21522 (N_21522,N_19203,N_19218);
or U21523 (N_21523,N_18393,N_18027);
or U21524 (N_21524,N_18874,N_19478);
nand U21525 (N_21525,N_18463,N_19020);
xor U21526 (N_21526,N_18508,N_19347);
nand U21527 (N_21527,N_19495,N_18139);
nor U21528 (N_21528,N_19818,N_19651);
xor U21529 (N_21529,N_19549,N_19224);
and U21530 (N_21530,N_18549,N_18551);
xnor U21531 (N_21531,N_19597,N_18757);
or U21532 (N_21532,N_19182,N_19119);
or U21533 (N_21533,N_18235,N_19551);
nor U21534 (N_21534,N_19284,N_18577);
nor U21535 (N_21535,N_18537,N_18349);
and U21536 (N_21536,N_18700,N_18377);
xnor U21537 (N_21537,N_18675,N_19433);
nor U21538 (N_21538,N_19955,N_18497);
or U21539 (N_21539,N_18877,N_19575);
xor U21540 (N_21540,N_19015,N_18050);
nand U21541 (N_21541,N_19864,N_19931);
nand U21542 (N_21542,N_18364,N_19165);
and U21543 (N_21543,N_19016,N_18018);
or U21544 (N_21544,N_18029,N_18184);
xnor U21545 (N_21545,N_19875,N_18879);
and U21546 (N_21546,N_18467,N_19698);
and U21547 (N_21547,N_19089,N_19315);
or U21548 (N_21548,N_18436,N_19035);
nor U21549 (N_21549,N_18828,N_18334);
nand U21550 (N_21550,N_18646,N_19860);
nand U21551 (N_21551,N_18145,N_19578);
nor U21552 (N_21552,N_18812,N_18728);
xor U21553 (N_21553,N_18658,N_19756);
or U21554 (N_21554,N_19025,N_18984);
or U21555 (N_21555,N_18686,N_18847);
nand U21556 (N_21556,N_19092,N_18885);
or U21557 (N_21557,N_19393,N_18475);
or U21558 (N_21558,N_19144,N_19126);
nand U21559 (N_21559,N_18326,N_19179);
or U21560 (N_21560,N_18176,N_18964);
xor U21561 (N_21561,N_18613,N_18428);
and U21562 (N_21562,N_19545,N_19941);
or U21563 (N_21563,N_18762,N_19411);
and U21564 (N_21564,N_19844,N_19782);
nor U21565 (N_21565,N_18954,N_19486);
and U21566 (N_21566,N_19146,N_19616);
and U21567 (N_21567,N_18294,N_19628);
or U21568 (N_21568,N_19858,N_18537);
xnor U21569 (N_21569,N_18283,N_19355);
xnor U21570 (N_21570,N_18141,N_18204);
nor U21571 (N_21571,N_18663,N_19839);
and U21572 (N_21572,N_18868,N_18700);
xor U21573 (N_21573,N_18297,N_19910);
nor U21574 (N_21574,N_19423,N_18792);
or U21575 (N_21575,N_19957,N_19270);
nand U21576 (N_21576,N_18599,N_19217);
or U21577 (N_21577,N_19912,N_18644);
nor U21578 (N_21578,N_18814,N_18905);
nor U21579 (N_21579,N_19375,N_19701);
xnor U21580 (N_21580,N_19553,N_19083);
nor U21581 (N_21581,N_19984,N_18593);
nand U21582 (N_21582,N_19588,N_19609);
and U21583 (N_21583,N_18050,N_18964);
or U21584 (N_21584,N_18954,N_18080);
xnor U21585 (N_21585,N_18604,N_19641);
xnor U21586 (N_21586,N_18807,N_19713);
nand U21587 (N_21587,N_19119,N_19748);
and U21588 (N_21588,N_19832,N_19976);
and U21589 (N_21589,N_19591,N_18892);
nand U21590 (N_21590,N_19659,N_18392);
xor U21591 (N_21591,N_19283,N_18887);
and U21592 (N_21592,N_19695,N_19266);
and U21593 (N_21593,N_19992,N_19759);
xor U21594 (N_21594,N_19054,N_18437);
nor U21595 (N_21595,N_18610,N_18387);
or U21596 (N_21596,N_18580,N_18081);
nor U21597 (N_21597,N_18889,N_19459);
or U21598 (N_21598,N_18413,N_18451);
nor U21599 (N_21599,N_18587,N_18471);
and U21600 (N_21600,N_19959,N_19875);
or U21601 (N_21601,N_18789,N_19082);
nor U21602 (N_21602,N_19550,N_18762);
nor U21603 (N_21603,N_18511,N_18279);
or U21604 (N_21604,N_19206,N_18519);
nor U21605 (N_21605,N_18431,N_18564);
or U21606 (N_21606,N_19029,N_18785);
or U21607 (N_21607,N_19848,N_18906);
nand U21608 (N_21608,N_18282,N_18104);
xnor U21609 (N_21609,N_18068,N_18942);
nand U21610 (N_21610,N_18352,N_18334);
nand U21611 (N_21611,N_19213,N_19657);
or U21612 (N_21612,N_19690,N_19107);
or U21613 (N_21613,N_18298,N_18777);
and U21614 (N_21614,N_18150,N_19825);
nor U21615 (N_21615,N_18725,N_19255);
nand U21616 (N_21616,N_19992,N_19348);
and U21617 (N_21617,N_18343,N_18465);
nand U21618 (N_21618,N_18786,N_19976);
nor U21619 (N_21619,N_19132,N_18656);
nor U21620 (N_21620,N_19370,N_18287);
nand U21621 (N_21621,N_18592,N_18397);
xor U21622 (N_21622,N_19188,N_18705);
or U21623 (N_21623,N_19664,N_18088);
and U21624 (N_21624,N_19883,N_19980);
xor U21625 (N_21625,N_19146,N_19064);
or U21626 (N_21626,N_18398,N_19483);
nand U21627 (N_21627,N_18097,N_18070);
nand U21628 (N_21628,N_19128,N_19191);
or U21629 (N_21629,N_19735,N_19284);
or U21630 (N_21630,N_18311,N_19589);
and U21631 (N_21631,N_19991,N_18255);
and U21632 (N_21632,N_19907,N_19008);
xnor U21633 (N_21633,N_19640,N_18707);
nor U21634 (N_21634,N_19168,N_18707);
xor U21635 (N_21635,N_18326,N_19187);
nor U21636 (N_21636,N_19918,N_18395);
nand U21637 (N_21637,N_19834,N_18889);
nand U21638 (N_21638,N_19031,N_19416);
xnor U21639 (N_21639,N_18338,N_19272);
nor U21640 (N_21640,N_18075,N_18789);
or U21641 (N_21641,N_19034,N_18239);
xor U21642 (N_21642,N_18376,N_18699);
xor U21643 (N_21643,N_19794,N_19513);
nor U21644 (N_21644,N_19220,N_19791);
and U21645 (N_21645,N_19147,N_19229);
nand U21646 (N_21646,N_18137,N_19837);
nand U21647 (N_21647,N_18336,N_18398);
nand U21648 (N_21648,N_18084,N_19877);
xnor U21649 (N_21649,N_18995,N_18758);
xnor U21650 (N_21650,N_19652,N_19561);
nor U21651 (N_21651,N_18489,N_18163);
nor U21652 (N_21652,N_18924,N_18411);
nand U21653 (N_21653,N_19744,N_19597);
xnor U21654 (N_21654,N_19275,N_18975);
or U21655 (N_21655,N_18532,N_18975);
xor U21656 (N_21656,N_18533,N_18774);
nor U21657 (N_21657,N_18036,N_19265);
nor U21658 (N_21658,N_19809,N_19020);
xor U21659 (N_21659,N_19504,N_18147);
or U21660 (N_21660,N_19104,N_19477);
or U21661 (N_21661,N_18110,N_18849);
nand U21662 (N_21662,N_19716,N_19862);
nand U21663 (N_21663,N_19645,N_19966);
and U21664 (N_21664,N_19501,N_18498);
nand U21665 (N_21665,N_19699,N_19000);
and U21666 (N_21666,N_18689,N_18082);
nor U21667 (N_21667,N_18661,N_18107);
nor U21668 (N_21668,N_19089,N_19286);
and U21669 (N_21669,N_18905,N_19008);
nor U21670 (N_21670,N_18787,N_19517);
or U21671 (N_21671,N_19180,N_19234);
or U21672 (N_21672,N_18916,N_18375);
nor U21673 (N_21673,N_18598,N_19666);
nor U21674 (N_21674,N_18206,N_19456);
xor U21675 (N_21675,N_18222,N_18456);
and U21676 (N_21676,N_19280,N_19684);
or U21677 (N_21677,N_18606,N_19919);
xnor U21678 (N_21678,N_19161,N_18857);
nor U21679 (N_21679,N_18722,N_18949);
xnor U21680 (N_21680,N_19490,N_18255);
nor U21681 (N_21681,N_18229,N_18519);
xor U21682 (N_21682,N_18275,N_19394);
and U21683 (N_21683,N_18697,N_18183);
xor U21684 (N_21684,N_19359,N_19012);
xor U21685 (N_21685,N_19410,N_18015);
and U21686 (N_21686,N_18885,N_18634);
and U21687 (N_21687,N_18262,N_19634);
nand U21688 (N_21688,N_18619,N_19321);
and U21689 (N_21689,N_19348,N_18098);
and U21690 (N_21690,N_18874,N_19596);
xnor U21691 (N_21691,N_19510,N_18457);
nor U21692 (N_21692,N_19495,N_18628);
and U21693 (N_21693,N_18240,N_18372);
or U21694 (N_21694,N_19637,N_19550);
nor U21695 (N_21695,N_19368,N_18385);
xnor U21696 (N_21696,N_19874,N_18171);
nand U21697 (N_21697,N_18206,N_19543);
xnor U21698 (N_21698,N_18142,N_19051);
xnor U21699 (N_21699,N_18514,N_18420);
nand U21700 (N_21700,N_19421,N_19246);
nand U21701 (N_21701,N_19592,N_19402);
or U21702 (N_21702,N_19635,N_18972);
or U21703 (N_21703,N_18529,N_19922);
nand U21704 (N_21704,N_19307,N_18863);
xnor U21705 (N_21705,N_19999,N_19531);
xnor U21706 (N_21706,N_18985,N_19868);
nor U21707 (N_21707,N_18144,N_18467);
xnor U21708 (N_21708,N_18777,N_19318);
and U21709 (N_21709,N_18554,N_18868);
nor U21710 (N_21710,N_18581,N_19240);
nand U21711 (N_21711,N_18580,N_18451);
xnor U21712 (N_21712,N_19325,N_18783);
and U21713 (N_21713,N_18103,N_19552);
xor U21714 (N_21714,N_18435,N_18668);
nor U21715 (N_21715,N_18706,N_19717);
nor U21716 (N_21716,N_18997,N_19860);
or U21717 (N_21717,N_19170,N_19012);
and U21718 (N_21718,N_18317,N_19145);
and U21719 (N_21719,N_18829,N_19809);
nor U21720 (N_21720,N_19893,N_19082);
nand U21721 (N_21721,N_18748,N_18558);
xor U21722 (N_21722,N_18760,N_19326);
nor U21723 (N_21723,N_19633,N_19650);
or U21724 (N_21724,N_18859,N_19410);
or U21725 (N_21725,N_18720,N_19463);
xor U21726 (N_21726,N_19177,N_19597);
xnor U21727 (N_21727,N_19775,N_18235);
nor U21728 (N_21728,N_18293,N_19980);
nor U21729 (N_21729,N_18725,N_19773);
nand U21730 (N_21730,N_19218,N_18259);
or U21731 (N_21731,N_19229,N_18177);
nand U21732 (N_21732,N_18427,N_19595);
or U21733 (N_21733,N_19028,N_18887);
nor U21734 (N_21734,N_18518,N_19761);
and U21735 (N_21735,N_19057,N_19639);
or U21736 (N_21736,N_19867,N_19411);
or U21737 (N_21737,N_19575,N_18860);
nand U21738 (N_21738,N_18317,N_19756);
xor U21739 (N_21739,N_19513,N_18814);
and U21740 (N_21740,N_19787,N_19575);
nand U21741 (N_21741,N_19983,N_18948);
nor U21742 (N_21742,N_18159,N_18495);
nand U21743 (N_21743,N_19993,N_19452);
and U21744 (N_21744,N_18114,N_18167);
xor U21745 (N_21745,N_19689,N_18560);
xor U21746 (N_21746,N_18294,N_18864);
and U21747 (N_21747,N_18488,N_19605);
nand U21748 (N_21748,N_18931,N_19809);
and U21749 (N_21749,N_19302,N_19065);
nand U21750 (N_21750,N_19713,N_19771);
or U21751 (N_21751,N_18160,N_18815);
nand U21752 (N_21752,N_18731,N_18551);
nor U21753 (N_21753,N_18949,N_18153);
nand U21754 (N_21754,N_19954,N_19380);
nor U21755 (N_21755,N_18988,N_18626);
nand U21756 (N_21756,N_19459,N_19013);
nor U21757 (N_21757,N_19982,N_18442);
nor U21758 (N_21758,N_19199,N_19444);
and U21759 (N_21759,N_19228,N_19142);
nor U21760 (N_21760,N_19672,N_19860);
xor U21761 (N_21761,N_18683,N_18705);
and U21762 (N_21762,N_18643,N_18060);
nand U21763 (N_21763,N_19274,N_19334);
or U21764 (N_21764,N_19549,N_18655);
or U21765 (N_21765,N_19897,N_19836);
xnor U21766 (N_21766,N_19528,N_18371);
and U21767 (N_21767,N_18198,N_19076);
or U21768 (N_21768,N_19501,N_18908);
nor U21769 (N_21769,N_19199,N_19999);
nor U21770 (N_21770,N_18215,N_19834);
xor U21771 (N_21771,N_19939,N_18144);
xor U21772 (N_21772,N_19263,N_18957);
or U21773 (N_21773,N_19999,N_19687);
and U21774 (N_21774,N_18397,N_19727);
nor U21775 (N_21775,N_19205,N_18542);
xor U21776 (N_21776,N_19250,N_19192);
nor U21777 (N_21777,N_18983,N_18283);
nor U21778 (N_21778,N_19998,N_19629);
and U21779 (N_21779,N_19867,N_19943);
xnor U21780 (N_21780,N_18727,N_18892);
or U21781 (N_21781,N_18512,N_18052);
nor U21782 (N_21782,N_18609,N_18760);
xnor U21783 (N_21783,N_19289,N_19635);
or U21784 (N_21784,N_19036,N_19233);
nor U21785 (N_21785,N_18584,N_19192);
and U21786 (N_21786,N_18821,N_18895);
nand U21787 (N_21787,N_19500,N_19671);
xnor U21788 (N_21788,N_18402,N_19897);
nand U21789 (N_21789,N_19808,N_18366);
or U21790 (N_21790,N_18677,N_18755);
nand U21791 (N_21791,N_19037,N_18878);
or U21792 (N_21792,N_19842,N_19871);
xor U21793 (N_21793,N_18168,N_19299);
or U21794 (N_21794,N_19840,N_18907);
nor U21795 (N_21795,N_18903,N_18221);
xor U21796 (N_21796,N_18581,N_19507);
xnor U21797 (N_21797,N_18775,N_18298);
or U21798 (N_21798,N_19518,N_18400);
xnor U21799 (N_21799,N_18733,N_19605);
or U21800 (N_21800,N_19917,N_19760);
and U21801 (N_21801,N_18036,N_18346);
xor U21802 (N_21802,N_19712,N_19242);
nor U21803 (N_21803,N_19146,N_18062);
and U21804 (N_21804,N_19635,N_19584);
nor U21805 (N_21805,N_19870,N_18746);
nor U21806 (N_21806,N_19418,N_18987);
xnor U21807 (N_21807,N_18677,N_18276);
xnor U21808 (N_21808,N_19750,N_19727);
and U21809 (N_21809,N_18605,N_19010);
xnor U21810 (N_21810,N_19965,N_18237);
nor U21811 (N_21811,N_18007,N_19423);
and U21812 (N_21812,N_19485,N_18430);
or U21813 (N_21813,N_19960,N_19944);
nand U21814 (N_21814,N_19582,N_19334);
xnor U21815 (N_21815,N_18646,N_18655);
nor U21816 (N_21816,N_19588,N_19700);
and U21817 (N_21817,N_19167,N_18582);
xor U21818 (N_21818,N_19958,N_18802);
nand U21819 (N_21819,N_18120,N_19494);
nor U21820 (N_21820,N_18062,N_19486);
xnor U21821 (N_21821,N_19782,N_18893);
nand U21822 (N_21822,N_19515,N_18827);
nand U21823 (N_21823,N_18915,N_19019);
nor U21824 (N_21824,N_18184,N_19798);
xnor U21825 (N_21825,N_19138,N_19949);
or U21826 (N_21826,N_19991,N_19972);
nor U21827 (N_21827,N_18140,N_18541);
xnor U21828 (N_21828,N_18698,N_18478);
and U21829 (N_21829,N_18366,N_19870);
xnor U21830 (N_21830,N_18204,N_18398);
or U21831 (N_21831,N_19674,N_19190);
and U21832 (N_21832,N_19197,N_18934);
or U21833 (N_21833,N_18045,N_18525);
and U21834 (N_21834,N_19354,N_19180);
nor U21835 (N_21835,N_19643,N_19710);
or U21836 (N_21836,N_18612,N_18344);
and U21837 (N_21837,N_18629,N_19667);
and U21838 (N_21838,N_18101,N_19320);
nor U21839 (N_21839,N_19681,N_19647);
nor U21840 (N_21840,N_18329,N_19314);
xor U21841 (N_21841,N_19738,N_18301);
and U21842 (N_21842,N_19730,N_18490);
nor U21843 (N_21843,N_18141,N_19809);
nand U21844 (N_21844,N_19724,N_19478);
nor U21845 (N_21845,N_18104,N_19205);
nand U21846 (N_21846,N_18269,N_19393);
nor U21847 (N_21847,N_19420,N_19751);
or U21848 (N_21848,N_18417,N_18835);
or U21849 (N_21849,N_18443,N_19381);
or U21850 (N_21850,N_19696,N_18148);
nor U21851 (N_21851,N_19377,N_19837);
nor U21852 (N_21852,N_19083,N_18359);
and U21853 (N_21853,N_19911,N_19811);
xnor U21854 (N_21854,N_18060,N_18085);
nor U21855 (N_21855,N_19257,N_19724);
nand U21856 (N_21856,N_19914,N_19777);
and U21857 (N_21857,N_19276,N_19615);
nand U21858 (N_21858,N_19769,N_19628);
xnor U21859 (N_21859,N_18982,N_19064);
or U21860 (N_21860,N_19966,N_19048);
or U21861 (N_21861,N_18822,N_19024);
or U21862 (N_21862,N_18689,N_19374);
xnor U21863 (N_21863,N_18227,N_18188);
xnor U21864 (N_21864,N_18518,N_18459);
and U21865 (N_21865,N_18471,N_19339);
and U21866 (N_21866,N_18655,N_19020);
or U21867 (N_21867,N_18862,N_19568);
nand U21868 (N_21868,N_19637,N_18808);
nor U21869 (N_21869,N_19236,N_18081);
nand U21870 (N_21870,N_18089,N_19919);
or U21871 (N_21871,N_18291,N_19111);
or U21872 (N_21872,N_18653,N_19287);
nor U21873 (N_21873,N_19233,N_18815);
xnor U21874 (N_21874,N_19446,N_19394);
or U21875 (N_21875,N_19631,N_19782);
and U21876 (N_21876,N_19288,N_19088);
nor U21877 (N_21877,N_19164,N_19227);
nor U21878 (N_21878,N_19062,N_18586);
or U21879 (N_21879,N_19206,N_19300);
or U21880 (N_21880,N_19668,N_18717);
or U21881 (N_21881,N_19670,N_18891);
nor U21882 (N_21882,N_19677,N_18424);
and U21883 (N_21883,N_19529,N_18488);
nand U21884 (N_21884,N_18916,N_19999);
xor U21885 (N_21885,N_19126,N_18110);
xnor U21886 (N_21886,N_19422,N_19038);
nand U21887 (N_21887,N_19345,N_18521);
xnor U21888 (N_21888,N_18051,N_19534);
nor U21889 (N_21889,N_18467,N_19905);
nand U21890 (N_21890,N_19959,N_18121);
and U21891 (N_21891,N_18357,N_18948);
nand U21892 (N_21892,N_19527,N_19649);
nor U21893 (N_21893,N_18462,N_18691);
and U21894 (N_21894,N_19703,N_18624);
nand U21895 (N_21895,N_18750,N_18308);
nor U21896 (N_21896,N_19330,N_18353);
nor U21897 (N_21897,N_19860,N_18671);
nor U21898 (N_21898,N_19541,N_19961);
nor U21899 (N_21899,N_18567,N_18438);
or U21900 (N_21900,N_18603,N_18238);
or U21901 (N_21901,N_18381,N_18535);
nand U21902 (N_21902,N_18452,N_19937);
and U21903 (N_21903,N_19515,N_18073);
or U21904 (N_21904,N_19071,N_19365);
nand U21905 (N_21905,N_18110,N_18488);
xor U21906 (N_21906,N_18338,N_18241);
and U21907 (N_21907,N_19211,N_19734);
nor U21908 (N_21908,N_19078,N_18300);
and U21909 (N_21909,N_19173,N_18915);
and U21910 (N_21910,N_19121,N_19167);
or U21911 (N_21911,N_18049,N_19484);
nor U21912 (N_21912,N_18323,N_19655);
or U21913 (N_21913,N_19097,N_18516);
xor U21914 (N_21914,N_19696,N_19895);
or U21915 (N_21915,N_18249,N_18652);
xor U21916 (N_21916,N_19874,N_18526);
nand U21917 (N_21917,N_18406,N_18745);
or U21918 (N_21918,N_18354,N_19332);
nor U21919 (N_21919,N_19238,N_19642);
xor U21920 (N_21920,N_19355,N_19461);
nor U21921 (N_21921,N_18467,N_18698);
or U21922 (N_21922,N_18049,N_18200);
nor U21923 (N_21923,N_18598,N_18201);
or U21924 (N_21924,N_19604,N_19286);
and U21925 (N_21925,N_19570,N_19869);
or U21926 (N_21926,N_18598,N_18590);
and U21927 (N_21927,N_18098,N_18685);
xor U21928 (N_21928,N_19626,N_18697);
and U21929 (N_21929,N_19622,N_18576);
and U21930 (N_21930,N_18830,N_19856);
nand U21931 (N_21931,N_18074,N_19355);
nor U21932 (N_21932,N_18356,N_18483);
nor U21933 (N_21933,N_18912,N_18130);
xnor U21934 (N_21934,N_18643,N_18188);
nor U21935 (N_21935,N_19009,N_19380);
nand U21936 (N_21936,N_19272,N_18355);
nor U21937 (N_21937,N_18108,N_18645);
and U21938 (N_21938,N_19085,N_19966);
xor U21939 (N_21939,N_19183,N_18853);
or U21940 (N_21940,N_18426,N_19641);
and U21941 (N_21941,N_19179,N_18522);
nand U21942 (N_21942,N_18614,N_18460);
nand U21943 (N_21943,N_18213,N_18345);
nand U21944 (N_21944,N_18045,N_19504);
and U21945 (N_21945,N_19250,N_18760);
nand U21946 (N_21946,N_18467,N_19206);
and U21947 (N_21947,N_18246,N_19037);
nor U21948 (N_21948,N_18911,N_19672);
and U21949 (N_21949,N_19167,N_18187);
and U21950 (N_21950,N_19390,N_19864);
and U21951 (N_21951,N_18002,N_19521);
nand U21952 (N_21952,N_18687,N_18709);
xor U21953 (N_21953,N_18068,N_18054);
nor U21954 (N_21954,N_19036,N_19901);
xor U21955 (N_21955,N_19813,N_19665);
nor U21956 (N_21956,N_19525,N_19242);
and U21957 (N_21957,N_18692,N_18757);
nand U21958 (N_21958,N_19122,N_18495);
and U21959 (N_21959,N_19398,N_18850);
nor U21960 (N_21960,N_18173,N_19226);
xnor U21961 (N_21961,N_19798,N_19976);
xnor U21962 (N_21962,N_19383,N_18902);
nand U21963 (N_21963,N_18787,N_18524);
xnor U21964 (N_21964,N_19260,N_18470);
or U21965 (N_21965,N_19139,N_18893);
nand U21966 (N_21966,N_18082,N_19919);
nor U21967 (N_21967,N_19032,N_18214);
nor U21968 (N_21968,N_18919,N_19205);
and U21969 (N_21969,N_18119,N_19133);
xnor U21970 (N_21970,N_18111,N_18917);
xor U21971 (N_21971,N_18442,N_19290);
nand U21972 (N_21972,N_19109,N_19973);
and U21973 (N_21973,N_18994,N_18469);
or U21974 (N_21974,N_18502,N_19745);
nand U21975 (N_21975,N_18633,N_18456);
nor U21976 (N_21976,N_18447,N_19527);
and U21977 (N_21977,N_19404,N_18390);
and U21978 (N_21978,N_18425,N_19791);
and U21979 (N_21979,N_19321,N_19618);
nor U21980 (N_21980,N_18786,N_18508);
xnor U21981 (N_21981,N_18235,N_18500);
xor U21982 (N_21982,N_19893,N_18963);
nor U21983 (N_21983,N_18721,N_19856);
nor U21984 (N_21984,N_18275,N_18492);
nand U21985 (N_21985,N_19199,N_18729);
xnor U21986 (N_21986,N_19071,N_19741);
or U21987 (N_21987,N_19527,N_18945);
and U21988 (N_21988,N_18764,N_19949);
and U21989 (N_21989,N_18994,N_18439);
nand U21990 (N_21990,N_19893,N_19378);
nand U21991 (N_21991,N_19402,N_18460);
and U21992 (N_21992,N_19242,N_18013);
or U21993 (N_21993,N_19101,N_18313);
and U21994 (N_21994,N_19427,N_19535);
xnor U21995 (N_21995,N_18792,N_19815);
and U21996 (N_21996,N_18996,N_19692);
nor U21997 (N_21997,N_19778,N_19392);
or U21998 (N_21998,N_18812,N_19243);
xnor U21999 (N_21999,N_18237,N_19275);
xor U22000 (N_22000,N_21914,N_21788);
nor U22001 (N_22001,N_21213,N_20829);
and U22002 (N_22002,N_20946,N_20218);
xor U22003 (N_22003,N_21892,N_21954);
and U22004 (N_22004,N_21774,N_21106);
nand U22005 (N_22005,N_20156,N_20446);
nand U22006 (N_22006,N_21725,N_21766);
or U22007 (N_22007,N_21399,N_20831);
nor U22008 (N_22008,N_21732,N_20095);
and U22009 (N_22009,N_21404,N_20406);
or U22010 (N_22010,N_21060,N_21228);
and U22011 (N_22011,N_20072,N_21207);
and U22012 (N_22012,N_20139,N_20165);
and U22013 (N_22013,N_21872,N_21628);
or U22014 (N_22014,N_21984,N_20726);
nand U22015 (N_22015,N_20339,N_20167);
or U22016 (N_22016,N_21898,N_21062);
nand U22017 (N_22017,N_21230,N_20252);
xnor U22018 (N_22018,N_21809,N_20659);
xnor U22019 (N_22019,N_20914,N_21359);
or U22020 (N_22020,N_21966,N_21490);
nand U22021 (N_22021,N_21688,N_20013);
nor U22022 (N_22022,N_20195,N_20382);
xor U22023 (N_22023,N_21524,N_20884);
nand U22024 (N_22024,N_20414,N_21654);
and U22025 (N_22025,N_20990,N_21812);
xnor U22026 (N_22026,N_21350,N_21697);
xnor U22027 (N_22027,N_21387,N_20492);
nor U22028 (N_22028,N_21367,N_21440);
xor U22029 (N_22029,N_21629,N_21990);
nor U22030 (N_22030,N_20038,N_21020);
nand U22031 (N_22031,N_20761,N_21454);
nor U22032 (N_22032,N_21423,N_21357);
or U22033 (N_22033,N_20225,N_21610);
or U22034 (N_22034,N_20904,N_21811);
or U22035 (N_22035,N_20314,N_21364);
nor U22036 (N_22036,N_21739,N_20424);
xnor U22037 (N_22037,N_20893,N_21283);
nor U22038 (N_22038,N_21846,N_20941);
nand U22039 (N_22039,N_20223,N_20454);
nor U22040 (N_22040,N_21791,N_20319);
nor U22041 (N_22041,N_20693,N_21355);
or U22042 (N_22042,N_20549,N_20898);
nor U22043 (N_22043,N_20330,N_21154);
and U22044 (N_22044,N_20459,N_20716);
xnor U22045 (N_22045,N_20355,N_21079);
nand U22046 (N_22046,N_20891,N_21082);
nand U22047 (N_22047,N_20912,N_20604);
nor U22048 (N_22048,N_20266,N_21940);
or U22049 (N_22049,N_20244,N_21613);
xor U22050 (N_22050,N_21602,N_21095);
nor U22051 (N_22051,N_21310,N_21088);
or U22052 (N_22052,N_20067,N_21836);
or U22053 (N_22053,N_21048,N_21176);
and U22054 (N_22054,N_21054,N_20079);
xnor U22055 (N_22055,N_20270,N_20516);
nand U22056 (N_22056,N_21152,N_20348);
nor U22057 (N_22057,N_21773,N_20438);
nor U22058 (N_22058,N_21273,N_20514);
or U22059 (N_22059,N_21127,N_21694);
or U22060 (N_22060,N_20626,N_20931);
xnor U22061 (N_22061,N_21757,N_21202);
nor U22062 (N_22062,N_21292,N_21280);
nand U22063 (N_22063,N_20572,N_21352);
xnor U22064 (N_22064,N_21869,N_20996);
and U22065 (N_22065,N_20276,N_21438);
and U22066 (N_22066,N_21566,N_20137);
and U22067 (N_22067,N_21470,N_21883);
xnor U22068 (N_22068,N_21320,N_20718);
nand U22069 (N_22069,N_20029,N_20034);
nand U22070 (N_22070,N_20151,N_20022);
and U22071 (N_22071,N_21923,N_20630);
and U22072 (N_22072,N_20674,N_20047);
or U22073 (N_22073,N_21449,N_20369);
nand U22074 (N_22074,N_21734,N_21445);
nand U22075 (N_22075,N_20159,N_21876);
nand U22076 (N_22076,N_20405,N_20080);
or U22077 (N_22077,N_20537,N_21264);
xor U22078 (N_22078,N_20986,N_20105);
xor U22079 (N_22079,N_20683,N_20526);
nand U22080 (N_22080,N_20471,N_21329);
nand U22081 (N_22081,N_21968,N_21815);
or U22082 (N_22082,N_20116,N_21887);
or U22083 (N_22083,N_21525,N_21414);
and U22084 (N_22084,N_20189,N_21483);
nand U22085 (N_22085,N_20363,N_21792);
nand U22086 (N_22086,N_20994,N_20593);
nor U22087 (N_22087,N_20863,N_21542);
and U22088 (N_22088,N_20240,N_21765);
or U22089 (N_22089,N_20714,N_21253);
nor U22090 (N_22090,N_21475,N_21021);
nor U22091 (N_22091,N_20612,N_21073);
nand U22092 (N_22092,N_21249,N_20852);
and U22093 (N_22093,N_20820,N_21850);
nand U22094 (N_22094,N_21004,N_20269);
nor U22095 (N_22095,N_21057,N_21056);
or U22096 (N_22096,N_20699,N_20963);
nor U22097 (N_22097,N_21536,N_20573);
xor U22098 (N_22098,N_20303,N_21282);
nor U22099 (N_22099,N_20608,N_20380);
and U22100 (N_22100,N_21903,N_21938);
nor U22101 (N_22101,N_21820,N_21879);
nor U22102 (N_22102,N_20848,N_20673);
nand U22103 (N_22103,N_20069,N_20379);
xor U22104 (N_22104,N_20345,N_21728);
and U22105 (N_22105,N_20190,N_20584);
and U22106 (N_22106,N_21810,N_20992);
nor U22107 (N_22107,N_20377,N_20478);
and U22108 (N_22108,N_20119,N_21341);
nor U22109 (N_22109,N_21917,N_21323);
or U22110 (N_22110,N_21169,N_21751);
or U22111 (N_22111,N_20425,N_21649);
nor U22112 (N_22112,N_21086,N_20388);
xor U22113 (N_22113,N_20408,N_20544);
or U22114 (N_22114,N_20474,N_21606);
or U22115 (N_22115,N_20551,N_21746);
nand U22116 (N_22116,N_20058,N_21698);
and U22117 (N_22117,N_21983,N_21556);
or U22118 (N_22118,N_21945,N_20725);
nand U22119 (N_22119,N_21240,N_20577);
or U22120 (N_22120,N_20463,N_21568);
xor U22121 (N_22121,N_20493,N_21199);
and U22122 (N_22122,N_20441,N_20274);
xor U22123 (N_22123,N_21922,N_20364);
nor U22124 (N_22124,N_20219,N_20410);
xor U22125 (N_22125,N_20136,N_20293);
nor U22126 (N_22126,N_21096,N_21242);
nand U22127 (N_22127,N_21370,N_20921);
and U22128 (N_22128,N_20158,N_20756);
xnor U22129 (N_22129,N_21593,N_21394);
xor U22130 (N_22130,N_21627,N_20563);
nand U22131 (N_22131,N_21172,N_21389);
nand U22132 (N_22132,N_20206,N_20403);
nand U22133 (N_22133,N_21999,N_21032);
nand U22134 (N_22134,N_21309,N_21306);
nand U22135 (N_22135,N_21499,N_20854);
or U22136 (N_22136,N_20899,N_20552);
nor U22137 (N_22137,N_21641,N_21011);
nor U22138 (N_22138,N_20569,N_21336);
xor U22139 (N_22139,N_21527,N_21117);
or U22140 (N_22140,N_21884,N_21797);
nor U22141 (N_22141,N_20669,N_21017);
or U22142 (N_22142,N_21582,N_20093);
nor U22143 (N_22143,N_20816,N_20130);
nor U22144 (N_22144,N_21078,N_20845);
or U22145 (N_22145,N_20827,N_20850);
nor U22146 (N_22146,N_21235,N_20596);
xnor U22147 (N_22147,N_20510,N_21795);
xor U22148 (N_22148,N_20332,N_20647);
or U22149 (N_22149,N_21551,N_20086);
nor U22150 (N_22150,N_21540,N_20582);
nor U22151 (N_22151,N_20028,N_21908);
xnor U22152 (N_22152,N_21175,N_21642);
xnor U22153 (N_22153,N_20114,N_21683);
xor U22154 (N_22154,N_21171,N_20987);
nor U22155 (N_22155,N_21581,N_21112);
or U22156 (N_22156,N_21772,N_21588);
nand U22157 (N_22157,N_21089,N_21248);
nand U22158 (N_22158,N_20457,N_21130);
xor U22159 (N_22159,N_21994,N_20228);
and U22160 (N_22160,N_20016,N_20295);
xnor U22161 (N_22161,N_21074,N_20880);
or U22162 (N_22162,N_20122,N_21347);
nand U22163 (N_22163,N_21959,N_20623);
nor U22164 (N_22164,N_20209,N_20800);
xor U22165 (N_22165,N_20634,N_20354);
xnor U22166 (N_22166,N_21436,N_20146);
and U22167 (N_22167,N_21519,N_20157);
nand U22168 (N_22168,N_20624,N_20595);
nor U22169 (N_22169,N_20064,N_20342);
and U22170 (N_22170,N_21194,N_20635);
nor U22171 (N_22171,N_20678,N_20692);
and U22172 (N_22172,N_21821,N_21245);
or U22173 (N_22173,N_21105,N_20654);
xnor U22174 (N_22174,N_20822,N_21114);
nand U22175 (N_22175,N_20886,N_21801);
and U22176 (N_22176,N_21302,N_20087);
nand U22177 (N_22177,N_21182,N_21743);
or U22178 (N_22178,N_21446,N_20541);
nor U22179 (N_22179,N_21433,N_21029);
and U22180 (N_22180,N_20025,N_20277);
and U22181 (N_22181,N_21794,N_20773);
or U22182 (N_22182,N_20389,N_21771);
xor U22183 (N_22183,N_21673,N_21687);
nand U22184 (N_22184,N_21702,N_20300);
and U22185 (N_22185,N_21951,N_21635);
nand U22186 (N_22186,N_21730,N_21873);
and U22187 (N_22187,N_21865,N_20422);
xor U22188 (N_22188,N_20394,N_21076);
and U22189 (N_22189,N_21948,N_20642);
and U22190 (N_22190,N_21197,N_20281);
nor U22191 (N_22191,N_20180,N_21374);
xor U22192 (N_22192,N_20603,N_20585);
nor U22193 (N_22193,N_20239,N_20063);
and U22194 (N_22194,N_20045,N_20134);
or U22195 (N_22195,N_21550,N_21521);
nor U22196 (N_22196,N_21888,N_20734);
and U22197 (N_22197,N_20755,N_21878);
xnor U22198 (N_22198,N_21224,N_21695);
and U22199 (N_22199,N_20702,N_21428);
xnor U22200 (N_22200,N_20580,N_21392);
or U22201 (N_22201,N_21612,N_21093);
nand U22202 (N_22202,N_20291,N_21344);
and U22203 (N_22203,N_21868,N_21885);
xnor U22204 (N_22204,N_20973,N_20217);
and U22205 (N_22205,N_21045,N_20766);
and U22206 (N_22206,N_20908,N_21987);
nand U22207 (N_22207,N_20535,N_21307);
nand U22208 (N_22208,N_20220,N_20231);
xor U22209 (N_22209,N_20943,N_20682);
or U22210 (N_22210,N_20280,N_21256);
xnor U22211 (N_22211,N_20201,N_21296);
or U22212 (N_22212,N_21901,N_20675);
and U22213 (N_22213,N_20708,N_20306);
or U22214 (N_22214,N_21488,N_21929);
and U22215 (N_22215,N_20507,N_21786);
nand U22216 (N_22216,N_21837,N_21961);
xnor U22217 (N_22217,N_21647,N_20315);
nor U22218 (N_22218,N_21462,N_20870);
nand U22219 (N_22219,N_20819,N_20125);
and U22220 (N_22220,N_21173,N_21972);
and U22221 (N_22221,N_20964,N_20103);
xnor U22222 (N_22222,N_21274,N_21150);
xnor U22223 (N_22223,N_21268,N_21996);
or U22224 (N_22224,N_20149,N_20468);
and U22225 (N_22225,N_20442,N_21388);
and U22226 (N_22226,N_21390,N_21395);
nand U22227 (N_22227,N_21431,N_20465);
xor U22228 (N_22228,N_20839,N_21376);
or U22229 (N_22229,N_21239,N_20002);
nand U22230 (N_22230,N_21149,N_21672);
nand U22231 (N_22231,N_20617,N_20041);
xor U22232 (N_22232,N_20937,N_21384);
or U22233 (N_22233,N_20476,N_21439);
nand U22234 (N_22234,N_20519,N_21886);
xor U22235 (N_22235,N_20836,N_21177);
nor U22236 (N_22236,N_21975,N_20932);
nor U22237 (N_22237,N_21978,N_21375);
and U22238 (N_22238,N_21121,N_21829);
nor U22239 (N_22239,N_21639,N_20609);
or U22240 (N_22240,N_20416,N_20186);
or U22241 (N_22241,N_20672,N_21552);
nand U22242 (N_22242,N_21759,N_21232);
xnor U22243 (N_22243,N_20719,N_20412);
nor U22244 (N_22244,N_21398,N_20030);
or U22245 (N_22245,N_20869,N_21301);
xnor U22246 (N_22246,N_20329,N_20411);
or U22247 (N_22247,N_20956,N_20031);
or U22248 (N_22248,N_21132,N_20823);
xor U22249 (N_22249,N_21825,N_21102);
nand U22250 (N_22250,N_20234,N_21158);
and U22251 (N_22251,N_21337,N_20288);
nor U22252 (N_22252,N_20779,N_21133);
nand U22253 (N_22253,N_20627,N_21616);
xnor U22254 (N_22254,N_20495,N_20444);
nand U22255 (N_22255,N_20920,N_21564);
nand U22256 (N_22256,N_20834,N_21382);
and U22257 (N_22257,N_21410,N_21690);
xnor U22258 (N_22258,N_20546,N_20343);
nor U22259 (N_22259,N_20333,N_21346);
or U22260 (N_22260,N_20715,N_20275);
nor U22261 (N_22261,N_21727,N_21510);
xnor U22262 (N_22262,N_20224,N_20916);
and U22263 (N_22263,N_20227,N_20088);
xor U22264 (N_22264,N_20575,N_20236);
xnor U22265 (N_22265,N_21035,N_20667);
xnor U22266 (N_22266,N_21981,N_21859);
and U22267 (N_22267,N_21162,N_21014);
nand U22268 (N_22268,N_20959,N_21682);
or U22269 (N_22269,N_20798,N_21135);
and U22270 (N_22270,N_21209,N_20808);
nor U22271 (N_22271,N_20538,N_21882);
and U22272 (N_22272,N_20062,N_21587);
and U22273 (N_22273,N_20824,N_21142);
xnor U22274 (N_22274,N_20074,N_20129);
nor U22275 (N_22275,N_20358,N_20974);
or U22276 (N_22276,N_21800,N_21024);
or U22277 (N_22277,N_20464,N_21650);
and U22278 (N_22278,N_20096,N_20110);
nor U22279 (N_22279,N_20109,N_20366);
nor U22280 (N_22280,N_20605,N_20525);
xnor U22281 (N_22281,N_21717,N_21247);
and U22282 (N_22282,N_21196,N_20501);
nand U22283 (N_22283,N_20795,N_20211);
nor U22284 (N_22284,N_20602,N_21779);
nor U22285 (N_22285,N_20371,N_20433);
or U22286 (N_22286,N_20940,N_21755);
nand U22287 (N_22287,N_20254,N_21049);
and U22288 (N_22288,N_20417,N_20243);
or U22289 (N_22289,N_21118,N_20090);
nor U22290 (N_22290,N_20668,N_21934);
and U22291 (N_22291,N_21441,N_20977);
xnor U22292 (N_22292,N_21385,N_20560);
or U22293 (N_22293,N_21509,N_20619);
xnor U22294 (N_22294,N_20326,N_21544);
and U22295 (N_22295,N_21862,N_21126);
xnor U22296 (N_22296,N_20196,N_21397);
xnor U22297 (N_22297,N_21339,N_20882);
and U22298 (N_22298,N_20607,N_20485);
or U22299 (N_22299,N_21071,N_21660);
nand U22300 (N_22300,N_21899,N_20426);
nand U22301 (N_22301,N_21806,N_20828);
nor U22302 (N_22302,N_21210,N_20771);
nand U22303 (N_22303,N_20531,N_21511);
xor U22304 (N_22304,N_21591,N_20840);
or U22305 (N_22305,N_21760,N_20737);
nor U22306 (N_22306,N_21457,N_21258);
or U22307 (N_22307,N_21895,N_20632);
and U22308 (N_22308,N_20311,N_21300);
xor U22309 (N_22309,N_21526,N_21512);
nor U22310 (N_22310,N_20688,N_21804);
xnor U22311 (N_22311,N_21645,N_20622);
and U22312 (N_22312,N_21281,N_20530);
and U22313 (N_22313,N_21492,N_21269);
or U22314 (N_22314,N_21030,N_21471);
xor U22315 (N_22315,N_20923,N_21824);
nor U22316 (N_22316,N_21299,N_21619);
or U22317 (N_22317,N_21770,N_20768);
nor U22318 (N_22318,N_20804,N_21776);
or U22319 (N_22319,N_20101,N_20078);
nand U22320 (N_22320,N_21195,N_20085);
xnor U22321 (N_22321,N_20500,N_21193);
and U22322 (N_22322,N_21855,N_20255);
or U22323 (N_22323,N_20184,N_20374);
nor U22324 (N_22324,N_21547,N_21167);
or U22325 (N_22325,N_21119,N_20427);
nor U22326 (N_22326,N_21379,N_21543);
xor U22327 (N_22327,N_20147,N_21603);
nand U22328 (N_22328,N_20684,N_20644);
or U22329 (N_22329,N_21001,N_20121);
nor U22330 (N_22330,N_21338,N_20302);
nor U22331 (N_22331,N_21580,N_20451);
nor U22332 (N_22332,N_21563,N_20133);
nand U22333 (N_22333,N_20356,N_20491);
nand U22334 (N_22334,N_20152,N_20955);
or U22335 (N_22335,N_21667,N_20076);
nor U22336 (N_22336,N_21129,N_20988);
and U22337 (N_22337,N_20655,N_21498);
nand U22338 (N_22338,N_20292,N_20806);
or U22339 (N_22339,N_20418,N_20154);
xnor U22340 (N_22340,N_20347,N_21317);
xnor U22341 (N_22341,N_20620,N_21799);
nand U22342 (N_22342,N_20318,N_21164);
nor U22343 (N_22343,N_21166,N_20599);
nor U22344 (N_22344,N_21992,N_20368);
or U22345 (N_22345,N_21244,N_21644);
and U22346 (N_22346,N_20749,N_20570);
xor U22347 (N_22347,N_21709,N_21830);
and U22348 (N_22348,N_21360,N_21085);
nor U22349 (N_22349,N_21700,N_21832);
nand U22350 (N_22350,N_21686,N_20375);
or U22351 (N_22351,N_20061,N_20046);
xor U22352 (N_22352,N_21617,N_20082);
nor U22353 (N_22353,N_20802,N_20203);
or U22354 (N_22354,N_20370,N_20140);
and U22355 (N_22355,N_20359,N_20504);
xor U22356 (N_22356,N_20173,N_20435);
nor U22357 (N_22357,N_21866,N_20975);
nor U22358 (N_22358,N_20689,N_21491);
xor U22359 (N_22359,N_20108,N_21960);
xnor U22360 (N_22360,N_21681,N_20037);
nand U22361 (N_22361,N_21289,N_21841);
nor U22362 (N_22362,N_20077,N_21002);
nand U22363 (N_22363,N_21015,N_20776);
nor U22364 (N_22364,N_20057,N_20349);
xor U22365 (N_22365,N_21116,N_21910);
nand U22366 (N_22366,N_21295,N_20968);
or U22367 (N_22367,N_20142,N_21377);
and U22368 (N_22368,N_21168,N_21493);
nor U22369 (N_22369,N_21924,N_20777);
and U22370 (N_22370,N_21936,N_20338);
nor U22371 (N_22371,N_20864,N_20871);
nor U22372 (N_22372,N_20202,N_20294);
xor U22373 (N_22373,N_21403,N_21600);
nor U22374 (N_22374,N_20498,N_21190);
and U22375 (N_22375,N_20008,N_20855);
nand U22376 (N_22376,N_21685,N_20600);
nand U22377 (N_22377,N_21615,N_20141);
nor U22378 (N_22378,N_21618,N_20767);
or U22379 (N_22379,N_20873,N_20743);
nor U22380 (N_22380,N_20232,N_21236);
nand U22381 (N_22381,N_21541,N_21270);
xnor U22382 (N_22382,N_21134,N_21051);
or U22383 (N_22383,N_21227,N_20543);
xnor U22384 (N_22384,N_21218,N_21170);
or U22385 (N_22385,N_21932,N_21065);
xor U22386 (N_22386,N_21533,N_21621);
xnor U22387 (N_22387,N_20738,N_20237);
and U22388 (N_22388,N_21037,N_20539);
or U22389 (N_22389,N_20948,N_21805);
and U22390 (N_22390,N_20327,N_21006);
nor U22391 (N_22391,N_21097,N_21448);
and U22392 (N_22392,N_21549,N_20488);
and U22393 (N_22393,N_21721,N_20534);
or U22394 (N_22394,N_21444,N_20246);
and U22395 (N_22395,N_20564,N_21894);
and U22396 (N_22396,N_20576,N_20759);
nand U22397 (N_22397,N_20128,N_20637);
or U22398 (N_22398,N_20872,N_20155);
or U22399 (N_22399,N_20657,N_20373);
nor U22400 (N_22400,N_20772,N_20790);
or U22401 (N_22401,N_21605,N_21442);
nand U22402 (N_22402,N_20594,N_20979);
xnor U22403 (N_22403,N_20399,N_20505);
nand U22404 (N_22404,N_21145,N_20296);
nand U22405 (N_22405,N_21070,N_21756);
nor U22406 (N_22406,N_21586,N_20331);
nand U22407 (N_22407,N_20470,N_20705);
nor U22408 (N_22408,N_20663,N_21677);
or U22409 (N_22409,N_21461,N_20258);
and U22410 (N_22410,N_20049,N_21816);
or U22411 (N_22411,N_21013,N_21583);
nor U22412 (N_22412,N_20976,N_20536);
xnor U22413 (N_22413,N_20409,N_21631);
xnor U22414 (N_22414,N_20443,N_21501);
and U22415 (N_22415,N_21189,N_20298);
and U22416 (N_22416,N_20351,N_20522);
or U22417 (N_22417,N_20520,N_20797);
xor U22418 (N_22418,N_21678,N_20928);
xor U22419 (N_22419,N_21955,N_20010);
nor U22420 (N_22420,N_21156,N_21557);
nand U22421 (N_22421,N_21704,N_20386);
and U22422 (N_22422,N_21502,N_21584);
xnor U22423 (N_22423,N_20739,N_20479);
nor U22424 (N_22424,N_20060,N_21326);
nor U22425 (N_22425,N_20229,N_21186);
nand U22426 (N_22426,N_21858,N_20307);
nor U22427 (N_22427,N_20467,N_20681);
and U22428 (N_22428,N_21560,N_21322);
nand U22429 (N_22429,N_21412,N_21098);
nor U22430 (N_22430,N_20111,N_20691);
nand U22431 (N_22431,N_21819,N_20264);
and U22432 (N_22432,N_21680,N_21092);
nand U22433 (N_22433,N_21831,N_21607);
and U22434 (N_22434,N_20018,N_20204);
and U22435 (N_22435,N_20760,N_21402);
nor U22436 (N_22436,N_20991,N_20769);
nor U22437 (N_22437,N_20949,N_21712);
xor U22438 (N_22438,N_20877,N_21211);
nor U22439 (N_22439,N_20353,N_21276);
or U22440 (N_22440,N_21084,N_21997);
and U22441 (N_22441,N_20023,N_21798);
and U22442 (N_22442,N_20117,N_20182);
or U22443 (N_22443,N_20911,N_21731);
xnor U22444 (N_22444,N_21405,N_20075);
nand U22445 (N_22445,N_20509,N_20094);
or U22446 (N_22446,N_20423,N_21467);
xor U22447 (N_22447,N_21450,N_21055);
and U22448 (N_22448,N_20287,N_21979);
nor U22449 (N_22449,N_21043,N_21646);
nor U22450 (N_22450,N_21316,N_20528);
xnor U22451 (N_22451,N_21919,N_20215);
and U22452 (N_22452,N_21304,N_21733);
nor U22453 (N_22453,N_21290,N_20826);
or U22454 (N_22454,N_21381,N_21918);
nand U22455 (N_22455,N_21161,N_21827);
and U22456 (N_22456,N_20717,N_21718);
nor U22457 (N_22457,N_21844,N_21622);
nand U22458 (N_22458,N_21109,N_21785);
nand U22459 (N_22459,N_20024,N_20462);
and U22460 (N_22460,N_20241,N_20562);
and U22461 (N_22461,N_21555,N_20508);
nand U22462 (N_22462,N_21763,N_21040);
and U22463 (N_22463,N_21003,N_21864);
or U22464 (N_22464,N_21986,N_20621);
or U22465 (N_22465,N_20671,N_20733);
nand U22466 (N_22466,N_20633,N_21921);
and U22467 (N_22467,N_21496,N_20936);
nand U22468 (N_22468,N_21148,N_21393);
nor U22469 (N_22469,N_21604,N_20922);
and U22470 (N_22470,N_20835,N_20091);
xnor U22471 (N_22471,N_20969,N_21880);
xor U22472 (N_22472,N_20550,N_21875);
and U22473 (N_22473,N_20200,N_21452);
nor U22474 (N_22474,N_20867,N_21203);
xnor U22475 (N_22475,N_21138,N_21008);
and U22476 (N_22476,N_20518,N_20833);
xnor U22477 (N_22477,N_21294,N_21447);
xnor U22478 (N_22478,N_21995,N_20282);
and U22479 (N_22479,N_21982,N_20497);
and U22480 (N_22480,N_20445,N_20053);
nor U22481 (N_22481,N_20253,N_21570);
and U22482 (N_22482,N_20178,N_21750);
nand U22483 (N_22483,N_20448,N_21146);
nand U22484 (N_22484,N_21719,N_21480);
and U22485 (N_22485,N_20006,N_20185);
nand U22486 (N_22486,N_21927,N_21851);
xnor U22487 (N_22487,N_21204,N_20557);
and U22488 (N_22488,N_21976,N_21005);
nand U22489 (N_22489,N_21159,N_20065);
xnor U22490 (N_22490,N_20611,N_20665);
nor U22491 (N_22491,N_21261,N_21857);
xor U22492 (N_22492,N_20192,N_20815);
or U22493 (N_22493,N_20701,N_20838);
nor U22494 (N_22494,N_20392,N_21184);
and U22495 (N_22495,N_21479,N_20837);
and U22496 (N_22496,N_20706,N_20529);
and U22497 (N_22497,N_21548,N_20106);
nor U22498 (N_22498,N_21971,N_20589);
or U22499 (N_22499,N_21692,N_20661);
or U22500 (N_22500,N_21928,N_21747);
or U22501 (N_22501,N_21468,N_20213);
or U22502 (N_22502,N_21522,N_21285);
nand U22503 (N_22503,N_21000,N_20793);
nor U22504 (N_22504,N_21577,N_21726);
nand U22505 (N_22505,N_21942,N_21155);
nand U22506 (N_22506,N_21072,N_20083);
nor U22507 (N_22507,N_21699,N_21340);
nand U22508 (N_22508,N_20758,N_20321);
and U22509 (N_22509,N_20316,N_21707);
xor U22510 (N_22510,N_21063,N_20614);
nand U22511 (N_22511,N_21590,N_21180);
nand U22512 (N_22512,N_21748,N_20279);
nand U22513 (N_22513,N_21291,N_21889);
or U22514 (N_22514,N_21980,N_21187);
and U22515 (N_22515,N_20805,N_21965);
or U22516 (N_22516,N_20162,N_20393);
or U22517 (N_22517,N_20641,N_21905);
nand U22518 (N_22518,N_20842,N_20014);
nor U22519 (N_22519,N_21991,N_20000);
nor U22520 (N_22520,N_20846,N_20262);
and U22521 (N_22521,N_20104,N_21250);
and U22522 (N_22522,N_21234,N_21046);
xnor U22523 (N_22523,N_21312,N_20044);
xnor U22524 (N_22524,N_21853,N_20565);
xor U22525 (N_22525,N_21506,N_20198);
and U22526 (N_22526,N_20272,N_21251);
and U22527 (N_22527,N_21443,N_20894);
xnor U22528 (N_22528,N_20325,N_20578);
or U22529 (N_22529,N_20547,N_21736);
and U22530 (N_22530,N_21693,N_21233);
and U22531 (N_22531,N_20748,N_21332);
or U22532 (N_22532,N_21953,N_20750);
or U22533 (N_22533,N_21315,N_21950);
nor U22534 (N_22534,N_20164,N_21663);
or U22535 (N_22535,N_20283,N_21874);
nor U22536 (N_22536,N_20753,N_20944);
and U22537 (N_22537,N_21424,N_21147);
nor U22538 (N_22538,N_20289,N_21077);
xor U22539 (N_22539,N_21313,N_20939);
nor U22540 (N_22540,N_21679,N_21599);
and U22541 (N_22541,N_21219,N_20460);
and U22542 (N_22542,N_21662,N_21396);
nand U22543 (N_22543,N_20700,N_20887);
or U22544 (N_22544,N_20161,N_21237);
nor U22545 (N_22545,N_20962,N_21897);
or U22546 (N_22546,N_20814,N_21188);
xor U22547 (N_22547,N_20740,N_20765);
nand U22548 (N_22548,N_20419,N_20794);
xnor U22549 (N_22549,N_21426,N_20452);
nand U22550 (N_22550,N_21254,N_21091);
and U22551 (N_22551,N_21260,N_20711);
or U22552 (N_22552,N_20197,N_20247);
nor U22553 (N_22553,N_20222,N_20420);
xnor U22554 (N_22554,N_20636,N_21411);
nor U22555 (N_22555,N_21041,N_21069);
or U22556 (N_22556,N_20163,N_21796);
nor U22557 (N_22557,N_21939,N_21066);
and U22558 (N_22558,N_21266,N_20927);
nand U22559 (N_22559,N_21453,N_20896);
and U22560 (N_22560,N_21460,N_20381);
nand U22561 (N_22561,N_21318,N_20774);
or U22562 (N_22562,N_21900,N_20561);
nand U22563 (N_22563,N_20746,N_20456);
nand U22564 (N_22564,N_21103,N_21674);
nor U22565 (N_22565,N_21417,N_21181);
xnor U22566 (N_22566,N_21368,N_21834);
nor U22567 (N_22567,N_21358,N_20817);
or U22568 (N_22568,N_20391,N_21275);
or U22569 (N_22569,N_21361,N_20704);
or U22570 (N_22570,N_20172,N_20984);
or U22571 (N_22571,N_21476,N_21231);
nand U22572 (N_22572,N_21803,N_21706);
and U22573 (N_22573,N_20512,N_20436);
xnor U22574 (N_22574,N_21226,N_20039);
nand U22575 (N_22575,N_20747,N_21061);
and U22576 (N_22576,N_21559,N_21861);
xor U22577 (N_22577,N_20763,N_20616);
and U22578 (N_22578,N_20881,N_21463);
nand U22579 (N_22579,N_21495,N_21775);
xor U22580 (N_22580,N_21022,N_20910);
nor U22581 (N_22581,N_20174,N_21601);
or U22582 (N_22582,N_20160,N_20764);
and U22583 (N_22583,N_20950,N_21331);
xor U22584 (N_22584,N_21125,N_20935);
and U22585 (N_22585,N_21516,N_21740);
xnor U22586 (N_22586,N_21518,N_21200);
nor U22587 (N_22587,N_21783,N_20066);
or U22588 (N_22588,N_20825,N_21474);
or U22589 (N_22589,N_20021,N_20450);
nand U22590 (N_22590,N_21425,N_21503);
xor U22591 (N_22591,N_21705,N_20148);
xnor U22592 (N_22592,N_20102,N_21325);
nor U22593 (N_22593,N_20513,N_20533);
nand U22594 (N_22594,N_21848,N_21205);
nor U22595 (N_22595,N_20628,N_21287);
and U22596 (N_22596,N_21241,N_20432);
or U22597 (N_22597,N_21691,N_20012);
nand U22598 (N_22598,N_20567,N_20489);
and U22599 (N_22599,N_21531,N_20906);
or U22600 (N_22600,N_20005,N_21123);
nand U22601 (N_22601,N_20801,N_20199);
xnor U22602 (N_22602,N_20284,N_21711);
nand U22603 (N_22603,N_21298,N_21342);
and U22604 (N_22604,N_21163,N_20131);
nand U22605 (N_22605,N_21016,N_21330);
nand U22606 (N_22606,N_20713,N_21598);
nor U22607 (N_22607,N_21572,N_20056);
xor U22608 (N_22608,N_21863,N_21949);
xnor U22609 (N_22609,N_21028,N_21137);
xor U22610 (N_22610,N_20727,N_21891);
or U22611 (N_22611,N_21335,N_21703);
or U22612 (N_22612,N_20340,N_20068);
xor U22613 (N_22613,N_21912,N_20484);
nand U22614 (N_22614,N_20050,N_20934);
or U22615 (N_22615,N_20554,N_21505);
xor U22616 (N_22616,N_20499,N_20810);
xor U22617 (N_22617,N_21140,N_20179);
or U22618 (N_22618,N_20144,N_21099);
nand U22619 (N_22619,N_21648,N_21482);
or U22620 (N_22620,N_21212,N_20588);
or U22621 (N_22621,N_21623,N_20360);
and U22622 (N_22622,N_21653,N_21589);
nor U22623 (N_22623,N_21321,N_21636);
xnor U22624 (N_22624,N_21802,N_20466);
and U22625 (N_22625,N_21174,N_21579);
nor U22626 (N_22626,N_20305,N_20558);
or U22627 (N_22627,N_20812,N_20397);
nor U22628 (N_22628,N_21787,N_20271);
or U22629 (N_22629,N_20791,N_20781);
and U22630 (N_22630,N_21539,N_20752);
or U22631 (N_22631,N_20517,N_20177);
or U22632 (N_22632,N_21745,N_20902);
xnor U22633 (N_22633,N_21489,N_21935);
xor U22634 (N_22634,N_21969,N_20084);
nand U22635 (N_22635,N_20789,N_20803);
or U22636 (N_22636,N_20242,N_21420);
nand U22637 (N_22637,N_20048,N_21345);
xnor U22638 (N_22638,N_20483,N_21023);
and U22639 (N_22639,N_21970,N_20187);
and U22640 (N_22640,N_21937,N_21749);
nand U22641 (N_22641,N_21497,N_20511);
and U22642 (N_22642,N_20590,N_21611);
xor U22643 (N_22643,N_20496,N_20112);
nand U22644 (N_22644,N_20267,N_20571);
and U22645 (N_22645,N_20322,N_21297);
xnor U22646 (N_22646,N_20653,N_20965);
xnor U22647 (N_22647,N_20751,N_21136);
xor U22648 (N_22648,N_21532,N_20120);
nand U22649 (N_22649,N_21666,N_21027);
and U22650 (N_22650,N_20744,N_21896);
xnor U22651 (N_22651,N_20469,N_20775);
and U22652 (N_22652,N_20615,N_20449);
nor U22653 (N_22653,N_21988,N_21523);
and U22654 (N_22654,N_21952,N_21380);
xnor U22655 (N_22655,N_20851,N_21752);
or U22656 (N_22656,N_20601,N_20866);
nand U22657 (N_22657,N_20532,N_21179);
and U22658 (N_22658,N_21416,N_20942);
or U22659 (N_22659,N_20957,N_20953);
or U22660 (N_22660,N_21514,N_21303);
and U22661 (N_22661,N_21789,N_20930);
nand U22662 (N_22662,N_20967,N_20004);
or U22663 (N_22663,N_20251,N_21573);
nor U22664 (N_22664,N_20960,N_20901);
xnor U22665 (N_22665,N_21090,N_21128);
xor U22666 (N_22666,N_21019,N_21664);
xor U22667 (N_22667,N_21034,N_21998);
nor U22668 (N_22668,N_21139,N_20506);
nand U22669 (N_22669,N_21255,N_21553);
xor U22670 (N_22670,N_20788,N_20915);
nand U22671 (N_22671,N_21363,N_21535);
nor U22672 (N_22672,N_20998,N_20650);
or U22673 (N_22673,N_21192,N_21401);
nor U22674 (N_22674,N_21545,N_21738);
xnor U22675 (N_22675,N_21277,N_20268);
or U22676 (N_22676,N_20703,N_20365);
nand U22677 (N_22677,N_21782,N_20579);
xnor U22678 (N_22678,N_21504,N_20334);
nand U22679 (N_22679,N_20115,N_20925);
and U22680 (N_22680,N_20421,N_20401);
and U22681 (N_22681,N_20900,N_20856);
nor U22682 (N_22682,N_20811,N_20261);
nor U22683 (N_22683,N_20376,N_20188);
nand U22684 (N_22684,N_21430,N_20431);
xor U22685 (N_22685,N_20807,N_21656);
nor U22686 (N_22686,N_20598,N_21638);
nand U22687 (N_22687,N_20384,N_20690);
or U22688 (N_22688,N_21407,N_21319);
or U22689 (N_22689,N_20337,N_20638);
nand U22690 (N_22690,N_20933,N_21151);
and U22691 (N_22691,N_21676,N_21478);
xor U22692 (N_22692,N_21620,N_21406);
nor U22693 (N_22693,N_21769,N_20892);
nor U22694 (N_22694,N_21354,N_21817);
and U22695 (N_22695,N_21630,N_20481);
or U22696 (N_22696,N_21201,N_21144);
xnor U22697 (N_22697,N_20707,N_21714);
nor U22698 (N_22698,N_20821,N_20770);
nor U22699 (N_22699,N_21500,N_20472);
or U22700 (N_22700,N_20841,N_20556);
or U22701 (N_22701,N_21068,N_20430);
nand U22702 (N_22702,N_20785,N_20553);
or U22703 (N_22703,N_21279,N_20145);
xnor U22704 (N_22704,N_20447,N_20978);
or U22705 (N_22705,N_21183,N_20631);
and U22706 (N_22706,N_20997,N_21508);
and U22707 (N_22707,N_21141,N_21465);
and U22708 (N_22708,N_21608,N_20404);
xor U22709 (N_22709,N_21413,N_20092);
and U22710 (N_22710,N_20778,N_20907);
xnor U22711 (N_22711,N_20081,N_21768);
nand U22712 (N_22712,N_21574,N_20043);
nor U22713 (N_22713,N_21349,N_21223);
xor U22714 (N_22714,N_21562,N_21486);
nor U22715 (N_22715,N_21124,N_21418);
nor U22716 (N_22716,N_20722,N_20032);
xnor U22717 (N_22717,N_21634,N_21909);
nor U22718 (N_22718,N_21758,N_20680);
nor U22719 (N_22719,N_20143,N_20361);
xnor U22720 (N_22720,N_21941,N_21484);
and U22721 (N_22721,N_20890,N_20677);
nand U22722 (N_22722,N_20487,N_21708);
xnor U22723 (N_22723,N_21534,N_20073);
nand U22724 (N_22724,N_21225,N_21569);
xor U22725 (N_22725,N_20336,N_21284);
or U22726 (N_22726,N_20954,N_21458);
nand U22727 (N_22727,N_20521,N_20226);
nor U22728 (N_22728,N_20309,N_20383);
and U22729 (N_22729,N_20730,N_20832);
or U22730 (N_22730,N_20679,N_20720);
xor U22731 (N_22731,N_20033,N_21947);
nor U22732 (N_22732,N_21429,N_21286);
nor U22733 (N_22733,N_20895,N_21383);
xor U22734 (N_22734,N_21867,N_21823);
nor U22735 (N_22735,N_20040,N_20876);
xor U22736 (N_22736,N_21537,N_20897);
xor U22737 (N_22737,N_20017,N_21920);
and U22738 (N_22738,N_20966,N_20741);
xnor U22739 (N_22739,N_20971,N_20862);
xor U22740 (N_22740,N_20475,N_21710);
or U22741 (N_22741,N_21643,N_20958);
nand U22742 (N_22742,N_20263,N_21050);
xor U22743 (N_22743,N_20256,N_21930);
xor U22744 (N_22744,N_21933,N_21437);
xnor U22745 (N_22745,N_21828,N_20429);
nand U22746 (N_22746,N_20745,N_20879);
nand U22747 (N_22747,N_20214,N_20754);
nand U22748 (N_22748,N_21856,N_20670);
xnor U22749 (N_22749,N_20118,N_20323);
nand U22750 (N_22750,N_20918,N_21852);
nor U22751 (N_22751,N_20656,N_21668);
nand U22752 (N_22752,N_21064,N_21288);
nor U22753 (N_22753,N_20883,N_20865);
nand U22754 (N_22754,N_21472,N_21915);
xor U22755 (N_22755,N_20909,N_21366);
and U22756 (N_22756,N_21716,N_20150);
and U22757 (N_22757,N_21962,N_20903);
or U22758 (N_22758,N_20183,N_20527);
or U22759 (N_22759,N_20818,N_20437);
nor U22760 (N_22760,N_21943,N_20868);
or U22761 (N_22761,N_20113,N_21944);
nor U22762 (N_22762,N_20171,N_21305);
xor U22763 (N_22763,N_21902,N_21115);
xor U22764 (N_22764,N_20297,N_20352);
xor U22765 (N_22765,N_20191,N_21963);
and U22766 (N_22766,N_20285,N_20055);
nor U22767 (N_22767,N_20993,N_20961);
and U22768 (N_22768,N_21308,N_21715);
and U22769 (N_22769,N_20099,N_20574);
nand U22770 (N_22770,N_20260,N_20153);
and U22771 (N_22771,N_21101,N_21671);
nand U22772 (N_22772,N_20221,N_20310);
nor U22773 (N_22773,N_21314,N_21080);
xor U22774 (N_22774,N_20015,N_21596);
xnor U22775 (N_22775,N_20736,N_20861);
nand U22776 (N_22776,N_21485,N_21293);
and U22777 (N_22777,N_20581,N_21371);
or U22778 (N_22778,N_21849,N_20723);
or U22779 (N_22779,N_21958,N_20857);
or U22780 (N_22780,N_20782,N_21780);
xor U22781 (N_22781,N_21753,N_20919);
nand U22782 (N_22782,N_21964,N_20132);
and U22783 (N_22783,N_21530,N_21538);
xnor U22784 (N_22784,N_21911,N_20696);
and U22785 (N_22785,N_21400,N_20729);
nor U22786 (N_22786,N_21893,N_20830);
nand U22787 (N_22787,N_20809,N_20341);
nand U22788 (N_22788,N_21778,N_20799);
or U22789 (N_22789,N_20646,N_20036);
nor U22790 (N_22790,N_21658,N_21839);
and U22791 (N_22791,N_21609,N_20721);
or U22792 (N_22792,N_20238,N_21735);
xor U22793 (N_22793,N_21432,N_20455);
xnor U22794 (N_22794,N_21520,N_20728);
nand U22795 (N_22795,N_21571,N_21640);
xnor U22796 (N_22796,N_20458,N_21575);
xnor U22797 (N_22797,N_20346,N_20257);
and U22798 (N_22798,N_21576,N_20888);
nor U22799 (N_22799,N_21554,N_20413);
nand U22800 (N_22800,N_20235,N_21257);
nor U22801 (N_22801,N_20929,N_20652);
nand U22802 (N_22802,N_21165,N_20362);
xor U22803 (N_22803,N_21956,N_20344);
nor U22804 (N_22804,N_21369,N_21221);
xor U22805 (N_22805,N_21661,N_21813);
nand U22806 (N_22806,N_20027,N_20999);
nand U22807 (N_22807,N_21026,N_20651);
nand U22808 (N_22808,N_21561,N_21160);
nand U22809 (N_22809,N_20985,N_20126);
nand U22810 (N_22810,N_20473,N_21110);
or U22811 (N_22811,N_20415,N_21348);
nand U22812 (N_22812,N_20540,N_20724);
nand U22813 (N_22813,N_21847,N_21100);
xor U22814 (N_22814,N_20193,N_20592);
nand U22815 (N_22815,N_20694,N_20490);
nand U22816 (N_22816,N_21333,N_20265);
xor U22817 (N_22817,N_21263,N_20878);
xor U22818 (N_22818,N_21993,N_21067);
nand U22819 (N_22819,N_21036,N_20390);
or U22820 (N_22820,N_20951,N_20009);
and U22821 (N_22821,N_21655,N_21267);
and U22822 (N_22822,N_21047,N_21826);
xnor U22823 (N_22823,N_20524,N_21094);
nor U22824 (N_22824,N_20098,N_20606);
nand U22825 (N_22825,N_20273,N_20402);
nand U22826 (N_22826,N_21652,N_20905);
or U22827 (N_22827,N_21632,N_20566);
xnor U22828 (N_22828,N_21422,N_20972);
nor U22829 (N_22829,N_20026,N_20385);
nor U22830 (N_22830,N_21926,N_20757);
nor U22831 (N_22831,N_21459,N_21989);
or U22832 (N_22832,N_21075,N_20230);
nor U22833 (N_22833,N_20613,N_21860);
or U22834 (N_22834,N_21957,N_20135);
xor U22835 (N_22835,N_20278,N_20732);
nor U22836 (N_22836,N_20643,N_21214);
xor U22837 (N_22837,N_20625,N_20780);
xnor U22838 (N_22838,N_21808,N_21271);
xor U22839 (N_22839,N_21637,N_21754);
xnor U22840 (N_22840,N_21845,N_20216);
and U22841 (N_22841,N_20917,N_20166);
and U22842 (N_22842,N_21372,N_21614);
or U22843 (N_22843,N_20054,N_21871);
xnor U22844 (N_22844,N_21010,N_20477);
nor U22845 (N_22845,N_21793,N_20658);
nor U22846 (N_22846,N_21624,N_21122);
nor U22847 (N_22847,N_20207,N_20317);
nor U22848 (N_22848,N_21822,N_20583);
nor U22849 (N_22849,N_20786,N_20889);
xor U22850 (N_22850,N_21818,N_20210);
or U22851 (N_22851,N_20194,N_20645);
or U22852 (N_22852,N_20301,N_20762);
xnor U22853 (N_22853,N_20697,N_21435);
xnor U22854 (N_22854,N_20502,N_20400);
nand U22855 (N_22855,N_20792,N_21513);
xnor U22856 (N_22856,N_21767,N_21907);
or U22857 (N_22857,N_21386,N_21042);
nand U22858 (N_22858,N_21104,N_20568);
xor U22859 (N_22859,N_20989,N_21713);
xnor U22860 (N_22860,N_20123,N_21843);
nand U22861 (N_22861,N_20324,N_20205);
nor U22862 (N_22862,N_21120,N_20019);
xnor U22863 (N_22863,N_20970,N_21216);
and U22864 (N_22864,N_20664,N_21262);
and U22865 (N_22865,N_21675,N_20859);
nor U22866 (N_22866,N_21724,N_21881);
or U22867 (N_22867,N_21565,N_21585);
xnor U22868 (N_22868,N_20731,N_21625);
and U22869 (N_22869,N_20523,N_21744);
and U22870 (N_22870,N_21456,N_20480);
nand U22871 (N_22871,N_21058,N_21722);
nand U22872 (N_22872,N_20350,N_20169);
and U22873 (N_22873,N_21870,N_21351);
or U22874 (N_22874,N_21311,N_21487);
and U22875 (N_22875,N_21729,N_21208);
nor U22876 (N_22876,N_21265,N_21973);
and U22877 (N_22877,N_21157,N_20698);
nand U22878 (N_22878,N_21324,N_20308);
nor U22879 (N_22879,N_21737,N_21784);
xnor U22880 (N_22880,N_20945,N_20853);
nand U22881 (N_22881,N_20742,N_20249);
and U22882 (N_22882,N_20245,N_21651);
or U22883 (N_22883,N_21373,N_21761);
and U22884 (N_22884,N_20618,N_21353);
and U22885 (N_22885,N_21854,N_21455);
and U22886 (N_22886,N_21529,N_20629);
nor U22887 (N_22887,N_21595,N_21153);
nand U22888 (N_22888,N_21108,N_21764);
and U22889 (N_22889,N_20127,N_21594);
nor U22890 (N_22890,N_20494,N_20461);
nand U22891 (N_22891,N_21217,N_21113);
nand U22892 (N_22892,N_20559,N_21025);
and U22893 (N_22893,N_21466,N_20597);
nand U22894 (N_22894,N_21083,N_21762);
nand U22895 (N_22895,N_20847,N_21415);
or U22896 (N_22896,N_20843,N_21835);
nand U22897 (N_22897,N_21272,N_20304);
xor U22898 (N_22898,N_21720,N_20335);
nor U22899 (N_22899,N_20849,N_20482);
xnor U22900 (N_22900,N_21362,N_21039);
nor U22901 (N_22901,N_20662,N_20059);
and U22902 (N_22902,N_21222,N_20070);
xor U22903 (N_22903,N_21777,N_21833);
nand U22904 (N_22904,N_20784,N_20947);
nand U22905 (N_22905,N_21178,N_20398);
nor U22906 (N_22906,N_20983,N_20170);
and U22907 (N_22907,N_20097,N_20610);
and U22908 (N_22908,N_21578,N_21464);
nor U22909 (N_22909,N_21742,N_20649);
and U22910 (N_22910,N_21328,N_21925);
and U22911 (N_22911,N_21626,N_21419);
xnor U22912 (N_22912,N_21528,N_20434);
nor U22913 (N_22913,N_20591,N_21906);
xnor U22914 (N_22914,N_20813,N_20003);
nor U22915 (N_22915,N_21477,N_20874);
or U22916 (N_22916,N_21111,N_20052);
or U22917 (N_22917,N_20648,N_21877);
xor U22918 (N_22918,N_20844,N_21409);
and U22919 (N_22919,N_20176,N_21840);
and U22920 (N_22920,N_21916,N_20396);
nand U22921 (N_22921,N_21259,N_21334);
xor U22922 (N_22922,N_21044,N_20407);
and U22923 (N_22923,N_20885,N_20555);
nor U22924 (N_22924,N_21967,N_20695);
nor U22925 (N_22925,N_20542,N_20687);
xnor U22926 (N_22926,N_20952,N_20320);
nand U22927 (N_22927,N_21107,N_21191);
xnor U22928 (N_22928,N_20328,N_20440);
and U22929 (N_22929,N_21081,N_20913);
and U22930 (N_22930,N_21974,N_21665);
nand U22931 (N_22931,N_20011,N_21904);
and U22932 (N_22932,N_21546,N_21633);
nor U22933 (N_22933,N_21059,N_21931);
xnor U22934 (N_22934,N_20486,N_20587);
nor U22935 (N_22935,N_21246,N_21427);
xnor U22936 (N_22936,N_20938,N_21592);
nor U22937 (N_22937,N_21515,N_20312);
or U22938 (N_22938,N_20735,N_20001);
xnor U22939 (N_22939,N_21494,N_21597);
and U22940 (N_22940,N_21238,N_20858);
xnor U22941 (N_22941,N_20100,N_21684);
nor U22942 (N_22942,N_20685,N_21220);
and U22943 (N_22943,N_20783,N_21481);
nor U22944 (N_22944,N_20453,N_21033);
nand U22945 (N_22945,N_21517,N_20372);
xor U22946 (N_22946,N_21378,N_21807);
nand U22947 (N_22947,N_21659,N_20138);
nand U22948 (N_22948,N_21558,N_20875);
nand U22949 (N_22949,N_21657,N_20515);
xor U22950 (N_22950,N_21408,N_20250);
nor U22951 (N_22951,N_20089,N_20395);
nor U22952 (N_22952,N_21507,N_21670);
nor U22953 (N_22953,N_20586,N_21278);
or U22954 (N_22954,N_21038,N_21890);
nor U22955 (N_22955,N_20860,N_20428);
or U22956 (N_22956,N_20367,N_21946);
xor U22957 (N_22957,N_21977,N_21018);
nor U22958 (N_22958,N_20168,N_20548);
or U22959 (N_22959,N_20686,N_20545);
nand U22960 (N_22960,N_21469,N_20233);
xnor U22961 (N_22961,N_21252,N_21781);
nor U22962 (N_22962,N_21009,N_20639);
or U22963 (N_22963,N_20259,N_20710);
nand U22964 (N_22964,N_20181,N_20212);
and U22965 (N_22965,N_20357,N_21229);
nor U22966 (N_22966,N_20035,N_20503);
nand U22967 (N_22967,N_20248,N_20709);
nor U22968 (N_22968,N_20042,N_20378);
nand U22969 (N_22969,N_20712,N_20981);
xnor U22970 (N_22970,N_20313,N_20290);
nand U22971 (N_22971,N_20208,N_20995);
nand U22972 (N_22972,N_21243,N_21143);
nor U22973 (N_22973,N_20982,N_20926);
nor U22974 (N_22974,N_20640,N_20387);
xnor U22975 (N_22975,N_20124,N_21473);
and U22976 (N_22976,N_21913,N_20107);
and U22977 (N_22977,N_21365,N_21567);
xnor U22978 (N_22978,N_21391,N_21696);
and U22979 (N_22979,N_21198,N_20051);
nor U22980 (N_22980,N_21185,N_21741);
xnor U22981 (N_22981,N_21343,N_20676);
and U22982 (N_22982,N_21052,N_20666);
xor U22983 (N_22983,N_21701,N_21053);
xor U22984 (N_22984,N_21451,N_20787);
and U22985 (N_22985,N_21087,N_20175);
or U22986 (N_22986,N_21421,N_21327);
nor U22987 (N_22987,N_20980,N_21012);
nand U22988 (N_22988,N_21669,N_21215);
or U22989 (N_22989,N_21434,N_20299);
and U22990 (N_22990,N_20796,N_20071);
nand U22991 (N_22991,N_21814,N_21131);
and U22992 (N_22992,N_21031,N_21985);
xnor U22993 (N_22993,N_20439,N_20286);
xor U22994 (N_22994,N_20660,N_21842);
nor U22995 (N_22995,N_21689,N_21838);
xnor U22996 (N_22996,N_21206,N_21356);
xnor U22997 (N_22997,N_20924,N_21790);
nand U22998 (N_22998,N_20020,N_21723);
or U22999 (N_22999,N_21007,N_20007);
nor U23000 (N_23000,N_20981,N_21610);
or U23001 (N_23001,N_20819,N_21314);
nor U23002 (N_23002,N_20669,N_21726);
xor U23003 (N_23003,N_20100,N_20865);
nand U23004 (N_23004,N_20981,N_21999);
and U23005 (N_23005,N_20551,N_20725);
or U23006 (N_23006,N_20975,N_20718);
or U23007 (N_23007,N_20813,N_21968);
nor U23008 (N_23008,N_21240,N_20443);
nor U23009 (N_23009,N_20409,N_20759);
nand U23010 (N_23010,N_21779,N_21439);
nor U23011 (N_23011,N_20866,N_21887);
nor U23012 (N_23012,N_20021,N_21091);
nor U23013 (N_23013,N_21688,N_21843);
or U23014 (N_23014,N_21258,N_21903);
nor U23015 (N_23015,N_20263,N_21752);
xnor U23016 (N_23016,N_21330,N_21509);
and U23017 (N_23017,N_20332,N_21189);
and U23018 (N_23018,N_20513,N_21768);
and U23019 (N_23019,N_20622,N_21988);
nor U23020 (N_23020,N_20757,N_20189);
and U23021 (N_23021,N_20182,N_21043);
nand U23022 (N_23022,N_21855,N_21640);
xnor U23023 (N_23023,N_20908,N_20578);
and U23024 (N_23024,N_21992,N_20692);
nor U23025 (N_23025,N_21449,N_21636);
xnor U23026 (N_23026,N_21979,N_20815);
or U23027 (N_23027,N_21879,N_20711);
or U23028 (N_23028,N_21360,N_20352);
and U23029 (N_23029,N_21225,N_21317);
nand U23030 (N_23030,N_20844,N_21463);
or U23031 (N_23031,N_21973,N_21063);
nand U23032 (N_23032,N_20260,N_20990);
nor U23033 (N_23033,N_21495,N_21972);
and U23034 (N_23034,N_21955,N_21614);
nand U23035 (N_23035,N_21074,N_21749);
nor U23036 (N_23036,N_20129,N_20215);
xor U23037 (N_23037,N_20357,N_21428);
or U23038 (N_23038,N_20543,N_20745);
or U23039 (N_23039,N_20453,N_20486);
nor U23040 (N_23040,N_21143,N_21057);
nand U23041 (N_23041,N_20891,N_20655);
xnor U23042 (N_23042,N_20103,N_21326);
nor U23043 (N_23043,N_20565,N_21604);
and U23044 (N_23044,N_20066,N_21328);
xor U23045 (N_23045,N_21667,N_21878);
nand U23046 (N_23046,N_21652,N_20147);
xor U23047 (N_23047,N_20761,N_21016);
nand U23048 (N_23048,N_20067,N_20142);
xnor U23049 (N_23049,N_20535,N_20913);
nor U23050 (N_23050,N_21116,N_21118);
and U23051 (N_23051,N_21942,N_21739);
xnor U23052 (N_23052,N_20305,N_20503);
xor U23053 (N_23053,N_20920,N_21546);
nand U23054 (N_23054,N_21960,N_20841);
nand U23055 (N_23055,N_20081,N_21755);
nor U23056 (N_23056,N_20753,N_21148);
xnor U23057 (N_23057,N_20568,N_20239);
or U23058 (N_23058,N_21204,N_20473);
or U23059 (N_23059,N_20863,N_21570);
and U23060 (N_23060,N_20504,N_20658);
nand U23061 (N_23061,N_21288,N_20695);
nor U23062 (N_23062,N_20062,N_21482);
nor U23063 (N_23063,N_20240,N_21905);
nor U23064 (N_23064,N_20392,N_20208);
and U23065 (N_23065,N_20631,N_21218);
xnor U23066 (N_23066,N_20308,N_21148);
or U23067 (N_23067,N_21831,N_21928);
nor U23068 (N_23068,N_21964,N_21312);
nand U23069 (N_23069,N_20744,N_20711);
nor U23070 (N_23070,N_21946,N_20621);
xnor U23071 (N_23071,N_20411,N_21438);
xnor U23072 (N_23072,N_21648,N_20780);
or U23073 (N_23073,N_20316,N_21573);
nor U23074 (N_23074,N_21752,N_21684);
or U23075 (N_23075,N_21538,N_20105);
xor U23076 (N_23076,N_21042,N_20729);
nor U23077 (N_23077,N_20505,N_20773);
xnor U23078 (N_23078,N_21837,N_20394);
nand U23079 (N_23079,N_20714,N_20380);
nor U23080 (N_23080,N_20408,N_21986);
and U23081 (N_23081,N_21166,N_21757);
xnor U23082 (N_23082,N_20152,N_20523);
and U23083 (N_23083,N_20891,N_20198);
or U23084 (N_23084,N_21897,N_21526);
nor U23085 (N_23085,N_20880,N_21265);
and U23086 (N_23086,N_20693,N_21607);
xnor U23087 (N_23087,N_21971,N_21052);
or U23088 (N_23088,N_20844,N_20408);
nor U23089 (N_23089,N_20568,N_21863);
or U23090 (N_23090,N_21329,N_20433);
and U23091 (N_23091,N_21319,N_20656);
and U23092 (N_23092,N_20972,N_21700);
and U23093 (N_23093,N_21020,N_20365);
or U23094 (N_23094,N_21699,N_21266);
nand U23095 (N_23095,N_21465,N_21363);
and U23096 (N_23096,N_20860,N_20639);
nand U23097 (N_23097,N_21684,N_20532);
xor U23098 (N_23098,N_20836,N_21000);
nand U23099 (N_23099,N_20103,N_20029);
nand U23100 (N_23100,N_20667,N_21118);
nand U23101 (N_23101,N_20541,N_20119);
and U23102 (N_23102,N_21084,N_21460);
or U23103 (N_23103,N_21199,N_21791);
nor U23104 (N_23104,N_21607,N_21541);
and U23105 (N_23105,N_21168,N_20489);
nor U23106 (N_23106,N_21203,N_21975);
xnor U23107 (N_23107,N_20627,N_20262);
and U23108 (N_23108,N_20449,N_20200);
xnor U23109 (N_23109,N_20442,N_21698);
xnor U23110 (N_23110,N_20874,N_21536);
xnor U23111 (N_23111,N_20817,N_21718);
or U23112 (N_23112,N_21293,N_21711);
or U23113 (N_23113,N_21296,N_21042);
and U23114 (N_23114,N_20037,N_20656);
and U23115 (N_23115,N_20988,N_21009);
or U23116 (N_23116,N_21373,N_20378);
and U23117 (N_23117,N_20734,N_20727);
xor U23118 (N_23118,N_20449,N_20100);
nor U23119 (N_23119,N_20679,N_20879);
or U23120 (N_23120,N_20315,N_21821);
or U23121 (N_23121,N_21821,N_21634);
nand U23122 (N_23122,N_20326,N_20875);
xor U23123 (N_23123,N_20509,N_21801);
nor U23124 (N_23124,N_20557,N_20550);
nor U23125 (N_23125,N_20566,N_20663);
and U23126 (N_23126,N_21082,N_20022);
nand U23127 (N_23127,N_20610,N_21401);
or U23128 (N_23128,N_21823,N_21561);
or U23129 (N_23129,N_21388,N_20350);
xor U23130 (N_23130,N_20384,N_20302);
nand U23131 (N_23131,N_20674,N_21397);
nand U23132 (N_23132,N_20354,N_20458);
xor U23133 (N_23133,N_20173,N_21501);
or U23134 (N_23134,N_20529,N_20970);
nor U23135 (N_23135,N_21297,N_21087);
and U23136 (N_23136,N_21314,N_20760);
nand U23137 (N_23137,N_20112,N_21700);
or U23138 (N_23138,N_20765,N_20860);
nor U23139 (N_23139,N_21206,N_20848);
nand U23140 (N_23140,N_21638,N_20680);
and U23141 (N_23141,N_21261,N_20502);
and U23142 (N_23142,N_21041,N_21980);
xor U23143 (N_23143,N_20368,N_20956);
and U23144 (N_23144,N_21341,N_21785);
xnor U23145 (N_23145,N_21444,N_21556);
or U23146 (N_23146,N_20403,N_20484);
nor U23147 (N_23147,N_20129,N_21782);
or U23148 (N_23148,N_20018,N_20821);
or U23149 (N_23149,N_21125,N_21517);
nor U23150 (N_23150,N_20014,N_20852);
or U23151 (N_23151,N_20243,N_21250);
and U23152 (N_23152,N_20509,N_21999);
nor U23153 (N_23153,N_20991,N_21329);
nor U23154 (N_23154,N_21929,N_21754);
or U23155 (N_23155,N_20568,N_21943);
or U23156 (N_23156,N_20145,N_20399);
nor U23157 (N_23157,N_21603,N_20448);
and U23158 (N_23158,N_20073,N_21147);
nor U23159 (N_23159,N_20280,N_21683);
and U23160 (N_23160,N_21539,N_20355);
nor U23161 (N_23161,N_20838,N_20038);
and U23162 (N_23162,N_20024,N_20400);
or U23163 (N_23163,N_21743,N_20832);
and U23164 (N_23164,N_21013,N_20443);
and U23165 (N_23165,N_20780,N_20302);
or U23166 (N_23166,N_20175,N_20487);
nor U23167 (N_23167,N_21422,N_20599);
nand U23168 (N_23168,N_20200,N_21095);
and U23169 (N_23169,N_21534,N_21807);
or U23170 (N_23170,N_20707,N_20611);
nor U23171 (N_23171,N_20609,N_20379);
nand U23172 (N_23172,N_20788,N_21852);
xnor U23173 (N_23173,N_21938,N_20903);
xnor U23174 (N_23174,N_21764,N_20077);
nor U23175 (N_23175,N_20867,N_20479);
xor U23176 (N_23176,N_21375,N_21244);
or U23177 (N_23177,N_21425,N_21804);
nor U23178 (N_23178,N_21190,N_21540);
or U23179 (N_23179,N_21860,N_21344);
xnor U23180 (N_23180,N_20922,N_20608);
nand U23181 (N_23181,N_21308,N_21674);
xnor U23182 (N_23182,N_20780,N_20338);
xnor U23183 (N_23183,N_20592,N_21577);
and U23184 (N_23184,N_21309,N_21230);
and U23185 (N_23185,N_21105,N_21875);
and U23186 (N_23186,N_21464,N_21190);
nor U23187 (N_23187,N_20186,N_20480);
or U23188 (N_23188,N_21591,N_20797);
nor U23189 (N_23189,N_21980,N_20515);
or U23190 (N_23190,N_20168,N_21261);
xnor U23191 (N_23191,N_21931,N_21518);
nand U23192 (N_23192,N_20438,N_20162);
nand U23193 (N_23193,N_21341,N_20071);
nor U23194 (N_23194,N_20231,N_20692);
xor U23195 (N_23195,N_20219,N_21263);
and U23196 (N_23196,N_20705,N_21230);
xor U23197 (N_23197,N_21463,N_21943);
nand U23198 (N_23198,N_20821,N_21123);
nand U23199 (N_23199,N_20223,N_20497);
and U23200 (N_23200,N_21386,N_20067);
nand U23201 (N_23201,N_20159,N_21202);
nand U23202 (N_23202,N_20861,N_20280);
nor U23203 (N_23203,N_20348,N_21868);
nor U23204 (N_23204,N_20594,N_20160);
and U23205 (N_23205,N_21532,N_20203);
nor U23206 (N_23206,N_21025,N_20104);
nor U23207 (N_23207,N_20088,N_21178);
nand U23208 (N_23208,N_21798,N_20503);
nand U23209 (N_23209,N_21350,N_20216);
nor U23210 (N_23210,N_21193,N_20738);
nand U23211 (N_23211,N_20566,N_20414);
or U23212 (N_23212,N_21677,N_21460);
nor U23213 (N_23213,N_20698,N_21265);
nor U23214 (N_23214,N_21465,N_21232);
nand U23215 (N_23215,N_21520,N_21096);
nor U23216 (N_23216,N_20801,N_20320);
xor U23217 (N_23217,N_20230,N_20144);
and U23218 (N_23218,N_20600,N_21959);
nor U23219 (N_23219,N_20316,N_21584);
and U23220 (N_23220,N_20618,N_21628);
xor U23221 (N_23221,N_20844,N_21649);
or U23222 (N_23222,N_21974,N_21303);
xnor U23223 (N_23223,N_20456,N_21839);
or U23224 (N_23224,N_20244,N_20454);
nor U23225 (N_23225,N_21492,N_20906);
nand U23226 (N_23226,N_20310,N_20538);
nor U23227 (N_23227,N_21993,N_21751);
xor U23228 (N_23228,N_20021,N_21567);
nor U23229 (N_23229,N_21522,N_20643);
or U23230 (N_23230,N_21794,N_20457);
xor U23231 (N_23231,N_20180,N_21455);
nand U23232 (N_23232,N_21513,N_21171);
xor U23233 (N_23233,N_21373,N_20849);
and U23234 (N_23234,N_20735,N_20639);
or U23235 (N_23235,N_20660,N_21807);
nor U23236 (N_23236,N_21546,N_20937);
or U23237 (N_23237,N_20695,N_20077);
xnor U23238 (N_23238,N_20519,N_20455);
or U23239 (N_23239,N_20863,N_20962);
nand U23240 (N_23240,N_21499,N_21454);
nor U23241 (N_23241,N_20484,N_20433);
and U23242 (N_23242,N_21578,N_20761);
xor U23243 (N_23243,N_21538,N_21485);
nand U23244 (N_23244,N_20272,N_20883);
nand U23245 (N_23245,N_21663,N_20221);
xnor U23246 (N_23246,N_21777,N_20700);
nor U23247 (N_23247,N_21945,N_20413);
nor U23248 (N_23248,N_20247,N_20223);
nand U23249 (N_23249,N_21840,N_20711);
xnor U23250 (N_23250,N_20640,N_20961);
nor U23251 (N_23251,N_20483,N_20927);
and U23252 (N_23252,N_21237,N_20277);
and U23253 (N_23253,N_21574,N_20329);
and U23254 (N_23254,N_20437,N_21557);
nor U23255 (N_23255,N_21535,N_20547);
and U23256 (N_23256,N_21573,N_20315);
nor U23257 (N_23257,N_20680,N_21989);
nand U23258 (N_23258,N_21686,N_21306);
nand U23259 (N_23259,N_20720,N_21025);
nand U23260 (N_23260,N_21416,N_21688);
nor U23261 (N_23261,N_21657,N_20752);
nor U23262 (N_23262,N_20010,N_20913);
or U23263 (N_23263,N_21669,N_21183);
and U23264 (N_23264,N_21584,N_20105);
or U23265 (N_23265,N_20789,N_21166);
or U23266 (N_23266,N_20184,N_20539);
xnor U23267 (N_23267,N_21357,N_20200);
or U23268 (N_23268,N_20866,N_20428);
nor U23269 (N_23269,N_20566,N_20058);
xor U23270 (N_23270,N_21164,N_21729);
xor U23271 (N_23271,N_20709,N_20331);
or U23272 (N_23272,N_21835,N_21185);
nand U23273 (N_23273,N_21835,N_20756);
and U23274 (N_23274,N_20866,N_21546);
nor U23275 (N_23275,N_21316,N_20542);
or U23276 (N_23276,N_21592,N_20815);
nor U23277 (N_23277,N_21800,N_20270);
nand U23278 (N_23278,N_20655,N_21971);
or U23279 (N_23279,N_21857,N_21017);
nand U23280 (N_23280,N_21997,N_20732);
nor U23281 (N_23281,N_20772,N_20361);
and U23282 (N_23282,N_20198,N_21409);
xnor U23283 (N_23283,N_20927,N_21978);
nand U23284 (N_23284,N_20028,N_20292);
and U23285 (N_23285,N_21052,N_20304);
nor U23286 (N_23286,N_21700,N_21467);
nand U23287 (N_23287,N_20393,N_21866);
nand U23288 (N_23288,N_20033,N_21708);
nor U23289 (N_23289,N_21356,N_21499);
nand U23290 (N_23290,N_20232,N_20271);
and U23291 (N_23291,N_20089,N_20156);
and U23292 (N_23292,N_21433,N_20363);
and U23293 (N_23293,N_20862,N_20818);
and U23294 (N_23294,N_20132,N_20723);
nand U23295 (N_23295,N_21593,N_21079);
or U23296 (N_23296,N_20422,N_20002);
nand U23297 (N_23297,N_21699,N_20169);
nor U23298 (N_23298,N_20257,N_21564);
and U23299 (N_23299,N_21321,N_20518);
nor U23300 (N_23300,N_20602,N_21896);
xnor U23301 (N_23301,N_21013,N_21096);
or U23302 (N_23302,N_20580,N_21231);
nor U23303 (N_23303,N_20846,N_21657);
and U23304 (N_23304,N_21071,N_20876);
nand U23305 (N_23305,N_20046,N_20059);
xnor U23306 (N_23306,N_20417,N_21509);
xnor U23307 (N_23307,N_20906,N_21598);
and U23308 (N_23308,N_21684,N_20794);
xnor U23309 (N_23309,N_20209,N_20722);
nand U23310 (N_23310,N_20887,N_20369);
nand U23311 (N_23311,N_20360,N_20901);
nor U23312 (N_23312,N_20721,N_21337);
nand U23313 (N_23313,N_21735,N_20893);
xor U23314 (N_23314,N_20716,N_20910);
xor U23315 (N_23315,N_20581,N_21276);
and U23316 (N_23316,N_21566,N_21076);
or U23317 (N_23317,N_21476,N_21965);
nor U23318 (N_23318,N_21884,N_20405);
xnor U23319 (N_23319,N_20138,N_20458);
xnor U23320 (N_23320,N_21768,N_21749);
or U23321 (N_23321,N_20306,N_21944);
nand U23322 (N_23322,N_20788,N_21702);
and U23323 (N_23323,N_20311,N_20038);
xnor U23324 (N_23324,N_21094,N_20587);
nand U23325 (N_23325,N_20208,N_20056);
and U23326 (N_23326,N_21102,N_20435);
xnor U23327 (N_23327,N_21413,N_20097);
nor U23328 (N_23328,N_21715,N_21593);
nor U23329 (N_23329,N_20734,N_20357);
nand U23330 (N_23330,N_21995,N_21210);
nor U23331 (N_23331,N_20241,N_21211);
and U23332 (N_23332,N_21692,N_20500);
nor U23333 (N_23333,N_20882,N_20852);
and U23334 (N_23334,N_20065,N_21264);
nand U23335 (N_23335,N_20490,N_21159);
xnor U23336 (N_23336,N_20340,N_21820);
nor U23337 (N_23337,N_20909,N_20216);
nor U23338 (N_23338,N_21683,N_20034);
and U23339 (N_23339,N_20916,N_20951);
and U23340 (N_23340,N_21973,N_20158);
xnor U23341 (N_23341,N_21092,N_21281);
nor U23342 (N_23342,N_20314,N_20605);
nor U23343 (N_23343,N_20646,N_20191);
xnor U23344 (N_23344,N_21256,N_21136);
nand U23345 (N_23345,N_20099,N_20468);
nor U23346 (N_23346,N_20347,N_21120);
xnor U23347 (N_23347,N_20584,N_21479);
nand U23348 (N_23348,N_20655,N_21838);
xor U23349 (N_23349,N_20635,N_20077);
nor U23350 (N_23350,N_21157,N_21062);
xnor U23351 (N_23351,N_21654,N_20591);
nor U23352 (N_23352,N_20241,N_20359);
or U23353 (N_23353,N_21497,N_21836);
nand U23354 (N_23354,N_21360,N_21303);
xor U23355 (N_23355,N_21282,N_21311);
nand U23356 (N_23356,N_20823,N_21855);
nand U23357 (N_23357,N_21795,N_21411);
and U23358 (N_23358,N_21167,N_20780);
xnor U23359 (N_23359,N_20308,N_20598);
xnor U23360 (N_23360,N_20797,N_21807);
nand U23361 (N_23361,N_21180,N_20568);
xor U23362 (N_23362,N_20826,N_21948);
xor U23363 (N_23363,N_21686,N_21725);
or U23364 (N_23364,N_20414,N_20620);
and U23365 (N_23365,N_20385,N_21509);
or U23366 (N_23366,N_20753,N_20826);
and U23367 (N_23367,N_20187,N_20424);
nand U23368 (N_23368,N_20984,N_20286);
nand U23369 (N_23369,N_21055,N_20275);
and U23370 (N_23370,N_21957,N_21282);
nor U23371 (N_23371,N_21983,N_20290);
xor U23372 (N_23372,N_21762,N_20189);
and U23373 (N_23373,N_20833,N_21434);
or U23374 (N_23374,N_21218,N_21567);
xnor U23375 (N_23375,N_21044,N_21271);
nor U23376 (N_23376,N_20976,N_21875);
and U23377 (N_23377,N_20258,N_20589);
nor U23378 (N_23378,N_21511,N_21046);
or U23379 (N_23379,N_20023,N_20179);
nor U23380 (N_23380,N_21551,N_20361);
and U23381 (N_23381,N_21755,N_20422);
or U23382 (N_23382,N_20707,N_21492);
xnor U23383 (N_23383,N_21954,N_21754);
nand U23384 (N_23384,N_21636,N_20519);
nor U23385 (N_23385,N_21828,N_20904);
nor U23386 (N_23386,N_21236,N_20271);
nor U23387 (N_23387,N_21172,N_20943);
nand U23388 (N_23388,N_21464,N_21784);
nor U23389 (N_23389,N_20621,N_20620);
nand U23390 (N_23390,N_20007,N_20469);
nand U23391 (N_23391,N_20629,N_21102);
or U23392 (N_23392,N_21428,N_21410);
or U23393 (N_23393,N_20815,N_20113);
nand U23394 (N_23394,N_21186,N_21609);
xor U23395 (N_23395,N_20596,N_20636);
nor U23396 (N_23396,N_21151,N_21227);
nor U23397 (N_23397,N_20853,N_21167);
nor U23398 (N_23398,N_21143,N_20328);
xnor U23399 (N_23399,N_21837,N_20668);
nor U23400 (N_23400,N_21292,N_21698);
nand U23401 (N_23401,N_21016,N_20704);
and U23402 (N_23402,N_20516,N_20172);
nand U23403 (N_23403,N_20878,N_20480);
or U23404 (N_23404,N_21127,N_21028);
xor U23405 (N_23405,N_20147,N_20512);
or U23406 (N_23406,N_21911,N_20187);
nor U23407 (N_23407,N_21512,N_20514);
nand U23408 (N_23408,N_21873,N_21659);
nor U23409 (N_23409,N_21001,N_21074);
and U23410 (N_23410,N_21438,N_21916);
or U23411 (N_23411,N_20903,N_21339);
or U23412 (N_23412,N_21070,N_20522);
xor U23413 (N_23413,N_21797,N_21008);
nor U23414 (N_23414,N_20875,N_21502);
nor U23415 (N_23415,N_21903,N_21518);
xnor U23416 (N_23416,N_20264,N_20591);
or U23417 (N_23417,N_20299,N_20702);
xnor U23418 (N_23418,N_21853,N_20445);
nor U23419 (N_23419,N_20864,N_20971);
and U23420 (N_23420,N_20370,N_20942);
and U23421 (N_23421,N_20602,N_21409);
nand U23422 (N_23422,N_20655,N_21475);
nand U23423 (N_23423,N_21510,N_21403);
and U23424 (N_23424,N_20721,N_21086);
or U23425 (N_23425,N_21394,N_21850);
nor U23426 (N_23426,N_20811,N_21207);
or U23427 (N_23427,N_21887,N_21048);
and U23428 (N_23428,N_21992,N_21787);
nand U23429 (N_23429,N_21826,N_21739);
or U23430 (N_23430,N_20914,N_20597);
or U23431 (N_23431,N_21192,N_20041);
and U23432 (N_23432,N_20031,N_20131);
nand U23433 (N_23433,N_20210,N_21717);
nand U23434 (N_23434,N_20936,N_20180);
xnor U23435 (N_23435,N_20934,N_21710);
xor U23436 (N_23436,N_21094,N_20623);
or U23437 (N_23437,N_21968,N_20083);
nor U23438 (N_23438,N_20645,N_20068);
nor U23439 (N_23439,N_20506,N_21839);
nand U23440 (N_23440,N_21024,N_20634);
or U23441 (N_23441,N_20269,N_20919);
xnor U23442 (N_23442,N_20296,N_20540);
and U23443 (N_23443,N_20028,N_21740);
xnor U23444 (N_23444,N_20384,N_20334);
xor U23445 (N_23445,N_20782,N_21535);
and U23446 (N_23446,N_21284,N_20871);
or U23447 (N_23447,N_21076,N_20702);
xor U23448 (N_23448,N_20754,N_20197);
nand U23449 (N_23449,N_21700,N_21307);
xnor U23450 (N_23450,N_21377,N_20630);
nor U23451 (N_23451,N_20539,N_21237);
nor U23452 (N_23452,N_20753,N_21582);
and U23453 (N_23453,N_21954,N_21776);
xnor U23454 (N_23454,N_21084,N_21321);
and U23455 (N_23455,N_20454,N_21324);
nand U23456 (N_23456,N_21862,N_20766);
or U23457 (N_23457,N_21718,N_21096);
nand U23458 (N_23458,N_20582,N_20117);
nor U23459 (N_23459,N_20204,N_20635);
nand U23460 (N_23460,N_21335,N_21510);
xor U23461 (N_23461,N_20076,N_21793);
nand U23462 (N_23462,N_21523,N_20440);
nand U23463 (N_23463,N_21948,N_21381);
and U23464 (N_23464,N_21452,N_20579);
and U23465 (N_23465,N_20140,N_21263);
and U23466 (N_23466,N_20573,N_20559);
xor U23467 (N_23467,N_21632,N_21469);
nor U23468 (N_23468,N_21497,N_21594);
xor U23469 (N_23469,N_20386,N_20172);
nor U23470 (N_23470,N_20710,N_20120);
nor U23471 (N_23471,N_21573,N_21111);
nor U23472 (N_23472,N_21386,N_20451);
nand U23473 (N_23473,N_21609,N_21921);
or U23474 (N_23474,N_20076,N_21373);
and U23475 (N_23475,N_20374,N_20739);
or U23476 (N_23476,N_21327,N_20878);
xor U23477 (N_23477,N_20959,N_20049);
or U23478 (N_23478,N_21683,N_21087);
nand U23479 (N_23479,N_21184,N_21374);
and U23480 (N_23480,N_20374,N_21352);
nor U23481 (N_23481,N_21423,N_20938);
or U23482 (N_23482,N_20459,N_21524);
nand U23483 (N_23483,N_20976,N_20428);
or U23484 (N_23484,N_20399,N_20082);
xnor U23485 (N_23485,N_21853,N_21225);
xnor U23486 (N_23486,N_21775,N_21883);
and U23487 (N_23487,N_20525,N_21454);
nand U23488 (N_23488,N_20764,N_21512);
or U23489 (N_23489,N_20904,N_20855);
and U23490 (N_23490,N_20943,N_20043);
and U23491 (N_23491,N_20278,N_21059);
xor U23492 (N_23492,N_21926,N_21021);
and U23493 (N_23493,N_21509,N_21229);
xor U23494 (N_23494,N_21500,N_21875);
xnor U23495 (N_23495,N_20997,N_21282);
xor U23496 (N_23496,N_21587,N_20330);
nor U23497 (N_23497,N_20231,N_20472);
nand U23498 (N_23498,N_20280,N_20615);
xor U23499 (N_23499,N_21370,N_20087);
nor U23500 (N_23500,N_20422,N_20349);
nor U23501 (N_23501,N_20084,N_21587);
and U23502 (N_23502,N_20975,N_21036);
and U23503 (N_23503,N_20802,N_21783);
nor U23504 (N_23504,N_21734,N_20986);
or U23505 (N_23505,N_21023,N_21697);
nand U23506 (N_23506,N_21808,N_21227);
nor U23507 (N_23507,N_21025,N_21031);
nand U23508 (N_23508,N_20688,N_20550);
or U23509 (N_23509,N_21013,N_20510);
and U23510 (N_23510,N_20581,N_21205);
xor U23511 (N_23511,N_21305,N_21829);
nor U23512 (N_23512,N_20830,N_20206);
and U23513 (N_23513,N_20737,N_20139);
xor U23514 (N_23514,N_21509,N_20810);
nor U23515 (N_23515,N_21498,N_20179);
and U23516 (N_23516,N_20051,N_20131);
or U23517 (N_23517,N_20294,N_21648);
or U23518 (N_23518,N_21881,N_20801);
nand U23519 (N_23519,N_21375,N_21989);
nand U23520 (N_23520,N_21302,N_20152);
or U23521 (N_23521,N_21783,N_21565);
nand U23522 (N_23522,N_20942,N_20027);
xor U23523 (N_23523,N_20255,N_21569);
or U23524 (N_23524,N_20679,N_20055);
xnor U23525 (N_23525,N_20428,N_21620);
and U23526 (N_23526,N_21039,N_21423);
xor U23527 (N_23527,N_20236,N_21086);
and U23528 (N_23528,N_20888,N_20153);
and U23529 (N_23529,N_21291,N_20372);
nor U23530 (N_23530,N_21170,N_21781);
nor U23531 (N_23531,N_21065,N_21048);
or U23532 (N_23532,N_20705,N_20592);
nor U23533 (N_23533,N_20378,N_20897);
nor U23534 (N_23534,N_20432,N_21211);
nor U23535 (N_23535,N_20325,N_21708);
xnor U23536 (N_23536,N_20761,N_21602);
nor U23537 (N_23537,N_20511,N_20487);
nand U23538 (N_23538,N_20678,N_21324);
nand U23539 (N_23539,N_21868,N_21682);
xor U23540 (N_23540,N_20239,N_21760);
and U23541 (N_23541,N_21051,N_21962);
xor U23542 (N_23542,N_21081,N_21815);
nor U23543 (N_23543,N_21830,N_21622);
xor U23544 (N_23544,N_20066,N_20969);
xor U23545 (N_23545,N_21974,N_20862);
nor U23546 (N_23546,N_21121,N_21615);
nand U23547 (N_23547,N_21362,N_20786);
and U23548 (N_23548,N_20707,N_21594);
nor U23549 (N_23549,N_21543,N_20619);
nor U23550 (N_23550,N_21634,N_20725);
nand U23551 (N_23551,N_21801,N_20262);
and U23552 (N_23552,N_21389,N_21412);
nor U23553 (N_23553,N_20176,N_21624);
nor U23554 (N_23554,N_20463,N_20781);
and U23555 (N_23555,N_21320,N_20248);
nand U23556 (N_23556,N_20525,N_21821);
xnor U23557 (N_23557,N_20474,N_20332);
nand U23558 (N_23558,N_20291,N_20374);
xnor U23559 (N_23559,N_20056,N_20233);
nand U23560 (N_23560,N_20671,N_20994);
or U23561 (N_23561,N_20189,N_21550);
nor U23562 (N_23562,N_21141,N_21368);
and U23563 (N_23563,N_20911,N_21906);
xor U23564 (N_23564,N_20700,N_21208);
nor U23565 (N_23565,N_21778,N_21484);
nor U23566 (N_23566,N_21234,N_21759);
nor U23567 (N_23567,N_21147,N_21785);
xnor U23568 (N_23568,N_21294,N_21502);
and U23569 (N_23569,N_20273,N_20455);
and U23570 (N_23570,N_20898,N_21941);
or U23571 (N_23571,N_21617,N_21995);
nor U23572 (N_23572,N_21574,N_20560);
nand U23573 (N_23573,N_21366,N_21815);
and U23574 (N_23574,N_21104,N_20130);
xor U23575 (N_23575,N_20099,N_21562);
or U23576 (N_23576,N_20348,N_20909);
nand U23577 (N_23577,N_20871,N_20215);
nor U23578 (N_23578,N_21919,N_21319);
nor U23579 (N_23579,N_21055,N_20455);
or U23580 (N_23580,N_21416,N_21597);
nor U23581 (N_23581,N_21671,N_20962);
xnor U23582 (N_23582,N_20876,N_21134);
nor U23583 (N_23583,N_20979,N_21095);
nand U23584 (N_23584,N_20866,N_20870);
or U23585 (N_23585,N_21885,N_20067);
xor U23586 (N_23586,N_21045,N_21585);
xnor U23587 (N_23587,N_21839,N_20312);
xor U23588 (N_23588,N_20014,N_20367);
and U23589 (N_23589,N_20156,N_21245);
and U23590 (N_23590,N_20239,N_21493);
or U23591 (N_23591,N_21604,N_21591);
or U23592 (N_23592,N_20477,N_20910);
nor U23593 (N_23593,N_20521,N_20868);
and U23594 (N_23594,N_20770,N_20257);
nand U23595 (N_23595,N_21863,N_20247);
nor U23596 (N_23596,N_21987,N_20254);
and U23597 (N_23597,N_21412,N_21073);
nand U23598 (N_23598,N_20950,N_21134);
nor U23599 (N_23599,N_20391,N_21209);
and U23600 (N_23600,N_21670,N_20769);
and U23601 (N_23601,N_21354,N_21349);
and U23602 (N_23602,N_21397,N_21814);
nor U23603 (N_23603,N_20402,N_21233);
or U23604 (N_23604,N_21526,N_21495);
or U23605 (N_23605,N_20968,N_20388);
or U23606 (N_23606,N_21376,N_20311);
and U23607 (N_23607,N_21562,N_21116);
and U23608 (N_23608,N_20518,N_20992);
nand U23609 (N_23609,N_20160,N_20399);
xor U23610 (N_23610,N_21366,N_20326);
xor U23611 (N_23611,N_21544,N_20627);
xnor U23612 (N_23612,N_21393,N_21171);
and U23613 (N_23613,N_21626,N_20795);
xor U23614 (N_23614,N_21472,N_21242);
nand U23615 (N_23615,N_21708,N_21691);
or U23616 (N_23616,N_20019,N_20845);
xor U23617 (N_23617,N_21485,N_21525);
nor U23618 (N_23618,N_20767,N_21983);
nand U23619 (N_23619,N_21357,N_20955);
xnor U23620 (N_23620,N_21519,N_21053);
xor U23621 (N_23621,N_20037,N_20962);
and U23622 (N_23622,N_21239,N_21058);
nand U23623 (N_23623,N_21728,N_20301);
nor U23624 (N_23624,N_21287,N_21949);
or U23625 (N_23625,N_20495,N_20317);
and U23626 (N_23626,N_20934,N_21918);
and U23627 (N_23627,N_20081,N_21698);
xor U23628 (N_23628,N_20637,N_20280);
xnor U23629 (N_23629,N_20173,N_21231);
nand U23630 (N_23630,N_20043,N_21426);
nand U23631 (N_23631,N_21138,N_21846);
nor U23632 (N_23632,N_20800,N_21867);
or U23633 (N_23633,N_21875,N_20361);
nand U23634 (N_23634,N_21574,N_20124);
or U23635 (N_23635,N_20876,N_21487);
and U23636 (N_23636,N_21704,N_20381);
nor U23637 (N_23637,N_20690,N_21436);
or U23638 (N_23638,N_20218,N_21398);
nor U23639 (N_23639,N_20283,N_21704);
or U23640 (N_23640,N_21167,N_21005);
nand U23641 (N_23641,N_20166,N_21690);
xnor U23642 (N_23642,N_20657,N_21546);
xor U23643 (N_23643,N_20636,N_20750);
nor U23644 (N_23644,N_21943,N_21316);
and U23645 (N_23645,N_21966,N_21621);
nand U23646 (N_23646,N_20595,N_20944);
xnor U23647 (N_23647,N_20215,N_21657);
nor U23648 (N_23648,N_20472,N_21322);
and U23649 (N_23649,N_21257,N_20607);
and U23650 (N_23650,N_21460,N_21143);
and U23651 (N_23651,N_20785,N_21362);
nand U23652 (N_23652,N_21769,N_21938);
and U23653 (N_23653,N_20249,N_21420);
or U23654 (N_23654,N_21512,N_21568);
xnor U23655 (N_23655,N_21490,N_20671);
and U23656 (N_23656,N_21060,N_20536);
nor U23657 (N_23657,N_20315,N_20450);
nand U23658 (N_23658,N_20765,N_20633);
or U23659 (N_23659,N_20827,N_21263);
and U23660 (N_23660,N_21727,N_20966);
nand U23661 (N_23661,N_20010,N_21325);
nor U23662 (N_23662,N_21271,N_20008);
or U23663 (N_23663,N_21426,N_21233);
and U23664 (N_23664,N_20641,N_21787);
xnor U23665 (N_23665,N_21772,N_21797);
xnor U23666 (N_23666,N_21836,N_21563);
nor U23667 (N_23667,N_21159,N_21662);
nand U23668 (N_23668,N_21827,N_20288);
xor U23669 (N_23669,N_20091,N_21437);
and U23670 (N_23670,N_21237,N_20252);
nor U23671 (N_23671,N_21857,N_21579);
nor U23672 (N_23672,N_20373,N_21959);
or U23673 (N_23673,N_20613,N_21040);
nor U23674 (N_23674,N_21636,N_21115);
and U23675 (N_23675,N_21472,N_20702);
xnor U23676 (N_23676,N_20763,N_20197);
and U23677 (N_23677,N_20889,N_21983);
or U23678 (N_23678,N_20390,N_20609);
nand U23679 (N_23679,N_21534,N_21112);
nand U23680 (N_23680,N_21976,N_20278);
nor U23681 (N_23681,N_20623,N_21954);
or U23682 (N_23682,N_20399,N_20408);
nor U23683 (N_23683,N_21746,N_21465);
xnor U23684 (N_23684,N_21324,N_20618);
or U23685 (N_23685,N_20856,N_21926);
nor U23686 (N_23686,N_20147,N_20283);
and U23687 (N_23687,N_21293,N_21645);
and U23688 (N_23688,N_20123,N_21348);
xnor U23689 (N_23689,N_20690,N_21384);
and U23690 (N_23690,N_20572,N_20501);
nand U23691 (N_23691,N_21699,N_21978);
xnor U23692 (N_23692,N_20382,N_20332);
nand U23693 (N_23693,N_21466,N_20787);
nor U23694 (N_23694,N_21232,N_21858);
or U23695 (N_23695,N_20122,N_21536);
nand U23696 (N_23696,N_20603,N_20750);
xnor U23697 (N_23697,N_21140,N_21361);
xnor U23698 (N_23698,N_20800,N_21812);
or U23699 (N_23699,N_21441,N_20832);
nand U23700 (N_23700,N_21490,N_21536);
and U23701 (N_23701,N_21185,N_20167);
nor U23702 (N_23702,N_20042,N_21112);
or U23703 (N_23703,N_21303,N_20038);
or U23704 (N_23704,N_21741,N_21698);
xor U23705 (N_23705,N_21043,N_21593);
nor U23706 (N_23706,N_21793,N_20988);
and U23707 (N_23707,N_21740,N_20503);
nand U23708 (N_23708,N_20252,N_21593);
and U23709 (N_23709,N_20729,N_21487);
and U23710 (N_23710,N_20515,N_20877);
or U23711 (N_23711,N_21560,N_21693);
xnor U23712 (N_23712,N_21848,N_20402);
or U23713 (N_23713,N_21130,N_21956);
xnor U23714 (N_23714,N_21412,N_20850);
nor U23715 (N_23715,N_21509,N_21230);
or U23716 (N_23716,N_20270,N_20359);
xnor U23717 (N_23717,N_20330,N_21084);
xnor U23718 (N_23718,N_21819,N_20931);
xor U23719 (N_23719,N_20936,N_20076);
and U23720 (N_23720,N_20961,N_20973);
or U23721 (N_23721,N_21909,N_21080);
nand U23722 (N_23722,N_20267,N_21973);
xor U23723 (N_23723,N_21160,N_20610);
xor U23724 (N_23724,N_21413,N_20351);
nand U23725 (N_23725,N_20857,N_20688);
and U23726 (N_23726,N_20509,N_20669);
or U23727 (N_23727,N_20318,N_20971);
or U23728 (N_23728,N_20025,N_21871);
xnor U23729 (N_23729,N_20069,N_21985);
nor U23730 (N_23730,N_20234,N_21984);
nor U23731 (N_23731,N_21565,N_21198);
or U23732 (N_23732,N_21671,N_20242);
nand U23733 (N_23733,N_20700,N_20933);
nand U23734 (N_23734,N_20750,N_20404);
nor U23735 (N_23735,N_20116,N_20956);
or U23736 (N_23736,N_20813,N_20643);
nor U23737 (N_23737,N_20043,N_20962);
nand U23738 (N_23738,N_20929,N_21381);
xor U23739 (N_23739,N_20890,N_21323);
nor U23740 (N_23740,N_21989,N_20076);
or U23741 (N_23741,N_20048,N_20046);
and U23742 (N_23742,N_21477,N_21944);
or U23743 (N_23743,N_20136,N_21102);
nand U23744 (N_23744,N_21541,N_20841);
xor U23745 (N_23745,N_21396,N_20640);
nor U23746 (N_23746,N_21389,N_21932);
or U23747 (N_23747,N_21462,N_21958);
nor U23748 (N_23748,N_20457,N_21785);
and U23749 (N_23749,N_20177,N_20449);
nand U23750 (N_23750,N_21035,N_21131);
xor U23751 (N_23751,N_20761,N_21803);
nand U23752 (N_23752,N_20242,N_20167);
and U23753 (N_23753,N_20581,N_20214);
or U23754 (N_23754,N_21086,N_20222);
and U23755 (N_23755,N_20398,N_21469);
and U23756 (N_23756,N_20175,N_21808);
xor U23757 (N_23757,N_21946,N_20624);
nor U23758 (N_23758,N_20311,N_21537);
and U23759 (N_23759,N_21829,N_21044);
nand U23760 (N_23760,N_20240,N_21623);
nand U23761 (N_23761,N_21851,N_21415);
and U23762 (N_23762,N_21280,N_21003);
nand U23763 (N_23763,N_20369,N_21996);
or U23764 (N_23764,N_20869,N_21414);
xor U23765 (N_23765,N_20067,N_20209);
nor U23766 (N_23766,N_20109,N_20941);
xor U23767 (N_23767,N_21356,N_21740);
nand U23768 (N_23768,N_20192,N_20447);
or U23769 (N_23769,N_20983,N_20710);
and U23770 (N_23770,N_20091,N_20978);
nand U23771 (N_23771,N_20858,N_21926);
or U23772 (N_23772,N_20726,N_20142);
nand U23773 (N_23773,N_20860,N_21227);
or U23774 (N_23774,N_20913,N_21738);
and U23775 (N_23775,N_20025,N_21093);
and U23776 (N_23776,N_20131,N_20500);
or U23777 (N_23777,N_21798,N_20260);
and U23778 (N_23778,N_21499,N_20071);
or U23779 (N_23779,N_20160,N_20685);
nand U23780 (N_23780,N_21071,N_21471);
or U23781 (N_23781,N_21102,N_21506);
or U23782 (N_23782,N_20130,N_20165);
nand U23783 (N_23783,N_21799,N_21643);
and U23784 (N_23784,N_20157,N_21249);
nor U23785 (N_23785,N_20266,N_21382);
or U23786 (N_23786,N_20226,N_20382);
xnor U23787 (N_23787,N_20165,N_20339);
nand U23788 (N_23788,N_20880,N_21664);
and U23789 (N_23789,N_21173,N_20862);
xnor U23790 (N_23790,N_21929,N_20021);
and U23791 (N_23791,N_20208,N_20510);
nand U23792 (N_23792,N_21968,N_20249);
nor U23793 (N_23793,N_20677,N_21129);
and U23794 (N_23794,N_20140,N_21739);
nand U23795 (N_23795,N_21976,N_21654);
nand U23796 (N_23796,N_20311,N_20905);
xnor U23797 (N_23797,N_20097,N_21714);
nand U23798 (N_23798,N_20187,N_21714);
nand U23799 (N_23799,N_20775,N_21969);
nor U23800 (N_23800,N_20482,N_20945);
and U23801 (N_23801,N_20706,N_20830);
and U23802 (N_23802,N_21155,N_21972);
nand U23803 (N_23803,N_21086,N_20129);
nor U23804 (N_23804,N_21973,N_20688);
xnor U23805 (N_23805,N_21810,N_20698);
nor U23806 (N_23806,N_21353,N_20298);
or U23807 (N_23807,N_21834,N_20995);
nor U23808 (N_23808,N_20604,N_20956);
nor U23809 (N_23809,N_21927,N_20789);
xor U23810 (N_23810,N_21466,N_20002);
nor U23811 (N_23811,N_21893,N_20263);
and U23812 (N_23812,N_20928,N_20392);
and U23813 (N_23813,N_20946,N_20298);
nand U23814 (N_23814,N_20260,N_21884);
or U23815 (N_23815,N_20847,N_21151);
or U23816 (N_23816,N_20348,N_21197);
xor U23817 (N_23817,N_21965,N_20604);
xor U23818 (N_23818,N_20071,N_20320);
and U23819 (N_23819,N_20749,N_21744);
or U23820 (N_23820,N_21759,N_21365);
xor U23821 (N_23821,N_21104,N_21631);
xor U23822 (N_23822,N_21294,N_21584);
nor U23823 (N_23823,N_21499,N_21234);
xnor U23824 (N_23824,N_20905,N_21287);
and U23825 (N_23825,N_21025,N_20896);
and U23826 (N_23826,N_21470,N_20304);
or U23827 (N_23827,N_21421,N_21525);
and U23828 (N_23828,N_20248,N_20694);
and U23829 (N_23829,N_21611,N_20250);
nor U23830 (N_23830,N_21434,N_20767);
xor U23831 (N_23831,N_21394,N_20490);
or U23832 (N_23832,N_21130,N_20814);
xor U23833 (N_23833,N_20213,N_20673);
nor U23834 (N_23834,N_20825,N_21852);
nor U23835 (N_23835,N_20244,N_21442);
nor U23836 (N_23836,N_21961,N_20436);
and U23837 (N_23837,N_21147,N_21367);
or U23838 (N_23838,N_20601,N_21728);
nor U23839 (N_23839,N_21078,N_21759);
and U23840 (N_23840,N_20948,N_20538);
and U23841 (N_23841,N_21258,N_20186);
xnor U23842 (N_23842,N_20588,N_20234);
nor U23843 (N_23843,N_20855,N_21987);
or U23844 (N_23844,N_20656,N_21377);
and U23845 (N_23845,N_20338,N_20942);
xor U23846 (N_23846,N_20398,N_21336);
nand U23847 (N_23847,N_21529,N_21709);
xnor U23848 (N_23848,N_20163,N_21030);
or U23849 (N_23849,N_20275,N_21487);
and U23850 (N_23850,N_21069,N_21070);
and U23851 (N_23851,N_21088,N_20518);
xor U23852 (N_23852,N_21784,N_21699);
xor U23853 (N_23853,N_20883,N_20617);
nor U23854 (N_23854,N_21894,N_21090);
and U23855 (N_23855,N_21829,N_21706);
and U23856 (N_23856,N_20578,N_20957);
nor U23857 (N_23857,N_21827,N_20641);
nor U23858 (N_23858,N_20023,N_20104);
xnor U23859 (N_23859,N_20147,N_20071);
and U23860 (N_23860,N_21184,N_20515);
and U23861 (N_23861,N_21102,N_20679);
xor U23862 (N_23862,N_20653,N_21829);
or U23863 (N_23863,N_21827,N_20870);
nand U23864 (N_23864,N_21431,N_21410);
nand U23865 (N_23865,N_21053,N_20499);
xor U23866 (N_23866,N_20474,N_20339);
xor U23867 (N_23867,N_21306,N_20854);
nand U23868 (N_23868,N_20311,N_21472);
nand U23869 (N_23869,N_21052,N_20634);
and U23870 (N_23870,N_21331,N_20789);
and U23871 (N_23871,N_20293,N_21440);
and U23872 (N_23872,N_20422,N_21334);
nor U23873 (N_23873,N_21548,N_20815);
and U23874 (N_23874,N_20673,N_20365);
nand U23875 (N_23875,N_20556,N_21363);
xnor U23876 (N_23876,N_20029,N_21235);
xor U23877 (N_23877,N_21946,N_21045);
nand U23878 (N_23878,N_20930,N_20148);
xnor U23879 (N_23879,N_20210,N_21079);
xor U23880 (N_23880,N_20916,N_21957);
or U23881 (N_23881,N_20783,N_21007);
nor U23882 (N_23882,N_21008,N_21068);
nor U23883 (N_23883,N_20899,N_20524);
nor U23884 (N_23884,N_20441,N_21866);
nand U23885 (N_23885,N_21205,N_21207);
and U23886 (N_23886,N_21987,N_21018);
or U23887 (N_23887,N_21828,N_21116);
nand U23888 (N_23888,N_20648,N_20514);
or U23889 (N_23889,N_21532,N_20458);
xor U23890 (N_23890,N_21313,N_21595);
and U23891 (N_23891,N_21309,N_20844);
nand U23892 (N_23892,N_21902,N_20551);
nor U23893 (N_23893,N_20653,N_20169);
and U23894 (N_23894,N_21413,N_21541);
xor U23895 (N_23895,N_20526,N_21462);
or U23896 (N_23896,N_20374,N_21534);
xnor U23897 (N_23897,N_21184,N_21075);
nor U23898 (N_23898,N_21036,N_21851);
or U23899 (N_23899,N_21519,N_20644);
xnor U23900 (N_23900,N_20538,N_21578);
nor U23901 (N_23901,N_20849,N_21803);
and U23902 (N_23902,N_21405,N_20197);
nand U23903 (N_23903,N_21059,N_20263);
and U23904 (N_23904,N_20416,N_21756);
nand U23905 (N_23905,N_21011,N_21623);
nor U23906 (N_23906,N_21878,N_20061);
and U23907 (N_23907,N_20196,N_20846);
or U23908 (N_23908,N_20517,N_20625);
or U23909 (N_23909,N_21606,N_21510);
nor U23910 (N_23910,N_20149,N_21579);
or U23911 (N_23911,N_20334,N_21448);
xnor U23912 (N_23912,N_20476,N_21882);
xor U23913 (N_23913,N_20686,N_20441);
and U23914 (N_23914,N_21345,N_20853);
nor U23915 (N_23915,N_21510,N_21232);
and U23916 (N_23916,N_20387,N_20802);
nor U23917 (N_23917,N_21950,N_21706);
nor U23918 (N_23918,N_20060,N_21406);
xor U23919 (N_23919,N_21652,N_21783);
nand U23920 (N_23920,N_21738,N_21028);
or U23921 (N_23921,N_20643,N_21058);
nand U23922 (N_23922,N_20538,N_20816);
xnor U23923 (N_23923,N_20134,N_21054);
nand U23924 (N_23924,N_21378,N_20777);
and U23925 (N_23925,N_20028,N_20348);
or U23926 (N_23926,N_21125,N_20439);
xor U23927 (N_23927,N_20021,N_21313);
or U23928 (N_23928,N_21320,N_20558);
and U23929 (N_23929,N_20945,N_21392);
nand U23930 (N_23930,N_21572,N_20043);
or U23931 (N_23931,N_20301,N_21095);
nor U23932 (N_23932,N_20470,N_20972);
nand U23933 (N_23933,N_20944,N_20768);
nand U23934 (N_23934,N_21623,N_20063);
and U23935 (N_23935,N_20767,N_20690);
nand U23936 (N_23936,N_21983,N_21273);
nand U23937 (N_23937,N_21861,N_20709);
xnor U23938 (N_23938,N_21158,N_21116);
xnor U23939 (N_23939,N_20152,N_20619);
or U23940 (N_23940,N_21712,N_20860);
or U23941 (N_23941,N_21145,N_21865);
or U23942 (N_23942,N_20242,N_21782);
nand U23943 (N_23943,N_20177,N_20918);
nor U23944 (N_23944,N_21377,N_20448);
or U23945 (N_23945,N_21858,N_20998);
nor U23946 (N_23946,N_20158,N_21822);
xnor U23947 (N_23947,N_20619,N_21036);
nor U23948 (N_23948,N_21523,N_21433);
nand U23949 (N_23949,N_20384,N_21540);
or U23950 (N_23950,N_20182,N_20186);
or U23951 (N_23951,N_20873,N_21069);
nand U23952 (N_23952,N_20124,N_21488);
nand U23953 (N_23953,N_21824,N_21090);
nand U23954 (N_23954,N_20569,N_20674);
and U23955 (N_23955,N_21454,N_21249);
xnor U23956 (N_23956,N_21489,N_21875);
nor U23957 (N_23957,N_21282,N_20300);
or U23958 (N_23958,N_20457,N_20936);
nand U23959 (N_23959,N_20044,N_20487);
nand U23960 (N_23960,N_20336,N_21996);
nor U23961 (N_23961,N_20789,N_21597);
nand U23962 (N_23962,N_21793,N_20555);
or U23963 (N_23963,N_20613,N_20718);
or U23964 (N_23964,N_21609,N_20638);
and U23965 (N_23965,N_21542,N_21619);
or U23966 (N_23966,N_21066,N_20254);
and U23967 (N_23967,N_21238,N_21233);
nand U23968 (N_23968,N_20535,N_21977);
and U23969 (N_23969,N_21034,N_20443);
nand U23970 (N_23970,N_21231,N_20677);
or U23971 (N_23971,N_21829,N_21486);
xnor U23972 (N_23972,N_20962,N_20313);
and U23973 (N_23973,N_21247,N_21112);
nand U23974 (N_23974,N_20252,N_21436);
and U23975 (N_23975,N_21761,N_20924);
nor U23976 (N_23976,N_21948,N_21603);
nor U23977 (N_23977,N_20918,N_20361);
and U23978 (N_23978,N_20982,N_21392);
nand U23979 (N_23979,N_20524,N_21458);
nor U23980 (N_23980,N_21388,N_20398);
xnor U23981 (N_23981,N_20446,N_21161);
nor U23982 (N_23982,N_21590,N_20885);
nor U23983 (N_23983,N_20292,N_20341);
or U23984 (N_23984,N_20578,N_21298);
and U23985 (N_23985,N_20665,N_21696);
nand U23986 (N_23986,N_20215,N_20879);
nor U23987 (N_23987,N_21934,N_21565);
or U23988 (N_23988,N_21353,N_20691);
nand U23989 (N_23989,N_20200,N_21489);
xnor U23990 (N_23990,N_21438,N_21393);
and U23991 (N_23991,N_21163,N_21772);
and U23992 (N_23992,N_21063,N_20885);
or U23993 (N_23993,N_20794,N_21736);
nor U23994 (N_23994,N_21564,N_20484);
nand U23995 (N_23995,N_21080,N_20944);
nor U23996 (N_23996,N_20592,N_21211);
nand U23997 (N_23997,N_21124,N_21040);
or U23998 (N_23998,N_21043,N_20517);
nor U23999 (N_23999,N_21250,N_21314);
nand U24000 (N_24000,N_23888,N_23625);
and U24001 (N_24001,N_23808,N_23797);
nand U24002 (N_24002,N_23840,N_22640);
xor U24003 (N_24003,N_23597,N_23890);
or U24004 (N_24004,N_22485,N_22590);
or U24005 (N_24005,N_22778,N_23258);
or U24006 (N_24006,N_22619,N_23738);
nand U24007 (N_24007,N_23416,N_23837);
xnor U24008 (N_24008,N_23389,N_23197);
nand U24009 (N_24009,N_22612,N_22073);
and U24010 (N_24010,N_22569,N_22994);
nor U24011 (N_24011,N_22060,N_23380);
nor U24012 (N_24012,N_23792,N_22671);
xor U24013 (N_24013,N_22001,N_22470);
xnor U24014 (N_24014,N_23732,N_23291);
and U24015 (N_24015,N_22114,N_23278);
and U24016 (N_24016,N_23144,N_22055);
xnor U24017 (N_24017,N_23246,N_22704);
or U24018 (N_24018,N_23508,N_22685);
xnor U24019 (N_24019,N_23066,N_22582);
and U24020 (N_24020,N_22290,N_22875);
nand U24021 (N_24021,N_22996,N_23071);
nor U24022 (N_24022,N_23112,N_23742);
or U24023 (N_24023,N_23342,N_23406);
xor U24024 (N_24024,N_22100,N_22256);
or U24025 (N_24025,N_23984,N_22866);
xnor U24026 (N_24026,N_23567,N_22628);
nand U24027 (N_24027,N_23202,N_23214);
nor U24028 (N_24028,N_23233,N_22347);
nor U24029 (N_24029,N_22272,N_23968);
or U24030 (N_24030,N_23158,N_23675);
or U24031 (N_24031,N_23002,N_22145);
or U24032 (N_24032,N_23247,N_23515);
nand U24033 (N_24033,N_22969,N_23138);
or U24034 (N_24034,N_23566,N_22864);
or U24035 (N_24035,N_22963,N_23776);
and U24036 (N_24036,N_22607,N_22877);
xor U24037 (N_24037,N_23205,N_23286);
nor U24038 (N_24038,N_23726,N_23520);
and U24039 (N_24039,N_22561,N_22534);
nand U24040 (N_24040,N_22896,N_23412);
nand U24041 (N_24041,N_23501,N_22828);
and U24042 (N_24042,N_22756,N_23815);
xor U24043 (N_24043,N_23757,N_22647);
xor U24044 (N_24044,N_23404,N_23648);
xor U24045 (N_24045,N_23468,N_23407);
and U24046 (N_24046,N_23951,N_23062);
or U24047 (N_24047,N_23006,N_22511);
nor U24048 (N_24048,N_23419,N_23492);
and U24049 (N_24049,N_23834,N_23504);
and U24050 (N_24050,N_22317,N_23123);
nand U24051 (N_24051,N_23975,N_23737);
nand U24052 (N_24052,N_22108,N_22972);
and U24053 (N_24053,N_22935,N_22601);
or U24054 (N_24054,N_22509,N_22392);
nand U24055 (N_24055,N_22696,N_22116);
nand U24056 (N_24056,N_23836,N_22424);
and U24057 (N_24057,N_22960,N_23126);
nor U24058 (N_24058,N_22103,N_22901);
or U24059 (N_24059,N_22462,N_22128);
and U24060 (N_24060,N_23299,N_23616);
or U24061 (N_24061,N_23820,N_22023);
or U24062 (N_24062,N_23651,N_23403);
or U24063 (N_24063,N_22213,N_22542);
or U24064 (N_24064,N_23308,N_22384);
nor U24065 (N_24065,N_23230,N_23762);
xor U24066 (N_24066,N_23736,N_23098);
and U24067 (N_24067,N_23751,N_22414);
nor U24068 (N_24068,N_23064,N_22514);
nand U24069 (N_24069,N_23878,N_22596);
nor U24070 (N_24070,N_22927,N_22748);
xnor U24071 (N_24071,N_23476,N_22735);
xor U24072 (N_24072,N_22070,N_23718);
nor U24073 (N_24073,N_23816,N_22507);
or U24074 (N_24074,N_22217,N_22194);
nand U24075 (N_24075,N_22205,N_23946);
nor U24076 (N_24076,N_22147,N_23490);
nand U24077 (N_24077,N_23284,N_23856);
nand U24078 (N_24078,N_22107,N_23295);
xor U24079 (N_24079,N_22657,N_22312);
nor U24080 (N_24080,N_23601,N_22078);
nor U24081 (N_24081,N_22719,N_23541);
and U24082 (N_24082,N_22974,N_23459);
nand U24083 (N_24083,N_23473,N_22940);
and U24084 (N_24084,N_22769,N_23234);
nor U24085 (N_24085,N_22325,N_23640);
nand U24086 (N_24086,N_22483,N_22621);
nand U24087 (N_24087,N_23174,N_22587);
xor U24088 (N_24088,N_23188,N_22529);
xor U24089 (N_24089,N_23219,N_22228);
or U24090 (N_24090,N_23716,N_22495);
nor U24091 (N_24091,N_23485,N_22718);
and U24092 (N_24092,N_22936,N_22813);
xnor U24093 (N_24093,N_22500,N_22680);
nand U24094 (N_24094,N_22544,N_23210);
or U24095 (N_24095,N_23710,N_23220);
and U24096 (N_24096,N_22241,N_22439);
nor U24097 (N_24097,N_22859,N_22422);
xnor U24098 (N_24098,N_23790,N_23868);
nor U24099 (N_24099,N_23670,N_22929);
nand U24100 (N_24100,N_22123,N_22235);
or U24101 (N_24101,N_23912,N_22567);
or U24102 (N_24102,N_23899,N_22246);
nand U24103 (N_24103,N_22088,N_22221);
nor U24104 (N_24104,N_23615,N_23365);
xor U24105 (N_24105,N_23645,N_22860);
nand U24106 (N_24106,N_22588,N_23229);
nor U24107 (N_24107,N_22025,N_23740);
nor U24108 (N_24108,N_23239,N_22505);
and U24109 (N_24109,N_23019,N_22141);
nand U24110 (N_24110,N_22009,N_23654);
nor U24111 (N_24111,N_22665,N_22686);
nor U24112 (N_24112,N_22932,N_23594);
or U24113 (N_24113,N_23402,N_22703);
xnor U24114 (N_24114,N_22967,N_23417);
nand U24115 (N_24115,N_22789,N_23498);
nor U24116 (N_24116,N_23555,N_23578);
nor U24117 (N_24117,N_22081,N_23533);
nand U24118 (N_24118,N_22668,N_23216);
or U24119 (N_24119,N_22649,N_23829);
nand U24120 (N_24120,N_23510,N_23104);
nand U24121 (N_24121,N_23185,N_23125);
xor U24122 (N_24122,N_22785,N_22244);
xor U24123 (N_24123,N_23564,N_23032);
and U24124 (N_24124,N_23922,N_22597);
nand U24125 (N_24125,N_22034,N_22096);
and U24126 (N_24126,N_22386,N_23045);
or U24127 (N_24127,N_23761,N_22177);
nand U24128 (N_24128,N_23784,N_23956);
xor U24129 (N_24129,N_23558,N_22930);
or U24130 (N_24130,N_22068,N_22702);
nand U24131 (N_24131,N_23034,N_22402);
and U24132 (N_24132,N_23374,N_22399);
nor U24133 (N_24133,N_22800,N_23078);
xnor U24134 (N_24134,N_22618,N_23539);
xor U24135 (N_24135,N_22743,N_23785);
xnor U24136 (N_24136,N_22664,N_23712);
and U24137 (N_24137,N_23517,N_23474);
nand U24138 (N_24138,N_22822,N_23256);
and U24139 (N_24139,N_23979,N_22303);
xnor U24140 (N_24140,N_23409,N_23273);
nand U24141 (N_24141,N_22423,N_23580);
or U24142 (N_24142,N_23568,N_23522);
nand U24143 (N_24143,N_22315,N_22477);
xnor U24144 (N_24144,N_22302,N_23608);
nand U24145 (N_24145,N_22155,N_22636);
xor U24146 (N_24146,N_23181,N_23916);
or U24147 (N_24147,N_23854,N_22938);
nor U24148 (N_24148,N_23961,N_22982);
nand U24149 (N_24149,N_22045,N_23448);
or U24150 (N_24150,N_23176,N_22032);
xor U24151 (N_24151,N_23364,N_23546);
nor U24152 (N_24152,N_22188,N_22144);
or U24153 (N_24153,N_22682,N_22951);
nor U24154 (N_24154,N_23434,N_23772);
or U24155 (N_24155,N_22817,N_22455);
nand U24156 (N_24156,N_23363,N_23041);
or U24157 (N_24157,N_22053,N_22862);
xor U24158 (N_24158,N_23963,N_23162);
and U24159 (N_24159,N_22441,N_23186);
nand U24160 (N_24160,N_23664,N_23628);
xnor U24161 (N_24161,N_22202,N_22079);
nand U24162 (N_24162,N_23667,N_23074);
and U24163 (N_24163,N_23898,N_23068);
nor U24164 (N_24164,N_22799,N_23493);
xor U24165 (N_24165,N_22993,N_22486);
xnor U24166 (N_24166,N_23770,N_22513);
and U24167 (N_24167,N_23775,N_22566);
or U24168 (N_24168,N_23250,N_23788);
nor U24169 (N_24169,N_22924,N_23455);
nand U24170 (N_24170,N_22253,N_23845);
and U24171 (N_24171,N_22784,N_23551);
nor U24172 (N_24172,N_23189,N_22230);
nor U24173 (N_24173,N_22730,N_23149);
nand U24174 (N_24174,N_22091,N_22062);
nand U24175 (N_24175,N_22193,N_23631);
or U24176 (N_24176,N_22547,N_22454);
nor U24177 (N_24177,N_22069,N_23672);
nor U24178 (N_24178,N_22174,N_22678);
nand U24179 (N_24179,N_22178,N_22606);
or U24180 (N_24180,N_23987,N_23199);
or U24181 (N_24181,N_22129,N_23862);
or U24182 (N_24182,N_23766,N_22295);
and U24183 (N_24183,N_22964,N_22774);
nor U24184 (N_24184,N_22523,N_22432);
xor U24185 (N_24185,N_22706,N_22371);
or U24186 (N_24186,N_23613,N_23516);
nor U24187 (N_24187,N_23860,N_22987);
or U24188 (N_24188,N_23151,N_22989);
nor U24189 (N_24189,N_23894,N_23970);
or U24190 (N_24190,N_23549,N_22203);
or U24191 (N_24191,N_22175,N_23467);
and U24192 (N_24192,N_22641,N_22981);
and U24193 (N_24193,N_22268,N_23410);
and U24194 (N_24194,N_22200,N_22771);
nor U24195 (N_24195,N_22631,N_22157);
and U24196 (N_24196,N_22273,N_22809);
or U24197 (N_24197,N_23893,N_22843);
nor U24198 (N_24198,N_22627,N_22858);
or U24199 (N_24199,N_23122,N_23926);
nand U24200 (N_24200,N_23989,N_22440);
nor U24201 (N_24201,N_22979,N_23690);
and U24202 (N_24202,N_23128,N_23025);
or U24203 (N_24203,N_22975,N_22870);
or U24204 (N_24204,N_22388,N_22790);
nand U24205 (N_24205,N_22536,N_22834);
nand U24206 (N_24206,N_22017,N_22027);
nand U24207 (N_24207,N_23131,N_22707);
nand U24208 (N_24208,N_23662,N_22933);
nor U24209 (N_24209,N_22700,N_23428);
or U24210 (N_24210,N_23077,N_23787);
and U24211 (N_24211,N_23735,N_22459);
or U24212 (N_24212,N_22028,N_23966);
or U24213 (N_24213,N_22092,N_23702);
and U24214 (N_24214,N_23693,N_22267);
and U24215 (N_24215,N_22095,N_23620);
nand U24216 (N_24216,N_22797,N_23570);
xnor U24217 (N_24217,N_23084,N_23356);
or U24218 (N_24218,N_22435,N_22050);
xnor U24219 (N_24219,N_22443,N_23610);
nor U24220 (N_24220,N_23307,N_23336);
nand U24221 (N_24221,N_23604,N_23746);
nand U24222 (N_24222,N_23630,N_23629);
nor U24223 (N_24223,N_23418,N_23101);
and U24224 (N_24224,N_22180,N_23395);
nor U24225 (N_24225,N_23985,N_22265);
and U24226 (N_24226,N_23572,N_22321);
nand U24227 (N_24227,N_22442,N_23288);
nand U24228 (N_24228,N_22727,N_23942);
or U24229 (N_24229,N_23532,N_23769);
nor U24230 (N_24230,N_23014,N_22768);
or U24231 (N_24231,N_22620,N_23750);
xnor U24232 (N_24232,N_22097,N_22694);
xor U24233 (N_24233,N_23992,N_22844);
and U24234 (N_24234,N_22720,N_22660);
or U24235 (N_24235,N_23764,N_23925);
nand U24236 (N_24236,N_23838,N_22493);
and U24237 (N_24237,N_23777,N_23184);
and U24238 (N_24238,N_23782,N_22291);
or U24239 (N_24239,N_23324,N_23287);
and U24240 (N_24240,N_23312,N_22897);
nand U24241 (N_24241,N_23182,N_22824);
or U24242 (N_24242,N_23861,N_23626);
nand U24243 (N_24243,N_23298,N_23744);
xnor U24244 (N_24244,N_22146,N_22330);
nand U24245 (N_24245,N_23832,N_22254);
and U24246 (N_24246,N_23581,N_23323);
or U24247 (N_24247,N_22375,N_23279);
nor U24248 (N_24248,N_23110,N_23542);
nor U24249 (N_24249,N_22942,N_22250);
and U24250 (N_24250,N_22279,N_23146);
and U24251 (N_24251,N_22998,N_22074);
nor U24252 (N_24252,N_23754,N_22992);
nand U24253 (N_24253,N_23209,N_22830);
or U24254 (N_24254,N_22431,N_23261);
nand U24255 (N_24255,N_22489,N_22654);
nand U24256 (N_24256,N_23511,N_22506);
nand U24257 (N_24257,N_22338,N_22739);
xnor U24258 (N_24258,N_23683,N_23939);
or U24259 (N_24259,N_22595,N_22332);
nor U24260 (N_24260,N_23399,N_23132);
nand U24261 (N_24261,N_23573,N_22190);
or U24262 (N_24262,N_22447,N_23386);
nand U24263 (N_24263,N_22226,N_23526);
and U24264 (N_24264,N_22541,N_23571);
nand U24265 (N_24265,N_23907,N_23691);
nand U24266 (N_24266,N_22889,N_23315);
and U24267 (N_24267,N_22322,N_23505);
nand U24268 (N_24268,N_23431,N_22953);
nor U24269 (N_24269,N_23923,N_23130);
xor U24270 (N_24270,N_22808,N_23470);
nand U24271 (N_24271,N_22503,N_22015);
and U24272 (N_24272,N_23067,N_22658);
xnor U24273 (N_24273,N_22433,N_22363);
and U24274 (N_24274,N_22580,N_23408);
nand U24275 (N_24275,N_22840,N_22663);
and U24276 (N_24276,N_22258,N_23272);
or U24277 (N_24277,N_22342,N_22645);
nor U24278 (N_24278,N_23642,N_23663);
and U24279 (N_24279,N_23009,N_23060);
xor U24280 (N_24280,N_23269,N_22085);
nand U24281 (N_24281,N_22215,N_23348);
nor U24282 (N_24282,N_23618,N_22501);
or U24283 (N_24283,N_22818,N_22872);
nand U24284 (N_24284,N_23524,N_23668);
and U24285 (N_24285,N_22300,N_23357);
xor U24286 (N_24286,N_23812,N_22736);
xnor U24287 (N_24287,N_23495,N_23819);
nand U24288 (N_24288,N_23478,N_22555);
nand U24289 (N_24289,N_23429,N_22343);
or U24290 (N_24290,N_22684,N_22832);
or U24291 (N_24291,N_22584,N_23752);
and U24292 (N_24292,N_22943,N_22159);
and U24293 (N_24293,N_22122,N_23650);
or U24294 (N_24294,N_22810,N_22299);
xor U24295 (N_24295,N_22805,N_23852);
or U24296 (N_24296,N_23953,N_22754);
and U24297 (N_24297,N_23337,N_23947);
nand U24298 (N_24298,N_23634,N_22130);
or U24299 (N_24299,N_22031,N_23007);
and U24300 (N_24300,N_23392,N_23512);
nor U24301 (N_24301,N_23850,N_22170);
nor U24302 (N_24302,N_23557,N_23226);
or U24303 (N_24303,N_22276,N_23930);
nand U24304 (N_24304,N_22519,N_22950);
nor U24305 (N_24305,N_23183,N_23706);
and U24306 (N_24306,N_23413,N_23649);
nor U24307 (N_24307,N_22758,N_22398);
or U24308 (N_24308,N_22036,N_23767);
nand U24309 (N_24309,N_22233,N_23666);
nor U24310 (N_24310,N_22018,N_22357);
and U24311 (N_24311,N_23094,N_23698);
xnor U24312 (N_24312,N_23369,N_22054);
nand U24313 (N_24313,N_23822,N_22804);
or U24314 (N_24314,N_22731,N_22538);
nor U24315 (N_24315,N_22318,N_23240);
xnor U24316 (N_24316,N_23660,N_22775);
and U24317 (N_24317,N_23332,N_22187);
nand U24318 (N_24318,N_22655,N_22382);
and U24319 (N_24319,N_23266,N_23780);
nor U24320 (N_24320,N_22708,N_23910);
and U24321 (N_24321,N_22077,N_22653);
xor U24322 (N_24322,N_22562,N_23051);
or U24323 (N_24323,N_22478,N_22602);
and U24324 (N_24324,N_23056,N_23595);
xor U24325 (N_24325,N_23026,N_23367);
and U24326 (N_24326,N_23095,N_22494);
nand U24327 (N_24327,N_23282,N_22856);
or U24328 (N_24328,N_22554,N_23724);
nor U24329 (N_24329,N_22610,N_23316);
xor U24330 (N_24330,N_22038,N_22307);
nand U24331 (N_24331,N_22716,N_23606);
or U24332 (N_24332,N_23694,N_23786);
and U24333 (N_24333,N_22080,N_23534);
xnor U24334 (N_24334,N_22308,N_22126);
nor U24335 (N_24335,N_23321,N_22076);
nand U24336 (N_24336,N_23304,N_22183);
xor U24337 (N_24337,N_22356,N_23656);
xnor U24338 (N_24338,N_22344,N_23100);
xor U24339 (N_24339,N_23804,N_22568);
nor U24340 (N_24340,N_22851,N_22644);
and U24341 (N_24341,N_22037,N_23155);
nand U24342 (N_24342,N_23633,N_23243);
nor U24343 (N_24343,N_22301,N_22458);
nor U24344 (N_24344,N_23699,N_22520);
and U24345 (N_24345,N_23344,N_23781);
xor U24346 (N_24346,N_23089,N_22191);
xor U24347 (N_24347,N_23262,N_22586);
nand U24348 (N_24348,N_23749,N_23309);
nand U24349 (N_24349,N_22405,N_23795);
nand U24350 (N_24350,N_22777,N_23217);
xnor U24351 (N_24351,N_22101,N_22121);
and U24352 (N_24352,N_22359,N_23325);
xor U24353 (N_24353,N_23447,N_23129);
xnor U24354 (N_24354,N_23506,N_22229);
xnor U24355 (N_24355,N_22282,N_22354);
nor U24356 (N_24356,N_23867,N_23024);
nor U24357 (N_24357,N_22367,N_22624);
nand U24358 (N_24358,N_23998,N_22013);
or U24359 (N_24359,N_22259,N_22954);
nor U24360 (N_24360,N_23993,N_23994);
xor U24361 (N_24361,N_23603,N_23225);
nand U24362 (N_24362,N_23873,N_22890);
or U24363 (N_24363,N_23909,N_22581);
or U24364 (N_24364,N_23464,N_22029);
and U24365 (N_24365,N_22022,N_23658);
nor U24366 (N_24366,N_23345,N_23117);
nor U24367 (N_24367,N_22801,N_22537);
xor U24368 (N_24368,N_22182,N_23306);
nand U24369 (N_24369,N_22539,N_23143);
nand U24370 (N_24370,N_22977,N_22786);
and U24371 (N_24371,N_23954,N_22524);
nor U24372 (N_24372,N_22304,N_23167);
and U24373 (N_24373,N_22687,N_22556);
nor U24374 (N_24374,N_23294,N_23929);
nand U24375 (N_24375,N_22575,N_23591);
xnor U24376 (N_24376,N_23215,N_22886);
and U24377 (N_24377,N_22755,N_22614);
xnor U24378 (N_24378,N_23059,N_22196);
or U24379 (N_24379,N_23914,N_23015);
nand U24380 (N_24380,N_22946,N_23390);
or U24381 (N_24381,N_23465,N_23639);
nand U24382 (N_24382,N_22713,N_23164);
nor U24383 (N_24383,N_22089,N_23941);
and U24384 (N_24384,N_22361,N_22498);
or U24385 (N_24385,N_22915,N_23932);
nand U24386 (N_24386,N_22140,N_22849);
or U24387 (N_24387,N_23375,N_23713);
xnor U24388 (N_24388,N_23127,N_23612);
or U24389 (N_24389,N_22863,N_23887);
or U24390 (N_24390,N_23016,N_23538);
nor U24391 (N_24391,N_23343,N_23621);
nor U24392 (N_24392,N_23943,N_22289);
nor U24393 (N_24393,N_22421,N_23430);
nor U24394 (N_24394,N_22528,N_22156);
xnor U24395 (N_24395,N_22540,N_22512);
nor U24396 (N_24396,N_22873,N_22807);
and U24397 (N_24397,N_22094,N_23659);
or U24398 (N_24398,N_23647,N_22753);
and U24399 (N_24399,N_23688,N_22257);
and U24400 (N_24400,N_23244,N_22667);
xor U24401 (N_24401,N_23108,N_23013);
xnor U24402 (N_24402,N_22378,N_23673);
and U24403 (N_24403,N_23727,N_23696);
xor U24404 (N_24404,N_22585,N_23086);
xor U24405 (N_24405,N_22099,N_23685);
and U24406 (N_24406,N_23983,N_23397);
nand U24407 (N_24407,N_22571,N_22965);
or U24408 (N_24408,N_22340,N_22532);
xnor U24409 (N_24409,N_23935,N_23022);
xnor U24410 (N_24410,N_23228,N_23969);
and U24411 (N_24411,N_22803,N_23224);
xor U24412 (N_24412,N_22339,N_22016);
nor U24413 (N_24413,N_22161,N_23773);
nand U24414 (N_24414,N_23714,N_23384);
and U24415 (N_24415,N_22961,N_23160);
or U24416 (N_24416,N_22041,N_23759);
or U24417 (N_24417,N_22625,N_23988);
nand U24418 (N_24418,N_23807,N_22393);
xnor U24419 (N_24419,N_23454,N_23589);
or U24420 (N_24420,N_23318,N_23443);
and U24421 (N_24421,N_22823,N_23372);
nor U24422 (N_24422,N_22297,N_22728);
nand U24423 (N_24423,N_22725,N_22223);
and U24424 (N_24424,N_22364,N_22275);
nor U24425 (N_24425,N_23543,N_22066);
xnor U24426 (N_24426,N_23099,N_23358);
or U24427 (N_24427,N_23553,N_23438);
nand U24428 (N_24428,N_23119,N_23725);
nor U24429 (N_24429,N_22467,N_23297);
or U24430 (N_24430,N_22999,N_22966);
nor U24431 (N_24431,N_22412,N_23720);
nor U24432 (N_24432,N_22976,N_23267);
nand U24433 (N_24433,N_23072,N_22035);
or U24434 (N_24434,N_22115,N_23711);
xor U24435 (N_24435,N_22952,N_22444);
nor U24436 (N_24436,N_23801,N_22184);
nor U24437 (N_24437,N_22948,N_22594);
nor U24438 (N_24438,N_22868,N_22526);
xnor U24439 (N_24439,N_22829,N_23869);
and U24440 (N_24440,N_23163,N_22918);
or U24441 (N_24441,N_22238,N_22733);
and U24442 (N_24442,N_22779,N_23707);
xnor U24443 (N_24443,N_23341,N_22815);
or U24444 (N_24444,N_23602,N_22407);
nor U24445 (N_24445,N_22464,N_22417);
nand U24446 (N_24446,N_23643,N_22293);
xor U24447 (N_24447,N_22056,N_22030);
nor U24448 (N_24448,N_22331,N_23335);
and U24449 (N_24449,N_22535,N_23599);
nor U24450 (N_24450,N_23398,N_23846);
xor U24451 (N_24451,N_23415,N_23547);
nand U24452 (N_24452,N_23190,N_23142);
and U24453 (N_24453,N_22838,N_22437);
nor U24454 (N_24454,N_23020,N_23695);
xor U24455 (N_24455,N_23486,N_22024);
xor U24456 (N_24456,N_23135,N_23708);
or U24457 (N_24457,N_22236,N_23902);
and U24458 (N_24458,N_23376,N_22852);
or U24459 (N_24459,N_23196,N_22565);
nand U24460 (N_24460,N_23427,N_22689);
or U24461 (N_24461,N_22418,N_23913);
xnor U24462 (N_24462,N_22346,N_23882);
nor U24463 (N_24463,N_22613,N_22162);
nand U24464 (N_24464,N_22710,N_23168);
xnor U24465 (N_24465,N_22496,N_22349);
xor U24466 (N_24466,N_23715,N_22604);
nand U24467 (N_24467,N_22420,N_23824);
nand U24468 (N_24468,N_23521,N_22978);
or U24469 (N_24469,N_22676,N_23107);
or U24470 (N_24470,N_22484,N_22825);
xor U24471 (N_24471,N_22603,N_22427);
nand U24472 (N_24472,N_22212,N_22895);
and U24473 (N_24473,N_23133,N_22986);
or U24474 (N_24474,N_23268,N_22679);
nor U24475 (N_24475,N_22814,N_23687);
xor U24476 (N_24476,N_23611,N_22492);
nor U24477 (N_24477,N_23574,N_22881);
nor U24478 (N_24478,N_22884,N_22794);
or U24479 (N_24479,N_22543,N_22109);
xor U24480 (N_24480,N_22693,N_22481);
nor U24481 (N_24481,N_22124,N_22133);
xor U24482 (N_24482,N_23145,N_23171);
nand U24483 (N_24483,N_23000,N_23974);
and U24484 (N_24484,N_23484,N_23435);
or U24485 (N_24485,N_23069,N_23456);
xor U24486 (N_24486,N_22004,N_22119);
and U24487 (N_24487,N_23588,N_23980);
nor U24488 (N_24488,N_23895,N_22674);
and U24489 (N_24489,N_23191,N_23180);
xnor U24490 (N_24490,N_22061,N_23957);
and U24491 (N_24491,N_23791,N_23811);
xnor U24492 (N_24492,N_22173,N_22167);
nand U24493 (N_24493,N_23871,N_23497);
or U24494 (N_24494,N_23703,N_23326);
nand U24495 (N_24495,N_23140,N_22841);
nor U24496 (N_24496,N_22869,N_22583);
or U24497 (N_24497,N_23017,N_22083);
xnor U24498 (N_24498,N_23242,N_23257);
nor U24499 (N_24499,N_22006,N_22836);
and U24500 (N_24500,N_22324,N_22669);
nand U24501 (N_24501,N_22861,N_22600);
nand U24502 (N_24502,N_22522,N_23874);
or U24503 (N_24503,N_22138,N_23697);
or U24504 (N_24504,N_22909,N_23331);
nand U24505 (N_24505,N_23952,N_22894);
nand U24506 (N_24506,N_23891,N_22630);
and U24507 (N_24507,N_22376,N_23875);
or U24508 (N_24508,N_23187,N_22377);
xnor U24509 (N_24509,N_22717,N_22651);
and U24510 (N_24510,N_22310,N_23139);
and U24511 (N_24511,N_22591,N_23927);
nor U24512 (N_24512,N_23586,N_22698);
or U24513 (N_24513,N_22262,N_22749);
or U24514 (N_24514,N_22752,N_22898);
xnor U24515 (N_24515,N_22218,N_22745);
and U24516 (N_24516,N_22553,N_22734);
and U24517 (N_24517,N_23821,N_23115);
nand U24518 (N_24518,N_22005,N_23483);
nor U24519 (N_24519,N_22152,N_22237);
nor U24520 (N_24520,N_22787,N_22853);
xnor U24521 (N_24521,N_23959,N_23960);
and U24522 (N_24522,N_23756,N_22847);
xnor U24523 (N_24523,N_23560,N_23680);
nor U24524 (N_24524,N_23931,N_23050);
xnor U24525 (N_24525,N_22319,N_22504);
xnor U24526 (N_24526,N_23446,N_22883);
and U24527 (N_24527,N_22049,N_22350);
nor U24528 (N_24528,N_23030,N_22166);
xnor U24529 (N_24529,N_23886,N_22766);
and U24530 (N_24530,N_23378,N_22515);
xor U24531 (N_24531,N_23917,N_23705);
or U24532 (N_24532,N_22260,N_23093);
xor U24533 (N_24533,N_23479,N_22453);
nor U24534 (N_24534,N_22058,N_23254);
or U24535 (N_24535,N_23481,N_22906);
nand U24536 (N_24536,N_22373,N_22209);
xor U24537 (N_24537,N_22944,N_23806);
nor U24538 (N_24538,N_23371,N_22008);
xor U24539 (N_24539,N_22783,N_23999);
nor U24540 (N_24540,N_22239,N_22353);
or U24541 (N_24541,N_22970,N_22019);
or U24542 (N_24542,N_23502,N_23251);
nor U24543 (N_24543,N_22819,N_23919);
nor U24544 (N_24544,N_23905,N_22850);
nor U24545 (N_24545,N_22104,N_22198);
nor U24546 (N_24546,N_23346,N_23394);
and U24547 (N_24547,N_22902,N_22452);
or U24548 (N_24548,N_22286,N_22316);
and U24549 (N_24549,N_23136,N_22557);
or U24550 (N_24550,N_23665,N_22280);
nor U24551 (N_24551,N_22007,N_23730);
xor U24552 (N_24552,N_23768,N_23991);
nor U24553 (N_24553,N_23839,N_22186);
nand U24554 (N_24554,N_23042,N_23159);
or U24555 (N_24555,N_22533,N_23362);
xor U24556 (N_24556,N_23977,N_22118);
and U24557 (N_24557,N_22574,N_23884);
xnor U24558 (N_24558,N_23293,N_23355);
or U24559 (N_24559,N_22051,N_22502);
and U24560 (N_24560,N_23103,N_22131);
nor U24561 (N_24561,N_22920,N_23420);
nor U24562 (N_24562,N_22638,N_23350);
and U24563 (N_24563,N_22087,N_23432);
nand U24564 (N_24564,N_22248,N_23088);
nor U24565 (N_24565,N_23684,N_23889);
nor U24566 (N_24566,N_22003,N_23027);
xnor U24567 (N_24567,N_22479,N_22888);
and U24568 (N_24568,N_22955,N_23280);
nor U24569 (N_24569,N_22937,N_23972);
or U24570 (N_24570,N_22406,N_22106);
xor U24571 (N_24571,N_22154,N_22404);
xor U24572 (N_24572,N_22093,N_22907);
and U24573 (N_24573,N_22491,N_22210);
or U24574 (N_24574,N_23809,N_23609);
and U24575 (N_24575,N_23320,N_22617);
nand U24576 (N_24576,N_22593,N_22021);
nor U24577 (N_24577,N_22232,N_23881);
nand U24578 (N_24578,N_23583,N_23028);
and U24579 (N_24579,N_23877,N_22419);
and U24580 (N_24580,N_22499,N_23111);
or U24581 (N_24581,N_23460,N_23141);
nor U24582 (N_24582,N_22033,N_22910);
xnor U24583 (N_24583,N_22939,N_23598);
and U24584 (N_24584,N_23422,N_22527);
nand U24585 (N_24585,N_23052,N_23383);
or U24586 (N_24586,N_22476,N_22622);
and U24587 (N_24587,N_23039,N_22243);
nor U24588 (N_24588,N_23070,N_23270);
nand U24589 (N_24589,N_23121,N_23828);
nand U24590 (N_24590,N_23120,N_23864);
or U24591 (N_24591,N_23535,N_23271);
or U24592 (N_24592,N_22922,N_22714);
xor U24593 (N_24593,N_22374,N_23964);
or U24594 (N_24594,N_22681,N_22269);
or U24595 (N_24595,N_22163,N_22516);
xor U24596 (N_24596,N_22968,N_22980);
or U24597 (N_24597,N_22750,N_23729);
nor U24598 (N_24598,N_22185,N_23049);
xor U24599 (N_24599,N_23340,N_22043);
or U24600 (N_24600,N_22648,N_22995);
nor U24601 (N_24601,N_23653,N_23569);
xor U24602 (N_24602,N_22438,N_22928);
nand U24603 (N_24603,N_23008,N_23771);
xnor U24604 (N_24604,N_22487,N_23872);
or U24605 (N_24605,N_22632,N_22835);
nor U24606 (N_24606,N_22579,N_22067);
xnor U24607 (N_24607,N_22430,N_23385);
or U24608 (N_24608,N_23012,N_22833);
xor U24609 (N_24609,N_23800,N_22334);
xor U24610 (N_24610,N_23655,N_22737);
and U24611 (N_24611,N_22252,N_23276);
nand U24612 (N_24612,N_23528,N_22892);
nand U24613 (N_24613,N_23177,N_23285);
xor U24614 (N_24614,N_23632,N_23296);
nand U24615 (N_24615,N_22110,N_22400);
nor U24616 (N_24616,N_22169,N_22434);
xnor U24617 (N_24617,N_23563,N_23260);
and U24618 (N_24618,N_22098,N_23018);
and U24619 (N_24619,N_23023,N_22117);
nand U24620 (N_24620,N_23843,N_22530);
xnor U24621 (N_24621,N_23623,N_23934);
xor U24622 (N_24622,N_22288,N_22782);
nor U24623 (N_24623,N_23940,N_23424);
and U24624 (N_24624,N_22337,N_23116);
and U24625 (N_24625,N_22313,N_23166);
nand U24626 (N_24626,N_22401,N_23387);
nand U24627 (N_24627,N_23582,N_22589);
and U24628 (N_24628,N_22245,N_23944);
nor U24629 (N_24629,N_23081,N_23661);
nand U24630 (N_24630,N_23153,N_22634);
nor U24631 (N_24631,N_23789,N_23252);
nor U24632 (N_24632,N_22057,N_23311);
nor U24633 (N_24633,N_23997,N_23491);
nor U24634 (N_24634,N_23124,N_23031);
nand U24635 (N_24635,N_23218,N_22683);
and U24636 (N_24636,N_23265,N_22010);
nor U24637 (N_24637,N_22264,N_23055);
nor U24638 (N_24638,N_22102,N_23172);
xor U24639 (N_24639,N_23739,N_22450);
and U24640 (N_24640,N_23494,N_22712);
nand U24641 (N_24641,N_22211,N_22510);
or U24642 (N_24642,N_22292,N_22413);
nand U24643 (N_24643,N_22973,N_23554);
nor U24644 (N_24644,N_22277,N_23853);
xor U24645 (N_24645,N_22549,N_22837);
nor U24646 (N_24646,N_23671,N_23082);
or U24647 (N_24647,N_23841,N_23179);
nand U24648 (N_24648,N_22637,N_23593);
or U24649 (N_24649,N_22959,N_22842);
nor U24650 (N_24650,N_23489,N_23109);
xor U24651 (N_24651,N_22699,N_23118);
nor U24652 (N_24652,N_23227,N_22389);
and U24653 (N_24653,N_22020,N_23540);
or U24654 (N_24654,N_23208,N_22827);
or U24655 (N_24655,N_22287,N_22084);
and U24656 (N_24656,N_23814,N_23303);
xnor U24657 (N_24657,N_23445,N_22650);
xor U24658 (N_24658,N_23289,N_22742);
nand U24659 (N_24659,N_23328,N_23405);
and U24660 (N_24660,N_23855,N_23955);
xor U24661 (N_24661,N_23967,N_22314);
nand U24662 (N_24662,N_22921,N_23924);
xor U24663 (N_24663,N_23682,N_23503);
nor U24664 (N_24664,N_23401,N_22415);
or U24665 (N_24665,N_23674,N_22773);
and U24666 (N_24666,N_22390,N_23245);
or U24667 (N_24667,N_22675,N_23817);
nand U24668 (N_24668,N_23178,N_23263);
nand U24669 (N_24669,N_23054,N_22677);
and U24670 (N_24670,N_22064,N_23681);
xor U24671 (N_24671,N_22709,N_22871);
or U24672 (N_24672,N_22362,N_22878);
and U24673 (N_24673,N_23451,N_22759);
and U24674 (N_24674,N_22135,N_22887);
xor U24675 (N_24675,N_22723,N_23499);
nor U24676 (N_24676,N_22294,N_23865);
nand U24677 (N_24677,N_22283,N_23897);
nor U24678 (N_24678,N_23330,N_23848);
nor U24679 (N_24679,N_22379,N_23835);
or U24680 (N_24680,N_23466,N_22428);
nor U24681 (N_24681,N_23686,N_22461);
or U24682 (N_24682,N_23148,N_22468);
nor U24683 (N_24683,N_22355,N_22002);
xor U24684 (N_24684,N_23379,N_22072);
or U24685 (N_24685,N_23607,N_23461);
and U24686 (N_24686,N_23010,N_22688);
and U24687 (N_24687,N_23748,N_22105);
or U24688 (N_24688,N_22776,N_23590);
xor U24689 (N_24689,N_22429,N_23763);
or U24690 (N_24690,N_22812,N_23463);
or U24691 (N_24691,N_22284,N_22626);
nand U24692 (N_24692,N_22525,N_22416);
or U24693 (N_24693,N_23277,N_22931);
and U24694 (N_24694,N_23753,N_22643);
and U24695 (N_24695,N_22899,N_22381);
nand U24696 (N_24696,N_22652,N_22691);
or U24697 (N_24697,N_23904,N_23525);
nor U24698 (N_24698,N_22044,N_23314);
xnor U24699 (N_24699,N_23552,N_22788);
nand U24700 (N_24700,N_22806,N_22659);
and U24701 (N_24701,N_23400,N_23825);
or U24702 (N_24702,N_22219,N_22231);
and U24703 (N_24703,N_22426,N_23561);
nand U24704 (N_24704,N_23900,N_22111);
xor U24705 (N_24705,N_23388,N_22865);
nor U24706 (N_24706,N_22457,N_23921);
nor U24707 (N_24707,N_22059,N_23802);
xor U24708 (N_24708,N_22855,N_23165);
or U24709 (N_24709,N_23513,N_22947);
nand U24710 (N_24710,N_22366,N_23818);
nand U24711 (N_24711,N_23518,N_22148);
or U24712 (N_24712,N_23003,N_23805);
nand U24713 (N_24713,N_23290,N_23452);
and U24714 (N_24714,N_23783,N_22075);
or U24715 (N_24715,N_22199,N_23462);
xor U24716 (N_24716,N_23937,N_23198);
or U24717 (N_24717,N_22670,N_23600);
and U24718 (N_24718,N_22592,N_23469);
nor U24719 (N_24719,N_23765,N_22705);
nand U24720 (N_24720,N_23313,N_22791);
and U24721 (N_24721,N_23859,N_23734);
xor U24722 (N_24722,N_23950,N_22726);
xor U24723 (N_24723,N_22380,N_22802);
nor U24724 (N_24724,N_23529,N_23302);
nor U24725 (N_24725,N_22172,N_23235);
nand U24726 (N_24726,N_23641,N_23844);
or U24727 (N_24727,N_23507,N_23075);
nor U24728 (N_24728,N_22857,N_23556);
nand U24729 (N_24729,N_23500,N_22997);
and U24730 (N_24730,N_23936,N_23195);
xnor U24731 (N_24731,N_22826,N_23433);
xor U24732 (N_24732,N_22642,N_23774);
and U24733 (N_24733,N_22409,N_23636);
nand U24734 (N_24734,N_22274,N_22052);
or U24735 (N_24735,N_23657,N_23063);
or U24736 (N_24736,N_23962,N_23530);
nor U24737 (N_24737,N_23876,N_22905);
xnor U24738 (N_24738,N_23614,N_22962);
or U24739 (N_24739,N_22341,N_22880);
or U24740 (N_24740,N_23981,N_22224);
and U24741 (N_24741,N_22711,N_22065);
nor U24742 (N_24742,N_23396,N_23339);
or U24743 (N_24743,N_22249,N_23021);
nor U24744 (N_24744,N_23458,N_23437);
or U24745 (N_24745,N_22465,N_22798);
and U24746 (N_24746,N_22456,N_23305);
and U24747 (N_24747,N_23892,N_23366);
or U24748 (N_24748,N_22251,N_23689);
and U24749 (N_24749,N_23368,N_22270);
or U24750 (N_24750,N_22740,N_22573);
nor U24751 (N_24751,N_22517,N_23193);
nor U24752 (N_24752,N_23373,N_22171);
or U24753 (N_24753,N_22911,N_22153);
or U24754 (N_24754,N_23377,N_22548);
nor U24755 (N_24755,N_23264,N_23080);
nand U24756 (N_24756,N_22137,N_22662);
and U24757 (N_24757,N_23719,N_23353);
xnor U24758 (N_24758,N_23361,N_23079);
xnor U24759 (N_24759,N_22879,N_23514);
or U24760 (N_24760,N_22179,N_22666);
nor U24761 (N_24761,N_23425,N_23544);
xor U24762 (N_24762,N_23721,N_23053);
nor U24763 (N_24763,N_23241,N_22949);
or U24764 (N_24764,N_23996,N_23354);
and U24765 (N_24765,N_22991,N_23635);
or U24766 (N_24766,N_23995,N_23203);
or U24767 (N_24767,N_22195,N_22387);
xor U24768 (N_24768,N_23065,N_22761);
and U24769 (N_24769,N_22181,N_22482);
nand U24770 (N_24770,N_23096,N_23150);
nand U24771 (N_24771,N_22039,N_23928);
nand U24772 (N_24772,N_23442,N_22351);
or U24773 (N_24773,N_22164,N_22225);
and U24774 (N_24774,N_23232,N_23223);
xnor U24775 (N_24775,N_23134,N_22298);
xor U24776 (N_24776,N_23281,N_23029);
nand U24777 (N_24777,N_23259,N_23352);
and U24778 (N_24778,N_23152,N_23201);
or U24779 (N_24779,N_22560,N_23982);
or U24780 (N_24780,N_23624,N_23211);
and U24781 (N_24781,N_22158,N_22234);
xnor U24782 (N_24782,N_23073,N_23870);
or U24783 (N_24783,N_23161,N_22189);
xor U24784 (N_24784,N_23577,N_23349);
and U24785 (N_24785,N_22578,N_23531);
or U24786 (N_24786,N_23978,N_22445);
nor U24787 (N_24787,N_23920,N_23758);
nor U24788 (N_24788,N_23831,N_23319);
xor U24789 (N_24789,N_23679,N_22266);
nor U24790 (N_24790,N_23038,N_22348);
and U24791 (N_24791,N_23472,N_22113);
nand U24792 (N_24792,N_22309,N_22220);
and U24793 (N_24793,N_22903,N_23945);
xnor U24794 (N_24794,N_23584,N_22919);
and U24795 (N_24795,N_22469,N_23879);
xnor U24796 (N_24796,N_22552,N_23450);
and U24797 (N_24797,N_23471,N_23810);
xor U24798 (N_24798,N_22900,N_23085);
or U24799 (N_24799,N_22760,N_22781);
xnor U24800 (N_24800,N_23037,N_22985);
or U24801 (N_24801,N_22757,N_22891);
and U24802 (N_24802,N_23200,N_22508);
nand U24803 (N_24803,N_22764,N_23329);
xnor U24804 (N_24804,N_23156,N_22473);
xor U24805 (N_24805,N_23351,N_23709);
nand U24806 (N_24806,N_22741,N_22831);
nor U24807 (N_24807,N_23678,N_22762);
or U24808 (N_24808,N_22605,N_22990);
nor U24809 (N_24809,N_22214,N_22796);
xnor U24810 (N_24810,N_23915,N_23440);
xor U24811 (N_24811,N_23731,N_23076);
nand U24812 (N_24812,N_22451,N_22770);
or U24813 (N_24813,N_22410,N_22729);
or U24814 (N_24814,N_23058,N_23576);
xnor U24815 (N_24815,N_22914,N_23360);
xnor U24816 (N_24816,N_23488,N_23237);
and U24817 (N_24817,N_22328,N_23359);
xnor U24818 (N_24818,N_23170,N_22368);
xor U24819 (N_24819,N_22635,N_23370);
nand U24820 (N_24820,N_23596,N_23617);
nand U24821 (N_24821,N_22576,N_23637);
xor U24822 (N_24822,N_22490,N_23548);
and U24823 (N_24823,N_23948,N_23918);
nor U24824 (N_24824,N_23087,N_22925);
xnor U24825 (N_24825,N_23858,N_22792);
nand U24826 (N_24826,N_23238,N_23426);
and U24827 (N_24827,N_23550,N_23175);
nand U24828 (N_24828,N_22673,N_22397);
xnor U24829 (N_24829,N_23883,N_22984);
or U24830 (N_24830,N_22336,N_22385);
nor U24831 (N_24831,N_22365,N_22564);
and U24832 (N_24832,N_23537,N_23090);
nor U24833 (N_24833,N_22048,N_22772);
and U24834 (N_24834,N_22132,N_22326);
nor U24835 (N_24835,N_22271,N_22391);
or U24836 (N_24836,N_22192,N_22176);
nand U24837 (N_24837,N_23192,N_23842);
and U24838 (N_24838,N_23421,N_23114);
nand U24839 (N_24839,N_22722,N_22845);
nor U24840 (N_24840,N_23880,N_23480);
xor U24841 (N_24841,N_23249,N_22854);
or U24842 (N_24842,N_23036,N_23204);
nor U24843 (N_24843,N_22926,N_23102);
nand U24844 (N_24844,N_22278,N_23212);
nand U24845 (N_24845,N_23253,N_22306);
xnor U24846 (N_24846,N_23990,N_22071);
or U24847 (N_24847,N_23248,N_22608);
nor U24848 (N_24848,N_22372,N_23033);
nand U24849 (N_24849,N_22615,N_23441);
or U24850 (N_24850,N_22358,N_22816);
or U24851 (N_24851,N_23901,N_22296);
nand U24852 (N_24852,N_23677,N_23393);
or U24853 (N_24853,N_22165,N_22820);
or U24854 (N_24854,N_23194,N_23453);
nor U24855 (N_24855,N_22957,N_22408);
nor U24856 (N_24856,N_22197,N_23778);
or U24857 (N_24857,N_23083,N_22012);
and U24858 (N_24858,N_23300,N_23382);
or U24859 (N_24859,N_22261,N_23717);
and U24860 (N_24860,N_22559,N_22480);
xor U24861 (N_24861,N_23381,N_22821);
xor U24862 (N_24862,N_22474,N_23857);
or U24863 (N_24863,N_22208,N_23701);
nand U24864 (N_24864,N_23169,N_23903);
nand U24865 (N_24865,N_23575,N_23813);
xor U24866 (N_24866,N_23092,N_22369);
nor U24867 (N_24867,N_22323,N_22721);
nand U24868 (N_24868,N_22609,N_22876);
nor U24869 (N_24869,N_22026,N_22360);
and U24870 (N_24870,N_22497,N_23097);
or U24871 (N_24871,N_22000,N_22988);
xnor U24872 (N_24872,N_23035,N_23333);
and U24873 (N_24873,N_23796,N_23587);
xor U24874 (N_24874,N_23676,N_22793);
nor U24875 (N_24875,N_23646,N_23157);
xnor U24876 (N_24876,N_22082,N_22151);
xnor U24877 (N_24877,N_23700,N_22661);
xnor U24878 (N_24878,N_22247,N_22550);
nor U24879 (N_24879,N_22436,N_22846);
nor U24880 (N_24880,N_22134,N_23439);
nand U24881 (N_24881,N_23044,N_23847);
nor U24882 (N_24882,N_22327,N_23444);
or U24883 (N_24883,N_23347,N_22656);
nand U24884 (N_24884,N_23487,N_23334);
or U24885 (N_24885,N_23976,N_22370);
xor U24886 (N_24886,N_23105,N_22912);
xor U24887 (N_24887,N_23213,N_22460);
xor U24888 (N_24888,N_22599,N_22222);
nand U24889 (N_24889,N_22090,N_22916);
xor U24890 (N_24890,N_22611,N_22913);
nor U24891 (N_24891,N_22598,N_23477);
and U24892 (N_24892,N_22136,N_22046);
and U24893 (N_24893,N_23562,N_22811);
xnor U24894 (N_24894,N_22063,N_23173);
xnor U24895 (N_24895,N_23704,N_23011);
nor U24896 (N_24896,N_23001,N_22396);
xnor U24897 (N_24897,N_22697,N_23545);
xnor U24898 (N_24898,N_23523,N_23755);
or U24899 (N_24899,N_23565,N_22471);
nand U24900 (N_24900,N_23798,N_23579);
and U24901 (N_24901,N_22160,N_23849);
and U24902 (N_24902,N_23652,N_22885);
nand U24903 (N_24903,N_22411,N_23043);
and U24904 (N_24904,N_22570,N_23536);
and U24905 (N_24905,N_22425,N_22446);
or U24906 (N_24906,N_22383,N_22120);
or U24907 (N_24907,N_22042,N_23906);
xnor U24908 (N_24908,N_22242,N_22956);
nor U24909 (N_24909,N_23619,N_23047);
xnor U24910 (N_24910,N_22908,N_23113);
or U24911 (N_24911,N_23414,N_22475);
nor U24912 (N_24912,N_23482,N_23310);
or U24913 (N_24913,N_22014,N_22335);
or U24914 (N_24914,N_22701,N_22047);
nand U24915 (N_24915,N_22867,N_22616);
nand U24916 (N_24916,N_22563,N_23411);
xor U24917 (N_24917,N_23231,N_22747);
and U24918 (N_24918,N_22633,N_23559);
and U24919 (N_24919,N_22518,N_23496);
xnor U24920 (N_24920,N_23793,N_22695);
and U24921 (N_24921,N_22168,N_23292);
and U24922 (N_24922,N_23896,N_22958);
and U24923 (N_24923,N_23048,N_23745);
and U24924 (N_24924,N_23317,N_22127);
or U24925 (N_24925,N_22320,N_22692);
nor U24926 (N_24926,N_23733,N_23803);
xnor U24927 (N_24927,N_23605,N_23938);
nor U24928 (N_24928,N_22394,N_22639);
nor U24929 (N_24929,N_23274,N_23322);
nor U24930 (N_24930,N_23851,N_23638);
or U24931 (N_24931,N_23692,N_23057);
and U24932 (N_24932,N_22738,N_22112);
or U24933 (N_24933,N_22904,N_22558);
or U24934 (N_24934,N_22352,N_23866);
xnor U24935 (N_24935,N_22917,N_23723);
nor U24936 (N_24936,N_23644,N_22149);
or U24937 (N_24937,N_22206,N_22466);
xnor U24938 (N_24938,N_22463,N_22672);
or U24939 (N_24939,N_22848,N_22941);
nand U24940 (N_24940,N_23519,N_22216);
nand U24941 (N_24941,N_23391,N_23833);
xnor U24942 (N_24942,N_23061,N_22971);
nand U24943 (N_24943,N_22545,N_23760);
nand U24944 (N_24944,N_23743,N_23275);
or U24945 (N_24945,N_22281,N_22345);
nor U24946 (N_24946,N_23475,N_23509);
or U24947 (N_24947,N_22139,N_22240);
nor U24948 (N_24948,N_22767,N_23863);
xor U24949 (N_24949,N_22629,N_23423);
nor U24950 (N_24950,N_22305,N_22882);
or U24951 (N_24951,N_22646,N_22403);
nor U24952 (N_24952,N_23592,N_22874);
nand U24953 (N_24953,N_23046,N_23823);
nor U24954 (N_24954,N_22311,N_23255);
nand U24955 (N_24955,N_23207,N_22763);
and U24956 (N_24956,N_23747,N_23741);
xnor U24957 (N_24957,N_23005,N_23338);
or U24958 (N_24958,N_22329,N_23221);
and U24959 (N_24959,N_22893,N_22765);
xnor U24960 (N_24960,N_23986,N_23933);
nand U24961 (N_24961,N_22204,N_23222);
xor U24962 (N_24962,N_23794,N_22255);
nor U24963 (N_24963,N_23040,N_23154);
nor U24964 (N_24964,N_23911,N_22395);
or U24965 (N_24965,N_22744,N_23106);
xnor U24966 (N_24966,N_23885,N_23627);
and U24967 (N_24967,N_23585,N_23137);
xnor U24968 (N_24968,N_23827,N_22201);
or U24969 (N_24969,N_22531,N_22227);
xor U24970 (N_24970,N_22780,N_23283);
nor U24971 (N_24971,N_22143,N_22546);
nor U24972 (N_24972,N_22011,N_22263);
and U24973 (N_24973,N_22551,N_22839);
nand U24974 (N_24974,N_22724,N_23327);
or U24975 (N_24975,N_22945,N_23622);
nor U24976 (N_24976,N_22449,N_22983);
nor U24977 (N_24977,N_23449,N_23457);
xor U24978 (N_24978,N_22572,N_23669);
and U24979 (N_24979,N_23973,N_22488);
or U24980 (N_24980,N_23799,N_23004);
or U24981 (N_24981,N_23206,N_22521);
nor U24982 (N_24982,N_22448,N_23301);
xor U24983 (N_24983,N_22923,N_22690);
or U24984 (N_24984,N_22207,N_22746);
nand U24985 (N_24985,N_23826,N_22715);
nor U24986 (N_24986,N_23436,N_22577);
xor U24987 (N_24987,N_23527,N_22150);
xnor U24988 (N_24988,N_23236,N_22472);
xor U24989 (N_24989,N_23908,N_22333);
or U24990 (N_24990,N_23091,N_22285);
or U24991 (N_24991,N_23147,N_22934);
nor U24992 (N_24992,N_23971,N_23958);
or U24993 (N_24993,N_22125,N_22623);
or U24994 (N_24994,N_23965,N_22732);
xor U24995 (N_24995,N_22142,N_22086);
xnor U24996 (N_24996,N_23728,N_23830);
xor U24997 (N_24997,N_22795,N_22751);
or U24998 (N_24998,N_23722,N_23949);
xor U24999 (N_24999,N_23779,N_22040);
nor U25000 (N_25000,N_23655,N_22657);
nor U25001 (N_25001,N_22039,N_22916);
nand U25002 (N_25002,N_22767,N_23317);
and U25003 (N_25003,N_22899,N_22274);
xnor U25004 (N_25004,N_22198,N_22362);
and U25005 (N_25005,N_23778,N_22222);
xor U25006 (N_25006,N_23081,N_23936);
or U25007 (N_25007,N_22391,N_23039);
xnor U25008 (N_25008,N_22427,N_23729);
nand U25009 (N_25009,N_22989,N_22515);
or U25010 (N_25010,N_23945,N_23186);
nor U25011 (N_25011,N_23626,N_22056);
and U25012 (N_25012,N_22677,N_23192);
or U25013 (N_25013,N_22433,N_22458);
nor U25014 (N_25014,N_22402,N_22852);
and U25015 (N_25015,N_22911,N_22808);
or U25016 (N_25016,N_23188,N_22178);
and U25017 (N_25017,N_22714,N_22110);
and U25018 (N_25018,N_23903,N_22484);
xnor U25019 (N_25019,N_23661,N_22446);
nor U25020 (N_25020,N_22880,N_22959);
xor U25021 (N_25021,N_22650,N_22465);
and U25022 (N_25022,N_22380,N_22250);
nand U25023 (N_25023,N_22697,N_22512);
or U25024 (N_25024,N_23641,N_23644);
and U25025 (N_25025,N_23282,N_22571);
nor U25026 (N_25026,N_23427,N_22635);
nor U25027 (N_25027,N_22958,N_23387);
nand U25028 (N_25028,N_22814,N_22338);
nand U25029 (N_25029,N_22443,N_23103);
and U25030 (N_25030,N_22586,N_23469);
nor U25031 (N_25031,N_22406,N_23941);
and U25032 (N_25032,N_23670,N_23982);
or U25033 (N_25033,N_23833,N_22823);
and U25034 (N_25034,N_23056,N_23177);
xnor U25035 (N_25035,N_23850,N_22813);
nand U25036 (N_25036,N_23819,N_22494);
xnor U25037 (N_25037,N_22214,N_22157);
xor U25038 (N_25038,N_23186,N_22530);
nand U25039 (N_25039,N_23358,N_22435);
nor U25040 (N_25040,N_22495,N_22818);
nor U25041 (N_25041,N_22228,N_23970);
nand U25042 (N_25042,N_22038,N_22190);
nand U25043 (N_25043,N_23365,N_22467);
xnor U25044 (N_25044,N_23024,N_22334);
xnor U25045 (N_25045,N_22458,N_22997);
or U25046 (N_25046,N_22021,N_22307);
nor U25047 (N_25047,N_23381,N_23704);
xor U25048 (N_25048,N_22738,N_23095);
or U25049 (N_25049,N_22500,N_22746);
or U25050 (N_25050,N_22362,N_23442);
nand U25051 (N_25051,N_22790,N_23166);
or U25052 (N_25052,N_23627,N_23176);
xnor U25053 (N_25053,N_23815,N_22520);
or U25054 (N_25054,N_23271,N_23641);
xor U25055 (N_25055,N_23526,N_22604);
xnor U25056 (N_25056,N_22726,N_22813);
nand U25057 (N_25057,N_22224,N_23631);
and U25058 (N_25058,N_22219,N_22680);
and U25059 (N_25059,N_22188,N_22169);
nor U25060 (N_25060,N_23753,N_23799);
and U25061 (N_25061,N_23587,N_22700);
or U25062 (N_25062,N_22330,N_23206);
nand U25063 (N_25063,N_23504,N_22599);
nor U25064 (N_25064,N_23823,N_23767);
nand U25065 (N_25065,N_23540,N_22962);
nor U25066 (N_25066,N_22805,N_22588);
xor U25067 (N_25067,N_22068,N_23854);
xor U25068 (N_25068,N_22243,N_22062);
nor U25069 (N_25069,N_22396,N_23718);
nor U25070 (N_25070,N_23371,N_23194);
and U25071 (N_25071,N_23974,N_22790);
xnor U25072 (N_25072,N_23620,N_23473);
nor U25073 (N_25073,N_22998,N_22169);
nand U25074 (N_25074,N_22534,N_22711);
nor U25075 (N_25075,N_23578,N_22998);
xor U25076 (N_25076,N_23276,N_22259);
and U25077 (N_25077,N_22542,N_22971);
or U25078 (N_25078,N_22948,N_23967);
nand U25079 (N_25079,N_23646,N_23516);
or U25080 (N_25080,N_22459,N_22252);
xnor U25081 (N_25081,N_23750,N_23862);
nand U25082 (N_25082,N_22127,N_23810);
nor U25083 (N_25083,N_22525,N_22681);
nor U25084 (N_25084,N_23547,N_23232);
or U25085 (N_25085,N_23284,N_22076);
nor U25086 (N_25086,N_23217,N_22637);
or U25087 (N_25087,N_23040,N_22092);
nand U25088 (N_25088,N_22110,N_22570);
nor U25089 (N_25089,N_23988,N_23173);
and U25090 (N_25090,N_23067,N_23077);
nor U25091 (N_25091,N_22406,N_22263);
or U25092 (N_25092,N_22651,N_22742);
or U25093 (N_25093,N_23654,N_23738);
xnor U25094 (N_25094,N_23568,N_22382);
nor U25095 (N_25095,N_23415,N_22481);
nor U25096 (N_25096,N_22199,N_23845);
nand U25097 (N_25097,N_22909,N_22155);
nor U25098 (N_25098,N_23703,N_23640);
or U25099 (N_25099,N_23038,N_22816);
nand U25100 (N_25100,N_23136,N_23002);
nand U25101 (N_25101,N_23728,N_22215);
xor U25102 (N_25102,N_23466,N_23747);
nand U25103 (N_25103,N_22890,N_22715);
nor U25104 (N_25104,N_22083,N_23716);
xor U25105 (N_25105,N_22586,N_22679);
xnor U25106 (N_25106,N_22739,N_23684);
or U25107 (N_25107,N_23637,N_22035);
or U25108 (N_25108,N_22428,N_23612);
xor U25109 (N_25109,N_22747,N_22179);
and U25110 (N_25110,N_22721,N_23977);
xnor U25111 (N_25111,N_23983,N_22238);
xor U25112 (N_25112,N_23655,N_22168);
and U25113 (N_25113,N_22911,N_23645);
nor U25114 (N_25114,N_22597,N_23364);
or U25115 (N_25115,N_23569,N_23675);
nor U25116 (N_25116,N_22906,N_23622);
nor U25117 (N_25117,N_23892,N_23885);
xor U25118 (N_25118,N_22611,N_23292);
nand U25119 (N_25119,N_22456,N_23494);
nand U25120 (N_25120,N_23874,N_22139);
nor U25121 (N_25121,N_22720,N_23037);
and U25122 (N_25122,N_23678,N_22560);
xnor U25123 (N_25123,N_22770,N_22942);
or U25124 (N_25124,N_23370,N_22819);
nand U25125 (N_25125,N_22327,N_23821);
xor U25126 (N_25126,N_22916,N_22678);
and U25127 (N_25127,N_23100,N_23473);
and U25128 (N_25128,N_22663,N_23063);
or U25129 (N_25129,N_23426,N_23657);
and U25130 (N_25130,N_23855,N_22019);
and U25131 (N_25131,N_23454,N_23297);
xnor U25132 (N_25132,N_23173,N_23047);
nor U25133 (N_25133,N_22722,N_23146);
nand U25134 (N_25134,N_22574,N_23612);
xor U25135 (N_25135,N_23872,N_22792);
and U25136 (N_25136,N_22412,N_22541);
xor U25137 (N_25137,N_22456,N_23119);
and U25138 (N_25138,N_22476,N_23086);
or U25139 (N_25139,N_22457,N_23531);
nand U25140 (N_25140,N_23022,N_23665);
or U25141 (N_25141,N_22753,N_22585);
and U25142 (N_25142,N_22031,N_23612);
or U25143 (N_25143,N_22569,N_23182);
and U25144 (N_25144,N_23586,N_22920);
and U25145 (N_25145,N_22588,N_23594);
or U25146 (N_25146,N_22399,N_22245);
and U25147 (N_25147,N_22508,N_23570);
and U25148 (N_25148,N_22380,N_23493);
or U25149 (N_25149,N_23773,N_23109);
nand U25150 (N_25150,N_23497,N_22145);
xor U25151 (N_25151,N_22902,N_22281);
nor U25152 (N_25152,N_23488,N_22159);
xor U25153 (N_25153,N_22441,N_22611);
nand U25154 (N_25154,N_23475,N_23075);
nand U25155 (N_25155,N_23737,N_23468);
nor U25156 (N_25156,N_23566,N_23857);
xnor U25157 (N_25157,N_23732,N_23202);
and U25158 (N_25158,N_22683,N_23566);
or U25159 (N_25159,N_22143,N_23538);
xor U25160 (N_25160,N_22102,N_22672);
or U25161 (N_25161,N_22914,N_23011);
xor U25162 (N_25162,N_23822,N_22788);
nand U25163 (N_25163,N_23790,N_23802);
and U25164 (N_25164,N_23881,N_22460);
or U25165 (N_25165,N_22996,N_22991);
and U25166 (N_25166,N_23042,N_22161);
and U25167 (N_25167,N_23702,N_22391);
nand U25168 (N_25168,N_23685,N_23831);
or U25169 (N_25169,N_22006,N_23201);
xnor U25170 (N_25170,N_22069,N_23603);
nand U25171 (N_25171,N_23750,N_22617);
or U25172 (N_25172,N_22874,N_22796);
or U25173 (N_25173,N_22009,N_23305);
or U25174 (N_25174,N_22458,N_23977);
or U25175 (N_25175,N_23801,N_23322);
nand U25176 (N_25176,N_23170,N_23394);
or U25177 (N_25177,N_23084,N_23470);
or U25178 (N_25178,N_23756,N_23823);
nand U25179 (N_25179,N_23147,N_22354);
or U25180 (N_25180,N_23021,N_22295);
nor U25181 (N_25181,N_23444,N_23964);
or U25182 (N_25182,N_22811,N_23585);
nor U25183 (N_25183,N_22432,N_22111);
or U25184 (N_25184,N_22785,N_22416);
nor U25185 (N_25185,N_23662,N_23514);
nand U25186 (N_25186,N_22125,N_22106);
xor U25187 (N_25187,N_23772,N_23666);
xnor U25188 (N_25188,N_23757,N_22222);
and U25189 (N_25189,N_22368,N_22420);
xnor U25190 (N_25190,N_23166,N_22275);
nand U25191 (N_25191,N_23172,N_22185);
xnor U25192 (N_25192,N_22991,N_22242);
nand U25193 (N_25193,N_23072,N_22043);
and U25194 (N_25194,N_23220,N_22526);
nand U25195 (N_25195,N_22118,N_22993);
nor U25196 (N_25196,N_23396,N_22252);
nor U25197 (N_25197,N_23759,N_22625);
or U25198 (N_25198,N_22087,N_22220);
and U25199 (N_25199,N_22828,N_22394);
xor U25200 (N_25200,N_23035,N_23541);
nor U25201 (N_25201,N_23917,N_22882);
nor U25202 (N_25202,N_23786,N_23395);
nor U25203 (N_25203,N_23331,N_23598);
nand U25204 (N_25204,N_22845,N_23729);
and U25205 (N_25205,N_23021,N_22864);
nor U25206 (N_25206,N_23747,N_23293);
xor U25207 (N_25207,N_22196,N_23155);
nand U25208 (N_25208,N_22581,N_22420);
or U25209 (N_25209,N_23513,N_23276);
xnor U25210 (N_25210,N_23052,N_22374);
nand U25211 (N_25211,N_23020,N_23146);
xor U25212 (N_25212,N_23181,N_22973);
nor U25213 (N_25213,N_23237,N_22642);
xor U25214 (N_25214,N_23424,N_23328);
xor U25215 (N_25215,N_22559,N_22525);
xnor U25216 (N_25216,N_22966,N_23771);
or U25217 (N_25217,N_22292,N_22076);
nor U25218 (N_25218,N_23077,N_22867);
or U25219 (N_25219,N_23641,N_22377);
and U25220 (N_25220,N_22912,N_23672);
xor U25221 (N_25221,N_22850,N_23166);
nand U25222 (N_25222,N_22650,N_23409);
nand U25223 (N_25223,N_23578,N_22603);
and U25224 (N_25224,N_22186,N_23922);
or U25225 (N_25225,N_23605,N_22317);
nor U25226 (N_25226,N_23661,N_23189);
nor U25227 (N_25227,N_22512,N_22638);
or U25228 (N_25228,N_23889,N_23148);
nor U25229 (N_25229,N_23758,N_23685);
nand U25230 (N_25230,N_22578,N_22778);
nand U25231 (N_25231,N_23167,N_23028);
and U25232 (N_25232,N_22450,N_23452);
and U25233 (N_25233,N_22359,N_22611);
or U25234 (N_25234,N_23531,N_22380);
or U25235 (N_25235,N_22126,N_23337);
xor U25236 (N_25236,N_23157,N_23887);
nand U25237 (N_25237,N_23200,N_23490);
and U25238 (N_25238,N_22840,N_23569);
or U25239 (N_25239,N_23275,N_23198);
nor U25240 (N_25240,N_23055,N_23694);
nor U25241 (N_25241,N_22424,N_23071);
or U25242 (N_25242,N_23437,N_23913);
xnor U25243 (N_25243,N_23926,N_23111);
xor U25244 (N_25244,N_22728,N_23292);
nand U25245 (N_25245,N_22197,N_22069);
or U25246 (N_25246,N_22511,N_22877);
nor U25247 (N_25247,N_23541,N_23997);
or U25248 (N_25248,N_23027,N_22466);
nand U25249 (N_25249,N_22878,N_22820);
and U25250 (N_25250,N_22957,N_23812);
nand U25251 (N_25251,N_23972,N_23244);
xnor U25252 (N_25252,N_22649,N_22958);
and U25253 (N_25253,N_23635,N_22199);
nand U25254 (N_25254,N_22509,N_22900);
or U25255 (N_25255,N_22528,N_23787);
xor U25256 (N_25256,N_22273,N_23299);
and U25257 (N_25257,N_22563,N_22007);
nand U25258 (N_25258,N_23080,N_23034);
xnor U25259 (N_25259,N_22669,N_23570);
or U25260 (N_25260,N_23280,N_23577);
and U25261 (N_25261,N_23049,N_22681);
nor U25262 (N_25262,N_23334,N_22828);
or U25263 (N_25263,N_23472,N_22701);
or U25264 (N_25264,N_22119,N_22562);
and U25265 (N_25265,N_22034,N_22485);
or U25266 (N_25266,N_22004,N_22630);
nand U25267 (N_25267,N_23720,N_22052);
nand U25268 (N_25268,N_22371,N_22875);
and U25269 (N_25269,N_22087,N_22118);
nand U25270 (N_25270,N_23741,N_23340);
or U25271 (N_25271,N_22215,N_23649);
xor U25272 (N_25272,N_23730,N_22756);
nor U25273 (N_25273,N_22320,N_23081);
or U25274 (N_25274,N_23453,N_23312);
and U25275 (N_25275,N_22536,N_23472);
xnor U25276 (N_25276,N_22744,N_23317);
nor U25277 (N_25277,N_23864,N_23316);
nor U25278 (N_25278,N_23654,N_23618);
nor U25279 (N_25279,N_22487,N_22675);
nor U25280 (N_25280,N_22834,N_22183);
xnor U25281 (N_25281,N_23088,N_23011);
or U25282 (N_25282,N_23279,N_22424);
nor U25283 (N_25283,N_22980,N_22234);
nor U25284 (N_25284,N_23787,N_23864);
nor U25285 (N_25285,N_23927,N_22751);
and U25286 (N_25286,N_22771,N_22184);
or U25287 (N_25287,N_23248,N_22746);
and U25288 (N_25288,N_23658,N_22487);
and U25289 (N_25289,N_23708,N_22840);
nor U25290 (N_25290,N_22889,N_23404);
or U25291 (N_25291,N_22819,N_23460);
xnor U25292 (N_25292,N_22173,N_23267);
xnor U25293 (N_25293,N_23430,N_22738);
xnor U25294 (N_25294,N_22907,N_23823);
and U25295 (N_25295,N_22744,N_22828);
xor U25296 (N_25296,N_22647,N_23462);
nor U25297 (N_25297,N_22934,N_22448);
xnor U25298 (N_25298,N_23273,N_23144);
nor U25299 (N_25299,N_22845,N_23499);
xor U25300 (N_25300,N_22650,N_23482);
nor U25301 (N_25301,N_23096,N_23291);
or U25302 (N_25302,N_22912,N_22724);
nor U25303 (N_25303,N_23181,N_22472);
and U25304 (N_25304,N_22429,N_23442);
and U25305 (N_25305,N_22888,N_23100);
nand U25306 (N_25306,N_22517,N_22816);
nor U25307 (N_25307,N_22608,N_22243);
xor U25308 (N_25308,N_22991,N_23041);
nand U25309 (N_25309,N_22734,N_23070);
and U25310 (N_25310,N_23943,N_23536);
nor U25311 (N_25311,N_22331,N_22288);
xnor U25312 (N_25312,N_23941,N_23387);
nand U25313 (N_25313,N_23373,N_22135);
xor U25314 (N_25314,N_23820,N_22494);
xor U25315 (N_25315,N_22313,N_22440);
xnor U25316 (N_25316,N_22550,N_22621);
nor U25317 (N_25317,N_22633,N_22981);
xor U25318 (N_25318,N_22316,N_23977);
nor U25319 (N_25319,N_22673,N_23268);
nand U25320 (N_25320,N_23296,N_22784);
nand U25321 (N_25321,N_22740,N_23342);
xor U25322 (N_25322,N_22880,N_22217);
and U25323 (N_25323,N_23339,N_22311);
and U25324 (N_25324,N_22695,N_23636);
xor U25325 (N_25325,N_22229,N_22310);
or U25326 (N_25326,N_23639,N_22581);
and U25327 (N_25327,N_23366,N_22204);
nor U25328 (N_25328,N_23460,N_22508);
nor U25329 (N_25329,N_23931,N_23553);
and U25330 (N_25330,N_22105,N_23773);
xor U25331 (N_25331,N_22029,N_22117);
xnor U25332 (N_25332,N_22546,N_23731);
and U25333 (N_25333,N_22493,N_23759);
or U25334 (N_25334,N_22391,N_22317);
nor U25335 (N_25335,N_22883,N_22544);
or U25336 (N_25336,N_23927,N_23403);
xnor U25337 (N_25337,N_23966,N_22528);
nand U25338 (N_25338,N_23363,N_23780);
xnor U25339 (N_25339,N_23623,N_23969);
nand U25340 (N_25340,N_23354,N_23307);
nand U25341 (N_25341,N_22617,N_22521);
nand U25342 (N_25342,N_23044,N_23378);
or U25343 (N_25343,N_22269,N_22977);
and U25344 (N_25344,N_22619,N_22164);
nor U25345 (N_25345,N_23198,N_23758);
nor U25346 (N_25346,N_23952,N_23128);
nor U25347 (N_25347,N_22245,N_22417);
and U25348 (N_25348,N_23499,N_23970);
and U25349 (N_25349,N_23444,N_22953);
xor U25350 (N_25350,N_23706,N_22132);
xnor U25351 (N_25351,N_22889,N_22281);
and U25352 (N_25352,N_23383,N_22170);
and U25353 (N_25353,N_22034,N_23295);
xnor U25354 (N_25354,N_22069,N_22809);
and U25355 (N_25355,N_23163,N_23075);
or U25356 (N_25356,N_22635,N_23269);
xnor U25357 (N_25357,N_23428,N_22944);
xor U25358 (N_25358,N_23574,N_22534);
xor U25359 (N_25359,N_22771,N_22933);
nand U25360 (N_25360,N_23972,N_22452);
xnor U25361 (N_25361,N_23836,N_22245);
xnor U25362 (N_25362,N_22491,N_23314);
and U25363 (N_25363,N_23304,N_22606);
or U25364 (N_25364,N_23490,N_22677);
xnor U25365 (N_25365,N_22148,N_23997);
nand U25366 (N_25366,N_22224,N_23950);
and U25367 (N_25367,N_22257,N_23400);
and U25368 (N_25368,N_23168,N_22093);
nor U25369 (N_25369,N_23909,N_22730);
and U25370 (N_25370,N_22237,N_23108);
nor U25371 (N_25371,N_23057,N_22036);
nor U25372 (N_25372,N_23291,N_23172);
xnor U25373 (N_25373,N_22825,N_22434);
nand U25374 (N_25374,N_23877,N_23390);
and U25375 (N_25375,N_23705,N_22217);
nand U25376 (N_25376,N_23833,N_23537);
and U25377 (N_25377,N_23076,N_22096);
nand U25378 (N_25378,N_23695,N_22925);
and U25379 (N_25379,N_23037,N_22503);
and U25380 (N_25380,N_22810,N_22843);
or U25381 (N_25381,N_23290,N_23100);
or U25382 (N_25382,N_22340,N_23242);
and U25383 (N_25383,N_22921,N_23105);
nor U25384 (N_25384,N_23176,N_23204);
nor U25385 (N_25385,N_22923,N_23440);
nor U25386 (N_25386,N_23627,N_23927);
or U25387 (N_25387,N_22442,N_23144);
nor U25388 (N_25388,N_23475,N_23718);
or U25389 (N_25389,N_23443,N_22416);
and U25390 (N_25390,N_22110,N_22072);
xnor U25391 (N_25391,N_23895,N_22344);
or U25392 (N_25392,N_22337,N_22396);
or U25393 (N_25393,N_22236,N_23925);
nor U25394 (N_25394,N_22473,N_23315);
and U25395 (N_25395,N_23288,N_23952);
or U25396 (N_25396,N_23384,N_23822);
xnor U25397 (N_25397,N_22772,N_23531);
and U25398 (N_25398,N_22016,N_22543);
xor U25399 (N_25399,N_23609,N_22125);
and U25400 (N_25400,N_23640,N_22905);
xor U25401 (N_25401,N_22453,N_22242);
nand U25402 (N_25402,N_22287,N_23465);
nand U25403 (N_25403,N_23128,N_22137);
nor U25404 (N_25404,N_23779,N_23307);
or U25405 (N_25405,N_22402,N_22689);
and U25406 (N_25406,N_23084,N_22610);
or U25407 (N_25407,N_23501,N_23381);
xnor U25408 (N_25408,N_22491,N_22137);
xor U25409 (N_25409,N_23322,N_22104);
nand U25410 (N_25410,N_22914,N_22151);
nor U25411 (N_25411,N_23676,N_23263);
nand U25412 (N_25412,N_22676,N_22483);
nand U25413 (N_25413,N_22676,N_23593);
xor U25414 (N_25414,N_22303,N_22780);
nor U25415 (N_25415,N_23318,N_22186);
and U25416 (N_25416,N_23435,N_23261);
and U25417 (N_25417,N_22461,N_23913);
and U25418 (N_25418,N_23061,N_23547);
xnor U25419 (N_25419,N_23111,N_22091);
nand U25420 (N_25420,N_23938,N_23368);
nor U25421 (N_25421,N_23275,N_22559);
and U25422 (N_25422,N_22354,N_23334);
and U25423 (N_25423,N_22149,N_22155);
nand U25424 (N_25424,N_23019,N_22018);
nand U25425 (N_25425,N_22436,N_23706);
nor U25426 (N_25426,N_22945,N_22506);
and U25427 (N_25427,N_23085,N_22337);
and U25428 (N_25428,N_22352,N_23162);
nand U25429 (N_25429,N_23702,N_22458);
nor U25430 (N_25430,N_23074,N_23295);
xnor U25431 (N_25431,N_22543,N_23765);
xnor U25432 (N_25432,N_23906,N_22729);
xor U25433 (N_25433,N_22449,N_23093);
nor U25434 (N_25434,N_23870,N_22816);
or U25435 (N_25435,N_23681,N_23522);
and U25436 (N_25436,N_23501,N_22728);
nor U25437 (N_25437,N_22372,N_23759);
nor U25438 (N_25438,N_23644,N_23104);
nand U25439 (N_25439,N_23609,N_23089);
nand U25440 (N_25440,N_22753,N_23379);
or U25441 (N_25441,N_22067,N_23015);
and U25442 (N_25442,N_22897,N_23386);
and U25443 (N_25443,N_23595,N_23200);
or U25444 (N_25444,N_22478,N_22796);
nand U25445 (N_25445,N_22432,N_22565);
and U25446 (N_25446,N_22947,N_22367);
nor U25447 (N_25447,N_22820,N_23037);
xnor U25448 (N_25448,N_22595,N_22333);
and U25449 (N_25449,N_22849,N_22577);
nand U25450 (N_25450,N_22448,N_22095);
nor U25451 (N_25451,N_23166,N_23884);
xor U25452 (N_25452,N_23139,N_23445);
and U25453 (N_25453,N_22169,N_23173);
nand U25454 (N_25454,N_23244,N_23613);
xor U25455 (N_25455,N_22552,N_23000);
xnor U25456 (N_25456,N_23838,N_23804);
and U25457 (N_25457,N_23945,N_22815);
and U25458 (N_25458,N_22727,N_22308);
nor U25459 (N_25459,N_23881,N_23558);
nand U25460 (N_25460,N_22896,N_23413);
xor U25461 (N_25461,N_23044,N_22194);
xnor U25462 (N_25462,N_22616,N_22203);
or U25463 (N_25463,N_22519,N_23650);
and U25464 (N_25464,N_23906,N_23070);
xnor U25465 (N_25465,N_22052,N_22252);
nand U25466 (N_25466,N_23066,N_23504);
xor U25467 (N_25467,N_22444,N_23283);
xor U25468 (N_25468,N_22270,N_22201);
xnor U25469 (N_25469,N_22568,N_23959);
xor U25470 (N_25470,N_23135,N_22553);
nor U25471 (N_25471,N_22126,N_22475);
xor U25472 (N_25472,N_23218,N_22809);
xnor U25473 (N_25473,N_23746,N_22264);
nand U25474 (N_25474,N_23369,N_23843);
nand U25475 (N_25475,N_22883,N_23955);
and U25476 (N_25476,N_23581,N_23471);
nand U25477 (N_25477,N_23986,N_22990);
xnor U25478 (N_25478,N_23208,N_23032);
or U25479 (N_25479,N_23677,N_22173);
xor U25480 (N_25480,N_23366,N_23963);
nor U25481 (N_25481,N_22940,N_23568);
nand U25482 (N_25482,N_23105,N_23913);
xor U25483 (N_25483,N_22395,N_22023);
xor U25484 (N_25484,N_22832,N_22308);
nand U25485 (N_25485,N_22911,N_22497);
and U25486 (N_25486,N_22980,N_22055);
nand U25487 (N_25487,N_23022,N_22379);
nand U25488 (N_25488,N_23316,N_23615);
xor U25489 (N_25489,N_23047,N_23172);
and U25490 (N_25490,N_23223,N_23401);
or U25491 (N_25491,N_22767,N_22394);
nand U25492 (N_25492,N_22492,N_23610);
nand U25493 (N_25493,N_23605,N_22785);
and U25494 (N_25494,N_23461,N_22276);
nand U25495 (N_25495,N_22479,N_22315);
xnor U25496 (N_25496,N_22054,N_23085);
nand U25497 (N_25497,N_23863,N_23109);
and U25498 (N_25498,N_23527,N_23297);
xor U25499 (N_25499,N_22795,N_23095);
xor U25500 (N_25500,N_22539,N_22923);
xor U25501 (N_25501,N_22322,N_23760);
nand U25502 (N_25502,N_22066,N_22590);
nor U25503 (N_25503,N_23441,N_23518);
or U25504 (N_25504,N_22567,N_23780);
and U25505 (N_25505,N_22141,N_22969);
nand U25506 (N_25506,N_22763,N_23495);
and U25507 (N_25507,N_22507,N_22478);
nand U25508 (N_25508,N_22476,N_22483);
nand U25509 (N_25509,N_22058,N_22610);
nor U25510 (N_25510,N_23733,N_23945);
and U25511 (N_25511,N_23349,N_22776);
and U25512 (N_25512,N_22940,N_23671);
or U25513 (N_25513,N_22656,N_22437);
nor U25514 (N_25514,N_22148,N_22138);
and U25515 (N_25515,N_22022,N_23812);
nand U25516 (N_25516,N_23642,N_22596);
nand U25517 (N_25517,N_23489,N_22698);
nand U25518 (N_25518,N_23192,N_23026);
nor U25519 (N_25519,N_22029,N_23827);
xnor U25520 (N_25520,N_23863,N_23592);
nand U25521 (N_25521,N_22359,N_23639);
nand U25522 (N_25522,N_23463,N_22373);
nand U25523 (N_25523,N_23670,N_23836);
nand U25524 (N_25524,N_23179,N_22656);
nand U25525 (N_25525,N_22917,N_22084);
or U25526 (N_25526,N_23929,N_22149);
nand U25527 (N_25527,N_22034,N_22893);
nand U25528 (N_25528,N_22020,N_23648);
nor U25529 (N_25529,N_22890,N_22926);
or U25530 (N_25530,N_23004,N_23410);
or U25531 (N_25531,N_22127,N_22401);
nor U25532 (N_25532,N_22519,N_23161);
xor U25533 (N_25533,N_22596,N_22261);
xnor U25534 (N_25534,N_22126,N_23693);
xnor U25535 (N_25535,N_23575,N_22604);
xnor U25536 (N_25536,N_23438,N_23183);
and U25537 (N_25537,N_23364,N_23733);
nor U25538 (N_25538,N_22873,N_22060);
or U25539 (N_25539,N_22174,N_23371);
xor U25540 (N_25540,N_22099,N_23843);
nor U25541 (N_25541,N_22271,N_22689);
xnor U25542 (N_25542,N_23695,N_23573);
nor U25543 (N_25543,N_22685,N_23776);
xnor U25544 (N_25544,N_22503,N_23593);
xnor U25545 (N_25545,N_22386,N_22101);
xnor U25546 (N_25546,N_22508,N_23630);
xor U25547 (N_25547,N_22830,N_23324);
or U25548 (N_25548,N_22117,N_22086);
nor U25549 (N_25549,N_22915,N_22109);
nand U25550 (N_25550,N_22562,N_23004);
xnor U25551 (N_25551,N_22116,N_22527);
nand U25552 (N_25552,N_22441,N_23768);
nand U25553 (N_25553,N_22468,N_22766);
xor U25554 (N_25554,N_22658,N_22510);
or U25555 (N_25555,N_22617,N_22891);
nor U25556 (N_25556,N_23738,N_23963);
or U25557 (N_25557,N_22750,N_23332);
xor U25558 (N_25558,N_22184,N_23820);
or U25559 (N_25559,N_22593,N_22923);
nand U25560 (N_25560,N_22912,N_22893);
nor U25561 (N_25561,N_23866,N_22460);
xnor U25562 (N_25562,N_22076,N_23138);
nand U25563 (N_25563,N_23645,N_22338);
and U25564 (N_25564,N_22575,N_22831);
xnor U25565 (N_25565,N_23306,N_23666);
and U25566 (N_25566,N_23313,N_22271);
nand U25567 (N_25567,N_23576,N_22228);
xnor U25568 (N_25568,N_23298,N_23484);
nand U25569 (N_25569,N_22712,N_23443);
nand U25570 (N_25570,N_22945,N_22332);
xor U25571 (N_25571,N_22560,N_22687);
xnor U25572 (N_25572,N_22059,N_23759);
or U25573 (N_25573,N_22007,N_22976);
nor U25574 (N_25574,N_22526,N_23355);
nand U25575 (N_25575,N_22211,N_23677);
and U25576 (N_25576,N_23972,N_22159);
nand U25577 (N_25577,N_23894,N_22750);
xor U25578 (N_25578,N_23968,N_22227);
and U25579 (N_25579,N_22643,N_23085);
xor U25580 (N_25580,N_22683,N_22761);
or U25581 (N_25581,N_22945,N_23727);
nor U25582 (N_25582,N_22907,N_23915);
and U25583 (N_25583,N_23901,N_22451);
nor U25584 (N_25584,N_23052,N_22376);
or U25585 (N_25585,N_23606,N_23834);
or U25586 (N_25586,N_23964,N_22893);
nor U25587 (N_25587,N_23300,N_23848);
xor U25588 (N_25588,N_23945,N_22239);
and U25589 (N_25589,N_22505,N_23508);
or U25590 (N_25590,N_23789,N_22717);
and U25591 (N_25591,N_23307,N_22221);
nand U25592 (N_25592,N_23905,N_23103);
and U25593 (N_25593,N_22860,N_22591);
nor U25594 (N_25594,N_22369,N_23104);
or U25595 (N_25595,N_23927,N_23573);
nor U25596 (N_25596,N_22923,N_23030);
nand U25597 (N_25597,N_22953,N_23083);
and U25598 (N_25598,N_23218,N_22497);
nor U25599 (N_25599,N_22392,N_22928);
nand U25600 (N_25600,N_22755,N_22911);
nand U25601 (N_25601,N_23257,N_22262);
and U25602 (N_25602,N_23292,N_22889);
xnor U25603 (N_25603,N_23220,N_22956);
or U25604 (N_25604,N_23957,N_23886);
nand U25605 (N_25605,N_23358,N_23691);
and U25606 (N_25606,N_23886,N_23531);
or U25607 (N_25607,N_22463,N_22460);
nor U25608 (N_25608,N_22763,N_22723);
xnor U25609 (N_25609,N_22931,N_23409);
and U25610 (N_25610,N_22443,N_22600);
and U25611 (N_25611,N_22080,N_22248);
xor U25612 (N_25612,N_23952,N_23851);
nor U25613 (N_25613,N_22764,N_23165);
or U25614 (N_25614,N_23730,N_22090);
nor U25615 (N_25615,N_22830,N_23637);
xor U25616 (N_25616,N_23594,N_23408);
nor U25617 (N_25617,N_23981,N_22564);
xor U25618 (N_25618,N_23728,N_22093);
nor U25619 (N_25619,N_23381,N_22694);
and U25620 (N_25620,N_23933,N_23826);
nand U25621 (N_25621,N_23605,N_22732);
or U25622 (N_25622,N_23768,N_22433);
and U25623 (N_25623,N_22249,N_23987);
or U25624 (N_25624,N_22592,N_23657);
nand U25625 (N_25625,N_23614,N_23452);
or U25626 (N_25626,N_22653,N_22028);
and U25627 (N_25627,N_22821,N_22333);
nor U25628 (N_25628,N_23974,N_23882);
and U25629 (N_25629,N_22989,N_23546);
xor U25630 (N_25630,N_22913,N_22401);
and U25631 (N_25631,N_23619,N_22311);
and U25632 (N_25632,N_23738,N_23523);
nand U25633 (N_25633,N_23634,N_23511);
xor U25634 (N_25634,N_22486,N_23680);
and U25635 (N_25635,N_23928,N_22325);
and U25636 (N_25636,N_22596,N_23235);
nor U25637 (N_25637,N_23966,N_22629);
nand U25638 (N_25638,N_22142,N_23889);
and U25639 (N_25639,N_23417,N_23551);
or U25640 (N_25640,N_23486,N_22580);
nand U25641 (N_25641,N_23558,N_22960);
nor U25642 (N_25642,N_22390,N_23861);
nand U25643 (N_25643,N_22780,N_23414);
and U25644 (N_25644,N_22431,N_23615);
or U25645 (N_25645,N_23020,N_22358);
nand U25646 (N_25646,N_22947,N_23602);
nand U25647 (N_25647,N_22136,N_23574);
or U25648 (N_25648,N_23172,N_23763);
nor U25649 (N_25649,N_23798,N_22338);
nor U25650 (N_25650,N_22959,N_22549);
xnor U25651 (N_25651,N_23970,N_22188);
nor U25652 (N_25652,N_23497,N_22787);
nor U25653 (N_25653,N_23170,N_22758);
xnor U25654 (N_25654,N_23989,N_22706);
xor U25655 (N_25655,N_22617,N_23461);
nand U25656 (N_25656,N_23818,N_22549);
or U25657 (N_25657,N_23181,N_23515);
and U25658 (N_25658,N_23022,N_23967);
or U25659 (N_25659,N_23773,N_23907);
or U25660 (N_25660,N_23120,N_22520);
nand U25661 (N_25661,N_23999,N_23563);
nand U25662 (N_25662,N_23771,N_22710);
and U25663 (N_25663,N_22018,N_22084);
nand U25664 (N_25664,N_22159,N_23255);
nand U25665 (N_25665,N_23611,N_22797);
nand U25666 (N_25666,N_22896,N_22085);
or U25667 (N_25667,N_22634,N_22225);
nand U25668 (N_25668,N_22312,N_22495);
and U25669 (N_25669,N_22132,N_22089);
or U25670 (N_25670,N_22329,N_23956);
nand U25671 (N_25671,N_22562,N_23559);
nor U25672 (N_25672,N_22630,N_23631);
nor U25673 (N_25673,N_22388,N_23245);
xor U25674 (N_25674,N_23129,N_23445);
and U25675 (N_25675,N_22592,N_22799);
and U25676 (N_25676,N_23889,N_22084);
nand U25677 (N_25677,N_22376,N_22516);
or U25678 (N_25678,N_23916,N_23109);
nor U25679 (N_25679,N_22452,N_22167);
xor U25680 (N_25680,N_22338,N_23272);
nand U25681 (N_25681,N_22649,N_23362);
xor U25682 (N_25682,N_23756,N_22851);
nor U25683 (N_25683,N_22350,N_22769);
xor U25684 (N_25684,N_23533,N_22838);
and U25685 (N_25685,N_23303,N_23638);
and U25686 (N_25686,N_23902,N_23172);
and U25687 (N_25687,N_22126,N_23074);
and U25688 (N_25688,N_23037,N_22277);
or U25689 (N_25689,N_22303,N_22872);
and U25690 (N_25690,N_23173,N_22720);
nor U25691 (N_25691,N_23941,N_22685);
or U25692 (N_25692,N_23269,N_22526);
or U25693 (N_25693,N_23485,N_23845);
and U25694 (N_25694,N_22957,N_22313);
or U25695 (N_25695,N_23586,N_23061);
xnor U25696 (N_25696,N_23469,N_23968);
nand U25697 (N_25697,N_23490,N_22457);
or U25698 (N_25698,N_22272,N_23016);
and U25699 (N_25699,N_23123,N_22246);
or U25700 (N_25700,N_23231,N_22453);
and U25701 (N_25701,N_23482,N_23864);
and U25702 (N_25702,N_23406,N_22712);
nand U25703 (N_25703,N_23367,N_22681);
and U25704 (N_25704,N_23443,N_23413);
nor U25705 (N_25705,N_23549,N_22878);
nand U25706 (N_25706,N_22568,N_22651);
and U25707 (N_25707,N_22007,N_22613);
and U25708 (N_25708,N_22491,N_22725);
and U25709 (N_25709,N_22062,N_23984);
xnor U25710 (N_25710,N_22917,N_23757);
xnor U25711 (N_25711,N_23505,N_22924);
or U25712 (N_25712,N_23959,N_23048);
xnor U25713 (N_25713,N_23656,N_23016);
xor U25714 (N_25714,N_22315,N_22126);
nor U25715 (N_25715,N_22962,N_22369);
nor U25716 (N_25716,N_23871,N_23406);
nand U25717 (N_25717,N_23739,N_23884);
xor U25718 (N_25718,N_22035,N_23867);
xnor U25719 (N_25719,N_22724,N_23761);
and U25720 (N_25720,N_23523,N_23031);
nor U25721 (N_25721,N_22027,N_22659);
or U25722 (N_25722,N_22499,N_22955);
nand U25723 (N_25723,N_23876,N_23216);
nand U25724 (N_25724,N_22435,N_22240);
nor U25725 (N_25725,N_23297,N_22369);
xnor U25726 (N_25726,N_22385,N_23999);
and U25727 (N_25727,N_23836,N_22289);
nand U25728 (N_25728,N_23101,N_23442);
xnor U25729 (N_25729,N_22875,N_22176);
nor U25730 (N_25730,N_23743,N_22965);
or U25731 (N_25731,N_22052,N_23474);
xor U25732 (N_25732,N_22235,N_23062);
nor U25733 (N_25733,N_22518,N_23551);
xor U25734 (N_25734,N_23735,N_22711);
nand U25735 (N_25735,N_23151,N_22076);
or U25736 (N_25736,N_23200,N_23162);
nand U25737 (N_25737,N_22062,N_23494);
xor U25738 (N_25738,N_23307,N_22170);
nor U25739 (N_25739,N_23629,N_23155);
nand U25740 (N_25740,N_22498,N_22633);
or U25741 (N_25741,N_23846,N_23829);
or U25742 (N_25742,N_22958,N_22136);
and U25743 (N_25743,N_22189,N_23922);
nand U25744 (N_25744,N_23800,N_23921);
or U25745 (N_25745,N_23518,N_22056);
nor U25746 (N_25746,N_22635,N_23254);
xnor U25747 (N_25747,N_23946,N_23645);
or U25748 (N_25748,N_23526,N_22140);
and U25749 (N_25749,N_23697,N_22376);
xnor U25750 (N_25750,N_22029,N_22518);
nand U25751 (N_25751,N_22792,N_23654);
and U25752 (N_25752,N_23081,N_23193);
nand U25753 (N_25753,N_23164,N_23874);
nand U25754 (N_25754,N_22205,N_23593);
and U25755 (N_25755,N_22990,N_22830);
and U25756 (N_25756,N_23841,N_23646);
and U25757 (N_25757,N_23215,N_23109);
nand U25758 (N_25758,N_22287,N_22754);
nor U25759 (N_25759,N_23490,N_23267);
nor U25760 (N_25760,N_22376,N_22416);
xor U25761 (N_25761,N_23308,N_23692);
nand U25762 (N_25762,N_22715,N_23075);
nor U25763 (N_25763,N_23876,N_23371);
nand U25764 (N_25764,N_23016,N_23114);
or U25765 (N_25765,N_22764,N_22817);
nor U25766 (N_25766,N_22960,N_22888);
or U25767 (N_25767,N_23929,N_23229);
nor U25768 (N_25768,N_23927,N_23272);
nor U25769 (N_25769,N_23850,N_23220);
nand U25770 (N_25770,N_22211,N_23963);
or U25771 (N_25771,N_22139,N_22120);
xor U25772 (N_25772,N_22490,N_22826);
nor U25773 (N_25773,N_23094,N_23604);
xnor U25774 (N_25774,N_22180,N_22189);
nand U25775 (N_25775,N_23089,N_23383);
and U25776 (N_25776,N_22186,N_22707);
and U25777 (N_25777,N_22352,N_23619);
or U25778 (N_25778,N_23524,N_22925);
and U25779 (N_25779,N_22625,N_22873);
nand U25780 (N_25780,N_22401,N_22346);
or U25781 (N_25781,N_22826,N_23850);
nor U25782 (N_25782,N_23389,N_22154);
or U25783 (N_25783,N_22301,N_22605);
nand U25784 (N_25784,N_23450,N_22921);
and U25785 (N_25785,N_23134,N_22777);
or U25786 (N_25786,N_23587,N_22889);
or U25787 (N_25787,N_22064,N_23823);
nand U25788 (N_25788,N_23959,N_22615);
xor U25789 (N_25789,N_23828,N_22556);
nand U25790 (N_25790,N_23000,N_22957);
or U25791 (N_25791,N_23972,N_23393);
or U25792 (N_25792,N_22645,N_22154);
xor U25793 (N_25793,N_23414,N_23226);
and U25794 (N_25794,N_23003,N_23928);
and U25795 (N_25795,N_22048,N_23061);
and U25796 (N_25796,N_22373,N_22559);
and U25797 (N_25797,N_22768,N_23509);
nor U25798 (N_25798,N_23378,N_23035);
nor U25799 (N_25799,N_22636,N_22956);
nand U25800 (N_25800,N_22426,N_23032);
and U25801 (N_25801,N_22827,N_23751);
xnor U25802 (N_25802,N_23738,N_23257);
nand U25803 (N_25803,N_22993,N_23881);
nor U25804 (N_25804,N_22248,N_22296);
xor U25805 (N_25805,N_22772,N_22653);
xor U25806 (N_25806,N_23199,N_22322);
nand U25807 (N_25807,N_22185,N_22951);
nand U25808 (N_25808,N_22897,N_23762);
xnor U25809 (N_25809,N_23360,N_22361);
and U25810 (N_25810,N_23836,N_23869);
xnor U25811 (N_25811,N_23878,N_23799);
and U25812 (N_25812,N_22628,N_23879);
and U25813 (N_25813,N_23007,N_23260);
xnor U25814 (N_25814,N_23951,N_22317);
and U25815 (N_25815,N_22508,N_22481);
nor U25816 (N_25816,N_22399,N_22147);
nor U25817 (N_25817,N_23412,N_22160);
or U25818 (N_25818,N_23031,N_22205);
nand U25819 (N_25819,N_23197,N_23911);
nor U25820 (N_25820,N_22124,N_22617);
xor U25821 (N_25821,N_23263,N_23297);
xnor U25822 (N_25822,N_22111,N_22118);
nor U25823 (N_25823,N_22127,N_22599);
and U25824 (N_25824,N_23204,N_22227);
nor U25825 (N_25825,N_22469,N_23260);
nand U25826 (N_25826,N_23102,N_23921);
and U25827 (N_25827,N_22123,N_22438);
and U25828 (N_25828,N_23421,N_23711);
or U25829 (N_25829,N_23266,N_22751);
nor U25830 (N_25830,N_23660,N_22443);
and U25831 (N_25831,N_22577,N_22034);
nand U25832 (N_25832,N_23018,N_23463);
or U25833 (N_25833,N_23435,N_22161);
or U25834 (N_25834,N_22563,N_23941);
and U25835 (N_25835,N_22180,N_23683);
or U25836 (N_25836,N_22432,N_23031);
xor U25837 (N_25837,N_23325,N_23431);
xor U25838 (N_25838,N_22377,N_23830);
nand U25839 (N_25839,N_22019,N_23292);
and U25840 (N_25840,N_22428,N_22190);
nor U25841 (N_25841,N_23389,N_23567);
nand U25842 (N_25842,N_22517,N_22143);
nand U25843 (N_25843,N_23464,N_22338);
xor U25844 (N_25844,N_22369,N_22254);
nand U25845 (N_25845,N_22186,N_23513);
nor U25846 (N_25846,N_22111,N_22806);
and U25847 (N_25847,N_22370,N_22932);
and U25848 (N_25848,N_22248,N_23355);
nand U25849 (N_25849,N_22175,N_22942);
nand U25850 (N_25850,N_23811,N_22512);
nand U25851 (N_25851,N_23372,N_23251);
and U25852 (N_25852,N_22661,N_22396);
nor U25853 (N_25853,N_23316,N_22399);
nor U25854 (N_25854,N_22329,N_22363);
nor U25855 (N_25855,N_22891,N_22647);
nor U25856 (N_25856,N_23087,N_23570);
xnor U25857 (N_25857,N_22536,N_22135);
nor U25858 (N_25858,N_23669,N_23381);
xor U25859 (N_25859,N_23663,N_23969);
and U25860 (N_25860,N_22507,N_23688);
or U25861 (N_25861,N_23400,N_22139);
and U25862 (N_25862,N_22202,N_23405);
nor U25863 (N_25863,N_23821,N_22663);
nor U25864 (N_25864,N_22742,N_22718);
and U25865 (N_25865,N_22562,N_22280);
or U25866 (N_25866,N_23685,N_22706);
nand U25867 (N_25867,N_22538,N_22781);
nand U25868 (N_25868,N_22261,N_22862);
nand U25869 (N_25869,N_23647,N_22018);
xnor U25870 (N_25870,N_22696,N_23872);
or U25871 (N_25871,N_23969,N_22460);
or U25872 (N_25872,N_22525,N_23081);
nand U25873 (N_25873,N_22592,N_23458);
xnor U25874 (N_25874,N_22918,N_23795);
or U25875 (N_25875,N_23854,N_23531);
xnor U25876 (N_25876,N_22946,N_22155);
or U25877 (N_25877,N_23737,N_22041);
nand U25878 (N_25878,N_22917,N_22072);
or U25879 (N_25879,N_23236,N_22278);
nor U25880 (N_25880,N_22725,N_23385);
nand U25881 (N_25881,N_23446,N_23333);
or U25882 (N_25882,N_23757,N_23108);
nand U25883 (N_25883,N_22209,N_22440);
or U25884 (N_25884,N_22540,N_23222);
or U25885 (N_25885,N_22859,N_23338);
and U25886 (N_25886,N_22213,N_23103);
and U25887 (N_25887,N_22644,N_23206);
or U25888 (N_25888,N_22140,N_23250);
or U25889 (N_25889,N_22356,N_22412);
or U25890 (N_25890,N_23444,N_22146);
xnor U25891 (N_25891,N_23492,N_23660);
and U25892 (N_25892,N_22029,N_22628);
and U25893 (N_25893,N_23784,N_23515);
or U25894 (N_25894,N_22622,N_22092);
and U25895 (N_25895,N_23858,N_22948);
or U25896 (N_25896,N_23326,N_22796);
xnor U25897 (N_25897,N_23076,N_22444);
nand U25898 (N_25898,N_22839,N_23572);
nand U25899 (N_25899,N_22129,N_22488);
and U25900 (N_25900,N_22521,N_23159);
and U25901 (N_25901,N_23040,N_23941);
or U25902 (N_25902,N_22380,N_22404);
nor U25903 (N_25903,N_22379,N_22892);
and U25904 (N_25904,N_23625,N_23627);
nor U25905 (N_25905,N_23554,N_23956);
nand U25906 (N_25906,N_22171,N_22175);
xor U25907 (N_25907,N_23748,N_22201);
and U25908 (N_25908,N_22080,N_23063);
xor U25909 (N_25909,N_22927,N_23247);
or U25910 (N_25910,N_22213,N_22484);
and U25911 (N_25911,N_23739,N_23349);
xor U25912 (N_25912,N_23097,N_22196);
or U25913 (N_25913,N_22580,N_22734);
and U25914 (N_25914,N_23920,N_23834);
nor U25915 (N_25915,N_22020,N_22125);
nor U25916 (N_25916,N_23620,N_22846);
or U25917 (N_25917,N_22957,N_23637);
and U25918 (N_25918,N_23880,N_23371);
nand U25919 (N_25919,N_23953,N_22707);
xnor U25920 (N_25920,N_23690,N_22944);
nor U25921 (N_25921,N_23667,N_22914);
xnor U25922 (N_25922,N_22592,N_22706);
and U25923 (N_25923,N_23955,N_23926);
nor U25924 (N_25924,N_23866,N_22827);
or U25925 (N_25925,N_23709,N_22610);
or U25926 (N_25926,N_22047,N_22171);
and U25927 (N_25927,N_23295,N_22447);
nor U25928 (N_25928,N_23068,N_22263);
nand U25929 (N_25929,N_22335,N_22509);
or U25930 (N_25930,N_22811,N_22250);
and U25931 (N_25931,N_23957,N_23125);
nor U25932 (N_25932,N_22977,N_23872);
or U25933 (N_25933,N_22355,N_23183);
or U25934 (N_25934,N_22609,N_22374);
nor U25935 (N_25935,N_23225,N_23130);
xor U25936 (N_25936,N_23790,N_23258);
nand U25937 (N_25937,N_22118,N_22179);
and U25938 (N_25938,N_22050,N_22097);
nor U25939 (N_25939,N_22301,N_22252);
or U25940 (N_25940,N_22566,N_23697);
nor U25941 (N_25941,N_22197,N_23191);
nand U25942 (N_25942,N_23052,N_22883);
or U25943 (N_25943,N_23695,N_23613);
nor U25944 (N_25944,N_22530,N_22595);
xor U25945 (N_25945,N_23742,N_22014);
nor U25946 (N_25946,N_22425,N_22877);
nand U25947 (N_25947,N_22595,N_23387);
nor U25948 (N_25948,N_23117,N_22522);
xor U25949 (N_25949,N_22204,N_23957);
and U25950 (N_25950,N_22993,N_23612);
nand U25951 (N_25951,N_22718,N_22927);
nand U25952 (N_25952,N_22451,N_22304);
and U25953 (N_25953,N_23982,N_23037);
xnor U25954 (N_25954,N_23728,N_23262);
or U25955 (N_25955,N_23313,N_22594);
nor U25956 (N_25956,N_22233,N_23358);
nand U25957 (N_25957,N_22763,N_22708);
and U25958 (N_25958,N_22765,N_22639);
or U25959 (N_25959,N_22157,N_23893);
xor U25960 (N_25960,N_23030,N_22636);
nand U25961 (N_25961,N_23605,N_22041);
and U25962 (N_25962,N_23145,N_22199);
nor U25963 (N_25963,N_23587,N_22895);
or U25964 (N_25964,N_22100,N_22740);
and U25965 (N_25965,N_22297,N_22103);
and U25966 (N_25966,N_23511,N_22242);
xor U25967 (N_25967,N_23561,N_22086);
or U25968 (N_25968,N_22562,N_22163);
nor U25969 (N_25969,N_23068,N_22136);
nand U25970 (N_25970,N_22577,N_23144);
nand U25971 (N_25971,N_23069,N_23170);
or U25972 (N_25972,N_22913,N_23493);
nor U25973 (N_25973,N_22699,N_22731);
nand U25974 (N_25974,N_23146,N_22522);
xor U25975 (N_25975,N_23322,N_22959);
and U25976 (N_25976,N_22920,N_22201);
xor U25977 (N_25977,N_22568,N_22514);
and U25978 (N_25978,N_22692,N_23209);
nand U25979 (N_25979,N_23442,N_23522);
nor U25980 (N_25980,N_23829,N_22641);
and U25981 (N_25981,N_23005,N_23546);
nor U25982 (N_25982,N_23324,N_22115);
nand U25983 (N_25983,N_22508,N_22091);
and U25984 (N_25984,N_22742,N_23479);
or U25985 (N_25985,N_23620,N_22437);
and U25986 (N_25986,N_23650,N_22546);
and U25987 (N_25987,N_23573,N_23390);
nand U25988 (N_25988,N_23133,N_23248);
or U25989 (N_25989,N_23261,N_23232);
xor U25990 (N_25990,N_23628,N_22340);
nand U25991 (N_25991,N_23298,N_23634);
nand U25992 (N_25992,N_22295,N_23605);
or U25993 (N_25993,N_22589,N_22181);
xor U25994 (N_25994,N_23002,N_23645);
nor U25995 (N_25995,N_22987,N_22268);
xor U25996 (N_25996,N_23700,N_23263);
nand U25997 (N_25997,N_23113,N_23115);
nand U25998 (N_25998,N_22939,N_23841);
or U25999 (N_25999,N_22621,N_22309);
and U26000 (N_26000,N_24326,N_24951);
nand U26001 (N_26001,N_24687,N_25606);
nand U26002 (N_26002,N_25251,N_24035);
nand U26003 (N_26003,N_24046,N_25124);
nor U26004 (N_26004,N_25748,N_25696);
nand U26005 (N_26005,N_25485,N_25930);
nor U26006 (N_26006,N_24370,N_25872);
or U26007 (N_26007,N_24107,N_24066);
nand U26008 (N_26008,N_24462,N_25396);
or U26009 (N_26009,N_25732,N_25878);
nor U26010 (N_26010,N_25196,N_24501);
or U26011 (N_26011,N_24560,N_25900);
xnor U26012 (N_26012,N_24496,N_24784);
nand U26013 (N_26013,N_24682,N_25572);
or U26014 (N_26014,N_25404,N_24468);
xor U26015 (N_26015,N_25240,N_25136);
nand U26016 (N_26016,N_25645,N_24477);
nand U26017 (N_26017,N_24990,N_25583);
xnor U26018 (N_26018,N_25468,N_24328);
and U26019 (N_26019,N_25891,N_24313);
nor U26020 (N_26020,N_24242,N_25267);
nor U26021 (N_26021,N_24236,N_24371);
xnor U26022 (N_26022,N_24749,N_24243);
and U26023 (N_26023,N_25046,N_24667);
or U26024 (N_26024,N_24985,N_24886);
nor U26025 (N_26025,N_25208,N_25429);
nor U26026 (N_26026,N_25566,N_24546);
nor U26027 (N_26027,N_25321,N_24137);
and U26028 (N_26028,N_25083,N_25339);
nor U26029 (N_26029,N_24217,N_24769);
xor U26030 (N_26030,N_24524,N_24274);
and U26031 (N_26031,N_24516,N_24879);
and U26032 (N_26032,N_25436,N_24393);
xnor U26033 (N_26033,N_24513,N_24356);
nor U26034 (N_26034,N_24998,N_24644);
or U26035 (N_26035,N_24541,N_25184);
and U26036 (N_26036,N_24811,N_25264);
or U26037 (N_26037,N_25987,N_25159);
xor U26038 (N_26038,N_25706,N_24450);
xnor U26039 (N_26039,N_25305,N_25947);
nor U26040 (N_26040,N_25835,N_24821);
xor U26041 (N_26041,N_25307,N_25150);
nor U26042 (N_26042,N_25912,N_25420);
and U26043 (N_26043,N_25644,N_25996);
and U26044 (N_26044,N_25211,N_24453);
nand U26045 (N_26045,N_25178,N_24210);
or U26046 (N_26046,N_24744,N_25418);
and U26047 (N_26047,N_25460,N_24130);
and U26048 (N_26048,N_24936,N_24401);
and U26049 (N_26049,N_25304,N_24551);
or U26050 (N_26050,N_24658,N_24941);
nor U26051 (N_26051,N_25326,N_24799);
or U26052 (N_26052,N_25742,N_24089);
xnor U26053 (N_26053,N_24207,N_25683);
or U26054 (N_26054,N_24997,N_24613);
or U26055 (N_26055,N_25935,N_25260);
xor U26056 (N_26056,N_25509,N_25800);
nor U26057 (N_26057,N_24475,N_24659);
or U26058 (N_26058,N_24676,N_24818);
xor U26059 (N_26059,N_24752,N_25301);
xor U26060 (N_26060,N_25443,N_25920);
or U26061 (N_26061,N_25454,N_24686);
or U26062 (N_26062,N_24261,N_25517);
and U26063 (N_26063,N_24763,N_24669);
or U26064 (N_26064,N_25491,N_24014);
or U26065 (N_26065,N_25385,N_25607);
xnor U26066 (N_26066,N_25838,N_24023);
nor U26067 (N_26067,N_25831,N_25475);
xnor U26068 (N_26068,N_24467,N_25882);
nand U26069 (N_26069,N_24302,N_25245);
nor U26070 (N_26070,N_24798,N_25568);
or U26071 (N_26071,N_24090,N_24262);
xnor U26072 (N_26072,N_24947,N_25204);
xor U26073 (N_26073,N_24314,N_24160);
nor U26074 (N_26074,N_25833,N_24465);
and U26075 (N_26075,N_24753,N_25248);
xor U26076 (N_26076,N_25603,N_24322);
xor U26077 (N_26077,N_24754,N_25155);
xnor U26078 (N_26078,N_24479,N_25357);
or U26079 (N_26079,N_24995,N_25837);
or U26080 (N_26080,N_25777,N_25044);
and U26081 (N_26081,N_24052,N_24907);
nor U26082 (N_26082,N_24823,N_24643);
xnor U26083 (N_26083,N_25582,N_24797);
nor U26084 (N_26084,N_24257,N_24295);
nand U26085 (N_26085,N_25822,N_25378);
nand U26086 (N_26086,N_25598,N_25705);
and U26087 (N_26087,N_25259,N_25297);
xnor U26088 (N_26088,N_25537,N_24157);
nand U26089 (N_26089,N_25229,N_24306);
xor U26090 (N_26090,N_24151,N_24522);
nor U26091 (N_26091,N_24408,N_25788);
and U26092 (N_26092,N_24276,N_24665);
and U26093 (N_26093,N_25415,N_24204);
nor U26094 (N_26094,N_24645,N_25074);
and U26095 (N_26095,N_25678,N_25444);
nor U26096 (N_26096,N_24855,N_24525);
and U26097 (N_26097,N_24296,N_25254);
nand U26098 (N_26098,N_25423,N_25666);
xnor U26099 (N_26099,N_24115,N_25699);
nor U26100 (N_26100,N_24913,N_24367);
nor U26101 (N_26101,N_25463,N_25299);
nand U26102 (N_26102,N_25352,N_25309);
or U26103 (N_26103,N_24580,N_25702);
and U26104 (N_26104,N_25784,N_25981);
and U26105 (N_26105,N_25172,N_24238);
and U26106 (N_26106,N_25675,N_24374);
xnor U26107 (N_26107,N_24178,N_24869);
xnor U26108 (N_26108,N_25375,N_25275);
xnor U26109 (N_26109,N_25439,N_24901);
and U26110 (N_26110,N_24471,N_24171);
nor U26111 (N_26111,N_24535,N_25764);
nor U26112 (N_26112,N_24926,N_24868);
xnor U26113 (N_26113,N_24074,N_25232);
xnor U26114 (N_26114,N_24455,N_24846);
nor U26115 (N_26115,N_24149,N_24139);
and U26116 (N_26116,N_25745,N_25035);
xnor U26117 (N_26117,N_24768,N_25515);
and U26118 (N_26118,N_24632,N_24069);
nor U26119 (N_26119,N_24812,N_24668);
nand U26120 (N_26120,N_24215,N_25815);
xor U26121 (N_26121,N_25173,N_24838);
nor U26122 (N_26122,N_25048,N_24365);
xnor U26123 (N_26123,N_25661,N_25365);
and U26124 (N_26124,N_24590,N_24076);
nand U26125 (N_26125,N_25885,N_24950);
and U26126 (N_26126,N_24737,N_24033);
nand U26127 (N_26127,N_25697,N_25356);
or U26128 (N_26128,N_24542,N_24212);
and U26129 (N_26129,N_25962,N_24547);
and U26130 (N_26130,N_25290,N_25883);
and U26131 (N_26131,N_25113,N_24004);
nand U26132 (N_26132,N_25970,N_24954);
or U26133 (N_26133,N_24618,N_25643);
nor U26134 (N_26134,N_24241,N_24826);
and U26135 (N_26135,N_25968,N_24379);
and U26136 (N_26136,N_25410,N_24303);
or U26137 (N_26137,N_25589,N_24949);
and U26138 (N_26138,N_24427,N_25752);
xnor U26139 (N_26139,N_24728,N_24843);
or U26140 (N_26140,N_25343,N_25002);
xnor U26141 (N_26141,N_25556,N_25425);
and U26142 (N_26142,N_24445,N_25482);
nor U26143 (N_26143,N_24751,N_25999);
nand U26144 (N_26144,N_25668,N_25479);
nand U26145 (N_26145,N_24724,N_24860);
and U26146 (N_26146,N_24279,N_24042);
xnor U26147 (N_26147,N_24795,N_25462);
xnor U26148 (N_26148,N_24219,N_24121);
nand U26149 (N_26149,N_25544,N_25677);
and U26150 (N_26150,N_25819,N_24536);
nand U26151 (N_26151,N_24135,N_24267);
nor U26152 (N_26152,N_25632,N_24862);
xor U26153 (N_26153,N_25104,N_25709);
and U26154 (N_26154,N_25472,N_25789);
nor U26155 (N_26155,N_25669,N_25754);
nor U26156 (N_26156,N_24406,N_25862);
nor U26157 (N_26157,N_24452,N_25884);
nor U26158 (N_26158,N_24413,N_25262);
nor U26159 (N_26159,N_24248,N_24931);
or U26160 (N_26160,N_25353,N_24125);
nand U26161 (N_26161,N_25873,N_25653);
xnor U26162 (N_26162,N_25360,N_25899);
xor U26163 (N_26163,N_24189,N_25400);
or U26164 (N_26164,N_24266,N_24012);
nand U26165 (N_26165,N_24515,N_25198);
nor U26166 (N_26166,N_24589,N_25086);
xor U26167 (N_26167,N_25327,N_24310);
and U26168 (N_26168,N_24946,N_25183);
nand U26169 (N_26169,N_24109,N_25610);
xor U26170 (N_26170,N_25380,N_25160);
and U26171 (N_26171,N_25918,N_25836);
nor U26172 (N_26172,N_24581,N_24150);
nor U26173 (N_26173,N_25246,N_24593);
and U26174 (N_26174,N_25293,N_24654);
nor U26175 (N_26175,N_24308,N_25540);
xor U26176 (N_26176,N_24263,N_25016);
nor U26177 (N_26177,N_25413,N_24369);
or U26178 (N_26178,N_25757,N_24801);
xnor U26179 (N_26179,N_25006,N_25255);
and U26180 (N_26180,N_25521,N_24329);
xnor U26181 (N_26181,N_24509,N_24566);
xor U26182 (N_26182,N_24388,N_25256);
xnor U26183 (N_26183,N_25986,N_25909);
or U26184 (N_26184,N_24761,N_25477);
and U26185 (N_26185,N_25504,N_24316);
and U26186 (N_26186,N_25557,N_24113);
and U26187 (N_26187,N_24169,N_25488);
or U26188 (N_26188,N_25876,N_24773);
and U26189 (N_26189,N_24835,N_25421);
and U26190 (N_26190,N_24794,N_24389);
nand U26191 (N_26191,N_24019,N_25931);
and U26192 (N_26192,N_25648,N_25176);
and U26193 (N_26193,N_25871,N_25760);
nand U26194 (N_26194,N_25153,N_24483);
or U26195 (N_26195,N_24982,N_24853);
nor U26196 (N_26196,N_24214,N_24866);
nand U26197 (N_26197,N_25192,N_24372);
nor U26198 (N_26198,N_24832,N_25750);
and U26199 (N_26199,N_25126,N_24854);
nand U26200 (N_26200,N_25334,N_25059);
nand U26201 (N_26201,N_24143,N_25671);
and U26202 (N_26202,N_24670,N_25470);
or U26203 (N_26203,N_25503,N_25190);
nor U26204 (N_26204,N_25852,N_25547);
or U26205 (N_26205,N_25880,N_24146);
and U26206 (N_26206,N_25584,N_24619);
or U26207 (N_26207,N_24772,N_25977);
and U26208 (N_26208,N_25201,N_24786);
or U26209 (N_26209,N_24271,N_25657);
nand U26210 (N_26210,N_24708,N_25511);
nand U26211 (N_26211,N_25911,N_25199);
xnor U26212 (N_26212,N_24747,N_25573);
xor U26213 (N_26213,N_24384,N_24805);
xnor U26214 (N_26214,N_25213,N_25522);
xor U26215 (N_26215,N_24932,N_24544);
xor U26216 (N_26216,N_24474,N_25455);
xor U26217 (N_26217,N_25170,N_25816);
nor U26218 (N_26218,N_24063,N_24916);
nand U26219 (N_26219,N_24630,N_25386);
nand U26220 (N_26220,N_24079,N_25585);
nand U26221 (N_26221,N_24834,N_25938);
xor U26222 (N_26222,N_25019,N_24315);
nand U26223 (N_26223,N_25391,N_25285);
nand U26224 (N_26224,N_25805,N_24182);
or U26225 (N_26225,N_24284,N_25730);
nor U26226 (N_26226,N_25039,N_25781);
and U26227 (N_26227,N_24489,N_25793);
or U26228 (N_26228,N_24902,N_25801);
or U26229 (N_26229,N_24438,N_24918);
xnor U26230 (N_26230,N_24208,N_24681);
and U26231 (N_26231,N_25091,N_25771);
xor U26232 (N_26232,N_25839,N_24021);
or U26233 (N_26233,N_25261,N_24764);
nand U26234 (N_26234,N_25928,N_25227);
nand U26235 (N_26235,N_25561,N_24988);
and U26236 (N_26236,N_24221,N_24490);
xnor U26237 (N_26237,N_24195,N_24294);
or U26238 (N_26238,N_25372,N_24830);
nand U26239 (N_26239,N_24211,N_24173);
xor U26240 (N_26240,N_25650,N_24873);
or U26241 (N_26241,N_25973,N_24179);
nand U26242 (N_26242,N_25367,N_25137);
nand U26243 (N_26243,N_25052,N_25217);
xor U26244 (N_26244,N_24712,N_25207);
nand U26245 (N_26245,N_25944,N_24792);
nand U26246 (N_26246,N_24499,N_24337);
xor U26247 (N_26247,N_24549,N_24640);
nand U26248 (N_26248,N_24675,N_24165);
and U26249 (N_26249,N_25812,N_25181);
xor U26250 (N_26250,N_24904,N_24226);
or U26251 (N_26251,N_24819,N_25085);
nand U26252 (N_26252,N_25894,N_24914);
and U26253 (N_26253,N_25971,N_25577);
nand U26254 (N_26254,N_24937,N_24906);
and U26255 (N_26255,N_24766,N_24008);
and U26256 (N_26256,N_25925,N_25937);
xnor U26257 (N_26257,N_24603,N_24225);
nand U26258 (N_26258,N_25312,N_24973);
nor U26259 (N_26259,N_24258,N_25011);
nand U26260 (N_26260,N_25428,N_25924);
and U26261 (N_26261,N_25765,N_25737);
nor U26262 (N_26262,N_24230,N_25348);
or U26263 (N_26263,N_24694,N_24281);
nand U26264 (N_26264,N_25902,N_24697);
xnor U26265 (N_26265,N_24850,N_24105);
or U26266 (N_26266,N_24699,N_24131);
and U26267 (N_26267,N_25140,N_25276);
or U26268 (N_26268,N_25743,N_25412);
nand U26269 (N_26269,N_25791,N_25407);
nor U26270 (N_26270,N_24674,N_24441);
and U26271 (N_26271,N_25888,N_25711);
nand U26272 (N_26272,N_25594,N_25955);
xnor U26273 (N_26273,N_25203,N_24520);
nor U26274 (N_26274,N_24494,N_25629);
or U26275 (N_26275,N_25167,N_24086);
nand U26276 (N_26276,N_25234,N_25630);
or U26277 (N_26277,N_24354,N_24555);
nor U26278 (N_26278,N_24779,N_24880);
and U26279 (N_26279,N_25438,N_25338);
nand U26280 (N_26280,N_25775,N_25257);
xnor U26281 (N_26281,N_25693,N_25435);
xor U26282 (N_26282,N_25325,N_24426);
and U26283 (N_26283,N_25437,N_24975);
and U26284 (N_26284,N_25127,N_24703);
xnor U26285 (N_26285,N_24829,N_24053);
and U26286 (N_26286,N_25316,N_25717);
xor U26287 (N_26287,N_25218,N_25672);
or U26288 (N_26288,N_24177,N_24858);
or U26289 (N_26289,N_25851,N_25563);
nor U26290 (N_26290,N_24098,N_24299);
nand U26291 (N_26291,N_25965,N_24320);
nand U26292 (N_26292,N_24083,N_24287);
nor U26293 (N_26293,N_24085,N_24925);
nand U26294 (N_26294,N_24162,N_24614);
xnor U26295 (N_26295,N_25130,N_25419);
and U26296 (N_26296,N_24727,N_25067);
xnor U26297 (N_26297,N_25782,N_24533);
xor U26298 (N_26298,N_24561,N_24126);
nor U26299 (N_26299,N_25659,N_25692);
xor U26300 (N_26300,N_25111,N_24587);
nor U26301 (N_26301,N_24815,N_25753);
nand U26302 (N_26302,N_24734,N_24142);
and U26303 (N_26303,N_25335,N_25703);
nand U26304 (N_26304,N_24845,N_24748);
xnor U26305 (N_26305,N_25810,N_24220);
nor U26306 (N_26306,N_24391,N_25636);
and U26307 (N_26307,N_25710,N_24713);
and U26308 (N_26308,N_24193,N_24191);
and U26309 (N_26309,N_25623,N_24039);
xnor U26310 (N_26310,N_25725,N_25135);
xor U26311 (N_26311,N_24627,N_24881);
xor U26312 (N_26312,N_24383,N_25071);
and U26313 (N_26313,N_25186,N_24963);
nor U26314 (N_26314,N_24108,N_24222);
and U26315 (N_26315,N_24022,N_25053);
and U26316 (N_26316,N_25310,N_25341);
or U26317 (N_26317,N_24001,N_24203);
xor U26318 (N_26318,N_24335,N_24884);
and U26319 (N_26319,N_25060,N_24852);
or U26320 (N_26320,N_24447,N_24297);
nor U26321 (N_26321,N_25762,N_24404);
xnor U26322 (N_26322,N_24953,N_25690);
or U26323 (N_26323,N_25272,N_25570);
xnor U26324 (N_26324,N_24010,N_25950);
and U26325 (N_26325,N_24449,N_25088);
and U26326 (N_26326,N_25430,N_25179);
or U26327 (N_26327,N_24908,N_24800);
or U26328 (N_26328,N_24631,N_25652);
or U26329 (N_26329,N_25622,N_24205);
nor U26330 (N_26330,N_25593,N_24124);
or U26331 (N_26331,N_25551,N_25863);
nor U26332 (N_26332,N_25929,N_25656);
and U26333 (N_26333,N_25141,N_25721);
or U26334 (N_26334,N_25817,N_25294);
nor U26335 (N_26335,N_25904,N_25337);
and U26336 (N_26336,N_24382,N_25376);
and U26337 (N_26337,N_24293,N_24403);
nand U26338 (N_26338,N_25064,N_24473);
xnor U26339 (N_26339,N_25298,N_24756);
and U26340 (N_26340,N_25770,N_24319);
nor U26341 (N_26341,N_24060,N_24836);
nor U26342 (N_26342,N_25897,N_24414);
nand U26343 (N_26343,N_24332,N_24174);
and U26344 (N_26344,N_24093,N_25082);
and U26345 (N_26345,N_24964,N_25125);
nor U26346 (N_26346,N_25235,N_25646);
and U26347 (N_26347,N_25802,N_25626);
nand U26348 (N_26348,N_24508,N_24484);
and U26349 (N_26349,N_25874,N_24216);
nor U26350 (N_26350,N_24537,N_25003);
nand U26351 (N_26351,N_24806,N_24153);
and U26352 (N_26352,N_25487,N_25205);
nor U26353 (N_26353,N_24782,N_25535);
and U26354 (N_26354,N_25116,N_24478);
xor U26355 (N_26355,N_25118,N_25148);
or U26356 (N_26356,N_25342,N_24323);
or U26357 (N_26357,N_25528,N_24915);
xnor U26358 (N_26358,N_24013,N_24421);
and U26359 (N_26359,N_25004,N_25769);
xor U26360 (N_26360,N_24443,N_24776);
nand U26361 (N_26361,N_24896,N_25998);
nor U26362 (N_26362,N_25825,N_24726);
nand U26363 (N_26363,N_25808,N_24240);
nor U26364 (N_26364,N_24154,N_24428);
xnor U26365 (N_26365,N_25978,N_25156);
nand U26366 (N_26366,N_24094,N_25633);
and U26367 (N_26367,N_24837,N_25966);
xor U26368 (N_26368,N_25456,N_24929);
nor U26369 (N_26369,N_25579,N_24407);
xnor U26370 (N_26370,N_25030,N_25500);
nand U26371 (N_26371,N_24291,N_24698);
nor U26372 (N_26372,N_25489,N_24608);
nor U26373 (N_26373,N_25483,N_24523);
or U26374 (N_26374,N_24134,N_25431);
nand U26375 (N_26375,N_25302,N_25628);
nor U26376 (N_26376,N_24282,N_24650);
nand U26377 (N_26377,N_24605,N_24361);
xor U26378 (N_26378,N_25185,N_25890);
nand U26379 (N_26379,N_25480,N_25426);
or U26380 (N_26380,N_25506,N_25814);
or U26381 (N_26381,N_24984,N_24810);
nor U26382 (N_26382,N_25274,N_24000);
nand U26383 (N_26383,N_24571,N_25370);
xnor U26384 (N_26384,N_25796,N_24198);
and U26385 (N_26385,N_25107,N_24129);
xor U26386 (N_26386,N_24739,N_24857);
and U26387 (N_26387,N_25219,N_24706);
nor U26388 (N_26388,N_25054,N_25898);
nand U26389 (N_26389,N_25673,N_24470);
or U26390 (N_26390,N_24583,N_24788);
nor U26391 (N_26391,N_24395,N_25602);
or U26392 (N_26392,N_24199,N_24999);
and U26393 (N_26393,N_25783,N_25361);
nor U26394 (N_26394,N_25289,N_24935);
or U26395 (N_26395,N_25886,N_25036);
and U26396 (N_26396,N_24979,N_24298);
and U26397 (N_26397,N_25860,N_25225);
nand U26398 (N_26398,N_24759,N_25129);
xor U26399 (N_26399,N_24405,N_24209);
and U26400 (N_26400,N_24588,N_24064);
and U26401 (N_26401,N_24362,N_25571);
xor U26402 (N_26402,N_24288,N_25887);
or U26403 (N_26403,N_25322,N_24570);
and U26404 (N_26404,N_24187,N_25639);
or U26405 (N_26405,N_24342,N_24194);
or U26406 (N_26406,N_24285,N_25820);
and U26407 (N_26407,N_24133,N_25486);
or U26408 (N_26408,N_25383,N_25772);
or U26409 (N_26409,N_24624,N_24368);
nand U26410 (N_26410,N_24223,N_24062);
or U26411 (N_26411,N_25624,N_25457);
or U26412 (N_26412,N_25271,N_24700);
or U26413 (N_26413,N_24817,N_24715);
or U26414 (N_26414,N_25660,N_24009);
xor U26415 (N_26415,N_25247,N_24972);
and U26416 (N_26416,N_24026,N_24486);
or U26417 (N_26417,N_24557,N_25471);
or U26418 (N_26418,N_25993,N_24436);
nor U26419 (N_26419,N_25151,N_24202);
nor U26420 (N_26420,N_24092,N_25637);
nand U26421 (N_26421,N_24859,N_25040);
nand U26422 (N_26422,N_24307,N_25465);
or U26423 (N_26423,N_25027,N_24331);
nand U26424 (N_26424,N_25724,N_25168);
nor U26425 (N_26425,N_24265,N_24155);
and U26426 (N_26426,N_25013,N_24055);
or U26427 (N_26427,N_25662,N_24185);
and U26428 (N_26428,N_24604,N_25381);
or U26429 (N_26429,N_24638,N_25287);
and U26430 (N_26430,N_24943,N_24690);
and U26431 (N_26431,N_25490,N_25879);
nand U26432 (N_26432,N_24061,N_24188);
or U26433 (N_26433,N_24575,N_24777);
or U26434 (N_26434,N_24986,N_24967);
nor U26435 (N_26435,N_25923,N_24161);
or U26436 (N_26436,N_25450,N_25394);
nor U26437 (N_26437,N_24980,N_25362);
nor U26438 (N_26438,N_25138,N_25895);
nor U26439 (N_26439,N_25744,N_25231);
and U26440 (N_26440,N_24548,N_24987);
or U26441 (N_26441,N_25134,N_25065);
or U26442 (N_26442,N_24373,N_24793);
and U26443 (N_26443,N_24027,N_25829);
and U26444 (N_26444,N_25280,N_24492);
and U26445 (N_26445,N_24636,N_24920);
xor U26446 (N_26446,N_24623,N_25798);
nand U26447 (N_26447,N_24377,N_24924);
nor U26448 (N_26448,N_24635,N_25286);
xor U26449 (N_26449,N_25665,N_24218);
nand U26450 (N_26450,N_25020,N_24101);
xnor U26451 (N_26451,N_24529,N_25073);
or U26452 (N_26452,N_25214,N_25976);
nor U26453 (N_26453,N_24976,N_25530);
and U26454 (N_26454,N_25096,N_25242);
or U26455 (N_26455,N_25038,N_24305);
xnor U26456 (N_26456,N_25440,N_25516);
or U26457 (N_26457,N_24378,N_25574);
or U26458 (N_26458,N_24625,N_25452);
nand U26459 (N_26459,N_25007,N_25684);
nor U26460 (N_26460,N_25875,N_25761);
nand U26461 (N_26461,N_25842,N_24442);
nand U26462 (N_26462,N_25663,N_24360);
nand U26463 (N_26463,N_24729,N_25560);
and U26464 (N_26464,N_25514,N_25110);
nand U26465 (N_26465,N_25145,N_24289);
or U26466 (N_26466,N_24647,N_25499);
xor U26467 (N_26467,N_24420,N_25406);
or U26468 (N_26468,N_25519,N_25202);
nand U26469 (N_26469,N_24435,N_24190);
nand U26470 (N_26470,N_24965,N_25034);
xor U26471 (N_26471,N_24770,N_24132);
or U26472 (N_26472,N_24646,N_25171);
or U26473 (N_26473,N_24228,N_24045);
xor U26474 (N_26474,N_25344,N_25467);
and U26475 (N_26475,N_24273,N_25719);
and U26476 (N_26476,N_25680,N_24528);
xnor U26477 (N_26477,N_25569,N_25651);
nor U26478 (N_26478,N_25131,N_24419);
or U26479 (N_26479,N_25401,N_24424);
and U26480 (N_26480,N_24514,N_25114);
nor U26481 (N_26481,N_25609,N_25508);
and U26482 (N_26482,N_25278,N_25850);
or U26483 (N_26483,N_25809,N_25824);
xnor U26484 (N_26484,N_24292,N_24206);
and U26485 (N_26485,N_25913,N_24683);
nor U26486 (N_26486,N_25575,N_25994);
and U26487 (N_26487,N_24167,N_25910);
or U26488 (N_26488,N_25253,N_24321);
nand U26489 (N_26489,N_24497,N_25230);
nor U26490 (N_26490,N_24526,N_25269);
or U26491 (N_26491,N_24791,N_25857);
and U26492 (N_26492,N_25615,N_24876);
xnor U26493 (N_26493,N_24755,N_25492);
or U26494 (N_26494,N_25078,N_25000);
and U26495 (N_26495,N_25161,N_25854);
or U26496 (N_26496,N_25350,N_25300);
or U26497 (N_26497,N_25658,N_24184);
and U26498 (N_26498,N_24586,N_24550);
or U26499 (N_26499,N_25949,N_24084);
xor U26500 (N_26500,N_25513,N_25523);
and U26501 (N_26501,N_25476,N_25209);
and U26502 (N_26502,N_25984,N_25936);
and U26503 (N_26503,N_24741,N_25858);
xor U26504 (N_26504,N_24567,N_24485);
or U26505 (N_26505,N_24434,N_25712);
nand U26506 (N_26506,N_24011,N_24396);
xnor U26507 (N_26507,N_24096,N_24839);
nand U26508 (N_26508,N_24034,N_25466);
xnor U26509 (N_26509,N_24574,N_24410);
xnor U26510 (N_26510,N_25351,N_25823);
nand U26511 (N_26511,N_24231,N_24911);
and U26512 (N_26512,N_24981,N_25474);
nand U26513 (N_26513,N_24488,N_25635);
nor U26514 (N_26514,N_25333,N_25195);
and U26515 (N_26515,N_25731,N_24917);
nand U26516 (N_26516,N_25057,N_24164);
and U26517 (N_26517,N_24458,N_24140);
or U26518 (N_26518,N_25197,N_25591);
nor U26519 (N_26519,N_25451,N_25481);
or U26520 (N_26520,N_24530,N_24685);
and U26521 (N_26521,N_24970,N_24503);
nand U26522 (N_26522,N_24933,N_25933);
nor U26523 (N_26523,N_24343,N_24227);
nand U26524 (N_26524,N_25881,N_24390);
nor U26525 (N_26525,N_25713,N_25926);
xnor U26526 (N_26526,N_24969,N_25614);
nand U26527 (N_26527,N_24280,N_25283);
nor U26528 (N_26528,N_25258,N_25469);
xnor U26529 (N_26529,N_24927,N_24874);
or U26530 (N_26530,N_24849,N_25249);
and U26531 (N_26531,N_24464,N_24993);
and U26532 (N_26532,N_25548,N_24082);
nor U26533 (N_26533,N_25856,N_25206);
xnor U26534 (N_26534,N_25969,N_25042);
or U26535 (N_26535,N_24720,N_24259);
nor U26536 (N_26536,N_25893,N_25704);
or U26537 (N_26537,N_25080,N_25586);
nor U26538 (N_26538,N_24456,N_25273);
nor U26539 (N_26539,N_25346,N_25464);
nor U26540 (N_26540,N_24738,N_25964);
or U26541 (N_26541,N_24163,N_24606);
and U26542 (N_26542,N_24740,N_25414);
or U26543 (N_26543,N_25292,N_25022);
or U26544 (N_26544,N_24088,N_24730);
nor U26545 (N_26545,N_24938,N_24861);
nor U26546 (N_26546,N_24460,N_24887);
or U26547 (N_26547,N_25708,N_24312);
or U26548 (N_26548,N_24330,N_25954);
and U26549 (N_26549,N_25787,N_25539);
nor U26550 (N_26550,N_24781,N_25374);
and U26551 (N_26551,N_24017,N_24015);
xnor U26552 (N_26552,N_24928,N_24412);
xor U26553 (N_26553,N_24498,N_24695);
or U26554 (N_26554,N_25952,N_25432);
and U26555 (N_26555,N_24380,N_24582);
nor U26556 (N_26556,N_25832,N_25720);
or U26557 (N_26557,N_25821,N_24422);
xor U26558 (N_26558,N_25369,N_24357);
and U26559 (N_26559,N_24563,N_25728);
nand U26560 (N_26560,N_24192,N_25306);
or U26561 (N_26561,N_24318,N_25943);
and U26562 (N_26562,N_25459,N_24554);
or U26563 (N_26563,N_24693,N_25618);
or U26564 (N_26564,N_24003,N_24552);
nand U26565 (N_26565,N_24510,N_24816);
and U26566 (N_26566,N_25605,N_25371);
and U26567 (N_26567,N_24511,N_24930);
or U26568 (N_26568,N_25695,N_25921);
xnor U26569 (N_26569,N_25620,N_24651);
and U26570 (N_26570,N_24080,N_25473);
xor U26571 (N_26571,N_25021,N_25980);
or U26572 (N_26572,N_24504,N_24111);
xnor U26573 (N_26573,N_25616,N_25368);
or U26574 (N_26574,N_25433,N_24844);
nand U26575 (N_26575,N_25177,N_25600);
nand U26576 (N_26576,N_25580,N_25767);
xor U26577 (N_26577,N_25799,N_24648);
nand U26578 (N_26578,N_25087,N_24666);
nor U26579 (N_26579,N_25077,N_25484);
or U26580 (N_26580,N_25641,N_25510);
xor U26581 (N_26581,N_25097,N_25288);
or U26582 (N_26582,N_24716,N_25549);
nand U26583 (N_26583,N_25538,N_25552);
xor U26584 (N_26584,N_24783,N_25405);
nand U26585 (N_26585,N_25773,N_25101);
nor U26586 (N_26586,N_25967,N_25193);
nand U26587 (N_26587,N_24156,N_24607);
nand U26588 (N_26588,N_25093,N_25157);
or U26589 (N_26589,N_24123,N_24556);
and U26590 (N_26590,N_25688,N_25100);
xor U26591 (N_26591,N_24872,N_25152);
and U26592 (N_26592,N_25774,N_25296);
nand U26593 (N_26593,N_24100,N_25345);
nor U26594 (N_26594,N_25106,N_25018);
nand U26595 (N_26595,N_25281,N_24448);
nor U26596 (N_26596,N_24628,N_24024);
nor U26597 (N_26597,N_25252,N_24482);
or U26598 (N_26598,N_24041,N_25266);
xor U26599 (N_26599,N_24237,N_24903);
and U26600 (N_26600,N_24264,N_25942);
nor U26601 (N_26601,N_25389,N_25811);
or U26602 (N_26602,N_24431,N_25453);
nor U26603 (N_26603,N_25498,N_25595);
nor U26604 (N_26604,N_25449,N_24745);
nor U26605 (N_26605,N_24186,N_24359);
nand U26606 (N_26606,N_24025,N_24991);
and U26607 (N_26607,N_25961,N_24376);
nor U26608 (N_26608,N_24762,N_24059);
and U26609 (N_26609,N_25212,N_24594);
nor U26610 (N_26610,N_24506,N_25043);
or U26611 (N_26611,N_24275,N_25390);
nor U26612 (N_26612,N_25050,N_25682);
nand U26613 (N_26613,N_25117,N_24457);
xor U26614 (N_26614,N_24820,N_25045);
and U26615 (N_26615,N_25397,N_24346);
nor U26616 (N_26616,N_25953,N_24517);
nand U26617 (N_26617,N_25865,N_25109);
or U26618 (N_26618,N_24235,N_24057);
nor U26619 (N_26619,N_24112,N_24277);
and U26620 (N_26620,N_25983,N_24657);
or U26621 (N_26621,N_24742,N_24073);
or U26622 (N_26622,N_24599,N_24634);
and U26623 (N_26623,N_24591,N_24197);
and U26624 (N_26624,N_24145,N_24122);
nand U26625 (N_26625,N_24957,N_25495);
nand U26626 (N_26626,N_24775,N_25358);
and U26627 (N_26627,N_25914,N_25501);
nor U26628 (N_26628,N_24364,N_24717);
nand U26629 (N_26629,N_24244,N_25768);
xnor U26630 (N_26630,N_25716,N_24891);
or U26631 (N_26631,N_25102,N_25318);
xnor U26632 (N_26632,N_25237,N_25478);
nor U26633 (N_26633,N_25975,N_24956);
nor U26634 (N_26634,N_25939,N_25216);
nor U26635 (N_26635,N_25531,N_25359);
or U26636 (N_26636,N_24890,N_24002);
and U26637 (N_26637,N_24176,N_25869);
nand U26638 (N_26638,N_25051,N_25445);
nand U26639 (N_26639,N_25896,N_25543);
nor U26640 (N_26640,N_25840,N_24272);
nand U26641 (N_26641,N_24399,N_24573);
and U26642 (N_26642,N_25502,N_25447);
nand U26643 (N_26643,N_25578,N_24239);
xnor U26644 (N_26644,N_24333,N_24172);
nor U26645 (N_26645,N_25377,N_25363);
and U26646 (N_26646,N_25562,N_25069);
xnor U26647 (N_26647,N_25158,N_24680);
or U26648 (N_26648,N_24934,N_24558);
and U26649 (N_26649,N_24867,N_24596);
nor U26650 (N_26650,N_24097,N_24559);
and U26651 (N_26651,N_25032,N_24158);
xnor U26652 (N_26652,N_25149,N_25689);
nor U26653 (N_26653,N_24989,N_24334);
xor U26654 (N_26654,N_25903,N_24641);
xnor U26655 (N_26655,N_24543,N_25388);
xor U26656 (N_26656,N_24255,N_24679);
xor U26657 (N_26657,N_24611,N_24610);
xor U26658 (N_26658,N_24663,N_24592);
or U26659 (N_26659,N_25596,N_24180);
nor U26660 (N_26660,N_25989,N_25685);
xor U26661 (N_26661,N_24044,N_24181);
nand U26662 (N_26662,N_24743,N_25906);
nor U26663 (N_26663,N_25849,N_25354);
xnor U26664 (N_26664,N_25277,N_24521);
nand U26665 (N_26665,N_24507,N_24750);
nand U26666 (N_26666,N_24895,N_24353);
nor U26667 (N_26667,N_25625,N_24116);
nand U26668 (N_26668,N_25581,N_25324);
and U26669 (N_26669,N_24527,N_24653);
or U26670 (N_26670,N_25366,N_25393);
xor U26671 (N_26671,N_24723,N_25864);
nand U26672 (N_26672,N_24710,N_24400);
or U26673 (N_26673,N_25055,N_25529);
xor U26674 (N_26674,N_24067,N_25763);
xor U26675 (N_26675,N_24565,N_25681);
nor U26676 (N_26676,N_25755,N_24392);
nand U26677 (N_26677,N_24885,N_24958);
nor U26678 (N_26678,N_25759,N_25047);
xor U26679 (N_26679,N_24301,N_25014);
nand U26680 (N_26680,N_24796,N_25715);
nand U26681 (N_26681,N_24701,N_25619);
nand U26682 (N_26682,N_25988,N_24939);
nor U26683 (N_26683,N_25005,N_24091);
or U26684 (N_26684,N_25590,N_24616);
nand U26685 (N_26685,N_25103,N_24531);
nor U26686 (N_26686,N_25597,N_25340);
nor U26687 (N_26687,N_24397,N_25241);
and U26688 (N_26688,N_24444,N_25907);
nor U26689 (N_26689,N_24899,N_24758);
nor U26690 (N_26690,N_25210,N_25676);
nor U26691 (N_26691,N_24429,N_24028);
nor U26692 (N_26692,N_24341,N_24200);
xor U26693 (N_26693,N_25608,N_24833);
or U26694 (N_26694,N_24324,N_24856);
and U26695 (N_26695,N_25349,N_25518);
xnor U26696 (N_26696,N_24629,N_24688);
nor U26697 (N_26697,N_24883,N_25555);
nand U26698 (N_26698,N_25075,N_24278);
xnor U26699 (N_26699,N_24711,N_25139);
nor U26700 (N_26700,N_24840,N_25826);
nand U26701 (N_26701,N_24099,N_24300);
nor U26702 (N_26702,N_24787,N_25422);
nor U26703 (N_26703,N_25142,N_24851);
and U26704 (N_26704,N_24662,N_25861);
or U26705 (N_26705,N_25940,N_24677);
nand U26706 (N_26706,N_24336,N_25559);
or U26707 (N_26707,N_24898,N_24540);
nand U26708 (N_26708,N_24269,N_24725);
or U26709 (N_26709,N_24709,N_24348);
nor U26710 (N_26710,N_25105,N_24340);
and U26711 (N_26711,N_25601,N_25092);
nor U26712 (N_26712,N_24411,N_24168);
or U26713 (N_26713,N_25834,N_24040);
xor U26714 (N_26714,N_25997,N_24183);
or U26715 (N_26715,N_24036,N_24398);
xor U26716 (N_26716,N_25332,N_24942);
nand U26717 (N_26717,N_24601,N_25766);
and U26718 (N_26718,N_24409,N_25734);
or U26719 (N_26719,N_25576,N_24553);
nand U26720 (N_26720,N_25494,N_25402);
nand U26721 (N_26721,N_25200,N_24251);
and U26722 (N_26722,N_24808,N_25613);
or U26723 (N_26723,N_24472,N_25806);
xor U26724 (N_26724,N_25236,N_24661);
xor U26725 (N_26725,N_24807,N_25162);
xor U26726 (N_26726,N_25963,N_24254);
xor U26727 (N_26727,N_24809,N_24070);
nor U26728 (N_26728,N_24637,N_25461);
or U26729 (N_26729,N_24897,N_25941);
or U26730 (N_26730,N_24454,N_24119);
or U26731 (N_26731,N_25956,N_24358);
xnor U26732 (N_26732,N_25604,N_24102);
nand U26733 (N_26733,N_24945,N_24141);
nand U26734 (N_26734,N_25691,N_25025);
nor U26735 (N_26735,N_25664,N_25427);
and U26736 (N_26736,N_24234,N_24325);
or U26737 (N_26737,N_25037,N_25546);
nor U26738 (N_26738,N_24966,N_25587);
nand U26739 (N_26739,N_25617,N_25194);
and U26740 (N_26740,N_24983,N_24539);
nand U26741 (N_26741,N_25497,N_25945);
nand U26742 (N_26742,N_24481,N_25017);
and U26743 (N_26743,N_24138,N_24765);
nor U26744 (N_26744,N_25336,N_24612);
nand U26745 (N_26745,N_25319,N_24718);
xor U26746 (N_26746,N_24780,N_24311);
xnor U26747 (N_26747,N_24355,N_25959);
or U26748 (N_26748,N_25634,N_25794);
xnor U26749 (N_26749,N_24050,N_24774);
nand U26750 (N_26750,N_25532,N_25033);
and U26751 (N_26751,N_24534,N_25189);
or U26752 (N_26752,N_24863,N_24152);
and U26753 (N_26753,N_25403,N_24439);
xnor U26754 (N_26754,N_24948,N_24664);
nand U26755 (N_26755,N_25654,N_25686);
or U26756 (N_26756,N_25001,N_25934);
nand U26757 (N_26757,N_25747,N_24451);
nor U26758 (N_26758,N_24250,N_25553);
or U26759 (N_26759,N_25112,N_25424);
nand U26760 (N_26760,N_25133,N_24469);
xor U26761 (N_26761,N_25736,N_24117);
or U26762 (N_26762,N_24778,N_25847);
or U26763 (N_26763,N_24994,N_24018);
nor U26764 (N_26764,N_24476,N_25785);
xnor U26765 (N_26765,N_25029,N_24803);
nand U26766 (N_26766,N_25756,N_24095);
nor U26767 (N_26767,N_25175,N_25063);
nand U26768 (N_26768,N_24136,N_24038);
or U26769 (N_26769,N_24923,N_25946);
xor U26770 (N_26770,N_25778,N_25303);
nand U26771 (N_26771,N_25746,N_25056);
and U26772 (N_26772,N_24696,N_25417);
nand U26773 (N_26773,N_25442,N_25263);
nor U26774 (N_26774,N_25739,N_25222);
and U26775 (N_26775,N_25008,N_25979);
nand U26776 (N_26776,N_24127,N_24888);
or U26777 (N_26777,N_25070,N_25960);
nand U26778 (N_26778,N_24466,N_25524);
xnor U26779 (N_26779,N_24007,N_24912);
nand U26780 (N_26780,N_25848,N_24166);
nand U26781 (N_26781,N_24871,N_24043);
nor U26782 (N_26782,N_25146,N_24201);
or U26783 (N_26783,N_25015,N_24639);
and U26784 (N_26784,N_25434,N_24692);
xor U26785 (N_26785,N_25621,N_25841);
nor U26786 (N_26786,N_25076,N_25496);
xor U26787 (N_26787,N_24363,N_24961);
nor U26788 (N_26788,N_24992,N_24030);
nand U26789 (N_26789,N_24538,N_24345);
nor U26790 (N_26790,N_24595,N_25655);
or U26791 (N_26791,N_25991,N_24246);
or U26792 (N_26792,N_24955,N_25244);
nand U26793 (N_26793,N_25889,N_24005);
nor U26794 (N_26794,N_25163,N_25233);
and U26795 (N_26795,N_25166,N_24463);
nor U26796 (N_26796,N_24051,N_25187);
nand U26797 (N_26797,N_24016,N_25638);
nand U26798 (N_26798,N_24785,N_25536);
or U26799 (N_26799,N_24804,N_25009);
xor U26800 (N_26800,N_24600,N_25507);
or U26801 (N_26801,N_24350,N_24652);
and U26802 (N_26802,N_25012,N_24339);
or U26803 (N_26803,N_25957,N_24078);
nor U26804 (N_26804,N_25905,N_25411);
xnor U26805 (N_26805,N_24617,N_24344);
xor U26806 (N_26806,N_24626,N_25674);
nor U26807 (N_26807,N_24789,N_24381);
and U26808 (N_26808,N_24037,N_25095);
and U26809 (N_26809,N_24736,N_24072);
nand U26810 (N_26810,N_25182,N_24978);
or U26811 (N_26811,N_24425,N_25062);
nor U26812 (N_26812,N_25972,N_24620);
nor U26813 (N_26813,N_24921,N_25061);
nor U26814 (N_26814,N_25174,N_25512);
nor U26815 (N_26815,N_25908,N_24048);
or U26816 (N_26816,N_24579,N_25099);
xor U26817 (N_26817,N_25776,N_24684);
xor U26818 (N_26818,N_25119,N_24394);
nor U26819 (N_26819,N_24385,N_24633);
nand U26820 (N_26820,N_25010,N_24831);
nand U26821 (N_26821,N_25533,N_25079);
nand U26822 (N_26822,N_24996,N_25611);
nor U26823 (N_26823,N_24719,N_24564);
and U26824 (N_26824,N_24878,N_24366);
nor U26825 (N_26825,N_25373,N_25314);
xor U26826 (N_26826,N_24842,N_25859);
nor U26827 (N_26827,N_25550,N_25220);
xnor U26828 (N_26828,N_25317,N_25919);
nor U26829 (N_26829,N_25631,N_25108);
and U26830 (N_26830,N_24290,N_24375);
nand U26831 (N_26831,N_24317,N_24568);
or U26832 (N_26832,N_25416,N_25308);
and U26833 (N_26833,N_24224,N_24968);
or U26834 (N_26834,N_24502,N_24252);
nor U26835 (N_26835,N_24569,N_25387);
xor U26836 (N_26836,N_24847,N_24415);
nor U26837 (N_26837,N_25541,N_24865);
nand U26838 (N_26838,N_24196,N_24487);
xnor U26839 (N_26839,N_25165,N_25687);
or U26840 (N_26840,N_25877,N_25714);
or U26841 (N_26841,N_24491,N_25328);
and U26842 (N_26842,N_25827,N_25870);
or U26843 (N_26843,N_25031,N_24106);
or U26844 (N_26844,N_24656,N_24922);
nor U26845 (N_26845,N_25554,N_24232);
nor U26846 (N_26846,N_25722,N_24671);
and U26847 (N_26847,N_25121,N_25384);
nand U26848 (N_26848,N_24767,N_24075);
xor U26849 (N_26849,N_24678,N_24732);
xor U26850 (N_26850,N_24735,N_25855);
nand U26851 (N_26851,N_25243,N_25917);
nand U26852 (N_26852,N_25392,N_25382);
or U26853 (N_26853,N_25493,N_25313);
xnor U26854 (N_26854,N_24144,N_24500);
and U26855 (N_26855,N_25120,N_25948);
xnor U26856 (N_26856,N_25291,N_24351);
nor U26857 (N_26857,N_24602,N_25398);
xor U26858 (N_26858,N_24461,N_24721);
nor U26859 (N_26859,N_24875,N_24870);
nand U26860 (N_26860,N_24952,N_25786);
nand U26861 (N_26861,N_24813,N_24147);
nand U26862 (N_26862,N_24256,N_24822);
or U26863 (N_26863,N_24087,N_25525);
nor U26864 (N_26864,N_25331,N_24233);
xnor U26865 (N_26865,N_24418,N_24578);
or U26866 (N_26866,N_25740,N_25311);
xnor U26867 (N_26867,N_25558,N_25409);
nor U26868 (N_26868,N_25221,N_24814);
nor U26869 (N_26869,N_25347,N_25098);
nand U26870 (N_26870,N_24213,N_25542);
xor U26871 (N_26871,N_25853,N_25995);
nor U26872 (N_26872,N_25723,N_25395);
xor U26873 (N_26873,N_25818,N_25446);
nand U26874 (N_26874,N_24584,N_25779);
xnor U26875 (N_26875,N_25932,N_25505);
nor U26876 (N_26876,N_24848,N_25023);
and U26877 (N_26877,N_25599,N_24705);
or U26878 (N_26878,N_25028,N_25068);
nand U26879 (N_26879,N_24058,N_25279);
xor U26880 (N_26880,N_25828,N_24722);
nor U26881 (N_26881,N_25534,N_25084);
or U26882 (N_26882,N_25089,N_25527);
nor U26883 (N_26883,N_24495,N_24689);
xnor U26884 (N_26884,N_25188,N_25330);
and U26885 (N_26885,N_24054,N_24673);
xnor U26886 (N_26886,N_25807,N_24077);
and U26887 (N_26887,N_24104,N_24597);
and U26888 (N_26888,N_25951,N_24402);
xor U26889 (N_26889,N_24047,N_25081);
nand U26890 (N_26890,N_24349,N_25790);
or U26891 (N_26891,N_25974,N_24691);
nor U26892 (N_26892,N_24572,N_25797);
and U26893 (N_26893,N_25751,N_24148);
nand U26894 (N_26894,N_24841,N_24020);
and U26895 (N_26895,N_24029,N_24974);
and U26896 (N_26896,N_25592,N_24905);
xnor U26897 (N_26897,N_25698,N_24120);
xor U26898 (N_26898,N_24828,N_25901);
and U26899 (N_26899,N_24430,N_24889);
and U26900 (N_26900,N_24286,N_25627);
xor U26901 (N_26901,N_25545,N_24621);
or U26902 (N_26902,N_25667,N_25115);
or U26903 (N_26903,N_24440,N_24423);
nor U26904 (N_26904,N_25320,N_25868);
and U26905 (N_26905,N_25215,N_25892);
or U26906 (N_26906,N_25180,N_25458);
xor U26907 (N_26907,N_25647,N_24229);
or U26908 (N_26908,N_24577,N_24714);
xnor U26909 (N_26909,N_25564,N_25990);
or U26910 (N_26910,N_25122,N_24437);
xor U26911 (N_26911,N_25804,N_24505);
and U26912 (N_26912,N_24519,N_24245);
xnor U26913 (N_26913,N_24327,N_25694);
nor U26914 (N_26914,N_25749,N_24672);
xnor U26915 (N_26915,N_25448,N_24253);
nor U26916 (N_26916,N_25701,N_25726);
nor U26917 (N_26917,N_24827,N_24480);
nor U26918 (N_26918,N_24433,N_25024);
and U26919 (N_26919,N_25399,N_25565);
xnor U26920 (N_26920,N_25364,N_25164);
and U26921 (N_26921,N_24309,N_24446);
and U26922 (N_26922,N_24864,N_25520);
or U26923 (N_26923,N_24270,N_25191);
and U26924 (N_26924,N_25315,N_24562);
nor U26925 (N_26925,N_24900,N_25803);
and U26926 (N_26926,N_25700,N_24006);
nand U26927 (N_26927,N_24175,N_24493);
nor U26928 (N_26928,N_24352,N_25226);
and U26929 (N_26929,N_24910,N_24247);
and U26930 (N_26930,N_24893,N_24283);
nor U26931 (N_26931,N_24940,N_25927);
and U26932 (N_26932,N_24068,N_25642);
xor U26933 (N_26933,N_25355,N_25223);
xnor U26934 (N_26934,N_25143,N_25741);
and U26935 (N_26935,N_24733,N_24103);
nand U26936 (N_26936,N_24532,N_25649);
xnor U26937 (N_26937,N_25094,N_25228);
nor U26938 (N_26938,N_25844,N_25058);
and U26939 (N_26939,N_25985,N_24249);
xor U26940 (N_26940,N_25238,N_24802);
nor U26941 (N_26941,N_24660,N_25792);
nand U26942 (N_26942,N_25958,N_25323);
xnor U26943 (N_26943,N_25729,N_25670);
nor U26944 (N_26944,N_24771,N_25830);
and U26945 (N_26945,N_24268,N_24959);
or U26946 (N_26946,N_24609,N_24909);
or U26947 (N_26947,N_24545,N_25735);
nand U26948 (N_26948,N_25295,N_25916);
xnor U26949 (N_26949,N_24065,N_24877);
and U26950 (N_26950,N_25270,N_25795);
nor U26951 (N_26951,N_25250,N_24892);
and U26952 (N_26952,N_24731,N_24760);
and U26953 (N_26953,N_24110,N_24757);
nand U26954 (N_26954,N_25707,N_24704);
and U26955 (N_26955,N_25982,N_25813);
nand U26956 (N_26956,N_25379,N_24944);
or U26957 (N_26957,N_25612,N_24128);
and U26958 (N_26958,N_25846,N_25147);
xnor U26959 (N_26959,N_25567,N_24649);
nand U26960 (N_26960,N_25922,N_25132);
or U26961 (N_26961,N_25284,N_24585);
or U26962 (N_26962,N_24655,N_25867);
nand U26963 (N_26963,N_24260,N_25727);
and U26964 (N_26964,N_25679,N_25718);
nor U26965 (N_26965,N_24971,N_24049);
xor U26966 (N_26966,N_25026,N_25041);
nand U26967 (N_26967,N_24882,N_25329);
and U26968 (N_26968,N_25758,N_25072);
and U26969 (N_26969,N_24432,N_24416);
nor U26970 (N_26970,N_24114,N_24338);
nand U26971 (N_26971,N_25738,N_25066);
or U26972 (N_26972,N_25526,N_24702);
xor U26973 (N_26973,N_24576,N_25049);
or U26974 (N_26974,N_25265,N_24598);
or U26975 (N_26975,N_25733,N_24615);
nand U26976 (N_26976,N_24417,N_25866);
nand U26977 (N_26977,N_25640,N_24081);
xnor U26978 (N_26978,N_24459,N_24622);
nor U26979 (N_26979,N_24159,N_25090);
or U26980 (N_26980,N_24977,N_24031);
and U26981 (N_26981,N_25169,N_24387);
xnor U26982 (N_26982,N_24512,N_24056);
nand U26983 (N_26983,N_24642,N_25224);
xnor U26984 (N_26984,N_24304,N_25408);
and U26985 (N_26985,N_25239,N_24518);
nand U26986 (N_26986,N_25992,N_24746);
xor U26987 (N_26987,N_24707,N_24386);
nand U26988 (N_26988,N_25845,N_24347);
or U26989 (N_26989,N_24919,N_25588);
xor U26990 (N_26990,N_24825,N_25282);
xor U26991 (N_26991,N_25154,N_25843);
or U26992 (N_26992,N_24962,N_25128);
nor U26993 (N_26993,N_25144,N_24790);
and U26994 (N_26994,N_24824,N_24960);
nand U26995 (N_26995,N_24894,N_24118);
and U26996 (N_26996,N_24170,N_24032);
xnor U26997 (N_26997,N_24071,N_25780);
nor U26998 (N_26998,N_25123,N_25268);
nand U26999 (N_26999,N_25915,N_25441);
xnor U27000 (N_27000,N_24810,N_25652);
nor U27001 (N_27001,N_25390,N_24489);
or U27002 (N_27002,N_25453,N_25321);
xor U27003 (N_27003,N_24063,N_24032);
nand U27004 (N_27004,N_24034,N_25979);
and U27005 (N_27005,N_25514,N_25424);
and U27006 (N_27006,N_24481,N_24826);
nor U27007 (N_27007,N_25579,N_24204);
or U27008 (N_27008,N_25733,N_25097);
nand U27009 (N_27009,N_24006,N_25655);
nand U27010 (N_27010,N_24549,N_24649);
nand U27011 (N_27011,N_25995,N_25564);
or U27012 (N_27012,N_25667,N_24028);
nor U27013 (N_27013,N_25732,N_24973);
xnor U27014 (N_27014,N_25505,N_25836);
and U27015 (N_27015,N_24855,N_25580);
and U27016 (N_27016,N_25298,N_24498);
or U27017 (N_27017,N_25088,N_24023);
xnor U27018 (N_27018,N_24838,N_24874);
or U27019 (N_27019,N_25976,N_24134);
nand U27020 (N_27020,N_24849,N_25824);
or U27021 (N_27021,N_24397,N_24491);
nor U27022 (N_27022,N_24950,N_25215);
nand U27023 (N_27023,N_24097,N_25958);
and U27024 (N_27024,N_25315,N_24551);
nand U27025 (N_27025,N_24786,N_25159);
and U27026 (N_27026,N_24132,N_25313);
nand U27027 (N_27027,N_24032,N_24287);
nand U27028 (N_27028,N_25610,N_25960);
and U27029 (N_27029,N_25416,N_25457);
xor U27030 (N_27030,N_25994,N_24883);
xnor U27031 (N_27031,N_24246,N_24632);
nand U27032 (N_27032,N_25529,N_25034);
nor U27033 (N_27033,N_25981,N_25006);
and U27034 (N_27034,N_24220,N_24892);
nand U27035 (N_27035,N_25157,N_24618);
nand U27036 (N_27036,N_25227,N_25413);
nand U27037 (N_27037,N_24877,N_25586);
nor U27038 (N_27038,N_24163,N_25379);
and U27039 (N_27039,N_24124,N_25603);
and U27040 (N_27040,N_24128,N_25781);
nor U27041 (N_27041,N_25836,N_24798);
xnor U27042 (N_27042,N_25179,N_25056);
and U27043 (N_27043,N_24246,N_24739);
nand U27044 (N_27044,N_24197,N_24860);
and U27045 (N_27045,N_25863,N_24455);
nand U27046 (N_27046,N_25045,N_24844);
or U27047 (N_27047,N_25942,N_24822);
xnor U27048 (N_27048,N_25984,N_25207);
nand U27049 (N_27049,N_24578,N_24566);
nand U27050 (N_27050,N_25964,N_25232);
and U27051 (N_27051,N_25083,N_24914);
and U27052 (N_27052,N_24177,N_25424);
xnor U27053 (N_27053,N_25860,N_25133);
xor U27054 (N_27054,N_25687,N_25932);
xor U27055 (N_27055,N_24732,N_25399);
xnor U27056 (N_27056,N_25566,N_24657);
nor U27057 (N_27057,N_24316,N_24049);
or U27058 (N_27058,N_24907,N_25386);
nor U27059 (N_27059,N_25509,N_25614);
xor U27060 (N_27060,N_25290,N_24229);
xor U27061 (N_27061,N_24709,N_24026);
nand U27062 (N_27062,N_24035,N_24695);
or U27063 (N_27063,N_24941,N_25557);
and U27064 (N_27064,N_24123,N_25197);
nor U27065 (N_27065,N_25918,N_24514);
xor U27066 (N_27066,N_24591,N_25002);
and U27067 (N_27067,N_25039,N_24045);
and U27068 (N_27068,N_24937,N_24991);
nand U27069 (N_27069,N_25650,N_25565);
nor U27070 (N_27070,N_24924,N_24540);
nand U27071 (N_27071,N_25164,N_24233);
and U27072 (N_27072,N_25946,N_24918);
or U27073 (N_27073,N_24146,N_24868);
or U27074 (N_27074,N_25866,N_24775);
nor U27075 (N_27075,N_25277,N_25121);
and U27076 (N_27076,N_24106,N_25291);
xnor U27077 (N_27077,N_24077,N_25575);
nand U27078 (N_27078,N_25527,N_25302);
xnor U27079 (N_27079,N_25284,N_24753);
nor U27080 (N_27080,N_24396,N_24988);
nand U27081 (N_27081,N_24713,N_25749);
and U27082 (N_27082,N_25213,N_25046);
nor U27083 (N_27083,N_24662,N_25885);
nand U27084 (N_27084,N_25464,N_24455);
nor U27085 (N_27085,N_25066,N_25961);
nand U27086 (N_27086,N_24127,N_24987);
or U27087 (N_27087,N_25621,N_24569);
nand U27088 (N_27088,N_25510,N_24050);
nand U27089 (N_27089,N_25681,N_24590);
xor U27090 (N_27090,N_24502,N_25915);
or U27091 (N_27091,N_25485,N_24352);
and U27092 (N_27092,N_24143,N_24821);
nor U27093 (N_27093,N_25270,N_24299);
nor U27094 (N_27094,N_25149,N_25151);
nand U27095 (N_27095,N_24246,N_24979);
nand U27096 (N_27096,N_25513,N_24797);
xor U27097 (N_27097,N_24268,N_25102);
and U27098 (N_27098,N_25214,N_25705);
xor U27099 (N_27099,N_25867,N_25916);
and U27100 (N_27100,N_24655,N_25200);
xnor U27101 (N_27101,N_24342,N_24064);
nand U27102 (N_27102,N_24908,N_24927);
nor U27103 (N_27103,N_25591,N_24646);
nand U27104 (N_27104,N_25093,N_24528);
nand U27105 (N_27105,N_25474,N_25298);
or U27106 (N_27106,N_25170,N_25243);
nand U27107 (N_27107,N_24760,N_25667);
and U27108 (N_27108,N_24336,N_24224);
or U27109 (N_27109,N_25692,N_25895);
xor U27110 (N_27110,N_25000,N_24109);
and U27111 (N_27111,N_25564,N_24277);
or U27112 (N_27112,N_25793,N_25335);
or U27113 (N_27113,N_24314,N_24782);
and U27114 (N_27114,N_24678,N_25615);
nor U27115 (N_27115,N_25551,N_24433);
and U27116 (N_27116,N_25738,N_24709);
nand U27117 (N_27117,N_24820,N_25276);
nand U27118 (N_27118,N_24470,N_25062);
xnor U27119 (N_27119,N_25167,N_24396);
or U27120 (N_27120,N_24288,N_25837);
nor U27121 (N_27121,N_25878,N_25830);
nand U27122 (N_27122,N_24451,N_25735);
xor U27123 (N_27123,N_24468,N_25744);
nand U27124 (N_27124,N_24572,N_24001);
and U27125 (N_27125,N_25557,N_24083);
nand U27126 (N_27126,N_24691,N_25995);
or U27127 (N_27127,N_24197,N_25216);
xor U27128 (N_27128,N_25766,N_25308);
nand U27129 (N_27129,N_24916,N_24539);
nand U27130 (N_27130,N_24300,N_25052);
nand U27131 (N_27131,N_25843,N_24169);
or U27132 (N_27132,N_24542,N_25240);
and U27133 (N_27133,N_25790,N_25585);
and U27134 (N_27134,N_25324,N_25692);
nand U27135 (N_27135,N_24926,N_25112);
nand U27136 (N_27136,N_24859,N_25957);
xnor U27137 (N_27137,N_25207,N_24830);
and U27138 (N_27138,N_25357,N_25893);
or U27139 (N_27139,N_25793,N_24897);
and U27140 (N_27140,N_24943,N_25994);
or U27141 (N_27141,N_24313,N_24731);
nand U27142 (N_27142,N_24784,N_25247);
or U27143 (N_27143,N_24050,N_25404);
or U27144 (N_27144,N_24507,N_25152);
or U27145 (N_27145,N_24542,N_24958);
nor U27146 (N_27146,N_25801,N_25896);
xnor U27147 (N_27147,N_25018,N_25167);
xor U27148 (N_27148,N_24959,N_25146);
xnor U27149 (N_27149,N_25380,N_25926);
nor U27150 (N_27150,N_25025,N_24825);
and U27151 (N_27151,N_25518,N_25133);
xor U27152 (N_27152,N_25570,N_25826);
nand U27153 (N_27153,N_25212,N_25023);
nor U27154 (N_27154,N_24864,N_24274);
or U27155 (N_27155,N_25993,N_25517);
nor U27156 (N_27156,N_24327,N_24462);
nor U27157 (N_27157,N_24368,N_24703);
nand U27158 (N_27158,N_24289,N_25460);
nor U27159 (N_27159,N_24782,N_24592);
xor U27160 (N_27160,N_25634,N_24350);
xnor U27161 (N_27161,N_24654,N_25922);
and U27162 (N_27162,N_24250,N_25818);
nand U27163 (N_27163,N_24349,N_24755);
nor U27164 (N_27164,N_24863,N_24244);
nand U27165 (N_27165,N_24296,N_25481);
and U27166 (N_27166,N_24205,N_24014);
xnor U27167 (N_27167,N_24986,N_25397);
nor U27168 (N_27168,N_25071,N_24689);
xnor U27169 (N_27169,N_24256,N_24557);
and U27170 (N_27170,N_25385,N_25898);
or U27171 (N_27171,N_25329,N_24648);
or U27172 (N_27172,N_25671,N_25881);
xor U27173 (N_27173,N_25603,N_25782);
nand U27174 (N_27174,N_24791,N_24956);
nor U27175 (N_27175,N_25679,N_25687);
nand U27176 (N_27176,N_24969,N_24796);
xnor U27177 (N_27177,N_25596,N_24238);
and U27178 (N_27178,N_25179,N_24792);
xor U27179 (N_27179,N_25496,N_25507);
nor U27180 (N_27180,N_25491,N_25788);
or U27181 (N_27181,N_24319,N_24098);
nor U27182 (N_27182,N_25257,N_25553);
xor U27183 (N_27183,N_25290,N_24789);
or U27184 (N_27184,N_24852,N_25853);
nor U27185 (N_27185,N_25071,N_24629);
and U27186 (N_27186,N_24878,N_25704);
or U27187 (N_27187,N_25777,N_24743);
nor U27188 (N_27188,N_24763,N_25151);
xor U27189 (N_27189,N_24644,N_25504);
xor U27190 (N_27190,N_24110,N_25293);
xor U27191 (N_27191,N_25755,N_24408);
xor U27192 (N_27192,N_25399,N_25721);
nand U27193 (N_27193,N_24370,N_25751);
or U27194 (N_27194,N_24607,N_25621);
xor U27195 (N_27195,N_25640,N_25891);
nor U27196 (N_27196,N_25296,N_25570);
or U27197 (N_27197,N_25821,N_25198);
nand U27198 (N_27198,N_24081,N_24677);
xnor U27199 (N_27199,N_25839,N_25048);
nor U27200 (N_27200,N_24502,N_24360);
nor U27201 (N_27201,N_25942,N_24129);
or U27202 (N_27202,N_24930,N_25702);
and U27203 (N_27203,N_24110,N_24170);
or U27204 (N_27204,N_25585,N_24729);
or U27205 (N_27205,N_25046,N_25965);
nor U27206 (N_27206,N_25343,N_25317);
or U27207 (N_27207,N_25881,N_25723);
or U27208 (N_27208,N_25677,N_25352);
or U27209 (N_27209,N_24131,N_25301);
nand U27210 (N_27210,N_25744,N_25321);
nand U27211 (N_27211,N_24905,N_25059);
xnor U27212 (N_27212,N_24689,N_24435);
or U27213 (N_27213,N_25985,N_25726);
xnor U27214 (N_27214,N_24497,N_24435);
xnor U27215 (N_27215,N_24389,N_25916);
nand U27216 (N_27216,N_25683,N_24273);
nor U27217 (N_27217,N_24076,N_25772);
nor U27218 (N_27218,N_25262,N_24428);
or U27219 (N_27219,N_24103,N_24517);
nor U27220 (N_27220,N_25565,N_24423);
and U27221 (N_27221,N_24163,N_25087);
or U27222 (N_27222,N_25730,N_25673);
nor U27223 (N_27223,N_24227,N_25858);
nor U27224 (N_27224,N_24969,N_25273);
nand U27225 (N_27225,N_25450,N_24333);
nand U27226 (N_27226,N_25339,N_24486);
xor U27227 (N_27227,N_24329,N_25457);
and U27228 (N_27228,N_25806,N_25784);
or U27229 (N_27229,N_25389,N_25615);
nand U27230 (N_27230,N_25665,N_25094);
nor U27231 (N_27231,N_24859,N_24473);
and U27232 (N_27232,N_25088,N_25710);
or U27233 (N_27233,N_25811,N_24351);
or U27234 (N_27234,N_25295,N_24491);
or U27235 (N_27235,N_25148,N_25163);
nor U27236 (N_27236,N_24726,N_24060);
nor U27237 (N_27237,N_24613,N_24357);
and U27238 (N_27238,N_24690,N_25401);
nand U27239 (N_27239,N_25678,N_24654);
nand U27240 (N_27240,N_24412,N_25277);
nand U27241 (N_27241,N_25614,N_24021);
nor U27242 (N_27242,N_25285,N_24550);
or U27243 (N_27243,N_25524,N_24732);
nand U27244 (N_27244,N_25094,N_24371);
and U27245 (N_27245,N_25374,N_25127);
nand U27246 (N_27246,N_24458,N_25097);
or U27247 (N_27247,N_25259,N_24208);
or U27248 (N_27248,N_24655,N_24361);
nand U27249 (N_27249,N_24984,N_24446);
xor U27250 (N_27250,N_24601,N_25767);
nor U27251 (N_27251,N_25968,N_24034);
xnor U27252 (N_27252,N_25901,N_24338);
nand U27253 (N_27253,N_24429,N_24762);
and U27254 (N_27254,N_24729,N_25242);
nand U27255 (N_27255,N_24256,N_25885);
or U27256 (N_27256,N_24870,N_24120);
nand U27257 (N_27257,N_24275,N_25556);
nand U27258 (N_27258,N_24446,N_24368);
nand U27259 (N_27259,N_25724,N_24015);
nand U27260 (N_27260,N_24437,N_25618);
nand U27261 (N_27261,N_25103,N_24830);
and U27262 (N_27262,N_25391,N_24831);
xor U27263 (N_27263,N_25157,N_25611);
nor U27264 (N_27264,N_24246,N_24404);
nand U27265 (N_27265,N_24014,N_25326);
and U27266 (N_27266,N_24208,N_25262);
and U27267 (N_27267,N_25034,N_24380);
or U27268 (N_27268,N_25434,N_24164);
nor U27269 (N_27269,N_24828,N_24190);
nand U27270 (N_27270,N_25140,N_25190);
or U27271 (N_27271,N_25313,N_25943);
xor U27272 (N_27272,N_25055,N_24979);
or U27273 (N_27273,N_25721,N_25484);
or U27274 (N_27274,N_25090,N_25255);
nand U27275 (N_27275,N_25457,N_24071);
or U27276 (N_27276,N_24805,N_24213);
nand U27277 (N_27277,N_25550,N_25807);
or U27278 (N_27278,N_24176,N_25336);
xor U27279 (N_27279,N_24872,N_25510);
xnor U27280 (N_27280,N_24028,N_24869);
nor U27281 (N_27281,N_24555,N_25950);
or U27282 (N_27282,N_24954,N_24825);
nand U27283 (N_27283,N_25483,N_25602);
nand U27284 (N_27284,N_24384,N_24079);
nand U27285 (N_27285,N_24010,N_24952);
or U27286 (N_27286,N_24954,N_24880);
nand U27287 (N_27287,N_24556,N_24179);
nand U27288 (N_27288,N_24209,N_24985);
nor U27289 (N_27289,N_24899,N_24834);
nand U27290 (N_27290,N_25432,N_25413);
xnor U27291 (N_27291,N_25979,N_25735);
nand U27292 (N_27292,N_25921,N_25065);
xor U27293 (N_27293,N_25875,N_24884);
nor U27294 (N_27294,N_24515,N_25705);
nor U27295 (N_27295,N_24306,N_25442);
nand U27296 (N_27296,N_25229,N_25918);
and U27297 (N_27297,N_25879,N_24583);
nand U27298 (N_27298,N_25887,N_25424);
xor U27299 (N_27299,N_24557,N_25192);
and U27300 (N_27300,N_24569,N_24570);
and U27301 (N_27301,N_24552,N_24394);
nand U27302 (N_27302,N_25070,N_25219);
or U27303 (N_27303,N_25130,N_25354);
and U27304 (N_27304,N_25369,N_24484);
nor U27305 (N_27305,N_25396,N_25924);
and U27306 (N_27306,N_25291,N_24860);
or U27307 (N_27307,N_25145,N_25226);
nor U27308 (N_27308,N_24443,N_25677);
and U27309 (N_27309,N_24196,N_25401);
nand U27310 (N_27310,N_24040,N_25812);
or U27311 (N_27311,N_25602,N_24604);
and U27312 (N_27312,N_25196,N_25284);
and U27313 (N_27313,N_24737,N_25358);
or U27314 (N_27314,N_24677,N_24726);
and U27315 (N_27315,N_25371,N_24125);
or U27316 (N_27316,N_24024,N_24912);
nor U27317 (N_27317,N_25378,N_25951);
and U27318 (N_27318,N_24711,N_25803);
and U27319 (N_27319,N_25692,N_24778);
xor U27320 (N_27320,N_25405,N_24034);
or U27321 (N_27321,N_24889,N_24128);
and U27322 (N_27322,N_24421,N_24709);
and U27323 (N_27323,N_24135,N_24890);
nand U27324 (N_27324,N_24364,N_24940);
or U27325 (N_27325,N_25831,N_25328);
xnor U27326 (N_27326,N_24883,N_24015);
xnor U27327 (N_27327,N_24436,N_24935);
and U27328 (N_27328,N_24473,N_24592);
xor U27329 (N_27329,N_24831,N_24803);
nand U27330 (N_27330,N_24991,N_24821);
or U27331 (N_27331,N_25202,N_24001);
and U27332 (N_27332,N_25530,N_25813);
nand U27333 (N_27333,N_25322,N_24950);
and U27334 (N_27334,N_24700,N_25872);
xor U27335 (N_27335,N_25452,N_25671);
or U27336 (N_27336,N_25179,N_24022);
nand U27337 (N_27337,N_24208,N_25995);
or U27338 (N_27338,N_25229,N_25411);
xnor U27339 (N_27339,N_25052,N_24798);
nand U27340 (N_27340,N_25662,N_24749);
nand U27341 (N_27341,N_25487,N_25278);
xnor U27342 (N_27342,N_25751,N_24092);
xnor U27343 (N_27343,N_25319,N_25467);
or U27344 (N_27344,N_25062,N_24908);
xnor U27345 (N_27345,N_24580,N_24681);
or U27346 (N_27346,N_24649,N_24675);
xor U27347 (N_27347,N_25342,N_24979);
nand U27348 (N_27348,N_25068,N_25306);
nor U27349 (N_27349,N_25120,N_25016);
nor U27350 (N_27350,N_25238,N_25036);
or U27351 (N_27351,N_25578,N_24364);
xor U27352 (N_27352,N_25559,N_25218);
xor U27353 (N_27353,N_25628,N_25647);
xnor U27354 (N_27354,N_24761,N_25541);
and U27355 (N_27355,N_24966,N_25584);
xor U27356 (N_27356,N_24806,N_25294);
xor U27357 (N_27357,N_25421,N_24962);
nor U27358 (N_27358,N_25966,N_24812);
or U27359 (N_27359,N_25885,N_25704);
nand U27360 (N_27360,N_25978,N_24786);
xor U27361 (N_27361,N_25546,N_25352);
xnor U27362 (N_27362,N_25809,N_24520);
nand U27363 (N_27363,N_25087,N_25160);
nor U27364 (N_27364,N_24857,N_24345);
and U27365 (N_27365,N_25452,N_25256);
nand U27366 (N_27366,N_25337,N_25402);
nor U27367 (N_27367,N_25430,N_24286);
nand U27368 (N_27368,N_24838,N_25966);
xor U27369 (N_27369,N_25220,N_24207);
and U27370 (N_27370,N_24262,N_25440);
and U27371 (N_27371,N_25458,N_25232);
nand U27372 (N_27372,N_24865,N_25252);
nand U27373 (N_27373,N_25352,N_24987);
xnor U27374 (N_27374,N_24381,N_25447);
or U27375 (N_27375,N_25515,N_25317);
nand U27376 (N_27376,N_24471,N_24062);
and U27377 (N_27377,N_24169,N_24917);
and U27378 (N_27378,N_24716,N_24960);
or U27379 (N_27379,N_25513,N_24443);
xor U27380 (N_27380,N_24648,N_25044);
or U27381 (N_27381,N_25633,N_24571);
nand U27382 (N_27382,N_24471,N_24893);
nand U27383 (N_27383,N_24627,N_25872);
nand U27384 (N_27384,N_24100,N_24768);
xor U27385 (N_27385,N_24402,N_25297);
nand U27386 (N_27386,N_25150,N_25273);
and U27387 (N_27387,N_25477,N_24149);
nor U27388 (N_27388,N_25728,N_25309);
xnor U27389 (N_27389,N_25733,N_24027);
nand U27390 (N_27390,N_24845,N_25274);
nand U27391 (N_27391,N_25284,N_25037);
xnor U27392 (N_27392,N_25621,N_24879);
or U27393 (N_27393,N_25969,N_25749);
nand U27394 (N_27394,N_25223,N_25131);
nor U27395 (N_27395,N_24029,N_24897);
nor U27396 (N_27396,N_24783,N_24541);
or U27397 (N_27397,N_24804,N_25062);
xnor U27398 (N_27398,N_24031,N_24606);
xnor U27399 (N_27399,N_24498,N_24930);
and U27400 (N_27400,N_24796,N_24551);
nand U27401 (N_27401,N_24409,N_24651);
nand U27402 (N_27402,N_25937,N_24520);
or U27403 (N_27403,N_25178,N_24450);
xor U27404 (N_27404,N_24619,N_25401);
xnor U27405 (N_27405,N_24059,N_25808);
nor U27406 (N_27406,N_24110,N_25082);
xor U27407 (N_27407,N_25426,N_25852);
or U27408 (N_27408,N_25756,N_24002);
nor U27409 (N_27409,N_25701,N_24635);
nand U27410 (N_27410,N_24721,N_24596);
and U27411 (N_27411,N_24161,N_25970);
nand U27412 (N_27412,N_24531,N_25509);
nor U27413 (N_27413,N_24115,N_25150);
nor U27414 (N_27414,N_25262,N_25918);
or U27415 (N_27415,N_24461,N_24633);
and U27416 (N_27416,N_24803,N_25079);
xnor U27417 (N_27417,N_25789,N_24185);
xnor U27418 (N_27418,N_25394,N_24540);
xnor U27419 (N_27419,N_24926,N_25864);
nand U27420 (N_27420,N_25333,N_24699);
xor U27421 (N_27421,N_24760,N_25312);
nand U27422 (N_27422,N_24464,N_25367);
and U27423 (N_27423,N_25272,N_24637);
nor U27424 (N_27424,N_25892,N_25055);
xor U27425 (N_27425,N_25706,N_25877);
nand U27426 (N_27426,N_25367,N_24160);
xnor U27427 (N_27427,N_24199,N_24558);
or U27428 (N_27428,N_24752,N_24155);
nor U27429 (N_27429,N_24928,N_25585);
or U27430 (N_27430,N_24005,N_25171);
nand U27431 (N_27431,N_25478,N_24609);
xor U27432 (N_27432,N_25691,N_24308);
or U27433 (N_27433,N_25235,N_25022);
xor U27434 (N_27434,N_24166,N_25432);
xor U27435 (N_27435,N_25400,N_24069);
xor U27436 (N_27436,N_24489,N_24247);
nand U27437 (N_27437,N_25860,N_24928);
nand U27438 (N_27438,N_25063,N_24067);
nand U27439 (N_27439,N_24035,N_24690);
or U27440 (N_27440,N_25070,N_25105);
nand U27441 (N_27441,N_24244,N_25633);
xor U27442 (N_27442,N_25973,N_24762);
and U27443 (N_27443,N_25685,N_24369);
nor U27444 (N_27444,N_24143,N_24013);
nand U27445 (N_27445,N_25026,N_25223);
xnor U27446 (N_27446,N_24256,N_24282);
nand U27447 (N_27447,N_25209,N_25728);
or U27448 (N_27448,N_25247,N_24908);
or U27449 (N_27449,N_25589,N_24747);
or U27450 (N_27450,N_24056,N_24546);
and U27451 (N_27451,N_24270,N_24524);
or U27452 (N_27452,N_25930,N_24982);
or U27453 (N_27453,N_24985,N_24310);
or U27454 (N_27454,N_24562,N_25933);
nor U27455 (N_27455,N_25471,N_25698);
or U27456 (N_27456,N_25934,N_25820);
nor U27457 (N_27457,N_25314,N_24895);
or U27458 (N_27458,N_25464,N_25550);
or U27459 (N_27459,N_24196,N_24098);
or U27460 (N_27460,N_24803,N_24009);
nand U27461 (N_27461,N_24119,N_24875);
xnor U27462 (N_27462,N_25679,N_25337);
xnor U27463 (N_27463,N_24066,N_24374);
xnor U27464 (N_27464,N_25071,N_24069);
nor U27465 (N_27465,N_25672,N_24603);
xnor U27466 (N_27466,N_24327,N_24737);
nor U27467 (N_27467,N_24149,N_24696);
and U27468 (N_27468,N_24927,N_24641);
nand U27469 (N_27469,N_24263,N_24047);
or U27470 (N_27470,N_25526,N_24496);
nand U27471 (N_27471,N_25413,N_25311);
and U27472 (N_27472,N_24849,N_24321);
and U27473 (N_27473,N_25697,N_24811);
xnor U27474 (N_27474,N_25762,N_24802);
nand U27475 (N_27475,N_25197,N_24098);
or U27476 (N_27476,N_25839,N_25526);
xor U27477 (N_27477,N_24901,N_24976);
nand U27478 (N_27478,N_25312,N_25037);
xor U27479 (N_27479,N_25135,N_24232);
or U27480 (N_27480,N_24065,N_24367);
or U27481 (N_27481,N_24508,N_24003);
and U27482 (N_27482,N_24229,N_25504);
nor U27483 (N_27483,N_24861,N_24977);
nand U27484 (N_27484,N_25143,N_25270);
nand U27485 (N_27485,N_25057,N_25760);
nor U27486 (N_27486,N_25149,N_24007);
xor U27487 (N_27487,N_24458,N_25880);
or U27488 (N_27488,N_24265,N_24525);
nor U27489 (N_27489,N_25420,N_25801);
xor U27490 (N_27490,N_24016,N_24096);
nor U27491 (N_27491,N_25768,N_24843);
nor U27492 (N_27492,N_24162,N_24721);
and U27493 (N_27493,N_25424,N_25389);
and U27494 (N_27494,N_25182,N_25531);
nor U27495 (N_27495,N_25208,N_25161);
nor U27496 (N_27496,N_24632,N_25906);
nor U27497 (N_27497,N_25528,N_25565);
and U27498 (N_27498,N_25973,N_25675);
or U27499 (N_27499,N_24005,N_25627);
xnor U27500 (N_27500,N_24821,N_24878);
nor U27501 (N_27501,N_25022,N_24528);
nand U27502 (N_27502,N_24509,N_24985);
xnor U27503 (N_27503,N_24387,N_25867);
nor U27504 (N_27504,N_24076,N_25213);
nor U27505 (N_27505,N_25452,N_24555);
nor U27506 (N_27506,N_25856,N_25298);
and U27507 (N_27507,N_24145,N_25491);
nor U27508 (N_27508,N_25797,N_25105);
or U27509 (N_27509,N_24637,N_24500);
nor U27510 (N_27510,N_24327,N_25163);
and U27511 (N_27511,N_24571,N_24569);
nor U27512 (N_27512,N_24874,N_25193);
nand U27513 (N_27513,N_25791,N_24874);
and U27514 (N_27514,N_24303,N_25697);
or U27515 (N_27515,N_24212,N_24179);
or U27516 (N_27516,N_24437,N_25132);
or U27517 (N_27517,N_25434,N_24922);
nand U27518 (N_27518,N_24366,N_25660);
xor U27519 (N_27519,N_25874,N_24951);
nand U27520 (N_27520,N_24501,N_25219);
nor U27521 (N_27521,N_25295,N_24981);
nor U27522 (N_27522,N_24687,N_24964);
nor U27523 (N_27523,N_25737,N_25154);
nor U27524 (N_27524,N_24077,N_24231);
xor U27525 (N_27525,N_24477,N_25974);
nand U27526 (N_27526,N_24927,N_25167);
xor U27527 (N_27527,N_25728,N_25497);
and U27528 (N_27528,N_24189,N_25843);
nand U27529 (N_27529,N_24835,N_25320);
nand U27530 (N_27530,N_24966,N_24681);
xnor U27531 (N_27531,N_24859,N_24666);
nand U27532 (N_27532,N_24871,N_24255);
or U27533 (N_27533,N_24895,N_25806);
and U27534 (N_27534,N_24035,N_25528);
and U27535 (N_27535,N_25538,N_25773);
nand U27536 (N_27536,N_25803,N_25011);
or U27537 (N_27537,N_24420,N_24603);
nand U27538 (N_27538,N_25920,N_24861);
nor U27539 (N_27539,N_25477,N_24363);
nand U27540 (N_27540,N_25734,N_24980);
or U27541 (N_27541,N_24668,N_24784);
nand U27542 (N_27542,N_24137,N_25934);
xor U27543 (N_27543,N_25307,N_25179);
and U27544 (N_27544,N_24076,N_24817);
nand U27545 (N_27545,N_24402,N_24251);
nand U27546 (N_27546,N_24253,N_24905);
or U27547 (N_27547,N_24916,N_25671);
nor U27548 (N_27548,N_25190,N_24713);
nor U27549 (N_27549,N_25737,N_25386);
nor U27550 (N_27550,N_24337,N_24531);
or U27551 (N_27551,N_25571,N_24343);
and U27552 (N_27552,N_24010,N_25766);
nor U27553 (N_27553,N_24922,N_24658);
or U27554 (N_27554,N_25475,N_24957);
nand U27555 (N_27555,N_25988,N_24874);
xnor U27556 (N_27556,N_25521,N_24227);
nor U27557 (N_27557,N_24688,N_24168);
nand U27558 (N_27558,N_24996,N_24554);
or U27559 (N_27559,N_24352,N_24856);
nor U27560 (N_27560,N_24214,N_24546);
and U27561 (N_27561,N_24698,N_24758);
nor U27562 (N_27562,N_25767,N_25986);
xnor U27563 (N_27563,N_25556,N_24227);
nor U27564 (N_27564,N_24176,N_25858);
xor U27565 (N_27565,N_25849,N_25829);
and U27566 (N_27566,N_25917,N_24372);
and U27567 (N_27567,N_24940,N_25845);
nand U27568 (N_27568,N_25753,N_24336);
or U27569 (N_27569,N_25831,N_25710);
xor U27570 (N_27570,N_25691,N_24378);
nor U27571 (N_27571,N_24114,N_24310);
xor U27572 (N_27572,N_25939,N_25813);
nand U27573 (N_27573,N_25683,N_24161);
or U27574 (N_27574,N_24562,N_25796);
nor U27575 (N_27575,N_25350,N_24803);
nor U27576 (N_27576,N_25353,N_25468);
or U27577 (N_27577,N_25536,N_25589);
nand U27578 (N_27578,N_25390,N_24634);
nand U27579 (N_27579,N_24047,N_25997);
nand U27580 (N_27580,N_25178,N_25572);
nand U27581 (N_27581,N_25685,N_25114);
nand U27582 (N_27582,N_24829,N_25814);
nand U27583 (N_27583,N_25720,N_24994);
or U27584 (N_27584,N_24323,N_24017);
and U27585 (N_27585,N_24580,N_24435);
nand U27586 (N_27586,N_25643,N_24611);
nor U27587 (N_27587,N_25659,N_25181);
nor U27588 (N_27588,N_25349,N_24931);
xor U27589 (N_27589,N_24795,N_24832);
nor U27590 (N_27590,N_24594,N_25547);
nand U27591 (N_27591,N_25678,N_24936);
nor U27592 (N_27592,N_24101,N_24370);
xnor U27593 (N_27593,N_25914,N_24619);
and U27594 (N_27594,N_24947,N_24283);
and U27595 (N_27595,N_24671,N_24716);
or U27596 (N_27596,N_25625,N_24429);
nor U27597 (N_27597,N_25389,N_24279);
nor U27598 (N_27598,N_25037,N_24065);
xor U27599 (N_27599,N_24218,N_24984);
xnor U27600 (N_27600,N_24944,N_24481);
xnor U27601 (N_27601,N_24765,N_24767);
nand U27602 (N_27602,N_24867,N_24765);
nand U27603 (N_27603,N_24104,N_24117);
nand U27604 (N_27604,N_25546,N_24218);
or U27605 (N_27605,N_25296,N_25989);
or U27606 (N_27606,N_25048,N_24574);
nand U27607 (N_27607,N_25360,N_24313);
xor U27608 (N_27608,N_25242,N_25143);
and U27609 (N_27609,N_25783,N_25921);
and U27610 (N_27610,N_24804,N_25174);
nand U27611 (N_27611,N_24216,N_25085);
and U27612 (N_27612,N_25543,N_25152);
xnor U27613 (N_27613,N_25707,N_25519);
nand U27614 (N_27614,N_25115,N_24140);
nand U27615 (N_27615,N_24018,N_25481);
xor U27616 (N_27616,N_25216,N_25095);
nand U27617 (N_27617,N_25085,N_24831);
nand U27618 (N_27618,N_24204,N_25713);
and U27619 (N_27619,N_25970,N_24636);
nor U27620 (N_27620,N_25083,N_24195);
nand U27621 (N_27621,N_25359,N_25567);
nor U27622 (N_27622,N_24589,N_25697);
nor U27623 (N_27623,N_24530,N_24599);
and U27624 (N_27624,N_25209,N_24945);
nor U27625 (N_27625,N_25340,N_24291);
xnor U27626 (N_27626,N_25676,N_25273);
nor U27627 (N_27627,N_24954,N_24198);
and U27628 (N_27628,N_25132,N_24740);
or U27629 (N_27629,N_25302,N_25456);
nand U27630 (N_27630,N_24583,N_25459);
xnor U27631 (N_27631,N_25428,N_24459);
xor U27632 (N_27632,N_25403,N_25251);
nor U27633 (N_27633,N_25194,N_25930);
nand U27634 (N_27634,N_24877,N_24408);
nand U27635 (N_27635,N_24834,N_25611);
or U27636 (N_27636,N_25934,N_25093);
nor U27637 (N_27637,N_24128,N_24317);
or U27638 (N_27638,N_25693,N_25336);
and U27639 (N_27639,N_25629,N_25724);
nand U27640 (N_27640,N_24483,N_25108);
xnor U27641 (N_27641,N_25170,N_24973);
xor U27642 (N_27642,N_24230,N_25957);
nor U27643 (N_27643,N_25736,N_25963);
or U27644 (N_27644,N_25149,N_24112);
xor U27645 (N_27645,N_25824,N_24435);
nor U27646 (N_27646,N_25022,N_25940);
nor U27647 (N_27647,N_25324,N_24296);
or U27648 (N_27648,N_25486,N_24684);
nor U27649 (N_27649,N_24086,N_25497);
nor U27650 (N_27650,N_24871,N_25794);
nor U27651 (N_27651,N_24377,N_24118);
nor U27652 (N_27652,N_25850,N_24118);
or U27653 (N_27653,N_25182,N_24191);
or U27654 (N_27654,N_24691,N_25351);
or U27655 (N_27655,N_24692,N_24712);
nand U27656 (N_27656,N_24175,N_24814);
nor U27657 (N_27657,N_24123,N_24138);
nand U27658 (N_27658,N_25598,N_25125);
xnor U27659 (N_27659,N_24632,N_25069);
or U27660 (N_27660,N_25459,N_25172);
nand U27661 (N_27661,N_25724,N_25933);
xor U27662 (N_27662,N_25488,N_24918);
or U27663 (N_27663,N_24692,N_25094);
xor U27664 (N_27664,N_24549,N_25503);
nor U27665 (N_27665,N_24012,N_24130);
nor U27666 (N_27666,N_25850,N_25542);
nand U27667 (N_27667,N_24811,N_24021);
xnor U27668 (N_27668,N_25463,N_25709);
xor U27669 (N_27669,N_25193,N_24603);
nor U27670 (N_27670,N_25416,N_24557);
or U27671 (N_27671,N_25265,N_25617);
or U27672 (N_27672,N_25643,N_24855);
or U27673 (N_27673,N_25405,N_24692);
or U27674 (N_27674,N_25298,N_25561);
and U27675 (N_27675,N_24765,N_25541);
nand U27676 (N_27676,N_24944,N_25052);
nor U27677 (N_27677,N_25141,N_25045);
and U27678 (N_27678,N_24979,N_25790);
nand U27679 (N_27679,N_24671,N_24295);
or U27680 (N_27680,N_25072,N_25626);
xor U27681 (N_27681,N_25952,N_25446);
nand U27682 (N_27682,N_25698,N_24113);
nor U27683 (N_27683,N_25226,N_25097);
nor U27684 (N_27684,N_24491,N_25160);
or U27685 (N_27685,N_25044,N_25914);
or U27686 (N_27686,N_24092,N_25415);
nor U27687 (N_27687,N_25626,N_24633);
and U27688 (N_27688,N_25535,N_24699);
nor U27689 (N_27689,N_25791,N_25655);
xor U27690 (N_27690,N_25555,N_25284);
nand U27691 (N_27691,N_25466,N_24985);
and U27692 (N_27692,N_24903,N_24194);
xnor U27693 (N_27693,N_24183,N_24357);
xor U27694 (N_27694,N_24296,N_24426);
nand U27695 (N_27695,N_25750,N_25579);
and U27696 (N_27696,N_25566,N_24530);
or U27697 (N_27697,N_24503,N_24675);
or U27698 (N_27698,N_25851,N_25062);
and U27699 (N_27699,N_25848,N_25363);
or U27700 (N_27700,N_25789,N_25696);
nand U27701 (N_27701,N_24058,N_24237);
xnor U27702 (N_27702,N_24055,N_24353);
nand U27703 (N_27703,N_25835,N_25070);
or U27704 (N_27704,N_24260,N_25314);
and U27705 (N_27705,N_25410,N_25623);
and U27706 (N_27706,N_25672,N_25762);
or U27707 (N_27707,N_24048,N_24306);
xor U27708 (N_27708,N_25614,N_24067);
and U27709 (N_27709,N_25269,N_25900);
or U27710 (N_27710,N_25419,N_25515);
xor U27711 (N_27711,N_25745,N_25935);
nor U27712 (N_27712,N_25613,N_24650);
or U27713 (N_27713,N_25312,N_25378);
or U27714 (N_27714,N_25259,N_24447);
nor U27715 (N_27715,N_24683,N_24166);
nor U27716 (N_27716,N_25808,N_24456);
xnor U27717 (N_27717,N_25073,N_24414);
nand U27718 (N_27718,N_25220,N_24175);
nor U27719 (N_27719,N_25938,N_25425);
or U27720 (N_27720,N_24450,N_25447);
and U27721 (N_27721,N_25100,N_25657);
nand U27722 (N_27722,N_25754,N_25566);
xnor U27723 (N_27723,N_25533,N_25257);
and U27724 (N_27724,N_24057,N_24743);
nor U27725 (N_27725,N_24188,N_24607);
and U27726 (N_27726,N_24384,N_24820);
nor U27727 (N_27727,N_24023,N_25082);
xnor U27728 (N_27728,N_25211,N_24374);
and U27729 (N_27729,N_25477,N_25658);
and U27730 (N_27730,N_25636,N_24193);
or U27731 (N_27731,N_24066,N_24611);
nand U27732 (N_27732,N_25683,N_25788);
and U27733 (N_27733,N_24934,N_25642);
or U27734 (N_27734,N_25922,N_24736);
nand U27735 (N_27735,N_25328,N_24401);
or U27736 (N_27736,N_24597,N_24996);
xnor U27737 (N_27737,N_24967,N_25979);
nor U27738 (N_27738,N_25373,N_25080);
nor U27739 (N_27739,N_24294,N_25381);
and U27740 (N_27740,N_25185,N_24399);
and U27741 (N_27741,N_24960,N_24674);
xor U27742 (N_27742,N_24940,N_24873);
and U27743 (N_27743,N_25489,N_24356);
nand U27744 (N_27744,N_24378,N_25178);
or U27745 (N_27745,N_25948,N_25331);
or U27746 (N_27746,N_25558,N_24406);
xor U27747 (N_27747,N_24471,N_24973);
and U27748 (N_27748,N_24424,N_24179);
and U27749 (N_27749,N_25265,N_24918);
nor U27750 (N_27750,N_25527,N_24667);
or U27751 (N_27751,N_25786,N_24069);
nor U27752 (N_27752,N_24497,N_25968);
xnor U27753 (N_27753,N_24440,N_24877);
xor U27754 (N_27754,N_24161,N_25391);
nand U27755 (N_27755,N_25098,N_25999);
nand U27756 (N_27756,N_25501,N_25622);
nor U27757 (N_27757,N_25529,N_24859);
xor U27758 (N_27758,N_24865,N_25919);
and U27759 (N_27759,N_24440,N_24743);
xor U27760 (N_27760,N_25731,N_24530);
nor U27761 (N_27761,N_24377,N_25423);
xor U27762 (N_27762,N_25510,N_25201);
nand U27763 (N_27763,N_24355,N_24272);
and U27764 (N_27764,N_25402,N_24318);
xnor U27765 (N_27765,N_24865,N_24562);
xor U27766 (N_27766,N_25766,N_24481);
or U27767 (N_27767,N_24849,N_24356);
nor U27768 (N_27768,N_25381,N_25690);
nor U27769 (N_27769,N_24812,N_25301);
nor U27770 (N_27770,N_25828,N_25268);
and U27771 (N_27771,N_24272,N_25695);
or U27772 (N_27772,N_24942,N_25414);
and U27773 (N_27773,N_25985,N_25767);
or U27774 (N_27774,N_24953,N_25160);
or U27775 (N_27775,N_24291,N_24623);
or U27776 (N_27776,N_25889,N_25911);
xor U27777 (N_27777,N_25575,N_24131);
nor U27778 (N_27778,N_25579,N_24888);
xnor U27779 (N_27779,N_24823,N_24343);
nand U27780 (N_27780,N_24858,N_24683);
nor U27781 (N_27781,N_24743,N_25095);
xor U27782 (N_27782,N_25964,N_25014);
nand U27783 (N_27783,N_25283,N_25150);
xor U27784 (N_27784,N_24858,N_24501);
and U27785 (N_27785,N_24017,N_25093);
xnor U27786 (N_27786,N_24119,N_25924);
nand U27787 (N_27787,N_25490,N_25070);
nor U27788 (N_27788,N_24918,N_25640);
nor U27789 (N_27789,N_24270,N_24598);
or U27790 (N_27790,N_25088,N_24174);
or U27791 (N_27791,N_25057,N_24159);
or U27792 (N_27792,N_24601,N_25994);
and U27793 (N_27793,N_24958,N_24032);
nand U27794 (N_27794,N_25062,N_24916);
or U27795 (N_27795,N_25520,N_24741);
or U27796 (N_27796,N_25339,N_24996);
xor U27797 (N_27797,N_24177,N_24443);
xnor U27798 (N_27798,N_24526,N_24158);
and U27799 (N_27799,N_25828,N_24625);
and U27800 (N_27800,N_24091,N_24679);
xnor U27801 (N_27801,N_25727,N_24497);
nor U27802 (N_27802,N_25696,N_25417);
xor U27803 (N_27803,N_24921,N_24487);
and U27804 (N_27804,N_25376,N_25789);
xor U27805 (N_27805,N_24856,N_24417);
xor U27806 (N_27806,N_24050,N_25279);
nor U27807 (N_27807,N_24125,N_25794);
xnor U27808 (N_27808,N_25279,N_24806);
nor U27809 (N_27809,N_24586,N_25811);
nand U27810 (N_27810,N_24009,N_25071);
and U27811 (N_27811,N_25386,N_25117);
or U27812 (N_27812,N_25150,N_24580);
nor U27813 (N_27813,N_25001,N_25336);
nor U27814 (N_27814,N_25979,N_24943);
xnor U27815 (N_27815,N_24618,N_25786);
nand U27816 (N_27816,N_25344,N_24347);
and U27817 (N_27817,N_25476,N_24651);
and U27818 (N_27818,N_25178,N_25691);
or U27819 (N_27819,N_24123,N_25640);
nand U27820 (N_27820,N_24800,N_24171);
xnor U27821 (N_27821,N_24996,N_24202);
xnor U27822 (N_27822,N_24188,N_24941);
nand U27823 (N_27823,N_25703,N_24794);
xor U27824 (N_27824,N_24683,N_25610);
nand U27825 (N_27825,N_25994,N_25678);
and U27826 (N_27826,N_24357,N_24676);
xor U27827 (N_27827,N_25110,N_24892);
nand U27828 (N_27828,N_24374,N_25676);
and U27829 (N_27829,N_25681,N_25679);
and U27830 (N_27830,N_25479,N_25920);
nand U27831 (N_27831,N_25943,N_24311);
nor U27832 (N_27832,N_25312,N_25510);
nor U27833 (N_27833,N_25539,N_24001);
nor U27834 (N_27834,N_25177,N_24453);
nor U27835 (N_27835,N_25188,N_25429);
and U27836 (N_27836,N_24315,N_25199);
xor U27837 (N_27837,N_25927,N_24961);
xor U27838 (N_27838,N_24727,N_24173);
nand U27839 (N_27839,N_24134,N_25830);
nand U27840 (N_27840,N_25773,N_24058);
or U27841 (N_27841,N_24527,N_24872);
or U27842 (N_27842,N_25429,N_25696);
and U27843 (N_27843,N_24041,N_25354);
nor U27844 (N_27844,N_25261,N_24322);
or U27845 (N_27845,N_24303,N_24469);
and U27846 (N_27846,N_25691,N_25917);
nand U27847 (N_27847,N_24260,N_25848);
nand U27848 (N_27848,N_25672,N_24876);
or U27849 (N_27849,N_24459,N_25685);
or U27850 (N_27850,N_25234,N_24672);
and U27851 (N_27851,N_24280,N_24115);
xnor U27852 (N_27852,N_24372,N_25101);
nand U27853 (N_27853,N_24717,N_24439);
nand U27854 (N_27854,N_24833,N_24560);
nand U27855 (N_27855,N_25825,N_24178);
and U27856 (N_27856,N_24157,N_24287);
nor U27857 (N_27857,N_24724,N_24113);
nand U27858 (N_27858,N_24921,N_24689);
or U27859 (N_27859,N_24618,N_24155);
xor U27860 (N_27860,N_24361,N_24836);
and U27861 (N_27861,N_24990,N_24967);
or U27862 (N_27862,N_24258,N_24816);
nand U27863 (N_27863,N_25129,N_24340);
xnor U27864 (N_27864,N_24937,N_24549);
nor U27865 (N_27865,N_24835,N_24234);
xor U27866 (N_27866,N_24069,N_24613);
nor U27867 (N_27867,N_24096,N_24879);
nor U27868 (N_27868,N_24856,N_25141);
and U27869 (N_27869,N_24149,N_25859);
xnor U27870 (N_27870,N_25067,N_25454);
or U27871 (N_27871,N_25041,N_25022);
xnor U27872 (N_27872,N_24996,N_24248);
xor U27873 (N_27873,N_25083,N_25089);
nor U27874 (N_27874,N_24702,N_25612);
or U27875 (N_27875,N_24519,N_25067);
or U27876 (N_27876,N_24537,N_24263);
or U27877 (N_27877,N_24787,N_25443);
nor U27878 (N_27878,N_24675,N_25783);
or U27879 (N_27879,N_24957,N_24251);
nand U27880 (N_27880,N_24975,N_25671);
xnor U27881 (N_27881,N_24806,N_24624);
and U27882 (N_27882,N_25429,N_25488);
and U27883 (N_27883,N_25728,N_24792);
or U27884 (N_27884,N_24965,N_24759);
or U27885 (N_27885,N_25858,N_25049);
and U27886 (N_27886,N_25657,N_25337);
nor U27887 (N_27887,N_25046,N_25128);
or U27888 (N_27888,N_24926,N_24215);
nor U27889 (N_27889,N_24418,N_24879);
nor U27890 (N_27890,N_25109,N_24884);
nand U27891 (N_27891,N_24677,N_25218);
xor U27892 (N_27892,N_24860,N_24126);
and U27893 (N_27893,N_25704,N_25536);
nor U27894 (N_27894,N_24501,N_25099);
nor U27895 (N_27895,N_24074,N_25992);
or U27896 (N_27896,N_24910,N_24276);
or U27897 (N_27897,N_24457,N_25709);
nor U27898 (N_27898,N_25799,N_24083);
nor U27899 (N_27899,N_24577,N_24626);
or U27900 (N_27900,N_25770,N_25176);
or U27901 (N_27901,N_25753,N_25258);
nand U27902 (N_27902,N_25563,N_25204);
or U27903 (N_27903,N_24788,N_24502);
or U27904 (N_27904,N_25871,N_24401);
or U27905 (N_27905,N_25553,N_24949);
xnor U27906 (N_27906,N_25027,N_25755);
and U27907 (N_27907,N_24228,N_25296);
nand U27908 (N_27908,N_25971,N_24291);
xnor U27909 (N_27909,N_25811,N_25046);
nand U27910 (N_27910,N_25312,N_25051);
and U27911 (N_27911,N_25818,N_24153);
xnor U27912 (N_27912,N_24316,N_24838);
nand U27913 (N_27913,N_24043,N_24386);
xnor U27914 (N_27914,N_25500,N_25576);
or U27915 (N_27915,N_24317,N_24344);
nor U27916 (N_27916,N_24741,N_25324);
xnor U27917 (N_27917,N_25921,N_25146);
and U27918 (N_27918,N_24778,N_24722);
nand U27919 (N_27919,N_24257,N_24539);
or U27920 (N_27920,N_24494,N_24796);
and U27921 (N_27921,N_25821,N_25020);
nor U27922 (N_27922,N_25138,N_24769);
and U27923 (N_27923,N_24062,N_24534);
nand U27924 (N_27924,N_24978,N_24039);
or U27925 (N_27925,N_24023,N_24907);
nand U27926 (N_27926,N_24570,N_24455);
xor U27927 (N_27927,N_25021,N_25111);
nand U27928 (N_27928,N_24272,N_24884);
nor U27929 (N_27929,N_24357,N_25475);
nand U27930 (N_27930,N_24875,N_25878);
and U27931 (N_27931,N_24045,N_25101);
nor U27932 (N_27932,N_24091,N_25217);
xor U27933 (N_27933,N_25420,N_24020);
and U27934 (N_27934,N_24685,N_24622);
or U27935 (N_27935,N_25997,N_24289);
xnor U27936 (N_27936,N_25363,N_25728);
nand U27937 (N_27937,N_24173,N_24588);
nor U27938 (N_27938,N_25849,N_25948);
and U27939 (N_27939,N_24964,N_24135);
and U27940 (N_27940,N_24624,N_25860);
nor U27941 (N_27941,N_25298,N_25774);
or U27942 (N_27942,N_25071,N_24888);
xnor U27943 (N_27943,N_24122,N_25581);
xor U27944 (N_27944,N_25651,N_25066);
and U27945 (N_27945,N_25598,N_25484);
nand U27946 (N_27946,N_24186,N_24365);
and U27947 (N_27947,N_24280,N_24035);
nor U27948 (N_27948,N_25941,N_25914);
xor U27949 (N_27949,N_25769,N_24108);
and U27950 (N_27950,N_25169,N_25893);
xor U27951 (N_27951,N_24969,N_25868);
nand U27952 (N_27952,N_24383,N_25647);
or U27953 (N_27953,N_25211,N_25018);
nand U27954 (N_27954,N_24935,N_25836);
nor U27955 (N_27955,N_25437,N_24516);
and U27956 (N_27956,N_24000,N_24911);
and U27957 (N_27957,N_24004,N_24219);
or U27958 (N_27958,N_24000,N_24228);
nor U27959 (N_27959,N_24273,N_25137);
or U27960 (N_27960,N_24597,N_25083);
nor U27961 (N_27961,N_25931,N_24632);
nand U27962 (N_27962,N_25572,N_24988);
xnor U27963 (N_27963,N_25119,N_24918);
xor U27964 (N_27964,N_24559,N_25770);
nand U27965 (N_27965,N_24708,N_25455);
nand U27966 (N_27966,N_25004,N_24211);
nor U27967 (N_27967,N_24721,N_25780);
or U27968 (N_27968,N_25678,N_24897);
nand U27969 (N_27969,N_24439,N_24976);
nor U27970 (N_27970,N_24088,N_25208);
and U27971 (N_27971,N_25597,N_25241);
or U27972 (N_27972,N_25479,N_25748);
and U27973 (N_27973,N_24025,N_24548);
xnor U27974 (N_27974,N_25710,N_25489);
or U27975 (N_27975,N_24497,N_25791);
or U27976 (N_27976,N_24470,N_24384);
and U27977 (N_27977,N_25898,N_25855);
xnor U27978 (N_27978,N_25561,N_25310);
nor U27979 (N_27979,N_24752,N_24120);
or U27980 (N_27980,N_25402,N_25365);
xor U27981 (N_27981,N_25026,N_25091);
or U27982 (N_27982,N_25308,N_25840);
nand U27983 (N_27983,N_24401,N_25729);
nor U27984 (N_27984,N_24189,N_24894);
and U27985 (N_27985,N_25101,N_25910);
nor U27986 (N_27986,N_25194,N_24806);
xnor U27987 (N_27987,N_25409,N_25634);
nor U27988 (N_27988,N_24163,N_25945);
xor U27989 (N_27989,N_24658,N_25065);
nor U27990 (N_27990,N_24868,N_25577);
nand U27991 (N_27991,N_24160,N_24186);
and U27992 (N_27992,N_24419,N_24338);
and U27993 (N_27993,N_24271,N_25854);
or U27994 (N_27994,N_24687,N_24368);
nand U27995 (N_27995,N_25929,N_25576);
or U27996 (N_27996,N_24375,N_24141);
and U27997 (N_27997,N_24141,N_25397);
and U27998 (N_27998,N_24807,N_24880);
nor U27999 (N_27999,N_24239,N_24549);
and U28000 (N_28000,N_27451,N_26322);
nand U28001 (N_28001,N_26694,N_27550);
xor U28002 (N_28002,N_26085,N_27095);
nand U28003 (N_28003,N_27864,N_26363);
nand U28004 (N_28004,N_26937,N_27184);
nand U28005 (N_28005,N_26433,N_27420);
nor U28006 (N_28006,N_27945,N_27037);
and U28007 (N_28007,N_26313,N_27390);
nor U28008 (N_28008,N_27499,N_27595);
or U28009 (N_28009,N_26421,N_27818);
and U28010 (N_28010,N_27255,N_27099);
and U28011 (N_28011,N_27188,N_27944);
and U28012 (N_28012,N_26632,N_26470);
xor U28013 (N_28013,N_27040,N_26951);
nor U28014 (N_28014,N_27544,N_26780);
or U28015 (N_28015,N_26436,N_27872);
or U28016 (N_28016,N_26591,N_26958);
nand U28017 (N_28017,N_26430,N_27924);
xor U28018 (N_28018,N_26525,N_26760);
nor U28019 (N_28019,N_27505,N_26651);
nor U28020 (N_28020,N_26731,N_27498);
nor U28021 (N_28021,N_27116,N_26557);
xnor U28022 (N_28022,N_26110,N_26296);
nor U28023 (N_28023,N_26494,N_26209);
and U28024 (N_28024,N_26747,N_27738);
xor U28025 (N_28025,N_27190,N_26443);
or U28026 (N_28026,N_27983,N_27667);
nand U28027 (N_28027,N_26946,N_27853);
and U28028 (N_28028,N_27512,N_26208);
nor U28029 (N_28029,N_27982,N_26096);
nor U28030 (N_28030,N_26415,N_27039);
nand U28031 (N_28031,N_27584,N_26440);
or U28032 (N_28032,N_27901,N_26424);
and U28033 (N_28033,N_26051,N_27735);
xnor U28034 (N_28034,N_26707,N_27626);
nor U28035 (N_28035,N_27311,N_26770);
nor U28036 (N_28036,N_27699,N_27091);
or U28037 (N_28037,N_27297,N_27830);
nor U28038 (N_28038,N_27434,N_27432);
xnor U28039 (N_28039,N_27612,N_26510);
nor U28040 (N_28040,N_26699,N_26933);
nor U28041 (N_28041,N_27133,N_26175);
nor U28042 (N_28042,N_26767,N_27881);
xor U28043 (N_28043,N_27618,N_26043);
nor U28044 (N_28044,N_26716,N_27600);
and U28045 (N_28045,N_26092,N_26144);
nor U28046 (N_28046,N_26463,N_27663);
xnor U28047 (N_28047,N_26272,N_27679);
xor U28048 (N_28048,N_26864,N_26812);
nor U28049 (N_28049,N_26220,N_27791);
and U28050 (N_28050,N_26396,N_27737);
nor U28051 (N_28051,N_27020,N_26585);
and U28052 (N_28052,N_27340,N_27166);
xnor U28053 (N_28053,N_26229,N_27442);
xor U28054 (N_28054,N_27624,N_26969);
nand U28055 (N_28055,N_26180,N_26703);
xnor U28056 (N_28056,N_26631,N_27856);
and U28057 (N_28057,N_27517,N_26364);
xnor U28058 (N_28058,N_27752,N_27363);
xnor U28059 (N_28059,N_27633,N_27168);
nand U28060 (N_28060,N_26537,N_27024);
nor U28061 (N_28061,N_27873,N_26513);
or U28062 (N_28062,N_26927,N_26761);
nor U28063 (N_28063,N_27790,N_27497);
and U28064 (N_28064,N_26349,N_27829);
nor U28065 (N_28065,N_27060,N_26369);
xor U28066 (N_28066,N_26331,N_26682);
or U28067 (N_28067,N_27777,N_27565);
nor U28068 (N_28068,N_27963,N_27046);
or U28069 (N_28069,N_26393,N_26603);
or U28070 (N_28070,N_27545,N_27378);
nand U28071 (N_28071,N_27716,N_26615);
nand U28072 (N_28072,N_26750,N_27126);
nor U28073 (N_28073,N_26517,N_26612);
nand U28074 (N_28074,N_27660,N_27770);
or U28075 (N_28075,N_26875,N_26530);
nand U28076 (N_28076,N_26552,N_26865);
nand U28077 (N_28077,N_27939,N_26098);
nor U28078 (N_28078,N_27987,N_27478);
or U28079 (N_28079,N_26904,N_26219);
or U28080 (N_28080,N_27823,N_27365);
and U28081 (N_28081,N_27071,N_27984);
or U28082 (N_28082,N_27842,N_26057);
nand U28083 (N_28083,N_26045,N_26811);
nor U28084 (N_28084,N_27110,N_26497);
and U28085 (N_28085,N_26995,N_27609);
or U28086 (N_28086,N_26006,N_27892);
nand U28087 (N_28087,N_27414,N_27507);
nor U28088 (N_28088,N_26339,N_27286);
nand U28089 (N_28089,N_27681,N_27713);
xor U28090 (N_28090,N_26056,N_27635);
nor U28091 (N_28091,N_26214,N_26920);
or U28092 (N_28092,N_26985,N_26000);
nand U28093 (N_28093,N_27324,N_27468);
and U28094 (N_28094,N_27602,N_27177);
xor U28095 (N_28095,N_26225,N_26885);
or U28096 (N_28096,N_26926,N_26425);
or U28097 (N_28097,N_26599,N_27495);
and U28098 (N_28098,N_27366,N_26554);
xor U28099 (N_28099,N_26858,N_26207);
nand U28100 (N_28100,N_27292,N_27005);
nor U28101 (N_28101,N_27561,N_27100);
xnor U28102 (N_28102,N_27249,N_27433);
or U28103 (N_28103,N_26142,N_27016);
nor U28104 (N_28104,N_26534,N_27440);
and U28105 (N_28105,N_27923,N_26127);
nand U28106 (N_28106,N_27483,N_27233);
or U28107 (N_28107,N_27796,N_26261);
xor U28108 (N_28108,N_26444,N_27801);
xor U28109 (N_28109,N_26779,N_27774);
nor U28110 (N_28110,N_26674,N_27004);
xnor U28111 (N_28111,N_27562,N_27794);
nor U28112 (N_28112,N_26492,N_27396);
xnor U28113 (N_28113,N_27488,N_27840);
nor U28114 (N_28114,N_27530,N_27920);
xor U28115 (N_28115,N_26499,N_27282);
xor U28116 (N_28116,N_26792,N_26724);
xnor U28117 (N_28117,N_26059,N_26233);
and U28118 (N_28118,N_26107,N_26873);
and U28119 (N_28119,N_26439,N_27997);
nor U28120 (N_28120,N_26186,N_26447);
nor U28121 (N_28121,N_27410,N_26783);
xor U28122 (N_28122,N_27090,N_27041);
nand U28123 (N_28123,N_26341,N_26485);
nor U28124 (N_28124,N_26660,N_26388);
nand U28125 (N_28125,N_26979,N_27094);
nor U28126 (N_28126,N_27083,N_27405);
or U28127 (N_28127,N_27586,N_26519);
or U28128 (N_28128,N_27548,N_27583);
nor U28129 (N_28129,N_26224,N_27136);
nand U28130 (N_28130,N_26738,N_26104);
xnor U28131 (N_28131,N_27568,N_26125);
and U28132 (N_28132,N_27272,N_26505);
xnor U28133 (N_28133,N_26155,N_26457);
and U28134 (N_28134,N_26931,N_27025);
nor U28135 (N_28135,N_27620,N_26159);
nor U28136 (N_28136,N_26973,N_27228);
and U28137 (N_28137,N_27714,N_27192);
nand U28138 (N_28138,N_27551,N_26071);
xnor U28139 (N_28139,N_26165,N_26515);
nor U28140 (N_28140,N_26966,N_27865);
and U28141 (N_28141,N_27514,N_26735);
or U28142 (N_28142,N_27021,N_27002);
xnor U28143 (N_28143,N_26283,N_27310);
xor U28144 (N_28144,N_27211,N_26422);
and U28145 (N_28145,N_26702,N_26355);
or U28146 (N_28146,N_27811,N_27597);
xnor U28147 (N_28147,N_27700,N_26857);
nor U28148 (N_28148,N_26484,N_26638);
xnor U28149 (N_28149,N_27274,N_27809);
nor U28150 (N_28150,N_27773,N_26223);
nor U28151 (N_28151,N_26498,N_27447);
nand U28152 (N_28152,N_27367,N_26136);
and U28153 (N_28153,N_27156,N_26662);
xnor U28154 (N_28154,N_27320,N_27081);
xor U28155 (N_28155,N_26265,N_26807);
or U28156 (N_28156,N_26238,N_26458);
and U28157 (N_28157,N_27910,N_26902);
xor U28158 (N_28158,N_27869,N_27135);
nor U28159 (N_28159,N_26828,N_26482);
nand U28160 (N_28160,N_27788,N_26550);
nand U28161 (N_28161,N_26459,N_27105);
nand U28162 (N_28162,N_27132,N_27585);
or U28163 (N_28163,N_26883,N_27740);
and U28164 (N_28164,N_27208,N_26370);
nand U28165 (N_28165,N_27558,N_26996);
nor U28166 (N_28166,N_26500,N_27392);
or U28167 (N_28167,N_27375,N_27914);
nor U28168 (N_28168,N_26733,N_26154);
and U28169 (N_28169,N_26236,N_27833);
nand U28170 (N_28170,N_26167,N_27837);
and U28171 (N_28171,N_27121,N_26390);
xnor U28172 (N_28172,N_27117,N_26001);
and U28173 (N_28173,N_26614,N_27106);
or U28174 (N_28174,N_26262,N_27569);
xor U28175 (N_28175,N_26917,N_27129);
nor U28176 (N_28176,N_27294,N_27336);
xor U28177 (N_28177,N_27382,N_27130);
nand U28178 (N_28178,N_26976,N_26601);
nand U28179 (N_28179,N_26205,N_26289);
xor U28180 (N_28180,N_27769,N_26479);
nand U28181 (N_28181,N_26894,N_27250);
nand U28182 (N_28182,N_26846,N_27131);
or U28183 (N_28183,N_26508,N_26011);
nand U28184 (N_28184,N_27931,N_27425);
and U28185 (N_28185,N_27623,N_27921);
nor U28186 (N_28186,N_27812,N_26670);
and U28187 (N_28187,N_26771,N_26356);
nor U28188 (N_28188,N_26570,N_27338);
or U28189 (N_28189,N_26778,N_27902);
nand U28190 (N_28190,N_27076,N_26897);
xor U28191 (N_28191,N_27466,N_26970);
or U28192 (N_28192,N_27238,N_26252);
xnor U28193 (N_28193,N_26950,N_27759);
nor U28194 (N_28194,N_27330,N_27061);
nand U28195 (N_28195,N_27026,N_27372);
nand U28196 (N_28196,N_27143,N_27628);
nand U28197 (N_28197,N_27846,N_26183);
or U28198 (N_28198,N_26757,N_27523);
nand U28199 (N_28199,N_26354,N_27707);
xnor U28200 (N_28200,N_26898,N_26541);
nor U28201 (N_28201,N_26571,N_26122);
nor U28202 (N_28202,N_27528,N_26343);
and U28203 (N_28203,N_27047,N_27243);
nor U28204 (N_28204,N_26791,N_27161);
nand U28205 (N_28205,N_27154,N_27269);
xor U28206 (N_28206,N_27147,N_27401);
and U28207 (N_28207,N_27043,N_27891);
or U28208 (N_28208,N_27280,N_27947);
and U28209 (N_28209,N_26055,N_26816);
nor U28210 (N_28210,N_26376,N_26799);
or U28211 (N_28211,N_27832,N_27056);
nand U28212 (N_28212,N_27315,N_27825);
or U28213 (N_28213,N_27761,N_27955);
nand U28214 (N_28214,N_27539,N_27848);
or U28215 (N_28215,N_26473,N_27219);
or U28216 (N_28216,N_26764,N_26823);
and U28217 (N_28217,N_26910,N_27671);
or U28218 (N_28218,N_27141,N_27547);
nand U28219 (N_28219,N_27867,N_26914);
nor U28220 (N_28220,N_26989,N_27408);
and U28221 (N_28221,N_27151,N_26407);
nor U28222 (N_28222,N_26701,N_26299);
or U28223 (N_28223,N_27651,N_26793);
xor U28224 (N_28224,N_27974,N_26972);
xnor U28225 (N_28225,N_27072,N_26635);
nand U28226 (N_28226,N_26467,N_26187);
xor U28227 (N_28227,N_26477,N_26414);
nor U28228 (N_28228,N_26538,N_26290);
xor U28229 (N_28229,N_27319,N_27746);
nor U28230 (N_28230,N_27463,N_26768);
xnor U28231 (N_28231,N_26560,N_26986);
and U28232 (N_28232,N_26244,N_27698);
nand U28233 (N_28233,N_27167,N_27464);
xor U28234 (N_28234,N_27007,N_26622);
and U28235 (N_28235,N_27666,N_27937);
and U28236 (N_28236,N_26941,N_26604);
nor U28237 (N_28237,N_27265,N_27082);
xnor U28238 (N_28238,N_26901,N_26395);
nor U28239 (N_28239,N_26113,N_27430);
or U28240 (N_28240,N_26271,N_27419);
nand U28241 (N_28241,N_27975,N_26173);
and U28242 (N_28242,N_27875,N_27234);
or U28243 (N_28243,N_27127,N_27959);
and U28244 (N_28244,N_26545,N_27028);
nor U28245 (N_28245,N_27764,N_26474);
nor U28246 (N_28246,N_27019,N_27075);
and U28247 (N_28247,N_26661,N_26139);
nand U28248 (N_28248,N_27101,N_27178);
nand U28249 (N_28249,N_26629,N_27515);
and U28250 (N_28250,N_26551,N_26977);
xnor U28251 (N_28251,N_26052,N_27938);
and U28252 (N_28252,N_26714,N_26041);
or U28253 (N_28253,N_27789,N_26608);
nor U28254 (N_28254,N_26956,N_26520);
nor U28255 (N_28255,N_26833,N_27346);
nand U28256 (N_28256,N_27221,N_27854);
nor U28257 (N_28257,N_27510,N_26569);
or U28258 (N_28258,N_26908,N_26023);
or U28259 (N_28259,N_27058,N_27631);
and U28260 (N_28260,N_27915,N_26678);
nor U28261 (N_28261,N_26297,N_26621);
and U28262 (N_28262,N_27760,N_27461);
xnor U28263 (N_28263,N_27073,N_26636);
and U28264 (N_28264,N_26679,N_26563);
nor U28265 (N_28265,N_27306,N_26624);
xor U28266 (N_28266,N_27971,N_26086);
and U28267 (N_28267,N_26751,N_26247);
and U28268 (N_28268,N_26382,N_27500);
and U28269 (N_28269,N_26308,N_26063);
or U28270 (N_28270,N_27819,N_27018);
or U28271 (N_28271,N_27560,N_27240);
nand U28272 (N_28272,N_26143,N_26533);
and U28273 (N_28273,N_26392,N_26556);
or U28274 (N_28274,N_26192,N_26486);
nand U28275 (N_28275,N_27493,N_27749);
and U28276 (N_28276,N_27590,N_27446);
or U28277 (N_28277,N_26021,N_27617);
or U28278 (N_28278,N_27036,N_26184);
xor U28279 (N_28279,N_27772,N_27202);
nand U28280 (N_28280,N_27150,N_26460);
or U28281 (N_28281,N_27383,N_26166);
nand U28282 (N_28282,N_26562,N_27653);
nand U28283 (N_28283,N_27606,N_26020);
or U28284 (N_28284,N_26705,N_26665);
xor U28285 (N_28285,N_27448,N_27031);
xor U28286 (N_28286,N_26350,N_26212);
nor U28287 (N_28287,N_27538,N_27407);
or U28288 (N_28288,N_27756,N_26344);
nor U28289 (N_28289,N_27035,N_27262);
nor U28290 (N_28290,N_27077,N_26118);
and U28291 (N_28291,N_26836,N_26069);
or U28292 (N_28292,N_27727,N_26254);
or U28293 (N_28293,N_27122,N_27967);
nor U28294 (N_28294,N_27525,N_26060);
or U28295 (N_28295,N_26548,N_26531);
or U28296 (N_28296,N_27137,N_27899);
or U28297 (N_28297,N_27103,N_26025);
nor U28298 (N_28298,N_27844,N_26991);
nor U28299 (N_28299,N_27828,N_26964);
and U28300 (N_28300,N_26191,N_27946);
xor U28301 (N_28301,N_27256,N_26790);
and U28302 (N_28302,N_26347,N_27387);
nand U28303 (N_28303,N_26162,N_26945);
xnor U28304 (N_28304,N_27301,N_26925);
xnor U28305 (N_28305,N_26275,N_27710);
and U28306 (N_28306,N_27787,N_27755);
nor U28307 (N_28307,N_26955,N_27153);
nand U28308 (N_28308,N_27010,N_27180);
xor U28309 (N_28309,N_26137,N_26961);
or U28310 (N_28310,N_27332,N_27919);
and U28311 (N_28311,N_26853,N_27098);
or U28312 (N_28312,N_26365,N_26772);
nand U28313 (N_28313,N_27717,N_27456);
and U28314 (N_28314,N_26423,N_27496);
nand U28315 (N_28315,N_27765,N_26765);
and U28316 (N_28316,N_27348,N_26709);
nor U28317 (N_28317,N_26659,N_26366);
xor U28318 (N_28318,N_27403,N_26642);
xor U28319 (N_28319,N_26867,N_27996);
xnor U28320 (N_28320,N_26361,N_27339);
nand U28321 (N_28321,N_27044,N_26164);
and U28322 (N_28322,N_27352,N_27596);
xnor U28323 (N_28323,N_27278,N_27647);
nor U28324 (N_28324,N_26801,N_26687);
xor U28325 (N_28325,N_27033,N_26116);
nand U28326 (N_28326,N_27397,N_27066);
and U28327 (N_28327,N_27251,N_26639);
nand U28328 (N_28328,N_26911,N_27267);
and U28329 (N_28329,N_26708,N_26524);
xor U28330 (N_28330,N_26685,N_27976);
nand U28331 (N_28331,N_27785,N_26481);
nand U28332 (N_28332,N_26826,N_26417);
nor U28333 (N_28333,N_27798,N_27692);
and U28334 (N_28334,N_27260,N_27157);
xor U28335 (N_28335,N_27501,N_27943);
or U28336 (N_28336,N_26256,N_27344);
and U28337 (N_28337,N_27013,N_26362);
nand U28338 (N_28338,N_27855,N_26882);
or U28339 (N_28339,N_26786,N_26371);
xor U28340 (N_28340,N_27664,N_26013);
and U28341 (N_28341,N_26400,N_26692);
xor U28342 (N_28342,N_27201,N_26321);
nand U28343 (N_28343,N_26586,N_26960);
and U28344 (N_28344,N_27231,N_27629);
and U28345 (N_28345,N_27406,N_26215);
nor U28346 (N_28346,N_26762,N_27068);
or U28347 (N_28347,N_26597,N_27490);
nand U28348 (N_28348,N_26856,N_26564);
xor U28349 (N_28349,N_26402,N_26048);
nand U28350 (N_28350,N_26487,N_26928);
xnor U28351 (N_28351,N_27815,N_26711);
and U28352 (N_28352,N_26269,N_26704);
xor U28353 (N_28353,N_26461,N_27171);
and U28354 (N_28354,N_27309,N_27045);
or U28355 (N_28355,N_26146,N_26311);
and U28356 (N_28356,N_27549,N_27668);
nand U28357 (N_28357,N_26042,N_27793);
nor U28358 (N_28358,N_27702,N_26516);
and U28359 (N_28359,N_26044,N_27563);
or U28360 (N_28360,N_26452,N_27334);
xor U28361 (N_28361,N_27128,N_26938);
xor U28362 (N_28362,N_27017,N_26633);
xnor U28363 (N_28363,N_26903,N_27032);
nand U28364 (N_28364,N_26197,N_26234);
nor U28365 (N_28365,N_27688,N_27655);
xnor U28366 (N_28366,N_26610,N_26583);
nor U28367 (N_28367,N_27476,N_26835);
nor U28368 (N_28368,N_27246,N_26844);
nor U28369 (N_28369,N_26346,N_26849);
nand U28370 (N_28370,N_26932,N_27841);
nand U28371 (N_28371,N_26666,N_26231);
and U28372 (N_28372,N_26884,N_27908);
xor U28373 (N_28373,N_27443,N_26009);
or U28374 (N_28374,N_26243,N_26005);
nand U28375 (N_28375,N_27198,N_26553);
or U28376 (N_28376,N_27593,N_27200);
and U28377 (N_28377,N_27989,N_26766);
or U28378 (N_28378,N_26909,N_26386);
and U28379 (N_28379,N_26158,N_26426);
xor U28380 (N_28380,N_27729,N_26198);
and U28381 (N_28381,N_26605,N_26302);
nand U28382 (N_28382,N_26852,N_26859);
xor U28383 (N_28383,N_27680,N_26333);
nand U28384 (N_28384,N_27465,N_26404);
xor U28385 (N_28385,N_26522,N_26310);
and U28386 (N_28386,N_27070,N_27564);
and U28387 (N_28387,N_26948,N_26352);
nor U28388 (N_28388,N_27162,N_27285);
and U28389 (N_28389,N_27535,N_26129);
nor U28390 (N_28390,N_26834,N_27380);
xnor U28391 (N_28391,N_26451,N_26874);
or U28392 (N_28392,N_27532,N_26646);
xnor U28393 (N_28393,N_26869,N_26468);
xor U28394 (N_28394,N_26230,N_27395);
nand U28395 (N_28395,N_26758,N_27588);
or U28396 (N_28396,N_27196,N_27369);
nor U28397 (N_28397,N_27592,N_27754);
nor U28398 (N_28398,N_27429,N_27927);
and U28399 (N_28399,N_27067,N_27308);
nor U28400 (N_28400,N_27988,N_26843);
xor U28401 (N_28401,N_27086,N_27723);
nor U28402 (N_28402,N_26070,N_27325);
nor U28403 (N_28403,N_27907,N_26030);
nand U28404 (N_28404,N_26743,N_27942);
nand U28405 (N_28405,N_26734,N_26115);
or U28406 (N_28406,N_26035,N_26915);
xor U28407 (N_28407,N_27870,N_27731);
and U28408 (N_28408,N_26745,N_26962);
and U28409 (N_28409,N_26282,N_26181);
nor U28410 (N_28410,N_27480,N_27805);
or U28411 (N_28411,N_26157,N_27916);
xor U28412 (N_28412,N_27102,N_26871);
and U28413 (N_28413,N_26300,N_26432);
nand U28414 (N_28414,N_26334,N_27062);
nand U28415 (N_28415,N_27437,N_26002);
and U28416 (N_28416,N_26434,N_26291);
nor U28417 (N_28417,N_27889,N_27165);
nand U28418 (N_28418,N_27054,N_27268);
xor U28419 (N_28419,N_26540,N_27107);
or U28420 (N_28420,N_27199,N_26431);
xor U28421 (N_28421,N_27566,N_27925);
nand U28422 (N_28422,N_26942,N_26377);
or U28423 (N_28423,N_26528,N_26547);
nor U28424 (N_28424,N_27096,N_27802);
nand U28425 (N_28425,N_26076,N_26145);
or U28426 (N_28426,N_27720,N_27615);
and U28427 (N_28427,N_26940,N_27894);
nand U28428 (N_28428,N_26640,N_26566);
nand U28429 (N_28429,N_27636,N_26637);
nand U28430 (N_28430,N_26881,N_26891);
nand U28431 (N_28431,N_26890,N_26304);
nor U28432 (N_28432,N_27264,N_26161);
nand U28433 (N_28433,N_26373,N_26831);
and U28434 (N_28434,N_26729,N_27784);
and U28435 (N_28435,N_27935,N_26993);
nand U28436 (N_28436,N_27415,N_26172);
nor U28437 (N_28437,N_27640,N_27504);
and U28438 (N_28438,N_26128,N_26489);
xor U28439 (N_28439,N_27457,N_26698);
xnor U28440 (N_28440,N_27775,N_27650);
nand U28441 (N_28441,N_27694,N_27423);
xnor U28442 (N_28442,N_26987,N_26575);
and U28443 (N_28443,N_27085,N_27581);
or U28444 (N_28444,N_27678,N_27730);
and U28445 (N_28445,N_27783,N_26453);
nor U28446 (N_28446,N_27516,N_26980);
nand U28447 (N_28447,N_27404,N_27299);
xor U28448 (N_28448,N_27259,N_27413);
xor U28449 (N_28449,N_27814,N_26316);
or U28450 (N_28450,N_26007,N_27176);
or U28451 (N_28451,N_26700,N_26267);
and U28452 (N_28452,N_26824,N_27999);
and U28453 (N_28453,N_26217,N_27424);
xnor U28454 (N_28454,N_27574,N_27155);
nand U28455 (N_28455,N_27470,N_26188);
and U28456 (N_28456,N_27722,N_26878);
or U28457 (N_28457,N_27797,N_26706);
or U28458 (N_28458,N_27537,N_26285);
and U28459 (N_28459,N_26880,N_26886);
or U28460 (N_28460,N_26804,N_27236);
nand U28461 (N_28461,N_27485,N_26131);
or U28462 (N_28462,N_26102,N_26755);
nor U28463 (N_28463,N_27627,N_26815);
or U28464 (N_28464,N_27934,N_27768);
nor U28465 (N_28465,N_26036,N_26509);
nand U28466 (N_28466,N_27642,N_26133);
nor U28467 (N_28467,N_26740,N_26527);
and U28468 (N_28468,N_26323,N_27972);
nor U28469 (N_28469,N_26596,N_26837);
nor U28470 (N_28470,N_27863,N_27683);
or U28471 (N_28471,N_27993,N_27006);
xor U28472 (N_28472,N_26465,N_27994);
nor U28473 (N_28473,N_26669,N_26776);
nor U28474 (N_28474,N_26163,N_27522);
or U28475 (N_28475,N_27092,N_26024);
or U28476 (N_28476,N_27933,N_27486);
nor U28477 (N_28477,N_27318,N_26084);
nand U28478 (N_28478,N_27771,N_26822);
nor U28479 (N_28479,N_27347,N_27649);
nor U28480 (N_28480,N_26016,N_26620);
nor U28481 (N_28481,N_26213,N_26710);
nand U28482 (N_28482,N_26809,N_27123);
or U28483 (N_28483,N_27567,N_27209);
and U28484 (N_28484,N_26368,N_26561);
or U28485 (N_28485,N_26190,N_26978);
and U28486 (N_28486,N_27069,N_26658);
nand U28487 (N_28487,N_26312,N_27521);
and U28488 (N_28488,N_26337,N_27816);
xnor U28489 (N_28489,N_26462,N_26454);
nand U28490 (N_28490,N_26242,N_26105);
nor U28491 (N_28491,N_26268,N_26120);
and U28492 (N_28492,N_27217,N_27850);
and U28493 (N_28493,N_27824,N_26775);
nor U28494 (N_28494,N_27589,N_26934);
and U28495 (N_28495,N_27529,N_26691);
xnor U28496 (N_28496,N_27810,N_27619);
and U28497 (N_28497,N_27445,N_26730);
nand U28498 (N_28498,N_27244,N_27956);
or U28499 (N_28499,N_27489,N_27290);
nand U28500 (N_28500,N_26029,N_26464);
xnor U28501 (N_28501,N_26542,N_27630);
or U28502 (N_28502,N_27140,N_27641);
nor U28503 (N_28503,N_27822,N_27441);
and U28504 (N_28504,N_27985,N_27898);
and U28505 (N_28505,N_27661,N_26359);
xor U28506 (N_28506,N_26838,N_26054);
or U28507 (N_28507,N_27323,N_27582);
nor U28508 (N_28508,N_27333,N_27374);
nor U28509 (N_28509,N_26251,N_27422);
nor U28510 (N_28510,N_27859,N_26012);
nand U28511 (N_28511,N_27603,N_26568);
nor U28512 (N_28512,N_27218,N_27479);
and U28513 (N_28513,N_26854,N_26263);
and U28514 (N_28514,N_27053,N_27471);
nor U28515 (N_28515,N_27360,N_26412);
nor U28516 (N_28516,N_26655,N_27232);
or U28517 (N_28517,N_27050,N_26039);
and U28518 (N_28518,N_27453,N_27358);
or U28519 (N_28519,N_26739,N_26073);
and U28520 (N_28520,N_27598,N_27475);
nor U28521 (N_28521,N_26336,N_26672);
and U28522 (N_28522,N_27962,N_26046);
xnor U28523 (N_28523,N_26315,N_27029);
nand U28524 (N_28524,N_26360,N_26478);
and U28525 (N_28525,N_27049,N_27242);
xor U28526 (N_28526,N_27652,N_26889);
xnor U28527 (N_28527,N_27492,N_27743);
or U28528 (N_28528,N_27377,N_26502);
and U28529 (N_28529,N_26003,N_27871);
and U28530 (N_28530,N_26375,N_27109);
and U28531 (N_28531,N_27173,N_26957);
nor U28532 (N_28532,N_26749,N_27146);
xor U28533 (N_28533,N_27543,N_26851);
or U28534 (N_28534,N_26781,N_26090);
nand U28535 (N_28535,N_27271,N_27351);
and U28536 (N_28536,N_27546,N_26328);
xnor U28537 (N_28537,N_26803,N_27065);
xor U28538 (N_28538,N_27861,N_27838);
or U28539 (N_28539,N_27115,N_26279);
nand U28540 (N_28540,N_27860,N_26839);
nand U28541 (N_28541,N_27876,N_27302);
nor U28542 (N_28542,N_27701,N_26982);
and U28543 (N_28543,N_26967,N_26171);
nor U28544 (N_28544,N_27473,N_26959);
nor U28545 (N_28545,N_26255,N_26984);
nand U28546 (N_28546,N_26936,N_26318);
nand U28547 (N_28547,N_27313,N_27940);
nor U28548 (N_28548,N_26626,N_27736);
or U28549 (N_28549,N_26680,N_26182);
nor U28550 (N_28550,N_26345,N_27911);
or U28551 (N_28551,N_27273,N_26543);
xnor U28552 (N_28552,N_26589,N_27181);
nand U28553 (N_28553,N_26744,N_27185);
nand U28554 (N_28554,N_26018,N_26994);
or U28555 (N_28555,N_27462,N_26820);
or U28556 (N_28556,N_27051,N_26195);
nor U28557 (N_28557,N_27594,N_27638);
xor U28558 (N_28558,N_26990,N_27534);
nor U28559 (N_28559,N_27158,N_27703);
nand U28560 (N_28560,N_26442,N_26712);
nor U28561 (N_28561,N_26286,N_27089);
and U28562 (N_28562,N_27317,N_26472);
xor U28563 (N_28563,N_27125,N_26893);
and U28564 (N_28564,N_26949,N_26095);
nand U28565 (N_28565,N_27957,N_26868);
nor U28566 (N_28566,N_27682,N_27469);
nand U28567 (N_28567,N_26998,N_26913);
nor U28568 (N_28568,N_27163,N_26916);
nand U28569 (N_28569,N_26523,N_26789);
nand U28570 (N_28570,N_27421,N_26860);
xor U28571 (N_28571,N_26935,N_26032);
xnor U28572 (N_28572,N_26602,N_26132);
xor U28573 (N_28573,N_27477,N_26004);
nor U28574 (N_28574,N_27227,N_26794);
and U28575 (N_28575,N_27675,N_26121);
xnor U28576 (N_28576,N_27733,N_27291);
or U28577 (N_28577,N_26080,N_26419);
nor U28578 (N_28578,N_27857,N_26576);
nand U28579 (N_28579,N_26257,N_26306);
and U28580 (N_28580,N_27426,N_27326);
xor U28581 (N_28581,N_26097,N_27148);
xor U28582 (N_28582,N_27757,N_27964);
xor U28583 (N_28583,N_27275,N_26693);
nor U28584 (N_28584,N_26899,N_27454);
nor U28585 (N_28585,N_27966,N_27444);
nor U28586 (N_28586,N_27969,N_27487);
nor U28587 (N_28587,N_27063,N_27930);
or U28588 (N_28588,N_26715,N_26773);
nand U28589 (N_28589,N_26249,N_27079);
or U28590 (N_28590,N_26429,N_26968);
nand U28591 (N_28591,N_26152,N_26253);
nor U28592 (N_28592,N_27038,N_27718);
and U28593 (N_28593,N_26999,N_27646);
or U28594 (N_28594,N_27287,N_27741);
nor U28595 (N_28595,N_26332,N_27393);
xor U28596 (N_28596,N_27834,N_27929);
nor U28597 (N_28597,N_26841,N_26536);
nand U28598 (N_28598,N_26677,N_27526);
nand U28599 (N_28599,N_27254,N_27000);
nand U28600 (N_28600,N_27918,N_27747);
and U28601 (N_28601,N_27684,N_26469);
or U28602 (N_28602,N_27527,N_26870);
xnor U28603 (N_28603,N_26319,N_26420);
nand U28604 (N_28604,N_27175,N_27482);
xor U28605 (N_28605,N_27762,N_26277);
or U28606 (N_28606,N_27665,N_26848);
or U28607 (N_28607,N_26153,N_26038);
nor U28608 (N_28608,N_27506,N_27831);
nor U28609 (N_28609,N_26293,N_26695);
xor U28610 (N_28610,N_27893,N_27961);
nor U28611 (N_28611,N_26546,N_27928);
and U28612 (N_28612,N_27048,N_27885);
or U28613 (N_28613,N_26618,N_27977);
nand U28614 (N_28614,N_27370,N_26455);
nor U28615 (N_28615,N_26549,N_26221);
nor U28616 (N_28616,N_27973,N_26061);
or U28617 (N_28617,N_26065,N_26109);
and U28618 (N_28618,N_26174,N_27239);
nand U28619 (N_28619,N_26123,N_27342);
and U28620 (N_28620,N_27843,N_26567);
nor U28621 (N_28621,N_26559,N_27542);
nand U28622 (N_28622,N_27182,N_27362);
nand U28623 (N_28623,N_26441,N_26921);
xnor U28624 (N_28624,N_26717,N_27335);
nor U28625 (N_28625,N_27235,N_26689);
nor U28626 (N_28626,N_26684,N_27763);
or U28627 (N_28627,N_26203,N_26033);
nand U28628 (N_28628,N_26049,N_26264);
nor U28629 (N_28629,N_27659,N_26387);
nor U28630 (N_28630,N_26027,N_26150);
nor U28631 (N_28631,N_27608,N_26748);
nand U28632 (N_28632,N_26028,N_26877);
and U28633 (N_28633,N_26594,N_26456);
xor U28634 (N_28634,N_27224,N_27536);
or U28635 (N_28635,N_27559,N_26544);
nand U28636 (N_28636,N_26273,N_26138);
and U28637 (N_28637,N_26235,N_26294);
and U28638 (N_28638,N_26924,N_26314);
xnor U28639 (N_28639,N_26992,N_27614);
nor U28640 (N_28640,N_27874,N_27695);
xnor U28641 (N_28641,N_27022,N_26532);
nor U28642 (N_28642,N_27909,N_26383);
nand U28643 (N_28643,N_26199,N_26609);
nor U28644 (N_28644,N_27767,N_26713);
nor U28645 (N_28645,N_26653,N_26135);
and U28646 (N_28646,N_27174,N_26521);
xor U28647 (N_28647,N_27950,N_27625);
nor U28648 (N_28648,N_27808,N_26746);
xnor U28649 (N_28649,N_26081,N_26342);
xor U28650 (N_28650,N_26876,N_27884);
xnor U28651 (N_28651,N_26216,N_27968);
or U28652 (N_28652,N_27686,N_27879);
and U28653 (N_28653,N_26667,N_27354);
nand U28654 (N_28654,N_26450,N_26611);
nor U28655 (N_28655,N_27697,N_27288);
nor U28656 (N_28656,N_26149,N_26276);
or U28657 (N_28657,N_27104,N_26493);
nand U28658 (N_28658,N_27298,N_27995);
or U28659 (N_28659,N_27386,N_26401);
or U28660 (N_28660,N_26284,N_27186);
and U28661 (N_28661,N_27936,N_26829);
and U28662 (N_28662,N_27331,N_27293);
xor U28663 (N_28663,N_26077,N_27391);
nand U28664 (N_28664,N_26117,N_26280);
nand U28665 (N_28665,N_27979,N_27748);
and U28666 (N_28666,N_26912,N_26736);
or U28667 (N_28667,N_26378,N_27751);
nor U28668 (N_28668,N_26613,N_27436);
or U28669 (N_28669,N_27992,N_27949);
or U28670 (N_28670,N_26850,N_26329);
xor U28671 (N_28671,N_26558,N_27712);
nor U28672 (N_28672,N_27316,N_26168);
nand U28673 (N_28673,N_27305,N_26491);
xnor U28674 (N_28674,N_26475,N_27394);
and U28675 (N_28675,N_27042,N_27277);
nand U28676 (N_28676,N_27080,N_27804);
xnor U28677 (N_28677,N_26134,N_27687);
and U28678 (N_28678,N_27229,N_27304);
nor U28679 (N_28679,N_26606,N_27644);
nor U28680 (N_28680,N_27511,N_26325);
or U28681 (N_28681,N_27611,N_27990);
xor U28682 (N_28682,N_26292,N_26079);
and U28683 (N_28683,N_27689,N_27591);
nor U28684 (N_28684,N_27225,N_27577);
nor U28685 (N_28685,N_26064,N_27289);
xor U28686 (N_28686,N_27905,N_26845);
xor U28687 (N_28687,N_27124,N_26628);
nand U28688 (N_28688,N_27303,N_27965);
and U28689 (N_28689,N_26650,N_27195);
nand U28690 (N_28690,N_27986,N_27622);
xor U28691 (N_28691,N_26278,N_27693);
nor U28692 (N_28692,N_26196,N_27508);
and U28693 (N_28693,N_26584,N_27890);
nand U28694 (N_28694,N_27520,N_27587);
nand U28695 (N_28695,N_27719,N_26722);
xnor U28696 (N_28696,N_26017,N_26842);
nand U28697 (N_28697,N_27012,N_26726);
or U28698 (N_28698,N_27059,N_26201);
xor U28699 (N_28699,N_26496,N_27877);
xor U28700 (N_28700,N_26019,N_27835);
nor U28701 (N_28701,N_26409,N_27203);
and U28702 (N_28702,N_27578,N_26696);
nor U28703 (N_28703,N_26721,N_26657);
nor U28704 (N_28704,N_27709,N_26448);
nor U28705 (N_28705,N_26119,N_27398);
or U28706 (N_28706,N_27119,N_27220);
nor U28707 (N_28707,N_26222,N_27839);
and U28708 (N_28708,N_26050,N_27074);
xnor U28709 (N_28709,N_27194,N_26384);
nor U28710 (N_28710,N_27144,N_26830);
nand U28711 (N_28711,N_27296,N_27690);
nand U28712 (N_28712,N_26483,N_26565);
nand U28713 (N_28713,N_27570,N_27895);
xor U28714 (N_28714,N_27954,N_26327);
nand U28715 (N_28715,N_27795,N_26075);
xnor U28716 (N_28716,N_27807,N_26952);
nor U28717 (N_28717,N_26697,N_26399);
xor U28718 (N_28718,N_27350,N_26806);
or U28719 (N_28719,N_26324,N_27170);
nand U28720 (N_28720,N_27704,N_27300);
or U28721 (N_28721,N_27247,N_26403);
nand U28722 (N_28722,N_27706,N_26930);
or U28723 (N_28723,N_26445,N_26385);
and U28724 (N_28724,N_27887,N_26919);
nor U28725 (N_28725,N_26178,N_27160);
nand U28726 (N_28726,N_26381,N_26617);
or U28727 (N_28727,N_27455,N_27645);
nand U28728 (N_28728,N_27779,N_26555);
or U28729 (N_28729,N_26754,N_27806);
nor U28730 (N_28730,N_27817,N_26607);
or U28731 (N_28731,N_27030,N_26418);
xor U28732 (N_28732,N_27353,N_27732);
nor U28733 (N_28733,N_26728,N_27112);
or U28734 (N_28734,N_27223,N_26258);
xnor U28735 (N_28735,N_26796,N_26176);
xnor U28736 (N_28736,N_27108,N_26922);
nor U28737 (N_28737,N_26818,N_26087);
or U28738 (N_28738,N_26641,N_26647);
and U28739 (N_28739,N_27991,N_26177);
nand U28740 (N_28740,N_26923,N_27786);
and U28741 (N_28741,N_27205,N_26983);
xor U28742 (N_28742,N_26582,N_26185);
or U28743 (N_28743,N_27981,N_27120);
or U28744 (N_28744,N_26805,N_27191);
and U28745 (N_28745,N_26900,N_27866);
xor U28746 (N_28746,N_27724,N_26529);
nand U28747 (N_28747,N_27820,N_27556);
and U28748 (N_28748,N_27978,N_27179);
xor U28749 (N_28749,N_27803,N_27312);
xor U28750 (N_28750,N_27502,N_26892);
or U28751 (N_28751,N_27328,N_27183);
nor U28752 (N_28752,N_26798,N_27474);
nand U28753 (N_28753,N_26572,N_27093);
or U28754 (N_28754,N_27237,N_27134);
xor U28755 (N_28755,N_26810,N_27009);
xnor U28756 (N_28756,N_27145,N_26066);
nand U28757 (N_28757,N_26788,N_26539);
nor U28758 (N_28758,N_26507,N_26742);
nand U28759 (N_28759,N_27266,N_27952);
and U28760 (N_28760,N_26014,N_27753);
xor U28761 (N_28761,N_27897,N_27998);
and U28762 (N_28762,N_27677,N_26593);
xnor U28763 (N_28763,N_27654,N_27368);
nand U28764 (N_28764,N_26504,N_26305);
nand U28765 (N_28765,N_26855,N_27206);
xor U28766 (N_28766,N_26827,N_27868);
or U28767 (N_28767,N_26088,N_26727);
and U28768 (N_28768,N_26408,N_27409);
nand U28769 (N_28769,N_27579,N_26652);
nor U28770 (N_28770,N_26449,N_26947);
or U28771 (N_28771,N_26026,N_26237);
nor U28772 (N_28772,N_26861,N_26241);
and U28773 (N_28773,N_26888,N_26295);
or U28774 (N_28774,N_27673,N_26394);
and U28775 (N_28775,N_26082,N_27064);
or U28776 (N_28776,N_26397,N_27257);
xor U28777 (N_28777,N_26574,N_26975);
xnor U28778 (N_28778,N_27427,N_26795);
and U28779 (N_28779,N_26690,N_27903);
xor U28780 (N_28780,N_27359,N_27721);
nand U28781 (N_28781,N_27886,N_27057);
nand U28782 (N_28782,N_26259,N_27458);
and U28783 (N_28783,N_26379,N_27052);
nand U28784 (N_28784,N_26671,N_26226);
nor U28785 (N_28785,N_26752,N_27845);
nor U28786 (N_28786,N_27613,N_27355);
xor U28787 (N_28787,N_27416,N_27571);
xor U28788 (N_28788,N_27097,N_27214);
nand U28789 (N_28789,N_26232,N_26503);
and U28790 (N_28790,N_27904,N_26246);
xnor U28791 (N_28791,N_27922,N_26506);
nor U28792 (N_28792,N_26053,N_26072);
xnor U28793 (N_28793,N_26266,N_26590);
and U28794 (N_28794,N_27023,N_26988);
nand U28795 (N_28795,N_27245,N_26141);
nor U28796 (N_28796,N_27572,N_27388);
xor U28797 (N_28797,N_26944,N_26787);
nand U28798 (N_28798,N_27385,N_27555);
xor U28799 (N_28799,N_27139,N_27601);
xor U28800 (N_28800,N_27742,N_27676);
and U28801 (N_28801,N_27821,N_27472);
or U28802 (N_28802,N_26981,N_26428);
or U28803 (N_28803,N_26147,N_26100);
and U28804 (N_28804,N_26619,N_26260);
xnor U28805 (N_28805,N_27011,N_27708);
or U28806 (N_28806,N_26200,N_26668);
or U28807 (N_28807,N_27481,N_26022);
xor U28808 (N_28808,N_26338,N_27452);
xnor U28809 (N_28809,N_26673,N_26895);
nor U28810 (N_28810,N_27953,N_27634);
or U28811 (N_28811,N_26808,N_26438);
xnor U28812 (N_28812,N_26476,N_27113);
xor U28813 (N_28813,N_27739,N_26340);
or U28814 (N_28814,N_27435,N_27210);
xor U28815 (N_28815,N_26644,N_27836);
nor U28816 (N_28816,N_27980,N_27580);
and U28817 (N_28817,N_27364,N_26965);
or U28818 (N_28818,N_27379,N_26686);
nand U28819 (N_28819,N_27766,N_26248);
and U28820 (N_28820,N_26648,N_26840);
xnor U28821 (N_28821,N_27172,N_26896);
or U28822 (N_28822,N_26866,N_26103);
nand U28823 (N_28823,N_26759,N_27215);
nand U28824 (N_28824,N_26535,N_27411);
or U28825 (N_28825,N_26769,N_27252);
xor U28826 (N_28826,N_26625,N_27518);
nand U28827 (N_28827,N_26763,N_26953);
or U28828 (N_28828,N_27605,N_27212);
nor U28829 (N_28829,N_26179,N_26616);
nor U28830 (N_28830,N_26782,N_26466);
xor U28831 (N_28831,N_26194,N_27276);
nor U28832 (N_28832,N_27263,N_27573);
or U28833 (N_28833,N_26270,N_26501);
or U28834 (N_28834,N_26227,N_27459);
nor U28835 (N_28835,N_26309,N_26863);
nor U28836 (N_28836,N_27913,N_27656);
nand U28837 (N_28837,N_27008,N_26301);
or U28838 (N_28838,N_27932,N_27216);
and U28839 (N_28839,N_26078,N_27412);
or U28840 (N_28840,N_26573,N_27648);
nand U28841 (N_28841,N_27610,N_27621);
xor U28842 (N_28842,N_27114,N_26160);
nand U28843 (N_28843,N_26189,N_26630);
xnor U28844 (N_28844,N_27207,N_27639);
and U28845 (N_28845,N_27027,N_26250);
and U28846 (N_28846,N_26832,N_27883);
xor U28847 (N_28847,N_27381,N_26335);
nand U28848 (N_28848,N_27149,N_27715);
xnor U28849 (N_28849,N_27576,N_27327);
and U28850 (N_28850,N_26681,N_27193);
nor U28851 (N_28851,N_27691,N_27734);
xor U28852 (N_28852,N_27658,N_26357);
xor U28853 (N_28853,N_27552,N_26847);
nor U28854 (N_28854,N_26654,N_27948);
and U28855 (N_28855,N_26737,N_27880);
and U28856 (N_28856,N_26093,N_27882);
and U28857 (N_28857,N_26240,N_27519);
xnor U28858 (N_28858,N_27906,N_27376);
and U28859 (N_28859,N_27213,N_27159);
xor U28860 (N_28860,N_26906,N_27467);
nor U28861 (N_28861,N_26320,N_26330);
xnor U28862 (N_28862,N_26954,N_26413);
and U28863 (N_28863,N_26511,N_27438);
nand U28864 (N_28864,N_27279,N_26623);
xor U28865 (N_28865,N_26592,N_26108);
and U28866 (N_28866,N_26643,N_27494);
nand U28867 (N_28867,N_26862,N_27524);
nand U28868 (N_28868,N_27138,N_26939);
or U28869 (N_28869,N_27222,N_27389);
nand U28870 (N_28870,N_27725,N_27087);
or U28871 (N_28871,N_27484,N_27792);
nand U28872 (N_28872,N_26732,N_27314);
nand U28873 (N_28873,N_26169,N_27847);
nor U28874 (N_28874,N_26800,N_27321);
nor U28875 (N_28875,N_26518,N_27361);
nor U28876 (N_28876,N_27357,N_26514);
xor U28877 (N_28877,N_27253,N_26719);
and U28878 (N_28878,N_27705,N_27674);
and U28879 (N_28879,N_26074,N_26211);
nor U28880 (N_28880,N_27827,N_27696);
or U28881 (N_28881,N_26228,N_27657);
or U28882 (N_28882,N_26753,N_26380);
xnor U28883 (N_28883,N_26298,N_27849);
and U28884 (N_28884,N_26372,N_27745);
xor U28885 (N_28885,N_27643,N_26367);
and U28886 (N_28886,N_26099,N_26645);
xnor U28887 (N_28887,N_26303,N_27553);
xnor U28888 (N_28888,N_27226,N_27862);
xor U28889 (N_28889,N_26206,N_27960);
or U28890 (N_28890,N_26512,N_26411);
and U28891 (N_28891,N_27337,N_26218);
nand U28892 (N_28892,N_26047,N_27900);
and U28893 (N_28893,N_26348,N_26094);
and U28894 (N_28894,N_26676,N_26034);
or U28895 (N_28895,N_26587,N_27204);
nor U28896 (N_28896,N_26202,N_26720);
nor U28897 (N_28897,N_26446,N_27428);
nand U28898 (N_28898,N_26410,N_27270);
nor U28899 (N_28899,N_27230,N_26688);
and U28900 (N_28900,N_26718,N_27307);
xor U28901 (N_28901,N_26204,N_27858);
nor U28902 (N_28902,N_27460,N_27758);
nand U28903 (N_28903,N_27189,N_26427);
or U28904 (N_28904,N_27616,N_26151);
nor U28905 (N_28905,N_26406,N_26274);
or U28906 (N_28906,N_27111,N_26943);
or U28907 (N_28907,N_26062,N_27258);
nand U28908 (N_28908,N_26997,N_27449);
nand U28909 (N_28909,N_27776,N_27015);
or U28910 (N_28910,N_27744,N_27778);
nor U28911 (N_28911,N_26111,N_27084);
or U28912 (N_28912,N_27607,N_26114);
nand U28913 (N_28913,N_26819,N_26471);
nand U28914 (N_28914,N_27034,N_26015);
nand U28915 (N_28915,N_26391,N_26239);
xnor U28916 (N_28916,N_26488,N_26649);
or U28917 (N_28917,N_27750,N_27001);
nor U28918 (N_28918,N_27439,N_27491);
nand U28919 (N_28919,N_27912,N_26774);
and U28920 (N_28920,N_27637,N_26656);
or U28921 (N_28921,N_26353,N_26887);
and U28922 (N_28922,N_26918,N_26741);
nand U28923 (N_28923,N_27540,N_27356);
or U28924 (N_28924,N_26580,N_26777);
nand U28925 (N_28925,N_27781,N_26140);
or U28926 (N_28926,N_27003,N_27941);
nor U28927 (N_28927,N_26578,N_26193);
or U28928 (N_28928,N_27780,N_26784);
nand U28929 (N_28929,N_26627,N_27014);
nor U28930 (N_28930,N_27295,N_26435);
nor U28931 (N_28931,N_27557,N_26351);
nor U28932 (N_28932,N_26040,N_27281);
nor U28933 (N_28933,N_26210,N_27958);
nand U28934 (N_28934,N_27450,N_27531);
nor U28935 (N_28935,N_27575,N_26595);
or U28936 (N_28936,N_26579,N_26101);
and U28937 (N_28937,N_26067,N_26437);
nand U28938 (N_28938,N_26929,N_26907);
and U28939 (N_28939,N_27341,N_26675);
and U28940 (N_28940,N_26281,N_26813);
nor U28941 (N_28941,N_26089,N_26756);
nand U28942 (N_28942,N_26288,N_26358);
nand U28943 (N_28943,N_26398,N_26879);
nor U28944 (N_28944,N_26083,N_27896);
nor U28945 (N_28945,N_27533,N_27197);
and U28946 (N_28946,N_26037,N_26130);
xor U28947 (N_28947,N_27164,N_27055);
or U28948 (N_28948,N_26307,N_26495);
and U28949 (N_28949,N_27726,N_27187);
nand U28950 (N_28950,N_27371,N_26872);
nand U28951 (N_28951,N_26683,N_27509);
xnor U28952 (N_28952,N_26664,N_27670);
and U28953 (N_28953,N_27503,N_27322);
and U28954 (N_28954,N_27917,N_27248);
and U28955 (N_28955,N_27169,N_26963);
nor U28956 (N_28956,N_26821,N_27400);
or U28957 (N_28957,N_26148,N_27800);
nand U28958 (N_28958,N_27728,N_26598);
nand U28959 (N_28959,N_26905,N_27541);
or U28960 (N_28960,N_27554,N_27852);
and U28961 (N_28961,N_26124,N_26008);
xor U28962 (N_28962,N_26389,N_27329);
nor U28963 (N_28963,N_26416,N_27283);
nor U28964 (N_28964,N_27813,N_27662);
and U28965 (N_28965,N_26797,N_26245);
and U28966 (N_28966,N_27632,N_26010);
xnor U28967 (N_28967,N_26577,N_26405);
or U28968 (N_28968,N_26058,N_26156);
nor U28969 (N_28969,N_27672,N_27826);
nand U28970 (N_28970,N_27402,N_27152);
and U28971 (N_28971,N_26031,N_26971);
or U28972 (N_28972,N_27418,N_27926);
or U28973 (N_28973,N_26091,N_27142);
or U28974 (N_28974,N_26600,N_27513);
xor U28975 (N_28975,N_26326,N_26817);
or U28976 (N_28976,N_27417,N_26802);
and U28977 (N_28977,N_27431,N_26825);
nand U28978 (N_28978,N_26068,N_27851);
xnor U28979 (N_28979,N_26170,N_27604);
and U28980 (N_28980,N_27284,N_26374);
and U28981 (N_28981,N_27782,N_27343);
and U28982 (N_28982,N_26663,N_27345);
or U28983 (N_28983,N_27878,N_26480);
and U28984 (N_28984,N_27599,N_26785);
and U28985 (N_28985,N_26588,N_27373);
xnor U28986 (N_28986,N_26723,N_26581);
nor U28987 (N_28987,N_27118,N_27669);
or U28988 (N_28988,N_26112,N_26106);
and U28989 (N_28989,N_26634,N_27241);
and U28990 (N_28990,N_27970,N_27951);
or U28991 (N_28991,N_26126,N_26317);
and U28992 (N_28992,N_27261,N_27384);
xnor U28993 (N_28993,N_26490,N_27685);
and U28994 (N_28994,N_26814,N_27088);
and U28995 (N_28995,N_27711,N_26287);
nor U28996 (N_28996,N_27399,N_26974);
nand U28997 (N_28997,N_27078,N_26526);
xor U28998 (N_28998,N_27799,N_27888);
nor U28999 (N_28999,N_26725,N_27349);
or U29000 (N_29000,N_26045,N_26406);
xor U29001 (N_29001,N_26942,N_27537);
nand U29002 (N_29002,N_27728,N_26442);
xnor U29003 (N_29003,N_27633,N_27514);
or U29004 (N_29004,N_26968,N_27231);
and U29005 (N_29005,N_27747,N_26383);
or U29006 (N_29006,N_27165,N_26465);
xor U29007 (N_29007,N_26864,N_26210);
nand U29008 (N_29008,N_27207,N_26257);
or U29009 (N_29009,N_27979,N_26933);
and U29010 (N_29010,N_26470,N_26169);
nand U29011 (N_29011,N_27136,N_26623);
and U29012 (N_29012,N_27682,N_26200);
nor U29013 (N_29013,N_27411,N_27140);
and U29014 (N_29014,N_27613,N_27460);
or U29015 (N_29015,N_27066,N_27144);
nor U29016 (N_29016,N_27493,N_26998);
xor U29017 (N_29017,N_27259,N_27486);
nand U29018 (N_29018,N_27951,N_26242);
xnor U29019 (N_29019,N_27368,N_27138);
nor U29020 (N_29020,N_26823,N_26021);
nor U29021 (N_29021,N_27750,N_26775);
xnor U29022 (N_29022,N_26392,N_27588);
and U29023 (N_29023,N_27052,N_27371);
nor U29024 (N_29024,N_27441,N_26185);
nand U29025 (N_29025,N_26012,N_27949);
or U29026 (N_29026,N_26467,N_26660);
xnor U29027 (N_29027,N_27375,N_27329);
and U29028 (N_29028,N_26062,N_27666);
xor U29029 (N_29029,N_27932,N_27354);
or U29030 (N_29030,N_27294,N_26090);
or U29031 (N_29031,N_26404,N_27254);
and U29032 (N_29032,N_26776,N_27579);
nand U29033 (N_29033,N_26106,N_26542);
and U29034 (N_29034,N_26814,N_27865);
or U29035 (N_29035,N_27729,N_26006);
or U29036 (N_29036,N_27217,N_27549);
or U29037 (N_29037,N_26534,N_27678);
nor U29038 (N_29038,N_27777,N_26110);
xor U29039 (N_29039,N_27004,N_26763);
nor U29040 (N_29040,N_27091,N_27727);
nor U29041 (N_29041,N_27270,N_27752);
xnor U29042 (N_29042,N_26065,N_26159);
and U29043 (N_29043,N_27190,N_27778);
xnor U29044 (N_29044,N_27284,N_27665);
and U29045 (N_29045,N_26970,N_26193);
nand U29046 (N_29046,N_26468,N_26382);
nor U29047 (N_29047,N_27967,N_26531);
nor U29048 (N_29048,N_26449,N_26471);
nand U29049 (N_29049,N_26017,N_26629);
xnor U29050 (N_29050,N_27513,N_27415);
xnor U29051 (N_29051,N_27334,N_26088);
and U29052 (N_29052,N_27985,N_26955);
xor U29053 (N_29053,N_26414,N_26302);
and U29054 (N_29054,N_27802,N_26470);
and U29055 (N_29055,N_26647,N_26687);
nor U29056 (N_29056,N_26394,N_26359);
nor U29057 (N_29057,N_27758,N_26959);
xor U29058 (N_29058,N_26059,N_27776);
xnor U29059 (N_29059,N_27644,N_26992);
nand U29060 (N_29060,N_27596,N_27867);
nand U29061 (N_29061,N_27994,N_27946);
xor U29062 (N_29062,N_27589,N_26137);
nor U29063 (N_29063,N_27953,N_26194);
xor U29064 (N_29064,N_27609,N_26018);
and U29065 (N_29065,N_26884,N_27843);
xor U29066 (N_29066,N_26888,N_26881);
or U29067 (N_29067,N_26099,N_27684);
or U29068 (N_29068,N_27982,N_26127);
xor U29069 (N_29069,N_26906,N_27395);
or U29070 (N_29070,N_27785,N_27467);
nor U29071 (N_29071,N_27284,N_26288);
or U29072 (N_29072,N_27035,N_27282);
xor U29073 (N_29073,N_26450,N_26251);
and U29074 (N_29074,N_27025,N_27430);
xnor U29075 (N_29075,N_27964,N_27752);
and U29076 (N_29076,N_27790,N_27674);
and U29077 (N_29077,N_27540,N_27870);
nor U29078 (N_29078,N_26250,N_26683);
nand U29079 (N_29079,N_26722,N_26407);
and U29080 (N_29080,N_26265,N_27328);
and U29081 (N_29081,N_26818,N_27665);
xor U29082 (N_29082,N_27368,N_26133);
nand U29083 (N_29083,N_27750,N_26068);
nand U29084 (N_29084,N_27191,N_27566);
and U29085 (N_29085,N_27126,N_26498);
or U29086 (N_29086,N_27297,N_27907);
nor U29087 (N_29087,N_27627,N_27156);
nor U29088 (N_29088,N_26167,N_26339);
nand U29089 (N_29089,N_27421,N_26457);
nand U29090 (N_29090,N_27888,N_27793);
or U29091 (N_29091,N_26553,N_26923);
nand U29092 (N_29092,N_26311,N_26866);
and U29093 (N_29093,N_27839,N_26121);
nor U29094 (N_29094,N_27002,N_27166);
xor U29095 (N_29095,N_27114,N_27074);
and U29096 (N_29096,N_26893,N_27251);
nor U29097 (N_29097,N_26919,N_27305);
xor U29098 (N_29098,N_27364,N_26897);
xor U29099 (N_29099,N_26329,N_27462);
nor U29100 (N_29100,N_27493,N_26016);
or U29101 (N_29101,N_27886,N_26844);
xnor U29102 (N_29102,N_26211,N_26448);
and U29103 (N_29103,N_26284,N_26182);
nand U29104 (N_29104,N_27971,N_26940);
and U29105 (N_29105,N_26199,N_26864);
nand U29106 (N_29106,N_26025,N_27056);
xor U29107 (N_29107,N_26680,N_26712);
nor U29108 (N_29108,N_26617,N_26245);
nand U29109 (N_29109,N_27512,N_27005);
or U29110 (N_29110,N_26923,N_27152);
nor U29111 (N_29111,N_26844,N_26508);
nor U29112 (N_29112,N_27000,N_27589);
nor U29113 (N_29113,N_27227,N_27285);
xnor U29114 (N_29114,N_27064,N_27442);
or U29115 (N_29115,N_26291,N_26143);
nand U29116 (N_29116,N_26643,N_26775);
or U29117 (N_29117,N_26987,N_26809);
xnor U29118 (N_29118,N_27003,N_26423);
nand U29119 (N_29119,N_27251,N_26868);
nor U29120 (N_29120,N_26423,N_26633);
or U29121 (N_29121,N_27381,N_27095);
nand U29122 (N_29122,N_26544,N_27751);
and U29123 (N_29123,N_26628,N_26639);
nor U29124 (N_29124,N_26955,N_27238);
xnor U29125 (N_29125,N_26355,N_27793);
or U29126 (N_29126,N_27302,N_26775);
nand U29127 (N_29127,N_26044,N_26249);
nor U29128 (N_29128,N_27820,N_27940);
and U29129 (N_29129,N_27280,N_26091);
nor U29130 (N_29130,N_27503,N_27377);
and U29131 (N_29131,N_27379,N_26873);
and U29132 (N_29132,N_26235,N_27335);
or U29133 (N_29133,N_26254,N_26145);
xor U29134 (N_29134,N_26315,N_26389);
and U29135 (N_29135,N_27110,N_26367);
nand U29136 (N_29136,N_27686,N_26064);
or U29137 (N_29137,N_26644,N_27003);
nand U29138 (N_29138,N_26522,N_26321);
xor U29139 (N_29139,N_26080,N_27311);
xor U29140 (N_29140,N_27655,N_26869);
xnor U29141 (N_29141,N_27088,N_26108);
or U29142 (N_29142,N_27743,N_26914);
nor U29143 (N_29143,N_26358,N_26553);
and U29144 (N_29144,N_27363,N_27624);
nor U29145 (N_29145,N_27601,N_27356);
and U29146 (N_29146,N_26217,N_27443);
xnor U29147 (N_29147,N_26461,N_27757);
nand U29148 (N_29148,N_27503,N_26293);
or U29149 (N_29149,N_26295,N_27497);
nor U29150 (N_29150,N_27188,N_27095);
nand U29151 (N_29151,N_26414,N_27330);
nand U29152 (N_29152,N_27630,N_27312);
nand U29153 (N_29153,N_27067,N_26183);
nand U29154 (N_29154,N_26766,N_26031);
nand U29155 (N_29155,N_26030,N_27131);
or U29156 (N_29156,N_26359,N_27769);
xnor U29157 (N_29157,N_27392,N_26091);
and U29158 (N_29158,N_27965,N_27630);
nor U29159 (N_29159,N_26904,N_27939);
and U29160 (N_29160,N_26083,N_26157);
or U29161 (N_29161,N_26230,N_26059);
nand U29162 (N_29162,N_27440,N_26117);
and U29163 (N_29163,N_27105,N_27311);
nand U29164 (N_29164,N_27679,N_26660);
nand U29165 (N_29165,N_26645,N_27404);
xor U29166 (N_29166,N_26883,N_26835);
or U29167 (N_29167,N_27242,N_27198);
nor U29168 (N_29168,N_27401,N_27841);
and U29169 (N_29169,N_27966,N_26182);
nor U29170 (N_29170,N_27609,N_27052);
nor U29171 (N_29171,N_27235,N_26756);
nand U29172 (N_29172,N_26764,N_26015);
nand U29173 (N_29173,N_27554,N_27673);
nor U29174 (N_29174,N_27797,N_26373);
xor U29175 (N_29175,N_27052,N_27341);
nor U29176 (N_29176,N_27096,N_26353);
and U29177 (N_29177,N_26827,N_27005);
xnor U29178 (N_29178,N_26914,N_26586);
or U29179 (N_29179,N_27751,N_26497);
nor U29180 (N_29180,N_27732,N_26468);
or U29181 (N_29181,N_26562,N_26677);
or U29182 (N_29182,N_26587,N_26262);
xnor U29183 (N_29183,N_27266,N_27188);
and U29184 (N_29184,N_26461,N_26059);
nor U29185 (N_29185,N_26023,N_26565);
nand U29186 (N_29186,N_26950,N_26808);
nor U29187 (N_29187,N_27277,N_26707);
xor U29188 (N_29188,N_26312,N_27064);
and U29189 (N_29189,N_26639,N_27065);
and U29190 (N_29190,N_26225,N_27996);
nor U29191 (N_29191,N_27871,N_27691);
nand U29192 (N_29192,N_27172,N_27740);
or U29193 (N_29193,N_26007,N_27765);
xor U29194 (N_29194,N_26564,N_27196);
or U29195 (N_29195,N_26455,N_26319);
xor U29196 (N_29196,N_26606,N_26905);
nor U29197 (N_29197,N_27749,N_26426);
xnor U29198 (N_29198,N_26181,N_27374);
or U29199 (N_29199,N_27766,N_26484);
and U29200 (N_29200,N_27667,N_27077);
xor U29201 (N_29201,N_26607,N_27835);
nand U29202 (N_29202,N_26945,N_26526);
or U29203 (N_29203,N_27557,N_26527);
or U29204 (N_29204,N_26603,N_26048);
xnor U29205 (N_29205,N_26306,N_26031);
nand U29206 (N_29206,N_27044,N_27984);
nand U29207 (N_29207,N_27067,N_26264);
and U29208 (N_29208,N_27675,N_27912);
and U29209 (N_29209,N_26520,N_26539);
xnor U29210 (N_29210,N_26742,N_26896);
xor U29211 (N_29211,N_27032,N_27738);
nor U29212 (N_29212,N_26764,N_26111);
nor U29213 (N_29213,N_27987,N_26773);
nor U29214 (N_29214,N_26032,N_27135);
or U29215 (N_29215,N_27175,N_26649);
nor U29216 (N_29216,N_26955,N_26907);
nor U29217 (N_29217,N_27818,N_26919);
nor U29218 (N_29218,N_27832,N_27035);
and U29219 (N_29219,N_27469,N_27508);
and U29220 (N_29220,N_26590,N_26164);
or U29221 (N_29221,N_27155,N_27108);
and U29222 (N_29222,N_26842,N_27176);
or U29223 (N_29223,N_27091,N_26746);
or U29224 (N_29224,N_26268,N_26596);
xnor U29225 (N_29225,N_26728,N_27266);
or U29226 (N_29226,N_27111,N_26436);
and U29227 (N_29227,N_26406,N_27477);
nor U29228 (N_29228,N_27921,N_27355);
and U29229 (N_29229,N_27501,N_27406);
xnor U29230 (N_29230,N_26903,N_27280);
or U29231 (N_29231,N_26459,N_26300);
nor U29232 (N_29232,N_27567,N_26859);
and U29233 (N_29233,N_27394,N_26142);
xnor U29234 (N_29234,N_26557,N_26216);
xnor U29235 (N_29235,N_26664,N_26869);
and U29236 (N_29236,N_26105,N_27690);
or U29237 (N_29237,N_26614,N_27313);
or U29238 (N_29238,N_26066,N_26644);
or U29239 (N_29239,N_26225,N_27619);
nand U29240 (N_29240,N_26915,N_26545);
nand U29241 (N_29241,N_26391,N_26050);
or U29242 (N_29242,N_27855,N_26906);
xor U29243 (N_29243,N_26173,N_27390);
xnor U29244 (N_29244,N_26281,N_26873);
xor U29245 (N_29245,N_26673,N_26536);
xor U29246 (N_29246,N_26943,N_27186);
and U29247 (N_29247,N_26884,N_26617);
xnor U29248 (N_29248,N_26263,N_27715);
and U29249 (N_29249,N_26236,N_26680);
or U29250 (N_29250,N_27581,N_26892);
or U29251 (N_29251,N_26271,N_27523);
or U29252 (N_29252,N_27235,N_27634);
nor U29253 (N_29253,N_26239,N_26757);
nor U29254 (N_29254,N_27618,N_26654);
or U29255 (N_29255,N_27328,N_26740);
and U29256 (N_29256,N_26136,N_27238);
xor U29257 (N_29257,N_26226,N_26489);
xor U29258 (N_29258,N_26119,N_26166);
xnor U29259 (N_29259,N_27897,N_26207);
xnor U29260 (N_29260,N_27563,N_27911);
or U29261 (N_29261,N_27361,N_26394);
or U29262 (N_29262,N_26425,N_27901);
or U29263 (N_29263,N_27645,N_26489);
or U29264 (N_29264,N_26813,N_26788);
and U29265 (N_29265,N_26026,N_26263);
nor U29266 (N_29266,N_27953,N_26617);
nand U29267 (N_29267,N_27986,N_27743);
nor U29268 (N_29268,N_26090,N_26584);
nand U29269 (N_29269,N_26767,N_27149);
xor U29270 (N_29270,N_26686,N_26929);
nor U29271 (N_29271,N_26428,N_26733);
xnor U29272 (N_29272,N_27309,N_27357);
and U29273 (N_29273,N_27513,N_27442);
nor U29274 (N_29274,N_27529,N_26003);
nand U29275 (N_29275,N_26500,N_26730);
and U29276 (N_29276,N_26394,N_26991);
and U29277 (N_29277,N_26916,N_26221);
and U29278 (N_29278,N_27903,N_26851);
nor U29279 (N_29279,N_27843,N_26955);
nor U29280 (N_29280,N_27137,N_27792);
and U29281 (N_29281,N_26236,N_27800);
nor U29282 (N_29282,N_26000,N_27640);
and U29283 (N_29283,N_26792,N_27766);
xor U29284 (N_29284,N_26877,N_27558);
nand U29285 (N_29285,N_27101,N_26587);
nor U29286 (N_29286,N_27468,N_26533);
nand U29287 (N_29287,N_26697,N_27480);
xor U29288 (N_29288,N_26581,N_26343);
xnor U29289 (N_29289,N_26290,N_27697);
nor U29290 (N_29290,N_27046,N_26813);
nand U29291 (N_29291,N_26839,N_26458);
nor U29292 (N_29292,N_27306,N_26329);
and U29293 (N_29293,N_27765,N_27790);
and U29294 (N_29294,N_26308,N_26400);
and U29295 (N_29295,N_27720,N_27610);
and U29296 (N_29296,N_26495,N_26270);
nand U29297 (N_29297,N_26989,N_27670);
or U29298 (N_29298,N_26947,N_26858);
nor U29299 (N_29299,N_26446,N_27310);
or U29300 (N_29300,N_27494,N_27542);
nor U29301 (N_29301,N_26407,N_27744);
nor U29302 (N_29302,N_26030,N_27808);
xnor U29303 (N_29303,N_27127,N_26815);
and U29304 (N_29304,N_26070,N_26341);
nand U29305 (N_29305,N_26808,N_27340);
nor U29306 (N_29306,N_26842,N_27743);
nor U29307 (N_29307,N_27769,N_26547);
nand U29308 (N_29308,N_27557,N_27165);
xnor U29309 (N_29309,N_26695,N_26952);
nand U29310 (N_29310,N_26694,N_26730);
nand U29311 (N_29311,N_26115,N_26088);
xnor U29312 (N_29312,N_26077,N_26295);
or U29313 (N_29313,N_26781,N_26667);
nor U29314 (N_29314,N_27751,N_26969);
and U29315 (N_29315,N_26921,N_27212);
nand U29316 (N_29316,N_27150,N_26972);
nor U29317 (N_29317,N_26974,N_26999);
nor U29318 (N_29318,N_27042,N_27881);
nand U29319 (N_29319,N_26168,N_27302);
or U29320 (N_29320,N_26782,N_27693);
and U29321 (N_29321,N_27766,N_26818);
nor U29322 (N_29322,N_26207,N_27332);
nor U29323 (N_29323,N_26178,N_27145);
and U29324 (N_29324,N_27246,N_26809);
and U29325 (N_29325,N_26435,N_27205);
or U29326 (N_29326,N_26455,N_26510);
nor U29327 (N_29327,N_27393,N_27894);
or U29328 (N_29328,N_26853,N_27587);
or U29329 (N_29329,N_26138,N_27270);
nand U29330 (N_29330,N_26918,N_27530);
nor U29331 (N_29331,N_26512,N_27294);
and U29332 (N_29332,N_27184,N_26752);
nand U29333 (N_29333,N_26667,N_26763);
xor U29334 (N_29334,N_26584,N_27085);
nor U29335 (N_29335,N_27246,N_27586);
nor U29336 (N_29336,N_27318,N_26100);
nand U29337 (N_29337,N_26310,N_27870);
and U29338 (N_29338,N_26050,N_27779);
or U29339 (N_29339,N_26121,N_26595);
and U29340 (N_29340,N_27784,N_27783);
or U29341 (N_29341,N_26618,N_27327);
nand U29342 (N_29342,N_26184,N_27002);
xnor U29343 (N_29343,N_26665,N_27753);
and U29344 (N_29344,N_26915,N_26760);
nor U29345 (N_29345,N_27853,N_27587);
or U29346 (N_29346,N_27383,N_27522);
or U29347 (N_29347,N_27064,N_26544);
nand U29348 (N_29348,N_27685,N_27548);
xor U29349 (N_29349,N_27623,N_27248);
or U29350 (N_29350,N_26950,N_26554);
xnor U29351 (N_29351,N_27798,N_27650);
or U29352 (N_29352,N_27955,N_27886);
xor U29353 (N_29353,N_26276,N_26900);
nor U29354 (N_29354,N_27019,N_26411);
and U29355 (N_29355,N_26166,N_26533);
nand U29356 (N_29356,N_27824,N_27325);
nand U29357 (N_29357,N_26661,N_27378);
nor U29358 (N_29358,N_27584,N_26088);
nor U29359 (N_29359,N_27676,N_26818);
nor U29360 (N_29360,N_27048,N_27311);
nand U29361 (N_29361,N_27765,N_27961);
and U29362 (N_29362,N_27035,N_26315);
nand U29363 (N_29363,N_26392,N_27710);
xnor U29364 (N_29364,N_27542,N_26577);
or U29365 (N_29365,N_26889,N_26966);
nor U29366 (N_29366,N_26924,N_26648);
and U29367 (N_29367,N_26192,N_26257);
or U29368 (N_29368,N_27961,N_26056);
nand U29369 (N_29369,N_27580,N_26756);
and U29370 (N_29370,N_27098,N_26723);
nor U29371 (N_29371,N_27481,N_26683);
nand U29372 (N_29372,N_26347,N_27403);
nand U29373 (N_29373,N_27295,N_26233);
xnor U29374 (N_29374,N_27963,N_26125);
nor U29375 (N_29375,N_26819,N_26228);
and U29376 (N_29376,N_26995,N_27819);
and U29377 (N_29377,N_26381,N_27844);
or U29378 (N_29378,N_26846,N_26049);
nand U29379 (N_29379,N_27478,N_26307);
nor U29380 (N_29380,N_27951,N_26994);
nand U29381 (N_29381,N_27841,N_26890);
and U29382 (N_29382,N_27457,N_26187);
nor U29383 (N_29383,N_26365,N_26095);
or U29384 (N_29384,N_26952,N_27925);
xor U29385 (N_29385,N_26352,N_26244);
xnor U29386 (N_29386,N_26867,N_27065);
or U29387 (N_29387,N_26636,N_26584);
nor U29388 (N_29388,N_26262,N_27766);
xor U29389 (N_29389,N_27886,N_26741);
or U29390 (N_29390,N_27435,N_26427);
nand U29391 (N_29391,N_26065,N_26385);
and U29392 (N_29392,N_26930,N_26440);
or U29393 (N_29393,N_26672,N_27968);
xor U29394 (N_29394,N_27972,N_27612);
nor U29395 (N_29395,N_26253,N_26071);
xor U29396 (N_29396,N_26745,N_27644);
nor U29397 (N_29397,N_26760,N_27152);
xnor U29398 (N_29398,N_27408,N_27761);
or U29399 (N_29399,N_26205,N_26296);
nand U29400 (N_29400,N_26716,N_26157);
and U29401 (N_29401,N_26010,N_27004);
and U29402 (N_29402,N_26672,N_26996);
nor U29403 (N_29403,N_26637,N_26340);
xor U29404 (N_29404,N_26130,N_27929);
or U29405 (N_29405,N_27848,N_27338);
nor U29406 (N_29406,N_26708,N_27368);
nand U29407 (N_29407,N_26316,N_27140);
xnor U29408 (N_29408,N_27498,N_27919);
or U29409 (N_29409,N_26753,N_27428);
or U29410 (N_29410,N_27941,N_26241);
nand U29411 (N_29411,N_27370,N_26996);
nor U29412 (N_29412,N_27024,N_26176);
and U29413 (N_29413,N_26386,N_26721);
or U29414 (N_29414,N_27229,N_26734);
nor U29415 (N_29415,N_26863,N_27719);
and U29416 (N_29416,N_26943,N_27952);
xor U29417 (N_29417,N_27906,N_27157);
or U29418 (N_29418,N_27755,N_27308);
and U29419 (N_29419,N_26256,N_26399);
nor U29420 (N_29420,N_27441,N_27535);
nor U29421 (N_29421,N_27912,N_26797);
xor U29422 (N_29422,N_27553,N_26962);
xor U29423 (N_29423,N_26275,N_26485);
xor U29424 (N_29424,N_26085,N_26684);
nand U29425 (N_29425,N_26382,N_27866);
and U29426 (N_29426,N_27424,N_26673);
or U29427 (N_29427,N_27712,N_26826);
nand U29428 (N_29428,N_27679,N_26503);
nor U29429 (N_29429,N_27837,N_26758);
nor U29430 (N_29430,N_26238,N_27681);
nand U29431 (N_29431,N_26355,N_26899);
nor U29432 (N_29432,N_27224,N_27336);
and U29433 (N_29433,N_27913,N_27169);
or U29434 (N_29434,N_26589,N_27576);
or U29435 (N_29435,N_26217,N_27565);
or U29436 (N_29436,N_26906,N_26098);
nand U29437 (N_29437,N_26582,N_26773);
nand U29438 (N_29438,N_26234,N_26691);
or U29439 (N_29439,N_27270,N_27827);
nand U29440 (N_29440,N_27107,N_26977);
and U29441 (N_29441,N_27352,N_27708);
nor U29442 (N_29442,N_27502,N_27332);
xnor U29443 (N_29443,N_27926,N_26421);
nand U29444 (N_29444,N_26575,N_27246);
nand U29445 (N_29445,N_26641,N_27245);
xnor U29446 (N_29446,N_26097,N_27425);
nor U29447 (N_29447,N_26810,N_27061);
or U29448 (N_29448,N_27550,N_26756);
nand U29449 (N_29449,N_26797,N_26631);
xnor U29450 (N_29450,N_26399,N_26547);
nor U29451 (N_29451,N_26762,N_26098);
nor U29452 (N_29452,N_26310,N_26093);
xor U29453 (N_29453,N_26887,N_26825);
and U29454 (N_29454,N_27986,N_27860);
nand U29455 (N_29455,N_27012,N_27288);
or U29456 (N_29456,N_27840,N_26978);
xnor U29457 (N_29457,N_27700,N_26465);
nor U29458 (N_29458,N_27964,N_27274);
xnor U29459 (N_29459,N_26920,N_27139);
and U29460 (N_29460,N_26860,N_27901);
nand U29461 (N_29461,N_26785,N_26075);
xor U29462 (N_29462,N_26344,N_27357);
nand U29463 (N_29463,N_26697,N_26338);
nand U29464 (N_29464,N_26616,N_27517);
nand U29465 (N_29465,N_26470,N_26195);
and U29466 (N_29466,N_26147,N_26473);
nor U29467 (N_29467,N_27927,N_26198);
xor U29468 (N_29468,N_26935,N_26540);
nand U29469 (N_29469,N_26400,N_27931);
or U29470 (N_29470,N_27331,N_27498);
and U29471 (N_29471,N_26042,N_26426);
or U29472 (N_29472,N_26868,N_26893);
nand U29473 (N_29473,N_27820,N_26439);
or U29474 (N_29474,N_26212,N_26029);
nand U29475 (N_29475,N_27176,N_27966);
nor U29476 (N_29476,N_27389,N_26366);
and U29477 (N_29477,N_26925,N_27566);
nand U29478 (N_29478,N_26645,N_26199);
xor U29479 (N_29479,N_26025,N_27736);
or U29480 (N_29480,N_27101,N_27937);
nand U29481 (N_29481,N_26367,N_26674);
and U29482 (N_29482,N_26635,N_26082);
and U29483 (N_29483,N_27229,N_26770);
and U29484 (N_29484,N_26967,N_26016);
or U29485 (N_29485,N_26842,N_27045);
or U29486 (N_29486,N_27174,N_27669);
nand U29487 (N_29487,N_26610,N_27739);
and U29488 (N_29488,N_27612,N_26577);
and U29489 (N_29489,N_27149,N_26391);
nand U29490 (N_29490,N_27014,N_27880);
nand U29491 (N_29491,N_27458,N_27406);
or U29492 (N_29492,N_26440,N_26842);
nor U29493 (N_29493,N_27812,N_27321);
and U29494 (N_29494,N_26717,N_27547);
and U29495 (N_29495,N_26568,N_27139);
nor U29496 (N_29496,N_27756,N_27557);
nand U29497 (N_29497,N_27305,N_27134);
and U29498 (N_29498,N_26967,N_26053);
nand U29499 (N_29499,N_27906,N_26584);
nand U29500 (N_29500,N_27619,N_26197);
nand U29501 (N_29501,N_26154,N_26099);
xnor U29502 (N_29502,N_27567,N_27249);
and U29503 (N_29503,N_26869,N_27496);
or U29504 (N_29504,N_26617,N_26202);
or U29505 (N_29505,N_26095,N_26816);
nor U29506 (N_29506,N_27778,N_27555);
nor U29507 (N_29507,N_26605,N_27672);
xor U29508 (N_29508,N_27720,N_27413);
nand U29509 (N_29509,N_26720,N_26070);
or U29510 (N_29510,N_27761,N_27116);
and U29511 (N_29511,N_27034,N_26499);
nand U29512 (N_29512,N_27294,N_27020);
xnor U29513 (N_29513,N_26491,N_27843);
xnor U29514 (N_29514,N_27100,N_27165);
or U29515 (N_29515,N_26752,N_27558);
xor U29516 (N_29516,N_27784,N_26277);
nor U29517 (N_29517,N_27108,N_27901);
or U29518 (N_29518,N_26202,N_27843);
or U29519 (N_29519,N_27084,N_27451);
or U29520 (N_29520,N_27300,N_27983);
nor U29521 (N_29521,N_26436,N_26483);
xnor U29522 (N_29522,N_26389,N_26123);
and U29523 (N_29523,N_27929,N_26160);
and U29524 (N_29524,N_27676,N_27152);
xnor U29525 (N_29525,N_26886,N_27642);
or U29526 (N_29526,N_27282,N_27316);
or U29527 (N_29527,N_26056,N_27184);
xnor U29528 (N_29528,N_26023,N_27117);
and U29529 (N_29529,N_26043,N_27873);
nand U29530 (N_29530,N_26946,N_26392);
and U29531 (N_29531,N_27647,N_27513);
nor U29532 (N_29532,N_27253,N_26588);
nor U29533 (N_29533,N_27244,N_26066);
or U29534 (N_29534,N_26164,N_27098);
nand U29535 (N_29535,N_27008,N_26269);
nand U29536 (N_29536,N_26952,N_26521);
xnor U29537 (N_29537,N_27168,N_26648);
or U29538 (N_29538,N_27839,N_27587);
xor U29539 (N_29539,N_27729,N_27528);
and U29540 (N_29540,N_27265,N_26528);
xor U29541 (N_29541,N_26157,N_27877);
nand U29542 (N_29542,N_26983,N_26772);
nor U29543 (N_29543,N_27026,N_26731);
xor U29544 (N_29544,N_26086,N_26413);
or U29545 (N_29545,N_26967,N_27157);
or U29546 (N_29546,N_26798,N_27763);
or U29547 (N_29547,N_27899,N_27883);
xor U29548 (N_29548,N_27534,N_27752);
nor U29549 (N_29549,N_27307,N_26021);
and U29550 (N_29550,N_26613,N_26137);
nor U29551 (N_29551,N_26789,N_27147);
nand U29552 (N_29552,N_26085,N_27768);
nand U29553 (N_29553,N_27284,N_27560);
and U29554 (N_29554,N_26368,N_27078);
and U29555 (N_29555,N_27120,N_26969);
nor U29556 (N_29556,N_26575,N_27914);
xor U29557 (N_29557,N_26825,N_27361);
or U29558 (N_29558,N_26760,N_26785);
nand U29559 (N_29559,N_26846,N_27266);
nand U29560 (N_29560,N_26857,N_26740);
or U29561 (N_29561,N_27279,N_27504);
and U29562 (N_29562,N_26736,N_27456);
nor U29563 (N_29563,N_26542,N_26652);
nand U29564 (N_29564,N_27438,N_26428);
or U29565 (N_29565,N_26343,N_26901);
and U29566 (N_29566,N_27773,N_27654);
nand U29567 (N_29567,N_26164,N_27878);
or U29568 (N_29568,N_26531,N_27374);
xor U29569 (N_29569,N_27986,N_27584);
nor U29570 (N_29570,N_26747,N_26991);
and U29571 (N_29571,N_26526,N_26379);
and U29572 (N_29572,N_26676,N_27152);
nand U29573 (N_29573,N_26980,N_27698);
nand U29574 (N_29574,N_27295,N_27047);
or U29575 (N_29575,N_27165,N_27106);
and U29576 (N_29576,N_27522,N_27822);
nand U29577 (N_29577,N_27793,N_26723);
or U29578 (N_29578,N_26790,N_27490);
xnor U29579 (N_29579,N_27712,N_27704);
nor U29580 (N_29580,N_27328,N_26163);
nand U29581 (N_29581,N_27152,N_26203);
nor U29582 (N_29582,N_26050,N_27467);
or U29583 (N_29583,N_27631,N_27507);
xnor U29584 (N_29584,N_27904,N_26614);
nand U29585 (N_29585,N_27210,N_26645);
nand U29586 (N_29586,N_27855,N_26082);
and U29587 (N_29587,N_27743,N_27182);
nand U29588 (N_29588,N_27015,N_26076);
or U29589 (N_29589,N_27933,N_27367);
nand U29590 (N_29590,N_27500,N_27953);
or U29591 (N_29591,N_26209,N_26588);
nor U29592 (N_29592,N_26029,N_26739);
and U29593 (N_29593,N_27815,N_27787);
nor U29594 (N_29594,N_26383,N_27166);
or U29595 (N_29595,N_27437,N_27935);
and U29596 (N_29596,N_27816,N_26985);
or U29597 (N_29597,N_26631,N_26464);
and U29598 (N_29598,N_27736,N_27964);
or U29599 (N_29599,N_27463,N_27810);
nor U29600 (N_29600,N_27993,N_26945);
and U29601 (N_29601,N_27044,N_27503);
and U29602 (N_29602,N_27267,N_26026);
and U29603 (N_29603,N_27239,N_27177);
nand U29604 (N_29604,N_27278,N_26081);
nand U29605 (N_29605,N_26263,N_26920);
nand U29606 (N_29606,N_27901,N_27614);
or U29607 (N_29607,N_27669,N_26308);
and U29608 (N_29608,N_26434,N_27559);
or U29609 (N_29609,N_27676,N_26663);
xnor U29610 (N_29610,N_26184,N_26144);
nor U29611 (N_29611,N_26670,N_26823);
nor U29612 (N_29612,N_26389,N_26723);
nor U29613 (N_29613,N_27466,N_27588);
nand U29614 (N_29614,N_26197,N_26684);
xnor U29615 (N_29615,N_27166,N_27098);
nand U29616 (N_29616,N_26808,N_27506);
nand U29617 (N_29617,N_27321,N_27923);
nand U29618 (N_29618,N_27265,N_26838);
nand U29619 (N_29619,N_27854,N_26978);
nand U29620 (N_29620,N_26234,N_26448);
and U29621 (N_29621,N_27782,N_27771);
nand U29622 (N_29622,N_26093,N_26778);
and U29623 (N_29623,N_26113,N_27417);
xor U29624 (N_29624,N_26859,N_27815);
and U29625 (N_29625,N_26309,N_27032);
xor U29626 (N_29626,N_27022,N_27663);
xnor U29627 (N_29627,N_26214,N_26419);
nand U29628 (N_29628,N_26905,N_27743);
or U29629 (N_29629,N_26591,N_26002);
or U29630 (N_29630,N_27999,N_26660);
and U29631 (N_29631,N_26895,N_27188);
and U29632 (N_29632,N_26171,N_26598);
or U29633 (N_29633,N_26046,N_27688);
xnor U29634 (N_29634,N_26640,N_27459);
and U29635 (N_29635,N_26775,N_27848);
xor U29636 (N_29636,N_27782,N_26762);
xnor U29637 (N_29637,N_26734,N_26766);
or U29638 (N_29638,N_27762,N_26922);
nand U29639 (N_29639,N_26431,N_26291);
nor U29640 (N_29640,N_27120,N_26256);
and U29641 (N_29641,N_26315,N_26959);
or U29642 (N_29642,N_27806,N_27543);
and U29643 (N_29643,N_27825,N_26327);
and U29644 (N_29644,N_27823,N_27775);
and U29645 (N_29645,N_26277,N_27398);
and U29646 (N_29646,N_26180,N_27015);
xnor U29647 (N_29647,N_27363,N_27913);
and U29648 (N_29648,N_26092,N_26280);
xor U29649 (N_29649,N_26995,N_27347);
xor U29650 (N_29650,N_26236,N_26319);
and U29651 (N_29651,N_26735,N_27130);
xor U29652 (N_29652,N_26867,N_26099);
xor U29653 (N_29653,N_27899,N_27029);
nand U29654 (N_29654,N_27696,N_26653);
and U29655 (N_29655,N_26586,N_27571);
xnor U29656 (N_29656,N_26389,N_27553);
nand U29657 (N_29657,N_27220,N_26185);
nand U29658 (N_29658,N_26821,N_26097);
xor U29659 (N_29659,N_26630,N_26008);
xor U29660 (N_29660,N_26355,N_27654);
xnor U29661 (N_29661,N_26052,N_26939);
nand U29662 (N_29662,N_27787,N_26576);
and U29663 (N_29663,N_27564,N_27586);
and U29664 (N_29664,N_27079,N_27745);
xnor U29665 (N_29665,N_26467,N_26003);
nand U29666 (N_29666,N_27186,N_27429);
or U29667 (N_29667,N_26983,N_26531);
nor U29668 (N_29668,N_27592,N_27438);
nor U29669 (N_29669,N_27620,N_27122);
and U29670 (N_29670,N_26966,N_27120);
nand U29671 (N_29671,N_27850,N_27503);
nor U29672 (N_29672,N_27752,N_27371);
nor U29673 (N_29673,N_26867,N_27096);
nor U29674 (N_29674,N_27914,N_26097);
and U29675 (N_29675,N_27645,N_26260);
nand U29676 (N_29676,N_27832,N_27758);
nor U29677 (N_29677,N_27461,N_26559);
nand U29678 (N_29678,N_26928,N_27900);
or U29679 (N_29679,N_27368,N_27822);
nand U29680 (N_29680,N_26300,N_26407);
xor U29681 (N_29681,N_26182,N_27791);
xor U29682 (N_29682,N_26416,N_26570);
and U29683 (N_29683,N_26546,N_27629);
and U29684 (N_29684,N_27649,N_27218);
or U29685 (N_29685,N_27842,N_26619);
and U29686 (N_29686,N_27744,N_27598);
xor U29687 (N_29687,N_27799,N_27544);
or U29688 (N_29688,N_26679,N_26896);
nand U29689 (N_29689,N_27215,N_26068);
nand U29690 (N_29690,N_26419,N_27984);
or U29691 (N_29691,N_27048,N_27031);
xor U29692 (N_29692,N_27386,N_26254);
xnor U29693 (N_29693,N_27294,N_27123);
and U29694 (N_29694,N_26004,N_26307);
nor U29695 (N_29695,N_27532,N_27268);
or U29696 (N_29696,N_26581,N_27846);
nand U29697 (N_29697,N_26148,N_27039);
xnor U29698 (N_29698,N_27234,N_27622);
or U29699 (N_29699,N_26971,N_26946);
and U29700 (N_29700,N_26082,N_26837);
nand U29701 (N_29701,N_26763,N_26403);
xnor U29702 (N_29702,N_27819,N_27537);
nor U29703 (N_29703,N_27552,N_27884);
and U29704 (N_29704,N_26323,N_27537);
nor U29705 (N_29705,N_27067,N_26912);
or U29706 (N_29706,N_26627,N_27005);
or U29707 (N_29707,N_27218,N_26136);
and U29708 (N_29708,N_27345,N_27854);
or U29709 (N_29709,N_27525,N_27841);
and U29710 (N_29710,N_27750,N_26680);
nand U29711 (N_29711,N_26036,N_27395);
and U29712 (N_29712,N_27999,N_26296);
xor U29713 (N_29713,N_26250,N_26913);
nand U29714 (N_29714,N_27056,N_26127);
or U29715 (N_29715,N_27573,N_27477);
xor U29716 (N_29716,N_26900,N_27797);
nor U29717 (N_29717,N_26457,N_27432);
or U29718 (N_29718,N_26572,N_27394);
or U29719 (N_29719,N_26482,N_26397);
and U29720 (N_29720,N_27183,N_27050);
xor U29721 (N_29721,N_26102,N_26599);
or U29722 (N_29722,N_27100,N_26806);
or U29723 (N_29723,N_27333,N_27502);
and U29724 (N_29724,N_26491,N_26569);
and U29725 (N_29725,N_26035,N_26359);
nor U29726 (N_29726,N_27157,N_27334);
nor U29727 (N_29727,N_27389,N_27571);
xnor U29728 (N_29728,N_26192,N_27442);
or U29729 (N_29729,N_27751,N_26155);
nor U29730 (N_29730,N_27224,N_27425);
xnor U29731 (N_29731,N_26398,N_26763);
xor U29732 (N_29732,N_26392,N_26890);
or U29733 (N_29733,N_26804,N_26854);
nand U29734 (N_29734,N_27898,N_27458);
or U29735 (N_29735,N_26412,N_27880);
xnor U29736 (N_29736,N_26338,N_26559);
xor U29737 (N_29737,N_26536,N_26096);
nand U29738 (N_29738,N_26384,N_27852);
nor U29739 (N_29739,N_26305,N_26432);
and U29740 (N_29740,N_26410,N_26704);
or U29741 (N_29741,N_26150,N_27817);
nand U29742 (N_29742,N_26321,N_26767);
nor U29743 (N_29743,N_27890,N_26114);
or U29744 (N_29744,N_27084,N_26006);
nor U29745 (N_29745,N_26844,N_26705);
nand U29746 (N_29746,N_27618,N_26973);
nor U29747 (N_29747,N_27865,N_26617);
or U29748 (N_29748,N_26567,N_26787);
nor U29749 (N_29749,N_26593,N_26831);
or U29750 (N_29750,N_27357,N_27849);
nand U29751 (N_29751,N_26904,N_27962);
and U29752 (N_29752,N_27439,N_26980);
nand U29753 (N_29753,N_27605,N_27511);
and U29754 (N_29754,N_26670,N_27213);
or U29755 (N_29755,N_26573,N_27541);
nand U29756 (N_29756,N_26220,N_27348);
nand U29757 (N_29757,N_26701,N_26828);
nand U29758 (N_29758,N_26909,N_27016);
or U29759 (N_29759,N_27466,N_27853);
and U29760 (N_29760,N_26621,N_27137);
nand U29761 (N_29761,N_27644,N_26549);
and U29762 (N_29762,N_26703,N_26473);
or U29763 (N_29763,N_27254,N_27011);
or U29764 (N_29764,N_27821,N_27198);
xnor U29765 (N_29765,N_27389,N_27209);
and U29766 (N_29766,N_26147,N_27929);
and U29767 (N_29767,N_26955,N_27695);
xor U29768 (N_29768,N_26803,N_27485);
xnor U29769 (N_29769,N_27146,N_26925);
nand U29770 (N_29770,N_27652,N_27125);
and U29771 (N_29771,N_26677,N_27354);
xnor U29772 (N_29772,N_26736,N_26961);
nand U29773 (N_29773,N_27690,N_27594);
xor U29774 (N_29774,N_27856,N_27593);
nor U29775 (N_29775,N_27381,N_27725);
and U29776 (N_29776,N_27396,N_26854);
or U29777 (N_29777,N_27933,N_26693);
xnor U29778 (N_29778,N_27490,N_27310);
nand U29779 (N_29779,N_27705,N_27622);
nand U29780 (N_29780,N_26960,N_27853);
xor U29781 (N_29781,N_27684,N_26815);
or U29782 (N_29782,N_27213,N_27837);
xnor U29783 (N_29783,N_26033,N_27894);
nand U29784 (N_29784,N_26631,N_27444);
or U29785 (N_29785,N_27263,N_26611);
or U29786 (N_29786,N_27483,N_27786);
nor U29787 (N_29787,N_27918,N_27752);
nand U29788 (N_29788,N_27373,N_26142);
nand U29789 (N_29789,N_26809,N_27669);
nor U29790 (N_29790,N_27133,N_26308);
nand U29791 (N_29791,N_27642,N_26799);
or U29792 (N_29792,N_27280,N_26336);
or U29793 (N_29793,N_26201,N_27207);
nand U29794 (N_29794,N_27166,N_26205);
and U29795 (N_29795,N_27942,N_26838);
or U29796 (N_29796,N_26674,N_27952);
nand U29797 (N_29797,N_27661,N_27550);
nand U29798 (N_29798,N_27659,N_26219);
nor U29799 (N_29799,N_27490,N_27360);
or U29800 (N_29800,N_27421,N_27949);
and U29801 (N_29801,N_27347,N_26950);
nand U29802 (N_29802,N_27040,N_27162);
and U29803 (N_29803,N_27063,N_27887);
and U29804 (N_29804,N_27778,N_27601);
nor U29805 (N_29805,N_26885,N_27276);
nor U29806 (N_29806,N_26244,N_26928);
nor U29807 (N_29807,N_27314,N_27775);
xnor U29808 (N_29808,N_27245,N_27944);
xor U29809 (N_29809,N_27672,N_27518);
nor U29810 (N_29810,N_27993,N_26525);
xor U29811 (N_29811,N_26242,N_26549);
and U29812 (N_29812,N_27169,N_27957);
or U29813 (N_29813,N_27502,N_27187);
nand U29814 (N_29814,N_26619,N_27654);
nand U29815 (N_29815,N_27666,N_26186);
and U29816 (N_29816,N_27211,N_26877);
or U29817 (N_29817,N_27831,N_27499);
and U29818 (N_29818,N_27706,N_27003);
xnor U29819 (N_29819,N_27269,N_27388);
xor U29820 (N_29820,N_27313,N_27952);
nor U29821 (N_29821,N_26941,N_27733);
nor U29822 (N_29822,N_26856,N_27918);
and U29823 (N_29823,N_27572,N_27759);
or U29824 (N_29824,N_26597,N_27021);
xor U29825 (N_29825,N_27863,N_26776);
or U29826 (N_29826,N_26261,N_27115);
nand U29827 (N_29827,N_26957,N_27941);
xnor U29828 (N_29828,N_26714,N_27867);
xor U29829 (N_29829,N_26177,N_26179);
xor U29830 (N_29830,N_27412,N_27235);
nor U29831 (N_29831,N_27593,N_27866);
or U29832 (N_29832,N_27873,N_27720);
or U29833 (N_29833,N_26280,N_27343);
or U29834 (N_29834,N_27876,N_26622);
and U29835 (N_29835,N_26103,N_26274);
xnor U29836 (N_29836,N_27861,N_27842);
nand U29837 (N_29837,N_27771,N_27064);
nand U29838 (N_29838,N_26965,N_26164);
or U29839 (N_29839,N_26272,N_27484);
and U29840 (N_29840,N_26079,N_26513);
xor U29841 (N_29841,N_27985,N_27592);
xor U29842 (N_29842,N_26845,N_27594);
or U29843 (N_29843,N_27876,N_26845);
nand U29844 (N_29844,N_27324,N_26365);
nor U29845 (N_29845,N_26775,N_27545);
and U29846 (N_29846,N_26262,N_27513);
nor U29847 (N_29847,N_26030,N_26512);
xnor U29848 (N_29848,N_26433,N_26112);
and U29849 (N_29849,N_27420,N_27575);
nand U29850 (N_29850,N_27819,N_27441);
xor U29851 (N_29851,N_26530,N_27134);
and U29852 (N_29852,N_27545,N_27250);
and U29853 (N_29853,N_27108,N_26959);
xor U29854 (N_29854,N_27397,N_27606);
nor U29855 (N_29855,N_27513,N_27677);
xor U29856 (N_29856,N_27928,N_26637);
nor U29857 (N_29857,N_27076,N_26383);
nand U29858 (N_29858,N_26260,N_26224);
nor U29859 (N_29859,N_26251,N_26517);
and U29860 (N_29860,N_27410,N_26738);
xnor U29861 (N_29861,N_27441,N_26495);
nor U29862 (N_29862,N_27392,N_26195);
xor U29863 (N_29863,N_26746,N_27853);
nor U29864 (N_29864,N_27255,N_26975);
nor U29865 (N_29865,N_27184,N_27104);
and U29866 (N_29866,N_26367,N_26747);
or U29867 (N_29867,N_27201,N_27425);
xor U29868 (N_29868,N_26048,N_26347);
xor U29869 (N_29869,N_27143,N_27480);
xor U29870 (N_29870,N_27770,N_26819);
and U29871 (N_29871,N_26159,N_27565);
nand U29872 (N_29872,N_26449,N_27229);
xor U29873 (N_29873,N_26935,N_27996);
nor U29874 (N_29874,N_27143,N_27460);
xnor U29875 (N_29875,N_27640,N_26489);
xor U29876 (N_29876,N_26956,N_26152);
nor U29877 (N_29877,N_26079,N_26013);
xor U29878 (N_29878,N_27671,N_27698);
xor U29879 (N_29879,N_26837,N_27268);
xor U29880 (N_29880,N_26219,N_26892);
nand U29881 (N_29881,N_26434,N_27315);
nand U29882 (N_29882,N_26561,N_26824);
or U29883 (N_29883,N_27569,N_27589);
nor U29884 (N_29884,N_27169,N_26461);
xor U29885 (N_29885,N_26384,N_27386);
and U29886 (N_29886,N_27788,N_27400);
and U29887 (N_29887,N_26968,N_27578);
nor U29888 (N_29888,N_26324,N_27496);
nor U29889 (N_29889,N_26893,N_26108);
nor U29890 (N_29890,N_26735,N_27602);
xor U29891 (N_29891,N_27241,N_26091);
xor U29892 (N_29892,N_26994,N_26369);
nor U29893 (N_29893,N_26380,N_26177);
nor U29894 (N_29894,N_26498,N_26912);
or U29895 (N_29895,N_26666,N_27456);
or U29896 (N_29896,N_26313,N_27280);
or U29897 (N_29897,N_27218,N_27443);
or U29898 (N_29898,N_27969,N_27590);
nand U29899 (N_29899,N_26081,N_26533);
xor U29900 (N_29900,N_27640,N_27806);
nand U29901 (N_29901,N_26326,N_26789);
xnor U29902 (N_29902,N_26668,N_26329);
and U29903 (N_29903,N_26416,N_26079);
nand U29904 (N_29904,N_27729,N_26657);
nand U29905 (N_29905,N_26524,N_27552);
or U29906 (N_29906,N_26882,N_27671);
and U29907 (N_29907,N_27538,N_27457);
nor U29908 (N_29908,N_27724,N_27093);
or U29909 (N_29909,N_26196,N_27532);
or U29910 (N_29910,N_27191,N_27557);
or U29911 (N_29911,N_27296,N_27354);
nand U29912 (N_29912,N_26339,N_27964);
xnor U29913 (N_29913,N_27772,N_27623);
xor U29914 (N_29914,N_27386,N_26996);
nand U29915 (N_29915,N_27485,N_26140);
and U29916 (N_29916,N_27771,N_26459);
or U29917 (N_29917,N_26746,N_26147);
or U29918 (N_29918,N_27097,N_27483);
nand U29919 (N_29919,N_27430,N_26838);
or U29920 (N_29920,N_27314,N_27261);
xnor U29921 (N_29921,N_27602,N_27235);
and U29922 (N_29922,N_26187,N_26359);
nor U29923 (N_29923,N_26294,N_27955);
xor U29924 (N_29924,N_26059,N_27987);
or U29925 (N_29925,N_27405,N_26155);
nand U29926 (N_29926,N_26089,N_27957);
nor U29927 (N_29927,N_27360,N_26271);
or U29928 (N_29928,N_27429,N_26476);
nand U29929 (N_29929,N_27511,N_26382);
nand U29930 (N_29930,N_26006,N_26929);
nand U29931 (N_29931,N_27572,N_27914);
and U29932 (N_29932,N_26665,N_26946);
nor U29933 (N_29933,N_27164,N_26133);
xnor U29934 (N_29934,N_26049,N_27689);
nand U29935 (N_29935,N_26814,N_27779);
nand U29936 (N_29936,N_26378,N_27474);
nor U29937 (N_29937,N_26928,N_27329);
nor U29938 (N_29938,N_27459,N_26125);
nand U29939 (N_29939,N_27371,N_27010);
nand U29940 (N_29940,N_26851,N_26682);
nor U29941 (N_29941,N_26917,N_26829);
nor U29942 (N_29942,N_27797,N_26731);
xnor U29943 (N_29943,N_27358,N_27419);
nor U29944 (N_29944,N_26605,N_27406);
or U29945 (N_29945,N_27808,N_26962);
nor U29946 (N_29946,N_26472,N_27971);
xor U29947 (N_29947,N_26532,N_26895);
xor U29948 (N_29948,N_26771,N_27287);
and U29949 (N_29949,N_26571,N_27967);
nor U29950 (N_29950,N_27596,N_27500);
and U29951 (N_29951,N_27518,N_26979);
nor U29952 (N_29952,N_27811,N_27349);
xor U29953 (N_29953,N_26938,N_27396);
nand U29954 (N_29954,N_26294,N_26526);
xor U29955 (N_29955,N_26553,N_27000);
or U29956 (N_29956,N_26511,N_27193);
xnor U29957 (N_29957,N_26176,N_26955);
and U29958 (N_29958,N_26892,N_26099);
and U29959 (N_29959,N_27728,N_26486);
nand U29960 (N_29960,N_26138,N_27920);
and U29961 (N_29961,N_27161,N_27922);
nor U29962 (N_29962,N_26381,N_26204);
or U29963 (N_29963,N_26127,N_27008);
xor U29964 (N_29964,N_27140,N_26634);
or U29965 (N_29965,N_27551,N_26364);
xor U29966 (N_29966,N_26746,N_26687);
or U29967 (N_29967,N_26639,N_27194);
xor U29968 (N_29968,N_27041,N_26578);
and U29969 (N_29969,N_27265,N_27889);
or U29970 (N_29970,N_27595,N_27295);
nand U29971 (N_29971,N_27704,N_27606);
and U29972 (N_29972,N_26227,N_27582);
nor U29973 (N_29973,N_27322,N_26184);
or U29974 (N_29974,N_26260,N_27722);
xnor U29975 (N_29975,N_27202,N_26669);
or U29976 (N_29976,N_27651,N_27127);
and U29977 (N_29977,N_26600,N_27735);
nand U29978 (N_29978,N_26214,N_27915);
and U29979 (N_29979,N_26615,N_26559);
and U29980 (N_29980,N_26576,N_26409);
and U29981 (N_29981,N_27767,N_27593);
nor U29982 (N_29982,N_26095,N_27406);
nand U29983 (N_29983,N_27878,N_27561);
or U29984 (N_29984,N_26596,N_27624);
nand U29985 (N_29985,N_26224,N_27071);
xor U29986 (N_29986,N_27407,N_27219);
nand U29987 (N_29987,N_26504,N_27843);
nand U29988 (N_29988,N_27992,N_26892);
and U29989 (N_29989,N_27920,N_27877);
and U29990 (N_29990,N_26988,N_27612);
or U29991 (N_29991,N_27106,N_26058);
nand U29992 (N_29992,N_26688,N_26286);
nor U29993 (N_29993,N_27600,N_26266);
and U29994 (N_29994,N_27555,N_26671);
nor U29995 (N_29995,N_26734,N_26298);
and U29996 (N_29996,N_27449,N_27851);
nor U29997 (N_29997,N_26869,N_26240);
and U29998 (N_29998,N_26653,N_27783);
nand U29999 (N_29999,N_26730,N_26600);
or U30000 (N_30000,N_29439,N_28959);
or U30001 (N_30001,N_28301,N_29726);
nor U30002 (N_30002,N_29515,N_28886);
nor U30003 (N_30003,N_29608,N_29480);
xor U30004 (N_30004,N_29253,N_28958);
xnor U30005 (N_30005,N_29484,N_28269);
nand U30006 (N_30006,N_29375,N_28387);
and U30007 (N_30007,N_28827,N_28477);
and U30008 (N_30008,N_29891,N_28713);
nor U30009 (N_30009,N_28492,N_28235);
nand U30010 (N_30010,N_29872,N_28519);
or U30011 (N_30011,N_28773,N_29141);
and U30012 (N_30012,N_29202,N_29887);
nand U30013 (N_30013,N_28365,N_29045);
or U30014 (N_30014,N_29605,N_29348);
and U30015 (N_30015,N_28249,N_28098);
xnor U30016 (N_30016,N_29241,N_29532);
or U30017 (N_30017,N_28429,N_28044);
xnor U30018 (N_30018,N_29182,N_28094);
nor U30019 (N_30019,N_29128,N_29495);
xnor U30020 (N_30020,N_29155,N_29234);
and U30021 (N_30021,N_29819,N_28496);
nor U30022 (N_30022,N_29007,N_28270);
nand U30023 (N_30023,N_28470,N_29340);
nand U30024 (N_30024,N_28107,N_28495);
nand U30025 (N_30025,N_28005,N_28167);
or U30026 (N_30026,N_28523,N_29871);
or U30027 (N_30027,N_28454,N_29860);
nand U30028 (N_30028,N_28314,N_28358);
or U30029 (N_30029,N_29000,N_28381);
xnor U30030 (N_30030,N_28423,N_28146);
nand U30031 (N_30031,N_29972,N_29279);
nor U30032 (N_30032,N_28040,N_29077);
nand U30033 (N_30033,N_28086,N_29165);
nor U30034 (N_30034,N_28196,N_29440);
or U30035 (N_30035,N_28426,N_28979);
xnor U30036 (N_30036,N_29643,N_29514);
nor U30037 (N_30037,N_28517,N_28809);
xor U30038 (N_30038,N_28066,N_29276);
nand U30039 (N_30039,N_29689,N_29765);
nor U30040 (N_30040,N_28376,N_29893);
xnor U30041 (N_30041,N_28869,N_28710);
or U30042 (N_30042,N_28067,N_29042);
and U30043 (N_30043,N_29038,N_29199);
nor U30044 (N_30044,N_29858,N_29508);
and U30045 (N_30045,N_28821,N_28490);
nor U30046 (N_30046,N_29296,N_28219);
and U30047 (N_30047,N_28500,N_28360);
and U30048 (N_30048,N_29210,N_29470);
xor U30049 (N_30049,N_29846,N_28532);
or U30050 (N_30050,N_28109,N_28625);
and U30051 (N_30051,N_28138,N_28306);
nand U30052 (N_30052,N_28339,N_29447);
xnor U30053 (N_30053,N_29705,N_28475);
xor U30054 (N_30054,N_28925,N_29719);
xnor U30055 (N_30055,N_29506,N_28199);
nor U30056 (N_30056,N_29397,N_29131);
and U30057 (N_30057,N_29570,N_29637);
xor U30058 (N_30058,N_28753,N_29776);
or U30059 (N_30059,N_28291,N_28616);
nor U30060 (N_30060,N_28657,N_29333);
nor U30061 (N_30061,N_28079,N_29051);
nand U30062 (N_30062,N_28082,N_28168);
or U30063 (N_30063,N_29378,N_28284);
or U30064 (N_30064,N_29496,N_29524);
and U30065 (N_30065,N_28329,N_28722);
or U30066 (N_30066,N_28647,N_29729);
or U30067 (N_30067,N_28289,N_28231);
nand U30068 (N_30068,N_29980,N_28015);
nor U30069 (N_30069,N_29897,N_28046);
and U30070 (N_30070,N_28059,N_28414);
nor U30071 (N_30071,N_29099,N_28734);
nor U30072 (N_30072,N_28090,N_29256);
nor U30073 (N_30073,N_29335,N_28285);
or U30074 (N_30074,N_29625,N_28084);
xnor U30075 (N_30075,N_29271,N_29393);
and U30076 (N_30076,N_28917,N_28264);
xnor U30077 (N_30077,N_28355,N_29485);
nor U30078 (N_30078,N_28580,N_28891);
xor U30079 (N_30079,N_28161,N_28882);
nand U30080 (N_30080,N_28690,N_29391);
and U30081 (N_30081,N_28350,N_28608);
nand U30082 (N_30082,N_28293,N_28334);
nor U30083 (N_30083,N_29292,N_28451);
nand U30084 (N_30084,N_29629,N_28413);
and U30085 (N_30085,N_29807,N_29108);
or U30086 (N_30086,N_29794,N_29655);
nor U30087 (N_30087,N_28212,N_28184);
nand U30088 (N_30088,N_29682,N_29015);
nor U30089 (N_30089,N_29565,N_29908);
nand U30090 (N_30090,N_28754,N_28404);
xor U30091 (N_30091,N_28386,N_29760);
or U30092 (N_30092,N_28771,N_29394);
nand U30093 (N_30093,N_28650,N_29513);
nand U30094 (N_30094,N_29081,N_29146);
or U30095 (N_30095,N_29620,N_28745);
or U30096 (N_30096,N_29002,N_28210);
or U30097 (N_30097,N_28047,N_28998);
xnor U30098 (N_30098,N_29947,N_29774);
nand U30099 (N_30099,N_29139,N_28342);
xor U30100 (N_30100,N_28063,N_28839);
and U30101 (N_30101,N_28026,N_28361);
nor U30102 (N_30102,N_28707,N_29886);
xnor U30103 (N_30103,N_28845,N_29069);
or U30104 (N_30104,N_28461,N_29206);
nor U30105 (N_30105,N_28163,N_29057);
nor U30106 (N_30106,N_29536,N_28281);
nand U30107 (N_30107,N_29085,N_29788);
xor U30108 (N_30108,N_29553,N_28782);
nor U30109 (N_30109,N_28195,N_28551);
and U30110 (N_30110,N_29677,N_28788);
or U30111 (N_30111,N_29734,N_29597);
xor U30112 (N_30112,N_29992,N_29429);
nand U30113 (N_30113,N_29885,N_28427);
nand U30114 (N_30114,N_29066,N_28016);
xor U30115 (N_30115,N_29461,N_28397);
nand U30116 (N_30116,N_28106,N_29414);
or U30117 (N_30117,N_29670,N_29104);
nand U30118 (N_30118,N_29218,N_29534);
or U30119 (N_30119,N_29548,N_28250);
xnor U30120 (N_30120,N_28543,N_29159);
xor U30121 (N_30121,N_29387,N_28364);
nand U30122 (N_30122,N_28993,N_28525);
or U30123 (N_30123,N_28223,N_29631);
xor U30124 (N_30124,N_29347,N_29249);
nand U30125 (N_30125,N_28419,N_28145);
and U30126 (N_30126,N_28022,N_28966);
nor U30127 (N_30127,N_28021,N_28031);
or U30128 (N_30128,N_29328,N_28324);
xnor U30129 (N_30129,N_28858,N_29339);
and U30130 (N_30130,N_28879,N_29309);
nor U30131 (N_30131,N_28356,N_28649);
nand U30132 (N_30132,N_29849,N_29418);
and U30133 (N_30133,N_29476,N_28240);
nor U30134 (N_30134,N_29766,N_29715);
nand U30135 (N_30135,N_28946,N_28550);
or U30136 (N_30136,N_29315,N_29137);
nand U30137 (N_30137,N_28818,N_29147);
xnor U30138 (N_30138,N_29498,N_29733);
and U30139 (N_30139,N_29317,N_28279);
xor U30140 (N_30140,N_29435,N_28677);
and U30141 (N_30141,N_29410,N_28478);
nand U30142 (N_30142,N_28582,N_28510);
nor U30143 (N_30143,N_29351,N_28153);
or U30144 (N_30144,N_29436,N_28759);
nand U30145 (N_30145,N_28631,N_29289);
xor U30146 (N_30146,N_28081,N_28417);
xnor U30147 (N_30147,N_29178,N_29406);
and U30148 (N_30148,N_28348,N_29877);
or U30149 (N_30149,N_28230,N_28542);
nor U30150 (N_30150,N_29644,N_29260);
and U30151 (N_30151,N_29985,N_28033);
xnor U30152 (N_30152,N_28635,N_29583);
nor U30153 (N_30153,N_28133,N_29955);
xnor U30154 (N_30154,N_28598,N_29696);
nor U30155 (N_30155,N_29662,N_29923);
xnor U30156 (N_30156,N_28848,N_28989);
and U30157 (N_30157,N_29041,N_28157);
xor U30158 (N_30158,N_28290,N_29832);
and U30159 (N_30159,N_29905,N_29493);
nor U30160 (N_30160,N_29995,N_28203);
nand U30161 (N_30161,N_29721,N_28434);
or U30162 (N_30162,N_29477,N_28276);
xnor U30163 (N_30163,N_28405,N_28296);
or U30164 (N_30164,N_28910,N_29901);
nor U30165 (N_30165,N_28844,N_28069);
and U30166 (N_30166,N_28758,N_28586);
and U30167 (N_30167,N_28854,N_28257);
nand U30168 (N_30168,N_28992,N_28904);
and U30169 (N_30169,N_29049,N_29373);
or U30170 (N_30170,N_29143,N_29633);
nand U30171 (N_30171,N_28064,N_29842);
xnor U30172 (N_30172,N_28062,N_28486);
or U30173 (N_30173,N_29941,N_29599);
and U30174 (N_30174,N_28988,N_28847);
nor U30175 (N_30175,N_28905,N_28487);
and U30176 (N_30176,N_29195,N_28981);
nor U30177 (N_30177,N_29227,N_29748);
xnor U30178 (N_30178,N_28102,N_28703);
nor U30179 (N_30179,N_29295,N_29502);
or U30180 (N_30180,N_29857,N_29151);
or U30181 (N_30181,N_29213,N_28013);
or U30182 (N_30182,N_29806,N_28595);
or U30183 (N_30183,N_28795,N_28530);
and U30184 (N_30184,N_28114,N_28641);
nor U30185 (N_30185,N_29463,N_28406);
or U30186 (N_30186,N_29148,N_29505);
and U30187 (N_30187,N_29430,N_29713);
nand U30188 (N_30188,N_29097,N_29831);
xnor U30189 (N_30189,N_28627,N_29869);
nor U30190 (N_30190,N_29086,N_29065);
xnor U30191 (N_30191,N_28846,N_28328);
and U30192 (N_30192,N_28258,N_29672);
nor U30193 (N_30193,N_28842,N_29003);
nor U30194 (N_30194,N_29685,N_29878);
and U30195 (N_30195,N_29699,N_28126);
nor U30196 (N_30196,N_28855,N_28592);
xor U30197 (N_30197,N_28392,N_29545);
xnor U30198 (N_30198,N_29984,N_29230);
nor U30199 (N_30199,N_29198,N_29735);
nand U30200 (N_30200,N_28695,N_29243);
xor U30201 (N_30201,N_28148,N_28225);
nand U30202 (N_30202,N_29645,N_29327);
nor U30203 (N_30203,N_29910,N_28604);
nand U30204 (N_30204,N_28103,N_29755);
nor U30205 (N_30205,N_28460,N_28170);
and U30206 (N_30206,N_29674,N_28780);
or U30207 (N_30207,N_29044,N_29013);
nand U30208 (N_30208,N_29071,N_28325);
and U30209 (N_30209,N_29825,N_28778);
nand U30210 (N_30210,N_29883,N_28473);
xnor U30211 (N_30211,N_29456,N_28154);
and U30212 (N_30212,N_29314,N_29360);
or U30213 (N_30213,N_28048,N_28077);
nor U30214 (N_30214,N_28915,N_28574);
nor U30215 (N_30215,N_29889,N_29529);
nor U30216 (N_30216,N_28330,N_29591);
xnor U30217 (N_30217,N_29371,N_28131);
nand U30218 (N_30218,N_28733,N_28425);
or U30219 (N_30219,N_28554,N_28685);
xnor U30220 (N_30220,N_29092,N_29839);
and U30221 (N_30221,N_28714,N_28481);
nand U30222 (N_30222,N_29403,N_28171);
nand U30223 (N_30223,N_28036,N_28137);
nand U30224 (N_30224,N_28420,N_29744);
nand U30225 (N_30225,N_29105,N_29490);
xnor U30226 (N_30226,N_29337,N_29163);
nand U30227 (N_30227,N_29184,N_28516);
nor U30228 (N_30228,N_28765,N_29288);
nand U30229 (N_30229,N_29727,N_29422);
or U30230 (N_30230,N_29700,N_28372);
or U30231 (N_30231,N_29462,N_29455);
or U30232 (N_30232,N_28666,N_29464);
and U30233 (N_30233,N_28415,N_28252);
or U30234 (N_30234,N_28205,N_29268);
xor U30235 (N_30235,N_28180,N_29415);
and U30236 (N_30236,N_29356,N_29746);
xnor U30237 (N_30237,N_29121,N_29709);
nand U30238 (N_30238,N_28874,N_28508);
and U30239 (N_30239,N_28615,N_29522);
and U30240 (N_30240,N_28065,N_28876);
nor U30241 (N_30241,N_29659,N_29736);
and U30242 (N_30242,N_29623,N_28401);
nor U30243 (N_30243,N_29229,N_29789);
nor U30244 (N_30244,N_28468,N_28819);
or U30245 (N_30245,N_28441,N_29959);
xor U30246 (N_30246,N_28295,N_28136);
or U30247 (N_30247,N_29906,N_28605);
nand U30248 (N_30248,N_28341,N_29377);
nor U30249 (N_30249,N_28175,N_29982);
xnor U30250 (N_30250,N_29293,N_29158);
nand U30251 (N_30251,N_29123,N_29445);
nor U30252 (N_30252,N_28242,N_28499);
nand U30253 (N_30253,N_29718,N_28472);
and U30254 (N_30254,N_28172,N_28462);
and U30255 (N_30255,N_29988,N_28977);
nor U30256 (N_30256,N_28357,N_28318);
or U30257 (N_30257,N_29650,N_28061);
xor U30258 (N_30258,N_28880,N_29424);
xor U30259 (N_30259,N_28911,N_29413);
and U30260 (N_30260,N_28467,N_28370);
xor U30261 (N_30261,N_29177,N_29334);
or U30262 (N_30262,N_29343,N_29466);
nor U30263 (N_30263,N_28347,N_28345);
nand U30264 (N_30264,N_28980,N_29740);
xor U30265 (N_30265,N_29399,N_29060);
nor U30266 (N_30266,N_29585,N_28101);
or U30267 (N_30267,N_29575,N_29329);
and U30268 (N_30268,N_28453,N_29054);
and U30269 (N_30269,N_29639,N_29215);
and U30270 (N_30270,N_29921,N_29129);
nor U30271 (N_30271,N_29386,N_28158);
nand U30272 (N_30272,N_28315,N_29946);
nor U30273 (N_30273,N_28117,N_29795);
xnor U30274 (N_30274,N_28333,N_28561);
and U30275 (N_30275,N_29005,N_29683);
nor U30276 (N_30276,N_29636,N_28099);
xnor U30277 (N_30277,N_29528,N_29107);
xor U30278 (N_30278,N_28730,N_29568);
nor U30279 (N_30279,N_29714,N_29773);
or U30280 (N_30280,N_29813,N_28027);
nor U30281 (N_30281,N_28632,N_28897);
nor U30282 (N_30282,N_29702,N_29242);
and U30283 (N_30283,N_29126,N_29306);
or U30284 (N_30284,N_29196,N_29179);
nor U30285 (N_30285,N_28791,N_29366);
nor U30286 (N_30286,N_28783,N_28907);
or U30287 (N_30287,N_28379,N_28952);
xnor U30288 (N_30288,N_29628,N_29352);
or U30289 (N_30289,N_29176,N_28954);
and U30290 (N_30290,N_28676,N_28179);
xor U30291 (N_30291,N_29706,N_28590);
nand U30292 (N_30292,N_29257,N_29067);
or U30293 (N_30293,N_28058,N_29321);
or U30294 (N_30294,N_28121,N_28857);
or U30295 (N_30295,N_28929,N_29987);
and U30296 (N_30296,N_29364,N_28505);
nor U30297 (N_30297,N_29149,N_28964);
or U30298 (N_30298,N_29687,N_29106);
and U30299 (N_30299,N_29816,N_28150);
nor U30300 (N_30300,N_29757,N_28698);
nor U30301 (N_30301,N_28255,N_28803);
nor U30302 (N_30302,N_28007,N_28261);
nor U30303 (N_30303,N_29965,N_28883);
and U30304 (N_30304,N_28226,N_28008);
or U30305 (N_30305,N_28411,N_29688);
and U30306 (N_30306,N_29549,N_28866);
and U30307 (N_30307,N_28772,N_28200);
or U30308 (N_30308,N_28385,N_29226);
xnor U30309 (N_30309,N_29667,N_28262);
nor U30310 (N_30310,N_29861,N_29973);
and U30311 (N_30311,N_28458,N_28547);
or U30312 (N_30312,N_29142,N_29854);
nor U30313 (N_30313,N_28994,N_29324);
nand U30314 (N_30314,N_28972,N_28057);
or U30315 (N_30315,N_29465,N_28936);
and U30316 (N_30316,N_29547,N_29018);
or U30317 (N_30317,N_28321,N_28599);
or U30318 (N_30318,N_28237,N_28909);
nand U30319 (N_30319,N_28535,N_29815);
or U30320 (N_30320,N_29269,N_29826);
nor U30321 (N_30321,N_28719,N_28646);
nor U30322 (N_30322,N_28060,N_29516);
or U30323 (N_30323,N_28528,N_29050);
nand U30324 (N_30324,N_29951,N_29283);
xor U30325 (N_30325,N_29392,N_28840);
nor U30326 (N_30326,N_28366,N_29090);
nor U30327 (N_30327,N_28691,N_29187);
nand U30328 (N_30328,N_28924,N_29851);
nand U30329 (N_30329,N_28878,N_28752);
nand U30330 (N_30330,N_29879,N_29383);
nor U30331 (N_30331,N_29517,N_29952);
or U30332 (N_30332,N_29974,N_29473);
nand U30333 (N_30333,N_28524,N_29824);
nand U30334 (N_30334,N_28436,N_28667);
nand U30335 (N_30335,N_29079,N_29423);
or U30336 (N_30336,N_29244,N_28254);
nand U30337 (N_30337,N_28147,N_29856);
nor U30338 (N_30338,N_28684,N_29690);
and U30339 (N_30339,N_29847,N_29759);
or U30340 (N_30340,N_29023,N_28232);
or U30341 (N_30341,N_29938,N_28479);
and U30342 (N_30342,N_29953,N_28642);
nor U30343 (N_30343,N_28830,N_29061);
nand U30344 (N_30344,N_29053,N_28286);
or U30345 (N_30345,N_28618,N_28011);
nor U30346 (N_30346,N_28653,N_29821);
nand U30347 (N_30347,N_29040,N_29780);
and U30348 (N_30348,N_29494,N_28697);
and U30349 (N_30349,N_28004,N_29431);
nand U30350 (N_30350,N_28800,N_28159);
and U30351 (N_30351,N_28020,N_29103);
nor U30352 (N_30352,N_29501,N_29756);
and U30353 (N_30353,N_29267,N_29749);
or U30354 (N_30354,N_28430,N_28798);
and U30355 (N_30355,N_29619,N_28545);
nand U30356 (N_30356,N_28310,N_29512);
or U30357 (N_30357,N_29754,N_28645);
nand U30358 (N_30358,N_29595,N_28587);
and U30359 (N_30359,N_29338,N_29741);
nand U30360 (N_30360,N_28521,N_28579);
or U30361 (N_30361,N_28197,N_29072);
nand U30362 (N_30362,N_28828,N_28096);
nor U30363 (N_30363,N_29835,N_28444);
nand U30364 (N_30364,N_28287,N_28512);
or U30365 (N_30365,N_28997,N_29526);
nand U30366 (N_30366,N_29382,N_28322);
or U30367 (N_30367,N_28610,N_29991);
and U30368 (N_30368,N_28476,N_28566);
or U30369 (N_30369,N_28422,N_28556);
or U30370 (N_30370,N_29245,N_29312);
xor U30371 (N_30371,N_28999,N_28974);
and U30372 (N_30372,N_28089,N_28332);
nand U30373 (N_30373,N_28140,N_29634);
nand U30374 (N_30374,N_29036,N_29747);
and U30375 (N_30375,N_28811,N_29660);
and U30376 (N_30376,N_28198,N_29926);
and U30377 (N_30377,N_28820,N_29864);
and U30378 (N_30378,N_28326,N_29238);
xor U30379 (N_30379,N_29273,N_28921);
xor U30380 (N_30380,N_28841,N_29668);
and U30381 (N_30381,N_29745,N_29829);
xnor U30382 (N_30382,N_29302,N_29409);
nor U30383 (N_30383,N_28243,N_29627);
xor U30384 (N_30384,N_29875,N_29384);
xnor U30385 (N_30385,N_28045,N_28637);
nand U30386 (N_30386,N_28986,N_29350);
nand U30387 (N_30387,N_29913,N_29948);
or U30388 (N_30388,N_29262,N_28251);
nor U30389 (N_30389,N_29607,N_28307);
and U30390 (N_30390,N_28620,N_28459);
or U30391 (N_30391,N_28228,N_29618);
nor U30392 (N_30392,N_28894,N_28648);
and U30393 (N_30393,N_28097,N_28693);
nor U30394 (N_30394,N_29642,N_28544);
and U30395 (N_30395,N_28686,N_28678);
nand U30396 (N_30396,N_29914,N_29232);
or U30397 (N_30397,N_28786,N_28222);
xor U30398 (N_30398,N_28832,N_28456);
nand U30399 (N_30399,N_28041,N_28119);
xnor U30400 (N_30400,N_29786,N_29640);
nand U30401 (N_30401,N_28323,N_28626);
nor U30402 (N_30402,N_28211,N_28573);
nand U30403 (N_30403,N_29110,N_29311);
nand U30404 (N_30404,N_28527,N_29820);
nor U30405 (N_30405,N_28120,N_29400);
nand U30406 (N_30406,N_29657,N_29596);
or U30407 (N_30407,N_28278,N_28564);
and U30408 (N_30408,N_28633,N_28541);
or U30409 (N_30409,N_28629,N_28221);
and U30410 (N_30410,N_29589,N_28139);
nor U30411 (N_30411,N_29742,N_29222);
and U30412 (N_30412,N_28229,N_29421);
nor U30413 (N_30413,N_28263,N_28216);
nand U30414 (N_30414,N_29162,N_29100);
nor U30415 (N_30415,N_28607,N_28560);
xnor U30416 (N_30416,N_29573,N_28091);
nand U30417 (N_30417,N_29183,N_29963);
or U30418 (N_30418,N_28515,N_28283);
nor U30419 (N_30419,N_28070,N_29933);
and U30420 (N_30420,N_29303,N_29537);
nor U30421 (N_30421,N_29358,N_29758);
or U30422 (N_30422,N_29248,N_29033);
or U30423 (N_30423,N_29880,N_29566);
and U30424 (N_30424,N_28399,N_29446);
and U30425 (N_30425,N_29544,N_28142);
and U30426 (N_30426,N_28207,N_29250);
xor U30427 (N_30427,N_29937,N_29367);
and U30428 (N_30428,N_29792,N_29986);
nor U30429 (N_30429,N_29801,N_29161);
nand U30430 (N_30430,N_29658,N_28352);
and U30431 (N_30431,N_29990,N_28856);
nand U30432 (N_30432,N_29978,N_29876);
xnor U30433 (N_30433,N_29535,N_28054);
nor U30434 (N_30434,N_28680,N_28371);
xnor U30435 (N_30435,N_28639,N_28884);
xnor U30436 (N_30436,N_28968,N_29592);
xor U30437 (N_30437,N_29322,N_29433);
nand U30438 (N_30438,N_28944,N_29144);
and U30439 (N_30439,N_28751,N_28181);
nor U30440 (N_30440,N_28439,N_29388);
nor U30441 (N_30441,N_28937,N_28337);
nor U30442 (N_30442,N_29088,N_29127);
nor U30443 (N_30443,N_28973,N_28238);
and U30444 (N_30444,N_29428,N_28538);
xor U30445 (N_30445,N_29203,N_28449);
nor U30446 (N_30446,N_29796,N_28675);
nand U30447 (N_30447,N_29977,N_29345);
and U30448 (N_30448,N_28717,N_29219);
nand U30449 (N_30449,N_29381,N_29724);
and U30450 (N_30450,N_29416,N_28617);
or U30451 (N_30451,N_28012,N_29940);
nor U30452 (N_30452,N_28292,N_28087);
and U30453 (N_30453,N_28178,N_29174);
nor U30454 (N_30454,N_28890,N_28346);
nor U30455 (N_30455,N_28723,N_29481);
xor U30456 (N_30456,N_29453,N_28732);
nor U30457 (N_30457,N_28644,N_28398);
nand U30458 (N_30458,N_29584,N_29420);
and U30459 (N_30459,N_29220,N_29693);
xnor U30460 (N_30460,N_28234,N_28726);
and U30461 (N_30461,N_28578,N_29169);
and U30462 (N_30462,N_28881,N_29609);
and U30463 (N_30463,N_28002,N_29654);
xor U30464 (N_30464,N_29800,N_28735);
xnor U30465 (N_30465,N_28068,N_29679);
nand U30466 (N_30466,N_28297,N_28796);
or U30467 (N_30467,N_28768,N_29047);
xnor U30468 (N_30468,N_29647,N_28540);
and U30469 (N_30469,N_29027,N_28962);
nand U30470 (N_30470,N_29567,N_28493);
xnor U30471 (N_30471,N_29942,N_28038);
nor U30472 (N_30472,N_29703,N_29450);
nand U30473 (N_30473,N_29925,N_29945);
xnor U30474 (N_30474,N_28995,N_28849);
nor U30475 (N_30475,N_28851,N_29641);
xnor U30476 (N_30476,N_28706,N_29094);
nand U30477 (N_30477,N_29785,N_29207);
nor U30478 (N_30478,N_28437,N_28865);
or U30479 (N_30479,N_28961,N_29361);
and U30480 (N_30480,N_28491,N_29068);
xnor U30481 (N_30481,N_28764,N_29332);
nor U30482 (N_30482,N_29298,N_28185);
xnor U30483 (N_30483,N_28950,N_28236);
and U30484 (N_30484,N_29598,N_29770);
xor U30485 (N_30485,N_28665,N_29290);
xnor U30486 (N_30486,N_29474,N_29564);
nor U30487 (N_30487,N_29280,N_28447);
or U30488 (N_30488,N_29472,N_28656);
or U30489 (N_30489,N_29853,N_29852);
and U30490 (N_30490,N_28835,N_28770);
or U30491 (N_30491,N_28448,N_28265);
nand U30492 (N_30492,N_28017,N_28662);
or U30493 (N_30493,N_29927,N_28702);
nor U30494 (N_30494,N_29881,N_29855);
nand U30495 (N_30495,N_28509,N_28531);
and U30496 (N_30496,N_28721,N_28609);
nand U30497 (N_30497,N_29827,N_28930);
and U30498 (N_30498,N_29936,N_28497);
xor U30499 (N_30499,N_28025,N_29405);
and U30500 (N_30500,N_29622,N_29888);
xnor U30501 (N_30501,N_29153,N_28708);
or U30502 (N_30502,N_29771,N_28728);
nor U30503 (N_30503,N_29803,N_28947);
or U30504 (N_30504,N_28368,N_29114);
and U30505 (N_30505,N_29419,N_28400);
nor U30506 (N_30506,N_28450,N_29621);
xnor U30507 (N_30507,N_28034,N_28273);
xor U30508 (N_30508,N_29525,N_28867);
xnor U30509 (N_30509,N_28654,N_29095);
and U30510 (N_30510,N_29164,N_29379);
or U30511 (N_30511,N_29341,N_28100);
nand U30512 (N_30512,N_28926,N_29396);
xnor U30513 (N_30513,N_29611,N_28777);
xnor U30514 (N_30514,N_29080,N_29769);
nor U30515 (N_30515,N_28636,N_29102);
or U30516 (N_30516,N_28781,N_28571);
or U30517 (N_30517,N_29552,N_29768);
xor U30518 (N_30518,N_29848,N_29404);
or U30519 (N_30519,N_28789,N_29731);
or U30520 (N_30520,N_29542,N_29961);
nand U30521 (N_30521,N_29240,N_28836);
nor U30522 (N_30522,N_29009,N_29907);
nor U30523 (N_30523,N_29281,N_28155);
and U30524 (N_30524,N_29225,N_28567);
or U30525 (N_30525,N_29578,N_28124);
or U30526 (N_30526,N_29460,N_28369);
and U30527 (N_30527,N_28354,N_28990);
nor U30528 (N_30528,N_28888,N_28612);
nand U30529 (N_30529,N_28860,N_29818);
or U30530 (N_30530,N_29145,N_28670);
xor U30531 (N_30531,N_28963,N_29915);
nand U30532 (N_30532,N_28747,N_29943);
nor U30533 (N_30533,N_29574,N_29016);
xnor U30534 (N_30534,N_29581,N_29994);
or U30535 (N_30535,N_28746,N_28122);
nor U30536 (N_30536,N_28431,N_28187);
nand U30537 (N_30537,N_29263,N_29798);
nor U30538 (N_30538,N_29124,N_28001);
or U30539 (N_30539,N_28298,N_28331);
nor U30540 (N_30540,N_28042,N_29576);
and U30541 (N_30541,N_29438,N_29949);
nor U30542 (N_30542,N_29764,N_29037);
nor U30543 (N_30543,N_29530,N_28668);
nand U30544 (N_30544,N_29274,N_29212);
or U30545 (N_30545,N_28182,N_28435);
nand U30546 (N_30546,N_29082,N_28748);
nand U30547 (N_30547,N_29325,N_29287);
nand U30548 (N_30548,N_29666,N_28712);
xor U30549 (N_30549,N_29132,N_29594);
xor U30550 (N_30550,N_28577,N_29917);
and U30551 (N_30551,N_28651,N_28173);
xnor U30552 (N_30552,N_28032,N_28862);
xor U30553 (N_30553,N_28638,N_29055);
or U30554 (N_30554,N_29056,N_28319);
or U30555 (N_30555,N_29804,N_29550);
xor U30556 (N_30556,N_28919,N_29170);
xor U30557 (N_30557,N_28951,N_28716);
nor U30558 (N_30558,N_28596,N_28970);
xnor U30559 (N_30559,N_28696,N_29930);
and U30560 (N_30560,N_29722,N_28123);
nand U30561 (N_30561,N_28576,N_28681);
xnor U30562 (N_30562,N_28546,N_29385);
nor U30563 (N_30563,N_29790,N_29308);
or U30564 (N_30564,N_29882,N_28718);
xor U30565 (N_30565,N_29319,N_29701);
nor U30566 (N_30566,N_28520,N_28901);
or U30567 (N_30567,N_29012,N_28446);
nand U30568 (N_30568,N_28737,N_28559);
nand U30569 (N_30569,N_29491,N_29034);
and U30570 (N_30570,N_28344,N_29235);
nor U30571 (N_30571,N_28294,N_29500);
nand U30572 (N_30572,N_29395,N_28382);
nand U30573 (N_30573,N_28640,N_28898);
nor U30574 (N_30574,N_28850,N_28494);
or U30575 (N_30575,N_29078,N_28934);
xor U30576 (N_30576,N_29900,N_28621);
and U30577 (N_30577,N_29252,N_29737);
nor U30578 (N_30578,N_29320,N_29775);
and U30579 (N_30579,N_29336,N_28373);
xor U30580 (N_30580,N_29519,N_29663);
or U30581 (N_30581,N_29112,N_29793);
xnor U30582 (N_30582,N_28480,N_29929);
xor U30583 (N_30583,N_29355,N_28432);
nand U30584 (N_30584,N_28553,N_28051);
and U30585 (N_30585,N_29669,N_29073);
nand U30586 (N_30586,N_29264,N_28729);
nand U30587 (N_30587,N_29152,N_29538);
and U30588 (N_30588,N_29762,N_29427);
or U30589 (N_30589,N_29698,N_29615);
nor U30590 (N_30590,N_29499,N_29026);
or U30591 (N_30591,N_28797,N_29021);
and U30592 (N_30592,N_29753,N_29830);
nand U30593 (N_30593,N_29960,N_28938);
xor U30594 (N_30594,N_28469,N_28779);
nand U30595 (N_30595,N_28600,N_29282);
or U30596 (N_30596,N_29996,N_28805);
nand U30597 (N_30597,N_29032,N_29843);
xnor U30598 (N_30598,N_28762,N_29217);
and U30599 (N_30599,N_29452,N_28506);
nand U30600 (N_30600,N_29265,N_29076);
or U30601 (N_30601,N_28799,N_28316);
and U30602 (N_30602,N_29511,N_29118);
nor U30603 (N_30603,N_28601,N_28584);
nand U30604 (N_30604,N_29389,N_28859);
nand U30605 (N_30605,N_29305,N_28421);
nor U30606 (N_30606,N_28864,N_28239);
nor U30607 (N_30607,N_29417,N_29865);
and U30608 (N_30608,N_28701,N_28683);
xor U30609 (N_30609,N_28895,N_29904);
xor U30610 (N_30610,N_28914,N_29488);
or U30611 (N_30611,N_28108,N_29543);
xor U30612 (N_30612,N_28774,N_28166);
xor U30613 (N_30613,N_29837,N_28960);
nand U30614 (N_30614,N_28393,N_28362);
and U30615 (N_30615,N_29113,N_29272);
nand U30616 (N_30616,N_29751,N_28272);
or U30617 (N_30617,N_29014,N_28965);
nor U30618 (N_30618,N_29989,N_29380);
nand U30619 (N_30619,N_29894,N_28709);
and U30620 (N_30620,N_28834,N_29884);
nand U30621 (N_30621,N_28955,N_28704);
nor U30622 (N_30622,N_29001,N_29772);
xnor U30623 (N_30623,N_28389,N_28916);
and U30624 (N_30624,N_28940,N_28268);
and U30625 (N_30625,N_29261,N_29799);
or U30626 (N_30626,N_28873,N_28174);
nor U30627 (N_30627,N_29136,N_29997);
nand U30628 (N_30628,N_29600,N_28482);
xor U30629 (N_30629,N_28614,N_29134);
xor U30630 (N_30630,N_29365,N_29186);
nand U30631 (N_30631,N_29692,N_29708);
nor U30632 (N_30632,N_28613,N_28104);
nand U30633 (N_30633,N_28562,N_29029);
or U30634 (N_30634,N_28378,N_29369);
nand U30635 (N_30635,N_28463,N_28056);
xor U30636 (N_30636,N_28872,N_29192);
nand U30637 (N_30637,N_28003,N_29840);
or U30638 (N_30638,N_29291,N_29898);
or U30639 (N_30639,N_29779,N_28075);
or U30640 (N_30640,N_28014,N_28256);
nor U30641 (N_30641,N_28186,N_29850);
nor U30642 (N_30642,N_29442,N_29316);
nor U30643 (N_30643,N_28802,N_28870);
nand U30644 (N_30644,N_29138,N_28663);
nor U30645 (N_30645,N_29958,N_28568);
nor U30646 (N_30646,N_28374,N_28628);
nor U30647 (N_30647,N_29617,N_29310);
nand U30648 (N_30648,N_29750,N_29626);
nand U30649 (N_30649,N_29052,N_28889);
xor U30650 (N_30650,N_29173,N_28227);
nor U30651 (N_30651,N_28534,N_28391);
or U30652 (N_30652,N_28700,N_28942);
nand U30653 (N_30653,N_29304,N_29135);
or U30654 (N_30654,N_28489,N_29458);
nand U30655 (N_30655,N_28591,N_28739);
and U30656 (N_30656,N_29346,N_28679);
xor U30657 (N_30657,N_28711,N_28394);
xnor U30658 (N_30658,N_28165,N_28412);
xnor U30659 (N_30659,N_28565,N_28736);
nor U30660 (N_30660,N_29459,N_28409);
nand U30661 (N_30661,N_28705,N_28280);
or U30662 (N_30662,N_29902,N_28823);
nor U30663 (N_30663,N_29140,N_29471);
and U30664 (N_30664,N_28367,N_29010);
nand U30665 (N_30665,N_29237,N_29539);
nor U30666 (N_30666,N_29193,N_28118);
and U30667 (N_30667,N_28407,N_29993);
or U30668 (N_30668,N_29671,N_28829);
nand U30669 (N_30669,N_28130,N_28923);
xor U30670 (N_30670,N_28824,N_29783);
nand U30671 (N_30671,N_29486,N_28388);
nor U30672 (N_30672,N_28790,N_29372);
xor U30673 (N_30673,N_29150,N_28410);
and U30674 (N_30674,N_29732,N_29223);
xnor U30675 (N_30675,N_29812,N_28208);
and U30676 (N_30676,N_29300,N_29357);
or U30677 (N_30677,N_29221,N_28183);
and U30678 (N_30678,N_29070,N_28127);
xnor U30679 (N_30679,N_28055,N_29294);
nor U30680 (N_30680,N_28724,N_28976);
and U30681 (N_30681,N_28455,N_29483);
nand U30682 (N_30682,N_29968,N_29752);
and U30683 (N_30683,N_29353,N_29546);
nor U30684 (N_30684,N_29426,N_28727);
and U30685 (N_30685,N_28445,N_28931);
or U30686 (N_30686,N_28557,N_28010);
xor U30687 (N_30687,N_29912,N_29313);
xor U30688 (N_30688,N_28349,N_29407);
nand U30689 (N_30689,N_29167,N_28164);
nor U30690 (N_30690,N_29604,N_29646);
and U30691 (N_30691,N_28177,N_29362);
nor U30692 (N_30692,N_28804,N_28019);
nand U30693 (N_30693,N_28006,N_28029);
nor U30694 (N_30694,N_29918,N_28466);
and U30695 (N_30695,N_28624,N_29200);
nand U30696 (N_30696,N_29370,N_28502);
or U30697 (N_30697,N_28794,N_28784);
nand U30698 (N_30698,N_28000,N_28785);
or U30699 (N_30699,N_29035,N_28078);
nor U30700 (N_30700,N_29008,N_29189);
or U30701 (N_30701,N_28504,N_29168);
or U30702 (N_30702,N_29556,N_29063);
nand U30703 (N_30703,N_29868,N_29944);
nand U30704 (N_30704,N_29810,N_28760);
nor U30705 (N_30705,N_28035,N_29449);
xor U30706 (N_30706,N_28246,N_29979);
nand U30707 (N_30707,N_28215,N_28687);
xnor U30708 (N_30708,N_28320,N_29838);
nand U30709 (N_30709,N_28672,N_29603);
nor U30710 (N_30710,N_29307,N_29704);
xnor U30711 (N_30711,N_28111,N_28892);
xnor U30712 (N_30712,N_29540,N_29725);
or U30713 (N_30713,N_29204,N_28204);
xor U30714 (N_30714,N_29928,N_28767);
xnor U30715 (N_30715,N_29782,N_28630);
or U30716 (N_30716,N_29562,N_29444);
or U30717 (N_30717,N_29601,N_29828);
xor U30718 (N_30718,N_28887,N_29130);
nor U30719 (N_30719,N_28806,N_28340);
nor U30720 (N_30720,N_28526,N_29492);
and U30721 (N_30721,N_28971,N_28715);
xnor U30722 (N_30722,N_28699,N_29489);
or U30723 (N_30723,N_29649,N_28110);
xnor U30724 (N_30724,N_28740,N_28943);
or U30725 (N_30725,N_29673,N_28537);
or U30726 (N_30726,N_29967,N_29022);
nor U30727 (N_30727,N_28498,N_29624);
nor U30728 (N_30728,N_28311,N_28030);
nand U30729 (N_30729,N_29954,N_29572);
xor U30730 (N_30730,N_29208,N_29509);
xnor U30731 (N_30731,N_29122,N_29091);
nand U30732 (N_30732,N_29730,N_28112);
nand U30733 (N_30733,N_29593,N_29932);
nand U30734 (N_30734,N_28826,N_28043);
or U30735 (N_30735,N_28643,N_29157);
nand U30736 (N_30736,N_28588,N_28585);
nand U30737 (N_30737,N_29175,N_29020);
xnor U30738 (N_30738,N_29695,N_28813);
xor U30739 (N_30739,N_29101,N_29109);
xnor U30740 (N_30740,N_28939,N_28009);
nand U30741 (N_30741,N_29728,N_28743);
nor U30742 (N_30742,N_28555,N_29299);
nor U30743 (N_30743,N_29239,N_28810);
and U30744 (N_30744,N_28522,N_29482);
xnor U30745 (N_30745,N_29115,N_28485);
xor U30746 (N_30746,N_29098,N_29467);
and U30747 (N_30747,N_28151,N_29214);
and U30748 (N_30748,N_29432,N_29691);
nor U30749 (N_30749,N_29247,N_28991);
xor U30750 (N_30750,N_29019,N_28088);
and U30751 (N_30751,N_29723,N_29504);
or U30752 (N_30752,N_28569,N_29588);
nand U30753 (N_30753,N_29093,N_29318);
nand U30754 (N_30754,N_28202,N_28606);
nor U30755 (N_30755,N_29194,N_29454);
or U30756 (N_30756,N_29326,N_28024);
nand U30757 (N_30757,N_29802,N_28143);
or U30758 (N_30758,N_28935,N_29448);
nand U30759 (N_30759,N_28801,N_29181);
and U30760 (N_30760,N_28028,N_28282);
nand U30761 (N_30761,N_28808,N_28529);
nor U30762 (N_30762,N_28023,N_29043);
and U30763 (N_30763,N_29711,N_28928);
nor U30764 (N_30764,N_28822,N_28471);
or U30765 (N_30765,N_29651,N_29652);
nor U30766 (N_30766,N_28105,N_29059);
nand U30767 (N_30767,N_29216,N_28899);
or U30768 (N_30768,N_28634,N_28442);
nand U30769 (N_30769,N_28913,N_29919);
nand U30770 (N_30770,N_28220,N_28669);
nor U30771 (N_30771,N_28214,N_29408);
nor U30772 (N_30772,N_28125,N_29896);
or U30773 (N_30773,N_29777,N_28338);
xnor U30774 (N_30774,N_28156,N_28288);
or U30775 (N_30775,N_29209,N_29931);
or U30776 (N_30776,N_29558,N_29686);
and U30777 (N_30777,N_28266,N_28116);
nor U30778 (N_30778,N_28922,N_28383);
and U30779 (N_30779,N_28474,N_28918);
nand U30780 (N_30780,N_28259,N_28744);
nand U30781 (N_30781,N_29011,N_28408);
nor U30782 (N_30782,N_29231,N_28742);
nand U30783 (N_30783,N_29845,N_29834);
nand U30784 (N_30784,N_28749,N_28787);
nor U30785 (N_30785,N_29246,N_29048);
nand U30786 (N_30786,N_29890,N_29998);
nor U30787 (N_30787,N_28484,N_28831);
nor U30788 (N_30788,N_29616,N_28052);
nor U30789 (N_30789,N_28611,N_28418);
and U30790 (N_30790,N_28533,N_28552);
or U30791 (N_30791,N_28396,N_28945);
and U30792 (N_30792,N_29039,N_28501);
xor U30793 (N_30793,N_28304,N_29784);
nor U30794 (N_30794,N_28514,N_29475);
nand U30795 (N_30795,N_28074,N_29089);
nand U30796 (N_30796,N_29330,N_28191);
xnor U30797 (N_30797,N_29863,N_29903);
xor U30798 (N_30798,N_29363,N_28218);
and U30799 (N_30799,N_28241,N_29916);
xnor U30800 (N_30800,N_29520,N_28978);
and U30801 (N_30801,N_29266,N_29971);
and U30802 (N_30802,N_29635,N_29006);
nor U30803 (N_30803,N_28050,N_28539);
and U30804 (N_30804,N_29376,N_29559);
or U30805 (N_30805,N_28933,N_28825);
and U30806 (N_30806,N_29836,N_28967);
xor U30807 (N_30807,N_29630,N_29401);
xnor U30808 (N_30808,N_29236,N_29614);
nor U30809 (N_30809,N_28652,N_29859);
nand U30810 (N_30810,N_29557,N_29809);
and U30811 (N_30811,N_29797,N_29156);
or U30812 (N_30812,N_29017,N_29656);
xnor U30813 (N_30813,N_29441,N_29862);
and U30814 (N_30814,N_29920,N_29201);
nand U30815 (N_30815,N_29966,N_29062);
or U30816 (N_30816,N_28248,N_28317);
and U30817 (N_30817,N_29707,N_28755);
or U30818 (N_30818,N_28658,N_28861);
xnor U30819 (N_30819,N_28141,N_28351);
or U30820 (N_30820,N_29172,N_28674);
nor U30821 (N_30821,N_29197,N_29004);
nor U30822 (N_30822,N_29087,N_28661);
xnor U30823 (N_30823,N_28756,N_29411);
or U30824 (N_30824,N_29833,N_29638);
nand U30825 (N_30825,N_28549,N_28885);
and U30826 (N_30826,N_28275,N_29590);
or U30827 (N_30827,N_29125,N_28623);
nor U30828 (N_30828,N_28247,N_29211);
nand U30829 (N_30829,N_29083,N_28363);
xnor U30830 (N_30830,N_29096,N_29694);
xnor U30831 (N_30831,N_28093,N_28072);
nand U30832 (N_30832,N_28049,N_28903);
nor U30833 (N_30833,N_29286,N_29743);
xnor U30834 (N_30834,N_29437,N_29046);
or U30835 (N_30835,N_29554,N_28655);
nor U30836 (N_30836,N_29349,N_28071);
or U30837 (N_30837,N_28132,N_28906);
nand U30838 (N_30838,N_28095,N_28664);
or U30839 (N_30839,N_28896,N_29767);
and U30840 (N_30840,N_29964,N_29278);
or U30841 (N_30841,N_29678,N_28583);
and U30842 (N_30842,N_29981,N_29781);
nor U30843 (N_30843,N_29563,N_28206);
or U30844 (N_30844,N_28589,N_28503);
and U30845 (N_30845,N_28725,N_29255);
xor U30846 (N_30846,N_29251,N_28863);
or U30847 (N_30847,N_29297,N_29541);
nand U30848 (N_30848,N_28868,N_29390);
nor U30849 (N_30849,N_28563,N_28260);
nand U30850 (N_30850,N_29895,N_29412);
or U30851 (N_30851,N_28750,N_29555);
nand U30852 (N_30852,N_28018,N_28761);
and U30853 (N_30853,N_28312,N_28817);
or U30854 (N_30854,N_29064,N_28277);
or U30855 (N_30855,N_29924,N_29503);
or U30856 (N_30856,N_28076,N_28843);
and U30857 (N_30857,N_29275,N_29518);
nand U30858 (N_30858,N_28893,N_28053);
xor U30859 (N_30859,N_28464,N_28987);
nor U30860 (N_30860,N_28689,N_28253);
xor U30861 (N_30861,N_28039,N_29587);
xor U30862 (N_30862,N_29323,N_29814);
nor U30863 (N_30863,N_28149,N_29551);
xor U30864 (N_30864,N_28377,N_29533);
xor U30865 (N_30865,N_28190,N_29119);
nand U30866 (N_30866,N_29277,N_29841);
xnor U30867 (N_30867,N_29975,N_28134);
or U30868 (N_30868,N_28092,N_28244);
nand U30869 (N_30869,N_28720,N_29805);
or U30870 (N_30870,N_29342,N_29739);
nand U30871 (N_30871,N_28380,N_28483);
nor U30872 (N_30872,N_28622,N_28518);
nor U30873 (N_30873,N_29684,N_28488);
nand U30874 (N_30874,N_29028,N_29270);
or U30875 (N_30875,N_29787,N_29075);
or U30876 (N_30876,N_29569,N_28852);
xnor U30877 (N_30877,N_28188,N_29571);
nor U30878 (N_30878,N_28192,N_28129);
or U30879 (N_30879,N_29680,N_29665);
nor U30880 (N_30880,N_29284,N_28359);
xnor U30881 (N_30881,N_28213,N_28983);
or U30882 (N_30882,N_28738,N_29560);
and U30883 (N_30883,N_29154,N_28731);
and U30884 (N_30884,N_29613,N_28115);
or U30885 (N_30885,N_29521,N_29228);
or U30886 (N_30886,N_29873,N_29817);
and U30887 (N_30887,N_28982,N_29117);
xor U30888 (N_30888,N_29398,N_28384);
or U30889 (N_30889,N_29084,N_28327);
and U30890 (N_30890,N_28900,N_28871);
and U30891 (N_30891,N_29190,N_29586);
nand U30892 (N_30892,N_28309,N_29166);
nor U30893 (N_30893,N_29507,N_29510);
and U30894 (N_30894,N_28902,N_28201);
and U30895 (N_30895,N_29648,N_29180);
and U30896 (N_30896,N_29935,N_28511);
xor U30897 (N_30897,N_29285,N_28558);
nor U30898 (N_30898,N_29577,N_29434);
or U30899 (N_30899,N_28128,N_29451);
nor U30900 (N_30900,N_28245,N_29468);
or U30901 (N_30901,N_29632,N_28741);
and U30902 (N_30902,N_29527,N_28985);
nor U30903 (N_30903,N_29479,N_28144);
nand U30904 (N_30904,N_28303,N_29487);
and U30905 (N_30905,N_29185,N_28853);
nand U30906 (N_30906,N_28816,N_28233);
nand U30907 (N_30907,N_28428,N_29116);
and U30908 (N_30908,N_28113,N_28169);
nor U30909 (N_30909,N_28308,N_29716);
nor U30910 (N_30910,N_28941,N_29497);
nor U30911 (N_30911,N_28957,N_29844);
nor U30912 (N_30912,N_29870,N_28932);
or U30913 (N_30913,N_28572,N_29957);
nand U30914 (N_30914,N_28440,N_29233);
nor U30915 (N_30915,N_29374,N_29778);
xnor U30916 (N_30916,N_29956,N_29457);
nor U30917 (N_30917,N_29681,N_28194);
nand U30918 (N_30918,N_28536,N_29171);
and U30919 (N_30919,N_28176,N_29579);
nand U30920 (N_30920,N_29258,N_29425);
xnor U30921 (N_30921,N_28660,N_29983);
nand U30922 (N_30922,N_29653,N_29606);
nand U30923 (N_30923,N_28597,N_29191);
and U30924 (N_30924,N_28160,N_28659);
xor U30925 (N_30925,N_28343,N_28594);
or U30926 (N_30926,N_28375,N_29712);
and U30927 (N_30927,N_28673,N_28757);
xor U30928 (N_30928,N_28688,N_28336);
and U30929 (N_30929,N_29867,N_28513);
xnor U30930 (N_30930,N_28766,N_29478);
and U30931 (N_30931,N_29301,N_28299);
xor U30932 (N_30932,N_29811,N_28403);
and U30933 (N_30933,N_29120,N_29874);
xor U30934 (N_30934,N_28769,N_28593);
and U30935 (N_30935,N_28912,N_28193);
and U30936 (N_30936,N_28875,N_29331);
xnor U30937 (N_30937,N_29602,N_29259);
nand U30938 (N_30938,N_29531,N_28305);
and U30939 (N_30939,N_28457,N_28671);
nand U30940 (N_30940,N_29133,N_28581);
or U30941 (N_30941,N_29899,N_28313);
or U30942 (N_30942,N_28833,N_28274);
and U30943 (N_30943,N_28814,N_28619);
nor U30944 (N_30944,N_28602,N_28438);
or U30945 (N_30945,N_28152,N_28302);
xnor U30946 (N_30946,N_28395,N_29074);
nand U30947 (N_30947,N_28390,N_28953);
and U30948 (N_30948,N_29160,N_28775);
or U30949 (N_30949,N_29561,N_28424);
xor U30950 (N_30950,N_28335,N_28189);
xnor U30951 (N_30951,N_28948,N_29911);
and U30952 (N_30952,N_28838,N_29892);
and U30953 (N_30953,N_29761,N_28209);
xor U30954 (N_30954,N_28575,N_29697);
xnor U30955 (N_30955,N_28949,N_29808);
nand U30956 (N_30956,N_29823,N_29922);
or U30957 (N_30957,N_28353,N_29664);
xnor U30958 (N_30958,N_29030,N_29612);
or U30959 (N_30959,N_29469,N_28694);
xnor U30960 (N_30960,N_28927,N_29710);
nand U30961 (N_30961,N_28837,N_28433);
xor U30962 (N_30962,N_28080,N_28996);
and U30963 (N_30963,N_28224,N_28956);
or U30964 (N_30964,N_28452,N_29344);
and U30965 (N_30965,N_29402,N_29969);
and U30966 (N_30966,N_29582,N_29368);
or U30967 (N_30967,N_28975,N_29866);
xor U30968 (N_30968,N_28763,N_28465);
or U30969 (N_30969,N_29675,N_28877);
nor U30970 (N_30970,N_28682,N_29443);
or U30971 (N_30971,N_29354,N_28548);
nor U30972 (N_30972,N_29717,N_28300);
nor U30973 (N_30973,N_28507,N_29939);
nor U30974 (N_30974,N_29822,N_29791);
and U30975 (N_30975,N_29763,N_28402);
nor U30976 (N_30976,N_29025,N_29950);
xnor U30977 (N_30977,N_29934,N_28217);
nand U30978 (N_30978,N_29188,N_29031);
xnor U30979 (N_30979,N_29661,N_28812);
nor U30980 (N_30980,N_28037,N_28085);
nor U30981 (N_30981,N_28271,N_28969);
and U30982 (N_30982,N_29676,N_29024);
or U30983 (N_30983,N_28603,N_28815);
or U30984 (N_30984,N_28267,N_29580);
xor U30985 (N_30985,N_29720,N_28920);
or U30986 (N_30986,N_28570,N_28162);
and U30987 (N_30987,N_29999,N_28776);
nor U30988 (N_30988,N_29058,N_28807);
xnor U30989 (N_30989,N_28073,N_29111);
nor U30990 (N_30990,N_29976,N_28692);
nor U30991 (N_30991,N_29909,N_28416);
nor U30992 (N_30992,N_29970,N_28135);
nor U30993 (N_30993,N_29738,N_28792);
xnor U30994 (N_30994,N_29205,N_29359);
nor U30995 (N_30995,N_29962,N_28908);
nand U30996 (N_30996,N_29610,N_29224);
or U30997 (N_30997,N_28984,N_29254);
xnor U30998 (N_30998,N_28793,N_28443);
nand U30999 (N_30999,N_28083,N_29523);
nand U31000 (N_31000,N_28484,N_29660);
xnor U31001 (N_31001,N_29466,N_28494);
nor U31002 (N_31002,N_29963,N_29109);
nor U31003 (N_31003,N_29390,N_28024);
or U31004 (N_31004,N_28405,N_29698);
and U31005 (N_31005,N_29047,N_28348);
nand U31006 (N_31006,N_28953,N_28244);
and U31007 (N_31007,N_28230,N_29194);
or U31008 (N_31008,N_29895,N_29770);
xor U31009 (N_31009,N_29238,N_28898);
or U31010 (N_31010,N_29311,N_29622);
nor U31011 (N_31011,N_28142,N_28798);
or U31012 (N_31012,N_29365,N_29071);
nand U31013 (N_31013,N_28756,N_29725);
or U31014 (N_31014,N_29211,N_28142);
nand U31015 (N_31015,N_28426,N_28155);
or U31016 (N_31016,N_28738,N_29703);
xor U31017 (N_31017,N_29981,N_28569);
or U31018 (N_31018,N_29489,N_28721);
or U31019 (N_31019,N_28397,N_29660);
xor U31020 (N_31020,N_28563,N_28550);
xnor U31021 (N_31021,N_28526,N_28962);
nand U31022 (N_31022,N_28696,N_28876);
or U31023 (N_31023,N_28507,N_29270);
or U31024 (N_31024,N_28585,N_28150);
or U31025 (N_31025,N_29949,N_29425);
xor U31026 (N_31026,N_29043,N_29823);
or U31027 (N_31027,N_29066,N_28855);
and U31028 (N_31028,N_29161,N_28575);
xor U31029 (N_31029,N_29039,N_29558);
or U31030 (N_31030,N_29140,N_28294);
nand U31031 (N_31031,N_29454,N_29735);
nand U31032 (N_31032,N_28098,N_28006);
xor U31033 (N_31033,N_29721,N_28978);
nand U31034 (N_31034,N_28248,N_29516);
nor U31035 (N_31035,N_28473,N_29459);
xnor U31036 (N_31036,N_28271,N_28485);
nor U31037 (N_31037,N_29498,N_29962);
and U31038 (N_31038,N_29158,N_28467);
and U31039 (N_31039,N_28000,N_29638);
nor U31040 (N_31040,N_29913,N_29936);
or U31041 (N_31041,N_28571,N_29608);
nor U31042 (N_31042,N_29293,N_28440);
or U31043 (N_31043,N_29655,N_28235);
or U31044 (N_31044,N_29378,N_28898);
nor U31045 (N_31045,N_29114,N_28923);
xor U31046 (N_31046,N_29326,N_28417);
and U31047 (N_31047,N_28658,N_28002);
nand U31048 (N_31048,N_28212,N_29238);
nor U31049 (N_31049,N_29202,N_28349);
nor U31050 (N_31050,N_29269,N_28307);
nand U31051 (N_31051,N_29852,N_28608);
or U31052 (N_31052,N_29404,N_29264);
and U31053 (N_31053,N_29943,N_29858);
xor U31054 (N_31054,N_29129,N_28409);
xor U31055 (N_31055,N_28792,N_28341);
or U31056 (N_31056,N_29753,N_28997);
or U31057 (N_31057,N_28284,N_29809);
and U31058 (N_31058,N_29465,N_28591);
xnor U31059 (N_31059,N_28257,N_28248);
nand U31060 (N_31060,N_28749,N_28969);
or U31061 (N_31061,N_29311,N_28939);
or U31062 (N_31062,N_29697,N_28437);
nand U31063 (N_31063,N_29956,N_29969);
xor U31064 (N_31064,N_29512,N_28177);
nand U31065 (N_31065,N_29904,N_28985);
nand U31066 (N_31066,N_28067,N_28436);
and U31067 (N_31067,N_29395,N_29358);
and U31068 (N_31068,N_29603,N_29192);
nand U31069 (N_31069,N_29402,N_28024);
xnor U31070 (N_31070,N_28439,N_29638);
nor U31071 (N_31071,N_28990,N_28576);
nor U31072 (N_31072,N_29131,N_29068);
nor U31073 (N_31073,N_28744,N_28757);
nor U31074 (N_31074,N_28249,N_28443);
nand U31075 (N_31075,N_29302,N_29583);
nor U31076 (N_31076,N_29525,N_28849);
nor U31077 (N_31077,N_29406,N_29209);
xor U31078 (N_31078,N_29816,N_29003);
nand U31079 (N_31079,N_29633,N_28307);
xnor U31080 (N_31080,N_29694,N_28009);
and U31081 (N_31081,N_28164,N_28561);
nor U31082 (N_31082,N_28821,N_29910);
xor U31083 (N_31083,N_29668,N_29148);
and U31084 (N_31084,N_28721,N_29260);
nand U31085 (N_31085,N_29552,N_28444);
or U31086 (N_31086,N_28194,N_28694);
or U31087 (N_31087,N_29416,N_29940);
nor U31088 (N_31088,N_29870,N_28778);
nor U31089 (N_31089,N_29162,N_29114);
nand U31090 (N_31090,N_28045,N_28762);
nor U31091 (N_31091,N_28015,N_28683);
and U31092 (N_31092,N_28809,N_28184);
and U31093 (N_31093,N_29164,N_28023);
xor U31094 (N_31094,N_28148,N_28479);
and U31095 (N_31095,N_29152,N_29684);
nand U31096 (N_31096,N_29440,N_28844);
nor U31097 (N_31097,N_29669,N_29385);
and U31098 (N_31098,N_29145,N_29226);
xor U31099 (N_31099,N_28031,N_28134);
xnor U31100 (N_31100,N_28926,N_28226);
and U31101 (N_31101,N_29773,N_28493);
nand U31102 (N_31102,N_28140,N_28669);
or U31103 (N_31103,N_29967,N_29755);
nand U31104 (N_31104,N_28501,N_29928);
or U31105 (N_31105,N_29238,N_28595);
nor U31106 (N_31106,N_29697,N_29942);
nand U31107 (N_31107,N_28114,N_28482);
nand U31108 (N_31108,N_28355,N_29682);
xnor U31109 (N_31109,N_28188,N_29454);
and U31110 (N_31110,N_28866,N_29916);
and U31111 (N_31111,N_28744,N_28443);
nor U31112 (N_31112,N_29531,N_29109);
and U31113 (N_31113,N_28126,N_28017);
nor U31114 (N_31114,N_28703,N_28817);
or U31115 (N_31115,N_29128,N_29072);
or U31116 (N_31116,N_28452,N_29247);
and U31117 (N_31117,N_28228,N_29425);
xor U31118 (N_31118,N_28696,N_29379);
nor U31119 (N_31119,N_29756,N_28983);
xnor U31120 (N_31120,N_29797,N_29775);
nor U31121 (N_31121,N_28575,N_28089);
or U31122 (N_31122,N_28220,N_29192);
nor U31123 (N_31123,N_28319,N_29373);
nor U31124 (N_31124,N_28251,N_29770);
or U31125 (N_31125,N_28851,N_29753);
nor U31126 (N_31126,N_28536,N_29480);
nand U31127 (N_31127,N_29101,N_29322);
xor U31128 (N_31128,N_29484,N_29206);
or U31129 (N_31129,N_28259,N_29215);
nor U31130 (N_31130,N_28290,N_29543);
and U31131 (N_31131,N_28052,N_28904);
and U31132 (N_31132,N_28050,N_28077);
xor U31133 (N_31133,N_29061,N_29705);
nand U31134 (N_31134,N_28828,N_29533);
nor U31135 (N_31135,N_28174,N_29461);
and U31136 (N_31136,N_29709,N_28472);
xor U31137 (N_31137,N_29750,N_29346);
and U31138 (N_31138,N_28843,N_29173);
or U31139 (N_31139,N_29179,N_28202);
nor U31140 (N_31140,N_29127,N_29928);
nand U31141 (N_31141,N_29057,N_28127);
nor U31142 (N_31142,N_29634,N_29338);
or U31143 (N_31143,N_29126,N_28399);
nor U31144 (N_31144,N_29339,N_29774);
or U31145 (N_31145,N_28189,N_28186);
nor U31146 (N_31146,N_28558,N_28978);
nor U31147 (N_31147,N_28078,N_29613);
nand U31148 (N_31148,N_29512,N_29816);
nand U31149 (N_31149,N_28692,N_29145);
nor U31150 (N_31150,N_28736,N_28913);
nor U31151 (N_31151,N_29668,N_29750);
or U31152 (N_31152,N_28369,N_28110);
or U31153 (N_31153,N_29775,N_29052);
nor U31154 (N_31154,N_29415,N_29611);
xor U31155 (N_31155,N_28102,N_28387);
or U31156 (N_31156,N_28839,N_28782);
nand U31157 (N_31157,N_28363,N_28328);
and U31158 (N_31158,N_28603,N_29375);
or U31159 (N_31159,N_28177,N_29386);
or U31160 (N_31160,N_28310,N_29447);
or U31161 (N_31161,N_28440,N_29888);
nand U31162 (N_31162,N_29062,N_29434);
nand U31163 (N_31163,N_29923,N_29070);
xor U31164 (N_31164,N_29415,N_28990);
nand U31165 (N_31165,N_29067,N_29312);
nand U31166 (N_31166,N_29480,N_28355);
xnor U31167 (N_31167,N_29334,N_28758);
xnor U31168 (N_31168,N_29692,N_28052);
and U31169 (N_31169,N_29834,N_29003);
and U31170 (N_31170,N_29479,N_28914);
nand U31171 (N_31171,N_28002,N_29357);
and U31172 (N_31172,N_29050,N_28390);
nand U31173 (N_31173,N_29390,N_28716);
nor U31174 (N_31174,N_29822,N_28110);
and U31175 (N_31175,N_29209,N_28633);
or U31176 (N_31176,N_28462,N_29076);
nand U31177 (N_31177,N_29268,N_29156);
or U31178 (N_31178,N_28884,N_29538);
nor U31179 (N_31179,N_29782,N_29638);
xor U31180 (N_31180,N_29102,N_28141);
and U31181 (N_31181,N_29534,N_29144);
xnor U31182 (N_31182,N_29692,N_29223);
or U31183 (N_31183,N_28150,N_28036);
xnor U31184 (N_31184,N_29407,N_29733);
or U31185 (N_31185,N_29149,N_28794);
or U31186 (N_31186,N_29601,N_28503);
or U31187 (N_31187,N_28289,N_29783);
nand U31188 (N_31188,N_28290,N_29209);
nor U31189 (N_31189,N_29330,N_29847);
xnor U31190 (N_31190,N_28400,N_29063);
or U31191 (N_31191,N_28431,N_29047);
or U31192 (N_31192,N_28268,N_28160);
nor U31193 (N_31193,N_28058,N_29335);
and U31194 (N_31194,N_28340,N_29631);
or U31195 (N_31195,N_28888,N_29715);
and U31196 (N_31196,N_28527,N_28977);
or U31197 (N_31197,N_28385,N_28827);
xor U31198 (N_31198,N_28309,N_28965);
and U31199 (N_31199,N_28529,N_29434);
or U31200 (N_31200,N_28988,N_28999);
and U31201 (N_31201,N_28834,N_29687);
and U31202 (N_31202,N_28499,N_29337);
and U31203 (N_31203,N_28465,N_28004);
or U31204 (N_31204,N_29115,N_28908);
xor U31205 (N_31205,N_28190,N_28900);
and U31206 (N_31206,N_29639,N_29501);
nor U31207 (N_31207,N_29254,N_29856);
and U31208 (N_31208,N_28970,N_28290);
xor U31209 (N_31209,N_29258,N_29005);
or U31210 (N_31210,N_28898,N_29702);
and U31211 (N_31211,N_29506,N_28454);
nand U31212 (N_31212,N_28170,N_29801);
nand U31213 (N_31213,N_29224,N_29812);
nor U31214 (N_31214,N_29784,N_28881);
and U31215 (N_31215,N_28322,N_29739);
xnor U31216 (N_31216,N_28181,N_29446);
nor U31217 (N_31217,N_28473,N_28745);
and U31218 (N_31218,N_28814,N_29087);
nor U31219 (N_31219,N_29689,N_28607);
or U31220 (N_31220,N_29923,N_28217);
nor U31221 (N_31221,N_29084,N_29536);
nor U31222 (N_31222,N_28836,N_28940);
nand U31223 (N_31223,N_29038,N_28359);
and U31224 (N_31224,N_28970,N_28286);
and U31225 (N_31225,N_28105,N_29719);
nor U31226 (N_31226,N_29561,N_29643);
nor U31227 (N_31227,N_28952,N_28454);
nor U31228 (N_31228,N_28675,N_29613);
nor U31229 (N_31229,N_29393,N_28944);
xor U31230 (N_31230,N_28081,N_28134);
or U31231 (N_31231,N_28577,N_28647);
nand U31232 (N_31232,N_28629,N_29298);
nor U31233 (N_31233,N_28862,N_29358);
xor U31234 (N_31234,N_28738,N_28808);
and U31235 (N_31235,N_28769,N_28574);
nand U31236 (N_31236,N_28077,N_29743);
and U31237 (N_31237,N_28358,N_28795);
and U31238 (N_31238,N_28528,N_29288);
or U31239 (N_31239,N_29037,N_28218);
nor U31240 (N_31240,N_29303,N_29389);
and U31241 (N_31241,N_28182,N_29178);
or U31242 (N_31242,N_28639,N_29161);
nor U31243 (N_31243,N_28429,N_29310);
and U31244 (N_31244,N_28920,N_28446);
or U31245 (N_31245,N_29217,N_28283);
nand U31246 (N_31246,N_28260,N_29361);
nand U31247 (N_31247,N_29005,N_29514);
nor U31248 (N_31248,N_28720,N_28517);
xnor U31249 (N_31249,N_28841,N_28182);
or U31250 (N_31250,N_29516,N_28039);
nor U31251 (N_31251,N_28880,N_29628);
xor U31252 (N_31252,N_29981,N_28313);
and U31253 (N_31253,N_29881,N_28008);
xor U31254 (N_31254,N_28451,N_29499);
or U31255 (N_31255,N_29986,N_28304);
or U31256 (N_31256,N_29816,N_29281);
xnor U31257 (N_31257,N_29792,N_29869);
nand U31258 (N_31258,N_28487,N_29102);
or U31259 (N_31259,N_29347,N_29836);
nand U31260 (N_31260,N_28379,N_28482);
and U31261 (N_31261,N_29427,N_29275);
xnor U31262 (N_31262,N_28171,N_29136);
nor U31263 (N_31263,N_29452,N_28836);
nand U31264 (N_31264,N_29920,N_29134);
or U31265 (N_31265,N_28235,N_29405);
xnor U31266 (N_31266,N_28686,N_29849);
and U31267 (N_31267,N_29352,N_29357);
nand U31268 (N_31268,N_28721,N_28825);
and U31269 (N_31269,N_28376,N_28254);
nand U31270 (N_31270,N_29392,N_28241);
and U31271 (N_31271,N_29184,N_29668);
nor U31272 (N_31272,N_29897,N_28033);
xor U31273 (N_31273,N_28144,N_28003);
xor U31274 (N_31274,N_28281,N_29858);
nor U31275 (N_31275,N_29200,N_28541);
nand U31276 (N_31276,N_28626,N_29916);
and U31277 (N_31277,N_29596,N_29424);
and U31278 (N_31278,N_28403,N_28447);
nor U31279 (N_31279,N_29177,N_29724);
nor U31280 (N_31280,N_29167,N_28413);
or U31281 (N_31281,N_29079,N_29243);
xnor U31282 (N_31282,N_28456,N_28045);
xnor U31283 (N_31283,N_28657,N_29247);
or U31284 (N_31284,N_29594,N_29472);
xor U31285 (N_31285,N_28362,N_28834);
and U31286 (N_31286,N_29292,N_29684);
or U31287 (N_31287,N_29700,N_28925);
xnor U31288 (N_31288,N_29109,N_28543);
nand U31289 (N_31289,N_29372,N_29671);
xnor U31290 (N_31290,N_29013,N_29904);
xor U31291 (N_31291,N_29578,N_29327);
xnor U31292 (N_31292,N_29212,N_28164);
nor U31293 (N_31293,N_28126,N_28550);
and U31294 (N_31294,N_28780,N_29882);
nand U31295 (N_31295,N_29067,N_29545);
nor U31296 (N_31296,N_28759,N_29786);
nand U31297 (N_31297,N_29533,N_28057);
and U31298 (N_31298,N_28395,N_29459);
and U31299 (N_31299,N_28515,N_29822);
nand U31300 (N_31300,N_28102,N_29487);
nand U31301 (N_31301,N_28746,N_28629);
nand U31302 (N_31302,N_29085,N_29880);
and U31303 (N_31303,N_29340,N_28081);
or U31304 (N_31304,N_29179,N_29881);
xor U31305 (N_31305,N_29925,N_29300);
and U31306 (N_31306,N_28787,N_28698);
nor U31307 (N_31307,N_29064,N_28741);
or U31308 (N_31308,N_28414,N_29846);
nand U31309 (N_31309,N_28648,N_29654);
or U31310 (N_31310,N_28764,N_29783);
nor U31311 (N_31311,N_28795,N_28813);
nand U31312 (N_31312,N_29303,N_29464);
and U31313 (N_31313,N_29547,N_28296);
xor U31314 (N_31314,N_28559,N_28996);
xor U31315 (N_31315,N_29763,N_28838);
xnor U31316 (N_31316,N_28273,N_28240);
or U31317 (N_31317,N_29998,N_28419);
nor U31318 (N_31318,N_29198,N_29763);
or U31319 (N_31319,N_29380,N_29174);
xnor U31320 (N_31320,N_28769,N_29860);
xor U31321 (N_31321,N_28303,N_29390);
nor U31322 (N_31322,N_28230,N_29969);
or U31323 (N_31323,N_28714,N_28882);
nor U31324 (N_31324,N_29122,N_28774);
xnor U31325 (N_31325,N_28072,N_28930);
nand U31326 (N_31326,N_29007,N_29819);
nand U31327 (N_31327,N_29472,N_29138);
nor U31328 (N_31328,N_28183,N_29998);
nor U31329 (N_31329,N_28365,N_28152);
or U31330 (N_31330,N_29169,N_28535);
xor U31331 (N_31331,N_28665,N_28204);
xnor U31332 (N_31332,N_29389,N_28795);
and U31333 (N_31333,N_29597,N_29465);
nor U31334 (N_31334,N_28270,N_29708);
nand U31335 (N_31335,N_29046,N_28525);
or U31336 (N_31336,N_28359,N_29704);
or U31337 (N_31337,N_28654,N_28450);
xor U31338 (N_31338,N_28276,N_28051);
and U31339 (N_31339,N_28279,N_28648);
or U31340 (N_31340,N_29751,N_29165);
and U31341 (N_31341,N_29856,N_28806);
xnor U31342 (N_31342,N_29096,N_28529);
nor U31343 (N_31343,N_29362,N_28692);
or U31344 (N_31344,N_28277,N_29725);
or U31345 (N_31345,N_29813,N_29051);
or U31346 (N_31346,N_28057,N_29673);
and U31347 (N_31347,N_29689,N_29771);
or U31348 (N_31348,N_28340,N_28987);
or U31349 (N_31349,N_29634,N_28053);
xor U31350 (N_31350,N_29349,N_29867);
or U31351 (N_31351,N_28121,N_29920);
nand U31352 (N_31352,N_28779,N_28685);
nor U31353 (N_31353,N_29887,N_29473);
nand U31354 (N_31354,N_29704,N_28186);
nand U31355 (N_31355,N_28727,N_29448);
and U31356 (N_31356,N_28397,N_29914);
nor U31357 (N_31357,N_29615,N_29328);
xnor U31358 (N_31358,N_29637,N_29858);
nor U31359 (N_31359,N_29547,N_28074);
xor U31360 (N_31360,N_28904,N_28076);
nand U31361 (N_31361,N_29471,N_29485);
or U31362 (N_31362,N_29253,N_28697);
and U31363 (N_31363,N_29200,N_28360);
nand U31364 (N_31364,N_28187,N_29104);
or U31365 (N_31365,N_29336,N_28723);
xnor U31366 (N_31366,N_28398,N_28721);
nor U31367 (N_31367,N_29916,N_28323);
xor U31368 (N_31368,N_29136,N_29226);
nand U31369 (N_31369,N_29999,N_29672);
xnor U31370 (N_31370,N_29303,N_28615);
or U31371 (N_31371,N_28835,N_28544);
xor U31372 (N_31372,N_28475,N_29746);
nor U31373 (N_31373,N_28846,N_29354);
and U31374 (N_31374,N_28433,N_29197);
nor U31375 (N_31375,N_29061,N_28726);
and U31376 (N_31376,N_29407,N_28783);
nand U31377 (N_31377,N_28069,N_29843);
and U31378 (N_31378,N_28048,N_28227);
or U31379 (N_31379,N_28412,N_29030);
xor U31380 (N_31380,N_28719,N_28062);
and U31381 (N_31381,N_28061,N_29780);
xnor U31382 (N_31382,N_29905,N_29342);
nand U31383 (N_31383,N_28818,N_28554);
xor U31384 (N_31384,N_28167,N_29668);
nand U31385 (N_31385,N_29164,N_28900);
nand U31386 (N_31386,N_28852,N_28045);
xnor U31387 (N_31387,N_29045,N_29609);
xor U31388 (N_31388,N_29829,N_28618);
or U31389 (N_31389,N_29731,N_28937);
xor U31390 (N_31390,N_28388,N_28987);
xnor U31391 (N_31391,N_28182,N_29770);
and U31392 (N_31392,N_29126,N_29760);
nand U31393 (N_31393,N_28362,N_29692);
or U31394 (N_31394,N_28134,N_28242);
xor U31395 (N_31395,N_28748,N_29607);
xnor U31396 (N_31396,N_28711,N_29633);
nand U31397 (N_31397,N_29847,N_29664);
nor U31398 (N_31398,N_29781,N_29771);
nand U31399 (N_31399,N_28147,N_29755);
or U31400 (N_31400,N_28651,N_29305);
or U31401 (N_31401,N_28507,N_28462);
and U31402 (N_31402,N_28588,N_29776);
nand U31403 (N_31403,N_29819,N_28356);
nand U31404 (N_31404,N_29285,N_28874);
or U31405 (N_31405,N_29559,N_29314);
xor U31406 (N_31406,N_28334,N_29726);
and U31407 (N_31407,N_29231,N_29902);
and U31408 (N_31408,N_29329,N_28608);
nand U31409 (N_31409,N_29693,N_28001);
xor U31410 (N_31410,N_29259,N_29513);
nor U31411 (N_31411,N_28687,N_28775);
nand U31412 (N_31412,N_29580,N_29244);
and U31413 (N_31413,N_29114,N_28930);
nand U31414 (N_31414,N_29289,N_29804);
nor U31415 (N_31415,N_29088,N_28008);
xnor U31416 (N_31416,N_29726,N_29368);
nor U31417 (N_31417,N_28408,N_28943);
or U31418 (N_31418,N_29135,N_28956);
nor U31419 (N_31419,N_29708,N_29338);
nand U31420 (N_31420,N_29377,N_28330);
xnor U31421 (N_31421,N_28678,N_29020);
or U31422 (N_31422,N_28771,N_29023);
nor U31423 (N_31423,N_29768,N_28856);
xor U31424 (N_31424,N_28650,N_29232);
and U31425 (N_31425,N_28284,N_29671);
or U31426 (N_31426,N_28360,N_29864);
and U31427 (N_31427,N_28886,N_28559);
and U31428 (N_31428,N_29695,N_28431);
nor U31429 (N_31429,N_28933,N_28202);
nand U31430 (N_31430,N_28607,N_29843);
xnor U31431 (N_31431,N_29300,N_28675);
nor U31432 (N_31432,N_28281,N_29939);
xnor U31433 (N_31433,N_28016,N_29896);
or U31434 (N_31434,N_29477,N_29282);
xnor U31435 (N_31435,N_28192,N_28896);
nand U31436 (N_31436,N_29416,N_28789);
xnor U31437 (N_31437,N_28753,N_29240);
nor U31438 (N_31438,N_29504,N_29462);
or U31439 (N_31439,N_29861,N_28711);
or U31440 (N_31440,N_28628,N_29758);
nor U31441 (N_31441,N_28644,N_28144);
and U31442 (N_31442,N_29833,N_29734);
xor U31443 (N_31443,N_28735,N_29775);
nor U31444 (N_31444,N_29213,N_28224);
and U31445 (N_31445,N_28232,N_29701);
nor U31446 (N_31446,N_28907,N_29479);
nor U31447 (N_31447,N_28898,N_28371);
xnor U31448 (N_31448,N_28383,N_28612);
or U31449 (N_31449,N_29387,N_29245);
nor U31450 (N_31450,N_29564,N_29209);
nand U31451 (N_31451,N_28972,N_28613);
or U31452 (N_31452,N_29249,N_28041);
and U31453 (N_31453,N_29888,N_28465);
nor U31454 (N_31454,N_29860,N_28012);
or U31455 (N_31455,N_28009,N_28193);
nor U31456 (N_31456,N_29921,N_29029);
nand U31457 (N_31457,N_29708,N_29399);
and U31458 (N_31458,N_28253,N_28406);
and U31459 (N_31459,N_28054,N_29009);
and U31460 (N_31460,N_28497,N_28502);
nand U31461 (N_31461,N_29207,N_29904);
and U31462 (N_31462,N_28943,N_28554);
nor U31463 (N_31463,N_29750,N_28398);
and U31464 (N_31464,N_29420,N_29779);
and U31465 (N_31465,N_28363,N_29869);
xor U31466 (N_31466,N_28217,N_29815);
xnor U31467 (N_31467,N_29194,N_29909);
and U31468 (N_31468,N_28355,N_28420);
xor U31469 (N_31469,N_29244,N_28619);
xor U31470 (N_31470,N_29132,N_28306);
xor U31471 (N_31471,N_29817,N_29527);
or U31472 (N_31472,N_29388,N_29439);
and U31473 (N_31473,N_29117,N_29321);
nand U31474 (N_31474,N_28298,N_29166);
and U31475 (N_31475,N_29079,N_28056);
xnor U31476 (N_31476,N_29187,N_28984);
nand U31477 (N_31477,N_28864,N_29104);
nand U31478 (N_31478,N_29822,N_29212);
nor U31479 (N_31479,N_29546,N_28459);
and U31480 (N_31480,N_29838,N_28814);
nor U31481 (N_31481,N_29270,N_28897);
nand U31482 (N_31482,N_28596,N_28972);
xor U31483 (N_31483,N_28391,N_28036);
nor U31484 (N_31484,N_28482,N_29910);
and U31485 (N_31485,N_28953,N_28769);
nor U31486 (N_31486,N_29686,N_28785);
or U31487 (N_31487,N_28304,N_28062);
nor U31488 (N_31488,N_29789,N_29573);
xor U31489 (N_31489,N_29422,N_29639);
nand U31490 (N_31490,N_29680,N_29146);
and U31491 (N_31491,N_28259,N_29012);
nor U31492 (N_31492,N_29547,N_29099);
xnor U31493 (N_31493,N_29224,N_28163);
nand U31494 (N_31494,N_28844,N_29778);
nor U31495 (N_31495,N_29201,N_28629);
xor U31496 (N_31496,N_29819,N_28752);
xor U31497 (N_31497,N_29952,N_28142);
xor U31498 (N_31498,N_28036,N_29264);
nor U31499 (N_31499,N_28595,N_29086);
nor U31500 (N_31500,N_28580,N_28653);
nand U31501 (N_31501,N_28238,N_29090);
and U31502 (N_31502,N_28183,N_29105);
and U31503 (N_31503,N_29912,N_29873);
nand U31504 (N_31504,N_29250,N_29202);
nand U31505 (N_31505,N_29946,N_29770);
nor U31506 (N_31506,N_28020,N_28893);
nor U31507 (N_31507,N_28212,N_28573);
or U31508 (N_31508,N_28452,N_29627);
nor U31509 (N_31509,N_28766,N_29635);
nand U31510 (N_31510,N_28950,N_28712);
nand U31511 (N_31511,N_28937,N_28930);
and U31512 (N_31512,N_29521,N_28105);
nand U31513 (N_31513,N_28589,N_28942);
and U31514 (N_31514,N_28056,N_29487);
and U31515 (N_31515,N_29913,N_29843);
nand U31516 (N_31516,N_28463,N_29290);
xor U31517 (N_31517,N_28062,N_28308);
xor U31518 (N_31518,N_29625,N_29353);
xor U31519 (N_31519,N_28788,N_28860);
nand U31520 (N_31520,N_29759,N_28092);
nand U31521 (N_31521,N_28098,N_29970);
xor U31522 (N_31522,N_28557,N_29520);
and U31523 (N_31523,N_28517,N_29944);
and U31524 (N_31524,N_29474,N_28647);
nand U31525 (N_31525,N_28691,N_28186);
or U31526 (N_31526,N_29704,N_29232);
nor U31527 (N_31527,N_28647,N_29094);
nor U31528 (N_31528,N_28867,N_28581);
nor U31529 (N_31529,N_28869,N_29801);
and U31530 (N_31530,N_28678,N_29794);
nor U31531 (N_31531,N_29068,N_29635);
xor U31532 (N_31532,N_29128,N_28373);
nor U31533 (N_31533,N_28385,N_29378);
xor U31534 (N_31534,N_29617,N_28500);
nand U31535 (N_31535,N_29593,N_28231);
nand U31536 (N_31536,N_28170,N_28670);
and U31537 (N_31537,N_28134,N_28877);
or U31538 (N_31538,N_28475,N_29257);
or U31539 (N_31539,N_28749,N_29679);
and U31540 (N_31540,N_28301,N_29481);
nor U31541 (N_31541,N_29909,N_28730);
or U31542 (N_31542,N_29215,N_28936);
or U31543 (N_31543,N_28525,N_29727);
xor U31544 (N_31544,N_29927,N_29273);
or U31545 (N_31545,N_28675,N_29698);
and U31546 (N_31546,N_29112,N_29877);
and U31547 (N_31547,N_29039,N_28933);
xor U31548 (N_31548,N_28208,N_28848);
xnor U31549 (N_31549,N_28890,N_29787);
nand U31550 (N_31550,N_29567,N_29101);
and U31551 (N_31551,N_28674,N_28477);
or U31552 (N_31552,N_29574,N_28434);
nand U31553 (N_31553,N_28691,N_29940);
and U31554 (N_31554,N_28586,N_29699);
nor U31555 (N_31555,N_29715,N_28878);
nand U31556 (N_31556,N_28649,N_28157);
or U31557 (N_31557,N_29812,N_28739);
xnor U31558 (N_31558,N_28471,N_28484);
xnor U31559 (N_31559,N_28474,N_29724);
or U31560 (N_31560,N_29017,N_28518);
nand U31561 (N_31561,N_29197,N_29880);
and U31562 (N_31562,N_28816,N_28527);
nand U31563 (N_31563,N_29204,N_28795);
and U31564 (N_31564,N_29995,N_28309);
or U31565 (N_31565,N_29707,N_28870);
or U31566 (N_31566,N_28971,N_28171);
or U31567 (N_31567,N_28811,N_28587);
and U31568 (N_31568,N_29668,N_28519);
nor U31569 (N_31569,N_28773,N_28641);
or U31570 (N_31570,N_28678,N_28985);
or U31571 (N_31571,N_28834,N_28825);
or U31572 (N_31572,N_29986,N_29655);
nor U31573 (N_31573,N_29461,N_29162);
or U31574 (N_31574,N_29489,N_29307);
nor U31575 (N_31575,N_29013,N_29393);
xor U31576 (N_31576,N_29496,N_28257);
nand U31577 (N_31577,N_29932,N_28687);
nand U31578 (N_31578,N_28614,N_28441);
xor U31579 (N_31579,N_28528,N_28690);
xor U31580 (N_31580,N_29395,N_29610);
or U31581 (N_31581,N_28893,N_28972);
nor U31582 (N_31582,N_28815,N_28806);
xor U31583 (N_31583,N_29338,N_28903);
and U31584 (N_31584,N_29420,N_29412);
xor U31585 (N_31585,N_29542,N_28746);
nand U31586 (N_31586,N_28031,N_28263);
nor U31587 (N_31587,N_29594,N_29180);
and U31588 (N_31588,N_28392,N_28153);
nor U31589 (N_31589,N_29498,N_28644);
nand U31590 (N_31590,N_29858,N_29402);
or U31591 (N_31591,N_29553,N_28135);
or U31592 (N_31592,N_28838,N_28037);
nor U31593 (N_31593,N_29171,N_29393);
or U31594 (N_31594,N_29822,N_28916);
or U31595 (N_31595,N_28712,N_28174);
or U31596 (N_31596,N_28459,N_29335);
and U31597 (N_31597,N_29770,N_28829);
and U31598 (N_31598,N_29967,N_29261);
or U31599 (N_31599,N_29580,N_28578);
nor U31600 (N_31600,N_29403,N_28698);
nand U31601 (N_31601,N_29702,N_28700);
nor U31602 (N_31602,N_28108,N_29239);
xnor U31603 (N_31603,N_29445,N_28663);
xor U31604 (N_31604,N_29011,N_28384);
nor U31605 (N_31605,N_29994,N_29292);
nand U31606 (N_31606,N_28220,N_28815);
and U31607 (N_31607,N_28787,N_29891);
xnor U31608 (N_31608,N_29338,N_29639);
or U31609 (N_31609,N_29121,N_29838);
nand U31610 (N_31610,N_29007,N_28807);
xnor U31611 (N_31611,N_29757,N_28688);
and U31612 (N_31612,N_29704,N_28588);
or U31613 (N_31613,N_29410,N_29752);
and U31614 (N_31614,N_29936,N_29866);
nand U31615 (N_31615,N_28809,N_28697);
nor U31616 (N_31616,N_28133,N_29758);
xor U31617 (N_31617,N_29535,N_29979);
nor U31618 (N_31618,N_29006,N_28162);
or U31619 (N_31619,N_29176,N_29273);
nand U31620 (N_31620,N_28079,N_29465);
nor U31621 (N_31621,N_28323,N_29083);
xor U31622 (N_31622,N_29101,N_29612);
or U31623 (N_31623,N_29545,N_29732);
and U31624 (N_31624,N_29138,N_29357);
or U31625 (N_31625,N_28057,N_29810);
nor U31626 (N_31626,N_28750,N_28428);
xnor U31627 (N_31627,N_28771,N_29489);
nand U31628 (N_31628,N_28389,N_28078);
or U31629 (N_31629,N_28385,N_28214);
and U31630 (N_31630,N_28740,N_29320);
nor U31631 (N_31631,N_28986,N_29966);
xor U31632 (N_31632,N_28590,N_29188);
nand U31633 (N_31633,N_28265,N_28323);
nand U31634 (N_31634,N_28698,N_28369);
and U31635 (N_31635,N_28506,N_29264);
nand U31636 (N_31636,N_28616,N_29577);
nor U31637 (N_31637,N_29855,N_28716);
or U31638 (N_31638,N_29759,N_29973);
nand U31639 (N_31639,N_28932,N_29669);
xnor U31640 (N_31640,N_28894,N_29482);
or U31641 (N_31641,N_28780,N_29593);
or U31642 (N_31642,N_29845,N_28395);
nand U31643 (N_31643,N_29443,N_28389);
and U31644 (N_31644,N_28122,N_28390);
xor U31645 (N_31645,N_29323,N_29618);
and U31646 (N_31646,N_28596,N_29513);
xor U31647 (N_31647,N_28552,N_28589);
and U31648 (N_31648,N_28175,N_29928);
and U31649 (N_31649,N_29314,N_28315);
nand U31650 (N_31650,N_28797,N_29493);
nor U31651 (N_31651,N_28437,N_28110);
or U31652 (N_31652,N_29079,N_29876);
or U31653 (N_31653,N_28169,N_29081);
nand U31654 (N_31654,N_29391,N_29232);
nand U31655 (N_31655,N_28326,N_29936);
xnor U31656 (N_31656,N_28441,N_28982);
and U31657 (N_31657,N_29787,N_28573);
and U31658 (N_31658,N_29050,N_29023);
xor U31659 (N_31659,N_28468,N_29010);
or U31660 (N_31660,N_28376,N_28933);
and U31661 (N_31661,N_28705,N_29089);
nand U31662 (N_31662,N_29997,N_28817);
or U31663 (N_31663,N_29261,N_29178);
nor U31664 (N_31664,N_29332,N_28304);
xnor U31665 (N_31665,N_28958,N_28544);
nand U31666 (N_31666,N_28097,N_28028);
nor U31667 (N_31667,N_29860,N_29402);
nand U31668 (N_31668,N_29432,N_29520);
and U31669 (N_31669,N_28656,N_28533);
and U31670 (N_31670,N_28848,N_28604);
and U31671 (N_31671,N_28607,N_29636);
and U31672 (N_31672,N_29305,N_28474);
or U31673 (N_31673,N_29423,N_28226);
or U31674 (N_31674,N_29308,N_28989);
xor U31675 (N_31675,N_29393,N_28198);
nor U31676 (N_31676,N_29892,N_28438);
xnor U31677 (N_31677,N_28267,N_29545);
nor U31678 (N_31678,N_29055,N_29530);
nand U31679 (N_31679,N_28134,N_28204);
or U31680 (N_31680,N_29489,N_29592);
nor U31681 (N_31681,N_29070,N_28729);
and U31682 (N_31682,N_29525,N_28799);
or U31683 (N_31683,N_28613,N_28388);
and U31684 (N_31684,N_29327,N_28485);
nand U31685 (N_31685,N_29500,N_29305);
nand U31686 (N_31686,N_29674,N_28925);
or U31687 (N_31687,N_29240,N_28570);
or U31688 (N_31688,N_29114,N_28689);
xor U31689 (N_31689,N_29835,N_28880);
nor U31690 (N_31690,N_28406,N_28536);
nand U31691 (N_31691,N_29931,N_29211);
nand U31692 (N_31692,N_28813,N_29747);
xor U31693 (N_31693,N_29368,N_28099);
nand U31694 (N_31694,N_28858,N_29911);
or U31695 (N_31695,N_29429,N_28164);
nand U31696 (N_31696,N_28069,N_28139);
nor U31697 (N_31697,N_29055,N_29844);
nor U31698 (N_31698,N_29618,N_28612);
xnor U31699 (N_31699,N_29128,N_29638);
xnor U31700 (N_31700,N_28293,N_29661);
nor U31701 (N_31701,N_28977,N_28522);
nand U31702 (N_31702,N_28222,N_29371);
xnor U31703 (N_31703,N_28796,N_28930);
and U31704 (N_31704,N_28380,N_28240);
xnor U31705 (N_31705,N_28134,N_29503);
and U31706 (N_31706,N_29533,N_29137);
nand U31707 (N_31707,N_29625,N_28903);
or U31708 (N_31708,N_29542,N_29062);
or U31709 (N_31709,N_28793,N_29077);
or U31710 (N_31710,N_29963,N_28732);
xnor U31711 (N_31711,N_29263,N_29981);
or U31712 (N_31712,N_29341,N_29086);
xnor U31713 (N_31713,N_28209,N_28637);
and U31714 (N_31714,N_28806,N_29565);
and U31715 (N_31715,N_28823,N_28563);
nor U31716 (N_31716,N_29602,N_29085);
nor U31717 (N_31717,N_28390,N_28399);
and U31718 (N_31718,N_29514,N_29016);
and U31719 (N_31719,N_28939,N_28202);
nor U31720 (N_31720,N_29590,N_28592);
and U31721 (N_31721,N_28978,N_28812);
xor U31722 (N_31722,N_29284,N_28387);
and U31723 (N_31723,N_28067,N_28837);
nor U31724 (N_31724,N_28526,N_29605);
and U31725 (N_31725,N_29433,N_29931);
nand U31726 (N_31726,N_28814,N_28245);
nand U31727 (N_31727,N_29536,N_28874);
nor U31728 (N_31728,N_28311,N_29701);
nor U31729 (N_31729,N_29579,N_28620);
or U31730 (N_31730,N_28412,N_28846);
nor U31731 (N_31731,N_29780,N_28573);
and U31732 (N_31732,N_28616,N_28126);
nand U31733 (N_31733,N_29499,N_28043);
nor U31734 (N_31734,N_28162,N_28414);
xnor U31735 (N_31735,N_28814,N_28803);
or U31736 (N_31736,N_29251,N_28146);
and U31737 (N_31737,N_28057,N_28775);
and U31738 (N_31738,N_29615,N_29787);
nor U31739 (N_31739,N_28387,N_28452);
nand U31740 (N_31740,N_29727,N_29872);
nor U31741 (N_31741,N_29339,N_28045);
nand U31742 (N_31742,N_28452,N_29260);
and U31743 (N_31743,N_28815,N_28873);
nand U31744 (N_31744,N_28637,N_29036);
nand U31745 (N_31745,N_29430,N_29842);
and U31746 (N_31746,N_28187,N_28635);
nand U31747 (N_31747,N_28240,N_29159);
nand U31748 (N_31748,N_28865,N_29087);
and U31749 (N_31749,N_29358,N_28015);
xor U31750 (N_31750,N_29262,N_28019);
xor U31751 (N_31751,N_28662,N_28147);
nor U31752 (N_31752,N_29180,N_29122);
xnor U31753 (N_31753,N_29650,N_29492);
and U31754 (N_31754,N_29061,N_29978);
nand U31755 (N_31755,N_28091,N_28758);
nand U31756 (N_31756,N_29295,N_28135);
xor U31757 (N_31757,N_29329,N_29829);
nand U31758 (N_31758,N_28040,N_28982);
and U31759 (N_31759,N_28631,N_29638);
or U31760 (N_31760,N_29220,N_28611);
xor U31761 (N_31761,N_29967,N_28477);
nor U31762 (N_31762,N_29194,N_28113);
or U31763 (N_31763,N_29617,N_28911);
and U31764 (N_31764,N_29002,N_29839);
nor U31765 (N_31765,N_29075,N_28632);
nand U31766 (N_31766,N_28341,N_29520);
nand U31767 (N_31767,N_28340,N_28949);
and U31768 (N_31768,N_28189,N_29400);
nor U31769 (N_31769,N_28809,N_28956);
or U31770 (N_31770,N_29481,N_29090);
or U31771 (N_31771,N_28740,N_28187);
or U31772 (N_31772,N_29624,N_29501);
nand U31773 (N_31773,N_28735,N_29891);
nor U31774 (N_31774,N_28613,N_28830);
and U31775 (N_31775,N_28204,N_29898);
and U31776 (N_31776,N_28313,N_29529);
nand U31777 (N_31777,N_28657,N_28632);
nand U31778 (N_31778,N_29685,N_28505);
xor U31779 (N_31779,N_29171,N_29795);
xnor U31780 (N_31780,N_29323,N_29731);
and U31781 (N_31781,N_29122,N_29783);
xnor U31782 (N_31782,N_29076,N_29094);
or U31783 (N_31783,N_29029,N_29140);
nor U31784 (N_31784,N_28061,N_28472);
nor U31785 (N_31785,N_28044,N_29248);
xnor U31786 (N_31786,N_29290,N_29868);
xor U31787 (N_31787,N_29845,N_28423);
nand U31788 (N_31788,N_29262,N_28829);
or U31789 (N_31789,N_29927,N_28000);
xnor U31790 (N_31790,N_28760,N_28656);
xnor U31791 (N_31791,N_28525,N_29734);
and U31792 (N_31792,N_28141,N_28619);
nand U31793 (N_31793,N_29372,N_29303);
xor U31794 (N_31794,N_29202,N_29246);
or U31795 (N_31795,N_29404,N_29495);
or U31796 (N_31796,N_29925,N_29486);
nor U31797 (N_31797,N_28018,N_29416);
nor U31798 (N_31798,N_28013,N_28790);
nand U31799 (N_31799,N_28481,N_28386);
nor U31800 (N_31800,N_28668,N_28947);
and U31801 (N_31801,N_29198,N_29767);
and U31802 (N_31802,N_29923,N_28795);
and U31803 (N_31803,N_29338,N_29721);
or U31804 (N_31804,N_29193,N_28010);
nor U31805 (N_31805,N_29351,N_29436);
or U31806 (N_31806,N_28896,N_28932);
and U31807 (N_31807,N_29678,N_28572);
nor U31808 (N_31808,N_29810,N_28766);
or U31809 (N_31809,N_28227,N_29807);
nand U31810 (N_31810,N_28404,N_28267);
and U31811 (N_31811,N_29489,N_29188);
and U31812 (N_31812,N_29777,N_29446);
xor U31813 (N_31813,N_29954,N_28770);
or U31814 (N_31814,N_28679,N_29312);
xor U31815 (N_31815,N_28939,N_28382);
or U31816 (N_31816,N_28577,N_28196);
xnor U31817 (N_31817,N_29104,N_28140);
nor U31818 (N_31818,N_29755,N_28378);
xnor U31819 (N_31819,N_29145,N_28131);
nor U31820 (N_31820,N_29776,N_28090);
or U31821 (N_31821,N_29398,N_28080);
nand U31822 (N_31822,N_29896,N_28032);
and U31823 (N_31823,N_29831,N_28785);
and U31824 (N_31824,N_29683,N_28662);
and U31825 (N_31825,N_28482,N_28026);
nor U31826 (N_31826,N_28817,N_28096);
nand U31827 (N_31827,N_29188,N_28968);
nor U31828 (N_31828,N_29924,N_28456);
or U31829 (N_31829,N_29063,N_28701);
xor U31830 (N_31830,N_29632,N_29136);
or U31831 (N_31831,N_28840,N_28316);
or U31832 (N_31832,N_29747,N_28063);
nor U31833 (N_31833,N_28888,N_28188);
and U31834 (N_31834,N_29005,N_29643);
and U31835 (N_31835,N_28764,N_29597);
or U31836 (N_31836,N_29291,N_29578);
or U31837 (N_31837,N_28601,N_28369);
xor U31838 (N_31838,N_29285,N_29174);
and U31839 (N_31839,N_29515,N_28525);
nand U31840 (N_31840,N_29826,N_28597);
nor U31841 (N_31841,N_28946,N_29476);
nand U31842 (N_31842,N_28555,N_28308);
and U31843 (N_31843,N_28401,N_29753);
and U31844 (N_31844,N_28238,N_29577);
and U31845 (N_31845,N_29630,N_28319);
xnor U31846 (N_31846,N_29731,N_29405);
or U31847 (N_31847,N_29825,N_28881);
or U31848 (N_31848,N_28092,N_28527);
or U31849 (N_31849,N_29733,N_29748);
nand U31850 (N_31850,N_28057,N_29557);
nand U31851 (N_31851,N_28921,N_29899);
xor U31852 (N_31852,N_28563,N_28551);
nor U31853 (N_31853,N_29701,N_29770);
xor U31854 (N_31854,N_29704,N_29011);
or U31855 (N_31855,N_28081,N_29986);
or U31856 (N_31856,N_28680,N_29835);
nor U31857 (N_31857,N_28222,N_28236);
and U31858 (N_31858,N_29446,N_28891);
nand U31859 (N_31859,N_28855,N_29993);
nand U31860 (N_31860,N_29089,N_29687);
nor U31861 (N_31861,N_29953,N_28361);
and U31862 (N_31862,N_28946,N_28534);
nor U31863 (N_31863,N_28390,N_28949);
xnor U31864 (N_31864,N_29255,N_28463);
and U31865 (N_31865,N_29865,N_28616);
xor U31866 (N_31866,N_28855,N_29169);
and U31867 (N_31867,N_29181,N_29618);
xor U31868 (N_31868,N_29492,N_29153);
nand U31869 (N_31869,N_29948,N_28170);
or U31870 (N_31870,N_29813,N_29853);
or U31871 (N_31871,N_29069,N_28696);
or U31872 (N_31872,N_28348,N_29416);
and U31873 (N_31873,N_28434,N_29091);
and U31874 (N_31874,N_28123,N_29075);
or U31875 (N_31875,N_28649,N_29087);
nand U31876 (N_31876,N_29525,N_29609);
or U31877 (N_31877,N_28091,N_28321);
or U31878 (N_31878,N_29978,N_28866);
nand U31879 (N_31879,N_28057,N_28090);
or U31880 (N_31880,N_28560,N_28474);
nand U31881 (N_31881,N_28843,N_28787);
and U31882 (N_31882,N_29778,N_28804);
or U31883 (N_31883,N_29029,N_29834);
or U31884 (N_31884,N_29775,N_28173);
nand U31885 (N_31885,N_28392,N_28640);
xor U31886 (N_31886,N_29972,N_29339);
xor U31887 (N_31887,N_28797,N_28974);
xor U31888 (N_31888,N_29155,N_28078);
and U31889 (N_31889,N_28040,N_29984);
and U31890 (N_31890,N_29282,N_29430);
and U31891 (N_31891,N_29671,N_29283);
and U31892 (N_31892,N_28686,N_28227);
or U31893 (N_31893,N_28203,N_29304);
or U31894 (N_31894,N_29443,N_28898);
xnor U31895 (N_31895,N_29658,N_28965);
and U31896 (N_31896,N_28863,N_28246);
and U31897 (N_31897,N_28877,N_29801);
and U31898 (N_31898,N_28321,N_28456);
nor U31899 (N_31899,N_29657,N_29502);
or U31900 (N_31900,N_28895,N_28029);
or U31901 (N_31901,N_29909,N_28746);
nor U31902 (N_31902,N_28748,N_29434);
nand U31903 (N_31903,N_28053,N_28917);
nand U31904 (N_31904,N_28785,N_28754);
or U31905 (N_31905,N_29966,N_29687);
nand U31906 (N_31906,N_29717,N_28794);
and U31907 (N_31907,N_29108,N_29734);
or U31908 (N_31908,N_28411,N_28914);
and U31909 (N_31909,N_28021,N_29507);
xor U31910 (N_31910,N_29905,N_29669);
nor U31911 (N_31911,N_29230,N_29490);
xnor U31912 (N_31912,N_28092,N_29967);
xnor U31913 (N_31913,N_29940,N_28962);
nor U31914 (N_31914,N_29500,N_28762);
and U31915 (N_31915,N_29576,N_29280);
nand U31916 (N_31916,N_29182,N_28602);
nor U31917 (N_31917,N_28247,N_28096);
or U31918 (N_31918,N_29158,N_29285);
xor U31919 (N_31919,N_29894,N_29425);
nand U31920 (N_31920,N_28170,N_29146);
and U31921 (N_31921,N_29917,N_28477);
nand U31922 (N_31922,N_28834,N_29430);
or U31923 (N_31923,N_28754,N_29640);
and U31924 (N_31924,N_28436,N_28463);
nor U31925 (N_31925,N_28052,N_28139);
nand U31926 (N_31926,N_29254,N_29174);
and U31927 (N_31927,N_28824,N_29851);
nor U31928 (N_31928,N_28941,N_28067);
or U31929 (N_31929,N_29581,N_28646);
and U31930 (N_31930,N_28834,N_28398);
xnor U31931 (N_31931,N_28700,N_28150);
nand U31932 (N_31932,N_28075,N_29675);
nor U31933 (N_31933,N_29466,N_28736);
and U31934 (N_31934,N_28790,N_28521);
or U31935 (N_31935,N_29003,N_28721);
nor U31936 (N_31936,N_28325,N_29394);
nor U31937 (N_31937,N_29897,N_28094);
or U31938 (N_31938,N_29817,N_29251);
nand U31939 (N_31939,N_29813,N_29922);
nand U31940 (N_31940,N_28541,N_29696);
xnor U31941 (N_31941,N_29344,N_28929);
nor U31942 (N_31942,N_28997,N_28477);
nor U31943 (N_31943,N_28620,N_28234);
xnor U31944 (N_31944,N_28980,N_28552);
xnor U31945 (N_31945,N_29677,N_29688);
xnor U31946 (N_31946,N_28139,N_29488);
or U31947 (N_31947,N_29125,N_28005);
xnor U31948 (N_31948,N_29321,N_28846);
nor U31949 (N_31949,N_29934,N_28362);
nor U31950 (N_31950,N_28898,N_28395);
nand U31951 (N_31951,N_29414,N_28358);
xor U31952 (N_31952,N_29359,N_29943);
nor U31953 (N_31953,N_28428,N_28102);
and U31954 (N_31954,N_29672,N_28343);
and U31955 (N_31955,N_28122,N_29375);
and U31956 (N_31956,N_28777,N_28312);
nand U31957 (N_31957,N_29264,N_29448);
or U31958 (N_31958,N_28452,N_28795);
or U31959 (N_31959,N_28086,N_29548);
xnor U31960 (N_31960,N_28257,N_28642);
xnor U31961 (N_31961,N_29781,N_28741);
nand U31962 (N_31962,N_29231,N_29092);
xor U31963 (N_31963,N_29912,N_29238);
nor U31964 (N_31964,N_29340,N_28673);
nor U31965 (N_31965,N_28066,N_29045);
nor U31966 (N_31966,N_29915,N_29957);
nand U31967 (N_31967,N_29496,N_28185);
xnor U31968 (N_31968,N_28523,N_28712);
and U31969 (N_31969,N_28845,N_28569);
nor U31970 (N_31970,N_28245,N_28808);
nor U31971 (N_31971,N_29101,N_28651);
xor U31972 (N_31972,N_29598,N_28141);
xnor U31973 (N_31973,N_28334,N_28324);
nor U31974 (N_31974,N_28180,N_29897);
nand U31975 (N_31975,N_28479,N_29087);
and U31976 (N_31976,N_28169,N_28716);
xor U31977 (N_31977,N_29515,N_28873);
xnor U31978 (N_31978,N_28726,N_28293);
nand U31979 (N_31979,N_28404,N_29830);
or U31980 (N_31980,N_29258,N_28706);
nor U31981 (N_31981,N_28964,N_29731);
and U31982 (N_31982,N_29075,N_28538);
nor U31983 (N_31983,N_28690,N_29379);
or U31984 (N_31984,N_29183,N_29396);
and U31985 (N_31985,N_28752,N_29583);
nand U31986 (N_31986,N_29634,N_28439);
nand U31987 (N_31987,N_28379,N_28867);
xor U31988 (N_31988,N_29604,N_29449);
or U31989 (N_31989,N_29244,N_28153);
or U31990 (N_31990,N_28231,N_28776);
xnor U31991 (N_31991,N_29014,N_28772);
xor U31992 (N_31992,N_29902,N_28471);
xor U31993 (N_31993,N_29035,N_29884);
xor U31994 (N_31994,N_29091,N_29823);
or U31995 (N_31995,N_28753,N_28859);
nor U31996 (N_31996,N_29899,N_29581);
nand U31997 (N_31997,N_28813,N_28953);
xnor U31998 (N_31998,N_28792,N_29439);
nand U31999 (N_31999,N_28672,N_28810);
xnor U32000 (N_32000,N_31541,N_31102);
nand U32001 (N_32001,N_30000,N_31063);
xnor U32002 (N_32002,N_31349,N_30946);
xnor U32003 (N_32003,N_31828,N_30470);
xor U32004 (N_32004,N_30276,N_31153);
and U32005 (N_32005,N_31381,N_30612);
nand U32006 (N_32006,N_30977,N_30336);
or U32007 (N_32007,N_30052,N_30143);
nor U32008 (N_32008,N_30613,N_30347);
and U32009 (N_32009,N_31090,N_30845);
and U32010 (N_32010,N_30774,N_30150);
and U32011 (N_32011,N_30917,N_31181);
and U32012 (N_32012,N_31465,N_30211);
and U32013 (N_32013,N_30231,N_30723);
nor U32014 (N_32014,N_30679,N_30009);
nor U32015 (N_32015,N_31737,N_30584);
nand U32016 (N_32016,N_30408,N_31518);
nand U32017 (N_32017,N_30361,N_30323);
nor U32018 (N_32018,N_31348,N_30937);
or U32019 (N_32019,N_30273,N_30804);
and U32020 (N_32020,N_31680,N_31591);
nand U32021 (N_32021,N_30434,N_31879);
and U32022 (N_32022,N_31421,N_31072);
xnor U32023 (N_32023,N_30850,N_30081);
xor U32024 (N_32024,N_31599,N_31588);
or U32025 (N_32025,N_30746,N_31309);
or U32026 (N_32026,N_31075,N_31367);
xor U32027 (N_32027,N_30505,N_30084);
xor U32028 (N_32028,N_30939,N_31423);
or U32029 (N_32029,N_30809,N_31555);
or U32030 (N_32030,N_31960,N_31957);
or U32031 (N_32031,N_30496,N_31499);
nor U32032 (N_32032,N_30719,N_31903);
and U32033 (N_32033,N_30121,N_30979);
nor U32034 (N_32034,N_30127,N_31777);
and U32035 (N_32035,N_31846,N_30563);
nand U32036 (N_32036,N_30327,N_31410);
and U32037 (N_32037,N_30559,N_30521);
or U32038 (N_32038,N_31164,N_30913);
nor U32039 (N_32039,N_30439,N_30762);
xnor U32040 (N_32040,N_30138,N_31700);
and U32041 (N_32041,N_30447,N_31898);
xnor U32042 (N_32042,N_30697,N_31255);
xnor U32043 (N_32043,N_31459,N_30650);
nor U32044 (N_32044,N_31756,N_30145);
or U32045 (N_32045,N_31691,N_30824);
or U32046 (N_32046,N_30004,N_30634);
nand U32047 (N_32047,N_31058,N_30567);
nand U32048 (N_32048,N_31977,N_31498);
or U32049 (N_32049,N_31693,N_30418);
xnor U32050 (N_32050,N_31649,N_31368);
nor U32051 (N_32051,N_30806,N_30229);
and U32052 (N_32052,N_30090,N_31122);
nor U32053 (N_32053,N_31303,N_30486);
or U32054 (N_32054,N_30092,N_31475);
nor U32055 (N_32055,N_31138,N_30450);
and U32056 (N_32056,N_31037,N_31782);
nor U32057 (N_32057,N_31457,N_31572);
xnor U32058 (N_32058,N_31109,N_31483);
xor U32059 (N_32059,N_31187,N_30173);
or U32060 (N_32060,N_30670,N_30346);
xor U32061 (N_32061,N_31811,N_31234);
nand U32062 (N_32062,N_30528,N_31354);
xor U32063 (N_32063,N_30453,N_31748);
xnor U32064 (N_32064,N_30062,N_31794);
or U32065 (N_32065,N_31525,N_30390);
nand U32066 (N_32066,N_30272,N_31476);
xnor U32067 (N_32067,N_30947,N_30250);
xnor U32068 (N_32068,N_31858,N_30763);
or U32069 (N_32069,N_31194,N_30147);
nor U32070 (N_32070,N_31389,N_30732);
or U32071 (N_32071,N_31160,N_31983);
nor U32072 (N_32072,N_31820,N_30747);
xor U32073 (N_32073,N_30733,N_31590);
or U32074 (N_32074,N_31778,N_31694);
or U32075 (N_32075,N_30476,N_31824);
nor U32076 (N_32076,N_31647,N_30295);
xnor U32077 (N_32077,N_31031,N_31620);
nand U32078 (N_32078,N_31056,N_30543);
or U32079 (N_32079,N_31540,N_31258);
nand U32080 (N_32080,N_31472,N_31965);
nand U32081 (N_32081,N_31874,N_30951);
nor U32082 (N_32082,N_31297,N_30045);
and U32083 (N_32083,N_30619,N_31639);
xor U32084 (N_32084,N_31909,N_31026);
nand U32085 (N_32085,N_30233,N_31600);
nor U32086 (N_32086,N_30588,N_30638);
nand U32087 (N_32087,N_30134,N_31841);
nand U32088 (N_32088,N_31968,N_31652);
xor U32089 (N_32089,N_31670,N_30339);
nand U32090 (N_32090,N_31534,N_30226);
xnor U32091 (N_32091,N_31329,N_30862);
nand U32092 (N_32092,N_30247,N_31514);
nor U32093 (N_32093,N_30648,N_31463);
nor U32094 (N_32094,N_31688,N_31994);
or U32095 (N_32095,N_30545,N_31615);
or U32096 (N_32096,N_31361,N_30888);
nand U32097 (N_32097,N_30017,N_30088);
and U32098 (N_32098,N_30596,N_30483);
nor U32099 (N_32099,N_30105,N_31192);
nand U32100 (N_32100,N_31814,N_31485);
xnor U32101 (N_32101,N_31658,N_30717);
and U32102 (N_32102,N_30113,N_30050);
nor U32103 (N_32103,N_31034,N_30654);
or U32104 (N_32104,N_30256,N_31486);
nand U32105 (N_32105,N_30311,N_31195);
nor U32106 (N_32106,N_31139,N_30731);
or U32107 (N_32107,N_30963,N_31889);
nand U32108 (N_32108,N_30674,N_31071);
and U32109 (N_32109,N_31640,N_30886);
nor U32110 (N_32110,N_30421,N_30071);
nand U32111 (N_32111,N_31511,N_31614);
xor U32112 (N_32112,N_30512,N_31079);
xnor U32113 (N_32113,N_31871,N_30729);
nor U32114 (N_32114,N_31370,N_31251);
nor U32115 (N_32115,N_31964,N_30156);
nand U32116 (N_32116,N_31337,N_30368);
or U32117 (N_32117,N_30460,N_30383);
or U32118 (N_32118,N_31262,N_31044);
nor U32119 (N_32119,N_30086,N_30076);
xnor U32120 (N_32120,N_31531,N_31467);
nand U32121 (N_32121,N_31736,N_30793);
xor U32122 (N_32122,N_31808,N_30877);
and U32123 (N_32123,N_31931,N_30966);
nor U32124 (N_32124,N_30176,N_31107);
nand U32125 (N_32125,N_30915,N_30669);
nor U32126 (N_32126,N_30676,N_31307);
and U32127 (N_32127,N_31581,N_30645);
nand U32128 (N_32128,N_30234,N_30152);
or U32129 (N_32129,N_30974,N_31692);
nor U32130 (N_32130,N_30827,N_31461);
and U32131 (N_32131,N_30182,N_30309);
and U32132 (N_32132,N_31260,N_30270);
nor U32133 (N_32133,N_30644,N_31850);
nor U32134 (N_32134,N_30942,N_30474);
xor U32135 (N_32135,N_30290,N_31690);
xnor U32136 (N_32136,N_30403,N_31781);
and U32137 (N_32137,N_30277,N_31863);
nor U32138 (N_32138,N_31018,N_31506);
or U32139 (N_32139,N_30249,N_30056);
nand U32140 (N_32140,N_30704,N_31041);
or U32141 (N_32141,N_31395,N_31248);
xnor U32142 (N_32142,N_30195,N_31403);
nor U32143 (N_32143,N_31259,N_31628);
xnor U32144 (N_32144,N_30519,N_30328);
nand U32145 (N_32145,N_31594,N_31523);
or U32146 (N_32146,N_31356,N_31012);
or U32147 (N_32147,N_30712,N_31807);
xor U32148 (N_32148,N_31085,N_30938);
nor U32149 (N_32149,N_30819,N_31979);
xor U32150 (N_32150,N_31664,N_30627);
or U32151 (N_32151,N_30536,N_31972);
nand U32152 (N_32152,N_30794,N_30671);
nand U32153 (N_32153,N_31944,N_30223);
nand U32154 (N_32154,N_31171,N_30040);
and U32155 (N_32155,N_31415,N_30841);
or U32156 (N_32156,N_30203,N_31228);
nor U32157 (N_32157,N_31870,N_30666);
and U32158 (N_32158,N_31478,N_31733);
nand U32159 (N_32159,N_30769,N_31915);
and U32160 (N_32160,N_31891,N_30060);
and U32161 (N_32161,N_31646,N_30681);
or U32162 (N_32162,N_30139,N_31270);
or U32163 (N_32163,N_30049,N_30120);
xor U32164 (N_32164,N_30326,N_31491);
nand U32165 (N_32165,N_31509,N_30068);
nand U32166 (N_32166,N_31515,N_30271);
nand U32167 (N_32167,N_30986,N_30846);
nor U32168 (N_32168,N_31477,N_30266);
xnor U32169 (N_32169,N_30218,N_31721);
xnor U32170 (N_32170,N_31254,N_30950);
nand U32171 (N_32171,N_30401,N_31943);
or U32172 (N_32172,N_30192,N_30541);
xor U32173 (N_32173,N_31454,N_31460);
xnor U32174 (N_32174,N_31859,N_30611);
nand U32175 (N_32175,N_31150,N_30014);
and U32176 (N_32176,N_30789,N_30727);
nor U32177 (N_32177,N_30212,N_30167);
or U32178 (N_32178,N_30861,N_31050);
nand U32179 (N_32179,N_30910,N_30720);
nand U32180 (N_32180,N_30817,N_30659);
nand U32181 (N_32181,N_30236,N_31411);
nand U32182 (N_32182,N_31554,N_30464);
or U32183 (N_32183,N_30906,N_30059);
or U32184 (N_32184,N_30377,N_30924);
xor U32185 (N_32185,N_31273,N_30007);
xnor U32186 (N_32186,N_31645,N_30184);
nor U32187 (N_32187,N_31057,N_30854);
nand U32188 (N_32188,N_31180,N_30376);
and U32189 (N_32189,N_31978,N_30183);
xor U32190 (N_32190,N_31526,N_30716);
and U32191 (N_32191,N_30248,N_31047);
or U32192 (N_32192,N_31829,N_30481);
or U32193 (N_32193,N_30471,N_30998);
nand U32194 (N_32194,N_31559,N_30170);
and U32195 (N_32195,N_30207,N_30340);
and U32196 (N_32196,N_30655,N_30503);
nor U32197 (N_32197,N_30104,N_30750);
or U32198 (N_32198,N_31765,N_31970);
and U32199 (N_32199,N_31752,N_30061);
nor U32200 (N_32200,N_30604,N_31165);
nand U32201 (N_32201,N_30356,N_30829);
xnor U32202 (N_32202,N_31061,N_30482);
nand U32203 (N_32203,N_30085,N_31834);
xnor U32204 (N_32204,N_31785,N_30805);
or U32205 (N_32205,N_30119,N_30890);
or U32206 (N_32206,N_31685,N_30919);
xor U32207 (N_32207,N_31622,N_31104);
nand U32208 (N_32208,N_30055,N_31082);
or U32209 (N_32209,N_31267,N_31039);
xnor U32210 (N_32210,N_31113,N_31562);
xor U32211 (N_32211,N_30849,N_30527);
nor U32212 (N_32212,N_30653,N_31200);
nor U32213 (N_32213,N_31028,N_30435);
nand U32214 (N_32214,N_30948,N_31768);
or U32215 (N_32215,N_30180,N_31856);
or U32216 (N_32216,N_31636,N_30570);
nor U32217 (N_32217,N_31519,N_31009);
or U32218 (N_32218,N_31655,N_31576);
or U32219 (N_32219,N_31775,N_31504);
or U32220 (N_32220,N_31543,N_31470);
nor U32221 (N_32221,N_30770,N_30440);
and U32222 (N_32222,N_30590,N_30952);
nor U32223 (N_32223,N_30033,N_31967);
xor U32224 (N_32224,N_30251,N_31585);
nand U32225 (N_32225,N_31791,N_31015);
nand U32226 (N_32226,N_30530,N_31320);
nor U32227 (N_32227,N_30920,N_30832);
and U32228 (N_32228,N_31822,N_30870);
or U32229 (N_32229,N_31098,N_30691);
xnor U32230 (N_32230,N_31168,N_31278);
and U32231 (N_32231,N_30564,N_31738);
nand U32232 (N_32232,N_31637,N_31002);
xor U32233 (N_32233,N_31099,N_31582);
or U32234 (N_32234,N_31988,N_30808);
xor U32235 (N_32235,N_31346,N_30420);
xor U32236 (N_32236,N_31689,N_31656);
nor U32237 (N_32237,N_30131,N_31275);
nor U32238 (N_32238,N_31433,N_31631);
xnor U32239 (N_32239,N_30889,N_31535);
nand U32240 (N_32240,N_31607,N_31326);
xor U32241 (N_32241,N_30740,N_31265);
and U32242 (N_32242,N_31579,N_31793);
nand U32243 (N_32243,N_30518,N_30760);
nand U32244 (N_32244,N_31293,N_31608);
nor U32245 (N_32245,N_31017,N_30466);
nand U32246 (N_32246,N_30488,N_31351);
nand U32247 (N_32247,N_30546,N_30661);
xnor U32248 (N_32248,N_30607,N_31279);
or U32249 (N_32249,N_31862,N_31991);
nand U32250 (N_32250,N_31000,N_30244);
nand U32251 (N_32251,N_31431,N_30043);
nand U32252 (N_32252,N_30548,N_30856);
and U32253 (N_32253,N_31202,N_30359);
nor U32254 (N_32254,N_30199,N_30755);
xor U32255 (N_32255,N_30267,N_30191);
xor U32256 (N_32256,N_31705,N_30868);
or U32257 (N_32257,N_30433,N_31152);
nand U32258 (N_32258,N_31833,N_30316);
and U32259 (N_32259,N_31920,N_30773);
or U32260 (N_32260,N_31635,N_31767);
or U32261 (N_32261,N_30128,N_30269);
nor U32262 (N_32262,N_30949,N_31537);
xor U32263 (N_32263,N_31069,N_30100);
and U32264 (N_32264,N_31065,N_31634);
nor U32265 (N_32265,N_31735,N_30992);
xor U32266 (N_32266,N_30651,N_31289);
nor U32267 (N_32267,N_31819,N_31792);
nand U32268 (N_32268,N_30916,N_30903);
nor U32269 (N_32269,N_31040,N_31757);
and U32270 (N_32270,N_30578,N_31203);
nor U32271 (N_32271,N_31908,N_31023);
nand U32272 (N_32272,N_30204,N_31584);
nor U32273 (N_32273,N_31261,N_31449);
nor U32274 (N_32274,N_31276,N_31376);
or U32275 (N_32275,N_31740,N_31088);
xor U32276 (N_32276,N_31712,N_31038);
xnor U32277 (N_32277,N_30855,N_31352);
xor U32278 (N_32278,N_31698,N_30800);
nor U32279 (N_32279,N_31338,N_30324);
xnor U32280 (N_32280,N_30032,N_30767);
or U32281 (N_32281,N_31003,N_31512);
xnor U32282 (N_32282,N_31084,N_30175);
or U32283 (N_32283,N_30363,N_30737);
nand U32284 (N_32284,N_30797,N_30874);
and U32285 (N_32285,N_31042,N_31335);
and U32286 (N_32286,N_30605,N_30550);
and U32287 (N_32287,N_30451,N_31849);
nand U32288 (N_32288,N_31055,N_31216);
xor U32289 (N_32289,N_31215,N_31604);
nor U32290 (N_32290,N_30784,N_31547);
xnor U32291 (N_32291,N_30148,N_30109);
or U32292 (N_32292,N_31188,N_30053);
nor U32293 (N_32293,N_30853,N_30169);
nand U32294 (N_32294,N_30066,N_30102);
or U32295 (N_32295,N_30629,N_30703);
nor U32296 (N_32296,N_31105,N_30023);
and U32297 (N_32297,N_31847,N_30673);
xnor U32298 (N_32298,N_31126,N_31949);
nand U32299 (N_32299,N_31971,N_30446);
and U32300 (N_32300,N_30786,N_30608);
and U32301 (N_32301,N_30472,N_31306);
or U32302 (N_32302,N_31696,N_31049);
nor U32303 (N_32303,N_30414,N_30111);
nand U32304 (N_32304,N_31825,N_31115);
and U32305 (N_32305,N_31494,N_30279);
xnor U32306 (N_32306,N_30335,N_31976);
nor U32307 (N_32307,N_31810,N_30778);
or U32308 (N_32308,N_30477,N_31672);
and U32309 (N_32309,N_30502,N_30286);
nor U32310 (N_32310,N_30073,N_30840);
nand U32311 (N_32311,N_31035,N_31795);
nand U32312 (N_32312,N_31996,N_31663);
nor U32313 (N_32313,N_31837,N_30625);
xor U32314 (N_32314,N_30652,N_30308);
xnor U32315 (N_32315,N_31927,N_30338);
xor U32316 (N_32316,N_31861,N_30643);
nor U32317 (N_32317,N_30162,N_31953);
nor U32318 (N_32318,N_31893,N_30179);
xor U32319 (N_32319,N_31832,N_30662);
nand U32320 (N_32320,N_31360,N_31549);
nor U32321 (N_32321,N_30141,N_31148);
nor U32322 (N_32322,N_31448,N_31571);
and U32323 (N_32323,N_30372,N_31186);
nor U32324 (N_32324,N_30258,N_30364);
nand U32325 (N_32325,N_30198,N_30458);
xnor U32326 (N_32326,N_30771,N_31416);
and U32327 (N_32327,N_31157,N_31564);
or U32328 (N_32328,N_31106,N_31958);
and U32329 (N_32329,N_30798,N_31229);
nor U32330 (N_32330,N_30463,N_30161);
xor U32331 (N_32331,N_31391,N_30956);
nand U32332 (N_32332,N_30663,N_30900);
nor U32333 (N_32333,N_30686,N_30116);
and U32334 (N_32334,N_30557,N_31089);
or U32335 (N_32335,N_31173,N_31653);
xnor U32336 (N_32336,N_30260,N_31045);
or U32337 (N_32337,N_30394,N_30858);
and U32338 (N_32338,N_30219,N_31442);
or U32339 (N_32339,N_30415,N_31095);
or U32340 (N_32340,N_30304,N_30298);
and U32341 (N_32341,N_31166,N_31046);
or U32342 (N_32342,N_31169,N_31372);
xor U32343 (N_32343,N_31926,N_30475);
xnor U32344 (N_32344,N_30788,N_31678);
or U32345 (N_32345,N_31159,N_30738);
nor U32346 (N_32346,N_31539,N_31980);
or U32347 (N_32347,N_30254,N_31134);
or U32348 (N_32348,N_31438,N_30871);
or U32349 (N_32349,N_30754,N_30287);
and U32350 (N_32350,N_30351,N_31196);
or U32351 (N_32351,N_31995,N_30695);
nor U32352 (N_32352,N_30239,N_30454);
and U32353 (N_32353,N_30144,N_31342);
nor U32354 (N_32354,N_30264,N_30462);
and U32355 (N_32355,N_30558,N_31605);
nand U32356 (N_32356,N_31030,N_31008);
nor U32357 (N_32357,N_30407,N_30230);
xnor U32358 (N_32358,N_30668,N_31921);
or U32359 (N_32359,N_30801,N_31162);
or U32360 (N_32360,N_31884,N_31366);
xnor U32361 (N_32361,N_30715,N_31412);
nand U32362 (N_32362,N_30540,N_30744);
or U32363 (N_32363,N_30305,N_31630);
and U32364 (N_32364,N_31899,N_30772);
nand U32365 (N_32365,N_31742,N_31906);
nand U32366 (N_32366,N_30333,N_31144);
or U32367 (N_32367,N_30636,N_30030);
xor U32368 (N_32368,N_31311,N_30206);
nor U32369 (N_32369,N_31520,N_30021);
and U32370 (N_32370,N_31201,N_30334);
nor U32371 (N_32371,N_31211,N_31732);
or U32372 (N_32372,N_31238,N_30960);
nand U32373 (N_32373,N_31805,N_30107);
nor U32374 (N_32374,N_30628,N_31129);
or U32375 (N_32375,N_31789,N_30430);
xnor U32376 (N_32376,N_31172,N_30240);
nor U32377 (N_32377,N_31557,N_30884);
nand U32378 (N_32378,N_31827,N_30232);
and U32379 (N_32379,N_31660,N_31324);
or U32380 (N_32380,N_31932,N_31316);
xnor U32381 (N_32381,N_31638,N_30722);
or U32382 (N_32382,N_30424,N_30572);
or U32383 (N_32383,N_31219,N_31838);
and U32384 (N_32384,N_30555,N_31623);
and U32385 (N_32385,N_30523,N_31945);
nor U32386 (N_32386,N_31930,N_30097);
nor U32387 (N_32387,N_31569,N_30675);
or U32388 (N_32388,N_30278,N_31051);
nor U32389 (N_32389,N_31418,N_31242);
xnor U32390 (N_32390,N_30027,N_30125);
nand U32391 (N_32391,N_30469,N_31709);
nand U32392 (N_32392,N_31142,N_31546);
and U32393 (N_32393,N_31529,N_31632);
xnor U32394 (N_32394,N_30412,N_30114);
nand U32395 (N_32395,N_30549,N_31011);
or U32396 (N_32396,N_30765,N_30997);
and U32397 (N_32397,N_31568,N_31093);
nor U32398 (N_32398,N_31676,N_31365);
and U32399 (N_32399,N_31125,N_31493);
or U32400 (N_32400,N_30404,N_30422);
nor U32401 (N_32401,N_30885,N_30205);
nand U32402 (N_32402,N_31813,N_30489);
nor U32403 (N_32403,N_31052,N_30582);
and U32404 (N_32404,N_30766,N_31759);
xnor U32405 (N_32405,N_30498,N_31377);
nand U32406 (N_32406,N_31854,N_30132);
and U32407 (N_32407,N_31231,N_31441);
or U32408 (N_32408,N_31249,N_31116);
nor U32409 (N_32409,N_30830,N_31062);
nor U32410 (N_32410,N_30665,N_31675);
xnor U32411 (N_32411,N_31434,N_31388);
nor U32412 (N_32412,N_30796,N_30002);
xnor U32413 (N_32413,N_31758,N_30616);
or U32414 (N_32414,N_30379,N_31078);
xnor U32415 (N_32415,N_30994,N_30705);
or U32416 (N_32416,N_31016,N_30388);
and U32417 (N_32417,N_31386,N_30449);
nand U32418 (N_32418,N_31524,N_30525);
xnor U32419 (N_32419,N_30544,N_31161);
or U32420 (N_32420,N_31083,N_31176);
or U32421 (N_32421,N_31487,N_30042);
nor U32422 (N_32422,N_31703,N_31488);
xnor U32423 (N_32423,N_30089,N_30566);
or U32424 (N_32424,N_30930,N_31288);
nand U32425 (N_32425,N_30171,N_30151);
and U32426 (N_32426,N_31048,N_31885);
or U32427 (N_32427,N_30013,N_30079);
xor U32428 (N_32428,N_30358,N_30932);
and U32429 (N_32429,N_30431,N_30442);
and U32430 (N_32430,N_31182,N_30690);
xor U32431 (N_32431,N_31786,N_31521);
and U32432 (N_32432,N_30641,N_30136);
and U32433 (N_32433,N_31956,N_31390);
xor U32434 (N_32434,N_31801,N_30228);
and U32435 (N_32435,N_30243,N_31214);
or U32436 (N_32436,N_31745,N_30200);
or U32437 (N_32437,N_30350,N_30225);
nand U32438 (N_32438,N_31818,N_30553);
or U32439 (N_32439,N_30093,N_31277);
nand U32440 (N_32440,N_31866,N_31650);
and U32441 (N_32441,N_31193,N_30034);
or U32442 (N_32442,N_31916,N_31776);
xnor U32443 (N_32443,N_31292,N_31603);
and U32444 (N_32444,N_30678,N_31310);
and U32445 (N_32445,N_30208,N_30876);
xnor U32446 (N_32446,N_30314,N_31059);
nand U32447 (N_32447,N_31425,N_31671);
nand U32448 (N_32448,N_31140,N_31661);
and U32449 (N_32449,N_31385,N_31401);
xor U32450 (N_32450,N_31420,N_31235);
xor U32451 (N_32451,N_31986,N_31888);
or U32452 (N_32452,N_30516,N_31305);
xnor U32453 (N_32453,N_31806,N_31067);
and U32454 (N_32454,N_31127,N_31598);
and U32455 (N_32455,N_30293,N_30852);
or U32456 (N_32456,N_31206,N_30971);
nand U32457 (N_32457,N_30576,N_31981);
nor U32458 (N_32458,N_31674,N_30818);
and U32459 (N_32459,N_30702,N_30878);
and U32460 (N_32460,N_30063,N_31299);
nor U32461 (N_32461,N_31340,N_30560);
and U32462 (N_32462,N_31007,N_31677);
or U32463 (N_32463,N_30891,N_31302);
and U32464 (N_32464,N_31892,N_31704);
or U32465 (N_32465,N_31087,N_31923);
nor U32466 (N_32466,N_31816,N_31642);
nor U32467 (N_32467,N_30163,N_31706);
xor U32468 (N_32468,N_31803,N_30280);
or U32469 (N_32469,N_30713,N_30775);
and U32470 (N_32470,N_30494,N_30303);
and U32471 (N_32471,N_30756,N_31271);
xnor U32472 (N_32472,N_30217,N_31151);
or U32473 (N_32473,N_31984,N_30345);
or U32474 (N_32474,N_31120,N_31440);
nor U32475 (N_32475,N_30393,N_31882);
or U32476 (N_32476,N_30317,N_31618);
and U32477 (N_32477,N_31577,N_31779);
nor U32478 (N_32478,N_31332,N_31027);
or U32479 (N_32479,N_30904,N_31359);
nor U32480 (N_32480,N_30467,N_31496);
nor U32481 (N_32481,N_30301,N_31887);
xor U32482 (N_32482,N_30517,N_31734);
nor U32483 (N_32483,N_30133,N_31350);
or U32484 (N_32484,N_31300,N_30753);
and U32485 (N_32485,N_30640,N_30001);
nor U32486 (N_32486,N_30814,N_31341);
nor U32487 (N_32487,N_30416,N_31843);
and U32488 (N_32488,N_30759,N_30872);
nor U32489 (N_32489,N_30700,N_31597);
nand U32490 (N_32490,N_30480,N_30983);
nand U32491 (N_32491,N_30907,N_31408);
xnor U32492 (N_32492,N_30820,N_30378);
xnor U32493 (N_32493,N_31933,N_30851);
or U32494 (N_32494,N_31548,N_30583);
and U32495 (N_32495,N_30322,N_31596);
xnor U32496 (N_32496,N_31137,N_31054);
nand U32497 (N_32497,N_31840,N_31100);
and U32498 (N_32498,N_30255,N_30883);
and U32499 (N_32499,N_31240,N_31975);
nand U32500 (N_32500,N_31327,N_30826);
and U32501 (N_32501,N_31830,N_30689);
xor U32502 (N_32502,N_30010,N_31070);
or U32503 (N_32503,N_31823,N_31429);
and U32504 (N_32504,N_31405,N_30126);
xor U32505 (N_32505,N_31220,N_31955);
xor U32506 (N_32506,N_31753,N_30529);
and U32507 (N_32507,N_30776,N_31938);
nand U32508 (N_32508,N_31896,N_30365);
nand U32509 (N_32509,N_30658,N_30610);
xor U32510 (N_32510,N_30623,N_31298);
nor U32511 (N_32511,N_31301,N_31317);
xnor U32512 (N_32512,N_31333,N_31993);
nor U32513 (N_32513,N_31667,N_30098);
xor U32514 (N_32514,N_31595,N_30828);
or U32515 (N_32515,N_31924,N_31741);
or U32516 (N_32516,N_31602,N_30461);
nor U32517 (N_32517,N_30508,N_30539);
nand U32518 (N_32518,N_30058,N_30222);
xor U32519 (N_32519,N_30041,N_31112);
or U32520 (N_32520,N_30812,N_30914);
nor U32521 (N_32521,N_31130,N_30506);
nand U32522 (N_32522,N_30561,N_31189);
xor U32523 (N_32523,N_31178,N_30172);
and U32524 (N_32524,N_31713,N_31437);
xnor U32525 (N_32525,N_30898,N_30585);
xnor U32526 (N_32526,N_30693,N_30976);
nor U32527 (N_32527,N_31580,N_31839);
or U32528 (N_32528,N_31593,N_31729);
or U32529 (N_32529,N_30174,N_31005);
or U32530 (N_32530,N_30822,N_30005);
or U32531 (N_32531,N_30112,N_30321);
and U32532 (N_32532,N_30892,N_31252);
nor U32533 (N_32533,N_31029,N_31147);
nand U32534 (N_32534,N_30284,N_31681);
or U32535 (N_32535,N_30140,N_30815);
xnor U32536 (N_32536,N_31358,N_30902);
or U32537 (N_32537,N_30238,N_30875);
xnor U32538 (N_32538,N_31990,N_30709);
nand U32539 (N_32539,N_30288,N_30263);
nand U32540 (N_32540,N_30901,N_31804);
nand U32541 (N_32541,N_31852,N_31369);
nand U32542 (N_32542,N_31935,N_30387);
xor U32543 (N_32543,N_30984,N_30209);
and U32544 (N_32544,N_30777,N_31239);
and U32545 (N_32545,N_31154,N_30028);
or U32546 (N_32546,N_30757,N_31272);
or U32547 (N_32547,N_31019,N_31744);
and U32548 (N_32548,N_31118,N_31687);
or U32549 (N_32549,N_30562,N_30514);
nand U32550 (N_32550,N_31197,N_31722);
nor U32551 (N_32551,N_31780,N_30122);
or U32552 (N_32552,N_30070,N_31318);
or U32553 (N_32553,N_30554,N_30300);
or U32554 (N_32554,N_31175,N_31308);
and U32555 (N_32555,N_31469,N_31379);
xnor U32556 (N_32556,N_31424,N_31080);
nand U32557 (N_32557,N_31553,N_31396);
nand U32558 (N_32558,N_31191,N_31290);
nor U32559 (N_32559,N_31560,N_30265);
or U32560 (N_32560,N_31266,N_30108);
nor U32561 (N_32561,N_30310,N_30146);
nand U32562 (N_32562,N_31092,N_31682);
and U32563 (N_32563,N_30943,N_31077);
or U32564 (N_32564,N_30600,N_31263);
and U32565 (N_32565,N_31575,N_31330);
and U32566 (N_32566,N_30096,N_30593);
xor U32567 (N_32567,N_31679,N_30123);
or U32568 (N_32568,N_31146,N_30166);
nor U32569 (N_32569,N_30838,N_30707);
nand U32570 (N_32570,N_31947,N_31123);
xor U32571 (N_32571,N_30094,N_30577);
or U32572 (N_32572,N_31797,N_31245);
nand U32573 (N_32573,N_31627,N_31398);
or U32574 (N_32574,N_30510,N_31886);
and U32575 (N_32575,N_30373,N_30542);
nand U32576 (N_32576,N_30443,N_31336);
xor U32577 (N_32577,N_31136,N_31666);
and U32578 (N_32578,N_30432,N_31720);
nand U32579 (N_32579,N_30909,N_31445);
nor U32580 (N_32580,N_30428,N_31091);
xor U32581 (N_32581,N_30843,N_30513);
nand U32582 (N_32582,N_30398,N_30025);
xnor U32583 (N_32583,N_31545,N_30664);
xnor U32584 (N_32584,N_31387,N_31826);
or U32585 (N_32585,N_30501,N_30245);
nor U32586 (N_32586,N_30465,N_30745);
and U32587 (N_32587,N_31974,N_30315);
nor U32588 (N_32588,N_30833,N_31695);
xnor U32589 (N_32589,N_30402,N_31802);
nand U32590 (N_32590,N_30609,N_31668);
and U32591 (N_32591,N_30186,N_30580);
xor U32592 (N_32592,N_30614,N_30500);
and U32593 (N_32593,N_31257,N_30242);
nor U32594 (N_32594,N_31480,N_30395);
and U32595 (N_32595,N_30534,N_31589);
nor U32596 (N_32596,N_30455,N_31497);
nand U32597 (N_32597,N_30227,N_30618);
or U32598 (N_32598,N_30926,N_30893);
nand U32599 (N_32599,N_31353,N_31625);
nand U32600 (N_32600,N_30160,N_31371);
or U32601 (N_32601,N_31502,N_30425);
nor U32602 (N_32602,N_31185,N_31578);
and U32603 (N_32603,N_31728,N_31513);
nor U32604 (N_32604,N_31836,N_30741);
nor U32605 (N_32605,N_31948,N_31081);
nor U32606 (N_32606,N_31285,N_31533);
nor U32607 (N_32607,N_31724,N_31998);
xnor U32608 (N_32608,N_30135,N_31024);
nor U32609 (N_32609,N_30024,N_30399);
and U32610 (N_32610,N_30834,N_31264);
xnor U32611 (N_32611,N_30426,N_30202);
or U32612 (N_32612,N_30353,N_30294);
nor U32613 (N_32613,N_31914,N_30839);
and U32614 (N_32614,N_31436,N_31961);
nand U32615 (N_32615,N_30036,N_31362);
and U32616 (N_32616,N_31225,N_31959);
or U32617 (N_32617,N_30292,N_30688);
nand U32618 (N_32618,N_30999,N_30799);
and U32619 (N_32619,N_30711,N_31110);
or U32620 (N_32620,N_30241,N_30342);
and U32621 (N_32621,N_31426,N_31014);
or U32622 (N_32622,N_30831,N_30880);
xnor U32623 (N_32623,N_31458,N_31455);
nand U32624 (N_32624,N_31845,N_30331);
xor U32625 (N_32625,N_30982,N_31747);
or U32626 (N_32626,N_31339,N_30103);
and U32627 (N_32627,N_31177,N_31982);
nor U32628 (N_32628,N_31280,N_30635);
xnor U32629 (N_32629,N_31905,N_30473);
nor U32630 (N_32630,N_31707,N_30130);
nand U32631 (N_32631,N_31875,N_30057);
or U32632 (N_32632,N_30268,N_31821);
nand U32633 (N_32633,N_30193,N_31962);
or U32634 (N_32634,N_30779,N_31864);
xnor U32635 (N_32635,N_31274,N_30035);
and U32636 (N_32636,N_30253,N_30330);
nor U32637 (N_32637,N_31877,N_31626);
and U32638 (N_32638,N_30811,N_31925);
or U32639 (N_32639,N_30008,N_30499);
xnor U32640 (N_32640,N_31873,N_30468);
nand U32641 (N_32641,N_30594,N_30213);
and U32642 (N_32642,N_30923,N_30142);
xnor U32643 (N_32643,N_31556,N_31474);
and U32644 (N_32644,N_31243,N_30597);
nor U32645 (N_32645,N_30391,N_30620);
xor U32646 (N_32646,N_30406,N_31851);
and U32647 (N_32647,N_31612,N_31432);
xnor U32648 (N_32648,N_30887,N_31450);
xnor U32649 (N_32649,N_31209,N_31773);
nand U32650 (N_32650,N_30237,N_30348);
and U32651 (N_32651,N_30275,N_30369);
or U32652 (N_32652,N_31479,N_31815);
xor U32653 (N_32653,N_30190,N_30220);
and U32654 (N_32654,N_31281,N_31451);
and U32655 (N_32655,N_30896,N_31439);
nand U32656 (N_32656,N_31809,N_30694);
or U32657 (N_32657,N_30087,N_30758);
and U32658 (N_32658,N_30341,N_30929);
nand U32659 (N_32659,N_30781,N_31566);
nor U32660 (N_32660,N_30708,N_31587);
nand U32661 (N_32661,N_31783,N_30411);
xnor U32662 (N_32662,N_30046,N_30864);
xor U32663 (N_32663,N_30185,N_31244);
xnor U32664 (N_32664,N_31073,N_31314);
or U32665 (N_32665,N_31796,N_30721);
and U32666 (N_32666,N_31155,N_30410);
and U32667 (N_32667,N_31156,N_30687);
nand U32668 (N_32668,N_30297,N_31374);
nand U32669 (N_32669,N_31375,N_31880);
nor U32670 (N_32670,N_30285,N_30457);
nand U32671 (N_32671,N_31552,N_31328);
or U32672 (N_32672,N_30569,N_30165);
nand U32673 (N_32673,N_31609,N_31999);
and U32674 (N_32674,N_31895,N_30064);
xnor U32675 (N_32675,N_30785,N_31218);
nor U32676 (N_32676,N_31718,N_31223);
nand U32677 (N_32677,N_30989,N_30615);
nand U32678 (N_32678,N_30177,N_30187);
xor U32679 (N_32679,N_31912,N_30188);
nor U32680 (N_32680,N_31657,N_31384);
nor U32681 (N_32681,N_30624,N_30456);
or U32682 (N_32682,N_30621,N_31842);
nand U32683 (N_32683,N_30825,N_31881);
nor U32684 (N_32684,N_31236,N_31226);
and U32685 (N_32685,N_30224,N_30642);
nand U32686 (N_32686,N_30685,N_31997);
nand U32687 (N_32687,N_31939,N_31659);
nand U32688 (N_32688,N_31364,N_31743);
nor U32689 (N_32689,N_31701,N_30867);
and U32690 (N_32690,N_30730,N_31501);
and U32691 (N_32691,N_31022,N_30537);
nand U32692 (N_32692,N_30332,N_31253);
xnor U32693 (N_32693,N_30429,N_30441);
nor U32694 (N_32694,N_31158,N_31446);
and U32695 (N_32695,N_31505,N_30178);
xnor U32696 (N_32696,N_30925,N_31883);
xnor U32697 (N_32697,N_31787,N_30955);
nand U32698 (N_32698,N_31510,N_31283);
or U32699 (N_32699,N_31001,N_31357);
and U32700 (N_32700,N_30863,N_31101);
and U32701 (N_32701,N_31284,N_30633);
nor U32702 (N_32702,N_31500,N_30684);
xnor U32703 (N_32703,N_31710,N_30405);
or U32704 (N_32704,N_30724,N_31711);
nor U32705 (N_32705,N_30532,N_31522);
and U32706 (N_32706,N_30957,N_30319);
nand U32707 (N_32707,N_31068,N_31133);
and U32708 (N_32708,N_30296,N_30080);
xor U32709 (N_32709,N_31592,N_30099);
nand U32710 (N_32710,N_31686,N_30214);
or U32711 (N_32711,N_30389,N_30842);
or U32712 (N_32712,N_30459,N_30565);
and U32713 (N_32713,N_31619,N_31006);
and U32714 (N_32714,N_30988,N_30894);
or U32715 (N_32715,N_31853,N_30343);
xnor U32716 (N_32716,N_30735,N_30844);
nor U32717 (N_32717,N_30031,N_30291);
nand U32718 (N_32718,N_30787,N_30215);
nor U32719 (N_32719,N_31345,N_30495);
and U32720 (N_32720,N_30780,N_31563);
and U32721 (N_32721,N_30734,N_31462);
and U32722 (N_32722,N_31662,N_30329);
nand U32723 (N_32723,N_30970,N_31170);
nor U32724 (N_32724,N_31749,N_31902);
or U32725 (N_32725,N_31739,N_30810);
or U32726 (N_32726,N_30189,N_31227);
xor U32727 (N_32727,N_31043,N_30980);
or U32728 (N_32728,N_31492,N_31731);
nand U32729 (N_32729,N_31973,N_31199);
or U32730 (N_32730,N_31708,N_30159);
or U32731 (N_32731,N_31053,N_31613);
or U32732 (N_32732,N_30115,N_31936);
nand U32733 (N_32733,N_31869,N_30515);
and U32734 (N_32734,N_31917,N_31934);
xnor U32735 (N_32735,N_31772,N_31256);
or U32736 (N_32736,N_31919,N_30987);
nor U32737 (N_32737,N_31128,N_31210);
nor U32738 (N_32738,N_30996,N_31393);
and U32739 (N_32739,N_30936,N_31319);
xnor U32740 (N_32740,N_30680,N_30743);
and U32741 (N_32741,N_30344,N_30129);
nor U32742 (N_32742,N_30622,N_31643);
or U32743 (N_32743,N_30881,N_30307);
nor U32744 (N_32744,N_31241,N_31145);
nand U32745 (N_32745,N_30283,N_30065);
and U32746 (N_32746,N_30701,N_30967);
xnor U32747 (N_32747,N_31149,N_31183);
or U32748 (N_32748,N_30692,N_31985);
nand U32749 (N_32749,N_31184,N_31036);
and U32750 (N_32750,N_31900,N_30375);
nand U32751 (N_32751,N_30968,N_31761);
and U32752 (N_32752,N_31287,N_31746);
nor U32753 (N_32753,N_31855,N_30012);
xor U32754 (N_32754,N_30074,N_30444);
nor U32755 (N_32755,N_30157,N_30075);
or U32756 (N_32756,N_31532,N_31495);
nor U32757 (N_32757,N_30969,N_31074);
or U32758 (N_32758,N_31294,N_31530);
nor U32759 (N_32759,N_31282,N_30972);
nand U32760 (N_32760,N_31121,N_30531);
xnor U32761 (N_32761,N_30595,N_31727);
or U32762 (N_32762,N_31790,N_30973);
or U32763 (N_32763,N_31751,N_30978);
or U32764 (N_32764,N_31291,N_31878);
nor U32765 (N_32765,N_30101,N_30384);
or U32766 (N_32766,N_30934,N_31629);
xor U32767 (N_32767,N_30526,N_31528);
nor U32768 (N_32768,N_30039,N_30252);
xor U32769 (N_32769,N_30985,N_30579);
xor U32770 (N_32770,N_31784,N_30848);
nand U32771 (N_32771,N_30168,N_30490);
xor U32772 (N_32772,N_30397,N_31246);
or U32773 (N_32773,N_30164,N_31697);
nor U32774 (N_32774,N_31527,N_30991);
nand U32775 (N_32775,N_31946,N_30522);
nand U32776 (N_32776,N_30568,N_30091);
nand U32777 (N_32777,N_31135,N_30016);
or U32778 (N_32778,N_31373,N_30699);
nor U32779 (N_32779,N_30857,N_30400);
nand U32780 (N_32780,N_31750,N_30944);
nor U32781 (N_32781,N_31119,N_30385);
and U32782 (N_32782,N_30959,N_30149);
or U32783 (N_32783,N_30438,N_31452);
xor U32784 (N_32784,N_30941,N_30696);
and U32785 (N_32785,N_30006,N_31343);
and U32786 (N_32786,N_31890,N_30911);
nor U32787 (N_32787,N_31205,N_30922);
nand U32788 (N_32788,N_31910,N_31004);
xnor U32789 (N_32789,N_30413,N_31669);
or U32790 (N_32790,N_30742,N_30235);
and U32791 (N_32791,N_31617,N_30437);
nand U32792 (N_32792,N_30599,N_30048);
and U32793 (N_32793,N_30598,N_31167);
nand U32794 (N_32794,N_30601,N_31508);
xor U32795 (N_32795,N_31378,N_30382);
or U32796 (N_32796,N_31911,N_31076);
or U32797 (N_32797,N_31456,N_30320);
and U32798 (N_32798,N_30067,N_31969);
or U32799 (N_32799,N_30478,N_30606);
or U32800 (N_32800,N_31060,N_31918);
or U32801 (N_32801,N_31901,N_30194);
xor U32802 (N_32802,N_31132,N_31702);
nand U32803 (N_32803,N_31397,N_30632);
nor U32804 (N_32804,N_31963,N_31250);
xor U32805 (N_32805,N_31313,N_30492);
and U32806 (N_32806,N_30349,N_31673);
nor U32807 (N_32807,N_31417,N_31190);
or U32808 (N_32808,N_30371,N_31484);
nand U32809 (N_32809,N_31382,N_31606);
and U32810 (N_32810,N_31730,N_30918);
nor U32811 (N_32811,N_31860,N_30873);
xnor U32812 (N_32812,N_31831,N_30637);
xnor U32813 (N_32813,N_31096,N_31725);
xnor U32814 (N_32814,N_30381,N_30728);
xnor U32815 (N_32815,N_31762,N_31897);
and U32816 (N_32816,N_31344,N_30261);
nor U32817 (N_32817,N_31021,N_30158);
and U32818 (N_32818,N_30386,N_31844);
and U32819 (N_32819,N_30751,N_30274);
nand U32820 (N_32820,N_31771,N_30964);
and U32821 (N_32821,N_31952,N_30895);
nor U32822 (N_32822,N_30975,N_30313);
and U32823 (N_32823,N_31907,N_30299);
or U32824 (N_32824,N_31928,N_30602);
or U32825 (N_32825,N_31754,N_31481);
or U32826 (N_32826,N_30037,N_30631);
and U32827 (N_32827,N_30497,N_30575);
nand U32828 (N_32828,N_31654,N_31020);
or U32829 (N_32829,N_30325,N_30816);
xnor U32830 (N_32830,N_30491,N_30795);
and U32831 (N_32831,N_30306,N_30905);
and U32832 (N_32832,N_30367,N_30677);
nand U32833 (N_32833,N_31684,N_30026);
or U32834 (N_32834,N_31233,N_31086);
or U32835 (N_32835,N_31325,N_31716);
or U32836 (N_32836,N_30945,N_31430);
nand U32837 (N_32837,N_30015,N_30507);
and U32838 (N_32838,N_30366,N_31402);
nand U32839 (N_32839,N_31987,N_30524);
or U32840 (N_32840,N_31013,N_31788);
or U32841 (N_32841,N_30044,N_31409);
xnor U32842 (N_32842,N_31536,N_30448);
and U32843 (N_32843,N_31224,N_30865);
and U32844 (N_32844,N_31538,N_31464);
nor U32845 (N_32845,N_30082,N_31331);
and U32846 (N_32846,N_30682,N_30954);
or U32847 (N_32847,N_30392,N_30639);
and U32848 (N_32848,N_30538,N_30935);
or U32849 (N_32849,N_31857,N_31550);
or U32850 (N_32850,N_31954,N_30586);
nand U32851 (N_32851,N_31760,N_30484);
xor U32852 (N_32852,N_31868,N_30783);
and U32853 (N_32853,N_30051,N_31064);
nand U32854 (N_32854,N_30646,N_31296);
nor U32855 (N_32855,N_30782,N_30591);
and U32856 (N_32856,N_31117,N_30879);
nor U32857 (N_32857,N_30509,N_30312);
nor U32858 (N_32858,N_30445,N_31904);
xnor U32859 (N_32859,N_30485,N_30077);
nor U32860 (N_32860,N_30837,N_30589);
and U32861 (N_32861,N_30511,N_31770);
or U32862 (N_32862,N_31033,N_31473);
and U32863 (N_32863,N_30072,N_31295);
and U32864 (N_32864,N_30337,N_31392);
and U32865 (N_32865,N_30038,N_30452);
or U32866 (N_32866,N_30552,N_31482);
or U32867 (N_32867,N_31204,N_30981);
nand U32868 (N_32868,N_30958,N_31726);
nor U32869 (N_32869,N_31583,N_31466);
nor U32870 (N_32870,N_30520,N_31269);
nand U32871 (N_32871,N_31723,N_31032);
nand U32872 (N_32872,N_31913,N_30246);
xnor U32873 (N_32873,N_31010,N_30095);
and U32874 (N_32874,N_30940,N_31610);
or U32875 (N_32875,N_30281,N_30672);
xor U32876 (N_32876,N_31221,N_30417);
or U32877 (N_32877,N_31247,N_30020);
nand U32878 (N_32878,N_30352,N_31570);
and U32879 (N_32879,N_30153,N_31489);
nand U32880 (N_32880,N_31468,N_30201);
xnor U32881 (N_32881,N_30571,N_30262);
nor U32882 (N_32882,N_30221,N_31641);
nor U32883 (N_32883,N_31763,N_30587);
nand U32884 (N_32884,N_30813,N_30908);
nor U32885 (N_32885,N_31208,N_30029);
and U32886 (N_32886,N_31447,N_30019);
nand U32887 (N_32887,N_30953,N_31025);
or U32888 (N_32888,N_30912,N_31383);
nand U32889 (N_32889,N_31769,N_31799);
nor U32890 (N_32890,N_30592,N_31699);
xor U32891 (N_32891,N_30069,N_31648);
nor U32892 (N_32892,N_31835,N_31230);
and U32893 (N_32893,N_30995,N_30726);
nor U32894 (N_32894,N_31304,N_31312);
xor U32895 (N_32895,N_30018,N_31586);
xnor U32896 (N_32896,N_30698,N_30882);
nor U32897 (N_32897,N_30836,N_31414);
and U32898 (N_32898,N_30802,N_31507);
and U32899 (N_32899,N_31124,N_31621);
xnor U32900 (N_32900,N_31222,N_31992);
and U32901 (N_32901,N_30617,N_31817);
or U32902 (N_32902,N_31867,N_30118);
nor U32903 (N_32903,N_30423,N_30859);
xnor U32904 (N_32904,N_30427,N_31114);
xnor U32905 (N_32905,N_30706,N_31951);
xnor U32906 (N_32906,N_30054,N_30396);
or U32907 (N_32907,N_30897,N_31174);
and U32908 (N_32908,N_31865,N_31094);
nand U32909 (N_32909,N_30533,N_30931);
or U32910 (N_32910,N_31633,N_31428);
xnor U32911 (N_32911,N_31141,N_31198);
or U32912 (N_32912,N_31143,N_30927);
or U32913 (N_32913,N_30047,N_31108);
and U32914 (N_32914,N_30374,N_31066);
nor U32915 (N_32915,N_30993,N_31516);
or U32916 (N_32916,N_30380,N_31427);
nor U32917 (N_32917,N_30928,N_31766);
nand U32918 (N_32918,N_31363,N_31435);
nor U32919 (N_32919,N_30961,N_30419);
xor U32920 (N_32920,N_30718,N_30124);
or U32921 (N_32921,N_31404,N_30791);
and U32922 (N_32922,N_31334,N_31876);
or U32923 (N_32923,N_31719,N_31714);
xnor U32924 (N_32924,N_30022,N_31798);
and U32925 (N_32925,N_31131,N_30318);
nand U32926 (N_32926,N_31355,N_31232);
xor U32927 (N_32927,N_30302,N_31942);
xnor U32928 (N_32928,N_30210,N_30656);
nand U32929 (N_32929,N_31764,N_31213);
nand U32930 (N_32930,N_30573,N_30479);
xnor U32931 (N_32931,N_30370,N_30547);
and U32932 (N_32932,N_30847,N_31574);
or U32933 (N_32933,N_30739,N_31399);
or U32934 (N_32934,N_30078,N_31212);
xnor U32935 (N_32935,N_30574,N_31179);
or U32936 (N_32936,N_31966,N_30803);
nand U32937 (N_32937,N_31717,N_31651);
or U32938 (N_32938,N_31565,N_30821);
and U32939 (N_32939,N_30761,N_31103);
nand U32940 (N_32940,N_30764,N_30354);
or U32941 (N_32941,N_30649,N_31422);
or U32942 (N_32942,N_31400,N_31406);
nand U32943 (N_32943,N_30011,N_31413);
xor U32944 (N_32944,N_30683,N_30106);
xnor U32945 (N_32945,N_31207,N_31922);
and U32946 (N_32946,N_30535,N_30725);
nand U32947 (N_32947,N_31323,N_30869);
or U32948 (N_32948,N_30117,N_31286);
or U32949 (N_32949,N_31940,N_30216);
and U32950 (N_32950,N_30110,N_31394);
xnor U32951 (N_32951,N_30504,N_31567);
or U32952 (N_32952,N_31573,N_31941);
or U32953 (N_32953,N_31715,N_30556);
and U32954 (N_32954,N_30137,N_31937);
nand U32955 (N_32955,N_30835,N_30355);
nor U32956 (N_32956,N_31800,N_31407);
and U32957 (N_32957,N_31453,N_31848);
xnor U32958 (N_32958,N_31872,N_30710);
and U32959 (N_32959,N_31774,N_31551);
xor U32960 (N_32960,N_30155,N_31812);
or U32961 (N_32961,N_30630,N_30257);
or U32962 (N_32962,N_31644,N_31611);
or U32963 (N_32963,N_30282,N_31616);
or U32964 (N_32964,N_31683,N_30790);
xor U32965 (N_32965,N_31237,N_30581);
or U32966 (N_32966,N_30083,N_30823);
and U32967 (N_32967,N_30807,N_30792);
xnor U32968 (N_32968,N_30626,N_31624);
and U32969 (N_32969,N_31503,N_31561);
or U32970 (N_32970,N_31544,N_30899);
and U32971 (N_32971,N_30197,N_30196);
nand U32972 (N_32972,N_31471,N_31950);
nand U32973 (N_32973,N_31542,N_30749);
or U32974 (N_32974,N_30660,N_31929);
nand U32975 (N_32975,N_30933,N_31315);
or U32976 (N_32976,N_31419,N_31111);
xor U32977 (N_32977,N_31268,N_30360);
and U32978 (N_32978,N_30657,N_30154);
xnor U32979 (N_32979,N_30768,N_30736);
or U32980 (N_32980,N_30409,N_30866);
and U32981 (N_32981,N_31490,N_30493);
or U32982 (N_32982,N_30003,N_30647);
xnor U32983 (N_32983,N_31894,N_30551);
xor U32984 (N_32984,N_30259,N_31517);
and U32985 (N_32985,N_31322,N_30487);
and U32986 (N_32986,N_30990,N_30965);
nand U32987 (N_32987,N_30860,N_31163);
nor U32988 (N_32988,N_30921,N_30752);
nor U32989 (N_32989,N_30289,N_31601);
and U32990 (N_32990,N_30181,N_31755);
nor U32991 (N_32991,N_31443,N_30357);
nor U32992 (N_32992,N_30362,N_31347);
nor U32993 (N_32993,N_31380,N_31989);
nand U32994 (N_32994,N_30603,N_31665);
and U32995 (N_32995,N_30667,N_31321);
and U32996 (N_32996,N_30436,N_31444);
or U32997 (N_32997,N_31558,N_31097);
xnor U32998 (N_32998,N_30714,N_31217);
or U32999 (N_32999,N_30748,N_30962);
or U33000 (N_33000,N_31674,N_30744);
nand U33001 (N_33001,N_31623,N_30876);
xnor U33002 (N_33002,N_30710,N_31843);
xnor U33003 (N_33003,N_31654,N_31650);
xnor U33004 (N_33004,N_31519,N_30014);
xor U33005 (N_33005,N_30755,N_31634);
nand U33006 (N_33006,N_31518,N_31187);
nor U33007 (N_33007,N_31406,N_31850);
or U33008 (N_33008,N_30415,N_31042);
and U33009 (N_33009,N_31771,N_30587);
nand U33010 (N_33010,N_30547,N_30263);
or U33011 (N_33011,N_31751,N_30341);
or U33012 (N_33012,N_30406,N_31405);
or U33013 (N_33013,N_30534,N_30302);
nand U33014 (N_33014,N_30427,N_31813);
xnor U33015 (N_33015,N_31910,N_31044);
xnor U33016 (N_33016,N_31160,N_31425);
nor U33017 (N_33017,N_31404,N_31647);
nand U33018 (N_33018,N_30678,N_30785);
xnor U33019 (N_33019,N_31526,N_30095);
and U33020 (N_33020,N_30089,N_31378);
nor U33021 (N_33021,N_30153,N_30939);
nand U33022 (N_33022,N_30374,N_31129);
or U33023 (N_33023,N_30896,N_31520);
xor U33024 (N_33024,N_30194,N_30589);
xor U33025 (N_33025,N_30323,N_31359);
or U33026 (N_33026,N_30041,N_31444);
or U33027 (N_33027,N_31833,N_30557);
nand U33028 (N_33028,N_30362,N_30754);
xor U33029 (N_33029,N_31713,N_31264);
nor U33030 (N_33030,N_30219,N_31140);
nor U33031 (N_33031,N_30764,N_30190);
xor U33032 (N_33032,N_30762,N_30979);
xnor U33033 (N_33033,N_31972,N_30731);
or U33034 (N_33034,N_31418,N_31407);
nand U33035 (N_33035,N_30379,N_31585);
xor U33036 (N_33036,N_30516,N_31104);
xnor U33037 (N_33037,N_30613,N_30619);
or U33038 (N_33038,N_30525,N_31713);
or U33039 (N_33039,N_31914,N_31078);
xnor U33040 (N_33040,N_31417,N_30674);
nor U33041 (N_33041,N_30091,N_31939);
and U33042 (N_33042,N_30488,N_31286);
and U33043 (N_33043,N_31581,N_31116);
nand U33044 (N_33044,N_30004,N_31550);
nand U33045 (N_33045,N_31137,N_31603);
xnor U33046 (N_33046,N_30344,N_30777);
nor U33047 (N_33047,N_31785,N_31467);
nor U33048 (N_33048,N_31746,N_30562);
xor U33049 (N_33049,N_30766,N_30472);
or U33050 (N_33050,N_31564,N_31130);
or U33051 (N_33051,N_31198,N_31785);
xor U33052 (N_33052,N_30003,N_31362);
nor U33053 (N_33053,N_30313,N_30530);
and U33054 (N_33054,N_30825,N_30399);
nand U33055 (N_33055,N_30064,N_31607);
or U33056 (N_33056,N_31680,N_31861);
nor U33057 (N_33057,N_30911,N_30031);
or U33058 (N_33058,N_31211,N_30819);
xnor U33059 (N_33059,N_30853,N_30560);
and U33060 (N_33060,N_31566,N_31121);
or U33061 (N_33061,N_30060,N_30267);
nand U33062 (N_33062,N_31949,N_30710);
or U33063 (N_33063,N_31667,N_30659);
and U33064 (N_33064,N_31924,N_31712);
and U33065 (N_33065,N_31353,N_30169);
or U33066 (N_33066,N_30161,N_31793);
and U33067 (N_33067,N_31495,N_31235);
nand U33068 (N_33068,N_30381,N_31821);
nor U33069 (N_33069,N_30855,N_31407);
and U33070 (N_33070,N_30523,N_31526);
and U33071 (N_33071,N_31078,N_31381);
nand U33072 (N_33072,N_30636,N_30950);
and U33073 (N_33073,N_31134,N_31831);
xor U33074 (N_33074,N_30547,N_30977);
nor U33075 (N_33075,N_30481,N_30035);
xnor U33076 (N_33076,N_30570,N_30959);
xor U33077 (N_33077,N_30709,N_30740);
and U33078 (N_33078,N_31644,N_31678);
xor U33079 (N_33079,N_30569,N_31053);
nor U33080 (N_33080,N_30034,N_30064);
and U33081 (N_33081,N_30782,N_31630);
nand U33082 (N_33082,N_31403,N_30593);
nor U33083 (N_33083,N_30601,N_30543);
xor U33084 (N_33084,N_31906,N_31237);
or U33085 (N_33085,N_31060,N_31078);
nand U33086 (N_33086,N_30890,N_30184);
xnor U33087 (N_33087,N_30497,N_31065);
nor U33088 (N_33088,N_30540,N_30960);
xnor U33089 (N_33089,N_30378,N_31256);
or U33090 (N_33090,N_31829,N_30631);
xor U33091 (N_33091,N_31522,N_30742);
xor U33092 (N_33092,N_30598,N_30813);
nand U33093 (N_33093,N_31539,N_30758);
nand U33094 (N_33094,N_31480,N_30865);
or U33095 (N_33095,N_30357,N_31782);
nor U33096 (N_33096,N_30071,N_30117);
xnor U33097 (N_33097,N_30740,N_31929);
nor U33098 (N_33098,N_30672,N_30980);
and U33099 (N_33099,N_30534,N_30818);
nand U33100 (N_33100,N_30568,N_30556);
and U33101 (N_33101,N_30228,N_30998);
and U33102 (N_33102,N_30780,N_31343);
nand U33103 (N_33103,N_31653,N_31398);
nand U33104 (N_33104,N_31053,N_30924);
or U33105 (N_33105,N_30473,N_31465);
or U33106 (N_33106,N_31928,N_30577);
nand U33107 (N_33107,N_31663,N_30464);
xnor U33108 (N_33108,N_31601,N_31618);
xnor U33109 (N_33109,N_30300,N_31280);
nor U33110 (N_33110,N_30248,N_30524);
or U33111 (N_33111,N_31349,N_31516);
xor U33112 (N_33112,N_31080,N_31144);
nand U33113 (N_33113,N_30059,N_31307);
or U33114 (N_33114,N_31896,N_31824);
nand U33115 (N_33115,N_31873,N_31946);
xor U33116 (N_33116,N_31397,N_30177);
nand U33117 (N_33117,N_30249,N_30281);
xor U33118 (N_33118,N_30200,N_31645);
or U33119 (N_33119,N_31561,N_31221);
nor U33120 (N_33120,N_31084,N_31230);
or U33121 (N_33121,N_30963,N_31858);
nand U33122 (N_33122,N_30100,N_30844);
or U33123 (N_33123,N_30024,N_30823);
or U33124 (N_33124,N_30286,N_30278);
or U33125 (N_33125,N_31966,N_30447);
xnor U33126 (N_33126,N_30879,N_30769);
or U33127 (N_33127,N_31322,N_31969);
xnor U33128 (N_33128,N_31191,N_31726);
or U33129 (N_33129,N_30569,N_30298);
nand U33130 (N_33130,N_31567,N_31507);
or U33131 (N_33131,N_31825,N_31637);
nor U33132 (N_33132,N_31064,N_31278);
or U33133 (N_33133,N_30789,N_30124);
and U33134 (N_33134,N_30930,N_30097);
xor U33135 (N_33135,N_31843,N_31221);
xnor U33136 (N_33136,N_30497,N_30523);
nand U33137 (N_33137,N_31874,N_30229);
xor U33138 (N_33138,N_30967,N_30855);
or U33139 (N_33139,N_31905,N_30848);
and U33140 (N_33140,N_31018,N_31573);
and U33141 (N_33141,N_31233,N_31977);
nor U33142 (N_33142,N_30687,N_31836);
and U33143 (N_33143,N_30357,N_31518);
or U33144 (N_33144,N_30127,N_30729);
xnor U33145 (N_33145,N_30485,N_30060);
xnor U33146 (N_33146,N_30723,N_30534);
xor U33147 (N_33147,N_31914,N_31911);
and U33148 (N_33148,N_31575,N_31750);
and U33149 (N_33149,N_30328,N_30973);
xnor U33150 (N_33150,N_31179,N_31030);
xor U33151 (N_33151,N_30089,N_30341);
or U33152 (N_33152,N_30647,N_30491);
nand U33153 (N_33153,N_30023,N_31898);
or U33154 (N_33154,N_31263,N_31476);
nor U33155 (N_33155,N_30170,N_30809);
xor U33156 (N_33156,N_30892,N_30161);
xnor U33157 (N_33157,N_31265,N_30368);
or U33158 (N_33158,N_30707,N_31115);
or U33159 (N_33159,N_31407,N_31082);
and U33160 (N_33160,N_31944,N_30387);
and U33161 (N_33161,N_30883,N_30412);
nand U33162 (N_33162,N_30929,N_30236);
nand U33163 (N_33163,N_30202,N_31135);
nand U33164 (N_33164,N_31794,N_31224);
and U33165 (N_33165,N_30434,N_30922);
and U33166 (N_33166,N_31225,N_30886);
and U33167 (N_33167,N_31988,N_30364);
xor U33168 (N_33168,N_31868,N_31390);
nand U33169 (N_33169,N_31886,N_30015);
or U33170 (N_33170,N_30958,N_30757);
or U33171 (N_33171,N_31394,N_30654);
xnor U33172 (N_33172,N_31480,N_31958);
nor U33173 (N_33173,N_31034,N_31079);
xnor U33174 (N_33174,N_31508,N_30344);
and U33175 (N_33175,N_31707,N_30948);
nand U33176 (N_33176,N_31046,N_30142);
nand U33177 (N_33177,N_30168,N_31313);
or U33178 (N_33178,N_31459,N_30162);
nand U33179 (N_33179,N_31933,N_30592);
nand U33180 (N_33180,N_30095,N_31395);
and U33181 (N_33181,N_31101,N_30141);
or U33182 (N_33182,N_31822,N_31799);
nand U33183 (N_33183,N_31333,N_30735);
xnor U33184 (N_33184,N_30168,N_31295);
nand U33185 (N_33185,N_30619,N_30251);
xor U33186 (N_33186,N_30184,N_30392);
and U33187 (N_33187,N_31946,N_30470);
or U33188 (N_33188,N_30855,N_31756);
nor U33189 (N_33189,N_30250,N_31002);
and U33190 (N_33190,N_31836,N_31172);
and U33191 (N_33191,N_30690,N_30693);
or U33192 (N_33192,N_31708,N_31962);
nand U33193 (N_33193,N_31458,N_31757);
nand U33194 (N_33194,N_31496,N_30092);
and U33195 (N_33195,N_31780,N_31193);
nand U33196 (N_33196,N_30425,N_30492);
nor U33197 (N_33197,N_31744,N_30236);
or U33198 (N_33198,N_30469,N_30654);
xnor U33199 (N_33199,N_30097,N_30078);
nand U33200 (N_33200,N_30343,N_31488);
nor U33201 (N_33201,N_31601,N_31578);
or U33202 (N_33202,N_30525,N_30420);
xor U33203 (N_33203,N_30368,N_31967);
and U33204 (N_33204,N_30567,N_31933);
and U33205 (N_33205,N_31234,N_30306);
xor U33206 (N_33206,N_31985,N_31852);
or U33207 (N_33207,N_31852,N_31074);
nor U33208 (N_33208,N_31883,N_30508);
nor U33209 (N_33209,N_31113,N_30431);
xnor U33210 (N_33210,N_30746,N_31843);
and U33211 (N_33211,N_31213,N_31030);
nand U33212 (N_33212,N_30100,N_30886);
nor U33213 (N_33213,N_30622,N_31374);
xor U33214 (N_33214,N_30913,N_31535);
xnor U33215 (N_33215,N_31150,N_31026);
nor U33216 (N_33216,N_31092,N_30837);
or U33217 (N_33217,N_31246,N_31786);
or U33218 (N_33218,N_30742,N_30963);
nor U33219 (N_33219,N_31827,N_31957);
or U33220 (N_33220,N_31189,N_30465);
and U33221 (N_33221,N_30948,N_30960);
nand U33222 (N_33222,N_30545,N_31041);
or U33223 (N_33223,N_30047,N_30744);
nor U33224 (N_33224,N_30164,N_30425);
nand U33225 (N_33225,N_31640,N_31575);
nor U33226 (N_33226,N_31552,N_31102);
nand U33227 (N_33227,N_31026,N_31884);
nand U33228 (N_33228,N_31782,N_30630);
or U33229 (N_33229,N_30885,N_31969);
nor U33230 (N_33230,N_30919,N_30864);
nor U33231 (N_33231,N_31675,N_31216);
xnor U33232 (N_33232,N_30817,N_31942);
and U33233 (N_33233,N_31422,N_31705);
nand U33234 (N_33234,N_31706,N_31109);
xor U33235 (N_33235,N_30763,N_31846);
and U33236 (N_33236,N_30545,N_30907);
nor U33237 (N_33237,N_30286,N_31666);
xor U33238 (N_33238,N_31877,N_31251);
nand U33239 (N_33239,N_30323,N_31087);
and U33240 (N_33240,N_31940,N_31833);
nor U33241 (N_33241,N_30758,N_30823);
xor U33242 (N_33242,N_31332,N_31815);
nand U33243 (N_33243,N_31488,N_30049);
nand U33244 (N_33244,N_30094,N_30154);
nand U33245 (N_33245,N_30052,N_30119);
nor U33246 (N_33246,N_30052,N_31131);
and U33247 (N_33247,N_31316,N_30551);
or U33248 (N_33248,N_31002,N_31370);
and U33249 (N_33249,N_31976,N_30006);
nor U33250 (N_33250,N_30125,N_30397);
nor U33251 (N_33251,N_31208,N_31023);
nor U33252 (N_33252,N_30743,N_30301);
nor U33253 (N_33253,N_30859,N_31458);
nor U33254 (N_33254,N_30369,N_31614);
nand U33255 (N_33255,N_31755,N_30871);
nor U33256 (N_33256,N_30124,N_31686);
or U33257 (N_33257,N_31678,N_31129);
or U33258 (N_33258,N_30096,N_30630);
or U33259 (N_33259,N_31163,N_30234);
nand U33260 (N_33260,N_30133,N_30441);
nand U33261 (N_33261,N_30003,N_30831);
nand U33262 (N_33262,N_30377,N_30944);
and U33263 (N_33263,N_30623,N_31972);
nor U33264 (N_33264,N_30070,N_31452);
nand U33265 (N_33265,N_31315,N_30298);
xnor U33266 (N_33266,N_30180,N_31749);
nand U33267 (N_33267,N_30247,N_31651);
xor U33268 (N_33268,N_30229,N_31352);
nand U33269 (N_33269,N_31387,N_30466);
nand U33270 (N_33270,N_30253,N_30916);
and U33271 (N_33271,N_30857,N_30251);
and U33272 (N_33272,N_31551,N_30165);
nand U33273 (N_33273,N_31891,N_30371);
nand U33274 (N_33274,N_30220,N_30893);
xor U33275 (N_33275,N_31673,N_30451);
xor U33276 (N_33276,N_30818,N_30011);
nand U33277 (N_33277,N_30491,N_31921);
or U33278 (N_33278,N_30680,N_31228);
xor U33279 (N_33279,N_31438,N_30329);
or U33280 (N_33280,N_30714,N_31142);
and U33281 (N_33281,N_31529,N_30310);
and U33282 (N_33282,N_30514,N_30108);
xnor U33283 (N_33283,N_31140,N_30909);
xnor U33284 (N_33284,N_30667,N_30991);
and U33285 (N_33285,N_31723,N_31845);
nand U33286 (N_33286,N_31402,N_30664);
nor U33287 (N_33287,N_30254,N_30154);
nand U33288 (N_33288,N_30013,N_30868);
and U33289 (N_33289,N_31565,N_31373);
nand U33290 (N_33290,N_30809,N_31040);
xor U33291 (N_33291,N_31873,N_31556);
nand U33292 (N_33292,N_31380,N_31977);
xor U33293 (N_33293,N_31472,N_30058);
nor U33294 (N_33294,N_31218,N_30157);
nand U33295 (N_33295,N_30240,N_30929);
xnor U33296 (N_33296,N_30808,N_30579);
nor U33297 (N_33297,N_30537,N_31699);
xor U33298 (N_33298,N_31170,N_31777);
and U33299 (N_33299,N_30898,N_30526);
nor U33300 (N_33300,N_31787,N_30137);
xor U33301 (N_33301,N_30383,N_31374);
xor U33302 (N_33302,N_31405,N_30204);
xor U33303 (N_33303,N_31908,N_30938);
and U33304 (N_33304,N_30269,N_31618);
nand U33305 (N_33305,N_31107,N_31153);
nor U33306 (N_33306,N_31452,N_31928);
nand U33307 (N_33307,N_31836,N_31342);
or U33308 (N_33308,N_31145,N_31262);
and U33309 (N_33309,N_30071,N_30081);
or U33310 (N_33310,N_31913,N_30249);
and U33311 (N_33311,N_30791,N_31935);
and U33312 (N_33312,N_30402,N_30911);
nor U33313 (N_33313,N_30551,N_31765);
nand U33314 (N_33314,N_30353,N_30545);
nand U33315 (N_33315,N_31690,N_30227);
nand U33316 (N_33316,N_30722,N_31988);
and U33317 (N_33317,N_30134,N_30020);
or U33318 (N_33318,N_31366,N_30274);
or U33319 (N_33319,N_30691,N_30851);
xor U33320 (N_33320,N_30469,N_30834);
nand U33321 (N_33321,N_30114,N_31401);
nor U33322 (N_33322,N_30383,N_30430);
nor U33323 (N_33323,N_30614,N_30406);
xnor U33324 (N_33324,N_30842,N_31819);
or U33325 (N_33325,N_30025,N_31370);
or U33326 (N_33326,N_31649,N_31390);
or U33327 (N_33327,N_31248,N_30888);
xor U33328 (N_33328,N_31504,N_31062);
or U33329 (N_33329,N_30503,N_31718);
nor U33330 (N_33330,N_30337,N_30794);
or U33331 (N_33331,N_31949,N_30608);
nand U33332 (N_33332,N_31403,N_31477);
or U33333 (N_33333,N_30360,N_31424);
xor U33334 (N_33334,N_31363,N_30904);
nor U33335 (N_33335,N_30139,N_30166);
nand U33336 (N_33336,N_31124,N_31724);
nor U33337 (N_33337,N_31504,N_30868);
nor U33338 (N_33338,N_31258,N_30462);
nor U33339 (N_33339,N_30653,N_31672);
and U33340 (N_33340,N_31453,N_31966);
and U33341 (N_33341,N_31768,N_31756);
nand U33342 (N_33342,N_31974,N_30433);
or U33343 (N_33343,N_31961,N_31508);
nor U33344 (N_33344,N_31867,N_31316);
nor U33345 (N_33345,N_30023,N_31583);
and U33346 (N_33346,N_31417,N_31022);
xnor U33347 (N_33347,N_30642,N_30388);
or U33348 (N_33348,N_31757,N_30669);
and U33349 (N_33349,N_30993,N_31400);
xnor U33350 (N_33350,N_30041,N_30721);
or U33351 (N_33351,N_30242,N_31536);
and U33352 (N_33352,N_31721,N_31545);
xor U33353 (N_33353,N_30495,N_31733);
xor U33354 (N_33354,N_30873,N_31651);
nand U33355 (N_33355,N_31696,N_30940);
xor U33356 (N_33356,N_31854,N_30139);
or U33357 (N_33357,N_31014,N_30631);
nor U33358 (N_33358,N_31502,N_30808);
and U33359 (N_33359,N_30889,N_31771);
nand U33360 (N_33360,N_31461,N_31998);
nor U33361 (N_33361,N_31652,N_31230);
or U33362 (N_33362,N_31997,N_30026);
and U33363 (N_33363,N_31373,N_30657);
nand U33364 (N_33364,N_30676,N_30277);
nand U33365 (N_33365,N_31206,N_30846);
and U33366 (N_33366,N_30355,N_31023);
xnor U33367 (N_33367,N_30756,N_31376);
and U33368 (N_33368,N_31747,N_31144);
xor U33369 (N_33369,N_31571,N_31907);
nor U33370 (N_33370,N_30813,N_31876);
nand U33371 (N_33371,N_30425,N_30750);
or U33372 (N_33372,N_31310,N_30266);
nand U33373 (N_33373,N_31402,N_31327);
or U33374 (N_33374,N_30776,N_31840);
or U33375 (N_33375,N_30461,N_30474);
or U33376 (N_33376,N_31418,N_31218);
nor U33377 (N_33377,N_31154,N_30060);
and U33378 (N_33378,N_30197,N_30831);
nand U33379 (N_33379,N_31756,N_30791);
nand U33380 (N_33380,N_31937,N_31800);
nor U33381 (N_33381,N_30568,N_31671);
and U33382 (N_33382,N_31597,N_31728);
and U33383 (N_33383,N_31985,N_30056);
and U33384 (N_33384,N_30366,N_31425);
nor U33385 (N_33385,N_30993,N_31306);
nand U33386 (N_33386,N_30178,N_31908);
nand U33387 (N_33387,N_31159,N_31482);
nor U33388 (N_33388,N_31249,N_30679);
or U33389 (N_33389,N_31756,N_30340);
or U33390 (N_33390,N_31029,N_30870);
xnor U33391 (N_33391,N_30591,N_30831);
and U33392 (N_33392,N_31099,N_31012);
nor U33393 (N_33393,N_31542,N_30931);
or U33394 (N_33394,N_31772,N_30235);
nor U33395 (N_33395,N_30927,N_30652);
nor U33396 (N_33396,N_30445,N_31889);
or U33397 (N_33397,N_31583,N_31527);
nand U33398 (N_33398,N_30891,N_31652);
or U33399 (N_33399,N_31816,N_30288);
and U33400 (N_33400,N_30007,N_31374);
nor U33401 (N_33401,N_31992,N_30201);
nor U33402 (N_33402,N_30278,N_30549);
nand U33403 (N_33403,N_31243,N_30423);
nor U33404 (N_33404,N_30928,N_30872);
xnor U33405 (N_33405,N_30250,N_30968);
and U33406 (N_33406,N_31058,N_31955);
xor U33407 (N_33407,N_30827,N_31759);
nand U33408 (N_33408,N_30579,N_31672);
xnor U33409 (N_33409,N_31384,N_30410);
or U33410 (N_33410,N_30395,N_30767);
and U33411 (N_33411,N_31604,N_30827);
nor U33412 (N_33412,N_31169,N_30662);
nor U33413 (N_33413,N_31444,N_31406);
xnor U33414 (N_33414,N_30340,N_30451);
xor U33415 (N_33415,N_31974,N_31775);
or U33416 (N_33416,N_31101,N_31669);
nor U33417 (N_33417,N_30886,N_30897);
xnor U33418 (N_33418,N_30504,N_31267);
xor U33419 (N_33419,N_31139,N_30362);
or U33420 (N_33420,N_30551,N_31347);
and U33421 (N_33421,N_31305,N_31864);
nor U33422 (N_33422,N_30825,N_30129);
and U33423 (N_33423,N_30458,N_31614);
nor U33424 (N_33424,N_30545,N_30888);
nand U33425 (N_33425,N_30169,N_30923);
xnor U33426 (N_33426,N_31787,N_30399);
xnor U33427 (N_33427,N_31847,N_31879);
or U33428 (N_33428,N_30225,N_31793);
nand U33429 (N_33429,N_31777,N_30839);
or U33430 (N_33430,N_31784,N_30469);
and U33431 (N_33431,N_30601,N_31149);
nand U33432 (N_33432,N_31115,N_30857);
and U33433 (N_33433,N_30059,N_30759);
and U33434 (N_33434,N_31531,N_31298);
xor U33435 (N_33435,N_31460,N_31935);
nand U33436 (N_33436,N_31746,N_31425);
nor U33437 (N_33437,N_31449,N_31200);
nor U33438 (N_33438,N_31845,N_31499);
nor U33439 (N_33439,N_30719,N_30580);
nand U33440 (N_33440,N_30063,N_31733);
or U33441 (N_33441,N_31663,N_31285);
nor U33442 (N_33442,N_31900,N_31518);
nand U33443 (N_33443,N_31637,N_31079);
or U33444 (N_33444,N_31898,N_31894);
or U33445 (N_33445,N_30879,N_30978);
nand U33446 (N_33446,N_30283,N_31642);
and U33447 (N_33447,N_31068,N_30608);
xnor U33448 (N_33448,N_31366,N_30003);
nor U33449 (N_33449,N_31637,N_30161);
and U33450 (N_33450,N_31296,N_31333);
nand U33451 (N_33451,N_31821,N_31674);
nand U33452 (N_33452,N_31899,N_30977);
nand U33453 (N_33453,N_31758,N_30215);
nor U33454 (N_33454,N_30838,N_31562);
and U33455 (N_33455,N_31745,N_31301);
xnor U33456 (N_33456,N_31956,N_31380);
or U33457 (N_33457,N_30900,N_31069);
and U33458 (N_33458,N_30533,N_30552);
xor U33459 (N_33459,N_30313,N_31513);
or U33460 (N_33460,N_31322,N_31480);
or U33461 (N_33461,N_31591,N_30880);
xor U33462 (N_33462,N_31698,N_31339);
and U33463 (N_33463,N_30349,N_31896);
xnor U33464 (N_33464,N_30925,N_31654);
and U33465 (N_33465,N_30857,N_31794);
nand U33466 (N_33466,N_30943,N_30231);
or U33467 (N_33467,N_31220,N_31335);
or U33468 (N_33468,N_30835,N_31648);
nor U33469 (N_33469,N_31466,N_31054);
or U33470 (N_33470,N_31823,N_31925);
and U33471 (N_33471,N_31222,N_30108);
xnor U33472 (N_33472,N_30431,N_31276);
nor U33473 (N_33473,N_30721,N_30161);
and U33474 (N_33474,N_30594,N_30985);
or U33475 (N_33475,N_30423,N_31928);
and U33476 (N_33476,N_31272,N_30169);
and U33477 (N_33477,N_30293,N_30354);
or U33478 (N_33478,N_30441,N_31513);
or U33479 (N_33479,N_31056,N_31338);
and U33480 (N_33480,N_31326,N_30717);
nor U33481 (N_33481,N_30050,N_31027);
xor U33482 (N_33482,N_31159,N_31399);
and U33483 (N_33483,N_31277,N_31238);
xnor U33484 (N_33484,N_31524,N_31489);
xnor U33485 (N_33485,N_30983,N_31595);
nor U33486 (N_33486,N_31882,N_30664);
nor U33487 (N_33487,N_31549,N_31668);
nor U33488 (N_33488,N_30508,N_31833);
or U33489 (N_33489,N_31225,N_31972);
xor U33490 (N_33490,N_31326,N_30498);
nand U33491 (N_33491,N_31656,N_31428);
nor U33492 (N_33492,N_31912,N_30605);
xnor U33493 (N_33493,N_30487,N_30744);
nor U33494 (N_33494,N_31743,N_31070);
nand U33495 (N_33495,N_31106,N_30940);
or U33496 (N_33496,N_30088,N_30112);
xor U33497 (N_33497,N_31754,N_30398);
or U33498 (N_33498,N_31090,N_31614);
and U33499 (N_33499,N_31286,N_31845);
and U33500 (N_33500,N_30310,N_31971);
nor U33501 (N_33501,N_31679,N_31422);
nor U33502 (N_33502,N_30830,N_30657);
nand U33503 (N_33503,N_30393,N_31641);
nand U33504 (N_33504,N_30142,N_31907);
nand U33505 (N_33505,N_31172,N_31213);
nand U33506 (N_33506,N_31735,N_31519);
or U33507 (N_33507,N_30595,N_31698);
nor U33508 (N_33508,N_31391,N_30985);
and U33509 (N_33509,N_30773,N_31450);
xor U33510 (N_33510,N_31223,N_31000);
nor U33511 (N_33511,N_30791,N_31836);
xor U33512 (N_33512,N_31860,N_30647);
xor U33513 (N_33513,N_31514,N_31615);
xor U33514 (N_33514,N_30710,N_30124);
or U33515 (N_33515,N_30664,N_30440);
or U33516 (N_33516,N_31800,N_31446);
xor U33517 (N_33517,N_31946,N_30007);
nor U33518 (N_33518,N_30812,N_31602);
and U33519 (N_33519,N_31510,N_31538);
xnor U33520 (N_33520,N_30348,N_30928);
xnor U33521 (N_33521,N_30316,N_31384);
nand U33522 (N_33522,N_30983,N_31463);
nand U33523 (N_33523,N_30918,N_30684);
xor U33524 (N_33524,N_30331,N_30017);
and U33525 (N_33525,N_30763,N_30694);
nor U33526 (N_33526,N_30398,N_30673);
nand U33527 (N_33527,N_30990,N_30038);
nand U33528 (N_33528,N_30451,N_30982);
nor U33529 (N_33529,N_30972,N_30045);
or U33530 (N_33530,N_30502,N_31557);
and U33531 (N_33531,N_31240,N_30129);
or U33532 (N_33532,N_31956,N_31742);
or U33533 (N_33533,N_31980,N_30322);
xor U33534 (N_33534,N_31585,N_30102);
nand U33535 (N_33535,N_30091,N_30616);
nand U33536 (N_33536,N_31141,N_31118);
and U33537 (N_33537,N_30363,N_31394);
or U33538 (N_33538,N_30677,N_31623);
nand U33539 (N_33539,N_31488,N_30491);
and U33540 (N_33540,N_31100,N_31660);
nor U33541 (N_33541,N_30864,N_30761);
xor U33542 (N_33542,N_31466,N_30650);
nor U33543 (N_33543,N_30484,N_31056);
xnor U33544 (N_33544,N_30464,N_31798);
and U33545 (N_33545,N_31726,N_31999);
nand U33546 (N_33546,N_31824,N_31754);
or U33547 (N_33547,N_31654,N_30513);
xor U33548 (N_33548,N_30940,N_30080);
nand U33549 (N_33549,N_31541,N_30507);
or U33550 (N_33550,N_30454,N_30445);
and U33551 (N_33551,N_31206,N_30331);
nand U33552 (N_33552,N_31204,N_30681);
and U33553 (N_33553,N_30154,N_30462);
xor U33554 (N_33554,N_30885,N_30424);
and U33555 (N_33555,N_30939,N_31870);
or U33556 (N_33556,N_30776,N_31336);
and U33557 (N_33557,N_30381,N_31150);
nor U33558 (N_33558,N_31289,N_30438);
or U33559 (N_33559,N_31776,N_30380);
and U33560 (N_33560,N_30745,N_30601);
xnor U33561 (N_33561,N_30215,N_30005);
or U33562 (N_33562,N_31171,N_30899);
nand U33563 (N_33563,N_31438,N_30366);
and U33564 (N_33564,N_31858,N_30398);
and U33565 (N_33565,N_30623,N_30791);
or U33566 (N_33566,N_31759,N_30399);
nor U33567 (N_33567,N_30163,N_30242);
nand U33568 (N_33568,N_30348,N_31434);
and U33569 (N_33569,N_30249,N_31159);
nor U33570 (N_33570,N_30429,N_31560);
and U33571 (N_33571,N_31457,N_31261);
nand U33572 (N_33572,N_31125,N_31956);
and U33573 (N_33573,N_31176,N_31179);
nand U33574 (N_33574,N_30722,N_30267);
nor U33575 (N_33575,N_31811,N_30605);
xnor U33576 (N_33576,N_30318,N_31505);
or U33577 (N_33577,N_30415,N_30742);
and U33578 (N_33578,N_30490,N_31360);
xor U33579 (N_33579,N_31845,N_30622);
nand U33580 (N_33580,N_30281,N_31316);
xnor U33581 (N_33581,N_30472,N_31604);
nand U33582 (N_33582,N_31925,N_31956);
nand U33583 (N_33583,N_30574,N_31677);
or U33584 (N_33584,N_30370,N_30556);
and U33585 (N_33585,N_30282,N_31975);
nor U33586 (N_33586,N_31671,N_31416);
or U33587 (N_33587,N_30270,N_31510);
nand U33588 (N_33588,N_31804,N_31002);
xor U33589 (N_33589,N_31417,N_31309);
xnor U33590 (N_33590,N_31853,N_31668);
and U33591 (N_33591,N_30689,N_31948);
and U33592 (N_33592,N_31462,N_31908);
nand U33593 (N_33593,N_30077,N_31927);
and U33594 (N_33594,N_30585,N_30271);
nor U33595 (N_33595,N_30198,N_31075);
nand U33596 (N_33596,N_30570,N_30345);
or U33597 (N_33597,N_31099,N_30617);
xor U33598 (N_33598,N_30455,N_31664);
and U33599 (N_33599,N_30549,N_30878);
nor U33600 (N_33600,N_31656,N_31014);
or U33601 (N_33601,N_31248,N_31857);
or U33602 (N_33602,N_31242,N_30820);
nor U33603 (N_33603,N_30971,N_30413);
and U33604 (N_33604,N_31382,N_31227);
nand U33605 (N_33605,N_31150,N_30600);
nand U33606 (N_33606,N_30592,N_30028);
nor U33607 (N_33607,N_31872,N_30153);
and U33608 (N_33608,N_31117,N_30893);
nand U33609 (N_33609,N_30072,N_31406);
or U33610 (N_33610,N_30593,N_31230);
xor U33611 (N_33611,N_31500,N_31787);
and U33612 (N_33612,N_31036,N_31406);
nor U33613 (N_33613,N_31720,N_30826);
and U33614 (N_33614,N_31817,N_31180);
and U33615 (N_33615,N_30853,N_31456);
nor U33616 (N_33616,N_31108,N_31066);
nand U33617 (N_33617,N_31304,N_31266);
nand U33618 (N_33618,N_30307,N_31691);
or U33619 (N_33619,N_30830,N_31656);
nor U33620 (N_33620,N_31846,N_31158);
nor U33621 (N_33621,N_31612,N_31087);
nor U33622 (N_33622,N_30811,N_30122);
xor U33623 (N_33623,N_31999,N_30532);
and U33624 (N_33624,N_30245,N_30166);
or U33625 (N_33625,N_30562,N_31827);
nand U33626 (N_33626,N_30434,N_31261);
nand U33627 (N_33627,N_30780,N_30785);
nor U33628 (N_33628,N_31483,N_31280);
nand U33629 (N_33629,N_30691,N_30267);
or U33630 (N_33630,N_30792,N_30512);
nor U33631 (N_33631,N_30931,N_30116);
or U33632 (N_33632,N_30194,N_30562);
and U33633 (N_33633,N_30950,N_30239);
xor U33634 (N_33634,N_31825,N_31355);
nand U33635 (N_33635,N_30805,N_31370);
and U33636 (N_33636,N_30240,N_30911);
nor U33637 (N_33637,N_30567,N_31934);
xnor U33638 (N_33638,N_30274,N_30240);
and U33639 (N_33639,N_31432,N_31841);
nor U33640 (N_33640,N_31541,N_31325);
and U33641 (N_33641,N_31140,N_30282);
or U33642 (N_33642,N_31009,N_31547);
nand U33643 (N_33643,N_30107,N_31961);
and U33644 (N_33644,N_30447,N_31055);
or U33645 (N_33645,N_31490,N_31191);
nor U33646 (N_33646,N_30749,N_30960);
and U33647 (N_33647,N_31493,N_30241);
nand U33648 (N_33648,N_30902,N_31150);
or U33649 (N_33649,N_31718,N_31001);
xor U33650 (N_33650,N_31655,N_31859);
nor U33651 (N_33651,N_30527,N_31880);
and U33652 (N_33652,N_30370,N_30884);
or U33653 (N_33653,N_31375,N_31614);
and U33654 (N_33654,N_31059,N_31581);
xnor U33655 (N_33655,N_30078,N_30835);
and U33656 (N_33656,N_31212,N_30410);
and U33657 (N_33657,N_30985,N_31397);
and U33658 (N_33658,N_31948,N_30890);
or U33659 (N_33659,N_30293,N_31537);
xnor U33660 (N_33660,N_30063,N_31710);
or U33661 (N_33661,N_31818,N_31263);
or U33662 (N_33662,N_31867,N_30857);
and U33663 (N_33663,N_31915,N_31129);
or U33664 (N_33664,N_30151,N_31030);
or U33665 (N_33665,N_31338,N_30651);
nand U33666 (N_33666,N_31326,N_30519);
and U33667 (N_33667,N_31661,N_31360);
nor U33668 (N_33668,N_30483,N_31744);
xor U33669 (N_33669,N_31466,N_31662);
xnor U33670 (N_33670,N_31630,N_30111);
nor U33671 (N_33671,N_31051,N_30555);
and U33672 (N_33672,N_31249,N_31213);
nor U33673 (N_33673,N_31595,N_30694);
or U33674 (N_33674,N_31001,N_31012);
xnor U33675 (N_33675,N_31621,N_31078);
or U33676 (N_33676,N_30703,N_30259);
nor U33677 (N_33677,N_30613,N_30056);
and U33678 (N_33678,N_31780,N_30877);
or U33679 (N_33679,N_31334,N_30189);
nand U33680 (N_33680,N_30137,N_30626);
or U33681 (N_33681,N_30684,N_30913);
and U33682 (N_33682,N_30086,N_30480);
xor U33683 (N_33683,N_30485,N_31734);
and U33684 (N_33684,N_31486,N_31538);
nor U33685 (N_33685,N_31124,N_30898);
xnor U33686 (N_33686,N_31445,N_30248);
nand U33687 (N_33687,N_31509,N_31608);
or U33688 (N_33688,N_30090,N_31032);
or U33689 (N_33689,N_30752,N_31399);
and U33690 (N_33690,N_31937,N_31256);
or U33691 (N_33691,N_30654,N_31260);
nand U33692 (N_33692,N_30388,N_31339);
and U33693 (N_33693,N_31171,N_30981);
nand U33694 (N_33694,N_31785,N_31157);
and U33695 (N_33695,N_30946,N_31195);
and U33696 (N_33696,N_30255,N_30202);
nand U33697 (N_33697,N_30301,N_31798);
nand U33698 (N_33698,N_30608,N_31630);
or U33699 (N_33699,N_31571,N_31781);
or U33700 (N_33700,N_31129,N_30141);
xnor U33701 (N_33701,N_31503,N_31490);
xor U33702 (N_33702,N_30066,N_30494);
nor U33703 (N_33703,N_31542,N_31128);
and U33704 (N_33704,N_31483,N_31821);
and U33705 (N_33705,N_30975,N_31847);
nand U33706 (N_33706,N_31358,N_31003);
nor U33707 (N_33707,N_31545,N_30925);
nand U33708 (N_33708,N_30046,N_31970);
or U33709 (N_33709,N_30979,N_30567);
nand U33710 (N_33710,N_30927,N_30232);
or U33711 (N_33711,N_30694,N_31613);
nor U33712 (N_33712,N_30428,N_31924);
nand U33713 (N_33713,N_31298,N_31190);
or U33714 (N_33714,N_30228,N_31132);
nand U33715 (N_33715,N_30981,N_31374);
or U33716 (N_33716,N_31581,N_31901);
or U33717 (N_33717,N_31905,N_31674);
nand U33718 (N_33718,N_30963,N_30119);
nand U33719 (N_33719,N_30503,N_30475);
xor U33720 (N_33720,N_31101,N_30658);
and U33721 (N_33721,N_31653,N_31340);
xnor U33722 (N_33722,N_30303,N_30628);
nor U33723 (N_33723,N_31354,N_31883);
nand U33724 (N_33724,N_30657,N_30988);
xor U33725 (N_33725,N_30532,N_30639);
and U33726 (N_33726,N_31642,N_30009);
or U33727 (N_33727,N_31230,N_30835);
nand U33728 (N_33728,N_30374,N_30590);
xor U33729 (N_33729,N_30010,N_30448);
and U33730 (N_33730,N_31254,N_31689);
or U33731 (N_33731,N_31710,N_31113);
xor U33732 (N_33732,N_31083,N_31717);
xor U33733 (N_33733,N_31268,N_31630);
nand U33734 (N_33734,N_31070,N_30803);
and U33735 (N_33735,N_31753,N_31431);
nor U33736 (N_33736,N_30310,N_31015);
nor U33737 (N_33737,N_31623,N_30909);
nand U33738 (N_33738,N_31460,N_31261);
nand U33739 (N_33739,N_31823,N_30946);
or U33740 (N_33740,N_30230,N_31821);
or U33741 (N_33741,N_30856,N_30807);
or U33742 (N_33742,N_30999,N_31649);
xor U33743 (N_33743,N_30909,N_31899);
and U33744 (N_33744,N_30645,N_30373);
nor U33745 (N_33745,N_30085,N_30730);
nand U33746 (N_33746,N_31130,N_31220);
nand U33747 (N_33747,N_31493,N_31641);
xnor U33748 (N_33748,N_30356,N_30353);
nand U33749 (N_33749,N_30533,N_31872);
nor U33750 (N_33750,N_30756,N_30926);
xor U33751 (N_33751,N_30121,N_31911);
or U33752 (N_33752,N_31954,N_31668);
nor U33753 (N_33753,N_31044,N_30635);
nor U33754 (N_33754,N_30901,N_31606);
nand U33755 (N_33755,N_31982,N_31949);
nand U33756 (N_33756,N_30708,N_30954);
nor U33757 (N_33757,N_30089,N_30186);
nor U33758 (N_33758,N_30772,N_30193);
or U33759 (N_33759,N_31917,N_30278);
nor U33760 (N_33760,N_31503,N_30077);
and U33761 (N_33761,N_31960,N_31286);
or U33762 (N_33762,N_31457,N_30391);
or U33763 (N_33763,N_31226,N_30398);
and U33764 (N_33764,N_30028,N_30603);
xnor U33765 (N_33765,N_30526,N_30268);
xor U33766 (N_33766,N_30231,N_31397);
and U33767 (N_33767,N_30228,N_30236);
or U33768 (N_33768,N_30606,N_31604);
nand U33769 (N_33769,N_31333,N_30893);
nor U33770 (N_33770,N_31323,N_30527);
nor U33771 (N_33771,N_30835,N_31973);
nor U33772 (N_33772,N_30620,N_31310);
and U33773 (N_33773,N_31342,N_31403);
or U33774 (N_33774,N_31345,N_30614);
xnor U33775 (N_33775,N_30465,N_31963);
nor U33776 (N_33776,N_31165,N_31285);
and U33777 (N_33777,N_30246,N_30748);
xor U33778 (N_33778,N_31609,N_30815);
or U33779 (N_33779,N_30744,N_30551);
xnor U33780 (N_33780,N_30963,N_31811);
or U33781 (N_33781,N_31204,N_30669);
xnor U33782 (N_33782,N_30676,N_30022);
xor U33783 (N_33783,N_31496,N_31642);
or U33784 (N_33784,N_31364,N_31224);
xor U33785 (N_33785,N_30733,N_31881);
and U33786 (N_33786,N_31127,N_31494);
nand U33787 (N_33787,N_30548,N_31102);
or U33788 (N_33788,N_31778,N_31522);
nand U33789 (N_33789,N_30651,N_30676);
nor U33790 (N_33790,N_31031,N_31124);
nand U33791 (N_33791,N_30856,N_31033);
nand U33792 (N_33792,N_30890,N_30746);
and U33793 (N_33793,N_31190,N_30623);
xor U33794 (N_33794,N_30669,N_31759);
or U33795 (N_33795,N_31142,N_31375);
and U33796 (N_33796,N_31938,N_31110);
nor U33797 (N_33797,N_31017,N_31258);
nand U33798 (N_33798,N_30333,N_31761);
nand U33799 (N_33799,N_30143,N_31055);
nand U33800 (N_33800,N_31652,N_31270);
and U33801 (N_33801,N_30271,N_31648);
or U33802 (N_33802,N_30954,N_30419);
nor U33803 (N_33803,N_31646,N_31322);
and U33804 (N_33804,N_30142,N_31656);
and U33805 (N_33805,N_31543,N_31179);
xnor U33806 (N_33806,N_31641,N_30277);
or U33807 (N_33807,N_30241,N_30137);
xor U33808 (N_33808,N_31065,N_30298);
nor U33809 (N_33809,N_30645,N_31911);
and U33810 (N_33810,N_31872,N_31574);
or U33811 (N_33811,N_30197,N_31837);
or U33812 (N_33812,N_30355,N_30566);
xnor U33813 (N_33813,N_30233,N_30114);
xor U33814 (N_33814,N_30568,N_30899);
and U33815 (N_33815,N_30300,N_31152);
nand U33816 (N_33816,N_31804,N_30884);
nand U33817 (N_33817,N_30695,N_30549);
nor U33818 (N_33818,N_31428,N_30547);
nor U33819 (N_33819,N_31463,N_30037);
or U33820 (N_33820,N_31114,N_30264);
or U33821 (N_33821,N_30246,N_30902);
nand U33822 (N_33822,N_31833,N_30332);
or U33823 (N_33823,N_30760,N_31337);
nand U33824 (N_33824,N_30402,N_31948);
nand U33825 (N_33825,N_31006,N_31897);
nand U33826 (N_33826,N_31991,N_31744);
or U33827 (N_33827,N_31951,N_31982);
and U33828 (N_33828,N_31149,N_31908);
nor U33829 (N_33829,N_31917,N_30593);
or U33830 (N_33830,N_31108,N_30267);
nor U33831 (N_33831,N_30346,N_31338);
nor U33832 (N_33832,N_31819,N_31681);
nand U33833 (N_33833,N_30268,N_31524);
and U33834 (N_33834,N_30067,N_31275);
and U33835 (N_33835,N_30568,N_30079);
nand U33836 (N_33836,N_30514,N_31062);
nor U33837 (N_33837,N_30272,N_30647);
and U33838 (N_33838,N_30339,N_31645);
nand U33839 (N_33839,N_31300,N_31514);
nand U33840 (N_33840,N_31010,N_30473);
and U33841 (N_33841,N_30923,N_30391);
nor U33842 (N_33842,N_31638,N_30447);
and U33843 (N_33843,N_31667,N_31155);
and U33844 (N_33844,N_31429,N_31135);
or U33845 (N_33845,N_30020,N_30958);
nand U33846 (N_33846,N_31966,N_31139);
nor U33847 (N_33847,N_30283,N_30976);
and U33848 (N_33848,N_31439,N_31619);
nand U33849 (N_33849,N_30346,N_30570);
xnor U33850 (N_33850,N_30105,N_31281);
and U33851 (N_33851,N_31499,N_30309);
or U33852 (N_33852,N_31066,N_31804);
nand U33853 (N_33853,N_30444,N_30196);
or U33854 (N_33854,N_30796,N_30958);
xor U33855 (N_33855,N_30366,N_31443);
nand U33856 (N_33856,N_30786,N_30527);
nor U33857 (N_33857,N_31731,N_30122);
and U33858 (N_33858,N_30009,N_31594);
or U33859 (N_33859,N_31011,N_30828);
and U33860 (N_33860,N_31206,N_31084);
nand U33861 (N_33861,N_30182,N_31814);
nor U33862 (N_33862,N_30933,N_30610);
nand U33863 (N_33863,N_30135,N_30915);
xnor U33864 (N_33864,N_31200,N_31758);
or U33865 (N_33865,N_31616,N_31576);
or U33866 (N_33866,N_31835,N_30589);
or U33867 (N_33867,N_31991,N_30118);
nand U33868 (N_33868,N_31606,N_31848);
or U33869 (N_33869,N_30866,N_30360);
xor U33870 (N_33870,N_30172,N_31706);
nand U33871 (N_33871,N_30125,N_31564);
nor U33872 (N_33872,N_31543,N_31550);
nand U33873 (N_33873,N_31049,N_31430);
nor U33874 (N_33874,N_31157,N_31210);
nor U33875 (N_33875,N_30870,N_30860);
xor U33876 (N_33876,N_31048,N_31425);
nor U33877 (N_33877,N_30173,N_30617);
xor U33878 (N_33878,N_30018,N_31335);
and U33879 (N_33879,N_31418,N_31051);
or U33880 (N_33880,N_31895,N_31908);
nor U33881 (N_33881,N_31493,N_30903);
nor U33882 (N_33882,N_30641,N_30059);
nor U33883 (N_33883,N_31615,N_31461);
nor U33884 (N_33884,N_31647,N_31886);
xor U33885 (N_33885,N_30767,N_31616);
and U33886 (N_33886,N_31890,N_30348);
and U33887 (N_33887,N_31208,N_31132);
nand U33888 (N_33888,N_30377,N_31550);
xnor U33889 (N_33889,N_31307,N_31642);
and U33890 (N_33890,N_31934,N_30510);
xnor U33891 (N_33891,N_31893,N_31301);
nand U33892 (N_33892,N_30579,N_31125);
nor U33893 (N_33893,N_30141,N_30976);
nand U33894 (N_33894,N_30895,N_30501);
nand U33895 (N_33895,N_30217,N_31880);
xnor U33896 (N_33896,N_30471,N_30879);
or U33897 (N_33897,N_31364,N_31398);
nor U33898 (N_33898,N_30351,N_30193);
or U33899 (N_33899,N_31802,N_31491);
nand U33900 (N_33900,N_31324,N_30030);
or U33901 (N_33901,N_30922,N_31496);
nand U33902 (N_33902,N_30494,N_31062);
nand U33903 (N_33903,N_30686,N_30993);
nor U33904 (N_33904,N_30200,N_30669);
and U33905 (N_33905,N_31702,N_31613);
and U33906 (N_33906,N_30189,N_30681);
or U33907 (N_33907,N_30182,N_31570);
or U33908 (N_33908,N_30896,N_31862);
nand U33909 (N_33909,N_30111,N_30528);
nor U33910 (N_33910,N_31234,N_31088);
or U33911 (N_33911,N_30841,N_31964);
xnor U33912 (N_33912,N_31159,N_31519);
and U33913 (N_33913,N_30626,N_30994);
xor U33914 (N_33914,N_30179,N_30929);
xor U33915 (N_33915,N_30526,N_30077);
nand U33916 (N_33916,N_30706,N_31960);
nand U33917 (N_33917,N_31810,N_31619);
nand U33918 (N_33918,N_30014,N_30885);
and U33919 (N_33919,N_30407,N_31699);
and U33920 (N_33920,N_30453,N_31501);
or U33921 (N_33921,N_31025,N_30318);
or U33922 (N_33922,N_30465,N_30587);
xor U33923 (N_33923,N_31799,N_30277);
or U33924 (N_33924,N_31122,N_31956);
and U33925 (N_33925,N_30606,N_31818);
nand U33926 (N_33926,N_31477,N_30245);
and U33927 (N_33927,N_30922,N_30446);
or U33928 (N_33928,N_31973,N_31897);
or U33929 (N_33929,N_30795,N_31267);
nand U33930 (N_33930,N_31682,N_31813);
xnor U33931 (N_33931,N_30495,N_31350);
or U33932 (N_33932,N_30112,N_31195);
or U33933 (N_33933,N_31035,N_31577);
xor U33934 (N_33934,N_30117,N_31420);
nor U33935 (N_33935,N_30879,N_31498);
xor U33936 (N_33936,N_31313,N_31075);
nand U33937 (N_33937,N_30017,N_30425);
nor U33938 (N_33938,N_30983,N_30000);
xnor U33939 (N_33939,N_30050,N_31878);
and U33940 (N_33940,N_30894,N_30810);
nand U33941 (N_33941,N_30389,N_31742);
or U33942 (N_33942,N_30662,N_31989);
and U33943 (N_33943,N_30892,N_30546);
nand U33944 (N_33944,N_30879,N_31062);
nor U33945 (N_33945,N_30088,N_31499);
nor U33946 (N_33946,N_30705,N_30632);
and U33947 (N_33947,N_30190,N_31725);
or U33948 (N_33948,N_30603,N_30572);
and U33949 (N_33949,N_31146,N_31332);
and U33950 (N_33950,N_30192,N_31499);
xnor U33951 (N_33951,N_30063,N_30170);
and U33952 (N_33952,N_31010,N_30204);
nand U33953 (N_33953,N_31599,N_30777);
nor U33954 (N_33954,N_30285,N_30006);
nand U33955 (N_33955,N_31349,N_30754);
nor U33956 (N_33956,N_30668,N_31402);
or U33957 (N_33957,N_30206,N_31938);
xnor U33958 (N_33958,N_30456,N_30509);
nor U33959 (N_33959,N_31672,N_31735);
xor U33960 (N_33960,N_31023,N_31836);
or U33961 (N_33961,N_31891,N_30271);
and U33962 (N_33962,N_31205,N_30925);
nand U33963 (N_33963,N_30596,N_31286);
nand U33964 (N_33964,N_30538,N_30493);
or U33965 (N_33965,N_30057,N_31305);
nand U33966 (N_33966,N_30891,N_31352);
nor U33967 (N_33967,N_30529,N_31951);
or U33968 (N_33968,N_30725,N_30653);
xnor U33969 (N_33969,N_31972,N_30865);
nand U33970 (N_33970,N_30353,N_31168);
and U33971 (N_33971,N_30872,N_30691);
nand U33972 (N_33972,N_31157,N_31745);
nand U33973 (N_33973,N_31645,N_30063);
and U33974 (N_33974,N_30653,N_30976);
and U33975 (N_33975,N_30621,N_31521);
and U33976 (N_33976,N_30224,N_31799);
xnor U33977 (N_33977,N_31295,N_31141);
or U33978 (N_33978,N_30987,N_30246);
and U33979 (N_33979,N_30739,N_30567);
xnor U33980 (N_33980,N_31707,N_30614);
and U33981 (N_33981,N_31915,N_31407);
nand U33982 (N_33982,N_30279,N_30486);
xnor U33983 (N_33983,N_30291,N_30022);
xor U33984 (N_33984,N_30268,N_31124);
xor U33985 (N_33985,N_31338,N_30463);
or U33986 (N_33986,N_31647,N_30671);
xnor U33987 (N_33987,N_31832,N_31885);
or U33988 (N_33988,N_31031,N_30630);
nand U33989 (N_33989,N_31458,N_31746);
and U33990 (N_33990,N_30367,N_30178);
or U33991 (N_33991,N_31808,N_30609);
nor U33992 (N_33992,N_31137,N_31256);
and U33993 (N_33993,N_30874,N_30462);
and U33994 (N_33994,N_31083,N_31858);
xnor U33995 (N_33995,N_31060,N_30283);
nor U33996 (N_33996,N_30124,N_30334);
and U33997 (N_33997,N_31614,N_31058);
nor U33998 (N_33998,N_31429,N_31021);
nand U33999 (N_33999,N_30656,N_31457);
and U34000 (N_34000,N_32712,N_33126);
nand U34001 (N_34001,N_32932,N_32920);
nand U34002 (N_34002,N_32427,N_33658);
nand U34003 (N_34003,N_32101,N_33896);
or U34004 (N_34004,N_32460,N_33285);
xnor U34005 (N_34005,N_32434,N_32172);
nor U34006 (N_34006,N_33268,N_32474);
or U34007 (N_34007,N_32835,N_32940);
nor U34008 (N_34008,N_33461,N_33601);
and U34009 (N_34009,N_32355,N_33237);
and U34010 (N_34010,N_33457,N_32408);
nand U34011 (N_34011,N_32989,N_32665);
nand U34012 (N_34012,N_33392,N_33982);
nor U34013 (N_34013,N_33222,N_33231);
nand U34014 (N_34014,N_32549,N_33241);
xor U34015 (N_34015,N_32952,N_33146);
nor U34016 (N_34016,N_33689,N_32093);
nand U34017 (N_34017,N_33438,N_33447);
nor U34018 (N_34018,N_32201,N_32797);
nor U34019 (N_34019,N_33611,N_32259);
nor U34020 (N_34020,N_33193,N_33225);
xor U34021 (N_34021,N_32609,N_32969);
or U34022 (N_34022,N_33736,N_32730);
or U34023 (N_34023,N_32195,N_33659);
or U34024 (N_34024,N_32241,N_32530);
nand U34025 (N_34025,N_33706,N_32176);
nor U34026 (N_34026,N_33933,N_32115);
or U34027 (N_34027,N_33833,N_33883);
or U34028 (N_34028,N_33105,N_33687);
nand U34029 (N_34029,N_33304,N_33489);
xnor U34030 (N_34030,N_33522,N_32888);
nor U34031 (N_34031,N_33725,N_32826);
and U34032 (N_34032,N_33542,N_32647);
or U34033 (N_34033,N_32412,N_33113);
or U34034 (N_34034,N_32454,N_33159);
xor U34035 (N_34035,N_33127,N_32145);
or U34036 (N_34036,N_33840,N_33204);
xor U34037 (N_34037,N_32187,N_33618);
or U34038 (N_34038,N_32563,N_32105);
and U34039 (N_34039,N_33936,N_32949);
or U34040 (N_34040,N_32983,N_32475);
and U34041 (N_34041,N_33995,N_33643);
and U34042 (N_34042,N_32126,N_33791);
nand U34043 (N_34043,N_32897,N_32857);
nand U34044 (N_34044,N_32527,N_32662);
nand U34045 (N_34045,N_32059,N_32253);
xnor U34046 (N_34046,N_32124,N_33320);
nor U34047 (N_34047,N_33321,N_33178);
xor U34048 (N_34048,N_32764,N_33900);
or U34049 (N_34049,N_32260,N_33600);
xor U34050 (N_34050,N_32581,N_33755);
nand U34051 (N_34051,N_32246,N_33265);
nor U34052 (N_34052,N_33115,N_32638);
and U34053 (N_34053,N_33869,N_33753);
xnor U34054 (N_34054,N_32502,N_32250);
nand U34055 (N_34055,N_32316,N_33514);
xnor U34056 (N_34056,N_32432,N_32671);
nor U34057 (N_34057,N_33297,N_32049);
or U34058 (N_34058,N_33001,N_33598);
nand U34059 (N_34059,N_32875,N_32675);
xor U34060 (N_34060,N_33575,N_32776);
xnor U34061 (N_34061,N_32303,N_33502);
nor U34062 (N_34062,N_32078,N_33016);
xor U34063 (N_34063,N_32541,N_33993);
and U34064 (N_34064,N_33850,N_32375);
nor U34065 (N_34065,N_32491,N_33131);
and U34066 (N_34066,N_32570,N_33423);
nand U34067 (N_34067,N_32467,N_32240);
and U34068 (N_34068,N_32242,N_32650);
and U34069 (N_34069,N_32330,N_32437);
nand U34070 (N_34070,N_32286,N_32083);
nand U34071 (N_34071,N_33814,N_32018);
nor U34072 (N_34072,N_32569,N_33721);
xnor U34073 (N_34073,N_32881,N_33120);
or U34074 (N_34074,N_32244,N_32235);
or U34075 (N_34075,N_32088,N_33289);
nor U34076 (N_34076,N_32080,N_33182);
or U34077 (N_34077,N_32894,N_33130);
xor U34078 (N_34078,N_33385,N_32986);
and U34079 (N_34079,N_32615,N_33244);
nor U34080 (N_34080,N_32008,N_33352);
or U34081 (N_34081,N_33141,N_32933);
and U34082 (N_34082,N_32511,N_33930);
and U34083 (N_34083,N_32339,N_33992);
nor U34084 (N_34084,N_33607,N_33411);
nor U34085 (N_34085,N_32977,N_32085);
xor U34086 (N_34086,N_33587,N_32655);
nand U34087 (N_34087,N_32545,N_33169);
nand U34088 (N_34088,N_33745,N_33345);
nor U34089 (N_34089,N_32370,N_33101);
xnor U34090 (N_34090,N_33813,N_32318);
nand U34091 (N_34091,N_33586,N_32081);
and U34092 (N_34092,N_33501,N_33625);
or U34093 (N_34093,N_33326,N_32923);
or U34094 (N_34094,N_32689,N_32030);
nand U34095 (N_34095,N_33991,N_32458);
nand U34096 (N_34096,N_32506,N_33458);
and U34097 (N_34097,N_33743,N_33531);
or U34098 (N_34098,N_32363,N_32700);
or U34099 (N_34099,N_32392,N_33367);
and U34100 (N_34100,N_33571,N_32440);
or U34101 (N_34101,N_32829,N_32902);
and U34102 (N_34102,N_32221,N_32291);
and U34103 (N_34103,N_33932,N_32684);
or U34104 (N_34104,N_33944,N_33094);
nor U34105 (N_34105,N_33842,N_32896);
nor U34106 (N_34106,N_32336,N_32783);
or U34107 (N_34107,N_32144,N_33556);
and U34108 (N_34108,N_33477,N_33221);
or U34109 (N_34109,N_32792,N_33012);
nor U34110 (N_34110,N_33901,N_32814);
or U34111 (N_34111,N_32086,N_32926);
xor U34112 (N_34112,N_33987,N_32677);
nor U34113 (N_34113,N_32074,N_33198);
nor U34114 (N_34114,N_32848,N_33639);
or U34115 (N_34115,N_33980,N_32775);
or U34116 (N_34116,N_32624,N_33647);
nor U34117 (N_34117,N_33621,N_32247);
nand U34118 (N_34118,N_32091,N_33748);
xor U34119 (N_34119,N_32343,N_33615);
or U34120 (N_34120,N_32271,N_32866);
nor U34121 (N_34121,N_32492,N_33952);
and U34122 (N_34122,N_32610,N_32180);
xnor U34123 (N_34123,N_33908,N_33986);
or U34124 (N_34124,N_33741,N_32519);
or U34125 (N_34125,N_33316,N_32514);
or U34126 (N_34126,N_33355,N_32041);
xor U34127 (N_34127,N_33811,N_33845);
and U34128 (N_34128,N_32297,N_32497);
or U34129 (N_34129,N_33638,N_33125);
and U34130 (N_34130,N_33123,N_32510);
nand U34131 (N_34131,N_33979,N_33533);
nand U34132 (N_34132,N_33319,N_33312);
or U34133 (N_34133,N_32140,N_32203);
nor U34134 (N_34134,N_32279,N_33242);
xnor U34135 (N_34135,N_32032,N_33894);
nor U34136 (N_34136,N_33603,N_32913);
nor U34137 (N_34137,N_33379,N_33313);
or U34138 (N_34138,N_33975,N_33938);
and U34139 (N_34139,N_33463,N_32646);
or U34140 (N_34140,N_33583,N_32155);
nand U34141 (N_34141,N_32064,N_32167);
xor U34142 (N_34142,N_32979,N_32660);
or U34143 (N_34143,N_33767,N_33035);
or U34144 (N_34144,N_33782,N_33527);
and U34145 (N_34145,N_33327,N_32236);
nor U34146 (N_34146,N_33965,N_33712);
and U34147 (N_34147,N_32205,N_32594);
nand U34148 (N_34148,N_32309,N_33255);
or U34149 (N_34149,N_33063,N_33181);
nor U34150 (N_34150,N_33253,N_33164);
nor U34151 (N_34151,N_33645,N_32114);
and U34152 (N_34152,N_32890,N_32395);
xnor U34153 (N_34153,N_33462,N_33346);
and U34154 (N_34154,N_33849,N_33910);
and U34155 (N_34155,N_32777,N_33314);
or U34156 (N_34156,N_32364,N_33128);
xnor U34157 (N_34157,N_33047,N_32191);
xor U34158 (N_34158,N_33545,N_32281);
xor U34159 (N_34159,N_33819,N_32351);
xnor U34160 (N_34160,N_32693,N_33261);
and U34161 (N_34161,N_32526,N_33860);
nor U34162 (N_34162,N_32625,N_33455);
xnor U34163 (N_34163,N_32914,N_33914);
or U34164 (N_34164,N_33177,N_32518);
and U34165 (N_34165,N_32404,N_33758);
nor U34166 (N_34166,N_32498,N_32982);
nand U34167 (N_34167,N_33673,N_33139);
xor U34168 (N_34168,N_32142,N_33072);
nor U34169 (N_34169,N_33688,N_33369);
or U34170 (N_34170,N_32354,N_33140);
or U34171 (N_34171,N_33990,N_32861);
nor U34172 (N_34172,N_33664,N_33570);
nor U34173 (N_34173,N_33719,N_33170);
nor U34174 (N_34174,N_32252,N_33051);
nand U34175 (N_34175,N_33613,N_33295);
or U34176 (N_34176,N_33796,N_33768);
nand U34177 (N_34177,N_33299,N_33300);
nor U34178 (N_34178,N_33847,N_32596);
nand U34179 (N_34179,N_33731,N_32739);
and U34180 (N_34180,N_33428,N_32716);
or U34181 (N_34181,N_33311,N_32143);
xnor U34182 (N_34182,N_33760,N_32346);
and U34183 (N_34183,N_33947,N_32729);
and U34184 (N_34184,N_33330,N_33812);
nand U34185 (N_34185,N_33494,N_33398);
and U34186 (N_34186,N_33949,N_32161);
and U34187 (N_34187,N_32299,N_33200);
and U34188 (N_34188,N_32870,N_32283);
and U34189 (N_34189,N_33946,N_32820);
xor U34190 (N_34190,N_32906,N_32277);
or U34191 (N_34191,N_33210,N_33629);
nor U34192 (N_34192,N_32543,N_32521);
xor U34193 (N_34193,N_32839,N_33276);
nor U34194 (N_34194,N_32500,N_33858);
or U34195 (N_34195,N_33523,N_32988);
nor U34196 (N_34196,N_32028,N_32159);
nor U34197 (N_34197,N_33358,N_32535);
xnor U34198 (N_34198,N_32054,N_33637);
nand U34199 (N_34199,N_32168,N_33623);
xor U34200 (N_34200,N_32342,N_32595);
and U34201 (N_34201,N_32052,N_32275);
or U34202 (N_34202,N_33715,N_32413);
and U34203 (N_34203,N_33082,N_32635);
nand U34204 (N_34204,N_33109,N_32925);
xor U34205 (N_34205,N_32889,N_33862);
nand U34206 (N_34206,N_33007,N_33493);
and U34207 (N_34207,N_33891,N_32048);
nor U34208 (N_34208,N_32555,N_33877);
and U34209 (N_34209,N_33310,N_32727);
nor U34210 (N_34210,N_33301,N_32778);
nor U34211 (N_34211,N_33927,N_32266);
nand U34212 (N_34212,N_33110,N_33260);
nand U34213 (N_34213,N_33735,N_32834);
and U34214 (N_34214,N_33165,N_32307);
or U34215 (N_34215,N_32770,N_33209);
or U34216 (N_34216,N_33716,N_33839);
and U34217 (N_34217,N_32269,N_32607);
nand U34218 (N_34218,N_32789,N_32606);
or U34219 (N_34219,N_33121,N_32760);
xor U34220 (N_34220,N_32181,N_33202);
or U34221 (N_34221,N_33981,N_33187);
or U34222 (N_34222,N_32189,N_32341);
nor U34223 (N_34223,N_33805,N_32466);
nand U34224 (N_34224,N_32488,N_33566);
and U34225 (N_34225,N_33642,N_32401);
nand U34226 (N_34226,N_33427,N_32423);
and U34227 (N_34227,N_33167,N_32153);
xor U34228 (N_34228,N_32938,N_32332);
xor U34229 (N_34229,N_32106,N_33046);
and U34230 (N_34230,N_33801,N_32453);
nand U34231 (N_34231,N_33377,N_33834);
and U34232 (N_34232,N_33400,N_33841);
nand U34233 (N_34233,N_33406,N_33405);
or U34234 (N_34234,N_33492,N_32016);
nor U34235 (N_34235,N_33614,N_32199);
nor U34236 (N_34236,N_33153,N_32072);
or U34237 (N_34237,N_32827,N_32495);
and U34238 (N_34238,N_32688,N_32053);
nor U34239 (N_34239,N_32382,N_33171);
nor U34240 (N_34240,N_33240,N_32991);
or U34241 (N_34241,N_33506,N_33386);
or U34242 (N_34242,N_33179,N_33835);
nor U34243 (N_34243,N_32147,N_33342);
nor U34244 (N_34244,N_33137,N_33983);
or U34245 (N_34245,N_33205,N_32691);
nor U34246 (N_34246,N_33283,N_32234);
nor U34247 (N_34247,N_33752,N_32941);
nand U34248 (N_34248,N_33157,N_33597);
nand U34249 (N_34249,N_33372,N_32865);
nor U34250 (N_34250,N_33609,N_33472);
nor U34251 (N_34251,N_32574,N_33925);
and U34252 (N_34252,N_33184,N_32046);
nand U34253 (N_34253,N_33953,N_32703);
xor U34254 (N_34254,N_32109,N_32715);
xnor U34255 (N_34255,N_33086,N_32702);
nor U34256 (N_34256,N_33911,N_33885);
nand U34257 (N_34257,N_33083,N_32780);
nor U34258 (N_34258,N_32674,N_33470);
or U34259 (N_34259,N_33878,N_33519);
or U34260 (N_34260,N_33680,N_33524);
nor U34261 (N_34261,N_32415,N_33696);
nand U34262 (N_34262,N_33665,N_32701);
or U34263 (N_34263,N_33703,N_33401);
or U34264 (N_34264,N_32999,N_32405);
nand U34265 (N_34265,N_32899,N_32451);
or U34266 (N_34266,N_32507,N_32024);
nor U34267 (N_34267,N_32344,N_32123);
xnor U34268 (N_34268,N_33194,N_32823);
xnor U34269 (N_34269,N_32695,N_33563);
nand U34270 (N_34270,N_32374,N_32171);
nor U34271 (N_34271,N_32350,N_33259);
nand U34272 (N_34272,N_33469,N_32044);
and U34273 (N_34273,N_32637,N_32146);
or U34274 (N_34274,N_33104,N_33449);
and U34275 (N_34275,N_33988,N_33905);
xnor U34276 (N_34276,N_33882,N_32748);
or U34277 (N_34277,N_33510,N_32393);
or U34278 (N_34278,N_33599,N_33433);
nor U34279 (N_34279,N_32591,N_33019);
xor U34280 (N_34280,N_32371,N_33871);
nand U34281 (N_34281,N_33360,N_32447);
and U34282 (N_34282,N_32619,N_33717);
and U34283 (N_34283,N_33430,N_32213);
nor U34284 (N_34284,N_33765,N_33818);
xor U34285 (N_34285,N_32978,N_32218);
nand U34286 (N_34286,N_32192,N_33776);
and U34287 (N_34287,N_33410,N_33854);
nand U34288 (N_34288,N_33906,N_32111);
or U34289 (N_34289,N_33544,N_33666);
nand U34290 (N_34290,N_32851,N_33008);
or U34291 (N_34291,N_32893,N_32904);
and U34292 (N_34292,N_33118,N_33266);
nor U34293 (N_34293,N_33511,N_33997);
or U34294 (N_34294,N_32939,N_32095);
xnor U34295 (N_34295,N_32485,N_33418);
nor U34296 (N_34296,N_33112,N_32104);
nand U34297 (N_34297,N_32622,N_32224);
nor U34298 (N_34298,N_33561,N_33678);
or U34299 (N_34299,N_33280,N_33577);
nor U34300 (N_34300,N_32504,N_33488);
nor U34301 (N_34301,N_32930,N_32854);
and U34302 (N_34302,N_32496,N_33790);
or U34303 (N_34303,N_32089,N_33568);
or U34304 (N_34304,N_33440,N_33339);
or U34305 (N_34305,N_33394,N_33507);
or U34306 (N_34306,N_33002,N_33432);
and U34307 (N_34307,N_32766,N_32821);
and U34308 (N_34308,N_32763,N_33770);
or U34309 (N_34309,N_33749,N_32166);
or U34310 (N_34310,N_32396,N_33234);
and U34311 (N_34311,N_32828,N_32464);
and U34312 (N_34312,N_32558,N_33567);
or U34313 (N_34313,N_32758,N_32924);
or U34314 (N_34314,N_32634,N_32811);
nor U34315 (N_34315,N_32002,N_33562);
and U34316 (N_34316,N_32931,N_33293);
and U34317 (N_34317,N_33889,N_32859);
nand U34318 (N_34318,N_32756,N_33453);
or U34319 (N_34319,N_33604,N_32333);
and U34320 (N_34320,N_33998,N_32749);
xnor U34321 (N_34321,N_32604,N_33294);
or U34322 (N_34322,N_33048,N_32338);
nor U34323 (N_34323,N_33864,N_32759);
and U34324 (N_34324,N_33122,N_33606);
and U34325 (N_34325,N_32628,N_33117);
and U34326 (N_34326,N_32314,N_33692);
and U34327 (N_34327,N_33174,N_32478);
xnor U34328 (N_34328,N_32833,N_32334);
nand U34329 (N_34329,N_32420,N_32233);
nand U34330 (N_34330,N_33956,N_32288);
or U34331 (N_34331,N_33709,N_33092);
nor U34332 (N_34332,N_32229,N_33846);
xnor U34333 (N_34333,N_32446,N_32562);
or U34334 (N_34334,N_32544,N_32482);
nor U34335 (N_34335,N_33484,N_32887);
and U34336 (N_34336,N_33413,N_32373);
or U34337 (N_34337,N_32304,N_32121);
nand U34338 (N_34338,N_33075,N_32694);
or U34339 (N_34339,N_32036,N_33341);
xnor U34340 (N_34340,N_33375,N_33150);
nand U34341 (N_34341,N_33694,N_32154);
xnor U34342 (N_34342,N_32225,N_33747);
nor U34343 (N_34343,N_32073,N_32540);
nand U34344 (N_34344,N_33976,N_33887);
xor U34345 (N_34345,N_32290,N_32974);
and U34346 (N_34346,N_33918,N_33388);
and U34347 (N_34347,N_32442,N_32282);
nor U34348 (N_34348,N_33274,N_32394);
nand U34349 (N_34349,N_32836,N_32965);
xor U34350 (N_34350,N_33649,N_32704);
xnor U34351 (N_34351,N_33421,N_32468);
xnor U34352 (N_34352,N_33160,N_32348);
and U34353 (N_34353,N_33508,N_32801);
and U34354 (N_34354,N_32377,N_32108);
xor U34355 (N_34355,N_32416,N_33547);
or U34356 (N_34356,N_32151,N_33628);
nand U34357 (N_34357,N_33435,N_33929);
nor U34358 (N_34358,N_32627,N_33409);
nor U34359 (N_34359,N_33710,N_32705);
and U34360 (N_34360,N_32084,N_33357);
and U34361 (N_34361,N_32360,N_33076);
and U34362 (N_34362,N_32559,N_32220);
xor U34363 (N_34363,N_33229,N_32597);
nand U34364 (N_34364,N_33924,N_33318);
xnor U34365 (N_34365,N_33926,N_33317);
xnor U34366 (N_34366,N_33837,N_33897);
or U34367 (N_34367,N_32238,N_33702);
nand U34368 (N_34368,N_33798,N_32868);
nor U34369 (N_34369,N_32964,N_32157);
and U34370 (N_34370,N_33009,N_33704);
xnor U34371 (N_34371,N_33403,N_32735);
and U34372 (N_34372,N_32556,N_32481);
xor U34373 (N_34373,N_33608,N_33359);
nand U34374 (N_34374,N_33161,N_32217);
and U34375 (N_34375,N_32156,N_32957);
and U34376 (N_34376,N_32422,N_32842);
nor U34377 (N_34377,N_32503,N_33505);
nor U34378 (N_34378,N_32568,N_32306);
nor U34379 (N_34379,N_33291,N_33366);
nor U34380 (N_34380,N_33464,N_33303);
or U34381 (N_34381,N_33579,N_32118);
and U34382 (N_34382,N_32648,N_32886);
nand U34383 (N_34383,N_33822,N_32287);
and U34384 (N_34384,N_32626,N_32517);
nor U34385 (N_34385,N_33196,N_33536);
nor U34386 (N_34386,N_32471,N_33857);
or U34387 (N_34387,N_33670,N_33152);
nand U34388 (N_34388,N_33496,N_33081);
nand U34389 (N_34389,N_33335,N_32910);
nor U34390 (N_34390,N_32672,N_33836);
and U34391 (N_34391,N_32973,N_32661);
nand U34392 (N_34392,N_33580,N_33348);
nand U34393 (N_34393,N_32582,N_33859);
nand U34394 (N_34394,N_33111,N_33296);
xor U34395 (N_34395,N_33351,N_33080);
and U34396 (N_34396,N_33077,N_32043);
or U34397 (N_34397,N_32548,N_32682);
nor U34398 (N_34398,N_32007,N_32090);
xnor U34399 (N_34399,N_32552,N_33968);
or U34400 (N_34400,N_33762,N_33381);
and U34401 (N_34401,N_33873,N_33480);
xnor U34402 (N_34402,N_32456,N_33751);
nand U34403 (N_34403,N_32403,N_32516);
nor U34404 (N_34404,N_33771,N_33500);
nor U34405 (N_34405,N_32365,N_33816);
nand U34406 (N_34406,N_32127,N_32680);
nor U34407 (N_34407,N_32633,N_32215);
nand U34408 (N_34408,N_32227,N_32034);
and U34409 (N_34409,N_33656,N_32577);
and U34410 (N_34410,N_32771,N_33957);
or U34411 (N_34411,N_33434,N_32152);
nor U34412 (N_34412,N_33399,N_32915);
and U34413 (N_34413,N_33920,N_33707);
xor U34414 (N_34414,N_32445,N_32566);
or U34415 (N_34415,N_32005,N_33984);
nand U34416 (N_34416,N_33044,N_32023);
and U34417 (N_34417,N_32476,N_33886);
nand U34418 (N_34418,N_33934,N_33476);
or U34419 (N_34419,N_32844,N_32321);
nand U34420 (N_34420,N_33955,N_33003);
nand U34421 (N_34421,N_33373,N_33939);
xor U34422 (N_34422,N_32305,N_33763);
nor U34423 (N_34423,N_33331,N_33509);
nor U34424 (N_34424,N_32872,N_32390);
xnor U34425 (N_34425,N_32096,N_33940);
or U34426 (N_34426,N_32216,N_33958);
and U34427 (N_34427,N_33677,N_32752);
nor U34428 (N_34428,N_32576,N_32862);
xor U34429 (N_34429,N_32177,N_32045);
xnor U34430 (N_34430,N_32493,N_33922);
xnor U34431 (N_34431,N_32200,N_32435);
nand U34432 (N_34432,N_32193,N_32818);
and U34433 (N_34433,N_32796,N_33041);
nand U34434 (N_34434,N_32676,N_33156);
nor U34435 (N_34435,N_33114,N_33393);
or U34436 (N_34436,N_32945,N_32232);
xnor U34437 (N_34437,N_32734,N_33067);
nand U34438 (N_34438,N_33228,N_33641);
xor U34439 (N_34439,N_33066,N_32173);
nand U34440 (N_34440,N_33784,N_32103);
or U34441 (N_34441,N_33328,N_33879);
nor U34442 (N_34442,N_32039,N_33256);
nand U34443 (N_34443,N_33057,N_32198);
nand U34444 (N_34444,N_33444,N_33419);
nand U34445 (N_34445,N_32357,N_33148);
xnor U34446 (N_34446,N_33416,N_32807);
xnor U34447 (N_34447,N_32956,N_33429);
and U34448 (N_34448,N_32264,N_32219);
nor U34449 (N_34449,N_32022,N_32919);
or U34450 (N_34450,N_32524,N_32840);
nand U34451 (N_34451,N_32838,N_33258);
nor U34452 (N_34452,N_32075,N_33652);
nand U34453 (N_34453,N_33807,N_32006);
or U34454 (N_34454,N_32825,N_33985);
nor U34455 (N_34455,N_32179,N_33460);
and U34456 (N_34456,N_33653,N_33828);
or U34457 (N_34457,N_32785,N_33970);
or U34458 (N_34458,N_32575,N_32391);
and U34459 (N_34459,N_32690,N_33068);
nand U34460 (N_34460,N_33088,N_32428);
nor U34461 (N_34461,N_33555,N_32981);
and U34462 (N_34462,N_32398,N_32239);
and U34463 (N_34463,N_33190,N_32593);
or U34464 (N_34464,N_32386,N_32958);
and U34465 (N_34465,N_32267,N_33340);
or U34466 (N_34466,N_33569,N_32614);
nand U34467 (N_34467,N_32572,N_33730);
nand U34468 (N_34468,N_33275,N_32328);
xor U34469 (N_34469,N_33902,N_33064);
xor U34470 (N_34470,N_33573,N_32629);
nand U34471 (N_34471,N_33578,N_33269);
nor U34472 (N_34472,N_33000,N_32900);
nand U34473 (N_34473,N_33551,N_32513);
xor U34474 (N_34474,N_32686,N_33868);
nand U34475 (N_34475,N_33271,N_33162);
nand U34476 (N_34476,N_33584,N_32733);
xor U34477 (N_34477,N_32533,N_32852);
nor U34478 (N_34478,N_32431,N_32951);
or U34479 (N_34479,N_32165,N_32137);
or U34480 (N_34480,N_32800,N_33916);
nand U34481 (N_34481,N_33049,N_32553);
nand U34482 (N_34482,N_32640,N_32697);
and U34483 (N_34483,N_32069,N_32786);
or U34484 (N_34484,N_32349,N_32211);
and U34485 (N_34485,N_33948,N_32550);
xor U34486 (N_34486,N_33912,N_32546);
and U34487 (N_34487,N_32831,N_32150);
or U34488 (N_34488,N_32055,N_33292);
or U34489 (N_34489,N_33633,N_32580);
and U34490 (N_34490,N_32347,N_33227);
or U34491 (N_34491,N_32469,N_33517);
nand U34492 (N_34492,N_32148,N_32295);
or U34493 (N_34493,N_33674,N_32141);
and U34494 (N_34494,N_33040,N_33943);
and U34495 (N_34495,N_33116,N_32289);
nor U34496 (N_34496,N_32094,N_33030);
nor U34497 (N_34497,N_33497,N_33091);
and U34498 (N_34498,N_32922,N_32790);
or U34499 (N_34499,N_32616,N_33230);
nand U34500 (N_34500,N_33740,N_33071);
xnor U34501 (N_34501,N_32813,N_33691);
or U34502 (N_34502,N_33226,N_33516);
nand U34503 (N_34503,N_33278,N_33754);
or U34504 (N_34504,N_33942,N_33277);
nor U34505 (N_34505,N_33350,N_33683);
nand U34506 (N_34506,N_32439,N_32056);
or U34507 (N_34507,N_32087,N_32194);
or U34508 (N_34508,N_33364,N_33954);
xnor U34509 (N_34509,N_33962,N_33535);
and U34510 (N_34510,N_32630,N_32565);
nand U34511 (N_34511,N_32183,N_33711);
or U34512 (N_34512,N_33826,N_33056);
nor U34513 (N_34513,N_32489,N_32322);
nor U34514 (N_34514,N_32256,N_33408);
nor U34515 (N_34515,N_33026,N_33616);
nand U34516 (N_34516,N_33052,N_33412);
nand U34517 (N_34517,N_32663,N_32803);
xnor U34518 (N_34518,N_33693,N_33695);
and U34519 (N_34519,N_32651,N_33972);
xor U34520 (N_34520,N_32912,N_32131);
nand U34521 (N_34521,N_32430,N_33098);
or U34522 (N_34522,N_33804,N_33761);
nand U34523 (N_34523,N_32107,N_32788);
nand U34524 (N_34524,N_33459,N_32934);
nor U34525 (N_34525,N_32313,N_33344);
or U34526 (N_34526,N_33465,N_32452);
xor U34527 (N_34527,N_33062,N_33053);
or U34528 (N_34528,N_32285,N_33324);
xor U34529 (N_34529,N_32998,N_33005);
nor U34530 (N_34530,N_33572,N_32158);
nor U34531 (N_34531,N_32047,N_32603);
and U34532 (N_34532,N_33336,N_32658);
xnor U34533 (N_34533,N_32381,N_32029);
and U34534 (N_34534,N_32943,N_33713);
nor U34535 (N_34535,N_33852,N_33808);
and U34536 (N_34536,N_32966,N_33699);
nor U34537 (N_34537,N_32280,N_32494);
nor U34538 (N_34538,N_32679,N_32501);
or U34539 (N_34539,N_33679,N_33451);
or U34540 (N_34540,N_32708,N_33334);
nor U34541 (N_34541,N_32751,N_33893);
nor U34542 (N_34542,N_32927,N_32869);
and U34543 (N_34543,N_33349,N_33168);
or U34544 (N_34544,N_32257,N_32812);
and U34545 (N_34545,N_33937,N_32169);
nor U34546 (N_34546,N_32678,N_32822);
xor U34547 (N_34547,N_32830,N_33437);
nand U34548 (N_34548,N_33967,N_32385);
nor U34549 (N_34549,N_32301,N_33923);
or U34550 (N_34550,N_33635,N_33264);
and U34551 (N_34551,N_33994,N_32644);
and U34552 (N_34552,N_33473,N_33823);
nor U34553 (N_34553,N_32726,N_33096);
or U34554 (N_34554,N_33726,N_32027);
xor U34555 (N_34555,N_32426,N_32642);
nor U34556 (N_34556,N_33592,N_33787);
nor U34557 (N_34557,N_32531,N_33591);
or U34558 (N_34558,N_32001,N_32402);
nand U34559 (N_34559,N_33728,N_32209);
xnor U34560 (N_34560,N_33027,N_32448);
xor U34561 (N_34561,N_32207,N_32190);
nor U34562 (N_34562,N_33415,N_32774);
and U34563 (N_34563,N_33903,N_33622);
nand U34564 (N_34564,N_33651,N_33945);
xnor U34565 (N_34565,N_33017,N_33960);
nand U34566 (N_34566,N_32639,N_33632);
or U34567 (N_34567,N_32465,N_33966);
nor U34568 (N_34568,N_32681,N_33426);
nand U34569 (N_34569,N_33028,N_33780);
or U34570 (N_34570,N_33108,N_33746);
or U34571 (N_34571,N_32149,N_32909);
nor U34572 (N_34572,N_33207,N_33876);
xor U34573 (N_34573,N_33337,N_32399);
xor U34574 (N_34574,N_33596,N_33185);
and U34575 (N_34575,N_32206,N_33099);
nand U34576 (N_34576,N_32534,N_33548);
nor U34577 (N_34577,N_33550,N_32905);
or U34578 (N_34578,N_33799,N_32673);
and U34579 (N_34579,N_32683,N_32669);
nor U34580 (N_34580,N_32611,N_32331);
xor U34581 (N_34581,N_32874,N_33362);
xnor U34582 (N_34582,N_33549,N_32362);
xnor U34583 (N_34583,N_33676,N_33376);
nor U34584 (N_34584,N_32936,N_32557);
or U34585 (N_34585,N_33391,N_32017);
or U34586 (N_34586,N_32025,N_32038);
and U34587 (N_34587,N_32885,N_32372);
xor U34588 (N_34588,N_32824,N_32898);
or U34589 (N_34589,N_33727,N_32685);
xnor U34590 (N_34590,N_32585,N_32128);
and U34591 (N_34591,N_33010,N_32806);
nand U34592 (N_34592,N_32174,N_33778);
xor U34593 (N_34593,N_33498,N_33395);
or U34594 (N_34594,N_32536,N_33238);
or U34595 (N_34595,N_32214,N_32656);
nor U34596 (N_34596,N_33619,N_32539);
nor U34597 (N_34597,N_33107,N_33773);
and U34598 (N_34598,N_33951,N_33084);
and U34599 (N_34599,N_32736,N_32584);
or U34600 (N_34600,N_33119,N_32122);
and U34601 (N_34601,N_33284,N_33195);
and U34602 (N_34602,N_32387,N_33546);
nand U34603 (N_34603,N_32061,N_33777);
nand U34604 (N_34604,N_33206,N_33772);
nor U34605 (N_34605,N_33779,N_33733);
nor U34606 (N_34606,N_32380,N_33329);
nand U34607 (N_34607,N_32102,N_32810);
and U34608 (N_34608,N_33921,N_32272);
or U34609 (N_34609,N_33581,N_33404);
xnor U34610 (N_34610,N_33838,N_32937);
or U34611 (N_34611,N_33738,N_33732);
or U34612 (N_34612,N_33201,N_32421);
nand U34613 (N_34613,N_32294,N_32479);
xor U34614 (N_34614,N_33909,N_32714);
nand U34615 (N_34615,N_32653,N_33701);
or U34616 (N_34616,N_33759,N_32325);
nand U34617 (N_34617,N_32707,N_32042);
nand U34618 (N_34618,N_32598,N_32163);
xnor U34619 (N_34619,N_33018,N_32960);
nand U34620 (N_34620,N_32414,N_33675);
nand U34621 (N_34621,N_32876,N_33183);
nor U34622 (N_34622,N_33559,N_32959);
xor U34623 (N_34623,N_32794,N_33031);
and U34624 (N_34624,N_32077,N_33034);
xnor U34625 (N_34625,N_33267,N_32459);
xor U34626 (N_34626,N_33655,N_32837);
xor U34627 (N_34627,N_32311,N_33060);
xor U34628 (N_34628,N_33543,N_32486);
xnor U34629 (N_34629,N_32858,N_32185);
xor U34630 (N_34630,N_32589,N_33038);
nor U34631 (N_34631,N_33332,N_33378);
or U34632 (N_34632,N_33173,N_33884);
and U34633 (N_34633,N_32532,N_33971);
nor U34634 (N_34634,N_32832,N_32003);
and U34635 (N_34635,N_32755,N_33058);
nor U34636 (N_34636,N_32916,N_32632);
nor U34637 (N_34637,N_33262,N_33197);
nor U34638 (N_34638,N_33690,N_32366);
xnor U34639 (N_34639,N_32608,N_32740);
or U34640 (N_34640,N_33214,N_33681);
and U34641 (N_34641,N_33786,N_32742);
or U34642 (N_34642,N_33396,N_32963);
nor U34643 (N_34643,N_32617,N_33895);
nor U34644 (N_34644,N_33757,N_33499);
or U34645 (N_34645,N_32444,N_33824);
or U34646 (N_34646,N_32962,N_32731);
xor U34647 (N_34647,N_33245,N_33093);
or U34648 (N_34648,N_32659,N_33552);
and U34649 (N_34649,N_32134,N_32587);
nor U34650 (N_34650,N_32769,N_32389);
nor U34651 (N_34651,N_32907,N_32262);
and U34652 (N_34652,N_33203,N_32652);
nor U34653 (N_34653,N_32228,N_33783);
xnor U34654 (N_34654,N_32573,N_32809);
and U34655 (N_34655,N_32196,N_33686);
nor U34656 (N_34656,N_33192,N_33588);
nor U34657 (N_34657,N_32612,N_33043);
nand U34658 (N_34658,N_33797,N_33750);
and U34659 (N_34659,N_32954,N_32062);
nand U34660 (N_34660,N_33103,N_32070);
xor U34661 (N_34661,N_32345,N_33243);
nand U34662 (N_34662,N_33087,N_32429);
nor U34663 (N_34663,N_33149,N_33302);
nor U34664 (N_34664,N_32120,N_32113);
and U34665 (N_34665,N_33931,N_32722);
nand U34666 (N_34666,N_33478,N_32747);
or U34667 (N_34667,N_32948,N_32138);
and U34668 (N_34668,N_32976,N_32011);
nand U34669 (N_34669,N_33425,N_33235);
xor U34670 (N_34670,N_33624,N_33919);
xnor U34671 (N_34671,N_32480,N_32706);
xor U34672 (N_34672,N_32184,N_32400);
xnor U34673 (N_34673,N_33466,N_32579);
and U34674 (N_34674,N_32738,N_32551);
xor U34675 (N_34675,N_33610,N_33907);
or U34676 (N_34676,N_33315,N_33070);
nor U34677 (N_34677,N_32720,N_33023);
or U34678 (N_34678,N_33417,N_32324);
nor U34679 (N_34679,N_32737,N_32098);
nand U34680 (N_34680,N_32268,N_33354);
nand U34681 (N_34681,N_32441,N_33530);
xor U34682 (N_34682,N_32746,N_32768);
xnor U34683 (N_34683,N_33263,N_32970);
xor U34684 (N_34684,N_33590,N_33079);
or U34685 (N_34685,N_32186,N_32119);
nand U34686 (N_34686,N_32721,N_33212);
xnor U34687 (N_34687,N_32878,N_33644);
xor U34688 (N_34688,N_33322,N_33368);
xor U34689 (N_34689,N_32197,N_32009);
xnor U34690 (N_34690,N_33347,N_33996);
or U34691 (N_34691,N_32641,N_33486);
xor U34692 (N_34692,N_33969,N_33538);
xnor U34693 (N_34693,N_33724,N_32164);
or U34694 (N_34694,N_33917,N_32019);
nand U34695 (N_34695,N_33729,N_32779);
and U34696 (N_34696,N_32529,N_32623);
nor U34697 (N_34697,N_33065,N_33021);
nand U34698 (N_34698,N_32254,N_32000);
or U34699 (N_34699,N_33802,N_32984);
and U34700 (N_34700,N_33282,N_33853);
or U34701 (N_34701,N_32877,N_33648);
xor U34702 (N_34702,N_32649,N_32050);
nand U34703 (N_34703,N_33420,N_33217);
nor U34704 (N_34704,N_33520,N_33085);
nand U34705 (N_34705,N_33904,N_32356);
and U34706 (N_34706,N_32378,N_33667);
or U34707 (N_34707,N_32512,N_32040);
and U34708 (N_34708,N_33881,N_32112);
or U34709 (N_34709,N_32696,N_33720);
nand U34710 (N_34710,N_32066,N_33036);
nor U34711 (N_34711,N_33353,N_32406);
xor U34712 (N_34712,N_32583,N_32315);
and U34713 (N_34713,N_33935,N_32578);
or U34714 (N_34714,N_33491,N_32419);
xor U34715 (N_34715,N_32160,N_32987);
and U34716 (N_34716,N_33220,N_33143);
or U34717 (N_34717,N_32805,N_32975);
nand U34718 (N_34718,N_33448,N_32586);
xnor U34719 (N_34719,N_32798,N_33504);
nor U34720 (N_34720,N_33325,N_33661);
nor U34721 (N_34721,N_33215,N_33769);
xor U34722 (N_34722,N_32856,N_33576);
xor U34723 (N_34723,N_33554,N_33697);
or U34724 (N_34724,N_32815,N_32621);
xnor U34725 (N_34725,N_33585,N_32182);
nor U34726 (N_34726,N_32515,N_33431);
xor U34727 (N_34727,N_32484,N_33513);
xnor U34728 (N_34728,N_33529,N_32741);
nor U34729 (N_34729,N_33147,N_33020);
xor U34730 (N_34730,N_32462,N_33154);
nor U34731 (N_34731,N_33663,N_32060);
nand U34732 (N_34732,N_33650,N_32026);
nor U34733 (N_34733,N_32895,N_32808);
or U34734 (N_34734,N_33880,N_32520);
or U34735 (N_34735,N_32483,N_32082);
nand U34736 (N_34736,N_32967,N_33142);
or U34737 (N_34737,N_32243,N_33443);
or U34738 (N_34738,N_33668,N_32961);
nand U34739 (N_34739,N_33380,N_32079);
or U34740 (N_34740,N_32433,N_32571);
xor U34741 (N_34741,N_33135,N_32202);
xnor U34742 (N_34742,N_33382,N_32368);
nand U34743 (N_34743,N_32772,N_32132);
nor U34744 (N_34744,N_32110,N_32525);
nor U34745 (N_34745,N_32352,N_33132);
and U34746 (N_34746,N_32170,N_32097);
and U34747 (N_34747,N_33815,N_33742);
or U34748 (N_34748,N_32645,N_32718);
nand U34749 (N_34749,N_32773,N_32509);
nand U34750 (N_34750,N_33323,N_32980);
xnor U34751 (N_34751,N_33672,N_32162);
and U34752 (N_34752,N_33795,N_33155);
nand U34753 (N_34753,N_32664,N_32058);
nand U34754 (N_34754,N_32804,N_33630);
xnor U34755 (N_34755,N_33574,N_32411);
or U34756 (N_34756,N_33756,N_33831);
nor U34757 (N_34757,N_32276,N_33482);
nand U34758 (N_34758,N_32463,N_33785);
or U34759 (N_34759,N_33033,N_33166);
or U34760 (N_34760,N_33384,N_33525);
or U34761 (N_34761,N_33471,N_33129);
nor U34762 (N_34762,N_32699,N_32249);
or U34763 (N_34763,N_33442,N_33698);
or U34764 (N_34764,N_33199,N_32237);
xor U34765 (N_34765,N_32505,N_32388);
xnor U34766 (N_34766,N_32744,N_33305);
or U34767 (N_34767,N_32523,N_32477);
or U34768 (N_34768,N_33281,N_33298);
nor U34769 (N_34769,N_32762,N_33356);
nand U34770 (N_34770,N_32883,N_32935);
nand U34771 (N_34771,N_33186,N_32996);
or U34772 (N_34772,N_32841,N_33999);
xnor U34773 (N_34773,N_33875,N_33407);
nand U34774 (N_34774,N_32068,N_33867);
and U34775 (N_34775,N_32719,N_33011);
xnor U34776 (N_34776,N_33863,N_33832);
and U34777 (N_34777,N_33055,N_32490);
nor U34778 (N_34778,N_32992,N_33809);
or U34779 (N_34779,N_32135,N_33387);
nor U34780 (N_34780,N_32139,N_33250);
nand U34781 (N_34781,N_32537,N_32226);
and U34782 (N_34782,N_32643,N_32329);
nor U34783 (N_34783,N_32994,N_33634);
or U34784 (N_34784,N_32561,N_33279);
xor U34785 (N_34785,N_33978,N_32470);
xor U34786 (N_34786,N_32410,N_32319);
xnor U34787 (N_34787,N_32732,N_33565);
xnor U34788 (N_34788,N_32130,N_33436);
or U34789 (N_34789,N_33307,N_33445);
nand U34790 (N_34790,N_32397,N_32302);
nand U34791 (N_34791,N_33456,N_33503);
nand U34792 (N_34792,N_32728,N_33133);
nand U34793 (N_34793,N_32560,N_33100);
or U34794 (N_34794,N_33553,N_32754);
nand U34795 (N_34795,N_32255,N_32620);
nor U34796 (N_34796,N_33025,N_33069);
or U34797 (N_34797,N_32968,N_33037);
or U34798 (N_34798,N_33532,N_33468);
xnor U34799 (N_34799,N_33806,N_33843);
and U34800 (N_34800,N_32031,N_33640);
xor U34801 (N_34801,N_33684,N_32099);
nand U34802 (N_34802,N_33254,N_32450);
nor U34803 (N_34803,N_33039,N_33208);
nor U34804 (N_34804,N_32717,N_33827);
nand U34805 (N_34805,N_33631,N_32947);
nand U34806 (N_34806,N_32407,N_33223);
or U34807 (N_34807,N_33708,N_33211);
or U34808 (N_34808,N_32667,N_33792);
nand U34809 (N_34809,N_32745,N_32317);
and U34810 (N_34810,N_33774,N_32037);
and U34811 (N_34811,N_32757,N_32767);
nor U34812 (N_34812,N_33251,N_32449);
and U34813 (N_34813,N_33539,N_32293);
nand U34814 (N_34814,N_33861,N_33989);
nand U34815 (N_34815,N_33671,N_32340);
and U34816 (N_34816,N_33095,N_33467);
or U34817 (N_34817,N_32817,N_32273);
and U34818 (N_34818,N_33825,N_32361);
xor U34819 (N_34819,N_33872,N_32864);
nor U34820 (N_34820,N_33582,N_33248);
nand U34821 (N_34821,N_32847,N_33888);
nor U34822 (N_34822,N_33402,N_32251);
or U34823 (N_34823,N_33662,N_33793);
nand U34824 (N_34824,N_32670,N_32358);
xnor U34825 (N_34825,N_32911,N_33479);
nand U34826 (N_34826,N_33343,N_33714);
xnor U34827 (N_34827,N_33594,N_32212);
nand U34828 (N_34828,N_33899,N_33006);
or U34829 (N_34829,N_32178,N_32522);
xor U34830 (N_34830,N_33308,N_33928);
and U34831 (N_34831,N_33855,N_32076);
nor U34832 (N_34832,N_33974,N_33657);
xnor U34833 (N_34833,N_32600,N_33487);
xnor U34834 (N_34834,N_32725,N_32971);
nor U34835 (N_34835,N_33188,N_32997);
or U34836 (N_34836,N_32296,N_33829);
nor U34837 (N_34837,N_32605,N_33363);
or U34838 (N_34838,N_32750,N_33050);
or U34839 (N_34839,N_32133,N_33973);
or U34840 (N_34840,N_33144,N_32487);
xor U34841 (N_34841,N_33247,N_33249);
and U34842 (N_34842,N_33483,N_33090);
nand U34843 (N_34843,N_32245,N_32547);
nor U34844 (N_34844,N_32880,N_33595);
nand U34845 (N_34845,N_32010,N_32542);
nand U34846 (N_34846,N_33073,N_32284);
and U34847 (N_34847,N_32849,N_32882);
nand U34848 (N_34848,N_32320,N_32698);
or U34849 (N_34849,N_33383,N_32892);
nand U34850 (N_34850,N_33163,N_32051);
xor U34851 (N_34851,N_32129,N_32222);
and U34852 (N_34852,N_32853,N_33817);
nor U34853 (N_34853,N_32298,N_32443);
and U34854 (N_34854,N_32845,N_33270);
nor U34855 (N_34855,N_32636,N_32292);
xnor U34856 (N_34856,N_33232,N_33977);
and U34857 (N_34857,N_33950,N_33821);
nor U34858 (N_34858,N_32944,N_33361);
xor U34859 (N_34859,N_33022,N_32274);
nand U34860 (N_34860,N_32602,N_32021);
nand U34861 (N_34861,N_33257,N_32613);
and U34862 (N_34862,N_32383,N_33180);
nor U34863 (N_34863,N_33830,N_33454);
and U34864 (N_34864,N_33941,N_33589);
and U34865 (N_34865,N_33422,N_33481);
xnor U34866 (N_34866,N_33788,N_32753);
nand U34867 (N_34867,N_32908,N_33612);
xor U34868 (N_34868,N_33540,N_32100);
nand U34869 (N_34869,N_33014,N_32791);
nand U34870 (N_34870,N_33913,N_32843);
nor U34871 (N_34871,N_32499,N_33626);
nor U34872 (N_34872,N_32795,N_32950);
nor U34873 (N_34873,N_32035,N_32993);
nor U34874 (N_34874,N_32188,N_32327);
or U34875 (N_34875,N_33059,N_33272);
nand U34876 (N_34876,N_32782,N_32990);
nor U34877 (N_34877,N_33617,N_32743);
and U34878 (N_34878,N_32033,N_32724);
and U34879 (N_34879,N_32554,N_32457);
nor U34880 (N_34880,N_32946,N_32942);
and U34881 (N_34881,N_32117,N_33789);
and U34882 (N_34882,N_33306,N_32418);
and U34883 (N_34883,N_32472,N_33734);
xor U34884 (N_34884,N_32588,N_32326);
and U34885 (N_34885,N_33892,N_32230);
and U34886 (N_34886,N_32015,N_33236);
nor U34887 (N_34887,N_33865,N_33176);
xnor U34888 (N_34888,N_33189,N_33794);
or U34889 (N_34889,N_33371,N_33191);
nand U34890 (N_34890,N_32455,N_32248);
xor U34891 (N_34891,N_32873,N_33744);
nand U34892 (N_34892,N_32846,N_33485);
nor U34893 (N_34893,N_32860,N_33309);
nor U34894 (N_34894,N_33737,N_33475);
nand U34895 (N_34895,N_33963,N_32972);
nor U34896 (N_34896,N_33526,N_32310);
or U34897 (N_34897,N_33074,N_32955);
nor U34898 (N_34898,N_32263,N_32409);
nand U34899 (N_34899,N_32335,N_32816);
xor U34900 (N_34900,N_32850,N_32538);
nor U34901 (N_34901,N_32323,N_33218);
nand U34902 (N_34902,N_33534,N_33439);
and U34903 (N_34903,N_33078,N_33669);
xor U34904 (N_34904,N_32376,N_32508);
or U34905 (N_34905,N_33042,N_32424);
or U34906 (N_34906,N_33106,N_33959);
nor U34907 (N_34907,N_33333,N_33273);
and U34908 (N_34908,N_32590,N_32921);
nand U34909 (N_34909,N_33061,N_33851);
and U34910 (N_34910,N_32668,N_32359);
and U34911 (N_34911,N_32278,N_33848);
or U34912 (N_34912,N_33870,N_32687);
nand U34913 (N_34913,N_32425,N_33224);
nor U34914 (N_34914,N_33866,N_33172);
nor U34915 (N_34915,N_33781,N_33605);
nand U34916 (N_34916,N_33288,N_33898);
and U34917 (N_34917,N_33844,N_32592);
nand U34918 (N_34918,N_33015,N_32761);
xnor U34919 (N_34919,N_32929,N_33233);
or U34920 (N_34920,N_32802,N_32781);
and U34921 (N_34921,N_33803,N_32709);
xnor U34922 (N_34922,N_33004,N_32723);
or U34923 (N_34923,N_32210,N_33216);
xor U34924 (N_34924,N_33029,N_32116);
or U34925 (N_34925,N_32567,N_32901);
xnor U34926 (N_34926,N_33089,N_32231);
nor U34927 (N_34927,N_32631,N_32784);
nor U34928 (N_34928,N_32063,N_32308);
xnor U34929 (N_34929,N_33287,N_33134);
and U34930 (N_34930,N_33660,N_33239);
nor U34931 (N_34931,N_33964,N_33102);
xnor U34932 (N_34932,N_32618,N_32057);
nand U34933 (N_34933,N_33374,N_33446);
nor U34934 (N_34934,N_32312,N_33654);
or U34935 (N_34935,N_32461,N_33338);
xnor U34936 (N_34936,N_33557,N_32384);
and U34937 (N_34937,N_33045,N_33219);
nand U34938 (N_34938,N_32417,N_33136);
nor U34939 (N_34939,N_32918,N_33627);
xnor U34940 (N_34940,N_33452,N_33537);
or U34941 (N_34941,N_33723,N_33700);
and U34942 (N_34942,N_32004,N_33441);
or U34943 (N_34943,N_32599,N_33515);
nor U34944 (N_34944,N_33290,N_32787);
xor U34945 (N_34945,N_33685,N_32270);
nor U34946 (N_34946,N_33518,N_32300);
and U34947 (N_34947,N_32223,N_33054);
nor U34948 (N_34948,N_32884,N_32136);
nand U34949 (N_34949,N_32601,N_33705);
xnor U34950 (N_34950,N_33722,N_32020);
nand U34951 (N_34951,N_32436,N_33602);
nand U34952 (N_34952,N_32175,N_33775);
nand U34953 (N_34953,N_32713,N_32367);
xnor U34954 (N_34954,N_32871,N_32657);
or U34955 (N_34955,N_32473,N_32855);
or U34956 (N_34956,N_32369,N_32863);
nand U34957 (N_34957,N_32819,N_32879);
and U34958 (N_34958,N_32891,N_32013);
xor U34959 (N_34959,N_32917,N_33138);
nand U34960 (N_34960,N_33560,N_33646);
nand U34961 (N_34961,N_33246,N_33175);
and U34962 (N_34962,N_33158,N_33450);
nor U34963 (N_34963,N_32065,N_33365);
or U34964 (N_34964,N_33145,N_32014);
or U34965 (N_34965,N_32092,N_33764);
or U34966 (N_34966,N_33636,N_33474);
nand U34967 (N_34967,N_32995,N_32379);
xor U34968 (N_34968,N_32265,N_33389);
and U34969 (N_34969,N_33874,N_33593);
nand U34970 (N_34970,N_33810,N_32666);
and U34971 (N_34971,N_32953,N_33558);
nand U34972 (N_34972,N_32985,N_32564);
nand U34973 (N_34973,N_33528,N_33286);
or U34974 (N_34974,N_32799,N_33013);
nand U34975 (N_34975,N_32208,N_32710);
nand U34976 (N_34976,N_33370,N_33213);
nand U34977 (N_34977,N_32528,N_33739);
xor U34978 (N_34978,N_32765,N_32711);
xnor U34979 (N_34979,N_33414,N_33512);
xor U34980 (N_34980,N_32067,N_32692);
or U34981 (N_34981,N_33397,N_32337);
nand U34982 (N_34982,N_32793,N_32928);
xnor U34983 (N_34983,N_33890,N_33495);
nand U34984 (N_34984,N_33718,N_33521);
or U34985 (N_34985,N_33682,N_33961);
nor U34986 (N_34986,N_32903,N_33424);
and U34987 (N_34987,N_32654,N_32867);
and U34988 (N_34988,N_33032,N_33097);
and U34989 (N_34989,N_33024,N_33151);
nor U34990 (N_34990,N_32261,N_33390);
xnor U34991 (N_34991,N_33766,N_33541);
or U34992 (N_34992,N_33800,N_32204);
nor U34993 (N_34993,N_33820,N_32071);
or U34994 (N_34994,N_33915,N_32012);
nor U34995 (N_34995,N_32353,N_33252);
xnor U34996 (N_34996,N_33490,N_32438);
or U34997 (N_34997,N_32125,N_33620);
or U34998 (N_34998,N_33564,N_32258);
and U34999 (N_34999,N_33124,N_33856);
nand U35000 (N_35000,N_32678,N_32321);
and U35001 (N_35001,N_32894,N_32674);
nand U35002 (N_35002,N_33320,N_32770);
nand U35003 (N_35003,N_33953,N_32857);
xor U35004 (N_35004,N_33090,N_33367);
xor U35005 (N_35005,N_33280,N_33582);
nor U35006 (N_35006,N_32880,N_32351);
xor U35007 (N_35007,N_32404,N_33241);
xor U35008 (N_35008,N_32763,N_32742);
nand U35009 (N_35009,N_33041,N_33093);
nand U35010 (N_35010,N_32713,N_32031);
xor U35011 (N_35011,N_32042,N_32251);
and U35012 (N_35012,N_32304,N_33675);
xnor U35013 (N_35013,N_32911,N_33327);
nand U35014 (N_35014,N_33449,N_33102);
nand U35015 (N_35015,N_33984,N_32796);
nor U35016 (N_35016,N_32158,N_33638);
nand U35017 (N_35017,N_33961,N_33293);
nand U35018 (N_35018,N_32553,N_32479);
nor U35019 (N_35019,N_32410,N_33218);
or U35020 (N_35020,N_33049,N_32397);
nand U35021 (N_35021,N_32727,N_33750);
and U35022 (N_35022,N_32387,N_32929);
nor U35023 (N_35023,N_33822,N_32501);
nor U35024 (N_35024,N_32959,N_33337);
xnor U35025 (N_35025,N_33425,N_33020);
or U35026 (N_35026,N_32598,N_32342);
nor U35027 (N_35027,N_33036,N_33284);
xor U35028 (N_35028,N_32542,N_32851);
and U35029 (N_35029,N_32619,N_33050);
xnor U35030 (N_35030,N_32845,N_33284);
nand U35031 (N_35031,N_32218,N_33819);
xnor U35032 (N_35032,N_33504,N_33051);
nand U35033 (N_35033,N_33969,N_32444);
or U35034 (N_35034,N_33704,N_32638);
nor U35035 (N_35035,N_32794,N_33656);
and U35036 (N_35036,N_33116,N_32431);
xor U35037 (N_35037,N_33509,N_32558);
or U35038 (N_35038,N_32935,N_32197);
nand U35039 (N_35039,N_32188,N_33591);
and U35040 (N_35040,N_33423,N_33439);
or U35041 (N_35041,N_32668,N_32804);
and U35042 (N_35042,N_32726,N_33940);
and U35043 (N_35043,N_32825,N_33091);
or U35044 (N_35044,N_32189,N_32333);
and U35045 (N_35045,N_33520,N_32959);
xnor U35046 (N_35046,N_32409,N_32808);
or U35047 (N_35047,N_33729,N_32539);
xnor U35048 (N_35048,N_32376,N_33861);
nor U35049 (N_35049,N_33813,N_33620);
nand U35050 (N_35050,N_33096,N_33992);
nand U35051 (N_35051,N_32077,N_32946);
and U35052 (N_35052,N_33557,N_33074);
nand U35053 (N_35053,N_32922,N_33818);
xor U35054 (N_35054,N_33757,N_33872);
nand U35055 (N_35055,N_33004,N_32550);
nor U35056 (N_35056,N_32868,N_32781);
nor U35057 (N_35057,N_32178,N_32179);
nand U35058 (N_35058,N_32912,N_32156);
nand U35059 (N_35059,N_33486,N_32001);
and U35060 (N_35060,N_33242,N_32800);
xnor U35061 (N_35061,N_33007,N_33247);
nor U35062 (N_35062,N_33206,N_32712);
xor U35063 (N_35063,N_33885,N_32663);
xor U35064 (N_35064,N_33031,N_32223);
xnor U35065 (N_35065,N_33459,N_33424);
nand U35066 (N_35066,N_32537,N_32639);
xnor U35067 (N_35067,N_32155,N_33261);
or U35068 (N_35068,N_33224,N_32057);
xnor U35069 (N_35069,N_33277,N_32515);
and U35070 (N_35070,N_33710,N_32492);
nor U35071 (N_35071,N_33514,N_32699);
nand U35072 (N_35072,N_33250,N_32484);
nand U35073 (N_35073,N_33625,N_32428);
and U35074 (N_35074,N_32263,N_33349);
and U35075 (N_35075,N_33166,N_32059);
and U35076 (N_35076,N_32833,N_32670);
or U35077 (N_35077,N_32310,N_32081);
nand U35078 (N_35078,N_33014,N_32338);
and U35079 (N_35079,N_33511,N_33692);
and U35080 (N_35080,N_33896,N_33088);
xnor U35081 (N_35081,N_33291,N_33523);
and U35082 (N_35082,N_33869,N_33665);
and U35083 (N_35083,N_33380,N_33699);
nor U35084 (N_35084,N_32044,N_32418);
and U35085 (N_35085,N_33295,N_32147);
xnor U35086 (N_35086,N_33670,N_33521);
nand U35087 (N_35087,N_33941,N_32233);
xnor U35088 (N_35088,N_33660,N_33527);
and U35089 (N_35089,N_32825,N_33501);
and U35090 (N_35090,N_33007,N_33686);
xnor U35091 (N_35091,N_32927,N_33643);
nand U35092 (N_35092,N_33403,N_32404);
and U35093 (N_35093,N_32394,N_33564);
and U35094 (N_35094,N_32119,N_32093);
or U35095 (N_35095,N_33203,N_33179);
xnor U35096 (N_35096,N_32555,N_32946);
xnor U35097 (N_35097,N_33793,N_33245);
nand U35098 (N_35098,N_33658,N_32806);
or U35099 (N_35099,N_33197,N_32995);
nand U35100 (N_35100,N_33214,N_32846);
xor U35101 (N_35101,N_33623,N_33088);
and U35102 (N_35102,N_33638,N_33901);
nor U35103 (N_35103,N_32536,N_33250);
xnor U35104 (N_35104,N_33268,N_32057);
and U35105 (N_35105,N_32066,N_32182);
or U35106 (N_35106,N_33832,N_32819);
xor U35107 (N_35107,N_33889,N_32370);
xnor U35108 (N_35108,N_32324,N_33824);
nor U35109 (N_35109,N_33596,N_32189);
xor U35110 (N_35110,N_33747,N_33617);
nor U35111 (N_35111,N_33656,N_33186);
or U35112 (N_35112,N_32361,N_32331);
nand U35113 (N_35113,N_32547,N_33608);
xor U35114 (N_35114,N_33140,N_32720);
xnor U35115 (N_35115,N_32353,N_32663);
or U35116 (N_35116,N_33708,N_32283);
nor U35117 (N_35117,N_32725,N_32772);
nand U35118 (N_35118,N_33221,N_33209);
or U35119 (N_35119,N_33212,N_32019);
or U35120 (N_35120,N_33277,N_33132);
xnor U35121 (N_35121,N_33969,N_33063);
or U35122 (N_35122,N_32537,N_32117);
nand U35123 (N_35123,N_33572,N_32834);
or U35124 (N_35124,N_32708,N_32279);
nand U35125 (N_35125,N_33812,N_32140);
nand U35126 (N_35126,N_33739,N_32975);
and U35127 (N_35127,N_33237,N_33142);
xnor U35128 (N_35128,N_33413,N_32403);
nor U35129 (N_35129,N_32486,N_32557);
and U35130 (N_35130,N_32369,N_32376);
and U35131 (N_35131,N_32912,N_32029);
or U35132 (N_35132,N_32190,N_33116);
nor U35133 (N_35133,N_33620,N_33383);
or U35134 (N_35134,N_33736,N_33883);
xor U35135 (N_35135,N_33849,N_32239);
or U35136 (N_35136,N_32905,N_33753);
nand U35137 (N_35137,N_32784,N_33780);
xnor U35138 (N_35138,N_32437,N_33668);
nor U35139 (N_35139,N_33625,N_33633);
or U35140 (N_35140,N_32408,N_33067);
nand U35141 (N_35141,N_32269,N_32166);
xnor U35142 (N_35142,N_33980,N_33482);
nand U35143 (N_35143,N_33657,N_33728);
xnor U35144 (N_35144,N_33194,N_33911);
nand U35145 (N_35145,N_33031,N_33112);
nor U35146 (N_35146,N_32884,N_33571);
and U35147 (N_35147,N_33890,N_33886);
or U35148 (N_35148,N_33798,N_33870);
nor U35149 (N_35149,N_32669,N_33136);
xnor U35150 (N_35150,N_33906,N_33717);
and U35151 (N_35151,N_32794,N_32132);
xor U35152 (N_35152,N_33248,N_33644);
nand U35153 (N_35153,N_32448,N_32148);
nand U35154 (N_35154,N_32395,N_32089);
xnor U35155 (N_35155,N_32058,N_32123);
or U35156 (N_35156,N_32111,N_32840);
and U35157 (N_35157,N_33842,N_32047);
nand U35158 (N_35158,N_32059,N_32128);
or U35159 (N_35159,N_33083,N_32840);
nor U35160 (N_35160,N_33674,N_33911);
and U35161 (N_35161,N_33012,N_32280);
xnor U35162 (N_35162,N_33730,N_33402);
and U35163 (N_35163,N_33756,N_32328);
or U35164 (N_35164,N_32097,N_32922);
or U35165 (N_35165,N_32581,N_33635);
and U35166 (N_35166,N_32435,N_32346);
and U35167 (N_35167,N_33182,N_32521);
and U35168 (N_35168,N_33594,N_33808);
xor U35169 (N_35169,N_32950,N_33503);
or U35170 (N_35170,N_33995,N_32664);
and U35171 (N_35171,N_33391,N_33499);
or U35172 (N_35172,N_33659,N_33755);
nand U35173 (N_35173,N_32256,N_33915);
nor U35174 (N_35174,N_32195,N_33670);
xnor U35175 (N_35175,N_32680,N_32924);
xnor U35176 (N_35176,N_33030,N_32550);
or U35177 (N_35177,N_33631,N_33225);
and U35178 (N_35178,N_32582,N_32713);
nand U35179 (N_35179,N_32120,N_33938);
nor U35180 (N_35180,N_33445,N_33562);
xor U35181 (N_35181,N_32670,N_33662);
nand U35182 (N_35182,N_32009,N_32817);
and U35183 (N_35183,N_33706,N_32019);
xnor U35184 (N_35184,N_33208,N_32859);
and U35185 (N_35185,N_32326,N_32702);
xnor U35186 (N_35186,N_33118,N_32624);
or U35187 (N_35187,N_32718,N_33411);
and U35188 (N_35188,N_33821,N_32408);
or U35189 (N_35189,N_33274,N_32923);
nor U35190 (N_35190,N_33004,N_33542);
xnor U35191 (N_35191,N_33752,N_33654);
and U35192 (N_35192,N_33791,N_32016);
xor U35193 (N_35193,N_33051,N_33409);
or U35194 (N_35194,N_32902,N_33993);
and U35195 (N_35195,N_33822,N_32591);
nand U35196 (N_35196,N_32654,N_32216);
nand U35197 (N_35197,N_32630,N_33113);
or U35198 (N_35198,N_32937,N_32034);
nor U35199 (N_35199,N_33638,N_32448);
nand U35200 (N_35200,N_33760,N_33168);
nand U35201 (N_35201,N_32752,N_32487);
or U35202 (N_35202,N_33135,N_33207);
and U35203 (N_35203,N_33249,N_33694);
xor U35204 (N_35204,N_32638,N_33306);
and U35205 (N_35205,N_33395,N_33769);
nor U35206 (N_35206,N_32734,N_33405);
and U35207 (N_35207,N_33818,N_32510);
and U35208 (N_35208,N_33157,N_33905);
nand U35209 (N_35209,N_32641,N_32650);
or U35210 (N_35210,N_33219,N_32117);
nand U35211 (N_35211,N_33194,N_32568);
xnor U35212 (N_35212,N_32716,N_32431);
nor U35213 (N_35213,N_32257,N_33641);
nor U35214 (N_35214,N_33184,N_32010);
nand U35215 (N_35215,N_33450,N_32891);
and U35216 (N_35216,N_33959,N_32031);
or U35217 (N_35217,N_32929,N_33920);
nand U35218 (N_35218,N_33633,N_32427);
nand U35219 (N_35219,N_32384,N_32629);
xor U35220 (N_35220,N_32126,N_33726);
and U35221 (N_35221,N_33676,N_33461);
xor U35222 (N_35222,N_33992,N_33075);
nand U35223 (N_35223,N_33276,N_33944);
xor U35224 (N_35224,N_33666,N_32468);
or U35225 (N_35225,N_33773,N_33120);
xnor U35226 (N_35226,N_32573,N_33595);
xnor U35227 (N_35227,N_32320,N_33186);
and U35228 (N_35228,N_32481,N_33701);
or U35229 (N_35229,N_32562,N_33134);
xor U35230 (N_35230,N_32675,N_32514);
xor U35231 (N_35231,N_32716,N_32253);
xnor U35232 (N_35232,N_32196,N_33603);
and U35233 (N_35233,N_32766,N_32248);
nor U35234 (N_35234,N_33284,N_32209);
xor U35235 (N_35235,N_33582,N_32799);
and U35236 (N_35236,N_32468,N_32105);
or U35237 (N_35237,N_32055,N_32529);
xor U35238 (N_35238,N_32360,N_32050);
or U35239 (N_35239,N_32037,N_33657);
and U35240 (N_35240,N_32365,N_33050);
nor U35241 (N_35241,N_32489,N_32819);
and U35242 (N_35242,N_33035,N_32630);
nor U35243 (N_35243,N_32247,N_33052);
or U35244 (N_35244,N_33676,N_33345);
nand U35245 (N_35245,N_33736,N_32013);
and U35246 (N_35246,N_32294,N_33458);
and U35247 (N_35247,N_33982,N_33254);
and U35248 (N_35248,N_32917,N_32067);
xor U35249 (N_35249,N_33456,N_32631);
nor U35250 (N_35250,N_33000,N_33458);
xor U35251 (N_35251,N_32678,N_33674);
xor U35252 (N_35252,N_33613,N_32230);
nor U35253 (N_35253,N_32005,N_33672);
nor U35254 (N_35254,N_33190,N_33035);
or U35255 (N_35255,N_32059,N_32628);
xnor U35256 (N_35256,N_33818,N_32491);
xnor U35257 (N_35257,N_33164,N_32736);
xor U35258 (N_35258,N_32393,N_32746);
xnor U35259 (N_35259,N_32230,N_33439);
nand U35260 (N_35260,N_32678,N_32052);
or U35261 (N_35261,N_33043,N_33674);
nor U35262 (N_35262,N_32523,N_33852);
xor U35263 (N_35263,N_33768,N_32294);
nand U35264 (N_35264,N_33547,N_33242);
nor U35265 (N_35265,N_32946,N_32358);
or U35266 (N_35266,N_33610,N_33398);
nand U35267 (N_35267,N_32084,N_33328);
nand U35268 (N_35268,N_33389,N_33902);
nand U35269 (N_35269,N_33484,N_33490);
xor U35270 (N_35270,N_33014,N_32240);
nor U35271 (N_35271,N_32880,N_32189);
or U35272 (N_35272,N_33996,N_32320);
nand U35273 (N_35273,N_32954,N_33782);
xor U35274 (N_35274,N_33963,N_33764);
xor U35275 (N_35275,N_33688,N_32725);
and U35276 (N_35276,N_33194,N_32215);
nand U35277 (N_35277,N_33455,N_32392);
or U35278 (N_35278,N_32368,N_32288);
or U35279 (N_35279,N_32712,N_32151);
and U35280 (N_35280,N_32464,N_33106);
nor U35281 (N_35281,N_33219,N_32781);
xor U35282 (N_35282,N_33453,N_32127);
nand U35283 (N_35283,N_33516,N_32866);
and U35284 (N_35284,N_32659,N_32041);
and U35285 (N_35285,N_32844,N_33414);
or U35286 (N_35286,N_32641,N_33089);
or U35287 (N_35287,N_33648,N_32871);
and U35288 (N_35288,N_33262,N_33045);
or U35289 (N_35289,N_33063,N_32487);
xor U35290 (N_35290,N_33201,N_33861);
and U35291 (N_35291,N_32776,N_33316);
nor U35292 (N_35292,N_32310,N_32530);
nor U35293 (N_35293,N_32372,N_32161);
nor U35294 (N_35294,N_33217,N_33033);
and U35295 (N_35295,N_32005,N_32717);
and U35296 (N_35296,N_32836,N_33183);
xnor U35297 (N_35297,N_33352,N_33191);
or U35298 (N_35298,N_33502,N_33067);
and U35299 (N_35299,N_33556,N_33933);
or U35300 (N_35300,N_32411,N_32595);
or U35301 (N_35301,N_32178,N_33796);
nor U35302 (N_35302,N_32331,N_33961);
or U35303 (N_35303,N_33036,N_32199);
nand U35304 (N_35304,N_32591,N_32266);
xnor U35305 (N_35305,N_33184,N_33331);
xnor U35306 (N_35306,N_32616,N_33014);
nand U35307 (N_35307,N_32705,N_33527);
and U35308 (N_35308,N_33396,N_33464);
nand U35309 (N_35309,N_33711,N_33043);
or U35310 (N_35310,N_32323,N_33187);
nor U35311 (N_35311,N_33633,N_33691);
and U35312 (N_35312,N_32446,N_32607);
nor U35313 (N_35313,N_32092,N_32807);
nand U35314 (N_35314,N_32727,N_33162);
xor U35315 (N_35315,N_32561,N_33218);
nand U35316 (N_35316,N_32848,N_32627);
xor U35317 (N_35317,N_33980,N_33363);
and U35318 (N_35318,N_32220,N_33179);
nand U35319 (N_35319,N_33367,N_33777);
nand U35320 (N_35320,N_32336,N_32333);
or U35321 (N_35321,N_33216,N_32303);
nor U35322 (N_35322,N_33193,N_33110);
nand U35323 (N_35323,N_33676,N_33133);
xor U35324 (N_35324,N_33291,N_33078);
or U35325 (N_35325,N_33964,N_32194);
and U35326 (N_35326,N_33850,N_32011);
nand U35327 (N_35327,N_32830,N_32608);
and U35328 (N_35328,N_33944,N_33090);
xor U35329 (N_35329,N_32766,N_32463);
nor U35330 (N_35330,N_33822,N_32145);
and U35331 (N_35331,N_33963,N_33207);
or U35332 (N_35332,N_33127,N_32811);
and U35333 (N_35333,N_33640,N_33398);
nor U35334 (N_35334,N_32904,N_32173);
and U35335 (N_35335,N_32470,N_32421);
and U35336 (N_35336,N_32455,N_32103);
or U35337 (N_35337,N_33357,N_32679);
nand U35338 (N_35338,N_32032,N_32645);
xor U35339 (N_35339,N_33022,N_33715);
and U35340 (N_35340,N_32320,N_32927);
nand U35341 (N_35341,N_33757,N_32671);
or U35342 (N_35342,N_33415,N_33438);
nor U35343 (N_35343,N_32311,N_33725);
nand U35344 (N_35344,N_32013,N_33784);
nor U35345 (N_35345,N_32076,N_32482);
nand U35346 (N_35346,N_33982,N_32846);
and U35347 (N_35347,N_32220,N_32027);
or U35348 (N_35348,N_32806,N_32031);
nor U35349 (N_35349,N_32114,N_33270);
or U35350 (N_35350,N_33604,N_32133);
nor U35351 (N_35351,N_32266,N_32301);
xor U35352 (N_35352,N_33092,N_33549);
and U35353 (N_35353,N_32429,N_33412);
or U35354 (N_35354,N_32197,N_33502);
or U35355 (N_35355,N_33047,N_33638);
or U35356 (N_35356,N_33716,N_32501);
and U35357 (N_35357,N_33325,N_33182);
nand U35358 (N_35358,N_33015,N_32016);
and U35359 (N_35359,N_33554,N_33884);
or U35360 (N_35360,N_33531,N_33622);
and U35361 (N_35361,N_33619,N_33720);
nor U35362 (N_35362,N_33437,N_32880);
xnor U35363 (N_35363,N_32158,N_32304);
or U35364 (N_35364,N_33947,N_32676);
or U35365 (N_35365,N_33262,N_32978);
nand U35366 (N_35366,N_33332,N_33703);
xnor U35367 (N_35367,N_33167,N_32936);
or U35368 (N_35368,N_33537,N_33259);
nor U35369 (N_35369,N_32827,N_32108);
and U35370 (N_35370,N_32965,N_32958);
nor U35371 (N_35371,N_33149,N_33731);
and U35372 (N_35372,N_33899,N_33944);
nor U35373 (N_35373,N_33219,N_32084);
xnor U35374 (N_35374,N_33463,N_32370);
and U35375 (N_35375,N_33237,N_32309);
nor U35376 (N_35376,N_32673,N_33334);
and U35377 (N_35377,N_33611,N_33468);
nand U35378 (N_35378,N_33314,N_32969);
or U35379 (N_35379,N_32059,N_32644);
and U35380 (N_35380,N_32231,N_33104);
nor U35381 (N_35381,N_32655,N_32489);
nor U35382 (N_35382,N_32009,N_33689);
xnor U35383 (N_35383,N_33071,N_32243);
or U35384 (N_35384,N_33078,N_33836);
xor U35385 (N_35385,N_33353,N_32693);
or U35386 (N_35386,N_32302,N_33308);
or U35387 (N_35387,N_33937,N_33221);
or U35388 (N_35388,N_32143,N_33339);
nor U35389 (N_35389,N_32288,N_33291);
nor U35390 (N_35390,N_33687,N_33294);
nand U35391 (N_35391,N_33859,N_32961);
nor U35392 (N_35392,N_32292,N_32326);
nor U35393 (N_35393,N_33384,N_33532);
or U35394 (N_35394,N_32674,N_33076);
or U35395 (N_35395,N_33770,N_32616);
nor U35396 (N_35396,N_33126,N_33077);
nor U35397 (N_35397,N_32120,N_33690);
or U35398 (N_35398,N_33699,N_32370);
nand U35399 (N_35399,N_33521,N_33254);
nand U35400 (N_35400,N_32342,N_32888);
xnor U35401 (N_35401,N_32496,N_33521);
nor U35402 (N_35402,N_32661,N_32452);
nand U35403 (N_35403,N_33042,N_32755);
nand U35404 (N_35404,N_32740,N_33711);
xor U35405 (N_35405,N_32662,N_32592);
nand U35406 (N_35406,N_33478,N_32119);
nand U35407 (N_35407,N_33638,N_32682);
and U35408 (N_35408,N_32107,N_32846);
and U35409 (N_35409,N_32353,N_32306);
nand U35410 (N_35410,N_32831,N_32554);
and U35411 (N_35411,N_33875,N_32154);
nor U35412 (N_35412,N_33262,N_33831);
and U35413 (N_35413,N_33584,N_32932);
or U35414 (N_35414,N_32203,N_32038);
nand U35415 (N_35415,N_32904,N_32683);
nand U35416 (N_35416,N_32395,N_32280);
or U35417 (N_35417,N_33492,N_32695);
and U35418 (N_35418,N_32027,N_32374);
xor U35419 (N_35419,N_32036,N_32271);
and U35420 (N_35420,N_33439,N_33015);
or U35421 (N_35421,N_32463,N_32681);
and U35422 (N_35422,N_33612,N_32627);
nand U35423 (N_35423,N_33878,N_33333);
and U35424 (N_35424,N_32299,N_32350);
xor U35425 (N_35425,N_32183,N_33233);
nand U35426 (N_35426,N_32901,N_33538);
and U35427 (N_35427,N_33921,N_32042);
or U35428 (N_35428,N_33999,N_32073);
nor U35429 (N_35429,N_33468,N_33579);
and U35430 (N_35430,N_32391,N_32102);
or U35431 (N_35431,N_32668,N_32805);
or U35432 (N_35432,N_32817,N_32174);
xnor U35433 (N_35433,N_33062,N_33806);
xor U35434 (N_35434,N_32165,N_33989);
xnor U35435 (N_35435,N_33087,N_32907);
and U35436 (N_35436,N_33833,N_33037);
nor U35437 (N_35437,N_32791,N_32272);
xor U35438 (N_35438,N_33090,N_33361);
xor U35439 (N_35439,N_33691,N_33442);
and U35440 (N_35440,N_32148,N_33687);
nand U35441 (N_35441,N_33537,N_33816);
xor U35442 (N_35442,N_32205,N_32772);
nand U35443 (N_35443,N_32447,N_32423);
nand U35444 (N_35444,N_32343,N_33118);
xnor U35445 (N_35445,N_33689,N_32636);
nand U35446 (N_35446,N_32823,N_33300);
and U35447 (N_35447,N_32688,N_33887);
nand U35448 (N_35448,N_32786,N_32325);
xor U35449 (N_35449,N_33266,N_32574);
and U35450 (N_35450,N_32982,N_33915);
and U35451 (N_35451,N_33129,N_32849);
nor U35452 (N_35452,N_32449,N_33105);
and U35453 (N_35453,N_32766,N_32142);
or U35454 (N_35454,N_32748,N_33966);
nor U35455 (N_35455,N_33823,N_32336);
nand U35456 (N_35456,N_32449,N_32181);
nor U35457 (N_35457,N_33202,N_33750);
or U35458 (N_35458,N_33371,N_32029);
nand U35459 (N_35459,N_33249,N_32281);
xnor U35460 (N_35460,N_33514,N_33337);
and U35461 (N_35461,N_32649,N_33837);
nand U35462 (N_35462,N_33215,N_32690);
or U35463 (N_35463,N_33592,N_32939);
and U35464 (N_35464,N_32693,N_32432);
nand U35465 (N_35465,N_32856,N_33087);
xnor U35466 (N_35466,N_33086,N_32959);
or U35467 (N_35467,N_32849,N_33275);
xor U35468 (N_35468,N_32819,N_33986);
xnor U35469 (N_35469,N_33307,N_32123);
or U35470 (N_35470,N_33126,N_32450);
and U35471 (N_35471,N_33742,N_33996);
nor U35472 (N_35472,N_33504,N_33949);
nand U35473 (N_35473,N_33049,N_33125);
nor U35474 (N_35474,N_33878,N_33294);
xnor U35475 (N_35475,N_33507,N_33131);
or U35476 (N_35476,N_33747,N_32082);
nand U35477 (N_35477,N_32201,N_32424);
or U35478 (N_35478,N_33135,N_32975);
nand U35479 (N_35479,N_32658,N_33786);
or U35480 (N_35480,N_32860,N_33414);
nor U35481 (N_35481,N_32059,N_32878);
xnor U35482 (N_35482,N_32708,N_32973);
and U35483 (N_35483,N_32428,N_32696);
nand U35484 (N_35484,N_32031,N_32938);
or U35485 (N_35485,N_32737,N_32931);
nand U35486 (N_35486,N_32845,N_32049);
or U35487 (N_35487,N_32290,N_32555);
nand U35488 (N_35488,N_33220,N_32205);
nand U35489 (N_35489,N_32986,N_33166);
nor U35490 (N_35490,N_32413,N_33122);
nand U35491 (N_35491,N_33388,N_32432);
or U35492 (N_35492,N_32523,N_32333);
and U35493 (N_35493,N_33823,N_32549);
or U35494 (N_35494,N_33159,N_33996);
and U35495 (N_35495,N_33914,N_32094);
nand U35496 (N_35496,N_32149,N_32619);
nand U35497 (N_35497,N_33200,N_33418);
and U35498 (N_35498,N_33278,N_33746);
nand U35499 (N_35499,N_33257,N_32629);
nand U35500 (N_35500,N_32949,N_32921);
nand U35501 (N_35501,N_32565,N_32695);
or U35502 (N_35502,N_33531,N_32564);
and U35503 (N_35503,N_32285,N_33989);
nor U35504 (N_35504,N_33871,N_32800);
nand U35505 (N_35505,N_32847,N_33731);
nand U35506 (N_35506,N_33521,N_33631);
and U35507 (N_35507,N_33706,N_32041);
nand U35508 (N_35508,N_32095,N_33797);
or U35509 (N_35509,N_32903,N_32542);
nand U35510 (N_35510,N_32424,N_33398);
xor U35511 (N_35511,N_33275,N_32152);
or U35512 (N_35512,N_32410,N_32134);
and U35513 (N_35513,N_32158,N_33213);
or U35514 (N_35514,N_33571,N_32812);
nor U35515 (N_35515,N_32754,N_33388);
nand U35516 (N_35516,N_32601,N_32577);
and U35517 (N_35517,N_33385,N_32120);
and U35518 (N_35518,N_33372,N_32729);
xnor U35519 (N_35519,N_33965,N_32824);
xnor U35520 (N_35520,N_32647,N_32033);
or U35521 (N_35521,N_32532,N_33440);
nor U35522 (N_35522,N_32992,N_32657);
or U35523 (N_35523,N_32285,N_32457);
nand U35524 (N_35524,N_32950,N_33694);
or U35525 (N_35525,N_32801,N_32986);
nand U35526 (N_35526,N_32082,N_32461);
nor U35527 (N_35527,N_32014,N_33059);
or U35528 (N_35528,N_32084,N_32150);
and U35529 (N_35529,N_32741,N_32314);
xnor U35530 (N_35530,N_33935,N_32168);
nand U35531 (N_35531,N_33347,N_32409);
or U35532 (N_35532,N_32009,N_33975);
and U35533 (N_35533,N_33089,N_32883);
and U35534 (N_35534,N_33024,N_33283);
xnor U35535 (N_35535,N_33438,N_33675);
xor U35536 (N_35536,N_33268,N_32740);
nand U35537 (N_35537,N_33757,N_33145);
xnor U35538 (N_35538,N_32075,N_32027);
or U35539 (N_35539,N_33776,N_32000);
xor U35540 (N_35540,N_33622,N_33472);
xor U35541 (N_35541,N_33891,N_32134);
nand U35542 (N_35542,N_33954,N_33705);
nor U35543 (N_35543,N_33662,N_32116);
nand U35544 (N_35544,N_32636,N_33021);
and U35545 (N_35545,N_32800,N_32923);
or U35546 (N_35546,N_32283,N_32331);
or U35547 (N_35547,N_32766,N_32461);
xnor U35548 (N_35548,N_32790,N_32477);
nand U35549 (N_35549,N_32807,N_32692);
nand U35550 (N_35550,N_33530,N_33803);
nor U35551 (N_35551,N_33208,N_32435);
or U35552 (N_35552,N_33308,N_32813);
and U35553 (N_35553,N_33365,N_32389);
or U35554 (N_35554,N_32920,N_33002);
and U35555 (N_35555,N_33287,N_32324);
xor U35556 (N_35556,N_32677,N_32905);
or U35557 (N_35557,N_32803,N_32115);
or U35558 (N_35558,N_33114,N_32147);
or U35559 (N_35559,N_32913,N_32063);
or U35560 (N_35560,N_33624,N_33716);
or U35561 (N_35561,N_32382,N_32268);
and U35562 (N_35562,N_32963,N_33595);
and U35563 (N_35563,N_32454,N_33469);
nand U35564 (N_35564,N_32967,N_33913);
or U35565 (N_35565,N_33539,N_33799);
xnor U35566 (N_35566,N_32130,N_33566);
nor U35567 (N_35567,N_33847,N_33955);
and U35568 (N_35568,N_33053,N_33716);
xor U35569 (N_35569,N_32605,N_32714);
nand U35570 (N_35570,N_33398,N_33773);
nor U35571 (N_35571,N_33288,N_32562);
and U35572 (N_35572,N_32732,N_32710);
xor U35573 (N_35573,N_32764,N_32928);
and U35574 (N_35574,N_33597,N_33453);
or U35575 (N_35575,N_32698,N_33162);
nand U35576 (N_35576,N_33065,N_33784);
and U35577 (N_35577,N_33126,N_32036);
nor U35578 (N_35578,N_32774,N_32826);
and U35579 (N_35579,N_32103,N_33124);
nor U35580 (N_35580,N_33435,N_32101);
and U35581 (N_35581,N_33009,N_33272);
or U35582 (N_35582,N_33517,N_33800);
and U35583 (N_35583,N_32755,N_32800);
nand U35584 (N_35584,N_33074,N_33669);
nor U35585 (N_35585,N_32881,N_33034);
nand U35586 (N_35586,N_32446,N_33848);
xor U35587 (N_35587,N_33351,N_32497);
xnor U35588 (N_35588,N_33128,N_33056);
and U35589 (N_35589,N_33583,N_32424);
nand U35590 (N_35590,N_32680,N_32341);
xor U35591 (N_35591,N_32890,N_32468);
and U35592 (N_35592,N_32120,N_33350);
nor U35593 (N_35593,N_32783,N_32423);
or U35594 (N_35594,N_33925,N_32949);
or U35595 (N_35595,N_33200,N_32555);
and U35596 (N_35596,N_33042,N_33579);
nor U35597 (N_35597,N_32235,N_33309);
xnor U35598 (N_35598,N_32587,N_33277);
xor U35599 (N_35599,N_32712,N_32669);
or U35600 (N_35600,N_33617,N_33975);
nor U35601 (N_35601,N_32938,N_32416);
or U35602 (N_35602,N_32658,N_33168);
and U35603 (N_35603,N_33235,N_32114);
nand U35604 (N_35604,N_33418,N_32436);
nor U35605 (N_35605,N_33040,N_32800);
and U35606 (N_35606,N_32628,N_33372);
xnor U35607 (N_35607,N_32990,N_32516);
or U35608 (N_35608,N_32815,N_33453);
xnor U35609 (N_35609,N_33157,N_33595);
nor U35610 (N_35610,N_33105,N_33707);
and U35611 (N_35611,N_32926,N_33921);
or U35612 (N_35612,N_32084,N_32281);
nand U35613 (N_35613,N_33795,N_33981);
or U35614 (N_35614,N_32273,N_33613);
nor U35615 (N_35615,N_33205,N_33754);
nand U35616 (N_35616,N_33121,N_32192);
or U35617 (N_35617,N_33058,N_33465);
nor U35618 (N_35618,N_32236,N_33642);
nor U35619 (N_35619,N_32408,N_32118);
or U35620 (N_35620,N_32025,N_32393);
or U35621 (N_35621,N_32326,N_32879);
xor U35622 (N_35622,N_32525,N_32972);
nor U35623 (N_35623,N_33249,N_33471);
nor U35624 (N_35624,N_32634,N_32276);
and U35625 (N_35625,N_33211,N_33394);
nor U35626 (N_35626,N_32122,N_33664);
and U35627 (N_35627,N_33301,N_32178);
nand U35628 (N_35628,N_32544,N_32862);
xnor U35629 (N_35629,N_32005,N_33704);
or U35630 (N_35630,N_33601,N_33962);
xor U35631 (N_35631,N_32712,N_32496);
xor U35632 (N_35632,N_33517,N_32487);
nor U35633 (N_35633,N_32998,N_33951);
nand U35634 (N_35634,N_33153,N_33986);
xor U35635 (N_35635,N_32831,N_32867);
or U35636 (N_35636,N_32627,N_32143);
xor U35637 (N_35637,N_33478,N_32441);
nor U35638 (N_35638,N_32997,N_33883);
and U35639 (N_35639,N_32026,N_33457);
xnor U35640 (N_35640,N_33380,N_32818);
nand U35641 (N_35641,N_33804,N_32812);
or U35642 (N_35642,N_33897,N_32267);
xor U35643 (N_35643,N_32888,N_33363);
nor U35644 (N_35644,N_32933,N_33753);
and U35645 (N_35645,N_33728,N_32131);
nand U35646 (N_35646,N_32336,N_32348);
or U35647 (N_35647,N_32898,N_33649);
nor U35648 (N_35648,N_33017,N_33085);
nand U35649 (N_35649,N_33318,N_32786);
or U35650 (N_35650,N_32519,N_32020);
and U35651 (N_35651,N_32456,N_32747);
or U35652 (N_35652,N_33315,N_33186);
or U35653 (N_35653,N_33779,N_33489);
and U35654 (N_35654,N_33101,N_32860);
and U35655 (N_35655,N_32156,N_33561);
nand U35656 (N_35656,N_33648,N_32425);
xnor U35657 (N_35657,N_32468,N_33116);
nor U35658 (N_35658,N_33722,N_33220);
xor U35659 (N_35659,N_33872,N_32893);
xnor U35660 (N_35660,N_32861,N_32074);
nor U35661 (N_35661,N_32800,N_33297);
and U35662 (N_35662,N_33162,N_32352);
nand U35663 (N_35663,N_32401,N_32649);
nand U35664 (N_35664,N_32509,N_33212);
or U35665 (N_35665,N_33424,N_32251);
nand U35666 (N_35666,N_33297,N_32188);
xnor U35667 (N_35667,N_33592,N_32219);
nor U35668 (N_35668,N_32356,N_32421);
or U35669 (N_35669,N_32028,N_32742);
nand U35670 (N_35670,N_33714,N_33879);
nand U35671 (N_35671,N_32085,N_32967);
nand U35672 (N_35672,N_33180,N_32742);
nand U35673 (N_35673,N_33746,N_32240);
nor U35674 (N_35674,N_32359,N_32844);
nor U35675 (N_35675,N_33225,N_33506);
or U35676 (N_35676,N_33176,N_33211);
or U35677 (N_35677,N_33384,N_33536);
and U35678 (N_35678,N_33266,N_33260);
and U35679 (N_35679,N_33324,N_32634);
xor U35680 (N_35680,N_32326,N_32673);
xor U35681 (N_35681,N_33670,N_33401);
nand U35682 (N_35682,N_33701,N_33897);
xnor U35683 (N_35683,N_32301,N_33885);
or U35684 (N_35684,N_33169,N_32686);
nand U35685 (N_35685,N_33389,N_33579);
nand U35686 (N_35686,N_33223,N_32197);
nor U35687 (N_35687,N_32414,N_33108);
xnor U35688 (N_35688,N_32304,N_32370);
or U35689 (N_35689,N_33375,N_33393);
nand U35690 (N_35690,N_32178,N_33197);
xnor U35691 (N_35691,N_32418,N_33356);
xor U35692 (N_35692,N_32869,N_33196);
and U35693 (N_35693,N_33211,N_33087);
nand U35694 (N_35694,N_33446,N_32527);
nand U35695 (N_35695,N_32116,N_32955);
nand U35696 (N_35696,N_33025,N_32280);
nor U35697 (N_35697,N_32078,N_32867);
xor U35698 (N_35698,N_32612,N_33703);
or U35699 (N_35699,N_32527,N_32251);
nand U35700 (N_35700,N_33729,N_32278);
or U35701 (N_35701,N_33145,N_33823);
xnor U35702 (N_35702,N_32615,N_33866);
xor U35703 (N_35703,N_33779,N_32782);
and U35704 (N_35704,N_33610,N_33840);
nor U35705 (N_35705,N_32798,N_32634);
nand U35706 (N_35706,N_32208,N_33769);
and U35707 (N_35707,N_32957,N_32894);
or U35708 (N_35708,N_33952,N_33559);
or U35709 (N_35709,N_33606,N_32805);
nand U35710 (N_35710,N_32122,N_33907);
or U35711 (N_35711,N_33890,N_32392);
nor U35712 (N_35712,N_32154,N_33206);
xor U35713 (N_35713,N_33727,N_33700);
and U35714 (N_35714,N_32292,N_33253);
xor U35715 (N_35715,N_32288,N_33145);
or U35716 (N_35716,N_32530,N_32600);
xor U35717 (N_35717,N_33650,N_33443);
or U35718 (N_35718,N_33187,N_32480);
xor U35719 (N_35719,N_33515,N_33487);
xor U35720 (N_35720,N_32632,N_32354);
and U35721 (N_35721,N_32647,N_33899);
nor U35722 (N_35722,N_33091,N_32605);
nand U35723 (N_35723,N_33869,N_33910);
or U35724 (N_35724,N_33108,N_33627);
nor U35725 (N_35725,N_33483,N_33041);
or U35726 (N_35726,N_32669,N_33134);
nor U35727 (N_35727,N_32590,N_33716);
nor U35728 (N_35728,N_33266,N_32498);
nor U35729 (N_35729,N_33759,N_32697);
and U35730 (N_35730,N_33929,N_32885);
nand U35731 (N_35731,N_32917,N_32269);
and U35732 (N_35732,N_32999,N_32746);
nand U35733 (N_35733,N_32424,N_32065);
and U35734 (N_35734,N_32402,N_32011);
and U35735 (N_35735,N_33947,N_33245);
nand U35736 (N_35736,N_32392,N_32009);
xor U35737 (N_35737,N_32741,N_32235);
nand U35738 (N_35738,N_32804,N_32795);
xor U35739 (N_35739,N_32213,N_33320);
nand U35740 (N_35740,N_33315,N_33999);
xnor U35741 (N_35741,N_32788,N_33284);
nor U35742 (N_35742,N_33162,N_33413);
xnor U35743 (N_35743,N_33073,N_32858);
or U35744 (N_35744,N_33980,N_32861);
or U35745 (N_35745,N_32680,N_33480);
or U35746 (N_35746,N_33650,N_32476);
nand U35747 (N_35747,N_32867,N_33184);
and U35748 (N_35748,N_32848,N_32326);
nand U35749 (N_35749,N_32275,N_32251);
nor U35750 (N_35750,N_33725,N_33346);
and U35751 (N_35751,N_33639,N_33666);
nor U35752 (N_35752,N_32663,N_33835);
and U35753 (N_35753,N_32400,N_32670);
xor U35754 (N_35754,N_32995,N_32338);
nor U35755 (N_35755,N_32244,N_32686);
nor U35756 (N_35756,N_33310,N_33093);
nand U35757 (N_35757,N_33372,N_32775);
or U35758 (N_35758,N_32993,N_33683);
nor U35759 (N_35759,N_33449,N_33935);
nand U35760 (N_35760,N_33671,N_32608);
nand U35761 (N_35761,N_32162,N_32491);
or U35762 (N_35762,N_33266,N_33388);
xnor U35763 (N_35763,N_33488,N_32352);
nand U35764 (N_35764,N_33619,N_33877);
or U35765 (N_35765,N_33837,N_32274);
nor U35766 (N_35766,N_32605,N_32483);
xnor U35767 (N_35767,N_33416,N_32193);
nand U35768 (N_35768,N_32456,N_32279);
and U35769 (N_35769,N_32141,N_32121);
and U35770 (N_35770,N_33633,N_33381);
xnor U35771 (N_35771,N_33031,N_32151);
xor U35772 (N_35772,N_32609,N_32909);
nor U35773 (N_35773,N_33225,N_32834);
or U35774 (N_35774,N_32162,N_32240);
xnor U35775 (N_35775,N_32044,N_33172);
nor U35776 (N_35776,N_32587,N_32182);
and U35777 (N_35777,N_33890,N_32911);
xor U35778 (N_35778,N_33097,N_33588);
nor U35779 (N_35779,N_33177,N_33646);
and U35780 (N_35780,N_32992,N_33763);
xor U35781 (N_35781,N_32729,N_33641);
nor U35782 (N_35782,N_33016,N_32564);
and U35783 (N_35783,N_33142,N_32362);
xor U35784 (N_35784,N_33373,N_33758);
nand U35785 (N_35785,N_33304,N_32530);
nand U35786 (N_35786,N_32364,N_32432);
xnor U35787 (N_35787,N_32094,N_32338);
nand U35788 (N_35788,N_33646,N_33745);
or U35789 (N_35789,N_32732,N_32153);
nand U35790 (N_35790,N_33102,N_32655);
nor U35791 (N_35791,N_32819,N_32003);
nor U35792 (N_35792,N_33204,N_33011);
and U35793 (N_35793,N_32439,N_33439);
xor U35794 (N_35794,N_32329,N_33538);
xnor U35795 (N_35795,N_32827,N_33841);
or U35796 (N_35796,N_33325,N_33736);
nor U35797 (N_35797,N_32716,N_32170);
xnor U35798 (N_35798,N_33165,N_33467);
nor U35799 (N_35799,N_33964,N_32002);
and U35800 (N_35800,N_32372,N_32956);
nor U35801 (N_35801,N_32820,N_33036);
xnor U35802 (N_35802,N_32201,N_32159);
or U35803 (N_35803,N_32004,N_33710);
and U35804 (N_35804,N_33253,N_32632);
xor U35805 (N_35805,N_33832,N_32195);
nor U35806 (N_35806,N_33321,N_33713);
xnor U35807 (N_35807,N_33737,N_32585);
nand U35808 (N_35808,N_32484,N_32432);
xnor U35809 (N_35809,N_32202,N_33311);
or U35810 (N_35810,N_33800,N_32778);
and U35811 (N_35811,N_33683,N_32012);
or U35812 (N_35812,N_33280,N_32007);
or U35813 (N_35813,N_32020,N_32159);
xnor U35814 (N_35814,N_32937,N_33050);
nand U35815 (N_35815,N_32599,N_32346);
and U35816 (N_35816,N_33311,N_32888);
nor U35817 (N_35817,N_32028,N_32394);
and U35818 (N_35818,N_33764,N_32308);
and U35819 (N_35819,N_32079,N_33172);
and U35820 (N_35820,N_32652,N_32681);
or U35821 (N_35821,N_32644,N_32377);
or U35822 (N_35822,N_32274,N_32579);
nand U35823 (N_35823,N_32068,N_32166);
xnor U35824 (N_35824,N_33742,N_33782);
and U35825 (N_35825,N_32978,N_33932);
nor U35826 (N_35826,N_33126,N_32424);
nand U35827 (N_35827,N_32358,N_32076);
xor U35828 (N_35828,N_33605,N_32754);
and U35829 (N_35829,N_33839,N_32410);
nand U35830 (N_35830,N_33018,N_32434);
or U35831 (N_35831,N_33387,N_33298);
nand U35832 (N_35832,N_33629,N_32808);
and U35833 (N_35833,N_32152,N_33311);
or U35834 (N_35834,N_32170,N_33363);
or U35835 (N_35835,N_33347,N_32299);
xnor U35836 (N_35836,N_32135,N_32641);
nand U35837 (N_35837,N_33437,N_33944);
or U35838 (N_35838,N_33545,N_32521);
xor U35839 (N_35839,N_33672,N_32736);
nand U35840 (N_35840,N_33665,N_32512);
nor U35841 (N_35841,N_33079,N_32068);
xnor U35842 (N_35842,N_33978,N_32296);
nor U35843 (N_35843,N_32545,N_33889);
and U35844 (N_35844,N_33468,N_32278);
or U35845 (N_35845,N_33457,N_32080);
or U35846 (N_35846,N_33627,N_32102);
nand U35847 (N_35847,N_32736,N_33894);
or U35848 (N_35848,N_32397,N_33031);
nor U35849 (N_35849,N_33187,N_33031);
and U35850 (N_35850,N_33725,N_32064);
or U35851 (N_35851,N_32607,N_32919);
nand U35852 (N_35852,N_32652,N_32264);
or U35853 (N_35853,N_32857,N_32477);
or U35854 (N_35854,N_32980,N_32707);
or U35855 (N_35855,N_33876,N_32761);
nand U35856 (N_35856,N_33683,N_33997);
xnor U35857 (N_35857,N_32803,N_32884);
and U35858 (N_35858,N_32665,N_33174);
and U35859 (N_35859,N_33821,N_33547);
xnor U35860 (N_35860,N_33526,N_32606);
and U35861 (N_35861,N_33302,N_32156);
or U35862 (N_35862,N_33571,N_33987);
nand U35863 (N_35863,N_32307,N_32250);
and U35864 (N_35864,N_32795,N_33160);
nor U35865 (N_35865,N_33850,N_32925);
or U35866 (N_35866,N_33813,N_33399);
or U35867 (N_35867,N_33920,N_32046);
nand U35868 (N_35868,N_32126,N_33408);
xor U35869 (N_35869,N_33843,N_32173);
or U35870 (N_35870,N_32553,N_33034);
nand U35871 (N_35871,N_33973,N_32011);
nand U35872 (N_35872,N_32710,N_33100);
or U35873 (N_35873,N_32976,N_32992);
and U35874 (N_35874,N_32161,N_32068);
or U35875 (N_35875,N_33352,N_33737);
or U35876 (N_35876,N_33947,N_33344);
nor U35877 (N_35877,N_33075,N_33947);
nand U35878 (N_35878,N_32456,N_32854);
nor U35879 (N_35879,N_33855,N_32911);
xnor U35880 (N_35880,N_33704,N_33827);
or U35881 (N_35881,N_33134,N_32698);
nand U35882 (N_35882,N_32596,N_32689);
and U35883 (N_35883,N_32742,N_33655);
or U35884 (N_35884,N_32757,N_32414);
and U35885 (N_35885,N_32039,N_32816);
nor U35886 (N_35886,N_32313,N_32559);
xor U35887 (N_35887,N_33386,N_33018);
nand U35888 (N_35888,N_33199,N_32394);
xnor U35889 (N_35889,N_33371,N_32493);
xnor U35890 (N_35890,N_33636,N_32770);
nor U35891 (N_35891,N_33505,N_32016);
xor U35892 (N_35892,N_32071,N_32646);
nor U35893 (N_35893,N_33954,N_32096);
nor U35894 (N_35894,N_33187,N_33610);
xnor U35895 (N_35895,N_33382,N_33194);
nor U35896 (N_35896,N_32848,N_33096);
nor U35897 (N_35897,N_32256,N_33157);
nand U35898 (N_35898,N_33273,N_33242);
or U35899 (N_35899,N_33887,N_33067);
xor U35900 (N_35900,N_33839,N_33543);
xor U35901 (N_35901,N_33740,N_32708);
nor U35902 (N_35902,N_32604,N_33661);
nor U35903 (N_35903,N_33960,N_32024);
and U35904 (N_35904,N_32349,N_33284);
or U35905 (N_35905,N_32889,N_33363);
or U35906 (N_35906,N_33283,N_32216);
xor U35907 (N_35907,N_33699,N_32063);
xor U35908 (N_35908,N_33688,N_33676);
nand U35909 (N_35909,N_33634,N_32828);
and U35910 (N_35910,N_33406,N_33260);
and U35911 (N_35911,N_32257,N_32241);
nand U35912 (N_35912,N_33384,N_33185);
or U35913 (N_35913,N_33975,N_33113);
or U35914 (N_35914,N_33764,N_32612);
nand U35915 (N_35915,N_33227,N_32977);
nor U35916 (N_35916,N_33121,N_32187);
nor U35917 (N_35917,N_33853,N_33752);
xnor U35918 (N_35918,N_33023,N_32374);
or U35919 (N_35919,N_33938,N_33626);
and U35920 (N_35920,N_33161,N_33922);
xnor U35921 (N_35921,N_33153,N_33938);
or U35922 (N_35922,N_32453,N_33001);
nand U35923 (N_35923,N_33561,N_33103);
or U35924 (N_35924,N_33066,N_32739);
or U35925 (N_35925,N_32182,N_33938);
nor U35926 (N_35926,N_32010,N_33298);
xnor U35927 (N_35927,N_33282,N_32860);
nand U35928 (N_35928,N_32772,N_32439);
xor U35929 (N_35929,N_33847,N_33350);
xor U35930 (N_35930,N_33754,N_33956);
xnor U35931 (N_35931,N_32939,N_32876);
nand U35932 (N_35932,N_32089,N_33242);
nor U35933 (N_35933,N_33797,N_33650);
or U35934 (N_35934,N_33724,N_32786);
nor U35935 (N_35935,N_33938,N_32253);
nand U35936 (N_35936,N_32465,N_33547);
and U35937 (N_35937,N_33281,N_33962);
nor U35938 (N_35938,N_32943,N_32635);
or U35939 (N_35939,N_32575,N_33181);
nor U35940 (N_35940,N_33915,N_32828);
nand U35941 (N_35941,N_33420,N_33429);
nor U35942 (N_35942,N_32765,N_33434);
nor U35943 (N_35943,N_33573,N_33115);
xnor U35944 (N_35944,N_32240,N_32696);
and U35945 (N_35945,N_32903,N_33119);
and U35946 (N_35946,N_32043,N_32634);
xnor U35947 (N_35947,N_32050,N_32362);
and U35948 (N_35948,N_32796,N_33819);
and U35949 (N_35949,N_33284,N_32614);
xor U35950 (N_35950,N_32758,N_33651);
xnor U35951 (N_35951,N_32338,N_33019);
nor U35952 (N_35952,N_32208,N_32152);
nor U35953 (N_35953,N_33091,N_33050);
and U35954 (N_35954,N_32271,N_32241);
and U35955 (N_35955,N_33033,N_32067);
nand U35956 (N_35956,N_33522,N_32098);
and U35957 (N_35957,N_32559,N_32642);
xnor U35958 (N_35958,N_32334,N_33179);
xnor U35959 (N_35959,N_32162,N_33214);
and U35960 (N_35960,N_33710,N_33959);
or U35961 (N_35961,N_32608,N_32333);
or U35962 (N_35962,N_33054,N_32454);
nand U35963 (N_35963,N_32097,N_33389);
nor U35964 (N_35964,N_32108,N_32306);
nor U35965 (N_35965,N_33003,N_32487);
xnor U35966 (N_35966,N_32425,N_33501);
or U35967 (N_35967,N_33301,N_33534);
or U35968 (N_35968,N_32620,N_33080);
nor U35969 (N_35969,N_33946,N_32611);
or U35970 (N_35970,N_32831,N_32568);
or U35971 (N_35971,N_33613,N_32372);
and U35972 (N_35972,N_32536,N_33755);
and U35973 (N_35973,N_32738,N_33155);
or U35974 (N_35974,N_33274,N_32356);
nor U35975 (N_35975,N_33681,N_32363);
nand U35976 (N_35976,N_33167,N_33317);
nand U35977 (N_35977,N_33157,N_32163);
nand U35978 (N_35978,N_32683,N_32939);
and U35979 (N_35979,N_33000,N_33488);
and U35980 (N_35980,N_32031,N_33088);
or U35981 (N_35981,N_32176,N_33657);
xor U35982 (N_35982,N_33232,N_33038);
and U35983 (N_35983,N_32353,N_32474);
or U35984 (N_35984,N_33989,N_32595);
nor U35985 (N_35985,N_33156,N_32061);
nor U35986 (N_35986,N_33255,N_32874);
and U35987 (N_35987,N_32101,N_32388);
nor U35988 (N_35988,N_33746,N_33972);
nand U35989 (N_35989,N_33159,N_33780);
xor U35990 (N_35990,N_33737,N_33748);
nor U35991 (N_35991,N_32394,N_32219);
and U35992 (N_35992,N_33449,N_32330);
xnor U35993 (N_35993,N_33759,N_33767);
or U35994 (N_35994,N_33240,N_32553);
or U35995 (N_35995,N_33065,N_32167);
and U35996 (N_35996,N_33545,N_33158);
nor U35997 (N_35997,N_32309,N_33947);
and U35998 (N_35998,N_33881,N_32320);
or U35999 (N_35999,N_32422,N_32294);
or U36000 (N_36000,N_34276,N_34546);
nand U36001 (N_36001,N_35917,N_34318);
xnor U36002 (N_36002,N_34360,N_35200);
nand U36003 (N_36003,N_34545,N_35783);
nor U36004 (N_36004,N_35034,N_35302);
xor U36005 (N_36005,N_34508,N_34895);
nand U36006 (N_36006,N_35657,N_34478);
xnor U36007 (N_36007,N_35022,N_35148);
nand U36008 (N_36008,N_35590,N_34373);
nor U36009 (N_36009,N_34523,N_35080);
nor U36010 (N_36010,N_34389,N_35384);
and U36011 (N_36011,N_35611,N_35266);
and U36012 (N_36012,N_34042,N_34942);
and U36013 (N_36013,N_35416,N_34715);
nand U36014 (N_36014,N_35788,N_34981);
nand U36015 (N_36015,N_35735,N_35252);
or U36016 (N_36016,N_35599,N_35125);
nor U36017 (N_36017,N_34149,N_34842);
or U36018 (N_36018,N_34882,N_34954);
or U36019 (N_36019,N_35988,N_34815);
nand U36020 (N_36020,N_34049,N_35989);
nand U36021 (N_36021,N_35708,N_34885);
nor U36022 (N_36022,N_34745,N_34470);
nor U36023 (N_36023,N_35824,N_34316);
xor U36024 (N_36024,N_35545,N_35315);
xor U36025 (N_36025,N_35334,N_34232);
nor U36026 (N_36026,N_35380,N_35793);
or U36027 (N_36027,N_34703,N_35679);
xnor U36028 (N_36028,N_35636,N_34811);
or U36029 (N_36029,N_34314,N_35616);
xor U36030 (N_36030,N_35860,N_35674);
xnor U36031 (N_36031,N_35179,N_35748);
or U36032 (N_36032,N_35591,N_35362);
xnor U36033 (N_36033,N_34940,N_35254);
nor U36034 (N_36034,N_34767,N_34562);
nand U36035 (N_36035,N_35291,N_35688);
nand U36036 (N_36036,N_35109,N_35535);
or U36037 (N_36037,N_35364,N_35191);
nand U36038 (N_36038,N_34972,N_34688);
and U36039 (N_36039,N_34177,N_34900);
nand U36040 (N_36040,N_35320,N_34302);
or U36041 (N_36041,N_34576,N_34266);
xor U36042 (N_36042,N_34747,N_34740);
and U36043 (N_36043,N_34469,N_35622);
and U36044 (N_36044,N_34691,N_34979);
nor U36045 (N_36045,N_35668,N_35787);
nand U36046 (N_36046,N_34072,N_35289);
nor U36047 (N_36047,N_34084,N_34456);
nor U36048 (N_36048,N_34352,N_34939);
xnor U36049 (N_36049,N_34629,N_34994);
nand U36050 (N_36050,N_34825,N_35300);
nor U36051 (N_36051,N_35982,N_34350);
or U36052 (N_36052,N_34174,N_35099);
and U36053 (N_36053,N_35028,N_35702);
and U36054 (N_36054,N_35634,N_35175);
or U36055 (N_36055,N_35219,N_34911);
and U36056 (N_36056,N_34856,N_34609);
nor U36057 (N_36057,N_35003,N_34116);
and U36058 (N_36058,N_34099,N_34261);
nand U36059 (N_36059,N_35001,N_35533);
nor U36060 (N_36060,N_35117,N_34441);
and U36061 (N_36061,N_35373,N_35999);
xor U36062 (N_36062,N_35433,N_35817);
nand U36063 (N_36063,N_34264,N_34066);
and U36064 (N_36064,N_35184,N_34887);
nor U36065 (N_36065,N_34105,N_34356);
nor U36066 (N_36066,N_34085,N_35934);
or U36067 (N_36067,N_35138,N_35071);
nor U36068 (N_36068,N_34847,N_35186);
nor U36069 (N_36069,N_35621,N_35163);
nand U36070 (N_36070,N_34416,N_34556);
nand U36071 (N_36071,N_34604,N_34566);
nand U36072 (N_36072,N_35531,N_35556);
or U36073 (N_36073,N_34769,N_34383);
xor U36074 (N_36074,N_35995,N_35948);
xor U36075 (N_36075,N_35093,N_35906);
xnor U36076 (N_36076,N_35007,N_34018);
nor U36077 (N_36077,N_35875,N_35804);
nand U36078 (N_36078,N_35346,N_34182);
nand U36079 (N_36079,N_34259,N_34789);
nor U36080 (N_36080,N_35032,N_34748);
nor U36081 (N_36081,N_35638,N_34283);
nand U36082 (N_36082,N_34484,N_35511);
xnor U36083 (N_36083,N_35724,N_35505);
or U36084 (N_36084,N_35968,N_35253);
nand U36085 (N_36085,N_35974,N_35276);
or U36086 (N_36086,N_34439,N_34152);
nand U36087 (N_36087,N_34357,N_34509);
nand U36088 (N_36088,N_34600,N_35810);
nand U36089 (N_36089,N_34483,N_34069);
xnor U36090 (N_36090,N_34025,N_35950);
nand U36091 (N_36091,N_35446,N_35233);
or U36092 (N_36092,N_34479,N_35976);
and U36093 (N_36093,N_34824,N_35108);
nor U36094 (N_36094,N_34423,N_34067);
xnor U36095 (N_36095,N_34570,N_34231);
xnor U36096 (N_36096,N_34816,N_34466);
or U36097 (N_36097,N_34550,N_34644);
nor U36098 (N_36098,N_34985,N_34662);
nand U36099 (N_36099,N_35326,N_35789);
and U36100 (N_36100,N_35197,N_34502);
nand U36101 (N_36101,N_34928,N_34415);
or U36102 (N_36102,N_35835,N_34068);
nand U36103 (N_36103,N_35297,N_34388);
or U36104 (N_36104,N_35943,N_34557);
or U36105 (N_36105,N_35360,N_35414);
xnor U36106 (N_36106,N_35514,N_35274);
and U36107 (N_36107,N_35598,N_35110);
and U36108 (N_36108,N_34201,N_34866);
xnor U36109 (N_36109,N_34516,N_34390);
nand U36110 (N_36110,N_35085,N_35541);
nand U36111 (N_36111,N_34327,N_35623);
or U36112 (N_36112,N_35872,N_35825);
or U36113 (N_36113,N_34980,N_34317);
nand U36114 (N_36114,N_34967,N_35229);
nand U36115 (N_36115,N_34250,N_35617);
and U36116 (N_36116,N_34706,N_34737);
nand U36117 (N_36117,N_35717,N_34658);
nor U36118 (N_36118,N_35646,N_35651);
xnor U36119 (N_36119,N_34473,N_35303);
nor U36120 (N_36120,N_34392,N_34973);
xor U36121 (N_36121,N_35418,N_35500);
xnor U36122 (N_36122,N_35056,N_35595);
nand U36123 (N_36123,N_35162,N_34238);
and U36124 (N_36124,N_35035,N_34716);
and U36125 (N_36125,N_34809,N_35673);
nand U36126 (N_36126,N_35236,N_34634);
nand U36127 (N_36127,N_35911,N_35070);
or U36128 (N_36128,N_35852,N_35608);
or U36129 (N_36129,N_34957,N_35214);
xor U36130 (N_36130,N_34082,N_35166);
nand U36131 (N_36131,N_34193,N_35938);
nand U36132 (N_36132,N_34134,N_34256);
and U36133 (N_36133,N_34349,N_35374);
nor U36134 (N_36134,N_35523,N_35648);
nor U36135 (N_36135,N_34059,N_34477);
nand U36136 (N_36136,N_35288,N_35115);
and U36137 (N_36137,N_34892,N_35164);
xnor U36138 (N_36138,N_35272,N_34571);
and U36139 (N_36139,N_34274,N_34035);
nor U36140 (N_36140,N_35192,N_35088);
nand U36141 (N_36141,N_34574,N_34111);
and U36142 (N_36142,N_35547,N_34241);
nor U36143 (N_36143,N_35750,N_35261);
or U36144 (N_36144,N_34062,N_34013);
nand U36145 (N_36145,N_35991,N_34914);
or U36146 (N_36146,N_34700,N_34301);
and U36147 (N_36147,N_35946,N_35493);
or U36148 (N_36148,N_34244,N_35068);
or U36149 (N_36149,N_35129,N_35935);
and U36150 (N_36150,N_35238,N_34958);
or U36151 (N_36151,N_35412,N_35415);
nor U36152 (N_36152,N_34646,N_34179);
nand U36153 (N_36153,N_35893,N_34180);
nor U36154 (N_36154,N_34409,N_35247);
or U36155 (N_36155,N_34095,N_34138);
nor U36156 (N_36156,N_35779,N_34625);
or U36157 (N_36157,N_35498,N_34043);
nand U36158 (N_36158,N_35421,N_35578);
and U36159 (N_36159,N_35024,N_35489);
nor U36160 (N_36160,N_35259,N_35987);
nor U36161 (N_36161,N_35201,N_34800);
or U36162 (N_36162,N_34590,N_35874);
nand U36163 (N_36163,N_34648,N_34262);
and U36164 (N_36164,N_34868,N_34890);
or U36165 (N_36165,N_35039,N_35468);
and U36166 (N_36166,N_34160,N_35121);
nor U36167 (N_36167,N_35894,N_35626);
xnor U36168 (N_36168,N_35361,N_35665);
nand U36169 (N_36169,N_35367,N_35880);
or U36170 (N_36170,N_35513,N_35728);
nor U36171 (N_36171,N_34313,N_35406);
or U36172 (N_36172,N_34398,N_35569);
xnor U36173 (N_36173,N_35086,N_35349);
and U36174 (N_36174,N_34157,N_35990);
and U36175 (N_36175,N_35849,N_35452);
xor U36176 (N_36176,N_35327,N_35019);
xor U36177 (N_36177,N_35153,N_35606);
nor U36178 (N_36178,N_34040,N_35966);
nand U36179 (N_36179,N_34873,N_34079);
nor U36180 (N_36180,N_34698,N_35543);
or U36181 (N_36181,N_34491,N_34130);
nor U36182 (N_36182,N_35747,N_35127);
xor U36183 (N_36183,N_34249,N_34652);
nand U36184 (N_36184,N_34290,N_35739);
nor U36185 (N_36185,N_35396,N_35399);
xor U36186 (N_36186,N_34781,N_34832);
or U36187 (N_36187,N_35185,N_35172);
nand U36188 (N_36188,N_34252,N_35321);
xnor U36189 (N_36189,N_35683,N_34229);
or U36190 (N_36190,N_35753,N_34493);
nor U36191 (N_36191,N_34270,N_35630);
and U36192 (N_36192,N_34382,N_34793);
or U36193 (N_36193,N_35478,N_35343);
and U36194 (N_36194,N_35706,N_35395);
nor U36195 (N_36195,N_35439,N_34480);
and U36196 (N_36196,N_35417,N_35246);
or U36197 (N_36197,N_34595,N_34253);
and U36198 (N_36198,N_34666,N_34204);
xnor U36199 (N_36199,N_34774,N_35216);
xnor U36200 (N_36200,N_35066,N_34552);
and U36201 (N_36201,N_34753,N_34826);
nor U36202 (N_36202,N_35993,N_34217);
nand U36203 (N_36203,N_34272,N_35487);
or U36204 (N_36204,N_34801,N_34225);
nand U36205 (N_36205,N_35832,N_34175);
and U36206 (N_36206,N_35660,N_35441);
nor U36207 (N_36207,N_35472,N_34504);
or U36208 (N_36208,N_35137,N_34185);
xnor U36209 (N_36209,N_34151,N_35741);
or U36210 (N_36210,N_34086,N_34880);
or U36211 (N_36211,N_35592,N_35637);
nand U36212 (N_36212,N_34210,N_34132);
nand U36213 (N_36213,N_34660,N_35503);
xnor U36214 (N_36214,N_34731,N_35152);
or U36215 (N_36215,N_35782,N_35432);
nand U36216 (N_36216,N_35521,N_34741);
xnor U36217 (N_36217,N_35018,N_35030);
nor U36218 (N_36218,N_35332,N_34092);
nand U36219 (N_36219,N_35037,N_34235);
nand U36220 (N_36220,N_34376,N_34533);
xor U36221 (N_36221,N_35700,N_34569);
or U36222 (N_36222,N_34943,N_34495);
and U36223 (N_36223,N_35405,N_35952);
nor U36224 (N_36224,N_34717,N_34281);
xor U36225 (N_36225,N_35562,N_34017);
xnor U36226 (N_36226,N_35806,N_34592);
nor U36227 (N_36227,N_34087,N_34923);
nor U36228 (N_36228,N_35366,N_35058);
or U36229 (N_36229,N_34777,N_34394);
and U36230 (N_36230,N_34341,N_35723);
nor U36231 (N_36231,N_34098,N_35359);
nor U36232 (N_36232,N_35839,N_34710);
nor U36233 (N_36233,N_34077,N_34366);
xnor U36234 (N_36234,N_34021,N_35695);
nand U36235 (N_36235,N_35925,N_35677);
nand U36236 (N_36236,N_35202,N_34678);
nand U36237 (N_36237,N_34788,N_35428);
nand U36238 (N_36238,N_34896,N_34447);
xnor U36239 (N_36239,N_35159,N_34517);
or U36240 (N_36240,N_35542,N_34915);
xor U36241 (N_36241,N_34864,N_34823);
xnor U36242 (N_36242,N_35784,N_35098);
nor U36243 (N_36243,N_34601,N_34853);
nand U36244 (N_36244,N_35554,N_35187);
and U36245 (N_36245,N_35838,N_35631);
or U36246 (N_36246,N_34221,N_34112);
or U36247 (N_36247,N_35102,N_34450);
nand U36248 (N_36248,N_34485,N_35927);
or U36249 (N_36249,N_34214,N_35467);
xor U36250 (N_36250,N_35407,N_35112);
xor U36251 (N_36251,N_35923,N_34547);
and U36252 (N_36252,N_35858,N_34459);
nor U36253 (N_36253,N_35701,N_35933);
xor U36254 (N_36254,N_35897,N_35814);
and U36255 (N_36255,N_34587,N_34258);
nand U36256 (N_36256,N_34831,N_35914);
nor U36257 (N_36257,N_35866,N_34454);
nor U36258 (N_36258,N_35996,N_35707);
nand U36259 (N_36259,N_34936,N_34430);
xor U36260 (N_36260,N_35530,N_34265);
and U36261 (N_36261,N_35287,N_35777);
nand U36262 (N_36262,N_35348,N_34119);
xor U36263 (N_36263,N_34818,N_35955);
or U36264 (N_36264,N_34291,N_34296);
xnor U36265 (N_36265,N_34778,N_34435);
and U36266 (N_36266,N_35699,N_34045);
or U36267 (N_36267,N_35819,N_35299);
xor U36268 (N_36268,N_35390,N_35869);
nor U36269 (N_36269,N_34093,N_35877);
nor U36270 (N_36270,N_34929,N_35566);
nand U36271 (N_36271,N_35083,N_34622);
nor U36272 (N_36272,N_34169,N_34154);
nor U36273 (N_36273,N_34050,N_35402);
or U36274 (N_36274,N_35444,N_35278);
or U36275 (N_36275,N_34344,N_34953);
and U36276 (N_36276,N_34707,N_34187);
nand U36277 (N_36277,N_34267,N_34878);
xor U36278 (N_36278,N_34061,N_35393);
or U36279 (N_36279,N_35292,N_34273);
and U36280 (N_36280,N_34670,N_35811);
or U36281 (N_36281,N_35563,N_34846);
and U36282 (N_36282,N_35628,N_34989);
xor U36283 (N_36283,N_35251,N_35907);
or U36284 (N_36284,N_35149,N_34694);
nor U36285 (N_36285,N_35241,N_35268);
or U36286 (N_36286,N_34791,N_35020);
nor U36287 (N_36287,N_34213,N_34080);
nand U36288 (N_36288,N_35460,N_35901);
nand U36289 (N_36289,N_35190,N_34400);
or U36290 (N_36290,N_35160,N_35675);
and U36291 (N_36291,N_35672,N_34839);
nor U36292 (N_36292,N_34729,N_34016);
nand U36293 (N_36293,N_35479,N_35799);
nand U36294 (N_36294,N_35855,N_35930);
nor U36295 (N_36295,N_34109,N_34089);
nor U36296 (N_36296,N_35884,N_35038);
and U36297 (N_36297,N_34287,N_34598);
or U36298 (N_36298,N_35802,N_35928);
nor U36299 (N_36299,N_35831,N_35208);
nand U36300 (N_36300,N_35520,N_35486);
and U36301 (N_36301,N_34310,N_34074);
and U36302 (N_36302,N_34792,N_35398);
xor U36303 (N_36303,N_34560,N_34063);
xor U36304 (N_36304,N_34538,N_34553);
and U36305 (N_36305,N_35977,N_35437);
or U36306 (N_36306,N_34408,N_35290);
nand U36307 (N_36307,N_35015,N_34207);
nand U36308 (N_36308,N_34630,N_34638);
nand U36309 (N_36309,N_35207,N_35309);
nand U36310 (N_36310,N_35044,N_35411);
nor U36311 (N_36311,N_35941,N_34676);
nand U36312 (N_36312,N_35703,N_34260);
xnor U36313 (N_36313,N_35009,N_35607);
xnor U36314 (N_36314,N_34934,N_34125);
or U36315 (N_36315,N_34156,N_34393);
xor U36316 (N_36316,N_35370,N_34875);
or U36317 (N_36317,N_35466,N_35639);
and U36318 (N_36318,N_35006,N_35087);
and U36319 (N_36319,N_34007,N_34499);
and U36320 (N_36320,N_34505,N_35945);
and U36321 (N_36321,N_34987,N_34775);
nand U36322 (N_36322,N_35775,N_35834);
xor U36323 (N_36323,N_34472,N_34257);
and U36324 (N_36324,N_35296,N_34926);
or U36325 (N_36325,N_34359,N_35453);
xor U36326 (N_36326,N_35565,N_34948);
xnor U36327 (N_36327,N_34996,N_35222);
or U36328 (N_36328,N_34860,N_35264);
or U36329 (N_36329,N_35409,N_34525);
nor U36330 (N_36330,N_34334,N_34367);
or U36331 (N_36331,N_35686,N_34143);
xnor U36332 (N_36332,N_35193,N_35659);
and U36333 (N_36333,N_34070,N_35386);
xnor U36334 (N_36334,N_35265,N_35213);
or U36335 (N_36335,N_34452,N_34127);
or U36336 (N_36336,N_35780,N_34656);
xor U36337 (N_36337,N_35603,N_35173);
xor U36338 (N_36338,N_35715,N_34088);
and U36339 (N_36339,N_35325,N_34462);
and U36340 (N_36340,N_35564,N_34404);
or U36341 (N_36341,N_34279,N_35026);
nand U36342 (N_36342,N_34186,N_34679);
and U36343 (N_36343,N_35188,N_35770);
and U36344 (N_36344,N_35859,N_35647);
xor U36345 (N_36345,N_35676,N_34835);
nand U36346 (N_36346,N_34924,N_34910);
or U36347 (N_36347,N_35536,N_34030);
or U36348 (N_36348,N_35499,N_34639);
and U36349 (N_36349,N_34969,N_35740);
xor U36350 (N_36350,N_35615,N_35998);
and U36351 (N_36351,N_35167,N_35786);
and U36352 (N_36352,N_34280,N_34346);
or U36353 (N_36353,N_34838,N_34236);
and U36354 (N_36354,N_35021,N_35336);
or U36355 (N_36355,N_35506,N_35368);
or U36356 (N_36356,N_34034,N_34512);
or U36357 (N_36357,N_34500,N_34162);
nand U36358 (N_36358,N_34812,N_35429);
nand U36359 (N_36359,N_34701,N_35377);
or U36360 (N_36360,N_35762,N_34100);
nand U36361 (N_36361,N_34022,N_35992);
xnor U36362 (N_36362,N_35760,N_34667);
and U36363 (N_36363,N_34937,N_34243);
nand U36364 (N_36364,N_35451,N_35641);
nor U36365 (N_36365,N_35571,N_34904);
or U36366 (N_36366,N_35601,N_35492);
xnor U36367 (N_36367,N_34849,N_35082);
nand U36368 (N_36368,N_35575,N_35633);
nor U36369 (N_36369,N_35400,N_35339);
or U36370 (N_36370,N_34668,N_35518);
nand U36371 (N_36371,N_35580,N_35146);
and U36372 (N_36372,N_35226,N_35481);
and U36373 (N_36373,N_34899,N_34837);
nor U36374 (N_36374,N_35174,N_34348);
nor U36375 (N_36375,N_34998,N_35932);
nand U36376 (N_36376,N_34411,N_35515);
and U36377 (N_36377,N_34369,N_35560);
nor U36378 (N_36378,N_35596,N_35338);
nor U36379 (N_36379,N_34921,N_34909);
or U36380 (N_36380,N_35862,N_35150);
xor U36381 (N_36381,N_35017,N_35625);
nand U36382 (N_36382,N_34075,N_35284);
and U36383 (N_36383,N_34126,N_35600);
and U36384 (N_36384,N_35781,N_34113);
and U36385 (N_36385,N_34399,N_35355);
nand U36386 (N_36386,N_35067,N_34510);
xnor U36387 (N_36387,N_34858,N_34714);
and U36388 (N_36388,N_35344,N_34681);
or U36389 (N_36389,N_34578,N_34877);
and U36390 (N_36390,N_34467,N_34199);
or U36391 (N_36391,N_35196,N_34732);
or U36392 (N_36392,N_35573,N_34836);
nor U36393 (N_36393,N_34573,N_34597);
xnor U36394 (N_36394,N_34857,N_35335);
nand U36395 (N_36395,N_34308,N_35358);
nor U36396 (N_36396,N_34006,N_34054);
and U36397 (N_36397,N_35820,N_34451);
or U36398 (N_36398,N_35795,N_34589);
nand U36399 (N_36399,N_35025,N_35275);
nand U36400 (N_36400,N_34032,N_34944);
nand U36401 (N_36401,N_35065,N_35837);
or U36402 (N_36402,N_35281,N_35450);
nor U36403 (N_36403,N_34616,N_34901);
and U36404 (N_36404,N_34329,N_34482);
and U36405 (N_36405,N_34364,N_35854);
nor U36406 (N_36406,N_35942,N_34817);
or U36407 (N_36407,N_35685,N_35589);
nand U36408 (N_36408,N_34725,N_34527);
nor U36409 (N_36409,N_35956,N_35951);
and U36410 (N_36410,N_35720,N_35132);
nor U36411 (N_36411,N_34284,N_34995);
xor U36412 (N_36412,N_35271,N_34228);
and U36413 (N_36413,N_35045,N_35796);
and U36414 (N_36414,N_34669,N_35342);
xor U36415 (N_36415,N_34671,N_35734);
and U36416 (N_36416,N_35937,N_35939);
and U36417 (N_36417,N_35729,N_34798);
nand U36418 (N_36418,N_35845,N_35234);
or U36419 (N_36419,N_35888,N_34894);
or U36420 (N_36420,N_34378,N_35277);
and U36421 (N_36421,N_35726,N_35372);
nor U36422 (N_36422,N_35610,N_34307);
or U36423 (N_36423,N_34719,N_35443);
nor U36424 (N_36424,N_34663,N_35763);
nand U36425 (N_36425,N_34437,N_35430);
nor U36426 (N_36426,N_34076,N_35885);
xnor U36427 (N_36427,N_34216,N_34397);
nor U36428 (N_36428,N_34593,N_35778);
xor U36429 (N_36429,N_34806,N_35871);
and U36430 (N_36430,N_35154,N_34759);
or U36431 (N_36431,N_35797,N_34405);
nand U36432 (N_36432,N_35435,N_35965);
nor U36433 (N_36433,N_35084,N_35661);
nand U36434 (N_36434,N_34602,N_34687);
nor U36435 (N_36435,N_35440,N_35408);
xnor U36436 (N_36436,N_35921,N_35232);
nand U36437 (N_36437,N_35738,N_34540);
and U36438 (N_36438,N_34246,N_35882);
xor U36439 (N_36439,N_35074,N_35331);
nor U36440 (N_36440,N_35718,N_35483);
xnor U36441 (N_36441,N_35091,N_34012);
nor U36442 (N_36442,N_34402,N_35594);
or U36443 (N_36443,N_35936,N_34403);
xnor U36444 (N_36444,N_34427,N_35667);
nor U36445 (N_36445,N_35484,N_34492);
or U36446 (N_36446,N_34146,N_35544);
xnor U36447 (N_36447,N_34102,N_34647);
and U36448 (N_36448,N_34370,N_35742);
xor U36449 (N_36449,N_35920,N_34766);
and U36450 (N_36450,N_35096,N_34561);
xnor U36451 (N_36451,N_34920,N_35279);
xnor U36452 (N_36452,N_34511,N_34565);
or U36453 (N_36453,N_34181,N_35997);
and U36454 (N_36454,N_34870,N_35161);
or U36455 (N_36455,N_35964,N_35260);
or U36456 (N_36456,N_34406,N_35051);
and U36457 (N_36457,N_34827,N_35267);
nor U36458 (N_36458,N_35126,N_35457);
and U36459 (N_36459,N_34607,N_35969);
and U36460 (N_36460,N_35761,N_34245);
nor U36461 (N_36461,N_34636,N_35510);
nand U36462 (N_36462,N_34804,N_35994);
xor U36463 (N_36463,N_35929,N_35559);
nand U36464 (N_36464,N_34654,N_35239);
nor U36465 (N_36465,N_34295,N_35256);
nand U36466 (N_36466,N_35949,N_35803);
xnor U36467 (N_36467,N_35857,N_34709);
nand U36468 (N_36468,N_34381,N_34758);
or U36469 (N_36469,N_34850,N_34821);
nand U36470 (N_36470,N_34693,N_35462);
nand U36471 (N_36471,N_35341,N_34726);
and U36472 (N_36472,N_34486,N_34705);
and U36473 (N_36473,N_35242,N_35847);
or U36474 (N_36474,N_34841,N_35204);
and U36475 (N_36475,N_34230,N_35687);
and U36476 (N_36476,N_35092,N_35328);
xnor U36477 (N_36477,N_35141,N_34918);
xnor U36478 (N_36478,N_34724,N_34263);
and U36479 (N_36479,N_34315,N_35539);
or U36480 (N_36480,N_35283,N_35961);
or U36481 (N_36481,N_34497,N_35389);
and U36482 (N_36482,N_34496,N_34463);
or U36483 (N_36483,N_34746,N_34611);
nand U36484 (N_36484,N_35900,N_34254);
and U36485 (N_36485,N_34713,N_34190);
or U36486 (N_36486,N_35262,N_35627);
xor U36487 (N_36487,N_34964,N_34541);
nor U36488 (N_36488,N_34783,N_35558);
and U36489 (N_36489,N_34129,N_34137);
and U36490 (N_36490,N_34702,N_34968);
or U36491 (N_36491,N_34448,N_34372);
or U36492 (N_36492,N_35000,N_35365);
nor U36493 (N_36493,N_34828,N_34723);
nor U36494 (N_36494,N_35094,N_34209);
nor U36495 (N_36495,N_34606,N_34977);
xor U36496 (N_36496,N_34884,N_35680);
nand U36497 (N_36497,N_35353,N_34927);
and U36498 (N_36498,N_34720,N_34722);
nor U36499 (N_36499,N_34288,N_34961);
and U36500 (N_36500,N_35089,N_34524);
and U36501 (N_36501,N_35519,N_35970);
xor U36502 (N_36502,N_34192,N_35744);
nor U36503 (N_36503,N_34321,N_34848);
or U36504 (N_36504,N_34277,N_35798);
nand U36505 (N_36505,N_35774,N_34874);
and U36506 (N_36506,N_35054,N_34487);
or U36507 (N_36507,N_35532,N_35546);
nor U36508 (N_36508,N_35392,N_34908);
or U36509 (N_36509,N_35438,N_35868);
nand U36510 (N_36510,N_35816,N_34577);
and U36511 (N_36511,N_35295,N_35751);
nand U36512 (N_36512,N_35712,N_34854);
nor U36513 (N_36513,N_35324,N_35602);
and U36514 (N_36514,N_35081,N_34941);
or U36515 (N_36515,N_35385,N_35691);
nand U36516 (N_36516,N_35012,N_35525);
xor U36517 (N_36517,N_34361,N_34649);
xnor U36518 (N_36518,N_34003,N_35549);
xnor U36519 (N_36519,N_35394,N_35801);
and U36520 (N_36520,N_35257,N_35759);
xnor U36521 (N_36521,N_34938,N_34037);
nand U36522 (N_36522,N_34488,N_34978);
and U36523 (N_36523,N_35892,N_35205);
or U36524 (N_36524,N_34428,N_34224);
and U36525 (N_36525,N_34682,N_34833);
nand U36526 (N_36526,N_34336,N_35864);
or U36527 (N_36527,N_35133,N_35985);
xnor U36528 (N_36528,N_34000,N_34771);
xor U36529 (N_36529,N_35652,N_34208);
nor U36530 (N_36530,N_34617,N_35049);
and U36531 (N_36531,N_34803,N_35419);
nand U36532 (N_36532,N_35329,N_35134);
and U36533 (N_36533,N_34564,N_35077);
nor U36534 (N_36534,N_35047,N_34686);
or U36535 (N_36535,N_35863,N_34387);
nand U36536 (N_36536,N_34289,N_35711);
nand U36537 (N_36537,N_35733,N_34328);
and U36538 (N_36538,N_35962,N_35553);
or U36539 (N_36539,N_34222,N_34956);
and U36540 (N_36540,N_34673,N_34993);
nand U36541 (N_36541,N_34696,N_34690);
xnor U36542 (N_36542,N_35318,N_35424);
xor U36543 (N_36543,N_34455,N_35629);
xnor U36544 (N_36544,N_35912,N_35757);
xnor U36545 (N_36545,N_35909,N_35572);
nand U36546 (N_36546,N_34358,N_34889);
or U36547 (N_36547,N_34782,N_34750);
and U36548 (N_36548,N_34907,N_34830);
and U36549 (N_36549,N_35371,N_34665);
nand U36550 (N_36550,N_35957,N_35870);
nand U36551 (N_36551,N_35768,N_34861);
and U36552 (N_36552,N_35567,N_34110);
nand U36553 (N_36553,N_35902,N_35570);
nor U36554 (N_36554,N_35106,N_35865);
nand U36555 (N_36555,N_34640,N_35609);
nand U36556 (N_36556,N_35209,N_34223);
and U36557 (N_36557,N_34628,N_34519);
and U36558 (N_36558,N_35016,N_34071);
nor U36559 (N_36559,N_35248,N_34865);
nand U36560 (N_36560,N_34935,N_35669);
nor U36561 (N_36561,N_35240,N_35114);
xnor U36562 (N_36562,N_35605,N_35593);
nor U36563 (N_36563,N_34990,N_35227);
and U36564 (N_36564,N_35846,N_35731);
and U36565 (N_36565,N_34015,N_34594);
or U36566 (N_36566,N_34294,N_35079);
xnor U36567 (N_36567,N_35710,N_34925);
nand U36568 (N_36568,N_34840,N_34761);
xnor U36569 (N_36569,N_35427,N_34773);
and U36570 (N_36570,N_34377,N_35476);
nor U36571 (N_36571,N_34251,N_35063);
nor U36572 (N_36572,N_35008,N_34871);
or U36573 (N_36573,N_34449,N_34651);
nor U36574 (N_36574,N_35075,N_34641);
nor U36575 (N_36575,N_35823,N_35458);
nor U36576 (N_36576,N_34103,N_35042);
or U36577 (N_36577,N_35449,N_35029);
xor U36578 (N_36578,N_35313,N_35908);
nor U36579 (N_36579,N_34684,N_35228);
nor U36580 (N_36580,N_34862,N_34549);
nor U36581 (N_36581,N_34886,N_34674);
or U36582 (N_36582,N_35095,N_34333);
nor U36583 (N_36583,N_34992,N_35496);
or U36584 (N_36584,N_35979,N_34822);
nor U36585 (N_36585,N_34536,N_34275);
nand U36586 (N_36586,N_35135,N_34083);
xor U36587 (N_36587,N_34756,N_34683);
nor U36588 (N_36588,N_35140,N_34419);
and U36589 (N_36589,N_34118,N_35585);
xnor U36590 (N_36590,N_35850,N_34422);
xor U36591 (N_36591,N_35524,N_35401);
and U36592 (N_36592,N_35250,N_34101);
xor U36593 (N_36593,N_34619,N_35800);
nand U36594 (N_36594,N_35656,N_34814);
nand U36595 (N_36595,N_34919,N_34718);
or U36596 (N_36596,N_35391,N_35064);
xnor U36597 (N_36597,N_35494,N_34581);
nor U36598 (N_36598,N_34401,N_34810);
or U36599 (N_36599,N_34170,N_35883);
and U36600 (N_36600,N_35245,N_35255);
xnor U36601 (N_36601,N_34966,N_35526);
nand U36602 (N_36602,N_35122,N_34114);
and U36603 (N_36603,N_34588,N_34677);
nor U36604 (N_36604,N_35243,N_35827);
or U36605 (N_36605,N_34064,N_34424);
or U36606 (N_36606,N_34052,N_34464);
or U36607 (N_36607,N_35828,N_35221);
nor U36608 (N_36608,N_34196,N_34418);
nor U36609 (N_36609,N_35919,N_35619);
nand U36610 (N_36610,N_35356,N_34239);
or U36611 (N_36611,N_34780,N_34445);
or U36612 (N_36612,N_34820,N_34465);
nor U36613 (N_36613,N_34551,N_35454);
nor U36614 (N_36614,N_34697,N_34991);
and U36615 (N_36615,N_34906,N_34727);
nor U36616 (N_36616,N_34903,N_35501);
nand U36617 (N_36617,N_34203,N_35931);
or U36618 (N_36618,N_35552,N_35794);
and U36619 (N_36619,N_34618,N_35754);
and U36620 (N_36620,N_34131,N_35078);
or U36621 (N_36621,N_35317,N_34881);
or U36622 (N_36622,N_34902,N_34443);
nor U36623 (N_36623,N_35423,N_35237);
nand U36624 (N_36624,N_34340,N_34395);
and U36625 (N_36625,N_34431,N_35851);
xnor U36626 (N_36626,N_34945,N_35387);
nand U36627 (N_36627,N_35791,N_34863);
nor U36628 (N_36628,N_34058,N_34528);
xor U36629 (N_36629,N_35100,N_34976);
xnor U36630 (N_36630,N_35655,N_34916);
nor U36631 (N_36631,N_34982,N_35808);
and U36632 (N_36632,N_35076,N_35972);
nor U36633 (N_36633,N_35716,N_35477);
nor U36634 (N_36634,N_35730,N_34247);
or U36635 (N_36635,N_34931,N_35732);
xor U36636 (N_36636,N_35061,N_34633);
nand U36637 (N_36637,N_35131,N_35597);
nand U36638 (N_36638,N_35199,N_35737);
nand U36639 (N_36639,N_34932,N_35767);
or U36640 (N_36640,N_35507,N_35670);
nor U36641 (N_36641,N_34829,N_34733);
nand U36642 (N_36642,N_34184,N_35792);
and U36643 (N_36643,N_35381,N_35168);
nand U36644 (N_36644,N_35471,N_34355);
or U36645 (N_36645,N_34612,N_34433);
xor U36646 (N_36646,N_35404,N_34286);
nor U36647 (N_36647,N_34807,N_34010);
or U36648 (N_36648,N_35363,N_34091);
nand U36649 (N_36649,N_34893,N_35971);
or U36650 (N_36650,N_35813,N_34115);
or U36651 (N_36651,N_34529,N_35480);
nor U36652 (N_36652,N_35456,N_34338);
xor U36653 (N_36653,N_35662,N_35818);
nand U36654 (N_36654,N_35534,N_35954);
and U36655 (N_36655,N_35983,N_35113);
nor U36656 (N_36656,N_34476,N_34354);
or U36657 (N_36657,N_35890,N_35527);
xnor U36658 (N_36658,N_35736,N_34432);
xor U36659 (N_36659,N_35981,N_34178);
xor U36660 (N_36660,N_34930,N_35642);
nor U36661 (N_36661,N_34786,N_34852);
and U36662 (N_36662,N_34580,N_35583);
xnor U36663 (N_36663,N_34624,N_34353);
and U36664 (N_36664,N_34742,N_34434);
nor U36665 (N_36665,N_35984,N_35551);
xnor U36666 (N_36666,N_35145,N_35210);
or U36667 (N_36667,N_35459,N_35383);
xnor U36668 (N_36668,N_34044,N_35036);
and U36669 (N_36669,N_35005,N_34046);
xor U36670 (N_36670,N_35183,N_34141);
or U36671 (N_36671,N_34202,N_35354);
xnor U36672 (N_36672,N_34951,N_34414);
nand U36673 (N_36673,N_34197,N_34563);
or U36674 (N_36674,N_35926,N_35517);
and U36675 (N_36675,N_34599,N_35123);
and U36676 (N_36676,N_34653,N_35182);
xor U36677 (N_36677,N_35203,N_34368);
xor U36678 (N_36678,N_34952,N_35958);
or U36679 (N_36679,N_34335,N_34164);
nor U36680 (N_36680,N_34999,N_35645);
and U36681 (N_36681,N_35944,N_34026);
nand U36682 (N_36682,N_35048,N_34147);
and U36683 (N_36683,N_34106,N_35650);
and U36684 (N_36684,N_34768,N_34960);
nand U36685 (N_36685,N_35014,N_34323);
xnor U36686 (N_36686,N_35822,N_35490);
nand U36687 (N_36687,N_34417,N_35643);
and U36688 (N_36688,N_35171,N_35143);
nand U36689 (N_36689,N_35013,N_35285);
and U36690 (N_36690,N_35689,N_34234);
nor U36691 (N_36691,N_34897,N_34764);
or U36692 (N_36692,N_34582,N_34205);
nand U36693 (N_36693,N_35198,N_35244);
nand U36694 (N_36694,N_35812,N_34107);
nor U36695 (N_36695,N_35050,N_34219);
nand U36696 (N_36696,N_35577,N_34002);
nor U36697 (N_36697,N_35046,N_34986);
nand U36698 (N_36698,N_35614,N_34471);
or U36699 (N_36699,N_34195,N_35561);
nor U36700 (N_36700,N_35529,N_35579);
or U36701 (N_36701,N_35705,N_34655);
nor U36702 (N_36702,N_35568,N_35225);
or U36703 (N_36703,N_35758,N_34150);
nand U36704 (N_36704,N_34028,N_35612);
xnor U36705 (N_36705,N_35413,N_34104);
nor U36706 (N_36706,N_35194,N_34757);
nor U36707 (N_36707,N_35840,N_35445);
or U36708 (N_36708,N_34955,N_34474);
or U36709 (N_36709,N_34912,N_34396);
nand U36710 (N_36710,N_34326,N_35574);
or U36711 (N_36711,N_34311,N_34365);
or U36712 (N_36712,N_34038,N_35886);
nand U36713 (N_36713,N_34166,N_34165);
nor U36714 (N_36714,N_34380,N_34554);
nand U36715 (N_36715,N_35905,N_35548);
nor U36716 (N_36716,N_34834,N_34971);
and U36717 (N_36717,N_34664,N_34056);
nor U36718 (N_36718,N_35181,N_34615);
and U36719 (N_36719,N_34004,N_34567);
nor U36720 (N_36720,N_35378,N_35397);
xnor U36721 (N_36721,N_35212,N_35136);
or U36722 (N_36722,N_35915,N_34031);
nor U36723 (N_36723,N_35766,N_34073);
xnor U36724 (N_36724,N_34988,N_34744);
and U36725 (N_36725,N_35347,N_35120);
nor U36726 (N_36726,N_35352,N_35713);
and U36727 (N_36727,N_34621,N_35144);
nor U36728 (N_36728,N_34743,N_35470);
and U36729 (N_36729,N_35682,N_35664);
nand U36730 (N_36730,N_34226,N_35913);
nand U36731 (N_36731,N_34384,N_35771);
nand U36732 (N_36732,N_34568,N_34772);
nor U36733 (N_36733,N_35853,N_34515);
and U36734 (N_36734,N_35898,N_35895);
nor U36735 (N_36735,N_34453,N_34297);
nand U36736 (N_36736,N_34330,N_34271);
nor U36737 (N_36737,N_35887,N_35624);
xor U36738 (N_36738,N_34739,N_34144);
or U36739 (N_36739,N_34632,N_35693);
or U36740 (N_36740,N_35790,N_34173);
nand U36741 (N_36741,N_34661,N_35495);
nor U36742 (N_36742,N_35809,N_34760);
nor U36743 (N_36743,N_34603,N_34255);
nand U36744 (N_36744,N_34959,N_34148);
xor U36745 (N_36745,N_34172,N_34331);
nor U36746 (N_36746,N_35940,N_35632);
and U36747 (N_36747,N_34876,N_35588);
nand U36748 (N_36748,N_35861,N_34047);
nor U36749 (N_36749,N_34057,N_35986);
nand U36750 (N_36750,N_35474,N_34096);
or U36751 (N_36751,N_35130,N_35273);
nand U36752 (N_36752,N_34819,N_35848);
nand U36753 (N_36753,N_35211,N_34591);
and U36754 (N_36754,N_34490,N_34794);
or U36755 (N_36755,N_35286,N_35475);
nand U36756 (N_36756,N_35856,N_34218);
nor U36757 (N_36757,N_35508,N_35764);
or U36758 (N_36758,N_34322,N_34458);
xnor U36759 (N_36759,N_34412,N_34332);
xor U36760 (N_36760,N_34120,N_34155);
or U36761 (N_36761,N_34721,N_34845);
xor U36762 (N_36762,N_34735,N_35055);
nor U36763 (N_36763,N_34446,N_35829);
nor U36764 (N_36764,N_35316,N_34438);
xnor U36765 (N_36765,N_34796,N_34642);
or U36766 (N_36766,N_35973,N_34094);
or U36767 (N_36767,N_35357,N_35350);
nor U36768 (N_36768,N_35714,N_34122);
nand U36769 (N_36769,N_34883,N_34555);
nand U36770 (N_36770,N_34468,N_34436);
nand U36771 (N_36771,N_35464,N_34051);
nand U36772 (N_36772,N_34211,N_35057);
nand U36773 (N_36773,N_34802,N_34014);
nor U36774 (N_36774,N_35722,N_35220);
xnor U36775 (N_36775,N_35550,N_34784);
nor U36776 (N_36776,N_34293,N_34543);
nand U36777 (N_36777,N_35721,N_35960);
nand U36778 (N_36778,N_35953,N_34233);
xnor U36779 (N_36779,N_34708,N_34117);
and U36780 (N_36780,N_34171,N_35557);
and U36781 (N_36781,N_34627,N_34776);
nand U36782 (N_36782,N_35436,N_35333);
xnor U36783 (N_36783,N_34167,N_34584);
or U36784 (N_36784,N_35528,N_34460);
and U36785 (N_36785,N_34730,N_34813);
or U36786 (N_36786,N_34020,N_35388);
xor U36787 (N_36787,N_35465,N_35833);
and U36788 (N_36788,N_35011,N_35282);
nand U36789 (N_36789,N_35043,N_35177);
and U36790 (N_36790,N_34650,N_34596);
and U36791 (N_36791,N_35671,N_35041);
nor U36792 (N_36792,N_35826,N_35206);
nand U36793 (N_36793,N_35899,N_34623);
or U36794 (N_36794,N_35473,N_35375);
or U36795 (N_36795,N_34613,N_34183);
or U36796 (N_36796,N_34530,N_35040);
xor U36797 (N_36797,N_34426,N_34188);
nand U36798 (N_36798,N_35666,N_35293);
nor U36799 (N_36799,N_35073,N_35653);
and U36800 (N_36800,N_34198,N_34362);
or U36801 (N_36801,N_35169,N_34558);
or U36802 (N_36802,N_35157,N_35319);
nor U36803 (N_36803,N_34521,N_35410);
and U36804 (N_36804,N_34513,N_34544);
and U36805 (N_36805,N_35704,N_35749);
or U36806 (N_36806,N_34905,N_34189);
xnor U36807 (N_36807,N_35916,N_35727);
or U36808 (N_36808,N_35217,N_34339);
or U36809 (N_36809,N_35218,N_35461);
nand U36810 (N_36810,N_34699,N_35463);
xor U36811 (N_36811,N_34153,N_34949);
nor U36812 (N_36812,N_35308,N_35448);
and U36813 (N_36813,N_35101,N_35910);
and U36814 (N_36814,N_35069,N_34375);
or U36815 (N_36815,N_34029,N_35224);
nand U36816 (N_36816,N_34374,N_34097);
xnor U36817 (N_36817,N_34292,N_35769);
or U36818 (N_36818,N_34041,N_35431);
nand U36819 (N_36819,N_35158,N_34498);
nand U36820 (N_36820,N_35337,N_34575);
or U36821 (N_36821,N_35697,N_34762);
and U36822 (N_36822,N_34005,N_34583);
or U36823 (N_36823,N_34501,N_34215);
and U36824 (N_36824,N_34728,N_34168);
and U36825 (N_36825,N_35881,N_34851);
or U36826 (N_36826,N_34489,N_35613);
xor U36827 (N_36827,N_35422,N_34191);
or U36828 (N_36828,N_35576,N_34379);
nand U36829 (N_36829,N_35189,N_34269);
nor U36830 (N_36830,N_35772,N_35620);
nand U36831 (N_36831,N_35842,N_35755);
nor U36832 (N_36832,N_35815,N_35841);
nor U36833 (N_36833,N_35447,N_35491);
and U36834 (N_36834,N_34008,N_34299);
nor U36835 (N_36835,N_34605,N_34159);
and U36836 (N_36836,N_34542,N_35215);
xnor U36837 (N_36837,N_34009,N_34312);
xnor U36838 (N_36838,N_34133,N_35644);
and U36839 (N_36839,N_34752,N_34751);
nand U36840 (N_36840,N_35280,N_34319);
and U36841 (N_36841,N_34506,N_34692);
xnor U36842 (N_36842,N_35010,N_34787);
xnor U36843 (N_36843,N_35978,N_35873);
or U36844 (N_36844,N_34090,N_35434);
nor U36845 (N_36845,N_35004,N_34481);
nand U36846 (N_36846,N_34736,N_34503);
xor U36847 (N_36847,N_34675,N_34444);
nand U36848 (N_36848,N_35258,N_35156);
xor U36849 (N_36849,N_34695,N_34635);
nor U36850 (N_36850,N_35151,N_34680);
xnor U36851 (N_36851,N_34643,N_34027);
xor U36852 (N_36852,N_34033,N_34343);
nand U36853 (N_36853,N_35230,N_35345);
nand U36854 (N_36854,N_35270,N_34440);
or U36855 (N_36855,N_34421,N_34765);
xor U36856 (N_36856,N_35959,N_34962);
xor U36857 (N_36857,N_34324,N_34194);
xnor U36858 (N_36858,N_35678,N_35830);
nor U36859 (N_36859,N_35512,N_34206);
and U36860 (N_36860,N_35305,N_34420);
and U36861 (N_36861,N_35323,N_35967);
nor U36862 (N_36862,N_34855,N_34036);
xor U36863 (N_36863,N_34532,N_34371);
nand U36864 (N_36864,N_34859,N_35376);
or U36865 (N_36865,N_35176,N_35776);
nand U36866 (N_36866,N_34898,N_35306);
or U36867 (N_36867,N_34711,N_34779);
and U36868 (N_36868,N_35663,N_34227);
and U36869 (N_36869,N_34539,N_35426);
or U36870 (N_36870,N_34805,N_34620);
nand U36871 (N_36871,N_35698,N_35649);
xor U36872 (N_36872,N_34785,N_35033);
nor U36873 (N_36873,N_35836,N_35060);
or U36874 (N_36874,N_34537,N_34325);
and U36875 (N_36875,N_34808,N_34128);
nand U36876 (N_36876,N_35023,N_35889);
nor U36877 (N_36877,N_35903,N_35170);
nor U36878 (N_36878,N_35178,N_35307);
and U36879 (N_36879,N_34145,N_34048);
or U36880 (N_36880,N_35195,N_34689);
nor U36881 (N_36881,N_34391,N_35581);
or U36882 (N_36882,N_35692,N_35180);
and U36883 (N_36883,N_35694,N_35249);
nand U36884 (N_36884,N_34345,N_35090);
or U36885 (N_36885,N_35382,N_34039);
and U36886 (N_36886,N_35105,N_35658);
xor U36887 (N_36887,N_35488,N_34200);
nand U36888 (N_36888,N_34586,N_35485);
nand U36889 (N_36889,N_35696,N_35263);
or U36890 (N_36890,N_35773,N_35072);
nor U36891 (N_36891,N_35062,N_35752);
and U36892 (N_36892,N_34442,N_35310);
nor U36893 (N_36893,N_34337,N_35403);
and U36894 (N_36894,N_34947,N_35584);
nor U36895 (N_36895,N_34268,N_35311);
and U36896 (N_36896,N_35922,N_34081);
nor U36897 (N_36897,N_34351,N_34282);
and U36898 (N_36898,N_35497,N_35425);
nand U36899 (N_36899,N_34136,N_34410);
nand U36900 (N_36900,N_35807,N_35690);
or U36901 (N_36901,N_34060,N_34799);
nor U36902 (N_36902,N_34867,N_34520);
nor U36903 (N_36903,N_34001,N_35294);
nand U36904 (N_36904,N_35963,N_34303);
xor U36905 (N_36905,N_34514,N_35516);
and U36906 (N_36906,N_34659,N_35235);
nor U36907 (N_36907,N_34300,N_34585);
nor U36908 (N_36908,N_34946,N_35053);
xor U36909 (N_36909,N_34712,N_34614);
xor U36910 (N_36910,N_34248,N_35103);
xnor U36911 (N_36911,N_34055,N_35604);
xor U36912 (N_36912,N_34139,N_34522);
or U36913 (N_36913,N_34970,N_34704);
and U36914 (N_36914,N_35509,N_34306);
nand U36915 (N_36915,N_34163,N_35537);
nand U36916 (N_36916,N_34763,N_34298);
and U36917 (N_36917,N_34548,N_35442);
and U36918 (N_36918,N_34386,N_35635);
nand U36919 (N_36919,N_34121,N_35027);
or U36920 (N_36920,N_35843,N_35586);
or U36921 (N_36921,N_35482,N_35746);
xnor U36922 (N_36922,N_35330,N_34342);
and U36923 (N_36923,N_34795,N_34738);
or U36924 (N_36924,N_34347,N_35745);
nor U36925 (N_36925,N_34770,N_35351);
or U36926 (N_36926,N_34645,N_34385);
or U36927 (N_36927,N_34535,N_34212);
nand U36928 (N_36928,N_35298,N_35111);
nand U36929 (N_36929,N_35165,N_35725);
xor U36930 (N_36930,N_34494,N_34922);
and U36931 (N_36931,N_34631,N_35147);
nand U36932 (N_36932,N_34019,N_35455);
xor U36933 (N_36933,N_34734,N_34872);
xnor U36934 (N_36934,N_34963,N_34278);
nor U36935 (N_36935,N_35128,N_35522);
nand U36936 (N_36936,N_35002,N_34754);
nand U36937 (N_36937,N_34176,N_35420);
or U36938 (N_36938,N_35555,N_34888);
and U36939 (N_36939,N_34657,N_35587);
and U36940 (N_36940,N_35116,N_35878);
xor U36941 (N_36941,N_34309,N_35223);
nand U36942 (N_36942,N_35904,N_35709);
xor U36943 (N_36943,N_34917,N_34790);
nand U36944 (N_36944,N_34237,N_34425);
or U36945 (N_36945,N_35821,N_35879);
xnor U36946 (N_36946,N_35301,N_34797);
or U36947 (N_36947,N_35805,N_35097);
and U36948 (N_36948,N_35844,N_35124);
xnor U36949 (N_36949,N_34407,N_35340);
nor U36950 (N_36950,N_35059,N_34933);
nor U36951 (N_36951,N_35322,N_34608);
xnor U36952 (N_36952,N_34161,N_34637);
or U36953 (N_36953,N_35540,N_34844);
and U36954 (N_36954,N_34320,N_34457);
and U36955 (N_36955,N_35867,N_35765);
or U36956 (N_36956,N_34285,N_35312);
nor U36957 (N_36957,N_35142,N_35304);
nand U36958 (N_36958,N_34685,N_35876);
xnor U36959 (N_36959,N_35681,N_34913);
nor U36960 (N_36960,N_34158,N_34429);
and U36961 (N_36961,N_34626,N_34242);
nand U36962 (N_36962,N_35918,N_35119);
and U36963 (N_36963,N_34572,N_34363);
or U36964 (N_36964,N_35896,N_34461);
nand U36965 (N_36965,N_34124,N_34997);
xor U36966 (N_36966,N_34135,N_34559);
xnor U36967 (N_36967,N_34123,N_35107);
and U36968 (N_36968,N_35756,N_35582);
and U36969 (N_36969,N_34579,N_35104);
or U36970 (N_36970,N_34475,N_35139);
or U36971 (N_36971,N_34078,N_34531);
xor U36972 (N_36972,N_34108,N_35379);
and U36973 (N_36973,N_34240,N_34304);
or U36974 (N_36974,N_34610,N_34755);
nor U36975 (N_36975,N_34983,N_35052);
nor U36976 (N_36976,N_34220,N_34507);
xor U36977 (N_36977,N_35980,N_35314);
nor U36978 (N_36978,N_34975,N_35924);
nand U36979 (N_36979,N_35469,N_34965);
xnor U36980 (N_36980,N_34879,N_35231);
nor U36981 (N_36981,N_35719,N_34869);
xnor U36982 (N_36982,N_35118,N_35269);
xnor U36983 (N_36983,N_35502,N_34413);
nand U36984 (N_36984,N_35538,N_34891);
xnor U36985 (N_36985,N_34011,N_34950);
and U36986 (N_36986,N_34749,N_34142);
nor U36987 (N_36987,N_34024,N_35684);
and U36988 (N_36988,N_35640,N_35947);
and U36989 (N_36989,N_35785,N_35618);
nand U36990 (N_36990,N_34053,N_34518);
and U36991 (N_36991,N_35975,N_34065);
nand U36992 (N_36992,N_35654,N_34140);
nand U36993 (N_36993,N_34534,N_35155);
nor U36994 (N_36994,N_35891,N_35031);
xor U36995 (N_36995,N_35743,N_34984);
nor U36996 (N_36996,N_35504,N_34974);
nor U36997 (N_36997,N_34305,N_35369);
and U36998 (N_36998,N_34672,N_34843);
nor U36999 (N_36999,N_34526,N_34023);
nand U37000 (N_37000,N_34076,N_35119);
xor U37001 (N_37001,N_35560,N_34198);
nand U37002 (N_37002,N_35597,N_35107);
xnor U37003 (N_37003,N_35174,N_34554);
and U37004 (N_37004,N_35900,N_35678);
and U37005 (N_37005,N_35779,N_35671);
xor U37006 (N_37006,N_35650,N_35094);
nor U37007 (N_37007,N_35644,N_34037);
nand U37008 (N_37008,N_35954,N_35463);
xnor U37009 (N_37009,N_35619,N_35570);
or U37010 (N_37010,N_34938,N_35675);
nand U37011 (N_37011,N_34792,N_34975);
nor U37012 (N_37012,N_34043,N_34624);
nor U37013 (N_37013,N_35111,N_35062);
xnor U37014 (N_37014,N_34026,N_34423);
or U37015 (N_37015,N_35448,N_35458);
or U37016 (N_37016,N_34471,N_35379);
or U37017 (N_37017,N_34138,N_35515);
or U37018 (N_37018,N_34063,N_35326);
nor U37019 (N_37019,N_34959,N_34414);
or U37020 (N_37020,N_35211,N_34624);
nor U37021 (N_37021,N_34685,N_34011);
nor U37022 (N_37022,N_35942,N_35431);
xor U37023 (N_37023,N_34935,N_34200);
and U37024 (N_37024,N_34286,N_34907);
xor U37025 (N_37025,N_34835,N_34083);
and U37026 (N_37026,N_34858,N_35059);
and U37027 (N_37027,N_34068,N_34822);
nand U37028 (N_37028,N_34664,N_34928);
or U37029 (N_37029,N_35135,N_34114);
xnor U37030 (N_37030,N_34212,N_34276);
nand U37031 (N_37031,N_34420,N_34489);
nor U37032 (N_37032,N_35465,N_35648);
or U37033 (N_37033,N_35048,N_34472);
and U37034 (N_37034,N_34566,N_34974);
nor U37035 (N_37035,N_35231,N_34493);
nand U37036 (N_37036,N_34858,N_35544);
xnor U37037 (N_37037,N_34778,N_35506);
xor U37038 (N_37038,N_35067,N_35706);
nor U37039 (N_37039,N_35072,N_34635);
or U37040 (N_37040,N_35867,N_34286);
or U37041 (N_37041,N_35978,N_35065);
nand U37042 (N_37042,N_35167,N_34061);
and U37043 (N_37043,N_35671,N_34923);
nor U37044 (N_37044,N_35548,N_35883);
nand U37045 (N_37045,N_35482,N_35974);
or U37046 (N_37046,N_34475,N_35536);
nand U37047 (N_37047,N_35569,N_35298);
nor U37048 (N_37048,N_34270,N_35108);
xnor U37049 (N_37049,N_35016,N_34023);
xor U37050 (N_37050,N_34557,N_34731);
and U37051 (N_37051,N_35804,N_34558);
xor U37052 (N_37052,N_34498,N_34497);
or U37053 (N_37053,N_34009,N_34593);
nor U37054 (N_37054,N_35524,N_35554);
or U37055 (N_37055,N_35554,N_35799);
or U37056 (N_37056,N_34561,N_35739);
and U37057 (N_37057,N_35766,N_35962);
nor U37058 (N_37058,N_35130,N_34404);
and U37059 (N_37059,N_34662,N_35980);
and U37060 (N_37060,N_35394,N_35823);
xor U37061 (N_37061,N_34061,N_34418);
nor U37062 (N_37062,N_35243,N_35123);
xnor U37063 (N_37063,N_35165,N_34290);
xor U37064 (N_37064,N_34091,N_35816);
xor U37065 (N_37065,N_34664,N_35007);
or U37066 (N_37066,N_35044,N_35161);
and U37067 (N_37067,N_34702,N_35459);
nand U37068 (N_37068,N_35192,N_34335);
or U37069 (N_37069,N_35492,N_34301);
xor U37070 (N_37070,N_35977,N_35822);
nand U37071 (N_37071,N_35793,N_34335);
or U37072 (N_37072,N_34593,N_34246);
or U37073 (N_37073,N_34979,N_35401);
nand U37074 (N_37074,N_34493,N_35005);
nor U37075 (N_37075,N_35997,N_34233);
nand U37076 (N_37076,N_35098,N_34100);
or U37077 (N_37077,N_34577,N_35527);
xor U37078 (N_37078,N_35542,N_35701);
and U37079 (N_37079,N_34321,N_34865);
or U37080 (N_37080,N_34238,N_34360);
nand U37081 (N_37081,N_34419,N_34981);
xnor U37082 (N_37082,N_34296,N_34894);
xor U37083 (N_37083,N_34769,N_35549);
nor U37084 (N_37084,N_34567,N_34892);
xor U37085 (N_37085,N_35227,N_34177);
and U37086 (N_37086,N_34080,N_34525);
xnor U37087 (N_37087,N_35452,N_35236);
and U37088 (N_37088,N_34505,N_34565);
xnor U37089 (N_37089,N_34337,N_35689);
and U37090 (N_37090,N_34820,N_34558);
and U37091 (N_37091,N_35469,N_34553);
and U37092 (N_37092,N_34132,N_35156);
nand U37093 (N_37093,N_34842,N_35563);
nand U37094 (N_37094,N_35361,N_35321);
nor U37095 (N_37095,N_35419,N_34120);
nand U37096 (N_37096,N_34262,N_34078);
xnor U37097 (N_37097,N_35774,N_35675);
xor U37098 (N_37098,N_34440,N_34712);
or U37099 (N_37099,N_34567,N_35848);
or U37100 (N_37100,N_35683,N_34770);
xor U37101 (N_37101,N_35929,N_35930);
nand U37102 (N_37102,N_35713,N_35593);
xor U37103 (N_37103,N_34738,N_34944);
nor U37104 (N_37104,N_35819,N_35105);
nor U37105 (N_37105,N_35248,N_34212);
xnor U37106 (N_37106,N_35178,N_35221);
and U37107 (N_37107,N_35411,N_35051);
nor U37108 (N_37108,N_35746,N_34748);
and U37109 (N_37109,N_35237,N_35957);
xor U37110 (N_37110,N_34123,N_34613);
nor U37111 (N_37111,N_34474,N_34254);
nand U37112 (N_37112,N_34633,N_35194);
or U37113 (N_37113,N_34568,N_34405);
xnor U37114 (N_37114,N_34470,N_34332);
and U37115 (N_37115,N_34494,N_34774);
or U37116 (N_37116,N_35983,N_35632);
or U37117 (N_37117,N_34636,N_35120);
nand U37118 (N_37118,N_34961,N_34485);
xnor U37119 (N_37119,N_34362,N_35137);
and U37120 (N_37120,N_35949,N_34530);
nand U37121 (N_37121,N_34049,N_34506);
and U37122 (N_37122,N_34733,N_35285);
or U37123 (N_37123,N_35828,N_35904);
xor U37124 (N_37124,N_34960,N_34607);
xnor U37125 (N_37125,N_34296,N_34385);
or U37126 (N_37126,N_35951,N_34298);
xnor U37127 (N_37127,N_35928,N_34424);
or U37128 (N_37128,N_35081,N_34799);
nand U37129 (N_37129,N_35240,N_34324);
nor U37130 (N_37130,N_34148,N_34708);
or U37131 (N_37131,N_35613,N_34869);
and U37132 (N_37132,N_35077,N_35218);
nand U37133 (N_37133,N_34458,N_34553);
or U37134 (N_37134,N_35942,N_34145);
and U37135 (N_37135,N_34276,N_35996);
xor U37136 (N_37136,N_35508,N_35749);
nand U37137 (N_37137,N_35751,N_34520);
or U37138 (N_37138,N_34755,N_35238);
nand U37139 (N_37139,N_34763,N_34624);
nand U37140 (N_37140,N_34648,N_34548);
or U37141 (N_37141,N_35519,N_34927);
xor U37142 (N_37142,N_34517,N_34363);
nor U37143 (N_37143,N_35746,N_35894);
nand U37144 (N_37144,N_35765,N_34950);
nor U37145 (N_37145,N_35009,N_35478);
nor U37146 (N_37146,N_34938,N_34540);
nand U37147 (N_37147,N_35126,N_34628);
and U37148 (N_37148,N_34503,N_35121);
xor U37149 (N_37149,N_34674,N_34457);
or U37150 (N_37150,N_34007,N_34209);
nor U37151 (N_37151,N_34550,N_35239);
or U37152 (N_37152,N_34688,N_35426);
nor U37153 (N_37153,N_34079,N_35149);
nor U37154 (N_37154,N_35166,N_34356);
xor U37155 (N_37155,N_34855,N_34838);
and U37156 (N_37156,N_34542,N_34366);
nand U37157 (N_37157,N_34495,N_34916);
or U37158 (N_37158,N_35622,N_34492);
nand U37159 (N_37159,N_34493,N_35616);
and U37160 (N_37160,N_35097,N_35581);
xor U37161 (N_37161,N_35398,N_35721);
nor U37162 (N_37162,N_35012,N_34144);
or U37163 (N_37163,N_35313,N_35776);
and U37164 (N_37164,N_34160,N_35154);
nand U37165 (N_37165,N_34818,N_34396);
nand U37166 (N_37166,N_35910,N_34498);
and U37167 (N_37167,N_35819,N_34123);
nand U37168 (N_37168,N_35232,N_34580);
and U37169 (N_37169,N_35368,N_35431);
or U37170 (N_37170,N_34426,N_34165);
xnor U37171 (N_37171,N_34395,N_35951);
or U37172 (N_37172,N_34812,N_35292);
nor U37173 (N_37173,N_35542,N_35069);
nor U37174 (N_37174,N_35789,N_34449);
or U37175 (N_37175,N_34662,N_35960);
nand U37176 (N_37176,N_35586,N_34382);
nand U37177 (N_37177,N_35344,N_34157);
nor U37178 (N_37178,N_34289,N_35578);
and U37179 (N_37179,N_35065,N_34174);
and U37180 (N_37180,N_35474,N_34645);
nand U37181 (N_37181,N_34901,N_34175);
nand U37182 (N_37182,N_35789,N_35467);
nor U37183 (N_37183,N_34570,N_35103);
xnor U37184 (N_37184,N_35532,N_34511);
nand U37185 (N_37185,N_34301,N_35101);
or U37186 (N_37186,N_35665,N_35659);
xor U37187 (N_37187,N_35151,N_35513);
nor U37188 (N_37188,N_34538,N_35847);
and U37189 (N_37189,N_34875,N_34574);
and U37190 (N_37190,N_34328,N_34936);
nor U37191 (N_37191,N_35228,N_35824);
nand U37192 (N_37192,N_34837,N_34445);
or U37193 (N_37193,N_35384,N_35380);
xor U37194 (N_37194,N_34678,N_35710);
nand U37195 (N_37195,N_34291,N_35155);
or U37196 (N_37196,N_35876,N_35583);
or U37197 (N_37197,N_35921,N_35018);
nor U37198 (N_37198,N_34978,N_35302);
nor U37199 (N_37199,N_34631,N_34974);
nor U37200 (N_37200,N_35766,N_35030);
nor U37201 (N_37201,N_34299,N_35529);
or U37202 (N_37202,N_35965,N_35212);
or U37203 (N_37203,N_35166,N_35361);
or U37204 (N_37204,N_34005,N_35790);
nor U37205 (N_37205,N_34731,N_34853);
nor U37206 (N_37206,N_35902,N_35133);
xnor U37207 (N_37207,N_35107,N_34130);
xor U37208 (N_37208,N_34106,N_35573);
and U37209 (N_37209,N_35227,N_35722);
nor U37210 (N_37210,N_34442,N_35413);
xnor U37211 (N_37211,N_35232,N_35629);
and U37212 (N_37212,N_34473,N_34328);
or U37213 (N_37213,N_34820,N_35811);
nor U37214 (N_37214,N_34642,N_34606);
nor U37215 (N_37215,N_35936,N_35182);
and U37216 (N_37216,N_35306,N_35340);
and U37217 (N_37217,N_34484,N_34095);
and U37218 (N_37218,N_34794,N_34928);
xnor U37219 (N_37219,N_35893,N_35568);
nand U37220 (N_37220,N_35186,N_34464);
nor U37221 (N_37221,N_34865,N_35522);
and U37222 (N_37222,N_34687,N_35861);
nor U37223 (N_37223,N_35419,N_34848);
or U37224 (N_37224,N_34366,N_35538);
or U37225 (N_37225,N_35025,N_34746);
nor U37226 (N_37226,N_34728,N_35848);
nand U37227 (N_37227,N_34021,N_34922);
xnor U37228 (N_37228,N_34833,N_35752);
or U37229 (N_37229,N_34569,N_35100);
or U37230 (N_37230,N_35015,N_35587);
xnor U37231 (N_37231,N_34112,N_34357);
nor U37232 (N_37232,N_34840,N_35628);
or U37233 (N_37233,N_34576,N_35090);
and U37234 (N_37234,N_35034,N_34049);
xnor U37235 (N_37235,N_34985,N_34041);
nand U37236 (N_37236,N_35186,N_34481);
nand U37237 (N_37237,N_35795,N_35703);
xor U37238 (N_37238,N_34256,N_35359);
nand U37239 (N_37239,N_35796,N_35061);
nor U37240 (N_37240,N_34696,N_35833);
and U37241 (N_37241,N_35180,N_35047);
or U37242 (N_37242,N_34522,N_35739);
nand U37243 (N_37243,N_35354,N_35373);
nor U37244 (N_37244,N_35495,N_34130);
xor U37245 (N_37245,N_35009,N_34518);
xor U37246 (N_37246,N_34266,N_35368);
or U37247 (N_37247,N_34612,N_34230);
or U37248 (N_37248,N_34374,N_35733);
and U37249 (N_37249,N_35412,N_34635);
and U37250 (N_37250,N_34396,N_35097);
nor U37251 (N_37251,N_35389,N_35633);
or U37252 (N_37252,N_35063,N_35771);
and U37253 (N_37253,N_35508,N_35766);
nand U37254 (N_37254,N_35441,N_35486);
nand U37255 (N_37255,N_34784,N_35352);
nor U37256 (N_37256,N_34664,N_34668);
nand U37257 (N_37257,N_34633,N_35596);
xnor U37258 (N_37258,N_34518,N_35344);
xnor U37259 (N_37259,N_34896,N_35198);
nor U37260 (N_37260,N_35051,N_34677);
or U37261 (N_37261,N_35035,N_34080);
nand U37262 (N_37262,N_34175,N_35470);
nand U37263 (N_37263,N_34506,N_35605);
xnor U37264 (N_37264,N_35831,N_34520);
or U37265 (N_37265,N_34242,N_34519);
xnor U37266 (N_37266,N_34688,N_35609);
nor U37267 (N_37267,N_35084,N_34711);
xnor U37268 (N_37268,N_35268,N_34627);
or U37269 (N_37269,N_35770,N_34921);
nor U37270 (N_37270,N_34540,N_35096);
nor U37271 (N_37271,N_35789,N_35476);
and U37272 (N_37272,N_35736,N_35222);
xnor U37273 (N_37273,N_35457,N_35435);
or U37274 (N_37274,N_35712,N_34477);
or U37275 (N_37275,N_34622,N_35236);
and U37276 (N_37276,N_34010,N_35696);
xor U37277 (N_37277,N_34140,N_35788);
and U37278 (N_37278,N_34064,N_35375);
xor U37279 (N_37279,N_35926,N_34354);
nand U37280 (N_37280,N_34687,N_35602);
nand U37281 (N_37281,N_34299,N_34420);
nor U37282 (N_37282,N_35462,N_34437);
nor U37283 (N_37283,N_35983,N_35644);
nor U37284 (N_37284,N_35524,N_34094);
xor U37285 (N_37285,N_35816,N_34793);
xor U37286 (N_37286,N_34470,N_34593);
xor U37287 (N_37287,N_34459,N_35854);
nand U37288 (N_37288,N_34398,N_35692);
and U37289 (N_37289,N_34017,N_34754);
or U37290 (N_37290,N_35823,N_34392);
xor U37291 (N_37291,N_35456,N_34123);
nand U37292 (N_37292,N_35219,N_34308);
or U37293 (N_37293,N_35320,N_35768);
and U37294 (N_37294,N_35871,N_35640);
nor U37295 (N_37295,N_34118,N_35810);
or U37296 (N_37296,N_34841,N_35194);
xnor U37297 (N_37297,N_34159,N_34620);
and U37298 (N_37298,N_34111,N_35586);
and U37299 (N_37299,N_35280,N_35080);
or U37300 (N_37300,N_35571,N_35638);
xor U37301 (N_37301,N_35946,N_35659);
nand U37302 (N_37302,N_34225,N_35148);
xnor U37303 (N_37303,N_35970,N_34604);
or U37304 (N_37304,N_34144,N_34884);
nand U37305 (N_37305,N_34228,N_34968);
xnor U37306 (N_37306,N_34477,N_35160);
xnor U37307 (N_37307,N_34689,N_34944);
nor U37308 (N_37308,N_35749,N_35686);
nor U37309 (N_37309,N_34214,N_34447);
and U37310 (N_37310,N_35532,N_34287);
xnor U37311 (N_37311,N_35520,N_35838);
nand U37312 (N_37312,N_35175,N_34632);
and U37313 (N_37313,N_35884,N_34437);
xnor U37314 (N_37314,N_35837,N_34900);
nor U37315 (N_37315,N_35847,N_34801);
or U37316 (N_37316,N_34228,N_35430);
and U37317 (N_37317,N_35566,N_35731);
or U37318 (N_37318,N_35401,N_34397);
and U37319 (N_37319,N_35808,N_34790);
and U37320 (N_37320,N_34631,N_34220);
or U37321 (N_37321,N_35774,N_34231);
or U37322 (N_37322,N_34552,N_34779);
nand U37323 (N_37323,N_35288,N_34689);
nor U37324 (N_37324,N_34734,N_34586);
nand U37325 (N_37325,N_34547,N_34421);
nand U37326 (N_37326,N_34489,N_34179);
nand U37327 (N_37327,N_34502,N_34084);
and U37328 (N_37328,N_35468,N_35979);
nand U37329 (N_37329,N_35194,N_34996);
nand U37330 (N_37330,N_34031,N_34405);
xor U37331 (N_37331,N_35047,N_34852);
or U37332 (N_37332,N_34263,N_35148);
nor U37333 (N_37333,N_35407,N_34551);
and U37334 (N_37334,N_34620,N_34331);
nor U37335 (N_37335,N_35288,N_34619);
nand U37336 (N_37336,N_34694,N_35074);
and U37337 (N_37337,N_35083,N_34212);
nor U37338 (N_37338,N_35660,N_35023);
or U37339 (N_37339,N_34602,N_35775);
xnor U37340 (N_37340,N_35157,N_35791);
nor U37341 (N_37341,N_35788,N_34069);
xor U37342 (N_37342,N_34574,N_35713);
xor U37343 (N_37343,N_34332,N_35962);
nor U37344 (N_37344,N_34961,N_34295);
xor U37345 (N_37345,N_34221,N_35620);
nor U37346 (N_37346,N_34544,N_34112);
nor U37347 (N_37347,N_35606,N_34785);
xnor U37348 (N_37348,N_34397,N_35556);
or U37349 (N_37349,N_34541,N_35951);
or U37350 (N_37350,N_35613,N_34640);
or U37351 (N_37351,N_34028,N_35779);
nand U37352 (N_37352,N_35974,N_35104);
and U37353 (N_37353,N_35223,N_34449);
nand U37354 (N_37354,N_34986,N_35759);
nor U37355 (N_37355,N_34638,N_34556);
nand U37356 (N_37356,N_34127,N_34581);
and U37357 (N_37357,N_34844,N_34670);
nor U37358 (N_37358,N_34678,N_34985);
and U37359 (N_37359,N_34060,N_34832);
nor U37360 (N_37360,N_34625,N_35530);
xnor U37361 (N_37361,N_34034,N_34252);
or U37362 (N_37362,N_34220,N_35389);
xor U37363 (N_37363,N_35069,N_34405);
or U37364 (N_37364,N_34342,N_34244);
and U37365 (N_37365,N_34832,N_34601);
xnor U37366 (N_37366,N_35527,N_34181);
xor U37367 (N_37367,N_34942,N_34018);
or U37368 (N_37368,N_34104,N_35160);
and U37369 (N_37369,N_34231,N_35621);
nand U37370 (N_37370,N_34509,N_35411);
xnor U37371 (N_37371,N_35776,N_34328);
nor U37372 (N_37372,N_34707,N_35902);
nand U37373 (N_37373,N_34898,N_34637);
nor U37374 (N_37374,N_35894,N_34302);
xor U37375 (N_37375,N_34889,N_35901);
and U37376 (N_37376,N_34864,N_34956);
xor U37377 (N_37377,N_35817,N_34893);
nand U37378 (N_37378,N_35945,N_35421);
or U37379 (N_37379,N_35958,N_35629);
or U37380 (N_37380,N_34262,N_34788);
or U37381 (N_37381,N_35813,N_34251);
xor U37382 (N_37382,N_34215,N_34674);
nand U37383 (N_37383,N_35684,N_35291);
or U37384 (N_37384,N_35750,N_35953);
nand U37385 (N_37385,N_34088,N_34976);
nor U37386 (N_37386,N_35518,N_34395);
nor U37387 (N_37387,N_34881,N_34444);
or U37388 (N_37388,N_34706,N_35850);
nor U37389 (N_37389,N_34961,N_34393);
nor U37390 (N_37390,N_34195,N_34958);
xnor U37391 (N_37391,N_35551,N_35610);
and U37392 (N_37392,N_35278,N_34791);
xor U37393 (N_37393,N_35187,N_35327);
and U37394 (N_37394,N_35086,N_34147);
nand U37395 (N_37395,N_35650,N_35179);
and U37396 (N_37396,N_34155,N_34911);
or U37397 (N_37397,N_34584,N_34627);
and U37398 (N_37398,N_35869,N_35627);
or U37399 (N_37399,N_35749,N_34670);
nand U37400 (N_37400,N_34838,N_35247);
and U37401 (N_37401,N_34594,N_35932);
and U37402 (N_37402,N_34402,N_34455);
and U37403 (N_37403,N_34844,N_34328);
nand U37404 (N_37404,N_35670,N_35164);
xnor U37405 (N_37405,N_35489,N_34527);
xnor U37406 (N_37406,N_34627,N_34032);
and U37407 (N_37407,N_34718,N_35251);
and U37408 (N_37408,N_35146,N_34767);
xor U37409 (N_37409,N_35849,N_35598);
and U37410 (N_37410,N_35896,N_35465);
nand U37411 (N_37411,N_34423,N_35891);
or U37412 (N_37412,N_35927,N_34508);
and U37413 (N_37413,N_35754,N_35101);
and U37414 (N_37414,N_34208,N_34993);
or U37415 (N_37415,N_35063,N_35078);
and U37416 (N_37416,N_35503,N_35231);
xor U37417 (N_37417,N_35139,N_34125);
nand U37418 (N_37418,N_35730,N_35366);
nand U37419 (N_37419,N_34627,N_35132);
nand U37420 (N_37420,N_34519,N_35523);
and U37421 (N_37421,N_34863,N_35147);
or U37422 (N_37422,N_35091,N_34633);
nand U37423 (N_37423,N_34737,N_35577);
or U37424 (N_37424,N_34235,N_35427);
nand U37425 (N_37425,N_34579,N_34907);
nor U37426 (N_37426,N_35785,N_35272);
and U37427 (N_37427,N_34928,N_34580);
and U37428 (N_37428,N_35161,N_34189);
xnor U37429 (N_37429,N_35850,N_35381);
or U37430 (N_37430,N_35728,N_35913);
or U37431 (N_37431,N_34431,N_34292);
or U37432 (N_37432,N_35318,N_34544);
nand U37433 (N_37433,N_35694,N_35803);
xnor U37434 (N_37434,N_35121,N_35969);
xnor U37435 (N_37435,N_34603,N_35249);
xnor U37436 (N_37436,N_34111,N_34093);
nand U37437 (N_37437,N_34657,N_34327);
and U37438 (N_37438,N_34376,N_34270);
and U37439 (N_37439,N_35301,N_34323);
or U37440 (N_37440,N_35840,N_34853);
nand U37441 (N_37441,N_34340,N_35796);
and U37442 (N_37442,N_34401,N_35420);
and U37443 (N_37443,N_35107,N_34998);
nand U37444 (N_37444,N_34133,N_34196);
and U37445 (N_37445,N_34757,N_35080);
nand U37446 (N_37446,N_34445,N_35637);
and U37447 (N_37447,N_35365,N_34975);
or U37448 (N_37448,N_34929,N_35004);
or U37449 (N_37449,N_34307,N_35003);
nand U37450 (N_37450,N_35144,N_35492);
nand U37451 (N_37451,N_35586,N_35324);
or U37452 (N_37452,N_35675,N_34553);
nand U37453 (N_37453,N_34385,N_35035);
nand U37454 (N_37454,N_34560,N_35572);
and U37455 (N_37455,N_35820,N_35628);
nand U37456 (N_37456,N_35797,N_35609);
nor U37457 (N_37457,N_35776,N_35957);
nand U37458 (N_37458,N_35156,N_35786);
nand U37459 (N_37459,N_34266,N_35261);
xnor U37460 (N_37460,N_35779,N_35433);
nand U37461 (N_37461,N_34324,N_34655);
or U37462 (N_37462,N_34601,N_34392);
nand U37463 (N_37463,N_35928,N_35589);
nand U37464 (N_37464,N_35609,N_35325);
nand U37465 (N_37465,N_34852,N_34702);
nor U37466 (N_37466,N_34017,N_35237);
or U37467 (N_37467,N_34919,N_35576);
or U37468 (N_37468,N_35973,N_34433);
and U37469 (N_37469,N_35288,N_35112);
and U37470 (N_37470,N_34584,N_35202);
xor U37471 (N_37471,N_35327,N_35809);
or U37472 (N_37472,N_34676,N_34509);
or U37473 (N_37473,N_34174,N_34817);
nand U37474 (N_37474,N_35245,N_34968);
nand U37475 (N_37475,N_35105,N_34971);
nor U37476 (N_37476,N_35986,N_35166);
or U37477 (N_37477,N_35718,N_35586);
nor U37478 (N_37478,N_34748,N_34272);
nor U37479 (N_37479,N_35493,N_34060);
nor U37480 (N_37480,N_35288,N_34810);
or U37481 (N_37481,N_34086,N_34981);
or U37482 (N_37482,N_34585,N_35247);
xor U37483 (N_37483,N_34358,N_34753);
and U37484 (N_37484,N_35832,N_34597);
nor U37485 (N_37485,N_34840,N_34240);
nand U37486 (N_37486,N_35851,N_34098);
and U37487 (N_37487,N_34758,N_35849);
and U37488 (N_37488,N_35812,N_34274);
and U37489 (N_37489,N_35776,N_35922);
and U37490 (N_37490,N_35816,N_34356);
or U37491 (N_37491,N_34928,N_35192);
nand U37492 (N_37492,N_35935,N_34887);
or U37493 (N_37493,N_35795,N_35444);
or U37494 (N_37494,N_34909,N_35691);
or U37495 (N_37495,N_34893,N_34125);
xnor U37496 (N_37496,N_35840,N_34868);
xor U37497 (N_37497,N_35167,N_35321);
xnor U37498 (N_37498,N_35060,N_34148);
nand U37499 (N_37499,N_34792,N_34945);
or U37500 (N_37500,N_35865,N_35931);
nand U37501 (N_37501,N_34639,N_35346);
and U37502 (N_37502,N_35495,N_35999);
and U37503 (N_37503,N_35270,N_34779);
or U37504 (N_37504,N_35892,N_34407);
or U37505 (N_37505,N_34119,N_35236);
and U37506 (N_37506,N_34405,N_35897);
and U37507 (N_37507,N_34173,N_35355);
or U37508 (N_37508,N_34882,N_34275);
or U37509 (N_37509,N_35369,N_34097);
nand U37510 (N_37510,N_35984,N_35520);
nand U37511 (N_37511,N_34108,N_34931);
nand U37512 (N_37512,N_34364,N_34954);
or U37513 (N_37513,N_35158,N_35645);
nor U37514 (N_37514,N_34635,N_34586);
xor U37515 (N_37515,N_34288,N_35931);
or U37516 (N_37516,N_34835,N_34011);
and U37517 (N_37517,N_34795,N_35943);
nand U37518 (N_37518,N_35222,N_35507);
nor U37519 (N_37519,N_35607,N_34934);
nor U37520 (N_37520,N_35547,N_35781);
nor U37521 (N_37521,N_35825,N_34177);
and U37522 (N_37522,N_35644,N_34010);
xor U37523 (N_37523,N_35842,N_34434);
xnor U37524 (N_37524,N_34854,N_34384);
nand U37525 (N_37525,N_35727,N_35296);
xnor U37526 (N_37526,N_34102,N_34656);
nand U37527 (N_37527,N_34597,N_35340);
nor U37528 (N_37528,N_35802,N_35033);
nand U37529 (N_37529,N_34183,N_35943);
nand U37530 (N_37530,N_34460,N_35676);
nand U37531 (N_37531,N_34017,N_35009);
and U37532 (N_37532,N_34070,N_34807);
or U37533 (N_37533,N_35476,N_35865);
and U37534 (N_37534,N_35268,N_34761);
xnor U37535 (N_37535,N_35261,N_35447);
xor U37536 (N_37536,N_34317,N_35776);
xor U37537 (N_37537,N_34056,N_34448);
and U37538 (N_37538,N_35428,N_34319);
and U37539 (N_37539,N_35283,N_35143);
nand U37540 (N_37540,N_34413,N_35259);
or U37541 (N_37541,N_34390,N_35203);
xor U37542 (N_37542,N_34482,N_34022);
xnor U37543 (N_37543,N_34457,N_35500);
nand U37544 (N_37544,N_34367,N_35069);
and U37545 (N_37545,N_34125,N_34986);
and U37546 (N_37546,N_34080,N_34276);
xor U37547 (N_37547,N_34445,N_35452);
nor U37548 (N_37548,N_34018,N_35789);
or U37549 (N_37549,N_35599,N_35131);
nand U37550 (N_37550,N_34417,N_34363);
nand U37551 (N_37551,N_35395,N_34223);
or U37552 (N_37552,N_35938,N_34482);
xnor U37553 (N_37553,N_35365,N_34701);
nand U37554 (N_37554,N_34805,N_34795);
nor U37555 (N_37555,N_34526,N_35641);
xor U37556 (N_37556,N_34583,N_34651);
xor U37557 (N_37557,N_34950,N_34734);
xnor U37558 (N_37558,N_34980,N_34246);
or U37559 (N_37559,N_35863,N_34625);
or U37560 (N_37560,N_34976,N_34344);
xnor U37561 (N_37561,N_34580,N_35642);
and U37562 (N_37562,N_34279,N_34289);
and U37563 (N_37563,N_35164,N_34972);
xor U37564 (N_37564,N_35723,N_34531);
and U37565 (N_37565,N_34018,N_34699);
nand U37566 (N_37566,N_35065,N_35730);
nand U37567 (N_37567,N_34235,N_35387);
xor U37568 (N_37568,N_34328,N_35710);
xnor U37569 (N_37569,N_34401,N_35177);
or U37570 (N_37570,N_35523,N_34859);
nor U37571 (N_37571,N_34030,N_35442);
nand U37572 (N_37572,N_34924,N_35015);
and U37573 (N_37573,N_34269,N_35956);
or U37574 (N_37574,N_34936,N_35258);
xor U37575 (N_37575,N_34842,N_35245);
nor U37576 (N_37576,N_35413,N_35820);
and U37577 (N_37577,N_35464,N_34428);
or U37578 (N_37578,N_34026,N_35064);
nand U37579 (N_37579,N_34854,N_35158);
nand U37580 (N_37580,N_35846,N_35222);
and U37581 (N_37581,N_34024,N_35768);
nand U37582 (N_37582,N_35712,N_34843);
and U37583 (N_37583,N_35100,N_34291);
nand U37584 (N_37584,N_34895,N_35762);
nand U37585 (N_37585,N_34876,N_34502);
xor U37586 (N_37586,N_35167,N_34218);
nor U37587 (N_37587,N_34044,N_34341);
and U37588 (N_37588,N_35190,N_35023);
nand U37589 (N_37589,N_34066,N_34418);
nor U37590 (N_37590,N_35979,N_34281);
nand U37591 (N_37591,N_35534,N_35940);
or U37592 (N_37592,N_35752,N_34459);
and U37593 (N_37593,N_35622,N_35201);
or U37594 (N_37594,N_35274,N_34004);
and U37595 (N_37595,N_34031,N_35850);
nand U37596 (N_37596,N_35234,N_35323);
nor U37597 (N_37597,N_35316,N_34842);
nand U37598 (N_37598,N_34502,N_34836);
xor U37599 (N_37599,N_35800,N_35368);
xnor U37600 (N_37600,N_34017,N_34992);
and U37601 (N_37601,N_35477,N_35687);
or U37602 (N_37602,N_35699,N_35293);
or U37603 (N_37603,N_34461,N_34816);
and U37604 (N_37604,N_34868,N_34027);
and U37605 (N_37605,N_34342,N_34734);
nor U37606 (N_37606,N_34409,N_34877);
and U37607 (N_37607,N_35594,N_35713);
nor U37608 (N_37608,N_34211,N_35092);
or U37609 (N_37609,N_35750,N_34393);
nand U37610 (N_37610,N_35045,N_35809);
nand U37611 (N_37611,N_34296,N_35155);
nor U37612 (N_37612,N_34066,N_34567);
nor U37613 (N_37613,N_35340,N_35569);
xor U37614 (N_37614,N_35336,N_34951);
nand U37615 (N_37615,N_34056,N_35852);
or U37616 (N_37616,N_35484,N_34381);
xor U37617 (N_37617,N_35853,N_34000);
nor U37618 (N_37618,N_35502,N_35563);
nor U37619 (N_37619,N_35428,N_34467);
xor U37620 (N_37620,N_34251,N_35354);
or U37621 (N_37621,N_34049,N_35267);
and U37622 (N_37622,N_35158,N_34492);
xnor U37623 (N_37623,N_34481,N_35811);
and U37624 (N_37624,N_34749,N_34770);
nor U37625 (N_37625,N_34697,N_34894);
and U37626 (N_37626,N_34337,N_34460);
nor U37627 (N_37627,N_35726,N_34809);
and U37628 (N_37628,N_35076,N_35890);
or U37629 (N_37629,N_35029,N_34844);
nor U37630 (N_37630,N_35875,N_34318);
nor U37631 (N_37631,N_35518,N_35092);
xnor U37632 (N_37632,N_35456,N_34052);
or U37633 (N_37633,N_34851,N_34980);
and U37634 (N_37634,N_34963,N_35118);
nand U37635 (N_37635,N_34965,N_35380);
and U37636 (N_37636,N_34026,N_34413);
or U37637 (N_37637,N_35412,N_34588);
xnor U37638 (N_37638,N_34511,N_34402);
and U37639 (N_37639,N_34150,N_35869);
xor U37640 (N_37640,N_34626,N_35649);
or U37641 (N_37641,N_35047,N_35725);
or U37642 (N_37642,N_34286,N_34413);
and U37643 (N_37643,N_35042,N_34800);
and U37644 (N_37644,N_34201,N_34056);
xor U37645 (N_37645,N_35562,N_35694);
nor U37646 (N_37646,N_35182,N_34167);
nor U37647 (N_37647,N_35007,N_35711);
xor U37648 (N_37648,N_35875,N_34633);
xor U37649 (N_37649,N_35042,N_34949);
xnor U37650 (N_37650,N_34302,N_34622);
nor U37651 (N_37651,N_34992,N_34150);
nor U37652 (N_37652,N_34426,N_35524);
xnor U37653 (N_37653,N_34022,N_35196);
xor U37654 (N_37654,N_34683,N_35171);
or U37655 (N_37655,N_35630,N_35278);
or U37656 (N_37656,N_34926,N_34778);
and U37657 (N_37657,N_34299,N_35755);
nand U37658 (N_37658,N_35451,N_35497);
or U37659 (N_37659,N_34805,N_35511);
and U37660 (N_37660,N_34038,N_34204);
nor U37661 (N_37661,N_35714,N_34160);
or U37662 (N_37662,N_34276,N_34180);
or U37663 (N_37663,N_34895,N_35014);
nand U37664 (N_37664,N_34430,N_35505);
nand U37665 (N_37665,N_35990,N_34840);
nand U37666 (N_37666,N_35517,N_35732);
or U37667 (N_37667,N_35203,N_35607);
xnor U37668 (N_37668,N_34904,N_35577);
xnor U37669 (N_37669,N_35440,N_34973);
xor U37670 (N_37670,N_35001,N_34062);
or U37671 (N_37671,N_35111,N_34374);
or U37672 (N_37672,N_34101,N_34636);
or U37673 (N_37673,N_34486,N_34525);
xor U37674 (N_37674,N_34522,N_34767);
nand U37675 (N_37675,N_35740,N_35830);
xnor U37676 (N_37676,N_35780,N_34316);
nor U37677 (N_37677,N_35612,N_35640);
nand U37678 (N_37678,N_34147,N_35977);
xnor U37679 (N_37679,N_34232,N_35015);
nand U37680 (N_37680,N_35249,N_34511);
nand U37681 (N_37681,N_34075,N_34806);
nand U37682 (N_37682,N_35031,N_35065);
nand U37683 (N_37683,N_34091,N_34473);
nor U37684 (N_37684,N_34247,N_35443);
nor U37685 (N_37685,N_35160,N_34346);
nand U37686 (N_37686,N_34365,N_34012);
nor U37687 (N_37687,N_35255,N_35783);
and U37688 (N_37688,N_34696,N_35837);
nor U37689 (N_37689,N_34040,N_35716);
nor U37690 (N_37690,N_34629,N_34027);
or U37691 (N_37691,N_35044,N_34526);
and U37692 (N_37692,N_35721,N_34993);
nand U37693 (N_37693,N_34383,N_34755);
nor U37694 (N_37694,N_34111,N_34479);
xnor U37695 (N_37695,N_34299,N_35356);
and U37696 (N_37696,N_35481,N_35110);
and U37697 (N_37697,N_34811,N_35533);
or U37698 (N_37698,N_35204,N_34080);
and U37699 (N_37699,N_34627,N_35872);
nand U37700 (N_37700,N_35600,N_35442);
nor U37701 (N_37701,N_34533,N_35255);
or U37702 (N_37702,N_35203,N_34184);
xnor U37703 (N_37703,N_35168,N_34699);
and U37704 (N_37704,N_34522,N_34981);
nand U37705 (N_37705,N_35688,N_34710);
or U37706 (N_37706,N_34730,N_35204);
nor U37707 (N_37707,N_35281,N_35280);
and U37708 (N_37708,N_35876,N_34136);
nand U37709 (N_37709,N_34601,N_34679);
and U37710 (N_37710,N_35986,N_35753);
and U37711 (N_37711,N_34185,N_34983);
xnor U37712 (N_37712,N_35966,N_34725);
nand U37713 (N_37713,N_35102,N_35001);
xor U37714 (N_37714,N_35158,N_34931);
or U37715 (N_37715,N_35339,N_35186);
and U37716 (N_37716,N_35911,N_34179);
nor U37717 (N_37717,N_35148,N_35404);
and U37718 (N_37718,N_34228,N_34510);
or U37719 (N_37719,N_34656,N_35665);
nor U37720 (N_37720,N_35760,N_35127);
and U37721 (N_37721,N_35972,N_34361);
xor U37722 (N_37722,N_35901,N_35871);
or U37723 (N_37723,N_34672,N_35637);
or U37724 (N_37724,N_35784,N_35132);
nor U37725 (N_37725,N_35493,N_35812);
nor U37726 (N_37726,N_34633,N_35558);
nor U37727 (N_37727,N_35306,N_35999);
xor U37728 (N_37728,N_35632,N_35168);
and U37729 (N_37729,N_34910,N_35040);
xnor U37730 (N_37730,N_34446,N_34007);
or U37731 (N_37731,N_34762,N_35356);
and U37732 (N_37732,N_34861,N_35294);
or U37733 (N_37733,N_34482,N_34768);
and U37734 (N_37734,N_34394,N_35828);
and U37735 (N_37735,N_34105,N_34798);
xor U37736 (N_37736,N_34512,N_35351);
nor U37737 (N_37737,N_35680,N_34552);
xor U37738 (N_37738,N_34595,N_35629);
or U37739 (N_37739,N_34221,N_35627);
xnor U37740 (N_37740,N_34529,N_34759);
and U37741 (N_37741,N_35837,N_34785);
and U37742 (N_37742,N_34389,N_35594);
nor U37743 (N_37743,N_34439,N_34144);
xor U37744 (N_37744,N_35542,N_35682);
nor U37745 (N_37745,N_35932,N_34066);
and U37746 (N_37746,N_35828,N_35527);
and U37747 (N_37747,N_35232,N_34222);
nand U37748 (N_37748,N_34478,N_34971);
and U37749 (N_37749,N_34075,N_35309);
or U37750 (N_37750,N_35784,N_35794);
nor U37751 (N_37751,N_35029,N_35609);
nor U37752 (N_37752,N_34365,N_35034);
or U37753 (N_37753,N_34425,N_34931);
nand U37754 (N_37754,N_35371,N_35508);
xor U37755 (N_37755,N_35195,N_35321);
nand U37756 (N_37756,N_35297,N_34852);
nor U37757 (N_37757,N_34419,N_35974);
nor U37758 (N_37758,N_35743,N_34626);
nand U37759 (N_37759,N_35745,N_34909);
nand U37760 (N_37760,N_34950,N_35466);
nor U37761 (N_37761,N_34275,N_34502);
and U37762 (N_37762,N_35123,N_35554);
nor U37763 (N_37763,N_34587,N_35399);
nor U37764 (N_37764,N_35818,N_35706);
nand U37765 (N_37765,N_35747,N_35168);
or U37766 (N_37766,N_35891,N_34625);
nand U37767 (N_37767,N_35039,N_35335);
xnor U37768 (N_37768,N_34431,N_35776);
xor U37769 (N_37769,N_34038,N_35107);
and U37770 (N_37770,N_35636,N_35987);
xor U37771 (N_37771,N_34861,N_35509);
or U37772 (N_37772,N_35873,N_34565);
nand U37773 (N_37773,N_35227,N_34850);
nor U37774 (N_37774,N_35957,N_35769);
nand U37775 (N_37775,N_35723,N_34499);
xor U37776 (N_37776,N_35681,N_35662);
nand U37777 (N_37777,N_34335,N_35657);
and U37778 (N_37778,N_35726,N_34639);
nand U37779 (N_37779,N_35295,N_34162);
nand U37780 (N_37780,N_35244,N_35107);
xor U37781 (N_37781,N_35238,N_35977);
nor U37782 (N_37782,N_35085,N_35919);
or U37783 (N_37783,N_34483,N_34070);
or U37784 (N_37784,N_34842,N_35656);
xor U37785 (N_37785,N_34663,N_35363);
or U37786 (N_37786,N_34038,N_34319);
and U37787 (N_37787,N_35424,N_35836);
xor U37788 (N_37788,N_35504,N_34646);
and U37789 (N_37789,N_34758,N_35131);
or U37790 (N_37790,N_34679,N_34547);
and U37791 (N_37791,N_34598,N_34273);
and U37792 (N_37792,N_35864,N_34091);
and U37793 (N_37793,N_35468,N_35464);
xnor U37794 (N_37794,N_35674,N_34579);
nand U37795 (N_37795,N_35395,N_35673);
or U37796 (N_37796,N_35943,N_34860);
nor U37797 (N_37797,N_35212,N_34925);
nand U37798 (N_37798,N_35357,N_35324);
and U37799 (N_37799,N_34427,N_35201);
xor U37800 (N_37800,N_35939,N_34902);
xor U37801 (N_37801,N_35665,N_35243);
xnor U37802 (N_37802,N_34045,N_34216);
or U37803 (N_37803,N_35422,N_34950);
or U37804 (N_37804,N_35530,N_34976);
nand U37805 (N_37805,N_35720,N_34546);
or U37806 (N_37806,N_35798,N_34834);
xor U37807 (N_37807,N_34490,N_35917);
nand U37808 (N_37808,N_34059,N_35571);
xor U37809 (N_37809,N_35604,N_35683);
nor U37810 (N_37810,N_34193,N_34848);
nor U37811 (N_37811,N_35070,N_35957);
nand U37812 (N_37812,N_34193,N_34367);
nand U37813 (N_37813,N_34956,N_34160);
nor U37814 (N_37814,N_34524,N_35248);
xnor U37815 (N_37815,N_34072,N_34163);
nor U37816 (N_37816,N_34555,N_35042);
nand U37817 (N_37817,N_35531,N_34294);
nor U37818 (N_37818,N_35329,N_35893);
or U37819 (N_37819,N_34471,N_34266);
or U37820 (N_37820,N_35489,N_34265);
and U37821 (N_37821,N_34162,N_35694);
and U37822 (N_37822,N_34019,N_35762);
nand U37823 (N_37823,N_34235,N_35323);
nor U37824 (N_37824,N_34655,N_35275);
nand U37825 (N_37825,N_35069,N_35418);
xor U37826 (N_37826,N_34538,N_34534);
nor U37827 (N_37827,N_35928,N_34701);
nand U37828 (N_37828,N_35246,N_34042);
nor U37829 (N_37829,N_34553,N_34935);
nand U37830 (N_37830,N_35008,N_34581);
nand U37831 (N_37831,N_35693,N_35561);
xnor U37832 (N_37832,N_34709,N_34246);
or U37833 (N_37833,N_35008,N_34951);
nand U37834 (N_37834,N_35331,N_35421);
nand U37835 (N_37835,N_34639,N_35988);
and U37836 (N_37836,N_35560,N_35438);
nand U37837 (N_37837,N_35495,N_35789);
and U37838 (N_37838,N_34490,N_35849);
and U37839 (N_37839,N_35170,N_35260);
nand U37840 (N_37840,N_35677,N_35960);
xnor U37841 (N_37841,N_34901,N_35178);
and U37842 (N_37842,N_35315,N_34111);
or U37843 (N_37843,N_34648,N_35747);
and U37844 (N_37844,N_35467,N_34371);
nand U37845 (N_37845,N_34096,N_34199);
and U37846 (N_37846,N_34356,N_35557);
nor U37847 (N_37847,N_35091,N_34070);
and U37848 (N_37848,N_34580,N_34785);
or U37849 (N_37849,N_35316,N_35230);
or U37850 (N_37850,N_35604,N_35241);
or U37851 (N_37851,N_35450,N_35932);
or U37852 (N_37852,N_34152,N_34894);
nand U37853 (N_37853,N_34859,N_34639);
and U37854 (N_37854,N_34699,N_34747);
nor U37855 (N_37855,N_35590,N_35454);
or U37856 (N_37856,N_35825,N_34099);
nand U37857 (N_37857,N_35833,N_35404);
nor U37858 (N_37858,N_35560,N_35841);
nor U37859 (N_37859,N_34507,N_35395);
or U37860 (N_37860,N_34271,N_34913);
nand U37861 (N_37861,N_35909,N_34017);
nor U37862 (N_37862,N_35333,N_35113);
xnor U37863 (N_37863,N_34475,N_34753);
or U37864 (N_37864,N_34195,N_34214);
xor U37865 (N_37865,N_35556,N_35602);
nor U37866 (N_37866,N_34295,N_35901);
xor U37867 (N_37867,N_34594,N_35507);
or U37868 (N_37868,N_34413,N_35999);
nand U37869 (N_37869,N_34520,N_34449);
xor U37870 (N_37870,N_35267,N_35171);
xnor U37871 (N_37871,N_34424,N_35749);
xnor U37872 (N_37872,N_35736,N_34412);
xnor U37873 (N_37873,N_34471,N_34881);
or U37874 (N_37874,N_34473,N_35960);
or U37875 (N_37875,N_35982,N_35952);
and U37876 (N_37876,N_35484,N_34329);
and U37877 (N_37877,N_35504,N_35469);
and U37878 (N_37878,N_34244,N_34192);
nand U37879 (N_37879,N_35670,N_34158);
and U37880 (N_37880,N_34130,N_34770);
or U37881 (N_37881,N_34501,N_34202);
or U37882 (N_37882,N_34521,N_34152);
nand U37883 (N_37883,N_34177,N_35733);
or U37884 (N_37884,N_35877,N_35048);
xor U37885 (N_37885,N_34632,N_35995);
and U37886 (N_37886,N_35148,N_34886);
nand U37887 (N_37887,N_34049,N_35335);
xnor U37888 (N_37888,N_34250,N_35283);
xor U37889 (N_37889,N_34274,N_34147);
nor U37890 (N_37890,N_35864,N_34525);
and U37891 (N_37891,N_34931,N_35364);
nor U37892 (N_37892,N_34564,N_34980);
and U37893 (N_37893,N_35572,N_34476);
xor U37894 (N_37894,N_35632,N_35385);
nor U37895 (N_37895,N_35653,N_35699);
or U37896 (N_37896,N_35472,N_35538);
nand U37897 (N_37897,N_34028,N_35869);
and U37898 (N_37898,N_34210,N_35473);
nand U37899 (N_37899,N_34194,N_35247);
nand U37900 (N_37900,N_34080,N_34103);
and U37901 (N_37901,N_34586,N_35016);
xnor U37902 (N_37902,N_34488,N_35792);
nor U37903 (N_37903,N_34080,N_35609);
nor U37904 (N_37904,N_34480,N_34680);
or U37905 (N_37905,N_34240,N_34802);
xor U37906 (N_37906,N_34105,N_35245);
and U37907 (N_37907,N_35778,N_34426);
nor U37908 (N_37908,N_34695,N_35753);
nor U37909 (N_37909,N_34807,N_35611);
xor U37910 (N_37910,N_35097,N_35971);
xnor U37911 (N_37911,N_35854,N_35277);
xnor U37912 (N_37912,N_34907,N_35711);
or U37913 (N_37913,N_34957,N_35684);
and U37914 (N_37914,N_34108,N_35264);
xor U37915 (N_37915,N_34689,N_34894);
or U37916 (N_37916,N_35706,N_34677);
xor U37917 (N_37917,N_34296,N_34170);
or U37918 (N_37918,N_34273,N_34091);
and U37919 (N_37919,N_35949,N_34890);
xor U37920 (N_37920,N_35765,N_34549);
nand U37921 (N_37921,N_35462,N_34470);
or U37922 (N_37922,N_34078,N_34915);
nor U37923 (N_37923,N_35349,N_34562);
nand U37924 (N_37924,N_34683,N_35027);
nand U37925 (N_37925,N_34575,N_35963);
nor U37926 (N_37926,N_34013,N_35183);
and U37927 (N_37927,N_35926,N_35152);
nor U37928 (N_37928,N_34556,N_34147);
xnor U37929 (N_37929,N_34023,N_35283);
xor U37930 (N_37930,N_34624,N_35152);
and U37931 (N_37931,N_34901,N_35794);
nor U37932 (N_37932,N_34630,N_34777);
nand U37933 (N_37933,N_35993,N_35422);
or U37934 (N_37934,N_35838,N_35248);
or U37935 (N_37935,N_35728,N_34908);
and U37936 (N_37936,N_34396,N_34830);
nor U37937 (N_37937,N_35071,N_35508);
nor U37938 (N_37938,N_35825,N_35849);
nand U37939 (N_37939,N_35492,N_34324);
and U37940 (N_37940,N_35323,N_34371);
and U37941 (N_37941,N_35801,N_34027);
nand U37942 (N_37942,N_35473,N_35072);
and U37943 (N_37943,N_35279,N_35125);
nand U37944 (N_37944,N_34568,N_34159);
and U37945 (N_37945,N_35948,N_35547);
nor U37946 (N_37946,N_35238,N_35938);
nand U37947 (N_37947,N_35460,N_34356);
nand U37948 (N_37948,N_34082,N_35147);
nor U37949 (N_37949,N_35503,N_34978);
or U37950 (N_37950,N_34975,N_35983);
nor U37951 (N_37951,N_34241,N_34659);
xor U37952 (N_37952,N_35055,N_34875);
nor U37953 (N_37953,N_34297,N_34849);
or U37954 (N_37954,N_35479,N_35347);
xor U37955 (N_37955,N_34988,N_34198);
xor U37956 (N_37956,N_34396,N_35473);
or U37957 (N_37957,N_34939,N_34026);
nor U37958 (N_37958,N_34913,N_34164);
nor U37959 (N_37959,N_34437,N_34861);
nand U37960 (N_37960,N_34330,N_34706);
and U37961 (N_37961,N_35101,N_34315);
and U37962 (N_37962,N_34330,N_34011);
and U37963 (N_37963,N_35249,N_34955);
nor U37964 (N_37964,N_34937,N_34180);
xnor U37965 (N_37965,N_35638,N_35579);
or U37966 (N_37966,N_34912,N_34457);
xor U37967 (N_37967,N_34540,N_35119);
xnor U37968 (N_37968,N_34752,N_34840);
and U37969 (N_37969,N_35379,N_34528);
nor U37970 (N_37970,N_35281,N_35929);
and U37971 (N_37971,N_34374,N_35381);
and U37972 (N_37972,N_35948,N_34547);
xnor U37973 (N_37973,N_34683,N_34269);
nand U37974 (N_37974,N_34151,N_35065);
nor U37975 (N_37975,N_34478,N_34236);
and U37976 (N_37976,N_35021,N_34327);
and U37977 (N_37977,N_34133,N_34851);
nor U37978 (N_37978,N_34040,N_34876);
or U37979 (N_37979,N_34498,N_35957);
and U37980 (N_37980,N_34261,N_35727);
and U37981 (N_37981,N_34320,N_35774);
or U37982 (N_37982,N_34089,N_35419);
nor U37983 (N_37983,N_35237,N_34886);
and U37984 (N_37984,N_35731,N_35367);
or U37985 (N_37985,N_34722,N_35361);
nor U37986 (N_37986,N_35724,N_35766);
nand U37987 (N_37987,N_34554,N_35295);
nor U37988 (N_37988,N_35600,N_35872);
nand U37989 (N_37989,N_34668,N_35022);
nor U37990 (N_37990,N_35245,N_34550);
and U37991 (N_37991,N_35145,N_35890);
xnor U37992 (N_37992,N_35314,N_34125);
nand U37993 (N_37993,N_34406,N_34449);
xnor U37994 (N_37994,N_35483,N_34148);
nand U37995 (N_37995,N_35261,N_34260);
and U37996 (N_37996,N_35665,N_34129);
nor U37997 (N_37997,N_35785,N_35397);
nor U37998 (N_37998,N_35677,N_35595);
nand U37999 (N_37999,N_35122,N_35352);
or U38000 (N_38000,N_37807,N_36673);
nor U38001 (N_38001,N_37446,N_37061);
nand U38002 (N_38002,N_37860,N_37110);
and U38003 (N_38003,N_36963,N_36439);
xnor U38004 (N_38004,N_36044,N_37408);
xnor U38005 (N_38005,N_36682,N_36042);
nor U38006 (N_38006,N_36412,N_36814);
xor U38007 (N_38007,N_37421,N_36718);
or U38008 (N_38008,N_36983,N_37868);
or U38009 (N_38009,N_37968,N_36293);
nand U38010 (N_38010,N_37808,N_36864);
xnor U38011 (N_38011,N_37412,N_36206);
nor U38012 (N_38012,N_37152,N_37322);
xnor U38013 (N_38013,N_37158,N_36394);
nand U38014 (N_38014,N_36062,N_37383);
nand U38015 (N_38015,N_36888,N_37320);
and U38016 (N_38016,N_36144,N_36286);
xor U38017 (N_38017,N_36798,N_36582);
nor U38018 (N_38018,N_36707,N_37688);
nand U38019 (N_38019,N_37019,N_36020);
and U38020 (N_38020,N_37715,N_36895);
xnor U38021 (N_38021,N_37148,N_36391);
nor U38022 (N_38022,N_36027,N_36744);
nor U38023 (N_38023,N_36498,N_37284);
or U38024 (N_38024,N_37310,N_37568);
or U38025 (N_38025,N_37083,N_36292);
nand U38026 (N_38026,N_37658,N_36843);
nand U38027 (N_38027,N_36420,N_37525);
nand U38028 (N_38028,N_36546,N_37800);
and U38029 (N_38029,N_37896,N_36052);
and U38030 (N_38030,N_36087,N_37544);
or U38031 (N_38031,N_37983,N_37269);
xnor U38032 (N_38032,N_37345,N_37413);
nand U38033 (N_38033,N_36540,N_37925);
and U38034 (N_38034,N_37793,N_37156);
nand U38035 (N_38035,N_36759,N_37393);
or U38036 (N_38036,N_36821,N_36926);
and U38037 (N_38037,N_36453,N_36897);
and U38038 (N_38038,N_36082,N_37614);
or U38039 (N_38039,N_37077,N_37048);
nor U38040 (N_38040,N_36916,N_37669);
or U38041 (N_38041,N_37832,N_36143);
nand U38042 (N_38042,N_37044,N_36681);
nand U38043 (N_38043,N_37670,N_36525);
nor U38044 (N_38044,N_37327,N_37580);
nand U38045 (N_38045,N_37897,N_37711);
or U38046 (N_38046,N_36696,N_36005);
xor U38047 (N_38047,N_37037,N_37713);
nor U38048 (N_38048,N_36088,N_37543);
nand U38049 (N_38049,N_36697,N_37536);
or U38050 (N_38050,N_36627,N_36162);
nand U38051 (N_38051,N_37623,N_37141);
xnor U38052 (N_38052,N_37861,N_36454);
and U38053 (N_38053,N_37038,N_36543);
nand U38054 (N_38054,N_36380,N_37557);
or U38055 (N_38055,N_37958,N_36428);
nand U38056 (N_38056,N_36958,N_37240);
nor U38057 (N_38057,N_37749,N_36830);
or U38058 (N_38058,N_37231,N_36319);
nor U38059 (N_38059,N_37755,N_36317);
xor U38060 (N_38060,N_36522,N_37782);
and U38061 (N_38061,N_37694,N_36155);
xnor U38062 (N_38062,N_36145,N_37729);
or U38063 (N_38063,N_37023,N_37654);
and U38064 (N_38064,N_36877,N_36616);
nand U38065 (N_38065,N_36652,N_36947);
nand U38066 (N_38066,N_37217,N_36887);
nor U38067 (N_38067,N_36995,N_37584);
xnor U38068 (N_38068,N_36869,N_37313);
and U38069 (N_38069,N_36692,N_37632);
and U38070 (N_38070,N_37407,N_37656);
and U38071 (N_38071,N_36844,N_37373);
nand U38072 (N_38072,N_36054,N_37912);
xor U38073 (N_38073,N_36743,N_37733);
and U38074 (N_38074,N_36306,N_37548);
xnor U38075 (N_38075,N_37066,N_36415);
nand U38076 (N_38076,N_37996,N_37640);
nor U38077 (N_38077,N_37503,N_36955);
xnor U38078 (N_38078,N_36418,N_37603);
nor U38079 (N_38079,N_36545,N_36621);
xnor U38080 (N_38080,N_37707,N_36429);
and U38081 (N_38081,N_37131,N_36819);
and U38082 (N_38082,N_37082,N_37053);
nand U38083 (N_38083,N_37326,N_37232);
and U38084 (N_38084,N_36960,N_36247);
nand U38085 (N_38085,N_36379,N_36455);
or U38086 (N_38086,N_37520,N_36303);
and U38087 (N_38087,N_37414,N_37368);
nor U38088 (N_38088,N_37797,N_37234);
xnor U38089 (N_38089,N_36185,N_36700);
nand U38090 (N_38090,N_37888,N_37224);
nand U38091 (N_38091,N_36631,N_37840);
and U38092 (N_38092,N_37325,N_36767);
xor U38093 (N_38093,N_36749,N_37559);
nor U38094 (N_38094,N_37831,N_37722);
and U38095 (N_38095,N_37033,N_36972);
xnor U38096 (N_38096,N_36358,N_36755);
nor U38097 (N_38097,N_37659,N_37998);
and U38098 (N_38098,N_36776,N_37975);
xor U38099 (N_38099,N_36867,N_36056);
nand U38100 (N_38100,N_37128,N_36261);
nand U38101 (N_38101,N_36126,N_37978);
or U38102 (N_38102,N_37646,N_36831);
xor U38103 (N_38103,N_36084,N_36530);
or U38104 (N_38104,N_36239,N_36297);
nor U38105 (N_38105,N_36740,N_37071);
and U38106 (N_38106,N_36721,N_36752);
nand U38107 (N_38107,N_36271,N_36413);
or U38108 (N_38108,N_36459,N_36290);
nor U38109 (N_38109,N_36851,N_36124);
nor U38110 (N_38110,N_37622,N_37505);
nand U38111 (N_38111,N_37389,N_37226);
xnor U38112 (N_38112,N_37332,N_36366);
nand U38113 (N_38113,N_37146,N_37428);
xor U38114 (N_38114,N_36966,N_37118);
nand U38115 (N_38115,N_36430,N_37261);
nor U38116 (N_38116,N_37067,N_36649);
nor U38117 (N_38117,N_36770,N_37573);
xnor U38118 (N_38118,N_36002,N_36702);
nor U38119 (N_38119,N_37107,N_36818);
and U38120 (N_38120,N_36160,N_36148);
and U38121 (N_38121,N_36985,N_37330);
and U38122 (N_38122,N_36894,N_36233);
and U38123 (N_38123,N_37369,N_37238);
nor U38124 (N_38124,N_37866,N_37171);
nand U38125 (N_38125,N_36528,N_36859);
and U38126 (N_38126,N_37180,N_37089);
xnor U38127 (N_38127,N_37305,N_36348);
nand U38128 (N_38128,N_36965,N_37449);
and U38129 (N_38129,N_36324,N_37980);
nor U38130 (N_38130,N_36092,N_37528);
or U38131 (N_38131,N_36023,N_37365);
and U38132 (N_38132,N_36167,N_37678);
or U38133 (N_38133,N_37040,N_37469);
and U38134 (N_38134,N_36884,N_36999);
nand U38135 (N_38135,N_36209,N_37161);
nor U38136 (N_38136,N_37982,N_37426);
xnor U38137 (N_38137,N_37781,N_36450);
or U38138 (N_38138,N_36009,N_37484);
and U38139 (N_38139,N_37768,N_36376);
or U38140 (N_38140,N_37395,N_36834);
nor U38141 (N_38141,N_37457,N_36706);
xnor U38142 (N_38142,N_36152,N_37168);
or U38143 (N_38143,N_37600,N_36437);
xor U38144 (N_38144,N_36769,N_36714);
nor U38145 (N_38145,N_37598,N_37579);
or U38146 (N_38146,N_36069,N_37386);
nor U38147 (N_38147,N_37164,N_36355);
nor U38148 (N_38148,N_37064,N_37283);
nor U38149 (N_38149,N_37054,N_36080);
and U38150 (N_38150,N_36774,N_36182);
nor U38151 (N_38151,N_36789,N_37836);
nand U38152 (N_38152,N_37361,N_37346);
nand U38153 (N_38153,N_36363,N_36795);
or U38154 (N_38154,N_37194,N_36125);
and U38155 (N_38155,N_37250,N_37591);
and U38156 (N_38156,N_37416,N_37576);
and U38157 (N_38157,N_36846,N_37889);
and U38158 (N_38158,N_36403,N_37092);
nand U38159 (N_38159,N_36733,N_36384);
nor U38160 (N_38160,N_37051,N_37055);
and U38161 (N_38161,N_37404,N_36989);
nand U38162 (N_38162,N_37069,N_37328);
nor U38163 (N_38163,N_36090,N_36485);
nor U38164 (N_38164,N_37550,N_37356);
xor U38165 (N_38165,N_37597,N_36328);
or U38166 (N_38166,N_36414,N_36529);
or U38167 (N_38167,N_37415,N_37956);
nand U38168 (N_38168,N_37561,N_36109);
xnor U38169 (N_38169,N_37186,N_37321);
nor U38170 (N_38170,N_37593,N_37191);
or U38171 (N_38171,N_37913,N_36077);
nor U38172 (N_38172,N_37391,N_37564);
nand U38173 (N_38173,N_37728,N_36745);
or U38174 (N_38174,N_37594,N_37621);
nor U38175 (N_38175,N_36663,N_36138);
xnor U38176 (N_38176,N_37792,N_37482);
xnor U38177 (N_38177,N_36557,N_36661);
or U38178 (N_38178,N_36093,N_37644);
nor U38179 (N_38179,N_37377,N_36256);
nor U38180 (N_38180,N_36189,N_37605);
xnor U38181 (N_38181,N_37318,N_36808);
or U38182 (N_38182,N_36288,N_36208);
xor U38183 (N_38183,N_36478,N_37878);
nand U38184 (N_38184,N_37466,N_36606);
and U38185 (N_38185,N_37075,N_37843);
and U38186 (N_38186,N_36953,N_36722);
and U38187 (N_38187,N_37085,N_36365);
xor U38188 (N_38188,N_36526,N_37298);
nand U38189 (N_38189,N_37279,N_36374);
and U38190 (N_38190,N_36875,N_36603);
or U38191 (N_38191,N_36460,N_37246);
and U38192 (N_38192,N_37296,N_36154);
xnor U38193 (N_38193,N_36600,N_37409);
nand U38194 (N_38194,N_37462,N_36993);
nand U38195 (N_38195,N_37572,N_36704);
and U38196 (N_38196,N_37215,N_37448);
nor U38197 (N_38197,N_36194,N_36248);
or U38198 (N_38198,N_37187,N_36572);
nand U38199 (N_38199,N_37166,N_37264);
or U38200 (N_38200,N_37645,N_36468);
or U38201 (N_38201,N_36514,N_37742);
nor U38202 (N_38202,N_36928,N_36510);
nor U38203 (N_38203,N_36624,N_36224);
or U38204 (N_38204,N_37617,N_37263);
or U38205 (N_38205,N_36619,N_36146);
nor U38206 (N_38206,N_36364,N_36784);
nor U38207 (N_38207,N_37304,N_37015);
nand U38208 (N_38208,N_36655,N_36939);
xor U38209 (N_38209,N_37629,N_36726);
nand U38210 (N_38210,N_37491,N_37714);
nor U38211 (N_38211,N_37828,N_37343);
nor U38212 (N_38212,N_37411,N_36198);
nand U38213 (N_38213,N_37074,N_36656);
nand U38214 (N_38214,N_37335,N_37891);
nor U38215 (N_38215,N_37222,N_37492);
nand U38216 (N_38216,N_36184,N_37043);
and U38217 (N_38217,N_36097,N_36866);
xor U38218 (N_38218,N_37753,N_36687);
and U38219 (N_38219,N_37811,N_37105);
or U38220 (N_38220,N_37435,N_36071);
xor U38221 (N_38221,N_36651,N_36738);
nand U38222 (N_38222,N_36541,N_37810);
and U38223 (N_38223,N_37760,N_37063);
nand U38224 (N_38224,N_37341,N_36728);
or U38225 (N_38225,N_36465,N_36486);
or U38226 (N_38226,N_37780,N_36754);
xnor U38227 (N_38227,N_36611,N_36799);
xnor U38228 (N_38228,N_36457,N_37959);
nand U38229 (N_38229,N_36284,N_36464);
nand U38230 (N_38230,N_37013,N_36367);
or U38231 (N_38231,N_36787,N_36272);
xnor U38232 (N_38232,N_36153,N_36667);
and U38233 (N_38233,N_36114,N_37702);
nor U38234 (N_38234,N_36730,N_37886);
and U38235 (N_38235,N_37006,N_37675);
xor U38236 (N_38236,N_37381,N_37995);
and U38237 (N_38237,N_37966,N_36564);
nor U38238 (N_38238,N_36570,N_37122);
or U38239 (N_38239,N_36796,N_37481);
and U38240 (N_38240,N_36236,N_37035);
nand U38241 (N_38241,N_36870,N_36724);
or U38242 (N_38242,N_37661,N_37287);
and U38243 (N_38243,N_36637,N_37057);
or U38244 (N_38244,N_36823,N_37964);
nand U38245 (N_38245,N_37767,N_36462);
nand U38246 (N_38246,N_36539,N_36797);
xnor U38247 (N_38247,N_36732,N_37652);
and U38248 (N_38248,N_37619,N_37850);
nor U38249 (N_38249,N_37929,N_37613);
nand U38250 (N_38250,N_36783,N_37689);
xnor U38251 (N_38251,N_37124,N_37697);
and U38252 (N_38252,N_36824,N_36312);
and U38253 (N_38253,N_36192,N_37560);
nand U38254 (N_38254,N_36142,N_36708);
nor U38255 (N_38255,N_36885,N_37917);
xor U38256 (N_38256,N_37954,N_37437);
xnor U38257 (N_38257,N_36320,N_37663);
and U38258 (N_38258,N_37639,N_37601);
and U38259 (N_38259,N_37851,N_36011);
or U38260 (N_38260,N_37885,N_37970);
or U38261 (N_38261,N_36008,N_36351);
nor U38262 (N_38262,N_37176,N_37522);
and U38263 (N_38263,N_36559,N_36676);
nand U38264 (N_38264,N_37265,N_36378);
nor U38265 (N_38265,N_37081,N_37200);
or U38266 (N_38266,N_36440,N_37739);
nand U38267 (N_38267,N_37101,N_37526);
and U38268 (N_38268,N_36130,N_36183);
xnor U38269 (N_38269,N_36969,N_36471);
xnor U38270 (N_38270,N_37672,N_37577);
or U38271 (N_38271,N_36852,N_37458);
nand U38272 (N_38272,N_36608,N_36477);
and U38273 (N_38273,N_37070,N_37143);
nor U38274 (N_38274,N_37422,N_37817);
and U38275 (N_38275,N_37216,N_36076);
and U38276 (N_38276,N_37993,N_36723);
or U38277 (N_38277,N_36369,N_36265);
nor U38278 (N_38278,N_37695,N_36251);
xor U38279 (N_38279,N_37147,N_37747);
and U38280 (N_38280,N_36640,N_36977);
or U38281 (N_38281,N_36193,N_37220);
nor U38282 (N_38282,N_37907,N_36173);
nand U38283 (N_38283,N_37869,N_37160);
xnor U38284 (N_38284,N_37551,N_36620);
nor U38285 (N_38285,N_36279,N_36501);
nor U38286 (N_38286,N_36442,N_37380);
xor U38287 (N_38287,N_37818,N_37257);
nor U38288 (N_38288,N_37424,N_36123);
or U38289 (N_38289,N_37531,N_36758);
nor U38290 (N_38290,N_36281,N_36100);
nand U38291 (N_38291,N_37034,N_36323);
nand U38292 (N_38292,N_36580,N_36187);
and U38293 (N_38293,N_36595,N_36492);
and U38294 (N_38294,N_37219,N_36409);
nor U38295 (N_38295,N_37104,N_37766);
and U38296 (N_38296,N_36405,N_37359);
xnor U38297 (N_38297,N_37438,N_37791);
nand U38298 (N_38298,N_37020,N_37615);
or U38299 (N_38299,N_36849,N_36028);
nand U38300 (N_38300,N_36003,N_36547);
or U38301 (N_38301,N_37943,N_37102);
xor U38302 (N_38302,N_36565,N_37403);
xnor U38303 (N_38303,N_37838,N_36695);
xor U38304 (N_38304,N_36555,N_36157);
nor U38305 (N_38305,N_36075,N_37839);
and U38306 (N_38306,N_36699,N_36370);
nor U38307 (N_38307,N_36277,N_37211);
or U38308 (N_38308,N_36536,N_37370);
or U38309 (N_38309,N_37685,N_36538);
xor U38310 (N_38310,N_36035,N_36961);
xnor U38311 (N_38311,N_36772,N_37510);
nor U38312 (N_38312,N_36120,N_37916);
and U38313 (N_38313,N_36927,N_37784);
nor U38314 (N_38314,N_36613,N_37881);
xnor U38315 (N_38315,N_36951,N_37884);
nand U38316 (N_38316,N_36871,N_37017);
and U38317 (N_38317,N_37001,N_36435);
and U38318 (N_38318,N_36504,N_36567);
or U38319 (N_38319,N_36404,N_36354);
nand U38320 (N_38320,N_37163,N_37465);
nand U38321 (N_38321,N_37280,N_37198);
xor U38322 (N_38322,N_37094,N_37230);
nand U38323 (N_38323,N_37677,N_37120);
or U38324 (N_38324,N_36805,N_37249);
nand U38325 (N_38325,N_37349,N_36195);
nand U38326 (N_38326,N_36036,N_37065);
nand U38327 (N_38327,N_37372,N_37692);
xor U38328 (N_38328,N_37779,N_37582);
xor U38329 (N_38329,N_37855,N_36489);
nor U38330 (N_38330,N_36562,N_36840);
xnor U38331 (N_38331,N_37350,N_37712);
or U38332 (N_38332,N_36742,N_36050);
xnor U38333 (N_38333,N_36618,N_36213);
or U38334 (N_38334,N_37653,N_36127);
nor U38335 (N_38335,N_36473,N_36779);
xor U38336 (N_38336,N_36643,N_36919);
and U38337 (N_38337,N_37820,N_37173);
nand U38338 (N_38338,N_36095,N_36105);
nand U38339 (N_38339,N_36932,N_36942);
and U38340 (N_38340,N_37521,N_36615);
nor U38341 (N_38341,N_37423,N_37440);
nand U38342 (N_38342,N_37690,N_36098);
or U38343 (N_38343,N_36747,N_36638);
xnor U38344 (N_38344,N_37933,N_37735);
xnor U38345 (N_38345,N_37049,N_36534);
nor U38346 (N_38346,N_36686,N_36214);
nand U38347 (N_38347,N_36889,N_37581);
nand U38348 (N_38348,N_36266,N_37047);
or U38349 (N_38349,N_36837,N_36861);
xor U38350 (N_38350,N_37073,N_36382);
xnor U38351 (N_38351,N_36907,N_36882);
xor U38352 (N_38352,N_36400,N_37292);
nor U38353 (N_38353,N_36280,N_36168);
or U38354 (N_38354,N_37880,N_37667);
and U38355 (N_38355,N_36968,N_37552);
xor U38356 (N_38356,N_37744,N_37461);
nand U38357 (N_38357,N_37575,N_37506);
or U38358 (N_38358,N_37442,N_37900);
nor U38359 (N_38359,N_37758,N_36149);
or U38360 (N_38360,N_37569,N_36978);
and U38361 (N_38361,N_37803,N_37827);
and U38362 (N_38362,N_36617,N_37445);
and U38363 (N_38363,N_37574,N_37202);
nand U38364 (N_38364,N_37399,N_37666);
and U38365 (N_38365,N_36186,N_36630);
and U38366 (N_38366,N_36204,N_37969);
nor U38367 (N_38367,N_36802,N_36734);
or U38368 (N_38368,N_37650,N_37532);
nor U38369 (N_38369,N_37227,N_37181);
and U38370 (N_38370,N_37301,N_36828);
nand U38371 (N_38371,N_36156,N_36101);
nand U38372 (N_38372,N_36135,N_37256);
nor U38373 (N_38373,N_37687,N_36548);
nand U38374 (N_38374,N_37170,N_36893);
nand U38375 (N_38375,N_36839,N_37825);
xor U38376 (N_38376,N_36267,N_37967);
or U38377 (N_38377,N_36339,N_36720);
xor U38378 (N_38378,N_36717,N_36503);
and U38379 (N_38379,N_36689,N_37425);
xor U38380 (N_38380,N_37333,N_37519);
or U38381 (N_38381,N_36234,N_37719);
and U38382 (N_38382,N_36967,N_37490);
xnor U38383 (N_38383,N_36719,N_36523);
nor U38384 (N_38384,N_37565,N_36480);
and U38385 (N_38385,N_36924,N_37028);
xnor U38386 (N_38386,N_37930,N_36452);
xnor U38387 (N_38387,N_37467,N_37400);
and U38388 (N_38388,N_36506,N_36902);
nor U38389 (N_38389,N_36646,N_37138);
nor U38390 (N_38390,N_37172,N_36377);
and U38391 (N_38391,N_36029,N_37530);
xnor U38392 (N_38392,N_36113,N_36253);
nand U38393 (N_38393,N_36739,N_37097);
xor U38394 (N_38394,N_37824,N_37329);
nor U38395 (N_38395,N_36984,N_36383);
nor U38396 (N_38396,N_36680,N_36811);
nand U38397 (N_38397,N_37595,N_36423);
nand U38398 (N_38398,N_36573,N_37939);
xnor U38399 (N_38399,N_36762,N_36933);
and U38400 (N_38400,N_36591,N_36596);
xor U38401 (N_38401,N_36847,N_36850);
nor U38402 (N_38402,N_37642,N_36026);
and U38403 (N_38403,N_36240,N_37934);
nand U38404 (N_38404,N_36636,N_36922);
nand U38405 (N_38405,N_36746,N_36604);
xor U38406 (N_38406,N_36931,N_36066);
nand U38407 (N_38407,N_36883,N_37979);
xnor U38408 (N_38408,N_37570,N_37981);
or U38409 (N_38409,N_37977,N_36019);
nand U38410 (N_38410,N_36679,N_36868);
and U38411 (N_38411,N_37463,N_37809);
xnor U38412 (N_38412,N_36842,N_37514);
or U38413 (N_38413,N_36031,N_36790);
and U38414 (N_38414,N_37516,N_36998);
and U38415 (N_38415,N_37949,N_36444);
and U38416 (N_38416,N_36586,N_37771);
nand U38417 (N_38417,N_36909,N_37628);
nand U38418 (N_38418,N_37245,N_36558);
nor U38419 (N_38419,N_36761,N_36016);
and U38420 (N_38420,N_36494,N_36289);
or U38421 (N_38421,N_37271,N_37756);
nor U38422 (N_38422,N_36302,N_36935);
nor U38423 (N_38423,N_37275,N_37854);
and U38424 (N_38424,N_37641,N_37681);
xnor U38425 (N_38425,N_37029,N_36110);
nor U38426 (N_38426,N_36048,N_37208);
and U38427 (N_38427,N_37014,N_37814);
nand U38428 (N_38428,N_36451,N_37799);
and U38429 (N_38429,N_37738,N_37431);
or U38430 (N_38430,N_37285,N_36359);
nor U38431 (N_38431,N_37145,N_37476);
nand U38432 (N_38432,N_37922,N_37655);
nor U38433 (N_38433,N_36181,N_36987);
or U38434 (N_38434,N_37253,N_37419);
nand U38435 (N_38435,N_36741,N_36322);
and U38436 (N_38436,N_37664,N_37306);
nor U38437 (N_38437,N_37115,N_37450);
or U38438 (N_38438,N_36801,N_36262);
nand U38439 (N_38439,N_36517,N_37347);
and U38440 (N_38440,N_36872,N_36357);
or U38441 (N_38441,N_36318,N_37274);
xor U38442 (N_38442,N_37849,N_36111);
nor U38443 (N_38443,N_36285,N_36254);
xor U38444 (N_38444,N_36491,N_37876);
xor U38445 (N_38445,N_37096,N_36314);
nor U38446 (N_38446,N_36352,N_37705);
nor U38447 (N_38447,N_36396,N_36032);
xnor U38448 (N_38448,N_36690,N_36013);
or U38449 (N_38449,N_37212,N_37489);
nand U38450 (N_38450,N_36693,N_36264);
and U38451 (N_38451,N_36915,N_36335);
nand U38452 (N_38452,N_36841,N_37512);
and U38453 (N_38453,N_36386,N_36488);
nand U38454 (N_38454,N_37025,N_36346);
and U38455 (N_38455,N_37862,N_36037);
xnor U38456 (N_38456,N_36419,N_36943);
nand U38457 (N_38457,N_36041,N_36857);
or U38458 (N_38458,N_37627,N_36858);
xnor U38459 (N_38459,N_36122,N_36007);
xnor U38460 (N_38460,N_37204,N_37798);
xnor U38461 (N_38461,N_37988,N_36677);
nor U38462 (N_38462,N_36107,N_37218);
xor U38463 (N_38463,N_36136,N_36301);
and U38464 (N_38464,N_37857,N_37473);
and U38465 (N_38465,N_36996,N_37633);
and U38466 (N_38466,N_37387,N_36350);
xor U38467 (N_38467,N_37355,N_36671);
nor U38468 (N_38468,N_36806,N_36448);
and U38469 (N_38469,N_37951,N_36258);
xnor U38470 (N_38470,N_36670,N_36668);
and U38471 (N_38471,N_36091,N_37870);
xnor U38472 (N_38472,N_37535,N_37882);
and U38473 (N_38473,N_37788,N_36777);
and U38474 (N_38474,N_36499,N_36873);
nand U38475 (N_38475,N_37761,N_36273);
nor U38476 (N_38476,N_36078,N_37267);
nor U38477 (N_38477,N_37348,N_36397);
nand U38478 (N_38478,N_36899,N_36211);
nand U38479 (N_38479,N_37451,N_36735);
and U38480 (N_38480,N_36197,N_37691);
nor U38481 (N_38481,N_36112,N_37478);
nand U38482 (N_38482,N_37207,N_36901);
nand U38483 (N_38483,N_36202,N_37875);
and U38484 (N_38484,N_37903,N_37717);
nand U38485 (N_38485,N_37201,N_36099);
nor U38486 (N_38486,N_37910,N_37611);
xnor U38487 (N_38487,N_36304,N_37802);
xor U38488 (N_38488,N_37938,N_36563);
xnor U38489 (N_38489,N_36361,N_36654);
nand U38490 (N_38490,N_36210,N_36691);
nor U38491 (N_38491,N_37342,N_36879);
nor U38492 (N_38492,N_37480,N_37371);
or U38493 (N_38493,N_37726,N_36766);
nand U38494 (N_38494,N_37139,N_36393);
nand U38495 (N_38495,N_36906,N_36001);
nor U38496 (N_38496,N_37363,N_36950);
xnor U38497 (N_38497,N_37926,N_37485);
nand U38498 (N_38498,N_36103,N_37390);
xor U38499 (N_38499,N_37209,N_37683);
or U38500 (N_38500,N_37162,N_37867);
or U38501 (N_38501,N_36298,N_37911);
nor U38502 (N_38502,N_37676,N_37783);
xnor U38503 (N_38503,N_37906,N_37398);
xor U38504 (N_38504,N_37357,N_36653);
and U38505 (N_38505,N_36644,N_36845);
and U38506 (N_38506,N_37087,N_37098);
nand U38507 (N_38507,N_37571,N_37904);
nand U38508 (N_38508,N_37474,N_36496);
nor U38509 (N_38509,N_36810,N_36096);
or U38510 (N_38510,N_36711,N_36432);
nand U38511 (N_38511,N_36338,N_36474);
and U38512 (N_38512,N_36326,N_37046);
or U38513 (N_38513,N_37294,N_37523);
and U38514 (N_38514,N_36633,N_36912);
nand U38515 (N_38515,N_37750,N_36827);
nand U38516 (N_38516,N_37010,N_36751);
nor U38517 (N_38517,N_36333,N_37007);
nor U38518 (N_38518,N_37498,N_36880);
nor U38519 (N_38519,N_37562,N_36180);
nand U38520 (N_38520,N_37863,N_37898);
nand U38521 (N_38521,N_37684,N_36660);
or U38522 (N_38522,N_36891,N_36245);
and U38523 (N_38523,N_36561,N_36217);
and U38524 (N_38524,N_37500,N_37157);
or U38525 (N_38525,N_36344,N_37859);
or U38526 (N_38526,N_36914,N_36736);
nand U38527 (N_38527,N_36863,N_36976);
nor U38528 (N_38528,N_36674,N_37239);
or U38529 (N_38529,N_37068,N_36399);
and U38530 (N_38530,N_36476,N_37763);
or U38531 (N_38531,N_37189,N_36664);
xor U38532 (N_38532,N_37923,N_36685);
nand U38533 (N_38533,N_37213,N_37950);
nor U38534 (N_38534,N_37117,N_36436);
nor U38535 (N_38535,N_36771,N_36662);
and U38536 (N_38536,N_37853,N_36447);
xor U38537 (N_38537,N_36578,N_37314);
or U38538 (N_38538,N_36137,N_36648);
xnor U38539 (N_38539,N_37625,N_36502);
xnor U38540 (N_38540,N_37515,N_37895);
nand U38541 (N_38541,N_36647,N_37541);
nand U38542 (N_38542,N_36634,N_37698);
or U38543 (N_38543,N_37030,N_37846);
nand U38544 (N_38544,N_36508,N_37554);
nor U38545 (N_38545,N_37251,N_37027);
or U38546 (N_38546,N_36763,N_36102);
and U38547 (N_38547,N_36282,N_37210);
nor U38548 (N_38548,N_37928,N_37608);
xnor U38549 (N_38549,N_37297,N_37472);
and U38550 (N_38550,N_36022,N_36625);
or U38551 (N_38551,N_37464,N_36238);
xnor U38552 (N_38552,N_37553,N_37723);
or U38553 (N_38553,N_36701,N_37920);
or U38554 (N_38554,N_36068,N_36853);
nand U38555 (N_38555,N_36119,N_37214);
or U38556 (N_38556,N_37344,N_36353);
and U38557 (N_38557,N_37734,N_37311);
nor U38558 (N_38558,N_36781,N_37674);
and U38559 (N_38559,N_36445,N_36310);
and U38560 (N_38560,N_36345,N_37538);
xnor U38561 (N_38561,N_36166,N_37353);
nor U38562 (N_38562,N_37273,N_37169);
and U38563 (N_38563,N_37657,N_37946);
or U38564 (N_38564,N_36014,N_36315);
nor U38565 (N_38565,N_36461,N_36073);
and U38566 (N_38566,N_37050,N_36039);
nor U38567 (N_38567,N_36513,N_36791);
or U38568 (N_38568,N_37759,N_36974);
or U38569 (N_38569,N_36949,N_37752);
or U38570 (N_38570,N_37185,N_36778);
nand U38571 (N_38571,N_36599,N_37529);
nand U38572 (N_38572,N_37801,N_37826);
xnor U38573 (N_38573,N_36516,N_37737);
xor U38574 (N_38574,N_37153,N_37455);
nand U38575 (N_38575,N_37765,N_36807);
or U38576 (N_38576,N_36063,N_37847);
nor U38577 (N_38577,N_36694,N_36085);
xor U38578 (N_38578,N_36550,N_36544);
xnor U38579 (N_38579,N_36809,N_36033);
nor U38580 (N_38580,N_37444,N_37036);
nand U38581 (N_38581,N_37291,N_37785);
xnor U38582 (N_38582,N_37337,N_37316);
and U38583 (N_38583,N_36765,N_36574);
nand U38584 (N_38584,N_36556,N_36244);
xor U38585 (N_38585,N_37796,N_36190);
nor U38586 (N_38586,N_37376,N_37103);
or U38587 (N_38587,N_37142,N_37319);
and U38588 (N_38588,N_37430,N_36579);
or U38589 (N_38589,N_36515,N_37487);
and U38590 (N_38590,N_36221,N_36389);
nand U38591 (N_38591,N_36487,N_37985);
or U38592 (N_38592,N_37660,N_37806);
xnor U38593 (N_38593,N_36268,N_37696);
nand U38594 (N_38594,N_37736,N_36051);
or U38595 (N_38595,N_36161,N_37460);
and U38596 (N_38596,N_36255,N_37225);
nor U38597 (N_38597,N_36274,N_37223);
nand U38598 (N_38598,N_36588,N_36356);
xnor U38599 (N_38599,N_36372,N_37447);
or U38600 (N_38600,N_37589,N_37718);
nand U38601 (N_38601,N_36908,N_37864);
xnor U38602 (N_38602,N_36201,N_36937);
xor U38603 (N_38603,N_36049,N_37721);
and U38604 (N_38604,N_36817,N_36948);
nor U38605 (N_38605,N_37534,N_37008);
or U38606 (N_38606,N_36585,N_36553);
nand U38607 (N_38607,N_36519,N_36467);
or U38608 (N_38608,N_37962,N_37366);
or U38609 (N_38609,N_36424,N_36043);
xor U38610 (N_38610,N_37392,N_37497);
xnor U38611 (N_38611,N_37704,N_36792);
nor U38612 (N_38612,N_37078,N_37079);
and U38613 (N_38613,N_37963,N_36118);
nand U38614 (N_38614,N_37991,N_36601);
nand U38615 (N_38615,N_36542,N_36941);
nand U38616 (N_38616,N_36583,N_36775);
and U38617 (N_38617,N_37242,N_37228);
and U38618 (N_38618,N_36252,N_37136);
xor U38619 (N_38619,N_37093,N_37024);
nor U38620 (N_38620,N_36300,N_37259);
or U38621 (N_38621,N_36176,N_36207);
nand U38622 (N_38622,N_37012,N_37848);
nand U38623 (N_38623,N_37151,N_36537);
nor U38624 (N_38624,N_36203,N_37427);
or U38625 (N_38625,N_37769,N_36566);
xnor U38626 (N_38626,N_37429,N_36472);
or U38627 (N_38627,N_36554,N_36470);
nor U38628 (N_38628,N_36228,N_36944);
or U38629 (N_38629,N_36276,N_37258);
xor U38630 (N_38630,N_36825,N_36709);
or U38631 (N_38631,N_36431,N_36590);
xnor U38632 (N_38632,N_36449,N_37724);
and U38633 (N_38633,N_37042,N_37039);
xor U38634 (N_38634,N_37812,N_37483);
xor U38635 (N_38635,N_36232,N_36316);
and U38636 (N_38636,N_36422,N_37730);
xor U38637 (N_38637,N_37665,N_37260);
nor U38638 (N_38638,N_36169,N_37134);
and U38639 (N_38639,N_37388,N_37362);
nand U38640 (N_38640,N_37443,N_37334);
and U38641 (N_38641,N_36368,N_36639);
and U38642 (N_38642,N_37237,N_36283);
nor U38643 (N_38643,N_36343,N_36177);
xor U38644 (N_38644,N_36237,N_36360);
nor U38645 (N_38645,N_36083,N_36004);
nand U38646 (N_38646,N_36179,N_37533);
nor U38647 (N_38647,N_36434,N_36986);
nand U38648 (N_38648,N_37109,N_37315);
and U38649 (N_38649,N_37693,N_37952);
or U38650 (N_38650,N_36665,N_37459);
nand U38651 (N_38651,N_36507,N_37794);
and U38652 (N_38652,N_36147,N_36527);
nand U38653 (N_38653,N_36862,N_36930);
and U38654 (N_38654,N_37127,N_36992);
and U38655 (N_38655,N_36151,N_37748);
and U38656 (N_38656,N_37302,N_37468);
nor U38657 (N_38657,N_36822,N_37555);
and U38658 (N_38658,N_36006,N_36220);
or U38659 (N_38659,N_36980,N_36911);
nand U38660 (N_38660,N_37563,N_37971);
nand U38661 (N_38661,N_36860,N_36712);
nor U38662 (N_38662,N_37453,N_36030);
or U38663 (N_38663,N_37790,N_37899);
or U38664 (N_38664,N_36395,N_37022);
nand U38665 (N_38665,N_36175,N_36331);
xnor U38666 (N_38666,N_36622,N_37990);
and U38667 (N_38667,N_37221,N_37493);
xor U38668 (N_38668,N_37140,N_37961);
and U38669 (N_38669,N_37965,N_37776);
nor U38670 (N_38670,N_36962,N_36521);
or U38671 (N_38671,N_37418,N_36385);
nor U38672 (N_38672,N_37003,N_37135);
and U38673 (N_38673,N_37309,N_36250);
and U38674 (N_38674,N_36785,N_36158);
and U38675 (N_38675,N_37494,N_36626);
or U38676 (N_38676,N_36576,N_37586);
and U38677 (N_38677,N_36133,N_36426);
nand U38678 (N_38678,N_36531,N_36940);
or U38679 (N_38679,N_36756,N_36216);
nand U38680 (N_38680,N_37307,N_37976);
xor U38681 (N_38681,N_36421,N_37137);
and U38682 (N_38682,N_37549,N_36737);
or U38683 (N_38683,N_37312,N_36313);
and U38684 (N_38684,N_36904,N_37454);
xnor U38685 (N_38685,N_37984,N_37770);
and U38686 (N_38686,N_37300,N_37420);
nand U38687 (N_38687,N_37874,N_37410);
nand U38688 (N_38688,N_37352,N_37125);
xor U38689 (N_38689,N_37299,N_36964);
or U38690 (N_38690,N_37339,N_36257);
or U38691 (N_38691,N_37084,N_37417);
nor U38692 (N_38692,N_36340,N_37130);
or U38693 (N_38693,N_36411,N_37317);
nand U38694 (N_38694,N_37609,N_37805);
and U38695 (N_38695,N_36408,N_36753);
xnor U38696 (N_38696,N_36602,N_36609);
nor U38697 (N_38697,N_36979,N_37486);
nor U38698 (N_38698,N_37578,N_36820);
nor U38699 (N_38699,N_36975,N_37835);
nand U38700 (N_38700,N_36053,N_37112);
nor U38701 (N_38701,N_37331,N_37195);
xnor U38702 (N_38702,N_36748,N_37757);
nand U38703 (N_38703,N_36241,N_37887);
nand U38704 (N_38704,N_36108,N_36878);
nand U38705 (N_38705,N_36410,N_36012);
nand U38706 (N_38706,N_37113,N_36981);
nor U38707 (N_38707,N_36141,N_36816);
and U38708 (N_38708,N_36903,N_37764);
xor U38709 (N_38709,N_37205,N_36094);
nand U38710 (N_38710,N_37255,N_36881);
or U38711 (N_38711,N_36191,N_37700);
xnor U38712 (N_38712,N_36199,N_36089);
and U38713 (N_38713,N_36757,N_36278);
nor U38714 (N_38714,N_36309,N_36900);
nand U38715 (N_38715,N_37973,N_36307);
nand U38716 (N_38716,N_37786,N_37354);
xor U38717 (N_38717,N_37720,N_36249);
nand U38718 (N_38718,N_37031,N_37821);
and U38719 (N_38719,N_36291,N_37901);
or U38720 (N_38720,N_37942,N_36938);
or U38721 (N_38721,N_37433,N_36381);
nand U38722 (N_38722,N_37374,N_37144);
nor U38723 (N_38723,N_36463,N_36560);
nor U38724 (N_38724,N_37193,N_36838);
xnor U38725 (N_38725,N_36055,N_37174);
nand U38726 (N_38726,N_36116,N_37539);
and U38727 (N_38727,N_36641,N_36605);
and U38728 (N_38728,N_37610,N_36024);
or U38729 (N_38729,N_36577,N_36549);
nor U38730 (N_38730,N_37927,N_37706);
xor U38731 (N_38731,N_36684,N_36991);
xor U38732 (N_38732,N_37754,N_36836);
nand U38733 (N_38733,N_37914,N_36227);
or U38734 (N_38734,N_36973,N_37822);
or U38735 (N_38735,N_37203,N_37470);
xor U38736 (N_38736,N_36493,N_36243);
or U38737 (N_38737,N_36079,N_37026);
or U38738 (N_38738,N_37647,N_36086);
or U38739 (N_38739,N_37000,N_37155);
nor U38740 (N_38740,N_37517,N_37682);
nor U38741 (N_38741,N_36000,N_37893);
and U38742 (N_38742,N_37732,N_36826);
and U38743 (N_38743,N_37631,N_36021);
and U38744 (N_38744,N_37932,N_37002);
nor U38745 (N_38745,N_36040,N_36509);
nor U38746 (N_38746,N_37877,N_36072);
nand U38747 (N_38747,N_36438,N_37183);
xor U38748 (N_38748,N_37507,N_37604);
and U38749 (N_38749,N_37804,N_37558);
nor U38750 (N_38750,N_36349,N_36375);
nor U38751 (N_38751,N_37360,N_36481);
or U38752 (N_38752,N_36325,N_36047);
nand U38753 (N_38753,N_37086,N_37585);
or U38754 (N_38754,N_36650,N_37167);
nand U38755 (N_38755,N_37841,N_36760);
and U38756 (N_38756,N_37777,N_36731);
nor U38757 (N_38757,N_36848,N_37679);
nand U38758 (N_38758,N_36997,N_37471);
or U38759 (N_38759,N_36165,N_36446);
xnor U38760 (N_38760,N_37596,N_36200);
and U38761 (N_38761,N_36970,N_37058);
or U38762 (N_38762,N_36296,N_37108);
nor U38763 (N_38763,N_37892,N_36275);
nand U38764 (N_38764,N_37662,N_36392);
or U38765 (N_38765,N_36855,N_37336);
or U38766 (N_38766,N_37637,N_36788);
xnor U38767 (N_38767,N_37106,N_36495);
nand U38768 (N_38768,N_37612,N_36341);
and U38769 (N_38769,N_37452,N_37272);
and U38770 (N_38770,N_36954,N_36416);
nand U38771 (N_38771,N_37367,N_37668);
nor U38772 (N_38772,N_36178,N_36067);
xor U38773 (N_38773,N_36854,N_36856);
or U38774 (N_38774,N_36390,N_37778);
or U38775 (N_38775,N_36263,N_37293);
nor U38776 (N_38776,N_36946,N_37262);
nand U38777 (N_38777,N_37546,N_37997);
or U38778 (N_38778,N_37241,N_37041);
nor U38779 (N_38779,N_36150,N_36773);
or U38780 (N_38780,N_37233,N_37479);
nand U38781 (N_38781,N_36713,N_37649);
nand U38782 (N_38782,N_37987,N_37671);
or U38783 (N_38783,N_37936,N_36971);
and U38784 (N_38784,N_37513,N_37100);
nor U38785 (N_38785,N_36230,N_37602);
or U38786 (N_38786,N_36896,N_37599);
nand U38787 (N_38787,N_37441,N_37052);
or U38788 (N_38788,N_37270,N_37397);
or U38789 (N_38789,N_37072,N_36174);
xnor U38790 (N_38790,N_36597,N_37091);
or U38791 (N_38791,N_37626,N_37908);
or U38792 (N_38792,N_37375,N_36594);
xor U38793 (N_38793,N_37475,N_36780);
and U38794 (N_38794,N_37248,N_37566);
nand U38795 (N_38795,N_37947,N_37018);
xor U38796 (N_38796,N_36518,N_36131);
xnor U38797 (N_38797,N_37746,N_37871);
nand U38798 (N_38798,N_36642,N_36552);
xnor U38799 (N_38799,N_37011,N_37725);
or U38800 (N_38800,N_37852,N_37190);
xnor U38801 (N_38801,N_37673,N_37150);
xnor U38802 (N_38802,N_37278,N_36669);
xnor U38803 (N_38803,N_37385,N_37948);
xnor U38804 (N_38804,N_36835,N_36260);
and U38805 (N_38805,N_36129,N_37643);
nand U38806 (N_38806,N_36215,N_37795);
nor U38807 (N_38807,N_37635,N_36433);
nand U38808 (N_38808,N_37192,N_37277);
nor U38809 (N_38809,N_37111,N_37518);
xor U38810 (N_38810,N_36793,N_37434);
and U38811 (N_38811,N_36417,N_36334);
or U38812 (N_38812,N_36132,N_37731);
nor U38813 (N_38813,N_36533,N_37762);
and U38814 (N_38814,N_36246,N_37323);
nor U38815 (N_38815,N_37175,N_36524);
and U38816 (N_38816,N_36387,N_37879);
nor U38817 (N_38817,N_36988,N_37741);
or U38818 (N_38818,N_37009,N_36270);
nand U38819 (N_38819,N_36934,N_37062);
nand U38820 (N_38820,N_37620,N_36106);
or U38821 (N_38821,N_37340,N_37126);
or U38822 (N_38822,N_36401,N_37590);
and U38823 (N_38823,N_37244,N_37282);
xor U38824 (N_38824,N_37123,N_36225);
xor U38825 (N_38825,N_36635,N_36672);
nor U38826 (N_38826,N_37935,N_36729);
nor U38827 (N_38827,N_36715,N_37114);
nor U38828 (N_38828,N_36458,N_36311);
nand U38829 (N_38829,N_36321,N_37303);
xor U38830 (N_38830,N_37236,N_37229);
nor U38831 (N_38831,N_37132,N_37179);
xor U38832 (N_38832,N_37699,N_36015);
xnor U38833 (N_38833,N_37989,N_37338);
nor U38834 (N_38834,N_36698,N_37833);
and U38835 (N_38835,N_37708,N_37941);
nand U38836 (N_38836,N_36406,N_36218);
xnor U38837 (N_38837,N_37196,N_36782);
xor U38838 (N_38838,N_37924,N_37957);
nor U38839 (N_38839,N_37436,N_37545);
nand U38840 (N_38840,N_37495,N_36678);
xnor U38841 (N_38841,N_37587,N_37992);
nand U38842 (N_38842,N_37972,N_36308);
nand U38843 (N_38843,N_36497,N_37556);
nand U38844 (N_38844,N_36046,N_36305);
or U38845 (N_38845,N_37624,N_37178);
xnor U38846 (N_38846,N_36832,N_37502);
nand U38847 (N_38847,N_36242,N_37606);
or U38848 (N_38848,N_36804,N_36929);
nor U38849 (N_38849,N_36017,N_37154);
nand U38850 (N_38850,N_36490,N_37630);
or U38851 (N_38851,N_36505,N_37944);
nor U38852 (N_38852,N_36128,N_37813);
and U38853 (N_38853,N_36159,N_37686);
nand U38854 (N_38854,N_37439,N_37149);
nand U38855 (N_38855,N_36059,N_36952);
nor U38856 (N_38856,N_36727,N_37501);
nor U38857 (N_38857,N_36623,N_36170);
nand U38858 (N_38858,N_37286,N_37945);
nor U38859 (N_38859,N_37184,N_37308);
xor U38860 (N_38860,N_36139,N_36956);
nand U38861 (N_38861,N_37206,N_37088);
or U38862 (N_38862,N_37709,N_36407);
nor U38863 (N_38863,N_37351,N_37740);
and U38864 (N_38864,N_37819,N_36569);
and U38865 (N_38865,N_36829,N_36892);
or U38866 (N_38866,N_36666,N_36342);
nor U38867 (N_38867,N_37815,N_37197);
xor U38868 (N_38868,N_36025,N_37583);
nand U38869 (N_38869,N_37844,N_36688);
or U38870 (N_38870,N_37456,N_36815);
and U38871 (N_38871,N_36658,N_36164);
xor U38872 (N_38872,N_36936,N_36443);
nor U38873 (N_38873,N_36581,N_36010);
xor U38874 (N_38874,N_36362,N_36571);
nand U38875 (N_38875,N_37651,N_36231);
nand U38876 (N_38876,N_37379,N_36675);
xor U38877 (N_38877,N_36990,N_37999);
and U38878 (N_38878,N_37499,N_37182);
or U38879 (N_38879,N_37940,N_36612);
xnor U38880 (N_38880,N_36725,N_36479);
xor U38881 (N_38881,N_37703,N_36923);
xnor U38882 (N_38882,N_36786,N_37394);
nor U38883 (N_38883,N_36484,N_37636);
or U38884 (N_38884,N_37378,N_37032);
nor U38885 (N_38885,N_37056,N_37496);
or U38886 (N_38886,N_37547,N_36918);
or U38887 (N_38887,N_36057,N_36921);
xor U38888 (N_38888,N_37716,N_37288);
xor U38889 (N_38889,N_37865,N_37076);
or U38890 (N_38890,N_36140,N_36034);
xor U38891 (N_38891,N_37268,N_37542);
nand U38892 (N_38892,N_37129,N_36188);
nor U38893 (N_38893,N_36592,N_36171);
or U38894 (N_38894,N_37537,N_36628);
or U38895 (N_38895,N_36212,N_37774);
nor U38896 (N_38896,N_37021,N_37829);
nand U38897 (N_38897,N_36045,N_36475);
or U38898 (N_38898,N_36172,N_36038);
and U38899 (N_38899,N_36945,N_36469);
and U38900 (N_38900,N_37890,N_36657);
nand U38901 (N_38901,N_37773,N_37902);
nand U38902 (N_38902,N_37918,N_36610);
xor U38903 (N_38903,N_36768,N_37177);
and U38904 (N_38904,N_37281,N_37540);
and U38905 (N_38905,N_36511,N_36800);
or U38906 (N_38906,N_36812,N_36764);
or U38907 (N_38907,N_36205,N_37974);
xnor U38908 (N_38908,N_36683,N_37080);
or U38909 (N_38909,N_36886,N_36994);
and U38910 (N_38910,N_36058,N_37937);
nand U38911 (N_38911,N_37384,N_37133);
or U38912 (N_38912,N_36425,N_37527);
and U38913 (N_38913,N_37243,N_37960);
xnor U38914 (N_38914,N_36121,N_36163);
nor U38915 (N_38915,N_36299,N_37618);
nand U38916 (N_38916,N_37235,N_36223);
and U38917 (N_38917,N_36520,N_37290);
xnor U38918 (N_38918,N_36876,N_37745);
xor U38919 (N_38919,N_37787,N_37789);
and U38920 (N_38920,N_37477,N_36794);
and U38921 (N_38921,N_37508,N_36074);
nor U38922 (N_38922,N_36716,N_36336);
and U38923 (N_38923,N_36865,N_36890);
and U38924 (N_38924,N_37165,N_37634);
and U38925 (N_38925,N_36104,N_36535);
xor U38926 (N_38926,N_36607,N_36913);
nand U38927 (N_38927,N_36500,N_36551);
nor U38928 (N_38928,N_36081,N_37364);
or U38929 (N_38929,N_37823,N_36813);
xnor U38930 (N_38930,N_37402,N_36235);
and U38931 (N_38931,N_37266,N_36512);
nor U38932 (N_38932,N_36347,N_37121);
xnor U38933 (N_38933,N_36589,N_36398);
xnor U38934 (N_38934,N_37837,N_36327);
nand U38935 (N_38935,N_36575,N_37567);
xnor U38936 (N_38936,N_36982,N_37382);
nor U38937 (N_38937,N_37509,N_37488);
nor U38938 (N_38938,N_37324,N_36388);
or U38939 (N_38939,N_37289,N_37834);
nand U38940 (N_38940,N_36295,N_36332);
or U38941 (N_38941,N_37188,N_36229);
or U38942 (N_38942,N_36917,N_37701);
nor U38943 (N_38943,N_36614,N_36064);
or U38944 (N_38944,N_37090,N_37638);
xnor U38945 (N_38945,N_37872,N_37405);
and U38946 (N_38946,N_37845,N_36898);
xnor U38947 (N_38947,N_37894,N_37953);
nor U38948 (N_38948,N_37772,N_37743);
xor U38949 (N_38949,N_37607,N_36337);
xnor U38950 (N_38950,N_36659,N_37873);
nand U38951 (N_38951,N_36920,N_37616);
or U38952 (N_38952,N_36957,N_37045);
xnor U38953 (N_38953,N_37504,N_37905);
nor U38954 (N_38954,N_37994,N_36330);
nand U38955 (N_38955,N_37005,N_37199);
nand U38956 (N_38956,N_36060,N_36833);
nand U38957 (N_38957,N_37060,N_37119);
or U38958 (N_38958,N_37986,N_37727);
nand U38959 (N_38959,N_36061,N_37592);
nand U38960 (N_38960,N_37432,N_37680);
and U38961 (N_38961,N_36703,N_37396);
nor U38962 (N_38962,N_37830,N_37095);
xor U38963 (N_38963,N_36959,N_37858);
and U38964 (N_38964,N_36584,N_36587);
xor U38965 (N_38965,N_37099,N_37016);
xor U38966 (N_38966,N_37751,N_37710);
xor U38967 (N_38967,N_37921,N_36269);
nor U38968 (N_38968,N_37116,N_36483);
xnor U38969 (N_38969,N_36065,N_37883);
nor U38970 (N_38970,N_37247,N_36402);
nand U38971 (N_38971,N_36441,N_37524);
and U38972 (N_38972,N_36222,N_36750);
nor U38973 (N_38973,N_37059,N_37816);
nor U38974 (N_38974,N_37648,N_36294);
nor U38975 (N_38975,N_37931,N_37358);
and U38976 (N_38976,N_37295,N_36117);
nor U38977 (N_38977,N_37919,N_36629);
nor U38978 (N_38978,N_37004,N_36645);
or U38979 (N_38979,N_36115,N_36070);
and U38980 (N_38980,N_36874,N_37955);
or U38981 (N_38981,N_36018,N_37252);
xor U38982 (N_38982,N_36632,N_36705);
and U38983 (N_38983,N_37511,N_36226);
nor U38984 (N_38984,N_36532,N_36710);
nand U38985 (N_38985,N_37159,N_37406);
xor U38986 (N_38986,N_36134,N_36568);
or U38987 (N_38987,N_37775,N_36925);
or U38988 (N_38988,N_37842,N_36259);
and U38989 (N_38989,N_36482,N_36910);
nand U38990 (N_38990,N_37276,N_36456);
and U38991 (N_38991,N_36196,N_37254);
or U38992 (N_38992,N_36373,N_37909);
nand U38993 (N_38993,N_36905,N_36287);
and U38994 (N_38994,N_37401,N_37856);
or U38995 (N_38995,N_36466,N_36329);
nor U38996 (N_38996,N_36593,N_36598);
nor U38997 (N_38997,N_37588,N_36219);
and U38998 (N_38998,N_36803,N_36427);
and U38999 (N_38999,N_37915,N_36371);
and U39000 (N_39000,N_36008,N_37741);
nor U39001 (N_39001,N_37924,N_36360);
xor U39002 (N_39002,N_37058,N_37748);
or U39003 (N_39003,N_36776,N_37019);
nor U39004 (N_39004,N_37922,N_36128);
or U39005 (N_39005,N_36520,N_36613);
xnor U39006 (N_39006,N_36216,N_36424);
or U39007 (N_39007,N_37313,N_37500);
xnor U39008 (N_39008,N_37488,N_36779);
xnor U39009 (N_39009,N_36170,N_37925);
or U39010 (N_39010,N_36761,N_36575);
nor U39011 (N_39011,N_37727,N_37107);
nand U39012 (N_39012,N_36057,N_36502);
nor U39013 (N_39013,N_37566,N_37845);
xnor U39014 (N_39014,N_36755,N_37050);
xnor U39015 (N_39015,N_37043,N_37694);
nand U39016 (N_39016,N_37329,N_36278);
nand U39017 (N_39017,N_36524,N_36674);
nand U39018 (N_39018,N_37598,N_37369);
nor U39019 (N_39019,N_37944,N_36192);
or U39020 (N_39020,N_37428,N_36924);
nor U39021 (N_39021,N_37988,N_36679);
xor U39022 (N_39022,N_37441,N_36574);
and U39023 (N_39023,N_36876,N_36613);
nand U39024 (N_39024,N_36545,N_37374);
nor U39025 (N_39025,N_36332,N_37756);
or U39026 (N_39026,N_37136,N_37446);
and U39027 (N_39027,N_36129,N_37480);
nand U39028 (N_39028,N_36189,N_36357);
nor U39029 (N_39029,N_37407,N_37914);
and U39030 (N_39030,N_36567,N_36353);
nand U39031 (N_39031,N_37302,N_36813);
nor U39032 (N_39032,N_37526,N_37642);
and U39033 (N_39033,N_36333,N_37549);
nand U39034 (N_39034,N_37430,N_36594);
xnor U39035 (N_39035,N_37728,N_36321);
nor U39036 (N_39036,N_37536,N_37774);
xor U39037 (N_39037,N_37443,N_36219);
xnor U39038 (N_39038,N_36885,N_37739);
nand U39039 (N_39039,N_37763,N_36642);
and U39040 (N_39040,N_37081,N_37447);
and U39041 (N_39041,N_37397,N_36043);
nor U39042 (N_39042,N_37850,N_36974);
nor U39043 (N_39043,N_37934,N_37057);
and U39044 (N_39044,N_36106,N_36972);
nand U39045 (N_39045,N_36654,N_36970);
and U39046 (N_39046,N_37082,N_36035);
xnor U39047 (N_39047,N_36724,N_37586);
xnor U39048 (N_39048,N_36666,N_36052);
xor U39049 (N_39049,N_36716,N_36902);
xor U39050 (N_39050,N_37392,N_37016);
nand U39051 (N_39051,N_36384,N_37012);
and U39052 (N_39052,N_36671,N_37699);
or U39053 (N_39053,N_37390,N_36356);
nor U39054 (N_39054,N_37466,N_37444);
nand U39055 (N_39055,N_37733,N_36394);
and U39056 (N_39056,N_37466,N_36270);
and U39057 (N_39057,N_37029,N_36608);
nor U39058 (N_39058,N_37100,N_36263);
xnor U39059 (N_39059,N_37265,N_37314);
or U39060 (N_39060,N_37730,N_36147);
xor U39061 (N_39061,N_36484,N_36715);
xor U39062 (N_39062,N_37349,N_37288);
nand U39063 (N_39063,N_36275,N_37319);
nand U39064 (N_39064,N_36540,N_37553);
nand U39065 (N_39065,N_37897,N_36290);
nor U39066 (N_39066,N_36705,N_36802);
or U39067 (N_39067,N_37242,N_37739);
nor U39068 (N_39068,N_36304,N_37604);
xnor U39069 (N_39069,N_37216,N_37632);
and U39070 (N_39070,N_36724,N_36365);
nor U39071 (N_39071,N_37778,N_37308);
nor U39072 (N_39072,N_37190,N_36045);
and U39073 (N_39073,N_37704,N_37097);
nand U39074 (N_39074,N_36593,N_36328);
nand U39075 (N_39075,N_37326,N_36986);
or U39076 (N_39076,N_36251,N_37623);
or U39077 (N_39077,N_36831,N_36918);
nor U39078 (N_39078,N_37467,N_36537);
and U39079 (N_39079,N_37004,N_36351);
nor U39080 (N_39080,N_37097,N_37241);
and U39081 (N_39081,N_37764,N_36636);
xnor U39082 (N_39082,N_36759,N_36417);
or U39083 (N_39083,N_36564,N_37291);
or U39084 (N_39084,N_36295,N_36635);
or U39085 (N_39085,N_36510,N_36595);
and U39086 (N_39086,N_37455,N_36950);
nand U39087 (N_39087,N_36844,N_37881);
or U39088 (N_39088,N_36604,N_36322);
and U39089 (N_39089,N_37708,N_37308);
nand U39090 (N_39090,N_36463,N_36229);
nand U39091 (N_39091,N_37323,N_36135);
or U39092 (N_39092,N_36037,N_36175);
and U39093 (N_39093,N_36184,N_36146);
xnor U39094 (N_39094,N_36722,N_37160);
nand U39095 (N_39095,N_37302,N_36545);
or U39096 (N_39096,N_36490,N_37637);
or U39097 (N_39097,N_36468,N_36623);
or U39098 (N_39098,N_36272,N_36155);
xor U39099 (N_39099,N_37921,N_37920);
and U39100 (N_39100,N_37195,N_37024);
and U39101 (N_39101,N_36749,N_37680);
nand U39102 (N_39102,N_36609,N_36608);
nor U39103 (N_39103,N_37855,N_37903);
nand U39104 (N_39104,N_36796,N_36905);
nand U39105 (N_39105,N_36578,N_36652);
or U39106 (N_39106,N_36428,N_36615);
or U39107 (N_39107,N_37222,N_36660);
or U39108 (N_39108,N_36271,N_36013);
nor U39109 (N_39109,N_36018,N_36638);
and U39110 (N_39110,N_37809,N_36922);
nor U39111 (N_39111,N_37986,N_37427);
nor U39112 (N_39112,N_37531,N_37005);
or U39113 (N_39113,N_36544,N_37717);
nor U39114 (N_39114,N_37278,N_36598);
and U39115 (N_39115,N_36150,N_36451);
or U39116 (N_39116,N_37268,N_37460);
nand U39117 (N_39117,N_36427,N_36614);
xor U39118 (N_39118,N_37109,N_37025);
nor U39119 (N_39119,N_37437,N_37110);
nand U39120 (N_39120,N_36911,N_36931);
xnor U39121 (N_39121,N_36671,N_36792);
or U39122 (N_39122,N_36417,N_36744);
xnor U39123 (N_39123,N_37255,N_37917);
or U39124 (N_39124,N_37846,N_37633);
or U39125 (N_39125,N_37569,N_37900);
nand U39126 (N_39126,N_36804,N_36615);
or U39127 (N_39127,N_36402,N_36000);
xor U39128 (N_39128,N_37434,N_37918);
and U39129 (N_39129,N_36658,N_37780);
or U39130 (N_39130,N_36249,N_36373);
xnor U39131 (N_39131,N_37973,N_37915);
or U39132 (N_39132,N_36014,N_37484);
nand U39133 (N_39133,N_36578,N_36935);
and U39134 (N_39134,N_37892,N_37146);
or U39135 (N_39135,N_37823,N_37392);
and U39136 (N_39136,N_37089,N_37800);
and U39137 (N_39137,N_36868,N_37181);
xnor U39138 (N_39138,N_37124,N_37392);
or U39139 (N_39139,N_37654,N_36316);
nor U39140 (N_39140,N_37975,N_36647);
or U39141 (N_39141,N_36070,N_36409);
or U39142 (N_39142,N_36483,N_37013);
nand U39143 (N_39143,N_37504,N_36706);
nor U39144 (N_39144,N_36549,N_36773);
nand U39145 (N_39145,N_37573,N_36356);
nand U39146 (N_39146,N_36348,N_36086);
and U39147 (N_39147,N_36324,N_37130);
nor U39148 (N_39148,N_36283,N_36858);
or U39149 (N_39149,N_37861,N_37678);
nor U39150 (N_39150,N_36531,N_37513);
and U39151 (N_39151,N_37111,N_37009);
xor U39152 (N_39152,N_36396,N_36139);
nor U39153 (N_39153,N_37602,N_37853);
and U39154 (N_39154,N_37075,N_37949);
or U39155 (N_39155,N_37674,N_36947);
nand U39156 (N_39156,N_36656,N_37510);
or U39157 (N_39157,N_36437,N_37380);
and U39158 (N_39158,N_36019,N_37208);
nor U39159 (N_39159,N_37575,N_36530);
nand U39160 (N_39160,N_36132,N_37822);
nor U39161 (N_39161,N_36841,N_36582);
nor U39162 (N_39162,N_37836,N_36183);
xor U39163 (N_39163,N_36541,N_36287);
xnor U39164 (N_39164,N_37112,N_36188);
nor U39165 (N_39165,N_36710,N_36231);
nor U39166 (N_39166,N_37840,N_37522);
or U39167 (N_39167,N_37666,N_36264);
nor U39168 (N_39168,N_37530,N_37470);
nand U39169 (N_39169,N_37136,N_36217);
or U39170 (N_39170,N_37014,N_36026);
nor U39171 (N_39171,N_37622,N_37646);
xor U39172 (N_39172,N_37603,N_37952);
or U39173 (N_39173,N_36167,N_37490);
nor U39174 (N_39174,N_36619,N_37128);
or U39175 (N_39175,N_36906,N_36131);
nor U39176 (N_39176,N_37891,N_36089);
and U39177 (N_39177,N_37660,N_36653);
and U39178 (N_39178,N_37924,N_37683);
nor U39179 (N_39179,N_37530,N_36920);
nand U39180 (N_39180,N_36606,N_37428);
or U39181 (N_39181,N_37089,N_37203);
nand U39182 (N_39182,N_36595,N_37258);
nand U39183 (N_39183,N_36121,N_37667);
xnor U39184 (N_39184,N_36031,N_36283);
or U39185 (N_39185,N_36798,N_36104);
or U39186 (N_39186,N_37628,N_37508);
or U39187 (N_39187,N_36546,N_36801);
and U39188 (N_39188,N_36943,N_36532);
nand U39189 (N_39189,N_36984,N_37729);
or U39190 (N_39190,N_37938,N_37429);
and U39191 (N_39191,N_36774,N_37344);
nor U39192 (N_39192,N_37085,N_36601);
and U39193 (N_39193,N_36761,N_36188);
xor U39194 (N_39194,N_36583,N_37830);
nand U39195 (N_39195,N_36486,N_37490);
and U39196 (N_39196,N_37132,N_37650);
nand U39197 (N_39197,N_36457,N_36823);
xor U39198 (N_39198,N_37771,N_36349);
nor U39199 (N_39199,N_36145,N_37764);
or U39200 (N_39200,N_37398,N_37339);
xor U39201 (N_39201,N_37454,N_36732);
or U39202 (N_39202,N_36029,N_37017);
and U39203 (N_39203,N_36091,N_37562);
xnor U39204 (N_39204,N_36928,N_37315);
nor U39205 (N_39205,N_36159,N_36908);
nand U39206 (N_39206,N_37245,N_37247);
xnor U39207 (N_39207,N_36512,N_36526);
xnor U39208 (N_39208,N_36196,N_37573);
xnor U39209 (N_39209,N_37164,N_37527);
and U39210 (N_39210,N_37917,N_37134);
or U39211 (N_39211,N_36052,N_37312);
or U39212 (N_39212,N_36208,N_37736);
nand U39213 (N_39213,N_37913,N_37249);
or U39214 (N_39214,N_36380,N_36352);
and U39215 (N_39215,N_37229,N_37255);
nand U39216 (N_39216,N_36254,N_36288);
xor U39217 (N_39217,N_36655,N_37096);
and U39218 (N_39218,N_37358,N_37056);
and U39219 (N_39219,N_37698,N_36577);
xnor U39220 (N_39220,N_37033,N_37670);
nor U39221 (N_39221,N_36759,N_37593);
xor U39222 (N_39222,N_37640,N_36362);
nor U39223 (N_39223,N_36037,N_36815);
nor U39224 (N_39224,N_36418,N_37508);
and U39225 (N_39225,N_37525,N_37089);
nor U39226 (N_39226,N_36391,N_36982);
and U39227 (N_39227,N_37279,N_37423);
and U39228 (N_39228,N_36028,N_37329);
and U39229 (N_39229,N_37719,N_36242);
nor U39230 (N_39230,N_36849,N_36490);
nor U39231 (N_39231,N_36568,N_36001);
xor U39232 (N_39232,N_37165,N_37974);
and U39233 (N_39233,N_36651,N_36680);
xnor U39234 (N_39234,N_36861,N_37720);
and U39235 (N_39235,N_37377,N_36912);
and U39236 (N_39236,N_37927,N_37931);
xor U39237 (N_39237,N_36510,N_36924);
xnor U39238 (N_39238,N_37488,N_36772);
nand U39239 (N_39239,N_37934,N_37917);
nor U39240 (N_39240,N_36633,N_37001);
xnor U39241 (N_39241,N_37599,N_37699);
nand U39242 (N_39242,N_36953,N_36586);
nor U39243 (N_39243,N_37637,N_36931);
nor U39244 (N_39244,N_36874,N_37112);
or U39245 (N_39245,N_37524,N_36651);
nand U39246 (N_39246,N_36230,N_37627);
nand U39247 (N_39247,N_37743,N_36241);
nor U39248 (N_39248,N_37735,N_36765);
and U39249 (N_39249,N_36812,N_37978);
xnor U39250 (N_39250,N_37017,N_36824);
nor U39251 (N_39251,N_37712,N_36468);
and U39252 (N_39252,N_36056,N_37426);
xor U39253 (N_39253,N_37009,N_37653);
or U39254 (N_39254,N_36888,N_37838);
nand U39255 (N_39255,N_36377,N_37003);
or U39256 (N_39256,N_36932,N_37680);
and U39257 (N_39257,N_36660,N_36463);
nor U39258 (N_39258,N_37131,N_37581);
or U39259 (N_39259,N_37175,N_36516);
nor U39260 (N_39260,N_36311,N_36084);
and U39261 (N_39261,N_37307,N_36174);
nand U39262 (N_39262,N_37403,N_37936);
xor U39263 (N_39263,N_37806,N_36058);
and U39264 (N_39264,N_36387,N_36534);
and U39265 (N_39265,N_36911,N_37683);
nor U39266 (N_39266,N_36350,N_36137);
xor U39267 (N_39267,N_37124,N_36290);
or U39268 (N_39268,N_37088,N_37946);
nor U39269 (N_39269,N_36812,N_36659);
xnor U39270 (N_39270,N_36191,N_36409);
and U39271 (N_39271,N_36796,N_37858);
nand U39272 (N_39272,N_37082,N_36192);
xnor U39273 (N_39273,N_37496,N_36073);
nand U39274 (N_39274,N_37067,N_37954);
xor U39275 (N_39275,N_36192,N_36379);
nand U39276 (N_39276,N_36198,N_37157);
nand U39277 (N_39277,N_36948,N_37280);
xor U39278 (N_39278,N_36385,N_37983);
or U39279 (N_39279,N_37845,N_36108);
nor U39280 (N_39280,N_36700,N_36654);
and U39281 (N_39281,N_36707,N_36741);
nand U39282 (N_39282,N_36482,N_37039);
nand U39283 (N_39283,N_37568,N_37716);
and U39284 (N_39284,N_36755,N_36594);
nand U39285 (N_39285,N_37198,N_37792);
nor U39286 (N_39286,N_37094,N_37202);
nand U39287 (N_39287,N_37029,N_36143);
or U39288 (N_39288,N_36177,N_36821);
nor U39289 (N_39289,N_37229,N_36567);
xor U39290 (N_39290,N_37384,N_36196);
nor U39291 (N_39291,N_36857,N_36333);
or U39292 (N_39292,N_37850,N_37965);
and U39293 (N_39293,N_36829,N_37783);
xor U39294 (N_39294,N_36948,N_36936);
xor U39295 (N_39295,N_36245,N_37732);
xor U39296 (N_39296,N_36736,N_36972);
and U39297 (N_39297,N_37192,N_37053);
or U39298 (N_39298,N_37876,N_36471);
xor U39299 (N_39299,N_37405,N_36073);
or U39300 (N_39300,N_36090,N_36855);
nor U39301 (N_39301,N_36943,N_37336);
or U39302 (N_39302,N_37527,N_37973);
or U39303 (N_39303,N_36841,N_36160);
and U39304 (N_39304,N_36250,N_36359);
and U39305 (N_39305,N_36146,N_37842);
xor U39306 (N_39306,N_36671,N_37305);
xnor U39307 (N_39307,N_36138,N_37663);
or U39308 (N_39308,N_36098,N_37682);
xor U39309 (N_39309,N_36939,N_37114);
or U39310 (N_39310,N_37613,N_36778);
or U39311 (N_39311,N_37866,N_37142);
nor U39312 (N_39312,N_37977,N_37622);
xor U39313 (N_39313,N_37637,N_37811);
or U39314 (N_39314,N_37716,N_36468);
nand U39315 (N_39315,N_36012,N_37154);
xor U39316 (N_39316,N_37812,N_37052);
or U39317 (N_39317,N_37667,N_37171);
or U39318 (N_39318,N_37244,N_36709);
and U39319 (N_39319,N_37221,N_36455);
or U39320 (N_39320,N_37812,N_37666);
xnor U39321 (N_39321,N_36241,N_36159);
xor U39322 (N_39322,N_36244,N_37259);
xnor U39323 (N_39323,N_36307,N_37589);
or U39324 (N_39324,N_36825,N_37263);
nor U39325 (N_39325,N_37604,N_36002);
nor U39326 (N_39326,N_37017,N_37459);
xnor U39327 (N_39327,N_37687,N_36052);
and U39328 (N_39328,N_37071,N_36878);
nand U39329 (N_39329,N_37758,N_37992);
and U39330 (N_39330,N_36729,N_36736);
or U39331 (N_39331,N_36186,N_37976);
or U39332 (N_39332,N_37446,N_37545);
or U39333 (N_39333,N_37094,N_36964);
nor U39334 (N_39334,N_36390,N_37851);
or U39335 (N_39335,N_37394,N_37784);
xor U39336 (N_39336,N_37833,N_37777);
nand U39337 (N_39337,N_36652,N_37141);
and U39338 (N_39338,N_36030,N_36054);
xnor U39339 (N_39339,N_37537,N_36885);
nand U39340 (N_39340,N_37849,N_37309);
xnor U39341 (N_39341,N_37552,N_36164);
nor U39342 (N_39342,N_36750,N_37978);
xnor U39343 (N_39343,N_36798,N_37897);
or U39344 (N_39344,N_37846,N_37357);
nor U39345 (N_39345,N_37543,N_37067);
nand U39346 (N_39346,N_36461,N_36915);
nand U39347 (N_39347,N_36947,N_37764);
xor U39348 (N_39348,N_37772,N_36565);
and U39349 (N_39349,N_37618,N_37673);
nor U39350 (N_39350,N_36895,N_36333);
or U39351 (N_39351,N_37993,N_36123);
and U39352 (N_39352,N_37109,N_36456);
xnor U39353 (N_39353,N_36654,N_36114);
or U39354 (N_39354,N_37098,N_37937);
nor U39355 (N_39355,N_36031,N_37402);
nand U39356 (N_39356,N_36684,N_37977);
nor U39357 (N_39357,N_36863,N_36265);
nor U39358 (N_39358,N_37765,N_37965);
xnor U39359 (N_39359,N_37253,N_37912);
or U39360 (N_39360,N_37854,N_36621);
xor U39361 (N_39361,N_36582,N_37979);
nor U39362 (N_39362,N_36717,N_36016);
and U39363 (N_39363,N_37175,N_36131);
xor U39364 (N_39364,N_37832,N_37630);
or U39365 (N_39365,N_37170,N_36426);
nand U39366 (N_39366,N_36452,N_36041);
nor U39367 (N_39367,N_36601,N_36050);
or U39368 (N_39368,N_36019,N_36172);
nor U39369 (N_39369,N_37306,N_37683);
xor U39370 (N_39370,N_37329,N_36735);
xnor U39371 (N_39371,N_37330,N_36822);
or U39372 (N_39372,N_37476,N_37668);
xnor U39373 (N_39373,N_37294,N_36910);
nor U39374 (N_39374,N_36566,N_36240);
nor U39375 (N_39375,N_37472,N_36927);
or U39376 (N_39376,N_36011,N_36360);
nor U39377 (N_39377,N_36286,N_36763);
or U39378 (N_39378,N_36644,N_37412);
nor U39379 (N_39379,N_36686,N_36400);
xnor U39380 (N_39380,N_37457,N_36838);
or U39381 (N_39381,N_37688,N_37144);
nand U39382 (N_39382,N_37338,N_36364);
or U39383 (N_39383,N_37224,N_36130);
xnor U39384 (N_39384,N_36670,N_36156);
nand U39385 (N_39385,N_37036,N_36325);
nor U39386 (N_39386,N_37691,N_37593);
or U39387 (N_39387,N_36815,N_36664);
nand U39388 (N_39388,N_36991,N_36125);
xnor U39389 (N_39389,N_36321,N_36891);
and U39390 (N_39390,N_37396,N_36022);
nand U39391 (N_39391,N_37253,N_36690);
nor U39392 (N_39392,N_36343,N_36605);
xor U39393 (N_39393,N_36542,N_36551);
or U39394 (N_39394,N_37966,N_37454);
xor U39395 (N_39395,N_37243,N_37428);
nor U39396 (N_39396,N_36792,N_37450);
nand U39397 (N_39397,N_37681,N_37977);
nand U39398 (N_39398,N_36873,N_36570);
nand U39399 (N_39399,N_37457,N_36202);
xnor U39400 (N_39400,N_36714,N_37210);
and U39401 (N_39401,N_36302,N_37242);
and U39402 (N_39402,N_37681,N_37565);
or U39403 (N_39403,N_37374,N_36454);
nand U39404 (N_39404,N_37893,N_36157);
nor U39405 (N_39405,N_37039,N_37346);
nand U39406 (N_39406,N_36489,N_37432);
xnor U39407 (N_39407,N_37480,N_36560);
and U39408 (N_39408,N_36262,N_36931);
and U39409 (N_39409,N_36179,N_36797);
and U39410 (N_39410,N_37307,N_37285);
and U39411 (N_39411,N_37307,N_36166);
and U39412 (N_39412,N_36343,N_36670);
or U39413 (N_39413,N_36462,N_36281);
and U39414 (N_39414,N_37727,N_37409);
and U39415 (N_39415,N_36119,N_37445);
nor U39416 (N_39416,N_37315,N_36187);
nor U39417 (N_39417,N_36204,N_36592);
or U39418 (N_39418,N_37786,N_36784);
and U39419 (N_39419,N_37198,N_37126);
and U39420 (N_39420,N_36699,N_37632);
and U39421 (N_39421,N_36462,N_36614);
xnor U39422 (N_39422,N_36415,N_36730);
nor U39423 (N_39423,N_36467,N_36203);
xnor U39424 (N_39424,N_36759,N_36810);
xnor U39425 (N_39425,N_37252,N_36732);
and U39426 (N_39426,N_37392,N_36183);
xor U39427 (N_39427,N_36497,N_36387);
nor U39428 (N_39428,N_36203,N_37361);
and U39429 (N_39429,N_36902,N_37752);
or U39430 (N_39430,N_37059,N_36511);
nand U39431 (N_39431,N_37365,N_37113);
nor U39432 (N_39432,N_37057,N_37294);
or U39433 (N_39433,N_36926,N_36196);
xnor U39434 (N_39434,N_37705,N_37778);
or U39435 (N_39435,N_37410,N_37427);
and U39436 (N_39436,N_37441,N_36310);
nand U39437 (N_39437,N_37549,N_36853);
or U39438 (N_39438,N_36696,N_36742);
or U39439 (N_39439,N_36702,N_37993);
nand U39440 (N_39440,N_36663,N_36266);
nand U39441 (N_39441,N_36303,N_37785);
nor U39442 (N_39442,N_37920,N_36009);
nand U39443 (N_39443,N_36587,N_37474);
nand U39444 (N_39444,N_36274,N_37354);
nand U39445 (N_39445,N_37812,N_37200);
nor U39446 (N_39446,N_36865,N_37490);
nand U39447 (N_39447,N_37084,N_37853);
xor U39448 (N_39448,N_37862,N_36147);
and U39449 (N_39449,N_37563,N_36332);
and U39450 (N_39450,N_37167,N_37282);
xnor U39451 (N_39451,N_36447,N_36668);
nor U39452 (N_39452,N_37098,N_37683);
xor U39453 (N_39453,N_37057,N_37550);
or U39454 (N_39454,N_37973,N_36823);
nor U39455 (N_39455,N_36043,N_37495);
xnor U39456 (N_39456,N_37826,N_37026);
nor U39457 (N_39457,N_37536,N_36880);
nor U39458 (N_39458,N_37826,N_36950);
xor U39459 (N_39459,N_36329,N_37247);
or U39460 (N_39460,N_37725,N_36354);
nor U39461 (N_39461,N_37683,N_36276);
or U39462 (N_39462,N_37839,N_36126);
or U39463 (N_39463,N_37772,N_37214);
and U39464 (N_39464,N_36087,N_36410);
nor U39465 (N_39465,N_36838,N_37844);
and U39466 (N_39466,N_36118,N_37595);
nor U39467 (N_39467,N_36285,N_36022);
xnor U39468 (N_39468,N_37278,N_36922);
xor U39469 (N_39469,N_36930,N_36495);
or U39470 (N_39470,N_37419,N_36621);
and U39471 (N_39471,N_36559,N_37348);
nor U39472 (N_39472,N_36845,N_36414);
nor U39473 (N_39473,N_36710,N_37673);
nor U39474 (N_39474,N_37519,N_36942);
or U39475 (N_39475,N_37474,N_36385);
and U39476 (N_39476,N_37352,N_37947);
nor U39477 (N_39477,N_36576,N_37040);
nor U39478 (N_39478,N_37397,N_36581);
nor U39479 (N_39479,N_36557,N_37167);
xor U39480 (N_39480,N_37608,N_37220);
and U39481 (N_39481,N_36927,N_37167);
and U39482 (N_39482,N_36911,N_37811);
and U39483 (N_39483,N_37353,N_36634);
nor U39484 (N_39484,N_37220,N_36019);
nand U39485 (N_39485,N_36402,N_36720);
or U39486 (N_39486,N_36020,N_37546);
or U39487 (N_39487,N_37098,N_37839);
and U39488 (N_39488,N_36917,N_36907);
nand U39489 (N_39489,N_37771,N_36078);
nor U39490 (N_39490,N_36540,N_37724);
nand U39491 (N_39491,N_37525,N_36595);
nor U39492 (N_39492,N_36203,N_36584);
or U39493 (N_39493,N_36047,N_37178);
and U39494 (N_39494,N_36942,N_37123);
or U39495 (N_39495,N_37057,N_36663);
xnor U39496 (N_39496,N_36920,N_37818);
and U39497 (N_39497,N_37627,N_36125);
and U39498 (N_39498,N_36160,N_36287);
or U39499 (N_39499,N_36251,N_37656);
nand U39500 (N_39500,N_36576,N_36938);
nand U39501 (N_39501,N_36348,N_37060);
and U39502 (N_39502,N_36578,N_37918);
or U39503 (N_39503,N_37865,N_36785);
nand U39504 (N_39504,N_36151,N_37348);
or U39505 (N_39505,N_37718,N_37771);
nand U39506 (N_39506,N_37414,N_37338);
and U39507 (N_39507,N_36075,N_36572);
nand U39508 (N_39508,N_36996,N_36810);
or U39509 (N_39509,N_37764,N_36254);
nand U39510 (N_39510,N_36415,N_37255);
or U39511 (N_39511,N_36815,N_36895);
nor U39512 (N_39512,N_36823,N_36308);
nand U39513 (N_39513,N_36683,N_37942);
xnor U39514 (N_39514,N_36552,N_37944);
nor U39515 (N_39515,N_36230,N_36172);
and U39516 (N_39516,N_37703,N_37097);
nand U39517 (N_39517,N_37679,N_36598);
nand U39518 (N_39518,N_36322,N_37139);
nor U39519 (N_39519,N_37985,N_36281);
nand U39520 (N_39520,N_36410,N_36771);
xnor U39521 (N_39521,N_36646,N_36001);
and U39522 (N_39522,N_36304,N_37986);
nand U39523 (N_39523,N_37883,N_37198);
nand U39524 (N_39524,N_37216,N_37950);
xor U39525 (N_39525,N_36773,N_37957);
xor U39526 (N_39526,N_37426,N_36375);
and U39527 (N_39527,N_37957,N_37138);
xor U39528 (N_39528,N_36969,N_36061);
or U39529 (N_39529,N_37099,N_37482);
and U39530 (N_39530,N_37249,N_37588);
or U39531 (N_39531,N_36745,N_36039);
and U39532 (N_39532,N_37386,N_36801);
nand U39533 (N_39533,N_36081,N_37894);
nand U39534 (N_39534,N_37859,N_37543);
or U39535 (N_39535,N_36098,N_36973);
xnor U39536 (N_39536,N_37184,N_37614);
xnor U39537 (N_39537,N_36963,N_36409);
nand U39538 (N_39538,N_37051,N_36956);
xnor U39539 (N_39539,N_36647,N_37670);
nor U39540 (N_39540,N_37768,N_37765);
and U39541 (N_39541,N_37347,N_36408);
or U39542 (N_39542,N_37748,N_36952);
xor U39543 (N_39543,N_37544,N_37857);
nor U39544 (N_39544,N_37134,N_36528);
nor U39545 (N_39545,N_36330,N_37696);
nor U39546 (N_39546,N_36438,N_37446);
nor U39547 (N_39547,N_37563,N_36747);
nand U39548 (N_39548,N_37313,N_37378);
nor U39549 (N_39549,N_36903,N_37126);
nand U39550 (N_39550,N_36302,N_36832);
and U39551 (N_39551,N_36327,N_36489);
and U39552 (N_39552,N_37094,N_36120);
nor U39553 (N_39553,N_36684,N_37158);
xnor U39554 (N_39554,N_37613,N_36996);
xnor U39555 (N_39555,N_37052,N_36379);
or U39556 (N_39556,N_36598,N_37041);
xnor U39557 (N_39557,N_36181,N_37073);
and U39558 (N_39558,N_37148,N_37743);
xor U39559 (N_39559,N_36152,N_37698);
xor U39560 (N_39560,N_37195,N_36075);
xnor U39561 (N_39561,N_37368,N_37380);
nor U39562 (N_39562,N_37793,N_37865);
and U39563 (N_39563,N_37418,N_36227);
nand U39564 (N_39564,N_36283,N_37220);
nand U39565 (N_39565,N_37978,N_36460);
xnor U39566 (N_39566,N_36533,N_37282);
or U39567 (N_39567,N_37199,N_37865);
nand U39568 (N_39568,N_37984,N_36940);
or U39569 (N_39569,N_37938,N_37675);
nand U39570 (N_39570,N_37955,N_36241);
nor U39571 (N_39571,N_37886,N_36252);
or U39572 (N_39572,N_36523,N_36227);
and U39573 (N_39573,N_37383,N_36473);
and U39574 (N_39574,N_37606,N_37261);
and U39575 (N_39575,N_37665,N_37151);
nand U39576 (N_39576,N_36315,N_36740);
nor U39577 (N_39577,N_37679,N_37807);
and U39578 (N_39578,N_36884,N_37887);
or U39579 (N_39579,N_37900,N_37585);
and U39580 (N_39580,N_37411,N_37583);
nor U39581 (N_39581,N_36439,N_37606);
nor U39582 (N_39582,N_36373,N_37337);
or U39583 (N_39583,N_36747,N_37360);
or U39584 (N_39584,N_36449,N_36073);
nor U39585 (N_39585,N_37145,N_37039);
nand U39586 (N_39586,N_37680,N_37637);
nand U39587 (N_39587,N_37510,N_37515);
and U39588 (N_39588,N_36361,N_36521);
xnor U39589 (N_39589,N_36913,N_36609);
or U39590 (N_39590,N_37095,N_37014);
nand U39591 (N_39591,N_36452,N_36723);
nand U39592 (N_39592,N_37148,N_37785);
xor U39593 (N_39593,N_37325,N_37515);
and U39594 (N_39594,N_37164,N_36683);
nor U39595 (N_39595,N_36725,N_36605);
or U39596 (N_39596,N_37327,N_36514);
and U39597 (N_39597,N_37448,N_37780);
xnor U39598 (N_39598,N_36820,N_36797);
and U39599 (N_39599,N_36002,N_36905);
nand U39600 (N_39600,N_36363,N_37557);
xor U39601 (N_39601,N_36314,N_37746);
nor U39602 (N_39602,N_36672,N_37957);
or U39603 (N_39603,N_36423,N_37778);
nor U39604 (N_39604,N_37712,N_37977);
and U39605 (N_39605,N_36663,N_36957);
and U39606 (N_39606,N_36394,N_36010);
or U39607 (N_39607,N_37862,N_36854);
xnor U39608 (N_39608,N_36802,N_36992);
nor U39609 (N_39609,N_37478,N_37283);
xor U39610 (N_39610,N_37970,N_37890);
and U39611 (N_39611,N_36437,N_36823);
or U39612 (N_39612,N_36327,N_37697);
nor U39613 (N_39613,N_36354,N_36800);
nand U39614 (N_39614,N_37003,N_37167);
and U39615 (N_39615,N_37389,N_37928);
nor U39616 (N_39616,N_37735,N_37641);
or U39617 (N_39617,N_37174,N_36206);
and U39618 (N_39618,N_36990,N_36703);
nor U39619 (N_39619,N_37882,N_37559);
or U39620 (N_39620,N_36186,N_36456);
or U39621 (N_39621,N_36020,N_37271);
nand U39622 (N_39622,N_36470,N_37191);
nand U39623 (N_39623,N_36303,N_37683);
or U39624 (N_39624,N_36531,N_37964);
nand U39625 (N_39625,N_37592,N_36208);
nand U39626 (N_39626,N_37983,N_37022);
nand U39627 (N_39627,N_37445,N_37108);
and U39628 (N_39628,N_37895,N_36047);
and U39629 (N_39629,N_36911,N_37933);
nand U39630 (N_39630,N_37911,N_36819);
xnor U39631 (N_39631,N_36051,N_37522);
or U39632 (N_39632,N_37540,N_36422);
nor U39633 (N_39633,N_37483,N_37318);
nor U39634 (N_39634,N_37239,N_36446);
nand U39635 (N_39635,N_36771,N_36613);
xnor U39636 (N_39636,N_36911,N_37343);
or U39637 (N_39637,N_37798,N_36567);
nor U39638 (N_39638,N_36915,N_37615);
and U39639 (N_39639,N_37836,N_37601);
xnor U39640 (N_39640,N_36565,N_37741);
nand U39641 (N_39641,N_37938,N_36311);
nand U39642 (N_39642,N_37897,N_37137);
and U39643 (N_39643,N_36466,N_36917);
nand U39644 (N_39644,N_37328,N_36345);
or U39645 (N_39645,N_36562,N_36674);
nand U39646 (N_39646,N_37356,N_36758);
nor U39647 (N_39647,N_36014,N_36666);
nand U39648 (N_39648,N_36907,N_37113);
nand U39649 (N_39649,N_36218,N_36330);
xnor U39650 (N_39650,N_36558,N_37999);
or U39651 (N_39651,N_37284,N_37222);
or U39652 (N_39652,N_37000,N_36265);
xnor U39653 (N_39653,N_36339,N_37930);
and U39654 (N_39654,N_37178,N_37359);
or U39655 (N_39655,N_37335,N_36939);
nand U39656 (N_39656,N_36421,N_37320);
xnor U39657 (N_39657,N_36530,N_36593);
or U39658 (N_39658,N_37196,N_36146);
or U39659 (N_39659,N_37916,N_36443);
nor U39660 (N_39660,N_36195,N_36173);
nor U39661 (N_39661,N_37580,N_36408);
xor U39662 (N_39662,N_37419,N_36415);
xor U39663 (N_39663,N_36366,N_36558);
and U39664 (N_39664,N_37103,N_37499);
or U39665 (N_39665,N_37272,N_37420);
xnor U39666 (N_39666,N_37411,N_37567);
nand U39667 (N_39667,N_36579,N_36963);
nand U39668 (N_39668,N_36002,N_36599);
nor U39669 (N_39669,N_36229,N_36614);
xnor U39670 (N_39670,N_36293,N_36935);
nand U39671 (N_39671,N_36346,N_36135);
or U39672 (N_39672,N_36954,N_37303);
nand U39673 (N_39673,N_37378,N_36672);
nand U39674 (N_39674,N_37194,N_37782);
or U39675 (N_39675,N_36043,N_37936);
and U39676 (N_39676,N_36135,N_36204);
nor U39677 (N_39677,N_36232,N_36585);
nand U39678 (N_39678,N_36559,N_36511);
nor U39679 (N_39679,N_36072,N_37974);
xor U39680 (N_39680,N_36306,N_36308);
and U39681 (N_39681,N_36905,N_37226);
xnor U39682 (N_39682,N_36666,N_37473);
and U39683 (N_39683,N_36757,N_36098);
nor U39684 (N_39684,N_37472,N_37188);
or U39685 (N_39685,N_37959,N_37902);
and U39686 (N_39686,N_36588,N_37683);
or U39687 (N_39687,N_36729,N_36064);
xor U39688 (N_39688,N_36440,N_37406);
nand U39689 (N_39689,N_37053,N_37463);
and U39690 (N_39690,N_36380,N_37584);
or U39691 (N_39691,N_37147,N_37995);
nor U39692 (N_39692,N_36040,N_36214);
and U39693 (N_39693,N_37523,N_37421);
nor U39694 (N_39694,N_36764,N_36822);
nand U39695 (N_39695,N_36669,N_36960);
or U39696 (N_39696,N_36960,N_37484);
nand U39697 (N_39697,N_37969,N_37447);
xnor U39698 (N_39698,N_36401,N_37090);
or U39699 (N_39699,N_37884,N_37453);
nor U39700 (N_39700,N_36339,N_37831);
xnor U39701 (N_39701,N_36981,N_36513);
or U39702 (N_39702,N_37289,N_37539);
or U39703 (N_39703,N_37048,N_36140);
or U39704 (N_39704,N_36647,N_36527);
xnor U39705 (N_39705,N_36987,N_36302);
nand U39706 (N_39706,N_36146,N_37021);
or U39707 (N_39707,N_36328,N_37528);
nor U39708 (N_39708,N_36958,N_37679);
or U39709 (N_39709,N_36175,N_37512);
xor U39710 (N_39710,N_37635,N_37295);
or U39711 (N_39711,N_37019,N_36958);
nand U39712 (N_39712,N_36096,N_37387);
or U39713 (N_39713,N_37475,N_36851);
or U39714 (N_39714,N_37942,N_37691);
nand U39715 (N_39715,N_36362,N_37136);
xnor U39716 (N_39716,N_36120,N_37134);
nand U39717 (N_39717,N_36274,N_37821);
nand U39718 (N_39718,N_36631,N_37833);
or U39719 (N_39719,N_37103,N_37082);
or U39720 (N_39720,N_36700,N_37476);
or U39721 (N_39721,N_37545,N_36340);
nand U39722 (N_39722,N_36029,N_36496);
nand U39723 (N_39723,N_36426,N_36787);
nor U39724 (N_39724,N_36766,N_37452);
and U39725 (N_39725,N_37923,N_36350);
and U39726 (N_39726,N_36160,N_36204);
or U39727 (N_39727,N_36144,N_37829);
or U39728 (N_39728,N_37738,N_37169);
or U39729 (N_39729,N_36959,N_37139);
nor U39730 (N_39730,N_36239,N_37327);
and U39731 (N_39731,N_37403,N_36419);
xor U39732 (N_39732,N_37177,N_36534);
nand U39733 (N_39733,N_36067,N_37150);
or U39734 (N_39734,N_36963,N_37845);
or U39735 (N_39735,N_36261,N_36634);
or U39736 (N_39736,N_37385,N_36125);
nor U39737 (N_39737,N_36996,N_37744);
nand U39738 (N_39738,N_36216,N_36603);
and U39739 (N_39739,N_36399,N_37682);
nor U39740 (N_39740,N_37480,N_36229);
nand U39741 (N_39741,N_37354,N_37542);
xnor U39742 (N_39742,N_36052,N_36373);
and U39743 (N_39743,N_37114,N_36196);
nor U39744 (N_39744,N_36542,N_37659);
and U39745 (N_39745,N_36765,N_36990);
and U39746 (N_39746,N_36360,N_36729);
nand U39747 (N_39747,N_36683,N_36486);
nand U39748 (N_39748,N_37480,N_36045);
and U39749 (N_39749,N_36053,N_36679);
and U39750 (N_39750,N_37331,N_36038);
nor U39751 (N_39751,N_36500,N_37974);
xor U39752 (N_39752,N_37964,N_37077);
or U39753 (N_39753,N_36438,N_37661);
xor U39754 (N_39754,N_36590,N_37529);
nand U39755 (N_39755,N_36544,N_37846);
or U39756 (N_39756,N_37169,N_37619);
xor U39757 (N_39757,N_36851,N_37929);
xnor U39758 (N_39758,N_37743,N_36592);
or U39759 (N_39759,N_37347,N_36684);
xor U39760 (N_39760,N_37361,N_36747);
and U39761 (N_39761,N_37507,N_36079);
nor U39762 (N_39762,N_37435,N_37529);
and U39763 (N_39763,N_36741,N_36234);
and U39764 (N_39764,N_36207,N_37253);
or U39765 (N_39765,N_37656,N_36625);
xnor U39766 (N_39766,N_37710,N_37119);
xnor U39767 (N_39767,N_37376,N_37246);
or U39768 (N_39768,N_36237,N_36614);
xor U39769 (N_39769,N_36418,N_36145);
nand U39770 (N_39770,N_37834,N_36319);
or U39771 (N_39771,N_37186,N_37283);
or U39772 (N_39772,N_36799,N_37514);
and U39773 (N_39773,N_37830,N_36492);
or U39774 (N_39774,N_36263,N_36670);
or U39775 (N_39775,N_37273,N_37159);
nor U39776 (N_39776,N_37942,N_37158);
nor U39777 (N_39777,N_36439,N_36254);
or U39778 (N_39778,N_36904,N_37565);
and U39779 (N_39779,N_36691,N_36800);
xnor U39780 (N_39780,N_36821,N_36130);
nand U39781 (N_39781,N_37181,N_37865);
or U39782 (N_39782,N_37916,N_36885);
and U39783 (N_39783,N_36473,N_36849);
or U39784 (N_39784,N_37876,N_36719);
nand U39785 (N_39785,N_36810,N_36526);
nand U39786 (N_39786,N_37822,N_37251);
nand U39787 (N_39787,N_36760,N_36995);
nor U39788 (N_39788,N_37276,N_37825);
xnor U39789 (N_39789,N_36334,N_37868);
and U39790 (N_39790,N_36790,N_37228);
xor U39791 (N_39791,N_37790,N_36659);
and U39792 (N_39792,N_37828,N_37763);
nand U39793 (N_39793,N_36770,N_36235);
nor U39794 (N_39794,N_37900,N_36614);
or U39795 (N_39795,N_37194,N_36744);
or U39796 (N_39796,N_36121,N_36233);
xor U39797 (N_39797,N_37976,N_36013);
xor U39798 (N_39798,N_36438,N_36339);
xor U39799 (N_39799,N_37928,N_36692);
nand U39800 (N_39800,N_37906,N_37806);
nand U39801 (N_39801,N_37120,N_37718);
xor U39802 (N_39802,N_37782,N_37495);
and U39803 (N_39803,N_36293,N_36601);
xnor U39804 (N_39804,N_37232,N_37144);
and U39805 (N_39805,N_37630,N_37211);
and U39806 (N_39806,N_37410,N_36292);
nor U39807 (N_39807,N_36206,N_37650);
xnor U39808 (N_39808,N_37335,N_36741);
or U39809 (N_39809,N_36218,N_37932);
nor U39810 (N_39810,N_37609,N_37506);
nor U39811 (N_39811,N_36571,N_36942);
nor U39812 (N_39812,N_37329,N_36493);
or U39813 (N_39813,N_37502,N_37988);
and U39814 (N_39814,N_37736,N_36813);
xor U39815 (N_39815,N_37652,N_36977);
nand U39816 (N_39816,N_37926,N_37858);
and U39817 (N_39817,N_37243,N_36902);
or U39818 (N_39818,N_36991,N_37260);
nand U39819 (N_39819,N_37685,N_36982);
nand U39820 (N_39820,N_37429,N_36789);
xor U39821 (N_39821,N_36763,N_36061);
nor U39822 (N_39822,N_37130,N_36455);
or U39823 (N_39823,N_37727,N_36043);
and U39824 (N_39824,N_37269,N_37851);
and U39825 (N_39825,N_37585,N_37355);
nand U39826 (N_39826,N_36367,N_37406);
nor U39827 (N_39827,N_37475,N_37565);
nand U39828 (N_39828,N_37144,N_37170);
or U39829 (N_39829,N_36860,N_36475);
or U39830 (N_39830,N_36981,N_37364);
nand U39831 (N_39831,N_37990,N_37579);
nor U39832 (N_39832,N_36363,N_37259);
and U39833 (N_39833,N_37496,N_36282);
and U39834 (N_39834,N_36287,N_36275);
nor U39835 (N_39835,N_37940,N_36849);
nand U39836 (N_39836,N_36779,N_37193);
and U39837 (N_39837,N_37780,N_37602);
and U39838 (N_39838,N_36169,N_37408);
and U39839 (N_39839,N_36306,N_37865);
and U39840 (N_39840,N_36155,N_36542);
and U39841 (N_39841,N_37661,N_37760);
or U39842 (N_39842,N_37044,N_37714);
xnor U39843 (N_39843,N_36956,N_37267);
or U39844 (N_39844,N_37970,N_37015);
xnor U39845 (N_39845,N_36193,N_37414);
nor U39846 (N_39846,N_36826,N_37299);
nor U39847 (N_39847,N_37017,N_37749);
nand U39848 (N_39848,N_37394,N_37631);
nand U39849 (N_39849,N_36510,N_37683);
nand U39850 (N_39850,N_37327,N_36395);
or U39851 (N_39851,N_36117,N_37323);
or U39852 (N_39852,N_36155,N_36364);
xor U39853 (N_39853,N_37444,N_36455);
or U39854 (N_39854,N_37572,N_37956);
nor U39855 (N_39855,N_36712,N_36997);
nand U39856 (N_39856,N_36700,N_36760);
and U39857 (N_39857,N_36370,N_36851);
and U39858 (N_39858,N_36656,N_37738);
xnor U39859 (N_39859,N_37634,N_36632);
nand U39860 (N_39860,N_37741,N_36055);
nor U39861 (N_39861,N_37675,N_36409);
and U39862 (N_39862,N_37575,N_37324);
xnor U39863 (N_39863,N_37573,N_36815);
nand U39864 (N_39864,N_36746,N_36030);
or U39865 (N_39865,N_37065,N_36939);
xnor U39866 (N_39866,N_37735,N_37102);
xor U39867 (N_39867,N_36015,N_36868);
and U39868 (N_39868,N_36410,N_37151);
or U39869 (N_39869,N_36695,N_36337);
nand U39870 (N_39870,N_37298,N_36107);
nor U39871 (N_39871,N_37551,N_37138);
nor U39872 (N_39872,N_37444,N_37552);
and U39873 (N_39873,N_36446,N_37956);
xnor U39874 (N_39874,N_37663,N_36483);
and U39875 (N_39875,N_37309,N_37965);
xor U39876 (N_39876,N_36042,N_36271);
and U39877 (N_39877,N_37667,N_36661);
and U39878 (N_39878,N_36424,N_36019);
nor U39879 (N_39879,N_37180,N_37980);
and U39880 (N_39880,N_37676,N_37501);
nand U39881 (N_39881,N_37401,N_36176);
xnor U39882 (N_39882,N_37622,N_37700);
and U39883 (N_39883,N_36941,N_36644);
xor U39884 (N_39884,N_36120,N_36712);
and U39885 (N_39885,N_37958,N_36835);
and U39886 (N_39886,N_36356,N_37612);
nand U39887 (N_39887,N_37118,N_36366);
or U39888 (N_39888,N_36986,N_36093);
xnor U39889 (N_39889,N_37684,N_37835);
and U39890 (N_39890,N_37380,N_36329);
or U39891 (N_39891,N_36218,N_37174);
nor U39892 (N_39892,N_36822,N_36235);
xor U39893 (N_39893,N_36478,N_37969);
and U39894 (N_39894,N_36765,N_36799);
and U39895 (N_39895,N_36986,N_36138);
or U39896 (N_39896,N_37437,N_37960);
nor U39897 (N_39897,N_36791,N_36543);
nor U39898 (N_39898,N_37418,N_37315);
nor U39899 (N_39899,N_36897,N_37747);
xor U39900 (N_39900,N_36225,N_37287);
and U39901 (N_39901,N_36125,N_37933);
nor U39902 (N_39902,N_37562,N_37488);
xnor U39903 (N_39903,N_36873,N_36920);
nand U39904 (N_39904,N_37779,N_36230);
nand U39905 (N_39905,N_36866,N_36275);
nand U39906 (N_39906,N_36618,N_36566);
and U39907 (N_39907,N_36802,N_36210);
xnor U39908 (N_39908,N_37490,N_36840);
or U39909 (N_39909,N_37162,N_36817);
xor U39910 (N_39910,N_37218,N_36729);
or U39911 (N_39911,N_37543,N_36116);
xor U39912 (N_39912,N_37610,N_37642);
and U39913 (N_39913,N_36915,N_36037);
nor U39914 (N_39914,N_37282,N_36201);
or U39915 (N_39915,N_36262,N_36463);
nand U39916 (N_39916,N_37661,N_37569);
nand U39917 (N_39917,N_36032,N_37463);
or U39918 (N_39918,N_36295,N_37928);
and U39919 (N_39919,N_36207,N_37620);
and U39920 (N_39920,N_37539,N_37177);
or U39921 (N_39921,N_37419,N_36205);
and U39922 (N_39922,N_37967,N_37272);
nand U39923 (N_39923,N_36645,N_36672);
nor U39924 (N_39924,N_37457,N_37312);
and U39925 (N_39925,N_37700,N_37657);
nor U39926 (N_39926,N_37334,N_36935);
and U39927 (N_39927,N_36399,N_37378);
xor U39928 (N_39928,N_37956,N_36191);
xnor U39929 (N_39929,N_37948,N_37029);
xor U39930 (N_39930,N_36059,N_37568);
and U39931 (N_39931,N_37429,N_37004);
or U39932 (N_39932,N_37960,N_37530);
and U39933 (N_39933,N_36419,N_36819);
and U39934 (N_39934,N_36601,N_36040);
xor U39935 (N_39935,N_36727,N_37599);
and U39936 (N_39936,N_36509,N_37957);
or U39937 (N_39937,N_37826,N_37650);
nor U39938 (N_39938,N_36744,N_36501);
or U39939 (N_39939,N_36290,N_37307);
nand U39940 (N_39940,N_36903,N_37809);
or U39941 (N_39941,N_36332,N_36506);
xor U39942 (N_39942,N_37200,N_36437);
xor U39943 (N_39943,N_37176,N_37670);
and U39944 (N_39944,N_36066,N_37875);
nor U39945 (N_39945,N_36459,N_36715);
xor U39946 (N_39946,N_36252,N_36980);
or U39947 (N_39947,N_37165,N_36126);
xnor U39948 (N_39948,N_36218,N_36414);
nor U39949 (N_39949,N_36222,N_36063);
xnor U39950 (N_39950,N_37608,N_36963);
or U39951 (N_39951,N_37800,N_37182);
or U39952 (N_39952,N_37350,N_37434);
nor U39953 (N_39953,N_37935,N_37192);
xor U39954 (N_39954,N_36436,N_36287);
or U39955 (N_39955,N_37450,N_37997);
nor U39956 (N_39956,N_36946,N_36300);
xor U39957 (N_39957,N_37950,N_37958);
xor U39958 (N_39958,N_37073,N_36863);
and U39959 (N_39959,N_37153,N_36218);
nor U39960 (N_39960,N_37962,N_36059);
or U39961 (N_39961,N_37444,N_36414);
and U39962 (N_39962,N_37026,N_37899);
xor U39963 (N_39963,N_37797,N_37166);
and U39964 (N_39964,N_37335,N_36756);
or U39965 (N_39965,N_37745,N_36896);
nor U39966 (N_39966,N_36301,N_36039);
nand U39967 (N_39967,N_37480,N_37462);
or U39968 (N_39968,N_37277,N_37536);
or U39969 (N_39969,N_37433,N_37874);
nor U39970 (N_39970,N_37768,N_37596);
nand U39971 (N_39971,N_37543,N_37269);
nor U39972 (N_39972,N_37784,N_36816);
and U39973 (N_39973,N_37629,N_36939);
nor U39974 (N_39974,N_36659,N_36421);
nand U39975 (N_39975,N_37426,N_37952);
or U39976 (N_39976,N_36077,N_36501);
or U39977 (N_39977,N_36022,N_37231);
xnor U39978 (N_39978,N_36825,N_36347);
and U39979 (N_39979,N_37567,N_36033);
or U39980 (N_39980,N_37645,N_37497);
nand U39981 (N_39981,N_37321,N_36552);
nor U39982 (N_39982,N_36004,N_36599);
and U39983 (N_39983,N_36050,N_37946);
nand U39984 (N_39984,N_37232,N_37224);
xnor U39985 (N_39985,N_36166,N_37655);
or U39986 (N_39986,N_37764,N_36883);
nand U39987 (N_39987,N_36386,N_36642);
nand U39988 (N_39988,N_37986,N_36897);
nand U39989 (N_39989,N_37017,N_37309);
nor U39990 (N_39990,N_37912,N_37482);
or U39991 (N_39991,N_36248,N_37866);
nand U39992 (N_39992,N_36554,N_37741);
nor U39993 (N_39993,N_36563,N_36952);
or U39994 (N_39994,N_36291,N_37182);
or U39995 (N_39995,N_36175,N_36222);
nor U39996 (N_39996,N_37770,N_36210);
and U39997 (N_39997,N_36098,N_37825);
nor U39998 (N_39998,N_37826,N_36021);
xor U39999 (N_39999,N_37395,N_37468);
nand U40000 (N_40000,N_38352,N_39277);
and U40001 (N_40001,N_39482,N_39317);
or U40002 (N_40002,N_39769,N_38771);
or U40003 (N_40003,N_39799,N_38971);
xor U40004 (N_40004,N_38322,N_39551);
nor U40005 (N_40005,N_38492,N_39547);
nor U40006 (N_40006,N_38877,N_39601);
xor U40007 (N_40007,N_38052,N_38676);
xnor U40008 (N_40008,N_39820,N_39921);
xnor U40009 (N_40009,N_38592,N_38516);
xor U40010 (N_40010,N_39886,N_38926);
or U40011 (N_40011,N_39285,N_38651);
nand U40012 (N_40012,N_39944,N_38759);
nand U40013 (N_40013,N_38143,N_38479);
nor U40014 (N_40014,N_38308,N_38266);
and U40015 (N_40015,N_38774,N_39696);
and U40016 (N_40016,N_39230,N_38998);
nand U40017 (N_40017,N_39902,N_39903);
and U40018 (N_40018,N_38122,N_39855);
nand U40019 (N_40019,N_39719,N_39890);
nand U40020 (N_40020,N_38001,N_39037);
nor U40021 (N_40021,N_39392,N_38554);
or U40022 (N_40022,N_39324,N_38798);
xnor U40023 (N_40023,N_39045,N_38329);
nor U40024 (N_40024,N_39202,N_39728);
and U40025 (N_40025,N_38232,N_38347);
nand U40026 (N_40026,N_39309,N_38591);
and U40027 (N_40027,N_39727,N_38723);
xor U40028 (N_40028,N_39917,N_38536);
nand U40029 (N_40029,N_39137,N_38740);
and U40030 (N_40030,N_38934,N_39621);
nor U40031 (N_40031,N_39009,N_39827);
nor U40032 (N_40032,N_39339,N_38870);
or U40033 (N_40033,N_39748,N_38303);
or U40034 (N_40034,N_39068,N_38588);
nand U40035 (N_40035,N_38027,N_38689);
and U40036 (N_40036,N_38099,N_39371);
xor U40037 (N_40037,N_38522,N_38396);
xor U40038 (N_40038,N_39969,N_38050);
nand U40039 (N_40039,N_39079,N_39311);
nand U40040 (N_40040,N_39543,N_38420);
and U40041 (N_40041,N_39821,N_38264);
and U40042 (N_40042,N_39489,N_39025);
nand U40043 (N_40043,N_38658,N_38355);
xor U40044 (N_40044,N_39826,N_38685);
or U40045 (N_40045,N_39987,N_38807);
xnor U40046 (N_40046,N_38333,N_39284);
or U40047 (N_40047,N_38278,N_39302);
or U40048 (N_40048,N_39367,N_39970);
or U40049 (N_40049,N_39138,N_38060);
or U40050 (N_40050,N_38924,N_38353);
nand U40051 (N_40051,N_39982,N_39135);
xnor U40052 (N_40052,N_38660,N_38513);
and U40053 (N_40053,N_39802,N_38974);
nor U40054 (N_40054,N_39542,N_39964);
nor U40055 (N_40055,N_39468,N_38416);
and U40056 (N_40056,N_39789,N_39618);
nand U40057 (N_40057,N_39851,N_38828);
xor U40058 (N_40058,N_38106,N_39548);
nand U40059 (N_40059,N_38512,N_38496);
or U40060 (N_40060,N_39117,N_38767);
or U40061 (N_40061,N_38571,N_38943);
xor U40062 (N_40062,N_38925,N_38020);
xnor U40063 (N_40063,N_38721,N_39130);
and U40064 (N_40064,N_39120,N_39654);
nor U40065 (N_40065,N_39262,N_39582);
xnor U40066 (N_40066,N_38640,N_38575);
and U40067 (N_40067,N_39775,N_38008);
and U40068 (N_40068,N_38917,N_39141);
xor U40069 (N_40069,N_39522,N_39749);
and U40070 (N_40070,N_38747,N_39761);
nand U40071 (N_40071,N_38968,N_38904);
nand U40072 (N_40072,N_38049,N_38922);
nor U40073 (N_40073,N_38059,N_38235);
and U40074 (N_40074,N_38826,N_39980);
xor U40075 (N_40075,N_39819,N_39013);
xor U40076 (N_40076,N_38582,N_38371);
or U40077 (N_40077,N_38775,N_38977);
nand U40078 (N_40078,N_38190,N_38247);
nand U40079 (N_40079,N_38734,N_38868);
or U40080 (N_40080,N_38984,N_38195);
nor U40081 (N_40081,N_38644,N_39810);
nor U40082 (N_40082,N_38800,N_39163);
xnor U40083 (N_40083,N_39579,N_39648);
nand U40084 (N_40084,N_39668,N_39145);
xor U40085 (N_40085,N_39707,N_39082);
and U40086 (N_40086,N_38490,N_38434);
nand U40087 (N_40087,N_39070,N_38538);
or U40088 (N_40088,N_39357,N_39513);
or U40089 (N_40089,N_39923,N_39467);
or U40090 (N_40090,N_38158,N_39104);
nand U40091 (N_40091,N_38900,N_39994);
or U40092 (N_40092,N_39651,N_39213);
nand U40093 (N_40093,N_39625,N_39047);
nor U40094 (N_40094,N_39714,N_39538);
and U40095 (N_40095,N_38550,N_39283);
or U40096 (N_40096,N_38577,N_39471);
xor U40097 (N_40097,N_39591,N_38441);
nor U40098 (N_40098,N_38350,N_39126);
nor U40099 (N_40099,N_39349,N_39729);
xnor U40100 (N_40100,N_38294,N_39111);
and U40101 (N_40101,N_38309,N_38526);
nor U40102 (N_40102,N_39927,N_38764);
nand U40103 (N_40103,N_38340,N_38555);
nand U40104 (N_40104,N_39530,N_38446);
or U40105 (N_40105,N_38908,N_38331);
and U40106 (N_40106,N_38220,N_38273);
nand U40107 (N_40107,N_39469,N_38482);
and U40108 (N_40108,N_39605,N_38817);
and U40109 (N_40109,N_38464,N_38346);
nand U40110 (N_40110,N_38727,N_38141);
xnor U40111 (N_40111,N_39377,N_38343);
xor U40112 (N_40112,N_38756,N_38992);
or U40113 (N_40113,N_39389,N_38657);
nand U40114 (N_40114,N_38123,N_38149);
xnor U40115 (N_40115,N_39143,N_39131);
and U40116 (N_40116,N_39878,N_38822);
xnor U40117 (N_40117,N_39912,N_38041);
nand U40118 (N_40118,N_39798,N_38722);
and U40119 (N_40119,N_38717,N_38988);
nor U40120 (N_40120,N_39694,N_38576);
xor U40121 (N_40121,N_39514,N_38133);
xor U40122 (N_40122,N_39448,N_38911);
nand U40123 (N_40123,N_39385,N_39107);
xor U40124 (N_40124,N_38259,N_38541);
and U40125 (N_40125,N_38091,N_38025);
nand U40126 (N_40126,N_39611,N_38458);
xnor U40127 (N_40127,N_38077,N_39937);
and U40128 (N_40128,N_39910,N_39843);
nor U40129 (N_40129,N_39140,N_38480);
nand U40130 (N_40130,N_38587,N_39847);
nor U40131 (N_40131,N_38944,N_38344);
nor U40132 (N_40132,N_39326,N_39413);
nand U40133 (N_40133,N_39716,N_38207);
and U40134 (N_40134,N_38426,N_39697);
and U40135 (N_40135,N_38489,N_38015);
nor U40136 (N_40136,N_39663,N_38214);
xor U40137 (N_40137,N_38750,N_38965);
and U40138 (N_40138,N_39331,N_38230);
nor U40139 (N_40139,N_39414,N_38138);
xnor U40140 (N_40140,N_39508,N_39372);
xnor U40141 (N_40141,N_38929,N_38384);
xor U40142 (N_40142,N_39444,N_38982);
xnor U40143 (N_40143,N_39201,N_38263);
and U40144 (N_40144,N_39406,N_38572);
and U40145 (N_40145,N_38578,N_38193);
and U40146 (N_40146,N_39315,N_38178);
or U40147 (N_40147,N_38947,N_39950);
and U40148 (N_40148,N_38405,N_38882);
nand U40149 (N_40149,N_39766,N_39680);
nand U40150 (N_40150,N_39273,N_38104);
and U40151 (N_40151,N_38056,N_38165);
nand U40152 (N_40152,N_39330,N_39614);
or U40153 (N_40153,N_38854,N_39184);
nand U40154 (N_40154,N_38859,N_39981);
and U40155 (N_40155,N_39175,N_39363);
and U40156 (N_40156,N_39046,N_38976);
nand U40157 (N_40157,N_38148,N_38810);
xor U40158 (N_40158,N_38906,N_39368);
nand U40159 (N_40159,N_39499,N_38137);
nand U40160 (N_40160,N_39110,N_38665);
nor U40161 (N_40161,N_39726,N_39279);
nor U40162 (N_40162,N_38370,N_39457);
or U40163 (N_40163,N_38184,N_39881);
xnor U40164 (N_40164,N_39039,N_38173);
and U40165 (N_40165,N_38291,N_39503);
nand U40166 (N_40166,N_39643,N_39752);
nor U40167 (N_40167,N_38799,N_39275);
nand U40168 (N_40168,N_38547,N_38830);
or U40169 (N_40169,N_38034,N_39822);
and U40170 (N_40170,N_38986,N_38629);
or U40171 (N_40171,N_39083,N_39091);
and U40172 (N_40172,N_38716,N_39825);
nand U40173 (N_40173,N_38975,N_38885);
or U40174 (N_40174,N_38829,N_38080);
nor U40175 (N_40175,N_38070,N_38853);
nand U40176 (N_40176,N_38670,N_39237);
or U40177 (N_40177,N_39196,N_38465);
xnor U40178 (N_40178,N_38210,N_39498);
and U40179 (N_40179,N_38873,N_38069);
and U40180 (N_40180,N_39801,N_39350);
and U40181 (N_40181,N_39760,N_38890);
nand U40182 (N_40182,N_38642,N_39777);
and U40183 (N_40183,N_39151,N_39021);
or U40184 (N_40184,N_39373,N_38607);
nand U40185 (N_40185,N_38633,N_39153);
nor U40186 (N_40186,N_39136,N_39195);
and U40187 (N_40187,N_39968,N_38811);
and U40188 (N_40188,N_38961,N_39312);
nor U40189 (N_40189,N_38702,N_38063);
or U40190 (N_40190,N_38487,N_39042);
nor U40191 (N_40191,N_39056,N_39174);
nor U40192 (N_40192,N_38602,N_38732);
or U40193 (N_40193,N_39666,N_38368);
or U40194 (N_40194,N_38762,N_39024);
nand U40195 (N_40195,N_39427,N_39018);
nor U40196 (N_40196,N_38560,N_38042);
nor U40197 (N_40197,N_39928,N_38816);
or U40198 (N_40198,N_38806,N_38401);
xor U40199 (N_40199,N_39767,N_38119);
and U40200 (N_40200,N_38525,N_39865);
or U40201 (N_40201,N_38394,N_38599);
nor U40202 (N_40202,N_38481,N_38517);
xnor U40203 (N_40203,N_38377,N_38098);
nor U40204 (N_40204,N_39405,N_39979);
xor U40205 (N_40205,N_39770,N_39484);
or U40206 (N_40206,N_39971,N_38175);
or U40207 (N_40207,N_39649,N_39002);
and U40208 (N_40208,N_39479,N_39099);
xnor U40209 (N_40209,N_38983,N_38736);
nor U40210 (N_40210,N_39329,N_38876);
nand U40211 (N_40211,N_38284,N_38215);
and U40212 (N_40212,N_39134,N_39124);
and U40213 (N_40213,N_39451,N_39840);
nand U40214 (N_40214,N_39308,N_38488);
and U40215 (N_40215,N_39828,N_39633);
and U40216 (N_40216,N_39177,N_39221);
or U40217 (N_40217,N_38079,N_39747);
nor U40218 (N_40218,N_38553,N_38166);
nor U40219 (N_40219,N_38742,N_39488);
or U40220 (N_40220,N_39250,N_39478);
nor U40221 (N_40221,N_39494,N_39845);
nand U40222 (N_40222,N_39022,N_38886);
nand U40223 (N_40223,N_39572,N_38696);
and U40224 (N_40224,N_39837,N_38501);
nand U40225 (N_40225,N_38095,N_39875);
or U40226 (N_40226,N_39112,N_39229);
nor U40227 (N_40227,N_39765,N_39269);
nor U40228 (N_40228,N_38239,N_38335);
or U40229 (N_40229,N_39695,N_39077);
and U40230 (N_40230,N_38760,N_39806);
xnor U40231 (N_40231,N_39270,N_39397);
and U40232 (N_40232,N_39071,N_39879);
and U40233 (N_40233,N_38018,N_38447);
nor U40234 (N_40234,N_38840,N_39526);
or U40235 (N_40235,N_38326,N_38037);
nor U40236 (N_40236,N_39790,N_39035);
nor U40237 (N_40237,N_39973,N_38625);
nand U40238 (N_40238,N_38978,N_38814);
or U40239 (N_40239,N_39988,N_38999);
xor U40240 (N_40240,N_39219,N_38227);
nor U40241 (N_40241,N_38515,N_39718);
xnor U40242 (N_40242,N_38545,N_38655);
nor U40243 (N_40243,N_39059,N_39282);
nor U40244 (N_40244,N_39620,N_38297);
or U40245 (N_40245,N_38005,N_39815);
nand U40246 (N_40246,N_39084,N_38423);
and U40247 (N_40247,N_39735,N_39090);
nand U40248 (N_40248,N_38144,N_39690);
nor U40249 (N_40249,N_38605,N_39824);
and U40250 (N_40250,N_38471,N_39604);
nor U40251 (N_40251,N_38495,N_38248);
or U40252 (N_40252,N_39856,N_39044);
and U40253 (N_40253,N_38867,N_38823);
nand U40254 (N_40254,N_39243,N_39733);
nor U40255 (N_40255,N_39209,N_39437);
or U40256 (N_40256,N_39787,N_38475);
xor U40257 (N_40257,N_39430,N_39390);
nand U40258 (N_40258,N_39528,N_38518);
nor U40259 (N_40259,N_38240,N_39688);
nand U40260 (N_40260,N_39300,N_39259);
nand U40261 (N_40261,N_39459,N_39561);
nand U40262 (N_40262,N_39656,N_39624);
xor U40263 (N_40263,N_39272,N_39412);
and U40264 (N_40264,N_38628,N_38542);
xor U40265 (N_40265,N_38187,N_39205);
or U40266 (N_40266,N_38425,N_39026);
or U40267 (N_40267,N_39383,N_39289);
xnor U40268 (N_40268,N_38073,N_38469);
nand U40269 (N_40269,N_38038,N_38649);
xor U40270 (N_40270,N_39382,N_38891);
nand U40271 (N_40271,N_38298,N_39835);
and U40272 (N_40272,N_39063,N_39720);
or U40273 (N_40273,N_39401,N_38274);
or U40274 (N_40274,N_39518,N_38902);
nor U40275 (N_40275,N_39612,N_39001);
or U40276 (N_40276,N_39408,N_38408);
and U40277 (N_40277,N_39816,N_39118);
or U40278 (N_40278,N_38786,N_39176);
xnor U40279 (N_40279,N_39757,N_38707);
nand U40280 (N_40280,N_39203,N_38903);
nand U40281 (N_40281,N_38780,N_39238);
nand U40282 (N_40282,N_39520,N_38745);
or U40283 (N_40283,N_38314,N_39938);
nor U40284 (N_40284,N_38535,N_38667);
nor U40285 (N_40285,N_38019,N_38110);
or U40286 (N_40286,N_39156,N_38580);
or U40287 (N_40287,N_38172,N_39570);
or U40288 (N_40288,N_38678,N_38463);
nand U40289 (N_40289,N_38251,N_38842);
nor U40290 (N_40290,N_39942,N_38889);
nor U40291 (N_40291,N_39318,N_38281);
nor U40292 (N_40292,N_38724,N_38321);
nand U40293 (N_40293,N_39731,N_38662);
and U40294 (N_40294,N_39653,N_39449);
nor U40295 (N_40295,N_39662,N_39480);
or U40296 (N_40296,N_38895,N_38679);
xnor U40297 (N_40297,N_38960,N_38045);
or U40298 (N_40298,N_39428,N_38815);
and U40299 (N_40299,N_38638,N_38939);
or U40300 (N_40300,N_39780,N_38595);
nand U40301 (N_40301,N_38228,N_38414);
nor U40302 (N_40302,N_39893,N_39951);
xnor U40303 (N_40303,N_38912,N_38221);
nor U40304 (N_40304,N_39355,N_38000);
nand U40305 (N_40305,N_39596,N_38409);
xor U40306 (N_40306,N_39545,N_39671);
and U40307 (N_40307,N_39294,N_38453);
nor U40308 (N_40308,N_39539,N_39303);
or U40309 (N_40309,N_38007,N_39686);
nor U40310 (N_40310,N_38341,N_38196);
xor U40311 (N_40311,N_39222,N_39256);
and U40312 (N_40312,N_39119,N_38156);
or U40313 (N_40313,N_39911,N_38494);
or U40314 (N_40314,N_38054,N_39281);
or U40315 (N_40315,N_39336,N_38684);
and U40316 (N_40316,N_38648,N_39028);
and U40317 (N_40317,N_39771,N_38801);
nand U40318 (N_40318,N_39506,N_38556);
nor U40319 (N_40319,N_39227,N_38872);
xor U40320 (N_40320,N_38439,N_39020);
nand U40321 (N_40321,N_39888,N_39603);
and U40322 (N_40322,N_38315,N_39916);
nor U40323 (N_40323,N_39316,N_39550);
or U40324 (N_40324,N_38935,N_38135);
nor U40325 (N_40325,N_38386,N_39212);
or U40326 (N_40326,N_38552,N_39580);
xnor U40327 (N_40327,N_39030,N_39832);
nand U40328 (N_40328,N_39005,N_39926);
or U40329 (N_40329,N_39636,N_38231);
or U40330 (N_40330,N_39246,N_39400);
nor U40331 (N_40331,N_39869,N_39533);
xor U40332 (N_40332,N_39475,N_39288);
nor U40333 (N_40333,N_39228,N_39080);
or U40334 (N_40334,N_39607,N_38708);
or U40335 (N_40335,N_39960,N_39876);
and U40336 (N_40336,N_38342,N_38874);
nor U40337 (N_40337,N_38654,N_38013);
or U40338 (N_40338,N_39431,N_38290);
nor U40339 (N_40339,N_39854,N_38508);
xnor U40340 (N_40340,N_39525,N_38506);
nand U40341 (N_40341,N_39419,N_38155);
nand U40342 (N_40342,N_39248,N_39681);
nand U40343 (N_40343,N_38850,N_38931);
or U40344 (N_40344,N_39635,N_39578);
nand U40345 (N_40345,N_38855,N_39299);
nor U40346 (N_40346,N_39129,N_38668);
nand U40347 (N_40347,N_39076,N_39340);
and U40348 (N_40348,N_39583,N_39081);
and U40349 (N_40349,N_39804,N_38838);
xor U40350 (N_40350,N_39023,N_38991);
nor U40351 (N_40351,N_39803,N_39337);
xnor U40352 (N_40352,N_39894,N_38851);
xor U40353 (N_40353,N_39168,N_38887);
xor U40354 (N_40354,N_39667,N_38746);
xor U40355 (N_40355,N_39573,N_38520);
nand U40356 (N_40356,N_38958,N_39711);
and U40357 (N_40357,N_38763,N_38834);
or U40358 (N_40358,N_38791,N_38307);
or U40359 (N_40359,N_38821,N_38404);
xnor U40360 (N_40360,N_38726,N_39493);
nand U40361 (N_40361,N_39391,N_39103);
or U40362 (N_40362,N_38082,N_39913);
or U40363 (N_40363,N_39008,N_39619);
and U40364 (N_40364,N_38688,N_39123);
xnor U40365 (N_40365,N_38613,N_38744);
and U40366 (N_40366,N_38219,N_39723);
or U40367 (N_40367,N_38897,N_39160);
nor U40368 (N_40368,N_39461,N_38932);
nor U40369 (N_40369,N_38336,N_38863);
xnor U40370 (N_40370,N_39225,N_39450);
or U40371 (N_40371,N_38626,N_38402);
xnor U40372 (N_40372,N_39516,N_38818);
xnor U40373 (N_40373,N_38254,N_38803);
nor U40374 (N_40374,N_38064,N_39705);
or U40375 (N_40375,N_38881,N_39818);
and U40376 (N_40376,N_38883,N_38624);
nor U40377 (N_40377,N_39904,N_39892);
nand U40378 (N_40378,N_38832,N_38354);
nor U40379 (N_40379,N_39193,N_38612);
and U40380 (N_40380,N_39057,N_38222);
xor U40381 (N_40381,N_38261,N_39795);
nand U40382 (N_40382,N_38406,N_38534);
and U40383 (N_40383,N_38301,N_38039);
nor U40384 (N_40384,N_39293,N_39346);
and U40385 (N_40385,N_38989,N_38693);
nor U40386 (N_40386,N_39433,N_38466);
nand U40387 (N_40387,N_39114,N_38435);
and U40388 (N_40388,N_38646,N_39872);
or U40389 (N_40389,N_39105,N_39632);
nand U40390 (N_40390,N_38743,N_39857);
xnor U40391 (N_40391,N_39096,N_39785);
nor U40392 (N_40392,N_39702,N_38271);
nor U40393 (N_40393,N_38009,N_38948);
nor U40394 (N_40394,N_38907,N_38269);
and U40395 (N_40395,N_38585,N_38250);
xor U40396 (N_40396,N_38705,N_39622);
or U40397 (N_40397,N_39584,N_38794);
nand U40398 (N_40398,N_38031,N_39657);
and U40399 (N_40399,N_39341,N_38440);
nor U40400 (N_40400,N_39884,N_39610);
nand U40401 (N_40401,N_39587,N_39496);
nand U40402 (N_40402,N_38093,N_38457);
or U40403 (N_40403,N_38083,N_39162);
or U40404 (N_40404,N_38524,N_38507);
xor U40405 (N_40405,N_38510,N_39362);
nor U40406 (N_40406,N_39575,N_38709);
xor U40407 (N_40407,N_38216,N_39715);
nor U40408 (N_40408,N_39447,N_39812);
nor U40409 (N_40409,N_38514,N_38127);
nor U40410 (N_40410,N_38164,N_38010);
nand U40411 (N_40411,N_38323,N_38398);
xnor U40412 (N_40412,N_38909,N_38604);
nand U40413 (N_40413,N_38637,N_38687);
nor U40414 (N_40414,N_39751,N_38381);
nand U40415 (N_40415,N_39121,N_39093);
and U40416 (N_40416,N_38061,N_38951);
nor U40417 (N_40417,N_38623,N_38076);
nor U40418 (N_40418,N_39905,N_39055);
nor U40419 (N_40419,N_39232,N_39850);
or U40420 (N_40420,N_39594,N_39356);
xor U40421 (N_40421,N_39199,N_39061);
and U40422 (N_40422,N_39388,N_38160);
xnor U40423 (N_40423,N_39764,N_38387);
nor U40424 (N_40424,N_39164,N_38875);
or U40425 (N_40425,N_39295,N_39567);
nand U40426 (N_40426,N_38692,N_39006);
or U40427 (N_40427,N_38390,N_39552);
xor U40428 (N_40428,N_38358,N_38531);
and U40429 (N_40429,N_38985,N_38017);
nor U40430 (N_40430,N_38836,N_38410);
xnor U40431 (N_40431,N_39509,N_38305);
and U40432 (N_40432,N_38088,N_38478);
nor U40433 (N_40433,N_39531,N_38781);
and U40434 (N_40434,N_39562,N_38739);
xor U40435 (N_40435,N_39863,N_38472);
and U40436 (N_40436,N_38997,N_38299);
and U40437 (N_40437,N_39935,N_39155);
and U40438 (N_40438,N_38120,N_38579);
or U40439 (N_40439,N_38788,N_39417);
nand U40440 (N_40440,N_38896,N_38433);
nor U40441 (N_40441,N_39344,N_38016);
xor U40442 (N_40442,N_39188,N_39639);
and U40443 (N_40443,N_39814,N_38226);
or U40444 (N_40444,N_38140,N_39019);
and U40445 (N_40445,N_39323,N_38711);
nor U40446 (N_40446,N_38246,N_38710);
nor U40447 (N_40447,N_38244,N_38036);
xnor U40448 (N_40448,N_38795,N_39952);
xor U40449 (N_40449,N_38325,N_38455);
nand U40450 (N_40450,N_39609,N_38936);
xnor U40451 (N_40451,N_38028,N_38940);
nor U40452 (N_40452,N_38030,N_38183);
xnor U40453 (N_40453,N_38672,N_38671);
nand U40454 (N_40454,N_39762,N_39053);
nor U40455 (N_40455,N_38610,N_38376);
or U40456 (N_40456,N_38622,N_39626);
xnor U40457 (N_40457,N_38972,N_39152);
and U40458 (N_40458,N_39504,N_38270);
and U40459 (N_40459,N_39946,N_39732);
xnor U40460 (N_40460,N_38530,N_39146);
nor U40461 (N_40461,N_39963,N_38601);
xor U40462 (N_40462,N_38540,N_38770);
xor U40463 (N_40463,N_39236,N_39590);
xor U40464 (N_40464,N_38635,N_39007);
or U40465 (N_40465,N_39178,N_39159);
nand U40466 (N_40466,N_38473,N_39483);
and U40467 (N_40467,N_38666,N_38113);
xnor U40468 (N_40468,N_38797,N_39298);
nor U40469 (N_40469,N_39031,N_38704);
xnor U40470 (N_40470,N_38682,N_39684);
nor U40471 (N_40471,N_38718,N_39703);
and U40472 (N_40472,N_39679,N_38092);
nor U40473 (N_40473,N_38669,N_39782);
and U40474 (N_40474,N_39858,N_39133);
or U40475 (N_40475,N_39352,N_38224);
nand U40476 (N_40476,N_38348,N_39713);
or U40477 (N_40477,N_38130,N_38167);
xor U40478 (N_40478,N_38177,N_38956);
nand U40479 (N_40479,N_39859,N_38391);
or U40480 (N_40480,N_39425,N_39692);
xor U40481 (N_40481,N_39954,N_38919);
and U40482 (N_40482,N_39965,N_38502);
nor U40483 (N_40483,N_39500,N_38369);
nand U40484 (N_40484,N_39640,N_38789);
and U40485 (N_40485,N_39544,N_39868);
nand U40486 (N_40486,N_38725,N_39836);
xnor U40487 (N_40487,N_38057,N_39348);
and U40488 (N_40488,N_38584,N_38608);
nand U40489 (N_40489,N_38674,N_38701);
or U40490 (N_40490,N_38966,N_39834);
nand U40491 (N_40491,N_38118,N_39333);
nor U40492 (N_40492,N_39194,N_38285);
nand U40493 (N_40493,N_38898,N_39805);
nor U40494 (N_40494,N_39320,N_38827);
nor U40495 (N_40495,N_38382,N_38606);
or U40496 (N_40496,N_39908,N_39515);
and U40497 (N_40497,N_39568,N_39452);
nor U40498 (N_40498,N_39549,N_38841);
nand U40499 (N_40499,N_38389,N_39998);
nor U40500 (N_40500,N_39930,N_38157);
or U40501 (N_40501,N_39197,N_39050);
nand U40502 (N_40502,N_38681,N_39698);
nand U40503 (N_40503,N_38700,N_39678);
or U40504 (N_40504,N_39010,N_38990);
or U40505 (N_40505,N_39784,N_39650);
or U40506 (N_40506,N_39943,N_38715);
xnor U40507 (N_40507,N_39485,N_39087);
nand U40508 (N_40508,N_39085,N_39701);
nor U40509 (N_40509,N_38243,N_39239);
nor U40510 (N_40510,N_39783,N_38497);
or U40511 (N_40511,N_39453,N_38197);
nand U40512 (N_40512,N_38758,N_39996);
and U40513 (N_40513,N_39877,N_39456);
nor U40514 (N_40514,N_39411,N_38385);
xnor U40515 (N_40515,N_38154,N_38621);
nor U40516 (N_40516,N_39793,N_39379);
nor U40517 (N_40517,N_38182,N_38287);
or U40518 (N_40518,N_39776,N_38706);
and U40519 (N_40519,N_38383,N_39186);
or U40520 (N_40520,N_39829,N_39510);
and U40521 (N_40521,N_38504,N_39924);
xor U40522 (N_40522,N_38448,N_39041);
xor U40523 (N_40523,N_39455,N_38981);
xor U40524 (N_40524,N_38089,N_38927);
nand U40525 (N_40525,N_38374,N_39613);
and U40526 (N_40526,N_38360,N_39440);
and U40527 (N_40527,N_39553,N_38046);
nor U40528 (N_40528,N_38505,N_39415);
nor U40529 (N_40529,N_38365,N_38320);
and U40530 (N_40530,N_38121,N_38749);
nor U40531 (N_40531,N_38139,N_39842);
xor U40532 (N_40532,N_38812,N_38349);
nand U40533 (N_40533,N_38955,N_39403);
or U40534 (N_40534,N_39676,N_38316);
or U40535 (N_40535,N_38040,N_38002);
and U40536 (N_40536,N_38430,N_39629);
xor U40537 (N_40537,N_39003,N_38852);
or U40538 (N_40538,N_39773,N_38793);
and U40539 (N_40539,N_39966,N_39149);
or U40540 (N_40540,N_38776,N_38286);
nand U40541 (N_40541,N_38432,N_38442);
xnor U40542 (N_40542,N_38549,N_38878);
xor U40543 (N_40543,N_38004,N_39883);
xor U40544 (N_40544,N_38361,N_38790);
and U40545 (N_40545,N_39245,N_38262);
xor U40546 (N_40546,N_38569,N_39170);
xnor U40547 (N_40547,N_39223,N_38825);
and U40548 (N_40548,N_39342,N_38209);
nand U40549 (N_40549,N_39418,N_39148);
xor U40550 (N_40550,N_38304,N_39290);
and U40551 (N_40551,N_38523,N_39873);
or U40552 (N_40552,N_39069,N_39861);
and U40553 (N_40553,N_39975,N_39953);
nand U40554 (N_40554,N_38544,N_39592);
xor U40555 (N_40555,N_38680,N_38921);
nand U40556 (N_40556,N_39669,N_38899);
or U40557 (N_40557,N_38639,N_39983);
and U40558 (N_40558,N_39477,N_39833);
or U40559 (N_40559,N_38731,N_38967);
and U40560 (N_40560,N_38598,N_38415);
or U40561 (N_40561,N_39693,N_38212);
nand U40562 (N_40562,N_39588,N_38573);
nor U40563 (N_40563,N_39541,N_38048);
nand U40564 (N_40564,N_39328,N_38289);
and U40565 (N_40565,N_38117,N_38831);
nand U40566 (N_40566,N_39384,N_39722);
xor U40567 (N_40567,N_39606,N_38620);
or U40568 (N_40568,N_38533,N_39345);
nand U40569 (N_40569,N_39252,N_38392);
nor U40570 (N_40570,N_38820,N_38973);
or U40571 (N_40571,N_39617,N_39661);
nand U40572 (N_40572,N_38737,N_38283);
or U40573 (N_40573,N_38199,N_39674);
xnor U40574 (N_40574,N_39589,N_39231);
nor U40575 (N_40575,N_38566,N_39310);
nor U40576 (N_40576,N_39347,N_39491);
and U40577 (N_40577,N_39127,N_38047);
nand U40578 (N_40578,N_38631,N_38597);
or U40579 (N_40579,N_38179,N_39637);
xor U40580 (N_40580,N_39585,N_39934);
or U40581 (N_40581,N_39278,N_39774);
nor U40582 (N_40582,N_39563,N_38869);
nor U40583 (N_40583,N_38630,N_39848);
or U40584 (N_40584,N_38914,N_38980);
nor U40585 (N_40585,N_39595,N_39746);
nor U40586 (N_40586,N_39673,N_39754);
nor U40587 (N_40587,N_39173,N_39423);
nand U40588 (N_40588,N_39933,N_39665);
or U40589 (N_40589,N_38094,N_39560);
nand U40590 (N_40590,N_38686,N_39991);
xnor U40591 (N_40591,N_38399,N_39254);
nand U40592 (N_40592,N_39738,N_39187);
xor U40593 (N_40593,N_39396,N_39458);
nand U40594 (N_40594,N_38615,N_38905);
xnor U40595 (N_40595,N_38950,N_39986);
or U40596 (N_40596,N_38265,N_38923);
xor U40597 (N_40597,N_39623,N_39032);
nand U40598 (N_40598,N_39659,N_38191);
and U40599 (N_40599,N_39257,N_39642);
and U40600 (N_40600,N_39839,N_38288);
xnor U40601 (N_40601,N_39796,N_39432);
nand U40602 (N_40602,N_39190,N_39486);
nor U40603 (N_40603,N_39495,N_39652);
nor U40604 (N_40604,N_38782,N_39380);
nand U40605 (N_40605,N_38436,N_38129);
nand U40606 (N_40606,N_39864,N_38930);
or U40607 (N_40607,N_38168,N_39395);
xnor U40608 (N_40608,N_38647,N_38162);
or U40609 (N_40609,N_38468,N_39078);
nand U40610 (N_40610,N_38954,N_39241);
nand U40611 (N_40611,N_39709,N_38856);
or U40612 (N_40612,N_39800,N_38835);
nand U40613 (N_40613,N_38043,N_38768);
xor U40614 (N_40614,N_38249,N_39420);
nor U40615 (N_40615,N_39936,N_39216);
xor U40616 (N_40616,N_39017,N_38362);
and U40617 (N_40617,N_39945,N_39577);
xnor U40618 (N_40618,N_39712,N_39327);
or U40619 (N_40619,N_38787,N_39376);
nand U40620 (N_40620,N_39529,N_39375);
nand U40621 (N_40621,N_39885,N_39683);
and U40622 (N_40622,N_39630,N_39139);
or U40623 (N_40623,N_39901,N_39849);
or U40624 (N_40624,N_39534,N_39307);
nand U40625 (N_40625,N_39100,N_39062);
nor U40626 (N_40626,N_39378,N_39106);
nand U40627 (N_40627,N_38528,N_38945);
or U40628 (N_40628,N_39882,N_39536);
nand U40629 (N_40629,N_39931,N_39753);
nand U40630 (N_40630,N_39993,N_39109);
nor U40631 (N_40631,N_39862,N_38395);
and U40632 (N_40632,N_39734,N_38683);
or U40633 (N_40633,N_39233,N_38467);
nand U40634 (N_40634,N_38310,N_39948);
or U40635 (N_40635,N_39366,N_38188);
or U40636 (N_40636,N_39215,N_39150);
xnor U40637 (N_40637,N_38116,N_38957);
nand U40638 (N_40638,N_39571,N_38963);
nor U40639 (N_40639,N_39354,N_38152);
xnor U40640 (N_40640,N_38499,N_39940);
nor U40641 (N_40641,N_39258,N_38952);
nor U40642 (N_40642,N_39291,N_38169);
nor U40643 (N_40643,N_39092,N_39523);
or U40644 (N_40644,N_38928,N_38345);
nand U40645 (N_40645,N_39557,N_38483);
or U40646 (N_40646,N_38022,N_38796);
and U40647 (N_40647,N_38084,N_39064);
nand U40648 (N_40648,N_39260,N_39144);
nor U40649 (N_40649,N_39909,N_39036);
xnor U40650 (N_40650,N_38238,N_38086);
xor U40651 (N_40651,N_38035,N_39165);
and U40652 (N_40652,N_39369,N_38450);
xnor U40653 (N_40653,N_38021,N_38754);
nand U40654 (N_40654,N_39999,N_38159);
nor U40655 (N_40655,N_38142,N_39004);
xnor U40656 (N_40656,N_38033,N_39407);
and U40657 (N_40657,N_39306,N_39505);
and U40658 (N_40658,N_38652,N_38777);
or U40659 (N_40659,N_38006,N_38107);
or U40660 (N_40660,N_38860,N_39255);
or U40661 (N_40661,N_39169,N_38115);
nand U40662 (N_40662,N_38186,N_39517);
or U40663 (N_40663,N_38847,N_38201);
and U40664 (N_40664,N_38074,N_38809);
or U40665 (N_40665,N_39616,N_38068);
nand U40666 (N_40666,N_39335,N_38011);
xor U40667 (N_40667,N_39370,N_38388);
and U40668 (N_40668,N_38833,N_38311);
xor U40669 (N_40669,N_39558,N_38942);
nand U40670 (N_40670,N_38880,N_38328);
nor U40671 (N_40671,N_39817,N_38632);
and U40672 (N_40672,N_38241,N_39161);
or U40673 (N_40673,N_39179,N_38675);
nand U40674 (N_40674,N_39235,N_39421);
xnor U40675 (N_40675,N_39758,N_38730);
xor U40676 (N_40676,N_38081,N_39670);
nand U40677 (N_40677,N_39313,N_38203);
or U40678 (N_40678,N_39874,N_38970);
and U40679 (N_40679,N_38915,N_38161);
nor U40680 (N_40680,N_39094,N_38839);
or U40681 (N_40681,N_39540,N_38493);
and U40682 (N_40682,N_39000,N_38996);
nor U40683 (N_40683,N_39602,N_39353);
or U40684 (N_40684,N_39074,N_39454);
and U40685 (N_40685,N_38857,N_39434);
xor U40686 (N_40686,N_38208,N_39939);
nor U40687 (N_40687,N_38486,N_38918);
nor U40688 (N_40688,N_38901,N_38373);
nand U40689 (N_40689,N_38920,N_39830);
nor U40690 (N_40690,N_38766,N_39217);
nor U40691 (N_40691,N_39460,N_38703);
and U40692 (N_40692,N_38543,N_39647);
and U40693 (N_40693,N_39967,N_38609);
nor U40694 (N_40694,N_39645,N_39900);
and U40695 (N_40695,N_38656,N_39206);
and U40696 (N_40696,N_39191,N_38114);
nand U40697 (N_40697,N_39204,N_38071);
nand U40698 (N_40698,N_39956,N_39961);
or U40699 (N_40699,N_39779,N_39073);
nor U40700 (N_40700,N_38712,N_39870);
and U40701 (N_40701,N_38090,N_39772);
nand U40702 (N_40702,N_39332,N_38987);
and U40703 (N_40703,N_39438,N_38229);
xor U40704 (N_40704,N_39297,N_39867);
or U40705 (N_40705,N_39244,N_39399);
and U40706 (N_40706,N_38275,N_38300);
or U40707 (N_40707,N_38330,N_39627);
nor U40708 (N_40708,N_39687,N_39441);
xor U40709 (N_40709,N_38618,N_39304);
xor U40710 (N_40710,N_39807,N_39422);
and U40711 (N_40711,N_38470,N_39338);
xor U40712 (N_40712,N_39424,N_39325);
nand U40713 (N_40713,N_38419,N_39439);
or U40714 (N_40714,N_38233,N_38979);
xor U40715 (N_40715,N_38521,N_39794);
and U40716 (N_40716,N_39122,N_38677);
nor U40717 (N_40717,N_39251,N_39435);
xnor U40718 (N_40718,N_38317,N_39708);
xnor U40719 (N_40719,N_39741,N_38527);
xor U40720 (N_40720,N_39240,N_39466);
xor U40721 (N_40721,N_39628,N_38147);
or U40722 (N_40722,N_39167,N_38202);
nor U40723 (N_40723,N_38586,N_39658);
xnor U40724 (N_40724,N_39116,N_38407);
nand U40725 (N_40725,N_39359,N_39844);
nand U40726 (N_40726,N_39198,N_39462);
nand U40727 (N_40727,N_38366,N_39402);
nand U40728 (N_40728,N_38422,N_38456);
xnor U40729 (N_40729,N_38170,N_38537);
nor U40730 (N_40730,N_38461,N_39891);
xor U40731 (N_40731,N_38367,N_38072);
nor U40732 (N_40732,N_38112,N_38128);
xor U40733 (N_40733,N_38462,N_39664);
and U40734 (N_40734,N_39985,N_38372);
xor U40735 (N_40735,N_38085,N_38444);
nand U40736 (N_40736,N_39490,N_38519);
and U40737 (N_40737,N_38252,N_38218);
xor U40738 (N_40738,N_38053,N_38772);
or U40739 (N_40739,N_38884,N_38282);
xor U40740 (N_40740,N_39638,N_38953);
or U40741 (N_40741,N_38424,N_38611);
nor U40742 (N_40742,N_39959,N_39016);
or U40743 (N_40743,N_39895,N_39097);
nand U40744 (N_40744,N_38146,N_39374);
and U40745 (N_40745,N_38096,N_39866);
and U40746 (N_40746,N_39564,N_39660);
or U40747 (N_40747,N_39266,N_38848);
or U40748 (N_40748,N_38837,N_39932);
and U40749 (N_40749,N_38378,N_38242);
nand U40750 (N_40750,N_39088,N_38332);
and U40751 (N_40751,N_38213,N_38783);
nor U40752 (N_40752,N_38864,N_39740);
nand U40753 (N_40753,N_39808,N_39871);
xnor U40754 (N_40754,N_39343,N_39095);
or U40755 (N_40755,N_38691,N_38995);
nand U40756 (N_40756,N_38593,N_39763);
nor U40757 (N_40757,N_38769,N_38272);
and U40758 (N_40758,N_39565,N_39267);
and U40759 (N_40759,N_39463,N_38634);
or U40760 (N_40760,N_39880,N_39101);
nand U40761 (N_40761,N_38589,N_39813);
nand U40762 (N_40762,N_39569,N_38206);
xnor U40763 (N_40763,N_38567,N_39242);
or U40764 (N_40764,N_39261,N_39737);
nand U40765 (N_40765,N_39990,N_38302);
nor U40766 (N_40766,N_38733,N_38012);
nand U40767 (N_40767,N_38843,N_38449);
and U40768 (N_40768,N_38650,N_38171);
or U40769 (N_40769,N_39689,N_39361);
xor U40770 (N_40770,N_38937,N_39296);
and U40771 (N_40771,N_38636,N_38779);
nand U40772 (N_40772,N_38459,N_39086);
nand U40773 (N_40773,N_38614,N_39113);
nand U40774 (N_40774,N_38663,N_39387);
nor U40775 (N_40775,N_39574,N_39487);
or U40776 (N_40776,N_39200,N_38189);
nor U40777 (N_40777,N_39997,N_38603);
nor U40778 (N_40778,N_39947,N_39593);
nor U40779 (N_40779,N_38411,N_39287);
xnor U40780 (N_40780,N_38032,N_38111);
xnor U40781 (N_40781,N_39791,N_39166);
xor U40782 (N_40782,N_38429,N_38334);
or U40783 (N_40783,N_39524,N_38204);
or U40784 (N_40784,N_39443,N_39052);
nor U40785 (N_40785,N_38101,N_38055);
xor U40786 (N_40786,N_39974,N_38645);
nand U40787 (N_40787,N_38044,N_38338);
or U40788 (N_40788,N_38428,N_39066);
nor U40789 (N_40789,N_39739,N_38363);
and U40790 (N_40790,N_38802,N_39512);
nor U40791 (N_40791,N_38561,N_38319);
or U40792 (N_40792,N_39446,N_39918);
xor U40793 (N_40793,N_39321,N_38893);
and U40794 (N_40794,N_39756,N_39108);
nand U40795 (N_40795,N_39492,N_39989);
and U40796 (N_40796,N_38454,N_39896);
xor U40797 (N_40797,N_39915,N_38023);
and U40798 (N_40798,N_38078,N_39147);
xor U40799 (N_40799,N_39416,N_39015);
and U40800 (N_40800,N_38277,N_38234);
and U40801 (N_40801,N_38198,N_39852);
xnor U40802 (N_40802,N_38596,N_38879);
nand U40803 (N_40803,N_38134,N_38150);
xor U40804 (N_40804,N_38318,N_39706);
or U40805 (N_40805,N_39476,N_39102);
nor U40806 (N_40806,N_38295,N_39264);
nand U40807 (N_40807,N_39597,N_39634);
nor U40808 (N_40808,N_38858,N_38757);
and U40809 (N_40809,N_39677,N_39730);
nand U40810 (N_40810,N_38962,N_38393);
nor U40811 (N_40811,N_39214,N_39700);
or U40812 (N_40812,N_39743,N_39887);
xnor U40813 (N_40813,N_39115,N_38491);
and U40814 (N_40814,N_38546,N_38484);
nor U40815 (N_40815,N_39811,N_39685);
nand U40816 (N_40816,N_38738,N_38752);
nand U40817 (N_40817,N_38695,N_38805);
nor U40818 (N_40818,N_38659,N_38949);
xnor U40819 (N_40819,N_38356,N_38051);
nand U40820 (N_40820,N_39364,N_39742);
nor U40821 (N_40821,N_38126,N_38180);
or U40822 (N_40822,N_39181,N_38938);
nand U40823 (N_40823,N_38477,N_38108);
or U40824 (N_40824,N_38888,N_39566);
or U40825 (N_40825,N_38253,N_38861);
or U40826 (N_40826,N_39301,N_39305);
nor U40827 (N_40827,N_39519,N_38200);
or U40828 (N_40828,N_39919,N_39051);
and U40829 (N_40829,N_39644,N_39768);
and U40830 (N_40830,N_38279,N_39792);
nor U40831 (N_40831,N_38427,N_39699);
nand U40832 (N_40832,N_38562,N_38600);
and U40833 (N_40833,N_38176,N_39704);
and U40834 (N_40834,N_39527,N_38728);
xnor U40835 (N_40835,N_38824,N_39208);
nand U40836 (N_40836,N_38946,N_39481);
or U40837 (N_40837,N_39992,N_39157);
or U40838 (N_40838,N_39672,N_39040);
or U40839 (N_40839,N_39220,N_39682);
or U40840 (N_40840,N_38563,N_38132);
nor U40841 (N_40841,N_39977,N_38024);
nand U40842 (N_40842,N_38778,N_39033);
xor U40843 (N_40843,N_38194,N_38564);
xor U40844 (N_40844,N_39060,N_38255);
nor U40845 (N_40845,N_38452,N_38397);
nor U40846 (N_40846,N_38916,N_38559);
or U40847 (N_40847,N_38306,N_38103);
nor U40848 (N_40848,N_38151,N_38445);
nor U40849 (N_40849,N_38804,N_38237);
or U40850 (N_40850,N_39889,N_38565);
or U40851 (N_40851,N_39853,N_38364);
xnor U40852 (N_40852,N_38773,N_39788);
xnor U40853 (N_40853,N_38412,N_38551);
nand U40854 (N_40854,N_38969,N_38994);
xnor U40855 (N_40855,N_38813,N_39608);
nand U40856 (N_40856,N_38617,N_39381);
nand U40857 (N_40857,N_39984,N_38570);
nand U40858 (N_40858,N_39280,N_38959);
or U40859 (N_40859,N_39314,N_39436);
xor U40860 (N_40860,N_38846,N_39914);
or U40861 (N_40861,N_38324,N_38699);
or U40862 (N_40862,N_39322,N_39029);
nand U40863 (N_40863,N_39470,N_39158);
nor U40864 (N_40864,N_38280,N_39183);
nor U40865 (N_40865,N_39472,N_39957);
nand U40866 (N_40866,N_39736,N_39048);
or U40867 (N_40867,N_39286,N_39897);
xor U40868 (N_40868,N_38735,N_39600);
or U40869 (N_40869,N_39559,N_38558);
nor U40870 (N_40870,N_39474,N_39172);
and U40871 (N_40871,N_39721,N_38529);
or U40872 (N_40872,N_39182,N_38964);
or U40873 (N_40873,N_38257,N_39398);
or U40874 (N_40874,N_39180,N_39226);
nand U40875 (N_40875,N_38581,N_38690);
and U40876 (N_40876,N_38100,N_39276);
or U40877 (N_40877,N_38866,N_39043);
xnor U40878 (N_40878,N_38065,N_39823);
nor U40879 (N_40879,N_38431,N_38643);
xnor U40880 (N_40880,N_39972,N_39786);
and U40881 (N_40881,N_39555,N_39185);
nor U40882 (N_40882,N_39537,N_38163);
or U40883 (N_40883,N_39710,N_38245);
or U40884 (N_40884,N_38357,N_39641);
xor U40885 (N_40885,N_39941,N_38421);
and U40886 (N_40886,N_39831,N_39556);
nor U40887 (N_40887,N_38574,N_39465);
xor U40888 (N_40888,N_39759,N_39442);
nand U40889 (N_40889,N_38359,N_39899);
nand U40890 (N_40890,N_38211,N_39922);
xor U40891 (N_40891,N_39207,N_39797);
or U40892 (N_40892,N_38124,N_38673);
nor U40893 (N_40893,N_38443,N_38616);
nor U40894 (N_40894,N_39247,N_39027);
xor U40895 (N_40895,N_38498,N_39067);
nand U40896 (N_40896,N_39507,N_39192);
or U40897 (N_40897,N_38438,N_38276);
nor U40898 (N_40898,N_39691,N_38594);
and U40899 (N_40899,N_39075,N_39351);
and U40900 (N_40900,N_38539,N_39511);
and U40901 (N_40901,N_38136,N_38503);
nand U40902 (N_40902,N_39125,N_39906);
nand U40903 (N_40903,N_38014,N_38849);
nor U40904 (N_40904,N_39386,N_38808);
xor U40905 (N_40905,N_38026,N_39089);
or U40906 (N_40906,N_39755,N_38845);
or U40907 (N_40907,N_38339,N_38714);
xnor U40908 (N_40908,N_38476,N_39744);
xnor U40909 (N_40909,N_39535,N_39949);
or U40910 (N_40910,N_38661,N_38403);
or U40911 (N_40911,N_38500,N_38511);
nor U40912 (N_40912,N_38087,N_38075);
nand U40913 (N_40913,N_38713,N_39907);
nand U40914 (N_40914,N_38418,N_38761);
nand U40915 (N_40915,N_39598,N_38097);
nand U40916 (N_40916,N_39210,N_39955);
xor U40917 (N_40917,N_38557,N_39265);
nand U40918 (N_40918,N_38698,N_39717);
and U40919 (N_40919,N_39393,N_39962);
xor U40920 (N_40920,N_39576,N_39409);
nand U40921 (N_40921,N_38755,N_39976);
or U40922 (N_40922,N_39249,N_38741);
nand U40923 (N_40923,N_38067,N_39334);
or U40924 (N_40924,N_38792,N_39426);
nor U40925 (N_40925,N_38892,N_39925);
nand U40926 (N_40926,N_38697,N_38993);
or U40927 (N_40927,N_38400,N_38145);
nand U40928 (N_40928,N_38417,N_38819);
or U40929 (N_40929,N_38548,N_39554);
nand U40930 (N_40930,N_39404,N_39034);
and U40931 (N_40931,N_38205,N_39189);
nor U40932 (N_40932,N_39038,N_38236);
nor U40933 (N_40933,N_38568,N_38785);
xor U40934 (N_40934,N_38351,N_39358);
or U40935 (N_40935,N_38375,N_38225);
or U40936 (N_40936,N_39065,N_39532);
xnor U40937 (N_40937,N_38720,N_38913);
nor U40938 (N_40938,N_38296,N_38619);
and U40939 (N_40939,N_39292,N_39445);
xor U40940 (N_40940,N_39860,N_38327);
nand U40941 (N_40941,N_38260,N_39502);
and U40942 (N_40942,N_38933,N_39631);
xnor U40943 (N_40943,N_38267,N_39011);
nand U40944 (N_40944,N_39464,N_38451);
nand U40945 (N_40945,N_39655,N_38313);
and U40946 (N_40946,N_38719,N_38413);
or U40947 (N_40947,N_38293,N_39920);
nand U40948 (N_40948,N_39581,N_38312);
nor U40949 (N_40949,N_38865,N_38653);
nor U40950 (N_40950,N_38583,N_39781);
xnor U40951 (N_40951,N_39958,N_39365);
nor U40952 (N_40952,N_38664,N_38337);
xnor U40953 (N_40953,N_39012,N_38784);
xor U40954 (N_40954,N_39171,N_39995);
and U40955 (N_40955,N_39072,N_38379);
and U40956 (N_40956,N_38102,N_38066);
or U40957 (N_40957,N_39132,N_39546);
nand U40958 (N_40958,N_38509,N_38641);
and U40959 (N_40959,N_38185,N_39521);
nor U40960 (N_40960,N_39724,N_38258);
nor U40961 (N_40961,N_39224,N_38485);
xor U40962 (N_40962,N_38223,N_39410);
nor U40963 (N_40963,N_38153,N_39058);
or U40964 (N_40964,N_38894,N_39014);
xor U40965 (N_40965,N_39978,N_39725);
nor U40966 (N_40966,N_39154,N_39234);
xnor U40967 (N_40967,N_39360,N_39497);
nand U40968 (N_40968,N_39319,N_39675);
xor U40969 (N_40969,N_39745,N_38029);
xor U40970 (N_40970,N_38105,N_39838);
xor U40971 (N_40971,N_38174,N_39599);
nand U40972 (N_40972,N_38862,N_39274);
and U40973 (N_40973,N_39429,N_39846);
and U40974 (N_40974,N_38125,N_39646);
and U40975 (N_40975,N_39218,N_38380);
nor U40976 (N_40976,N_38192,N_38058);
or U40977 (N_40977,N_39271,N_38437);
nor U40978 (N_40978,N_39054,N_38871);
or U40979 (N_40979,N_38627,N_39211);
nor U40980 (N_40980,N_38753,N_38729);
and U40981 (N_40981,N_38844,N_38217);
nor U40982 (N_40982,N_39253,N_39049);
xnor U40983 (N_40983,N_39473,N_38910);
or U40984 (N_40984,N_38292,N_39809);
or U40985 (N_40985,N_39778,N_38532);
and U40986 (N_40986,N_38256,N_38748);
nor U40987 (N_40987,N_39268,N_39501);
and U40988 (N_40988,N_39841,N_38751);
xnor U40989 (N_40989,N_39586,N_39098);
nand U40990 (N_40990,N_38765,N_38268);
or U40991 (N_40991,N_39394,N_38181);
and U40992 (N_40992,N_39142,N_39128);
nor U40993 (N_40993,N_38941,N_38003);
nand U40994 (N_40994,N_39615,N_38109);
nor U40995 (N_40995,N_38062,N_38590);
xnor U40996 (N_40996,N_38474,N_39750);
nand U40997 (N_40997,N_38460,N_39898);
and U40998 (N_40998,N_38131,N_39929);
or U40999 (N_40999,N_39263,N_38694);
xnor U41000 (N_41000,N_38474,N_38927);
nor U41001 (N_41001,N_39321,N_38422);
xor U41002 (N_41002,N_38160,N_39779);
nand U41003 (N_41003,N_39724,N_38381);
nand U41004 (N_41004,N_39960,N_38300);
and U41005 (N_41005,N_39676,N_39599);
nand U41006 (N_41006,N_39626,N_38002);
nor U41007 (N_41007,N_39458,N_38585);
nand U41008 (N_41008,N_38491,N_39951);
xnor U41009 (N_41009,N_38197,N_38146);
xor U41010 (N_41010,N_38363,N_39899);
xnor U41011 (N_41011,N_38997,N_38340);
nor U41012 (N_41012,N_39228,N_39744);
nor U41013 (N_41013,N_38992,N_39544);
and U41014 (N_41014,N_38577,N_39788);
or U41015 (N_41015,N_38503,N_39433);
nand U41016 (N_41016,N_39746,N_39196);
and U41017 (N_41017,N_39028,N_38558);
xor U41018 (N_41018,N_38903,N_38486);
xnor U41019 (N_41019,N_38527,N_38742);
or U41020 (N_41020,N_38562,N_38570);
nand U41021 (N_41021,N_38142,N_39575);
xor U41022 (N_41022,N_38908,N_38521);
or U41023 (N_41023,N_38445,N_38699);
nand U41024 (N_41024,N_39787,N_38638);
or U41025 (N_41025,N_39528,N_39859);
or U41026 (N_41026,N_38103,N_38948);
and U41027 (N_41027,N_39132,N_38609);
nand U41028 (N_41028,N_38993,N_39816);
nand U41029 (N_41029,N_39281,N_38340);
nand U41030 (N_41030,N_38189,N_39324);
xnor U41031 (N_41031,N_39928,N_39867);
nand U41032 (N_41032,N_38375,N_38870);
nand U41033 (N_41033,N_38790,N_39860);
nor U41034 (N_41034,N_39292,N_38651);
nor U41035 (N_41035,N_38757,N_38804);
xor U41036 (N_41036,N_39825,N_39756);
nand U41037 (N_41037,N_39514,N_39420);
and U41038 (N_41038,N_39690,N_39940);
xor U41039 (N_41039,N_38689,N_38328);
and U41040 (N_41040,N_39466,N_38273);
xnor U41041 (N_41041,N_38245,N_39634);
nand U41042 (N_41042,N_39367,N_39324);
and U41043 (N_41043,N_38295,N_38043);
and U41044 (N_41044,N_39325,N_39888);
nand U41045 (N_41045,N_38572,N_38141);
and U41046 (N_41046,N_38603,N_39270);
nand U41047 (N_41047,N_39711,N_38831);
or U41048 (N_41048,N_39688,N_38398);
nor U41049 (N_41049,N_38067,N_38828);
nor U41050 (N_41050,N_39393,N_39528);
xnor U41051 (N_41051,N_38861,N_38118);
nor U41052 (N_41052,N_39749,N_39183);
xor U41053 (N_41053,N_38640,N_39094);
and U41054 (N_41054,N_38871,N_38997);
nor U41055 (N_41055,N_39755,N_39445);
nor U41056 (N_41056,N_39647,N_39572);
and U41057 (N_41057,N_39422,N_38708);
or U41058 (N_41058,N_39306,N_38821);
and U41059 (N_41059,N_39549,N_39898);
nand U41060 (N_41060,N_39250,N_38178);
and U41061 (N_41061,N_38405,N_38473);
and U41062 (N_41062,N_39938,N_39029);
and U41063 (N_41063,N_39626,N_38809);
nand U41064 (N_41064,N_38346,N_38608);
nor U41065 (N_41065,N_38993,N_38282);
nand U41066 (N_41066,N_38272,N_39645);
nor U41067 (N_41067,N_38637,N_38997);
xor U41068 (N_41068,N_38287,N_39632);
or U41069 (N_41069,N_38915,N_38830);
nand U41070 (N_41070,N_39464,N_39634);
or U41071 (N_41071,N_38506,N_38903);
and U41072 (N_41072,N_39982,N_39683);
nor U41073 (N_41073,N_38706,N_38556);
and U41074 (N_41074,N_38004,N_38208);
nor U41075 (N_41075,N_38890,N_39303);
xnor U41076 (N_41076,N_38437,N_39584);
and U41077 (N_41077,N_39310,N_39703);
xor U41078 (N_41078,N_39116,N_39342);
or U41079 (N_41079,N_39851,N_38576);
and U41080 (N_41080,N_39190,N_39576);
or U41081 (N_41081,N_39556,N_39080);
xnor U41082 (N_41082,N_38373,N_38981);
nand U41083 (N_41083,N_39696,N_38005);
xor U41084 (N_41084,N_39781,N_38517);
xor U41085 (N_41085,N_38105,N_39009);
and U41086 (N_41086,N_39602,N_38676);
nand U41087 (N_41087,N_39703,N_39785);
and U41088 (N_41088,N_39744,N_38248);
nor U41089 (N_41089,N_39287,N_39739);
or U41090 (N_41090,N_39155,N_39972);
xor U41091 (N_41091,N_38881,N_39463);
nor U41092 (N_41092,N_39828,N_38529);
and U41093 (N_41093,N_39492,N_39781);
xor U41094 (N_41094,N_39983,N_39212);
xnor U41095 (N_41095,N_39778,N_38681);
xor U41096 (N_41096,N_38140,N_39048);
xor U41097 (N_41097,N_39550,N_39891);
nor U41098 (N_41098,N_39578,N_38320);
nand U41099 (N_41099,N_38034,N_38350);
or U41100 (N_41100,N_39479,N_38982);
and U41101 (N_41101,N_38910,N_39602);
nand U41102 (N_41102,N_39846,N_38499);
nand U41103 (N_41103,N_38939,N_39914);
and U41104 (N_41104,N_39102,N_38457);
nand U41105 (N_41105,N_39775,N_38287);
xor U41106 (N_41106,N_39697,N_38530);
and U41107 (N_41107,N_38346,N_39203);
and U41108 (N_41108,N_38141,N_38105);
or U41109 (N_41109,N_38435,N_39850);
or U41110 (N_41110,N_38703,N_39349);
nand U41111 (N_41111,N_39180,N_38517);
or U41112 (N_41112,N_39850,N_39727);
nand U41113 (N_41113,N_39020,N_38769);
xor U41114 (N_41114,N_39221,N_39867);
or U41115 (N_41115,N_38686,N_39193);
and U41116 (N_41116,N_38716,N_39446);
nand U41117 (N_41117,N_38646,N_39071);
xnor U41118 (N_41118,N_39242,N_39317);
nor U41119 (N_41119,N_39900,N_39297);
and U41120 (N_41120,N_39718,N_39205);
nand U41121 (N_41121,N_39599,N_38189);
nand U41122 (N_41122,N_39167,N_38661);
nand U41123 (N_41123,N_38576,N_39323);
nor U41124 (N_41124,N_38324,N_38537);
nand U41125 (N_41125,N_39838,N_39034);
xor U41126 (N_41126,N_38908,N_38448);
or U41127 (N_41127,N_38899,N_38377);
nand U41128 (N_41128,N_38256,N_39565);
nand U41129 (N_41129,N_39579,N_39656);
and U41130 (N_41130,N_39100,N_38928);
nor U41131 (N_41131,N_39042,N_39905);
or U41132 (N_41132,N_39570,N_39761);
or U41133 (N_41133,N_39975,N_39739);
nor U41134 (N_41134,N_38506,N_38571);
xnor U41135 (N_41135,N_39278,N_39226);
xor U41136 (N_41136,N_39506,N_39261);
nand U41137 (N_41137,N_38159,N_39711);
xnor U41138 (N_41138,N_38286,N_39407);
or U41139 (N_41139,N_38402,N_39788);
nand U41140 (N_41140,N_39097,N_39592);
or U41141 (N_41141,N_39193,N_38021);
or U41142 (N_41142,N_39210,N_38911);
or U41143 (N_41143,N_38254,N_39562);
or U41144 (N_41144,N_38951,N_38226);
nor U41145 (N_41145,N_38074,N_39918);
and U41146 (N_41146,N_38273,N_38994);
and U41147 (N_41147,N_38862,N_39268);
or U41148 (N_41148,N_38218,N_38485);
or U41149 (N_41149,N_38116,N_39807);
nand U41150 (N_41150,N_39240,N_39898);
nand U41151 (N_41151,N_38103,N_39024);
and U41152 (N_41152,N_39413,N_39857);
or U41153 (N_41153,N_39820,N_39542);
nand U41154 (N_41154,N_38831,N_39788);
nand U41155 (N_41155,N_38005,N_38935);
nand U41156 (N_41156,N_39367,N_38101);
nand U41157 (N_41157,N_39563,N_39070);
xnor U41158 (N_41158,N_38627,N_39450);
xnor U41159 (N_41159,N_39443,N_38471);
nor U41160 (N_41160,N_39491,N_39560);
or U41161 (N_41161,N_38163,N_39826);
and U41162 (N_41162,N_39629,N_38333);
and U41163 (N_41163,N_39303,N_39650);
xor U41164 (N_41164,N_39705,N_39004);
and U41165 (N_41165,N_38221,N_39806);
nor U41166 (N_41166,N_39767,N_39091);
or U41167 (N_41167,N_39595,N_39968);
nand U41168 (N_41168,N_39941,N_38651);
and U41169 (N_41169,N_38137,N_39204);
nand U41170 (N_41170,N_38178,N_38744);
nor U41171 (N_41171,N_39723,N_39182);
and U41172 (N_41172,N_39020,N_38324);
nor U41173 (N_41173,N_38386,N_39242);
nor U41174 (N_41174,N_39810,N_39342);
nand U41175 (N_41175,N_38184,N_38089);
nor U41176 (N_41176,N_38214,N_38687);
nand U41177 (N_41177,N_38939,N_38733);
xor U41178 (N_41178,N_39851,N_39162);
or U41179 (N_41179,N_38686,N_38059);
nand U41180 (N_41180,N_39208,N_38430);
xor U41181 (N_41181,N_39033,N_38734);
nor U41182 (N_41182,N_38180,N_39711);
and U41183 (N_41183,N_38389,N_38687);
and U41184 (N_41184,N_39633,N_39258);
nor U41185 (N_41185,N_38835,N_39652);
nand U41186 (N_41186,N_39902,N_39465);
xnor U41187 (N_41187,N_38074,N_38507);
or U41188 (N_41188,N_39526,N_38113);
nand U41189 (N_41189,N_38082,N_39932);
nand U41190 (N_41190,N_39928,N_39364);
xnor U41191 (N_41191,N_38779,N_38808);
and U41192 (N_41192,N_39208,N_39116);
or U41193 (N_41193,N_39186,N_39213);
nand U41194 (N_41194,N_39192,N_38833);
or U41195 (N_41195,N_38555,N_39597);
or U41196 (N_41196,N_39293,N_38859);
and U41197 (N_41197,N_39503,N_39931);
nor U41198 (N_41198,N_38977,N_39426);
or U41199 (N_41199,N_39583,N_39363);
or U41200 (N_41200,N_38696,N_39670);
nand U41201 (N_41201,N_39114,N_38678);
nand U41202 (N_41202,N_38944,N_38815);
or U41203 (N_41203,N_39291,N_38869);
or U41204 (N_41204,N_39177,N_39521);
nor U41205 (N_41205,N_38336,N_39565);
and U41206 (N_41206,N_39441,N_39961);
xor U41207 (N_41207,N_38474,N_39445);
nand U41208 (N_41208,N_39052,N_38420);
nand U41209 (N_41209,N_38188,N_38870);
and U41210 (N_41210,N_39820,N_38061);
xnor U41211 (N_41211,N_39674,N_39096);
xor U41212 (N_41212,N_38300,N_39275);
and U41213 (N_41213,N_38856,N_39679);
nor U41214 (N_41214,N_38010,N_38596);
nand U41215 (N_41215,N_39458,N_39798);
xor U41216 (N_41216,N_38726,N_39896);
nand U41217 (N_41217,N_39042,N_38726);
or U41218 (N_41218,N_38847,N_38036);
nand U41219 (N_41219,N_39229,N_38115);
nand U41220 (N_41220,N_38532,N_38127);
xor U41221 (N_41221,N_38097,N_38794);
and U41222 (N_41222,N_39216,N_39921);
or U41223 (N_41223,N_39906,N_39837);
nand U41224 (N_41224,N_39860,N_38525);
nand U41225 (N_41225,N_38726,N_38215);
or U41226 (N_41226,N_38814,N_39801);
nand U41227 (N_41227,N_39627,N_39329);
or U41228 (N_41228,N_38255,N_38537);
or U41229 (N_41229,N_38723,N_38173);
xnor U41230 (N_41230,N_39921,N_38448);
xor U41231 (N_41231,N_39155,N_39386);
or U41232 (N_41232,N_38981,N_38160);
nor U41233 (N_41233,N_39628,N_39278);
and U41234 (N_41234,N_39904,N_38799);
or U41235 (N_41235,N_38420,N_38224);
or U41236 (N_41236,N_39475,N_38413);
nand U41237 (N_41237,N_38054,N_38223);
and U41238 (N_41238,N_38206,N_39333);
xnor U41239 (N_41239,N_39916,N_38258);
nor U41240 (N_41240,N_38242,N_38100);
nor U41241 (N_41241,N_38959,N_38480);
or U41242 (N_41242,N_38833,N_38895);
nand U41243 (N_41243,N_39594,N_38745);
or U41244 (N_41244,N_39755,N_39147);
xnor U41245 (N_41245,N_39979,N_38235);
xor U41246 (N_41246,N_39204,N_39247);
nand U41247 (N_41247,N_38371,N_39141);
or U41248 (N_41248,N_39106,N_38794);
or U41249 (N_41249,N_39311,N_38787);
and U41250 (N_41250,N_38724,N_39846);
nand U41251 (N_41251,N_38280,N_38353);
nor U41252 (N_41252,N_38723,N_38205);
or U41253 (N_41253,N_38434,N_39452);
and U41254 (N_41254,N_39490,N_38299);
or U41255 (N_41255,N_38042,N_38611);
and U41256 (N_41256,N_38549,N_38951);
and U41257 (N_41257,N_39981,N_38893);
nor U41258 (N_41258,N_39501,N_38563);
nand U41259 (N_41259,N_39203,N_39430);
and U41260 (N_41260,N_39024,N_38614);
xor U41261 (N_41261,N_38159,N_38310);
and U41262 (N_41262,N_38094,N_38987);
nand U41263 (N_41263,N_38683,N_38150);
nor U41264 (N_41264,N_38764,N_39943);
or U41265 (N_41265,N_39050,N_39974);
nor U41266 (N_41266,N_38847,N_38736);
nand U41267 (N_41267,N_39821,N_39490);
xor U41268 (N_41268,N_39025,N_39876);
xnor U41269 (N_41269,N_39894,N_39572);
and U41270 (N_41270,N_39363,N_38578);
nand U41271 (N_41271,N_39918,N_38827);
xor U41272 (N_41272,N_38007,N_39131);
nand U41273 (N_41273,N_39020,N_38082);
xor U41274 (N_41274,N_39193,N_38072);
xnor U41275 (N_41275,N_39937,N_38263);
xor U41276 (N_41276,N_39412,N_39082);
nand U41277 (N_41277,N_38619,N_39916);
xor U41278 (N_41278,N_38606,N_38423);
nand U41279 (N_41279,N_39168,N_38677);
xnor U41280 (N_41280,N_39592,N_39282);
nor U41281 (N_41281,N_38552,N_39838);
nor U41282 (N_41282,N_39349,N_38228);
nor U41283 (N_41283,N_39419,N_39163);
or U41284 (N_41284,N_38546,N_38598);
or U41285 (N_41285,N_39463,N_39813);
nor U41286 (N_41286,N_39724,N_38608);
or U41287 (N_41287,N_39364,N_38173);
nand U41288 (N_41288,N_38568,N_39976);
xor U41289 (N_41289,N_39485,N_39670);
and U41290 (N_41290,N_38478,N_38922);
nand U41291 (N_41291,N_39875,N_38279);
and U41292 (N_41292,N_39868,N_38618);
and U41293 (N_41293,N_39963,N_38901);
or U41294 (N_41294,N_39361,N_38945);
xor U41295 (N_41295,N_38120,N_39313);
nor U41296 (N_41296,N_39847,N_38852);
and U41297 (N_41297,N_38336,N_39484);
or U41298 (N_41298,N_39151,N_39826);
nand U41299 (N_41299,N_38995,N_38114);
and U41300 (N_41300,N_39021,N_38834);
and U41301 (N_41301,N_38886,N_38519);
nor U41302 (N_41302,N_39026,N_38416);
and U41303 (N_41303,N_38839,N_38036);
nor U41304 (N_41304,N_39388,N_39192);
or U41305 (N_41305,N_39003,N_39969);
or U41306 (N_41306,N_39290,N_39123);
and U41307 (N_41307,N_39675,N_38217);
or U41308 (N_41308,N_39151,N_38850);
nand U41309 (N_41309,N_39145,N_38046);
nor U41310 (N_41310,N_38069,N_38469);
nand U41311 (N_41311,N_39253,N_38236);
or U41312 (N_41312,N_39577,N_39181);
xor U41313 (N_41313,N_39648,N_39137);
and U41314 (N_41314,N_39480,N_39618);
nand U41315 (N_41315,N_39741,N_38468);
nand U41316 (N_41316,N_38665,N_39150);
or U41317 (N_41317,N_38995,N_39281);
nor U41318 (N_41318,N_38286,N_38611);
nand U41319 (N_41319,N_39854,N_38772);
nand U41320 (N_41320,N_38383,N_38327);
and U41321 (N_41321,N_38575,N_39301);
nor U41322 (N_41322,N_38269,N_39904);
nor U41323 (N_41323,N_38015,N_38699);
and U41324 (N_41324,N_38048,N_39656);
or U41325 (N_41325,N_38761,N_39902);
or U41326 (N_41326,N_38303,N_39850);
nor U41327 (N_41327,N_39846,N_39813);
nor U41328 (N_41328,N_39303,N_39419);
or U41329 (N_41329,N_38922,N_38576);
xor U41330 (N_41330,N_38804,N_38672);
nor U41331 (N_41331,N_39127,N_39409);
nand U41332 (N_41332,N_39611,N_38973);
or U41333 (N_41333,N_39108,N_38086);
xnor U41334 (N_41334,N_39375,N_38101);
xnor U41335 (N_41335,N_39188,N_39993);
nand U41336 (N_41336,N_38330,N_39726);
or U41337 (N_41337,N_38328,N_38435);
or U41338 (N_41338,N_39964,N_39648);
and U41339 (N_41339,N_39089,N_39734);
xnor U41340 (N_41340,N_39092,N_39830);
and U41341 (N_41341,N_38863,N_39812);
nand U41342 (N_41342,N_39782,N_38356);
or U41343 (N_41343,N_38738,N_39022);
and U41344 (N_41344,N_38232,N_39095);
xor U41345 (N_41345,N_38537,N_38620);
nand U41346 (N_41346,N_38073,N_38625);
nor U41347 (N_41347,N_39757,N_38093);
nand U41348 (N_41348,N_38812,N_39934);
and U41349 (N_41349,N_39905,N_38170);
nor U41350 (N_41350,N_39058,N_38332);
or U41351 (N_41351,N_38347,N_39514);
and U41352 (N_41352,N_39347,N_38856);
xor U41353 (N_41353,N_39820,N_39752);
or U41354 (N_41354,N_38231,N_38684);
nor U41355 (N_41355,N_39045,N_38157);
and U41356 (N_41356,N_39647,N_39745);
nor U41357 (N_41357,N_38331,N_38573);
or U41358 (N_41358,N_38517,N_38522);
nor U41359 (N_41359,N_38229,N_39026);
nor U41360 (N_41360,N_39692,N_38557);
xor U41361 (N_41361,N_38640,N_39519);
nand U41362 (N_41362,N_38480,N_39692);
nand U41363 (N_41363,N_39577,N_39785);
or U41364 (N_41364,N_38996,N_39763);
and U41365 (N_41365,N_38904,N_39554);
and U41366 (N_41366,N_39235,N_38565);
and U41367 (N_41367,N_39191,N_38673);
or U41368 (N_41368,N_39524,N_38163);
or U41369 (N_41369,N_38392,N_38531);
xnor U41370 (N_41370,N_38496,N_38129);
nand U41371 (N_41371,N_38550,N_38995);
and U41372 (N_41372,N_38006,N_39273);
or U41373 (N_41373,N_39892,N_39243);
nor U41374 (N_41374,N_38432,N_38056);
nor U41375 (N_41375,N_39378,N_38135);
xnor U41376 (N_41376,N_38610,N_39220);
or U41377 (N_41377,N_38329,N_39526);
and U41378 (N_41378,N_38078,N_39384);
nand U41379 (N_41379,N_38552,N_38547);
and U41380 (N_41380,N_39525,N_38519);
and U41381 (N_41381,N_39653,N_39701);
xor U41382 (N_41382,N_39556,N_38537);
and U41383 (N_41383,N_39242,N_38075);
xnor U41384 (N_41384,N_38184,N_39430);
nand U41385 (N_41385,N_39058,N_39074);
nand U41386 (N_41386,N_39234,N_39002);
and U41387 (N_41387,N_38576,N_39530);
or U41388 (N_41388,N_38016,N_39325);
nand U41389 (N_41389,N_39609,N_39110);
nor U41390 (N_41390,N_39974,N_39448);
or U41391 (N_41391,N_38678,N_38217);
xnor U41392 (N_41392,N_39421,N_38805);
and U41393 (N_41393,N_38926,N_39092);
or U41394 (N_41394,N_38391,N_39386);
and U41395 (N_41395,N_38057,N_39709);
nand U41396 (N_41396,N_39023,N_39316);
and U41397 (N_41397,N_38851,N_39437);
xor U41398 (N_41398,N_38311,N_39281);
nand U41399 (N_41399,N_38690,N_39822);
and U41400 (N_41400,N_39194,N_39627);
nand U41401 (N_41401,N_39105,N_38494);
nand U41402 (N_41402,N_38035,N_39908);
nor U41403 (N_41403,N_39070,N_39337);
and U41404 (N_41404,N_38472,N_39789);
nand U41405 (N_41405,N_38985,N_39560);
nand U41406 (N_41406,N_38530,N_38150);
nor U41407 (N_41407,N_38612,N_39260);
nand U41408 (N_41408,N_39967,N_39337);
and U41409 (N_41409,N_38747,N_38107);
or U41410 (N_41410,N_38643,N_39752);
nor U41411 (N_41411,N_39649,N_38916);
xor U41412 (N_41412,N_39883,N_38300);
nand U41413 (N_41413,N_38441,N_39269);
nand U41414 (N_41414,N_38737,N_39919);
nor U41415 (N_41415,N_38352,N_38321);
nor U41416 (N_41416,N_39406,N_38325);
nand U41417 (N_41417,N_38618,N_38388);
and U41418 (N_41418,N_38975,N_38300);
xor U41419 (N_41419,N_38837,N_38581);
and U41420 (N_41420,N_39980,N_38259);
nand U41421 (N_41421,N_38791,N_39861);
and U41422 (N_41422,N_38842,N_38793);
nand U41423 (N_41423,N_39673,N_38263);
nand U41424 (N_41424,N_38690,N_39214);
xor U41425 (N_41425,N_39079,N_39125);
or U41426 (N_41426,N_38898,N_38440);
nand U41427 (N_41427,N_38094,N_38980);
xor U41428 (N_41428,N_38047,N_38230);
nand U41429 (N_41429,N_39606,N_38228);
and U41430 (N_41430,N_38977,N_38361);
xnor U41431 (N_41431,N_39970,N_39111);
nand U41432 (N_41432,N_39717,N_38985);
xnor U41433 (N_41433,N_39937,N_38783);
and U41434 (N_41434,N_39067,N_39469);
nor U41435 (N_41435,N_39769,N_39893);
xnor U41436 (N_41436,N_39039,N_39912);
and U41437 (N_41437,N_39478,N_38130);
and U41438 (N_41438,N_38811,N_38311);
and U41439 (N_41439,N_38056,N_38176);
nand U41440 (N_41440,N_38691,N_39612);
nor U41441 (N_41441,N_39802,N_38161);
nor U41442 (N_41442,N_39679,N_38992);
xnor U41443 (N_41443,N_38621,N_39541);
xnor U41444 (N_41444,N_39339,N_39472);
nand U41445 (N_41445,N_39102,N_38339);
nor U41446 (N_41446,N_38783,N_38556);
or U41447 (N_41447,N_38408,N_39201);
and U41448 (N_41448,N_39428,N_38071);
xor U41449 (N_41449,N_39781,N_38057);
nand U41450 (N_41450,N_39891,N_38751);
nand U41451 (N_41451,N_39441,N_39283);
nand U41452 (N_41452,N_38138,N_38152);
nor U41453 (N_41453,N_38985,N_39204);
or U41454 (N_41454,N_39250,N_39013);
nand U41455 (N_41455,N_38462,N_38018);
nand U41456 (N_41456,N_38124,N_38819);
nor U41457 (N_41457,N_38970,N_39429);
and U41458 (N_41458,N_39873,N_39261);
or U41459 (N_41459,N_39339,N_38123);
and U41460 (N_41460,N_38592,N_38252);
or U41461 (N_41461,N_38569,N_38919);
and U41462 (N_41462,N_39402,N_39875);
xor U41463 (N_41463,N_38266,N_39404);
or U41464 (N_41464,N_39768,N_39357);
nor U41465 (N_41465,N_39546,N_38019);
nand U41466 (N_41466,N_38772,N_38536);
xor U41467 (N_41467,N_39740,N_38634);
nor U41468 (N_41468,N_38208,N_38018);
and U41469 (N_41469,N_39691,N_38487);
xnor U41470 (N_41470,N_38492,N_39711);
nand U41471 (N_41471,N_39122,N_39080);
and U41472 (N_41472,N_38243,N_38350);
xnor U41473 (N_41473,N_38799,N_38120);
nand U41474 (N_41474,N_38311,N_39621);
nor U41475 (N_41475,N_38244,N_39920);
and U41476 (N_41476,N_38435,N_38015);
xor U41477 (N_41477,N_38074,N_38095);
nand U41478 (N_41478,N_39976,N_38372);
xnor U41479 (N_41479,N_39222,N_38852);
nand U41480 (N_41480,N_38996,N_39285);
nand U41481 (N_41481,N_39249,N_39652);
or U41482 (N_41482,N_38135,N_38889);
or U41483 (N_41483,N_38874,N_38982);
nor U41484 (N_41484,N_38169,N_38880);
xnor U41485 (N_41485,N_38178,N_38182);
or U41486 (N_41486,N_38707,N_38394);
and U41487 (N_41487,N_38357,N_38527);
and U41488 (N_41488,N_38464,N_38519);
nand U41489 (N_41489,N_39952,N_39150);
xor U41490 (N_41490,N_39214,N_39505);
xnor U41491 (N_41491,N_38181,N_38102);
or U41492 (N_41492,N_38282,N_38034);
nand U41493 (N_41493,N_38179,N_38816);
nand U41494 (N_41494,N_38599,N_39138);
xor U41495 (N_41495,N_39591,N_39414);
nor U41496 (N_41496,N_38252,N_39644);
or U41497 (N_41497,N_39302,N_38722);
or U41498 (N_41498,N_39651,N_38571);
xnor U41499 (N_41499,N_39035,N_38232);
or U41500 (N_41500,N_38145,N_38907);
xor U41501 (N_41501,N_38531,N_39987);
nand U41502 (N_41502,N_39980,N_38069);
and U41503 (N_41503,N_38358,N_39706);
nor U41504 (N_41504,N_38540,N_39127);
or U41505 (N_41505,N_39914,N_38102);
or U41506 (N_41506,N_38407,N_39862);
or U41507 (N_41507,N_39845,N_38241);
and U41508 (N_41508,N_38606,N_39930);
or U41509 (N_41509,N_39399,N_39993);
or U41510 (N_41510,N_39454,N_39330);
nor U41511 (N_41511,N_38637,N_38519);
nor U41512 (N_41512,N_38866,N_39135);
xnor U41513 (N_41513,N_39415,N_39246);
and U41514 (N_41514,N_39165,N_39643);
xnor U41515 (N_41515,N_38630,N_38545);
or U41516 (N_41516,N_38145,N_39259);
and U41517 (N_41517,N_39216,N_39700);
xor U41518 (N_41518,N_38152,N_38318);
and U41519 (N_41519,N_39983,N_39304);
and U41520 (N_41520,N_38247,N_39481);
xnor U41521 (N_41521,N_38308,N_38188);
or U41522 (N_41522,N_39092,N_39994);
nand U41523 (N_41523,N_39868,N_39114);
xor U41524 (N_41524,N_38235,N_38897);
xnor U41525 (N_41525,N_38646,N_38478);
nand U41526 (N_41526,N_39631,N_39929);
or U41527 (N_41527,N_39394,N_38738);
and U41528 (N_41528,N_39775,N_38089);
nor U41529 (N_41529,N_38617,N_38752);
nand U41530 (N_41530,N_38638,N_39681);
nand U41531 (N_41531,N_38747,N_38717);
and U41532 (N_41532,N_38357,N_39970);
and U41533 (N_41533,N_38742,N_38986);
nand U41534 (N_41534,N_38596,N_39336);
xnor U41535 (N_41535,N_38312,N_38498);
or U41536 (N_41536,N_38788,N_39590);
or U41537 (N_41537,N_39115,N_38057);
nand U41538 (N_41538,N_38899,N_39766);
or U41539 (N_41539,N_38037,N_39302);
or U41540 (N_41540,N_39423,N_39375);
nand U41541 (N_41541,N_39502,N_39557);
nand U41542 (N_41542,N_38431,N_39576);
xor U41543 (N_41543,N_39620,N_38700);
xor U41544 (N_41544,N_38201,N_39293);
xor U41545 (N_41545,N_38045,N_38923);
nor U41546 (N_41546,N_38876,N_38482);
nand U41547 (N_41547,N_39147,N_38100);
and U41548 (N_41548,N_38704,N_39453);
xor U41549 (N_41549,N_39580,N_38037);
xnor U41550 (N_41550,N_39313,N_38262);
nand U41551 (N_41551,N_38055,N_38140);
or U41552 (N_41552,N_39958,N_39045);
xor U41553 (N_41553,N_38712,N_39008);
or U41554 (N_41554,N_39240,N_38114);
nand U41555 (N_41555,N_39045,N_39396);
or U41556 (N_41556,N_38703,N_39108);
or U41557 (N_41557,N_38514,N_38921);
xor U41558 (N_41558,N_39603,N_38653);
nor U41559 (N_41559,N_39748,N_38077);
or U41560 (N_41560,N_38225,N_38578);
nor U41561 (N_41561,N_38748,N_38547);
nand U41562 (N_41562,N_38195,N_39677);
xor U41563 (N_41563,N_38106,N_38392);
xnor U41564 (N_41564,N_38493,N_39982);
nor U41565 (N_41565,N_39798,N_38142);
or U41566 (N_41566,N_38935,N_39721);
and U41567 (N_41567,N_39807,N_38326);
and U41568 (N_41568,N_38451,N_39611);
or U41569 (N_41569,N_39463,N_39947);
and U41570 (N_41570,N_38681,N_38257);
nand U41571 (N_41571,N_39688,N_39013);
or U41572 (N_41572,N_39734,N_39211);
nor U41573 (N_41573,N_39402,N_38417);
nor U41574 (N_41574,N_38714,N_39532);
nor U41575 (N_41575,N_39820,N_39312);
and U41576 (N_41576,N_39043,N_38463);
or U41577 (N_41577,N_38231,N_39785);
and U41578 (N_41578,N_39982,N_38899);
nor U41579 (N_41579,N_39790,N_38577);
nand U41580 (N_41580,N_39301,N_38697);
or U41581 (N_41581,N_38816,N_39697);
and U41582 (N_41582,N_39919,N_38907);
nand U41583 (N_41583,N_39938,N_39261);
and U41584 (N_41584,N_39767,N_38584);
nand U41585 (N_41585,N_39338,N_39774);
nand U41586 (N_41586,N_38835,N_39659);
or U41587 (N_41587,N_38643,N_38727);
or U41588 (N_41588,N_38237,N_38642);
and U41589 (N_41589,N_39355,N_38435);
xor U41590 (N_41590,N_38388,N_39442);
and U41591 (N_41591,N_39488,N_39728);
and U41592 (N_41592,N_39045,N_38786);
xor U41593 (N_41593,N_38043,N_38632);
nor U41594 (N_41594,N_38591,N_39402);
or U41595 (N_41595,N_39093,N_39428);
and U41596 (N_41596,N_38252,N_39065);
nand U41597 (N_41597,N_39631,N_39088);
nand U41598 (N_41598,N_38854,N_38186);
and U41599 (N_41599,N_38082,N_38060);
nor U41600 (N_41600,N_39916,N_39326);
xnor U41601 (N_41601,N_39828,N_38984);
nor U41602 (N_41602,N_38423,N_38109);
and U41603 (N_41603,N_38227,N_38501);
and U41604 (N_41604,N_38773,N_39227);
and U41605 (N_41605,N_38010,N_38858);
xor U41606 (N_41606,N_39636,N_39128);
or U41607 (N_41607,N_39735,N_39382);
nor U41608 (N_41608,N_38664,N_38004);
or U41609 (N_41609,N_39898,N_39327);
nor U41610 (N_41610,N_38207,N_39782);
xor U41611 (N_41611,N_38882,N_39658);
xnor U41612 (N_41612,N_38524,N_39053);
and U41613 (N_41613,N_39028,N_38826);
or U41614 (N_41614,N_38549,N_38285);
and U41615 (N_41615,N_38997,N_38923);
nand U41616 (N_41616,N_39757,N_38917);
xor U41617 (N_41617,N_39395,N_39072);
and U41618 (N_41618,N_39505,N_39935);
nand U41619 (N_41619,N_38421,N_39922);
and U41620 (N_41620,N_39992,N_38047);
and U41621 (N_41621,N_38765,N_39300);
and U41622 (N_41622,N_38247,N_38232);
and U41623 (N_41623,N_39977,N_39390);
nand U41624 (N_41624,N_39961,N_39509);
or U41625 (N_41625,N_39232,N_38366);
nand U41626 (N_41626,N_38601,N_39151);
and U41627 (N_41627,N_39856,N_38973);
nor U41628 (N_41628,N_39280,N_38934);
xnor U41629 (N_41629,N_38061,N_38903);
and U41630 (N_41630,N_38898,N_38476);
xor U41631 (N_41631,N_38640,N_39495);
and U41632 (N_41632,N_38216,N_38669);
and U41633 (N_41633,N_39663,N_39986);
or U41634 (N_41634,N_38590,N_38511);
nor U41635 (N_41635,N_38985,N_39974);
nor U41636 (N_41636,N_38507,N_39373);
xnor U41637 (N_41637,N_39103,N_39240);
and U41638 (N_41638,N_38278,N_38999);
xor U41639 (N_41639,N_38679,N_39130);
or U41640 (N_41640,N_39154,N_39347);
nor U41641 (N_41641,N_39538,N_39969);
nand U41642 (N_41642,N_38867,N_38713);
nand U41643 (N_41643,N_39962,N_38246);
and U41644 (N_41644,N_38150,N_39003);
xnor U41645 (N_41645,N_38240,N_39094);
and U41646 (N_41646,N_38896,N_38501);
nand U41647 (N_41647,N_39612,N_38100);
or U41648 (N_41648,N_38785,N_39386);
or U41649 (N_41649,N_39467,N_38044);
and U41650 (N_41650,N_39647,N_39279);
xor U41651 (N_41651,N_38280,N_39627);
and U41652 (N_41652,N_38742,N_39326);
or U41653 (N_41653,N_38057,N_38604);
nor U41654 (N_41654,N_38930,N_39506);
xnor U41655 (N_41655,N_38224,N_39068);
xnor U41656 (N_41656,N_39975,N_39256);
nand U41657 (N_41657,N_38647,N_39544);
nand U41658 (N_41658,N_38738,N_38572);
nor U41659 (N_41659,N_38142,N_38371);
or U41660 (N_41660,N_39845,N_39183);
nor U41661 (N_41661,N_39012,N_39325);
nand U41662 (N_41662,N_38198,N_38279);
and U41663 (N_41663,N_39544,N_38002);
and U41664 (N_41664,N_38910,N_39931);
and U41665 (N_41665,N_39340,N_39612);
and U41666 (N_41666,N_38266,N_39390);
or U41667 (N_41667,N_38946,N_39533);
or U41668 (N_41668,N_39991,N_38511);
and U41669 (N_41669,N_38165,N_39996);
nor U41670 (N_41670,N_39775,N_39439);
xnor U41671 (N_41671,N_38500,N_39439);
nor U41672 (N_41672,N_39493,N_39693);
nand U41673 (N_41673,N_39065,N_38064);
nand U41674 (N_41674,N_38401,N_38190);
or U41675 (N_41675,N_38143,N_38812);
xnor U41676 (N_41676,N_39157,N_39747);
and U41677 (N_41677,N_38189,N_39279);
and U41678 (N_41678,N_39957,N_39784);
and U41679 (N_41679,N_39398,N_39014);
xnor U41680 (N_41680,N_39237,N_38579);
nor U41681 (N_41681,N_39472,N_38345);
and U41682 (N_41682,N_39514,N_38328);
and U41683 (N_41683,N_39817,N_39335);
and U41684 (N_41684,N_38329,N_39666);
or U41685 (N_41685,N_39209,N_38014);
xnor U41686 (N_41686,N_38038,N_38787);
and U41687 (N_41687,N_39800,N_39367);
nor U41688 (N_41688,N_39289,N_39937);
nand U41689 (N_41689,N_39936,N_39582);
and U41690 (N_41690,N_39759,N_39371);
nor U41691 (N_41691,N_38394,N_39831);
xor U41692 (N_41692,N_39184,N_38943);
xnor U41693 (N_41693,N_38418,N_38247);
and U41694 (N_41694,N_39954,N_39028);
nor U41695 (N_41695,N_38667,N_39556);
or U41696 (N_41696,N_38568,N_39027);
xor U41697 (N_41697,N_39948,N_39888);
nor U41698 (N_41698,N_39465,N_39383);
nand U41699 (N_41699,N_38855,N_39710);
and U41700 (N_41700,N_39915,N_39344);
xor U41701 (N_41701,N_38964,N_39655);
nor U41702 (N_41702,N_38971,N_38334);
xor U41703 (N_41703,N_39077,N_38554);
nor U41704 (N_41704,N_39646,N_39996);
or U41705 (N_41705,N_38194,N_38021);
nor U41706 (N_41706,N_39306,N_38709);
nand U41707 (N_41707,N_39376,N_38728);
nand U41708 (N_41708,N_38064,N_39147);
xor U41709 (N_41709,N_38876,N_38739);
xnor U41710 (N_41710,N_38449,N_38121);
nand U41711 (N_41711,N_39019,N_38878);
or U41712 (N_41712,N_39099,N_39312);
nand U41713 (N_41713,N_39287,N_39453);
or U41714 (N_41714,N_39606,N_38523);
nor U41715 (N_41715,N_38465,N_38209);
nor U41716 (N_41716,N_39215,N_38141);
xnor U41717 (N_41717,N_39513,N_39478);
nand U41718 (N_41718,N_38078,N_39524);
xnor U41719 (N_41719,N_39858,N_39540);
nand U41720 (N_41720,N_38363,N_39110);
xnor U41721 (N_41721,N_39771,N_38673);
xor U41722 (N_41722,N_38934,N_39940);
xor U41723 (N_41723,N_39425,N_38826);
xnor U41724 (N_41724,N_39197,N_39051);
and U41725 (N_41725,N_38794,N_39021);
or U41726 (N_41726,N_38717,N_39455);
nand U41727 (N_41727,N_38543,N_38310);
xnor U41728 (N_41728,N_38730,N_39274);
and U41729 (N_41729,N_38040,N_38645);
nand U41730 (N_41730,N_39635,N_39619);
or U41731 (N_41731,N_38269,N_39810);
and U41732 (N_41732,N_39877,N_39305);
and U41733 (N_41733,N_39206,N_38354);
nor U41734 (N_41734,N_39469,N_38040);
or U41735 (N_41735,N_39139,N_38383);
xor U41736 (N_41736,N_39278,N_38321);
xor U41737 (N_41737,N_38282,N_38473);
or U41738 (N_41738,N_38783,N_39032);
and U41739 (N_41739,N_39354,N_38684);
nand U41740 (N_41740,N_38878,N_38432);
or U41741 (N_41741,N_39844,N_39198);
nand U41742 (N_41742,N_39936,N_39637);
or U41743 (N_41743,N_38083,N_38586);
and U41744 (N_41744,N_39218,N_38765);
nand U41745 (N_41745,N_38673,N_38928);
nor U41746 (N_41746,N_38305,N_38297);
nand U41747 (N_41747,N_39213,N_39612);
and U41748 (N_41748,N_39120,N_39052);
nand U41749 (N_41749,N_39662,N_38516);
or U41750 (N_41750,N_38920,N_39994);
nor U41751 (N_41751,N_39100,N_39506);
or U41752 (N_41752,N_39306,N_38970);
nor U41753 (N_41753,N_39547,N_38530);
nand U41754 (N_41754,N_39139,N_38636);
and U41755 (N_41755,N_39148,N_39977);
or U41756 (N_41756,N_38843,N_38564);
and U41757 (N_41757,N_38886,N_38222);
nand U41758 (N_41758,N_39765,N_39722);
nand U41759 (N_41759,N_39329,N_38794);
nand U41760 (N_41760,N_39435,N_39148);
xor U41761 (N_41761,N_38034,N_38402);
xnor U41762 (N_41762,N_39018,N_38006);
and U41763 (N_41763,N_38647,N_39752);
and U41764 (N_41764,N_38479,N_39795);
or U41765 (N_41765,N_38907,N_39943);
nand U41766 (N_41766,N_38324,N_38201);
xor U41767 (N_41767,N_38333,N_38048);
nand U41768 (N_41768,N_38847,N_39281);
and U41769 (N_41769,N_39621,N_39170);
and U41770 (N_41770,N_38063,N_38325);
nor U41771 (N_41771,N_39865,N_39800);
nor U41772 (N_41772,N_38617,N_39757);
nand U41773 (N_41773,N_39274,N_38624);
nand U41774 (N_41774,N_38601,N_39350);
xnor U41775 (N_41775,N_39246,N_39343);
and U41776 (N_41776,N_39771,N_39383);
xor U41777 (N_41777,N_39556,N_39553);
nor U41778 (N_41778,N_39972,N_39033);
nand U41779 (N_41779,N_39625,N_39675);
or U41780 (N_41780,N_39062,N_38858);
xnor U41781 (N_41781,N_39273,N_39745);
nand U41782 (N_41782,N_38556,N_39142);
or U41783 (N_41783,N_39697,N_38038);
or U41784 (N_41784,N_39762,N_38355);
or U41785 (N_41785,N_38266,N_39330);
nor U41786 (N_41786,N_38582,N_38438);
or U41787 (N_41787,N_39226,N_38002);
xnor U41788 (N_41788,N_38084,N_38092);
nor U41789 (N_41789,N_39688,N_39918);
nor U41790 (N_41790,N_38343,N_38169);
nand U41791 (N_41791,N_39973,N_39686);
nand U41792 (N_41792,N_39412,N_39726);
nor U41793 (N_41793,N_38265,N_39775);
nor U41794 (N_41794,N_39468,N_39553);
or U41795 (N_41795,N_39105,N_38967);
and U41796 (N_41796,N_39984,N_39536);
nor U41797 (N_41797,N_39509,N_38266);
xnor U41798 (N_41798,N_38842,N_39819);
xor U41799 (N_41799,N_39861,N_39801);
or U41800 (N_41800,N_38976,N_39807);
nor U41801 (N_41801,N_38096,N_39357);
and U41802 (N_41802,N_38046,N_39314);
nand U41803 (N_41803,N_39605,N_39406);
and U41804 (N_41804,N_39861,N_39775);
nand U41805 (N_41805,N_39686,N_38106);
xnor U41806 (N_41806,N_38159,N_39646);
and U41807 (N_41807,N_38993,N_39273);
xor U41808 (N_41808,N_39998,N_39091);
or U41809 (N_41809,N_39005,N_38594);
xor U41810 (N_41810,N_39401,N_38563);
xor U41811 (N_41811,N_39647,N_39646);
or U41812 (N_41812,N_39718,N_39436);
nand U41813 (N_41813,N_38881,N_38176);
or U41814 (N_41814,N_39461,N_38602);
nor U41815 (N_41815,N_38528,N_38453);
and U41816 (N_41816,N_38069,N_38028);
nand U41817 (N_41817,N_39342,N_38225);
xnor U41818 (N_41818,N_39557,N_39608);
nor U41819 (N_41819,N_38664,N_39444);
or U41820 (N_41820,N_38469,N_38471);
xnor U41821 (N_41821,N_38984,N_39063);
and U41822 (N_41822,N_38943,N_38522);
xnor U41823 (N_41823,N_39586,N_39977);
nand U41824 (N_41824,N_38100,N_39984);
and U41825 (N_41825,N_39342,N_38524);
xor U41826 (N_41826,N_38069,N_39410);
nor U41827 (N_41827,N_38917,N_39838);
xnor U41828 (N_41828,N_39644,N_39681);
and U41829 (N_41829,N_38232,N_38675);
nand U41830 (N_41830,N_38719,N_38487);
nor U41831 (N_41831,N_39545,N_39648);
and U41832 (N_41832,N_38213,N_39161);
nand U41833 (N_41833,N_39996,N_38383);
xor U41834 (N_41834,N_39306,N_39310);
nor U41835 (N_41835,N_39261,N_39788);
nor U41836 (N_41836,N_38286,N_38096);
and U41837 (N_41837,N_39835,N_39623);
xor U41838 (N_41838,N_38922,N_39702);
and U41839 (N_41839,N_39732,N_38879);
or U41840 (N_41840,N_39089,N_39482);
xor U41841 (N_41841,N_38726,N_38934);
or U41842 (N_41842,N_39354,N_38877);
and U41843 (N_41843,N_38614,N_39878);
xor U41844 (N_41844,N_39992,N_39801);
nand U41845 (N_41845,N_38705,N_38746);
xor U41846 (N_41846,N_38845,N_39987);
nor U41847 (N_41847,N_39433,N_39732);
nand U41848 (N_41848,N_39402,N_38214);
and U41849 (N_41849,N_39736,N_38325);
nand U41850 (N_41850,N_39761,N_39804);
nand U41851 (N_41851,N_39481,N_38412);
xor U41852 (N_41852,N_39253,N_39742);
or U41853 (N_41853,N_39880,N_38138);
and U41854 (N_41854,N_38799,N_39136);
or U41855 (N_41855,N_38507,N_38932);
or U41856 (N_41856,N_39406,N_38432);
xnor U41857 (N_41857,N_38892,N_38306);
and U41858 (N_41858,N_38723,N_38041);
and U41859 (N_41859,N_39976,N_39447);
and U41860 (N_41860,N_39256,N_39969);
and U41861 (N_41861,N_39649,N_39182);
xor U41862 (N_41862,N_39840,N_39763);
nand U41863 (N_41863,N_39690,N_38283);
and U41864 (N_41864,N_39336,N_39226);
nor U41865 (N_41865,N_39518,N_38571);
xnor U41866 (N_41866,N_39193,N_38894);
nand U41867 (N_41867,N_39565,N_38198);
and U41868 (N_41868,N_38589,N_38901);
xnor U41869 (N_41869,N_38001,N_39435);
or U41870 (N_41870,N_38226,N_38110);
xnor U41871 (N_41871,N_39375,N_38134);
nand U41872 (N_41872,N_38501,N_39117);
and U41873 (N_41873,N_39104,N_39789);
nand U41874 (N_41874,N_39402,N_38955);
nand U41875 (N_41875,N_39736,N_39665);
or U41876 (N_41876,N_38617,N_38085);
nor U41877 (N_41877,N_38606,N_38153);
nand U41878 (N_41878,N_39897,N_39891);
or U41879 (N_41879,N_39926,N_39514);
nand U41880 (N_41880,N_38143,N_39539);
nand U41881 (N_41881,N_38392,N_39283);
or U41882 (N_41882,N_39361,N_38870);
or U41883 (N_41883,N_39247,N_39532);
and U41884 (N_41884,N_38243,N_38421);
and U41885 (N_41885,N_39562,N_39276);
and U41886 (N_41886,N_39113,N_39837);
and U41887 (N_41887,N_39665,N_38269);
and U41888 (N_41888,N_39223,N_39692);
or U41889 (N_41889,N_38264,N_38351);
nand U41890 (N_41890,N_38381,N_39922);
xnor U41891 (N_41891,N_38534,N_39958);
xnor U41892 (N_41892,N_39269,N_38438);
or U41893 (N_41893,N_38503,N_39052);
nand U41894 (N_41894,N_39237,N_38349);
or U41895 (N_41895,N_38224,N_39016);
and U41896 (N_41896,N_38041,N_38628);
or U41897 (N_41897,N_39884,N_39775);
nand U41898 (N_41898,N_38952,N_39673);
nand U41899 (N_41899,N_39574,N_39721);
nand U41900 (N_41900,N_38168,N_38196);
or U41901 (N_41901,N_39666,N_38994);
or U41902 (N_41902,N_38705,N_38700);
or U41903 (N_41903,N_38612,N_38692);
nand U41904 (N_41904,N_39477,N_39659);
or U41905 (N_41905,N_38430,N_39349);
and U41906 (N_41906,N_38550,N_38031);
nand U41907 (N_41907,N_38352,N_38943);
or U41908 (N_41908,N_38753,N_39630);
nand U41909 (N_41909,N_39442,N_38968);
or U41910 (N_41910,N_38950,N_38716);
nor U41911 (N_41911,N_39670,N_39327);
nor U41912 (N_41912,N_38368,N_39161);
xor U41913 (N_41913,N_39554,N_38890);
and U41914 (N_41914,N_39334,N_39512);
nand U41915 (N_41915,N_39458,N_39385);
or U41916 (N_41916,N_39670,N_39455);
nor U41917 (N_41917,N_38988,N_38556);
or U41918 (N_41918,N_39874,N_39915);
nor U41919 (N_41919,N_39459,N_39852);
xnor U41920 (N_41920,N_39944,N_39638);
nand U41921 (N_41921,N_38433,N_39459);
and U41922 (N_41922,N_38312,N_38985);
nor U41923 (N_41923,N_38086,N_38325);
xor U41924 (N_41924,N_39115,N_39356);
or U41925 (N_41925,N_38501,N_38265);
and U41926 (N_41926,N_39707,N_38635);
and U41927 (N_41927,N_38953,N_39925);
nand U41928 (N_41928,N_39342,N_38758);
nand U41929 (N_41929,N_39778,N_39954);
or U41930 (N_41930,N_38930,N_39574);
and U41931 (N_41931,N_38846,N_39220);
nor U41932 (N_41932,N_38417,N_39185);
or U41933 (N_41933,N_38397,N_38373);
or U41934 (N_41934,N_39799,N_38168);
xnor U41935 (N_41935,N_38066,N_38630);
xor U41936 (N_41936,N_39314,N_38301);
xnor U41937 (N_41937,N_38287,N_38001);
nor U41938 (N_41938,N_38786,N_39173);
and U41939 (N_41939,N_38086,N_39668);
or U41940 (N_41940,N_39011,N_38983);
and U41941 (N_41941,N_38556,N_38674);
nor U41942 (N_41942,N_39903,N_38985);
xnor U41943 (N_41943,N_38193,N_38627);
or U41944 (N_41944,N_38212,N_38120);
nor U41945 (N_41945,N_38695,N_39391);
or U41946 (N_41946,N_39450,N_38251);
xnor U41947 (N_41947,N_38200,N_38243);
or U41948 (N_41948,N_39965,N_38539);
and U41949 (N_41949,N_39733,N_39483);
nand U41950 (N_41950,N_39507,N_39999);
nand U41951 (N_41951,N_39768,N_39874);
or U41952 (N_41952,N_39854,N_39298);
nand U41953 (N_41953,N_39300,N_38786);
nor U41954 (N_41954,N_39306,N_38847);
or U41955 (N_41955,N_39244,N_39178);
nand U41956 (N_41956,N_38352,N_38516);
and U41957 (N_41957,N_39719,N_38134);
nor U41958 (N_41958,N_38757,N_39281);
xor U41959 (N_41959,N_39918,N_38687);
and U41960 (N_41960,N_39096,N_38561);
and U41961 (N_41961,N_39982,N_38845);
nand U41962 (N_41962,N_39637,N_39769);
and U41963 (N_41963,N_38202,N_39003);
nor U41964 (N_41964,N_38260,N_39366);
xnor U41965 (N_41965,N_39829,N_38855);
nand U41966 (N_41966,N_39392,N_39170);
xnor U41967 (N_41967,N_38044,N_39216);
nor U41968 (N_41968,N_38372,N_38082);
nand U41969 (N_41969,N_39090,N_38568);
and U41970 (N_41970,N_38038,N_39238);
xor U41971 (N_41971,N_38949,N_39532);
or U41972 (N_41972,N_38867,N_38590);
and U41973 (N_41973,N_38395,N_39772);
nor U41974 (N_41974,N_39531,N_38963);
nor U41975 (N_41975,N_39913,N_38819);
and U41976 (N_41976,N_39134,N_38590);
nor U41977 (N_41977,N_39027,N_38284);
nor U41978 (N_41978,N_38750,N_39535);
and U41979 (N_41979,N_38274,N_39061);
xnor U41980 (N_41980,N_38998,N_38862);
xor U41981 (N_41981,N_38333,N_38165);
and U41982 (N_41982,N_39249,N_38962);
nor U41983 (N_41983,N_39262,N_38389);
nand U41984 (N_41984,N_39869,N_39465);
or U41985 (N_41985,N_38442,N_39929);
or U41986 (N_41986,N_38058,N_38733);
nand U41987 (N_41987,N_38074,N_39754);
nor U41988 (N_41988,N_38249,N_39058);
nor U41989 (N_41989,N_38143,N_38186);
xnor U41990 (N_41990,N_39558,N_39347);
or U41991 (N_41991,N_39068,N_39179);
xnor U41992 (N_41992,N_38526,N_39268);
or U41993 (N_41993,N_39277,N_38973);
and U41994 (N_41994,N_38589,N_38221);
nor U41995 (N_41995,N_38841,N_38169);
nor U41996 (N_41996,N_39651,N_38407);
nand U41997 (N_41997,N_38451,N_38835);
and U41998 (N_41998,N_38222,N_38193);
nor U41999 (N_41999,N_39234,N_38818);
nand U42000 (N_42000,N_41865,N_40332);
xor U42001 (N_42001,N_41915,N_40722);
or U42002 (N_42002,N_41960,N_40289);
nor U42003 (N_42003,N_40612,N_41552);
or U42004 (N_42004,N_40991,N_41634);
xor U42005 (N_42005,N_41427,N_41350);
or U42006 (N_42006,N_40620,N_40685);
xnor U42007 (N_42007,N_41135,N_41781);
xnor U42008 (N_42008,N_41625,N_41872);
xnor U42009 (N_42009,N_41644,N_40918);
xor U42010 (N_42010,N_40753,N_40400);
nor U42011 (N_42011,N_40598,N_41927);
xnor U42012 (N_42012,N_40968,N_41438);
xor U42013 (N_42013,N_40259,N_40125);
or U42014 (N_42014,N_41793,N_41816);
xor U42015 (N_42015,N_40187,N_41950);
or U42016 (N_42016,N_40497,N_40762);
and U42017 (N_42017,N_41904,N_41482);
and U42018 (N_42018,N_41606,N_40085);
nand U42019 (N_42019,N_40500,N_41340);
or U42020 (N_42020,N_41954,N_40978);
xor U42021 (N_42021,N_40727,N_41422);
or U42022 (N_42022,N_41263,N_41726);
or U42023 (N_42023,N_41504,N_40358);
nor U42024 (N_42024,N_41678,N_41367);
nor U42025 (N_42025,N_40269,N_40094);
and U42026 (N_42026,N_40290,N_40997);
nand U42027 (N_42027,N_41188,N_41985);
nor U42028 (N_42028,N_41250,N_40380);
nand U42029 (N_42029,N_40787,N_40329);
and U42030 (N_42030,N_40975,N_41683);
and U42031 (N_42031,N_41016,N_40051);
nand U42032 (N_42032,N_41624,N_40238);
or U42033 (N_42033,N_40814,N_41332);
and U42034 (N_42034,N_40169,N_41414);
and U42035 (N_42035,N_40297,N_40286);
nor U42036 (N_42036,N_40234,N_41609);
nor U42037 (N_42037,N_40650,N_40222);
nor U42038 (N_42038,N_40462,N_40314);
xor U42039 (N_42039,N_40256,N_40327);
or U42040 (N_42040,N_41903,N_40107);
nor U42041 (N_42041,N_40534,N_40247);
and U42042 (N_42042,N_40388,N_41021);
nand U42043 (N_42043,N_40793,N_41933);
nor U42044 (N_42044,N_40794,N_41913);
nand U42045 (N_42045,N_40424,N_40869);
and U42046 (N_42046,N_40890,N_41175);
nand U42047 (N_42047,N_40928,N_41205);
nand U42048 (N_42048,N_40111,N_41900);
or U42049 (N_42049,N_41009,N_41481);
or U42050 (N_42050,N_41527,N_41329);
and U42051 (N_42051,N_41444,N_40653);
and U42052 (N_42052,N_41256,N_40059);
nand U42053 (N_42053,N_40318,N_40830);
xnor U42054 (N_42054,N_40819,N_41529);
xnor U42055 (N_42055,N_40158,N_40344);
nand U42056 (N_42056,N_40970,N_41743);
nor U42057 (N_42057,N_41072,N_40265);
or U42058 (N_42058,N_40093,N_40356);
xor U42059 (N_42059,N_41592,N_40788);
and U42060 (N_42060,N_41584,N_41947);
nand U42061 (N_42061,N_41730,N_41354);
xnor U42062 (N_42062,N_40113,N_41233);
nand U42063 (N_42063,N_41020,N_41965);
nor U42064 (N_42064,N_41671,N_40150);
nor U42065 (N_42065,N_41884,N_40376);
and U42066 (N_42066,N_41699,N_40213);
xnor U42067 (N_42067,N_41631,N_41075);
or U42068 (N_42068,N_40527,N_40268);
nand U42069 (N_42069,N_40924,N_41964);
nor U42070 (N_42070,N_41496,N_40503);
nand U42071 (N_42071,N_41081,N_40707);
xor U42072 (N_42072,N_40601,N_40427);
nand U42073 (N_42073,N_40480,N_41610);
nor U42074 (N_42074,N_40235,N_41531);
nor U42075 (N_42075,N_41299,N_41269);
or U42076 (N_42076,N_41526,N_41126);
or U42077 (N_42077,N_41371,N_40022);
nand U42078 (N_42078,N_40197,N_40587);
and U42079 (N_42079,N_40525,N_40531);
and U42080 (N_42080,N_41387,N_41488);
or U42081 (N_42081,N_41017,N_41405);
xnor U42082 (N_42082,N_41105,N_40553);
nor U42083 (N_42083,N_40335,N_40846);
or U42084 (N_42084,N_41448,N_41499);
nor U42085 (N_42085,N_41877,N_41672);
nor U42086 (N_42086,N_41362,N_40824);
xnor U42087 (N_42087,N_41109,N_41291);
xnor U42088 (N_42088,N_41996,N_40694);
xor U42089 (N_42089,N_41807,N_40962);
nand U42090 (N_42090,N_41317,N_40431);
and U42091 (N_42091,N_41782,N_40764);
nand U42092 (N_42092,N_40073,N_40972);
nand U42093 (N_42093,N_41429,N_41944);
xor U42094 (N_42094,N_40743,N_41220);
nand U42095 (N_42095,N_41246,N_40837);
and U42096 (N_42096,N_41945,N_41948);
xnor U42097 (N_42097,N_41045,N_40360);
and U42098 (N_42098,N_41599,N_41923);
nor U42099 (N_42099,N_40446,N_40906);
nand U42100 (N_42100,N_40010,N_41612);
xnor U42101 (N_42101,N_40628,N_41648);
nor U42102 (N_42102,N_40457,N_40664);
nand U42103 (N_42103,N_40602,N_40331);
xor U42104 (N_42104,N_41452,N_41008);
nand U42105 (N_42105,N_40780,N_40087);
nand U42106 (N_42106,N_41809,N_41393);
nor U42107 (N_42107,N_41590,N_41617);
xor U42108 (N_42108,N_40378,N_41495);
and U42109 (N_42109,N_41171,N_40605);
nand U42110 (N_42110,N_40119,N_41554);
or U42111 (N_42111,N_40663,N_41304);
nor U42112 (N_42112,N_41757,N_41516);
and U42113 (N_42113,N_40956,N_40834);
nand U42114 (N_42114,N_40060,N_40145);
nand U42115 (N_42115,N_40648,N_40625);
nor U42116 (N_42116,N_41077,N_40563);
or U42117 (N_42117,N_40366,N_40210);
or U42118 (N_42118,N_40237,N_40752);
and U42119 (N_42119,N_40025,N_40634);
nor U42120 (N_42120,N_41788,N_41528);
nand U42121 (N_42121,N_40273,N_41180);
nand U42122 (N_42122,N_41776,N_40401);
xnor U42123 (N_42123,N_40039,N_41618);
or U42124 (N_42124,N_41472,N_40275);
nor U42125 (N_42125,N_41643,N_40382);
nand U42126 (N_42126,N_41335,N_41160);
nor U42127 (N_42127,N_41303,N_41064);
or U42128 (N_42128,N_40614,N_41640);
nor U42129 (N_42129,N_41176,N_41986);
xnor U42130 (N_42130,N_40325,N_41875);
and U42131 (N_42131,N_41031,N_41787);
and U42132 (N_42132,N_41321,N_40729);
nand U42133 (N_42133,N_41929,N_41379);
nor U42134 (N_42134,N_40985,N_40310);
and U42135 (N_42135,N_41149,N_40436);
nor U42136 (N_42136,N_40948,N_41254);
and U42137 (N_42137,N_40532,N_41028);
nand U42138 (N_42138,N_41187,N_40746);
or U42139 (N_42139,N_40546,N_40180);
xor U42140 (N_42140,N_40923,N_40294);
and U42141 (N_42141,N_40712,N_40671);
nand U42142 (N_42142,N_41675,N_40800);
xnor U42143 (N_42143,N_40960,N_41976);
xor U42144 (N_42144,N_41852,N_41984);
and U42145 (N_42145,N_41011,N_40930);
nand U42146 (N_42146,N_41076,N_41662);
or U42147 (N_42147,N_41356,N_40496);
xnor U42148 (N_42148,N_41858,N_41539);
or U42149 (N_42149,N_41853,N_40047);
or U42150 (N_42150,N_40134,N_40434);
xor U42151 (N_42151,N_41044,N_41423);
or U42152 (N_42152,N_41754,N_40422);
nand U42153 (N_42153,N_40166,N_40319);
and U42154 (N_42154,N_41748,N_41523);
and U42155 (N_42155,N_40742,N_41215);
nand U42156 (N_42156,N_41975,N_41869);
nand U42157 (N_42157,N_41883,N_40526);
or U42158 (N_42158,N_41403,N_40823);
nand U42159 (N_42159,N_41733,N_41722);
nor U42160 (N_42160,N_40175,N_41494);
and U42161 (N_42161,N_41421,N_40304);
xor U42162 (N_42162,N_40233,N_40790);
and U42163 (N_42163,N_41708,N_41719);
nor U42164 (N_42164,N_41078,N_41433);
xnor U42165 (N_42165,N_40364,N_40333);
or U42166 (N_42166,N_41407,N_41093);
nor U42167 (N_42167,N_41475,N_40441);
xor U42168 (N_42168,N_40285,N_41172);
or U42169 (N_42169,N_40139,N_41148);
and U42170 (N_42170,N_40672,N_41157);
nand U42171 (N_42171,N_40755,N_40528);
nor U42172 (N_42172,N_40915,N_41766);
nor U42173 (N_42173,N_40413,N_41661);
xor U42174 (N_42174,N_40866,N_41343);
or U42175 (N_42175,N_41633,N_41473);
or U42176 (N_42176,N_41588,N_41131);
and U42177 (N_42177,N_40399,N_41518);
nand U42178 (N_42178,N_41839,N_40581);
nor U42179 (N_42179,N_40556,N_40949);
xor U42180 (N_42180,N_41326,N_40698);
or U42181 (N_42181,N_41988,N_41843);
or U42182 (N_42182,N_41870,N_41847);
xor U42183 (N_42183,N_41514,N_40120);
or U42184 (N_42184,N_40683,N_41619);
or U42185 (N_42185,N_41166,N_40944);
xor U42186 (N_42186,N_40463,N_41502);
xnor U42187 (N_42187,N_41761,N_40179);
and U42188 (N_42188,N_40686,N_40008);
or U42189 (N_42189,N_40130,N_41555);
nor U42190 (N_42190,N_40882,N_40980);
and U42191 (N_42191,N_40088,N_40354);
or U42192 (N_42192,N_40161,N_40315);
and U42193 (N_42193,N_40410,N_40937);
and U42194 (N_42194,N_40293,N_40573);
xor U42195 (N_42195,N_41971,N_40146);
nor U42196 (N_42196,N_41165,N_41183);
nand U42197 (N_42197,N_41653,N_40435);
or U42198 (N_42198,N_41038,N_41795);
or U42199 (N_42199,N_41741,N_41258);
nand U42200 (N_42200,N_40765,N_40695);
nand U42201 (N_42201,N_40679,N_41363);
nand U42202 (N_42202,N_41380,N_40630);
xor U42203 (N_42203,N_41118,N_41124);
nor U42204 (N_42204,N_41731,N_41104);
and U42205 (N_42205,N_41132,N_40868);
nor U42206 (N_42206,N_41435,N_40321);
nand U42207 (N_42207,N_40377,N_41597);
xnor U42208 (N_42208,N_40543,N_41336);
nand U42209 (N_42209,N_40056,N_40043);
or U42210 (N_42210,N_41202,N_41576);
nand U42211 (N_42211,N_40836,N_40456);
and U42212 (N_42212,N_41247,N_40542);
nand U42213 (N_42213,N_41533,N_41614);
nor U42214 (N_42214,N_40163,N_41510);
and U42215 (N_42215,N_41701,N_40078);
or U42216 (N_42216,N_40189,N_41979);
and U42217 (N_42217,N_41121,N_40292);
or U42218 (N_42218,N_40362,N_40375);
and U42219 (N_42219,N_40969,N_41241);
or U42220 (N_42220,N_41301,N_41096);
or U42221 (N_42221,N_40629,N_40328);
xnor U42222 (N_42222,N_41394,N_41308);
xnor U42223 (N_42223,N_40384,N_40407);
xor U42224 (N_42224,N_40552,N_40618);
nor U42225 (N_42225,N_40555,N_40839);
nand U42226 (N_42226,N_40444,N_40582);
and U42227 (N_42227,N_40034,N_40004);
or U42228 (N_42228,N_40943,N_41899);
xor U42229 (N_42229,N_41251,N_41377);
nor U42230 (N_42230,N_41449,N_41656);
xor U42231 (N_42231,N_41441,N_40693);
nor U42232 (N_42232,N_41764,N_41264);
nor U42233 (N_42233,N_40308,N_41862);
nor U42234 (N_42234,N_41928,N_41265);
or U42235 (N_42235,N_40263,N_40149);
nor U42236 (N_42236,N_41320,N_41842);
xor U42237 (N_42237,N_41262,N_40498);
or U42238 (N_42238,N_40749,N_40826);
nand U42239 (N_42239,N_40028,N_41231);
and U42240 (N_42240,N_41602,N_40964);
nand U42241 (N_42241,N_40536,N_40363);
nor U42242 (N_42242,N_41805,N_41637);
xnor U42243 (N_42243,N_40501,N_40522);
or U42244 (N_42244,N_40853,N_41818);
or U42245 (N_42245,N_41994,N_40430);
nor U42246 (N_42246,N_41092,N_40350);
or U42247 (N_42247,N_40639,N_40852);
or U42248 (N_42248,N_40517,N_41506);
xnor U42249 (N_42249,N_40876,N_40425);
nand U42250 (N_42250,N_41242,N_41874);
xor U42251 (N_42251,N_41322,N_40768);
and U42252 (N_42252,N_40061,N_40816);
xnor U42253 (N_42253,N_40880,N_41147);
xnor U42254 (N_42254,N_40505,N_41497);
nand U42255 (N_42255,N_41003,N_40433);
or U42256 (N_42256,N_41159,N_41706);
and U42257 (N_42257,N_40908,N_41015);
and U42258 (N_42258,N_40661,N_41574);
or U42259 (N_42259,N_40284,N_40603);
nor U42260 (N_42260,N_40954,N_41228);
nor U42261 (N_42261,N_41866,N_41930);
and U42262 (N_42262,N_40781,N_41978);
xor U42263 (N_42263,N_40984,N_41997);
and U42264 (N_42264,N_41673,N_40981);
or U42265 (N_42265,N_40894,N_41211);
xnor U42266 (N_42266,N_40044,N_41134);
nand U42267 (N_42267,N_41755,N_40224);
nor U42268 (N_42268,N_40538,N_41848);
or U42269 (N_42269,N_41418,N_41400);
or U42270 (N_42270,N_41562,N_40758);
xor U42271 (N_42271,N_40586,N_40223);
and U42272 (N_42272,N_40218,N_40607);
and U42273 (N_42273,N_41926,N_40696);
xnor U42274 (N_42274,N_41519,N_40005);
xnor U42275 (N_42275,N_41999,N_41342);
or U42276 (N_42276,N_40281,N_40334);
or U42277 (N_42277,N_41345,N_41738);
or U42278 (N_42278,N_40815,N_40127);
and U42279 (N_42279,N_40104,N_40253);
xnor U42280 (N_42280,N_40106,N_41829);
nand U42281 (N_42281,N_40348,N_40006);
nand U42282 (N_42282,N_40521,N_40231);
or U42283 (N_42283,N_40706,N_40476);
nor U42284 (N_42284,N_41388,N_41587);
nand U42285 (N_42285,N_41920,N_41060);
nor U42286 (N_42286,N_40792,N_40718);
xor U42287 (N_42287,N_40379,N_41910);
or U42288 (N_42288,N_40151,N_41995);
xnor U42289 (N_42289,N_41810,N_41613);
or U42290 (N_42290,N_40575,N_40799);
xor U42291 (N_42291,N_40199,N_40907);
xor U42292 (N_42292,N_40075,N_40458);
and U42293 (N_42293,N_41358,N_41245);
nand U42294 (N_42294,N_40646,N_41040);
nand U42295 (N_42295,N_41989,N_41991);
nor U42296 (N_42296,N_41550,N_40961);
xnor U42297 (N_42297,N_41981,N_40137);
and U42298 (N_42298,N_41477,N_40267);
nor U42299 (N_42299,N_40885,N_40099);
nand U42300 (N_42300,N_41703,N_40579);
nor U42301 (N_42301,N_40050,N_40188);
xnor U42302 (N_42302,N_41771,N_40979);
or U42303 (N_42303,N_40109,N_41218);
and U42304 (N_42304,N_41445,N_40802);
nand U42305 (N_42305,N_41668,N_40771);
xnor U42306 (N_42306,N_41275,N_41177);
or U42307 (N_42307,N_41049,N_40174);
nor U42308 (N_42308,N_40214,N_41556);
and U42309 (N_42309,N_41993,N_40687);
and U42310 (N_42310,N_40156,N_40867);
and U42311 (N_42311,N_40699,N_41549);
and U42312 (N_42312,N_41489,N_41143);
and U42313 (N_42313,N_41749,N_40609);
nor U42314 (N_42314,N_40029,N_40515);
nand U42315 (N_42315,N_40030,N_41714);
or U42316 (N_42316,N_40535,N_41416);
nand U42317 (N_42317,N_41398,N_40881);
nor U42318 (N_42318,N_40772,N_40019);
and U42319 (N_42319,N_41774,N_41838);
xnor U42320 (N_42320,N_40927,N_40323);
or U42321 (N_42321,N_40662,N_40838);
and U42322 (N_42322,N_41314,N_40805);
xnor U42323 (N_42323,N_40903,N_41718);
xnor U42324 (N_42324,N_41369,N_40668);
nand U42325 (N_42325,N_40225,N_40776);
xnor U42326 (N_42326,N_41088,N_41271);
and U42327 (N_42327,N_41669,N_41337);
nand U42328 (N_42328,N_41144,N_41911);
xnor U42329 (N_42329,N_41036,N_40829);
nand U42330 (N_42330,N_41541,N_41811);
nor U42331 (N_42331,N_40299,N_40529);
nor U42332 (N_42332,N_40052,N_41067);
xnor U42333 (N_42333,N_40596,N_40467);
and U42334 (N_42334,N_41392,N_41267);
xor U42335 (N_42335,N_40647,N_41626);
and U42336 (N_42336,N_40549,N_41952);
nor U42337 (N_42337,N_41545,N_40066);
nor U42338 (N_42338,N_40057,N_40511);
or U42339 (N_42339,N_41420,N_40254);
and U42340 (N_42340,N_40089,N_41660);
nor U42341 (N_42341,N_40578,N_41074);
nand U42342 (N_42342,N_41199,N_40658);
or U42343 (N_42343,N_40250,N_40568);
or U42344 (N_42344,N_40572,N_41799);
nor U42345 (N_42345,N_40420,N_41413);
or U42346 (N_42346,N_41227,N_40688);
nand U42347 (N_42347,N_40847,N_41492);
xnor U42348 (N_42348,N_41191,N_40390);
nand U42349 (N_42349,N_41977,N_40121);
and U42350 (N_42350,N_41447,N_40063);
and U42351 (N_42351,N_41066,N_40919);
and U42352 (N_42352,N_41879,N_40701);
and U42353 (N_42353,N_41068,N_41351);
xor U42354 (N_42354,N_40545,N_40888);
xor U42355 (N_42355,N_40081,N_41399);
xnor U42356 (N_42356,N_41462,N_41294);
nor U42357 (N_42357,N_41410,N_40198);
and U42358 (N_42358,N_41864,N_41917);
nand U42359 (N_42359,N_41750,N_41744);
nand U42360 (N_42360,N_40172,N_41470);
nand U42361 (N_42361,N_41196,N_41521);
nor U42362 (N_42362,N_41601,N_41374);
or U42363 (N_42363,N_41773,N_40372);
xnor U42364 (N_42364,N_40177,N_40370);
nand U42365 (N_42365,N_41747,N_41001);
or U42366 (N_42366,N_41130,N_41697);
xor U42367 (N_42367,N_40053,N_40351);
xor U42368 (N_42368,N_40404,N_40725);
and U42369 (N_42369,N_41270,N_40450);
nor U42370 (N_42370,N_40840,N_40822);
and U42371 (N_42371,N_40453,N_41295);
and U42372 (N_42372,N_40616,N_40655);
nand U42373 (N_42373,N_41006,N_40635);
and U42374 (N_42374,N_41004,N_41168);
and U42375 (N_42375,N_40872,N_41082);
and U42376 (N_42376,N_41098,N_41876);
xnor U42377 (N_42377,N_41658,N_40442);
and U42378 (N_42378,N_41501,N_40565);
xor U42379 (N_42379,N_40484,N_41953);
and U42380 (N_42380,N_40076,N_41779);
nand U42381 (N_42381,N_41179,N_40091);
nor U42382 (N_42382,N_40958,N_40443);
xor U42383 (N_42383,N_41107,N_41302);
or U42384 (N_42384,N_41902,N_41224);
nor U42385 (N_42385,N_41408,N_41146);
xor U42386 (N_42386,N_41959,N_41957);
and U42387 (N_42387,N_41012,N_40593);
and U42388 (N_42388,N_41834,N_40588);
or U42389 (N_42389,N_40623,N_40873);
and U42390 (N_42390,N_41801,N_41479);
nand U42391 (N_42391,N_41980,N_40103);
nand U42392 (N_42392,N_41663,N_41728);
or U42393 (N_42393,N_40312,N_40986);
xor U42394 (N_42394,N_40249,N_41353);
nand U42395 (N_42395,N_41820,N_40296);
nand U42396 (N_42396,N_41459,N_40574);
xnor U42397 (N_42397,N_40619,N_40295);
and U42398 (N_42398,N_40957,N_41288);
or U42399 (N_42399,N_41136,N_41305);
or U42400 (N_42400,N_40072,N_41182);
xnor U42401 (N_42401,N_41798,N_41682);
nor U42402 (N_42402,N_40719,N_41279);
nor U42403 (N_42403,N_41666,N_41559);
or U42404 (N_42404,N_40309,N_40313);
xnor U42405 (N_42405,N_41192,N_41649);
or U42406 (N_42406,N_40232,N_40606);
or U42407 (N_42407,N_41893,N_41327);
or U42408 (N_42408,N_41306,N_40406);
and U42409 (N_42409,N_40914,N_41936);
or U42410 (N_42410,N_40411,N_40395);
and U42411 (N_42411,N_40564,N_41992);
and U42412 (N_42412,N_40773,N_41282);
nor U42413 (N_42413,N_40054,N_41882);
nor U42414 (N_42414,N_41822,N_41232);
nor U42415 (N_42415,N_41628,N_40007);
nor U42416 (N_42416,N_40692,N_40064);
nand U42417 (N_42417,N_41156,N_41100);
nor U42418 (N_42418,N_41970,N_40069);
and U42419 (N_42419,N_41710,N_41101);
and U42420 (N_42420,N_40750,N_40717);
xnor U42421 (N_42421,N_41277,N_41513);
or U42422 (N_42422,N_41446,N_41384);
and U42423 (N_42423,N_41164,N_41832);
or U42424 (N_42424,N_40303,N_41402);
nor U42425 (N_42425,N_41286,N_40262);
and U42426 (N_42426,N_40058,N_40396);
nor U42427 (N_42427,N_41712,N_40594);
or U42428 (N_42428,N_41785,N_41013);
or U42429 (N_42429,N_41571,N_41208);
nor U42430 (N_42430,N_41128,N_40205);
nor U42431 (N_42431,N_40939,N_40864);
nand U42432 (N_42432,N_41700,N_41646);
and U42433 (N_42433,N_41434,N_41524);
or U42434 (N_42434,N_41690,N_40715);
nand U42435 (N_42435,N_41517,N_41162);
or U42436 (N_42436,N_40239,N_40394);
and U42437 (N_42437,N_41257,N_40080);
nand U42438 (N_42438,N_40541,N_41709);
nor U42439 (N_42439,N_40624,N_41688);
and U42440 (N_42440,N_41152,N_40920);
xor U42441 (N_42441,N_41824,N_40514);
and U42442 (N_42442,N_40946,N_40942);
nand U42443 (N_42443,N_40167,N_40935);
and U42444 (N_42444,N_40763,N_41685);
or U42445 (N_42445,N_40913,N_41087);
nor U42446 (N_42446,N_40381,N_40015);
xor U42447 (N_42447,N_40490,N_41018);
nand U42448 (N_42448,N_41907,N_41850);
or U42449 (N_42449,N_41558,N_40035);
nand U42450 (N_42450,N_41716,N_40176);
and U42451 (N_42451,N_41914,N_40341);
xnor U42452 (N_42452,N_41752,N_41827);
nand U42453 (N_42453,N_40708,N_41909);
nor U42454 (N_42454,N_41024,N_40155);
nor U42455 (N_42455,N_41505,N_40641);
or U42456 (N_42456,N_41207,N_40951);
nor U42457 (N_42457,N_40455,N_40898);
nor U42458 (N_42458,N_41620,N_40610);
nand U42459 (N_42459,N_41888,N_40633);
nand U42460 (N_42460,N_41347,N_41095);
or U42461 (N_42461,N_40468,N_41585);
nor U42462 (N_42462,N_41687,N_41276);
and U42463 (N_42463,N_40896,N_41339);
or U42464 (N_42464,N_40518,N_41278);
xnor U42465 (N_42465,N_40720,N_41361);
and U42466 (N_42466,N_40336,N_40181);
nor U42467 (N_42467,N_41789,N_40845);
xor U42468 (N_42468,N_40803,N_40482);
and U42469 (N_42469,N_41577,N_40649);
or U42470 (N_42470,N_40206,N_41823);
xnor U42471 (N_42471,N_41222,N_40544);
or U42472 (N_42472,N_40084,N_41120);
and U42473 (N_42473,N_40576,N_40171);
or U42474 (N_42474,N_41835,N_41652);
and U42475 (N_42475,N_40832,N_41490);
or U42476 (N_42476,N_41209,N_40797);
and U42477 (N_42477,N_41564,N_41670);
nor U42478 (N_42478,N_41071,N_40902);
nand U42479 (N_42479,N_41110,N_41840);
nand U42480 (N_42480,N_40105,N_40300);
or U42481 (N_42481,N_41775,N_40808);
and U42482 (N_42482,N_41050,N_41509);
and U42483 (N_42483,N_41252,N_41122);
and U42484 (N_42484,N_40392,N_41476);
nand U42485 (N_42485,N_40317,N_40884);
xor U42486 (N_42486,N_41255,N_41198);
or U42487 (N_42487,N_40809,N_40194);
nor U42488 (N_42488,N_40571,N_40703);
nor U42489 (N_42489,N_40361,N_41627);
or U42490 (N_42490,N_41760,N_40818);
or U42491 (N_42491,N_41603,N_40138);
and U42492 (N_42492,N_41963,N_40055);
or U42493 (N_42493,N_41515,N_40012);
nor U42494 (N_42494,N_41005,N_40813);
and U42495 (N_42495,N_41141,N_40494);
or U42496 (N_42496,N_41217,N_41027);
nor U42497 (N_42497,N_40812,N_40767);
nor U42498 (N_42498,N_40856,N_40676);
nand U42499 (N_42499,N_40251,N_41061);
nand U42500 (N_42500,N_41695,N_41319);
xnor U42501 (N_42501,N_41962,N_41943);
and U42502 (N_42502,N_40021,N_40516);
xnor U42503 (N_42503,N_41238,N_40897);
or U42504 (N_42504,N_40257,N_40759);
or U42505 (N_42505,N_40011,N_40128);
and U42506 (N_42506,N_41778,N_41841);
xor U42507 (N_42507,N_40569,N_40682);
nor U42508 (N_42508,N_41958,N_41234);
xnor U42509 (N_42509,N_41804,N_41151);
nand U42510 (N_42510,N_40841,N_41537);
xor U42511 (N_42511,N_40472,N_41696);
nand U42512 (N_42512,N_41906,N_41593);
nand U42513 (N_42513,N_40821,N_41540);
xnor U42514 (N_42514,N_40745,N_40895);
nor U42515 (N_42515,N_41137,N_40770);
nor U42516 (N_42516,N_40353,N_40154);
nand U42517 (N_42517,N_41113,N_41193);
or U42518 (N_42518,N_41751,N_41355);
or U42519 (N_42519,N_40959,N_41551);
nand U42520 (N_42520,N_40638,N_41032);
xnor U42521 (N_42521,N_41503,N_41578);
xnor U42522 (N_42522,N_40114,N_41034);
or U42523 (N_42523,N_41535,N_40673);
nand U42524 (N_42524,N_41333,N_41404);
xor U42525 (N_42525,N_41376,N_40416);
nor U42526 (N_42526,N_41635,N_40524);
nor U42527 (N_42527,N_41419,N_40347);
nand U42528 (N_42528,N_41905,N_40850);
and U42529 (N_42529,N_40548,N_41935);
and U42530 (N_42530,N_40402,N_41925);
xnor U42531 (N_42531,N_41328,N_40977);
xor U42532 (N_42532,N_40074,N_41694);
or U42533 (N_42533,N_40626,N_40855);
nor U42534 (N_42534,N_40615,N_40849);
nand U42535 (N_42535,N_40368,N_40611);
or U42536 (N_42536,N_40530,N_40164);
or U42537 (N_42537,N_41014,N_40240);
and U42538 (N_42538,N_40827,N_41129);
and U42539 (N_42539,N_41463,N_40561);
or U42540 (N_42540,N_40669,N_40389);
nor U42541 (N_42541,N_40711,N_41916);
nor U42542 (N_42542,N_41341,N_40448);
or U42543 (N_42543,N_41051,N_40403);
and U42544 (N_42544,N_41154,N_41777);
or U42545 (N_42545,N_40018,N_41591);
nand U42546 (N_42546,N_40660,N_41029);
or U42547 (N_42547,N_40804,N_41186);
and U42548 (N_42548,N_40412,N_40398);
and U42549 (N_42549,N_41451,N_40989);
xnor U42550 (N_42550,N_41868,N_40900);
nor U42551 (N_42551,N_40140,N_41063);
nand U42552 (N_42552,N_40512,N_41431);
xnor U42553 (N_42553,N_40426,N_41507);
and U42554 (N_42554,N_40993,N_41145);
nor U42555 (N_42555,N_41062,N_41813);
and U42556 (N_42556,N_40326,N_40971);
nor U42557 (N_42557,N_41069,N_40831);
xor U42558 (N_42558,N_40994,N_41534);
and U42559 (N_42559,N_41090,N_41794);
or U42560 (N_42560,N_40734,N_40493);
nor U42561 (N_42561,N_41546,N_41498);
nor U42562 (N_42562,N_41030,N_41885);
or U42563 (N_42563,N_40726,N_40631);
nor U42564 (N_42564,N_40143,N_40242);
nand U42565 (N_42565,N_40371,N_40666);
and U42566 (N_42566,N_40567,N_40854);
nor U42567 (N_42567,N_41924,N_41629);
nor U42568 (N_42568,N_40097,N_41439);
nor U42569 (N_42569,N_40270,N_41406);
xor U42570 (N_42570,N_40252,N_41312);
nor U42571 (N_42571,N_41912,N_40168);
or U42572 (N_42572,N_40474,N_40700);
nor U42573 (N_42573,N_41742,N_41396);
nand U42574 (N_42574,N_41594,N_40724);
and U42575 (N_42575,N_40191,N_40651);
nor U42576 (N_42576,N_41698,N_40036);
and U42577 (N_42577,N_41210,N_41892);
nor U42578 (N_42578,N_41575,N_41582);
nand U42579 (N_42579,N_40133,N_40118);
xnor U42580 (N_42580,N_40953,N_41365);
xnor U42581 (N_42581,N_41511,N_40226);
nor U42582 (N_42582,N_40879,N_40190);
and U42583 (N_42583,N_40481,N_40945);
or U42584 (N_42584,N_40990,N_41676);
xnor U42585 (N_42585,N_40122,N_41973);
nand U42586 (N_42586,N_40784,N_40112);
xnor U42587 (N_42587,N_41244,N_41762);
xor U42588 (N_42588,N_40657,N_40769);
and U42589 (N_42589,N_40744,N_40513);
and U42590 (N_42590,N_41287,N_40933);
nand U42591 (N_42591,N_41659,N_40667);
nand U42592 (N_42592,N_40428,N_40201);
xnor U42593 (N_42593,N_41941,N_41240);
nor U42594 (N_42594,N_40550,N_40280);
xor U42595 (N_42595,N_40709,N_41491);
nor U42596 (N_42596,N_40040,N_40116);
or U42597 (N_42597,N_41280,N_40533);
nor U42598 (N_42598,N_40045,N_41583);
and U42599 (N_42599,N_41898,N_40941);
or U42600 (N_42600,N_41967,N_41125);
nand U42601 (N_42601,N_40032,N_41806);
or U42602 (N_42602,N_40385,N_40246);
nand U42603 (N_42603,N_41411,N_40159);
or U42604 (N_42604,N_40184,N_41204);
xnor U42605 (N_42605,N_41324,N_41142);
or U42606 (N_42606,N_40298,N_40678);
nor U42607 (N_42607,N_41615,N_40738);
and U42608 (N_42608,N_41607,N_41520);
nor U42609 (N_42609,N_40857,N_40539);
or U42610 (N_42610,N_41881,N_40090);
and U42611 (N_42611,N_40966,N_40048);
or U42612 (N_42612,N_40537,N_40681);
xor U42613 (N_42613,N_41385,N_41642);
or U42614 (N_42614,N_41378,N_41657);
nand U42615 (N_42615,N_40405,N_41746);
nand U42616 (N_42616,N_40917,N_40491);
or U42617 (N_42617,N_41849,N_41735);
or U42618 (N_42618,N_40316,N_41195);
xor U42619 (N_42619,N_41586,N_41316);
xor U42620 (N_42620,N_41780,N_40485);
nor U42621 (N_42621,N_41249,N_40230);
nand U42622 (N_42622,N_41863,N_41041);
nand U42623 (N_42623,N_40551,N_41665);
and U42624 (N_42624,N_41679,N_40912);
nor U42625 (N_42625,N_41454,N_41391);
nand U42626 (N_42626,N_41225,N_41831);
nor U42627 (N_42627,N_40186,N_40883);
and U42628 (N_42628,N_40228,N_41604);
nor U42629 (N_42629,N_41102,N_40451);
or U42630 (N_42630,N_41230,N_40483);
xor U42631 (N_42631,N_41455,N_41127);
nand U42632 (N_42632,N_40608,N_40136);
and U42633 (N_42633,N_41056,N_40271);
nand U42634 (N_42634,N_41825,N_40892);
nand U42635 (N_42635,N_41616,N_41284);
nand U42636 (N_42636,N_41854,N_40674);
xnor U42637 (N_42637,N_40477,N_40068);
nand U42638 (N_42638,N_40182,N_40504);
or U42639 (N_42639,N_41099,N_41372);
and U42640 (N_42640,N_40340,N_41309);
or U42641 (N_42641,N_41073,N_41630);
and U42642 (N_42642,N_40733,N_40600);
nor U42643 (N_42643,N_40878,N_41456);
xor U42644 (N_42644,N_41206,N_41784);
or U42645 (N_42645,N_41019,N_41123);
and U42646 (N_42646,N_41457,N_40965);
nand U42647 (N_42647,N_40282,N_41382);
xnor U42648 (N_42648,N_40735,N_40301);
nor U42649 (N_42649,N_40419,N_41260);
xnor U42650 (N_42650,N_41266,N_41052);
nor U42651 (N_42651,N_41543,N_40033);
nand U42652 (N_42652,N_40162,N_40324);
and U42653 (N_42653,N_41493,N_41880);
nor U42654 (N_42654,N_40613,N_40492);
or U42655 (N_42655,N_41150,N_41566);
nor U42656 (N_42656,N_41048,N_41522);
nor U42657 (N_42657,N_40737,N_40659);
xor U42658 (N_42658,N_41346,N_41538);
and U42659 (N_42659,N_40835,N_41972);
or U42660 (N_42660,N_41114,N_40098);
and U42661 (N_42661,N_41480,N_41111);
nor U42662 (N_42662,N_40432,N_40778);
nand U42663 (N_42663,N_41383,N_41815);
nor U42664 (N_42664,N_40973,N_40875);
xnor U42665 (N_42665,N_41800,N_40974);
or U42666 (N_42666,N_41213,N_40373);
nand U42667 (N_42667,N_40478,N_41856);
xnor U42668 (N_42668,N_41023,N_41119);
or U42669 (N_42669,N_41440,N_40345);
or U42670 (N_42670,N_40779,N_40645);
nand U42671 (N_42671,N_40570,N_41803);
or U42672 (N_42672,N_41315,N_41821);
and U42673 (N_42673,N_41572,N_40470);
xor U42674 (N_42674,N_40466,N_40691);
nor U42675 (N_42675,N_40675,N_41007);
and U42676 (N_42676,N_41460,N_41290);
nor U42677 (N_42677,N_41732,N_40786);
nand U42678 (N_42678,N_41650,N_40858);
and U42679 (N_42679,N_41373,N_41772);
nor U42680 (N_42680,N_40110,N_41458);
or U42681 (N_42681,N_40255,N_40757);
xor U42682 (N_42682,N_40987,N_41138);
nand U42683 (N_42683,N_40142,N_40196);
or U42684 (N_42684,N_40020,N_40266);
and U42685 (N_42685,N_40024,N_41037);
and U42686 (N_42686,N_41289,N_41474);
nand U42687 (N_42687,N_40046,N_40642);
xor U42688 (N_42688,N_40071,N_41921);
nand U42689 (N_42689,N_40215,N_41808);
nand U42690 (N_42690,N_40967,N_40147);
or U42691 (N_42691,N_40487,N_41375);
nand U42692 (N_42692,N_40554,N_41786);
nand U42693 (N_42693,N_40248,N_40449);
nand U42694 (N_42694,N_40245,N_40644);
and U42695 (N_42695,N_40077,N_40346);
or U42696 (N_42696,N_41595,N_41724);
or U42697 (N_42697,N_40844,N_40848);
and U42698 (N_42698,N_41645,N_41106);
and U42699 (N_42699,N_41639,N_41221);
xnor U42700 (N_42700,N_41079,N_41998);
or U42701 (N_42701,N_41395,N_40473);
xor U42702 (N_42702,N_40916,N_40216);
xor U42703 (N_42703,N_40931,N_41859);
or U42704 (N_42704,N_41261,N_41908);
xor U42705 (N_42705,N_40023,N_40665);
nand U42706 (N_42706,N_40558,N_41968);
nor U42707 (N_42707,N_41542,N_41573);
nand U42708 (N_42708,N_40899,N_40070);
nand U42709 (N_42709,N_41797,N_41686);
xor U42710 (N_42710,N_40108,N_40349);
nor U42711 (N_42711,N_40747,N_40865);
and U42712 (N_42712,N_41727,N_41837);
nor U42713 (N_42713,N_41486,N_41368);
and U42714 (N_42714,N_40207,N_41466);
or U42715 (N_42715,N_41560,N_41974);
xor U42716 (N_42716,N_40863,N_40026);
or U42717 (N_42717,N_41058,N_41465);
or U42718 (N_42718,N_40798,N_40092);
nand U42719 (N_42719,N_41323,N_41563);
nor U42720 (N_42720,N_40096,N_41366);
and U42721 (N_42721,N_41053,N_41693);
nor U42722 (N_42722,N_40409,N_40730);
nand U42723 (N_42723,N_40590,N_40891);
and U42724 (N_42724,N_40870,N_41283);
or U42725 (N_42725,N_40739,N_41623);
and U42726 (N_42726,N_40322,N_41201);
nor U42727 (N_42727,N_41605,N_40721);
nand U42728 (N_42728,N_40429,N_41737);
and U42729 (N_42729,N_40599,N_40387);
and U42730 (N_42730,N_41717,N_41237);
xnor U42731 (N_42731,N_41891,N_40095);
xnor U42732 (N_42732,N_40192,N_40632);
or U42733 (N_42733,N_40825,N_40585);
and U42734 (N_42734,N_41765,N_41739);
or U42735 (N_42735,N_41641,N_41691);
or U42736 (N_42736,N_40421,N_41178);
and U42737 (N_42737,N_41983,N_40287);
nor U42738 (N_42738,N_41293,N_41412);
or U42739 (N_42739,N_40643,N_40785);
and U42740 (N_42740,N_41116,N_41937);
xnor U42741 (N_42741,N_40067,N_41817);
and U42742 (N_42742,N_41415,N_40636);
and U42743 (N_42743,N_41409,N_41181);
nand U42744 (N_42744,N_41812,N_41352);
and U42745 (N_42745,N_40791,N_40288);
and U42746 (N_42746,N_40236,N_41938);
nand U42747 (N_42747,N_41464,N_40654);
nand U42748 (N_42748,N_40461,N_41861);
xnor U42749 (N_42749,N_40016,N_40102);
or U42750 (N_42750,N_41956,N_41702);
xor U42751 (N_42751,N_40640,N_40486);
or U42752 (N_42752,N_40135,N_41338);
xnor U42753 (N_42753,N_40909,N_40440);
or U42754 (N_42754,N_41756,N_40756);
nand U42755 (N_42755,N_40170,N_40000);
nand U42756 (N_42756,N_41163,N_41942);
nand U42757 (N_42757,N_41873,N_41229);
xor U42758 (N_42758,N_40031,N_41525);
and U42759 (N_42759,N_40355,N_40604);
nor U42760 (N_42760,N_41194,N_41310);
nand U42761 (N_42761,N_40934,N_41939);
and U42762 (N_42762,N_41934,N_41570);
and U42763 (N_42763,N_41401,N_40464);
xor U42764 (N_42764,N_40220,N_40277);
nand U42765 (N_42765,N_41243,N_41033);
or U42766 (N_42766,N_40383,N_41042);
xnor U42767 (N_42767,N_41897,N_41680);
nand U42768 (N_42768,N_41768,N_40795);
or U42769 (N_42769,N_41235,N_41530);
or U42770 (N_42770,N_41059,N_41297);
xnor U42771 (N_42771,N_41389,N_41197);
nand U42772 (N_42772,N_40393,N_41855);
xnor U42773 (N_42773,N_40859,N_41397);
or U42774 (N_42774,N_40983,N_40495);
xor U42775 (N_42775,N_40843,N_40343);
nand U42776 (N_42776,N_40049,N_40507);
xor U42777 (N_42777,N_41239,N_40921);
nor U42778 (N_42778,N_40597,N_41185);
xor U42779 (N_42779,N_40276,N_41568);
or U42780 (N_42780,N_40922,N_41878);
nand U42781 (N_42781,N_40806,N_40279);
nand U42782 (N_42782,N_41483,N_41386);
nor U42783 (N_42783,N_40460,N_40479);
nor U42784 (N_42784,N_41103,N_41248);
nor U42785 (N_42785,N_41561,N_41330);
or U42786 (N_42786,N_40760,N_40766);
or U42787 (N_42787,N_40452,N_40320);
xor U42788 (N_42788,N_40027,N_40352);
xor U42789 (N_42789,N_40195,N_41895);
and U42790 (N_42790,N_40714,N_41871);
nor U42791 (N_42791,N_40062,N_40212);
or U42792 (N_42792,N_41684,N_40851);
xnor U42793 (N_42793,N_41357,N_41608);
or U42794 (N_42794,N_41035,N_40132);
nand U42795 (N_42795,N_40041,N_41589);
and U42796 (N_42796,N_40520,N_41814);
and U42797 (N_42797,N_40911,N_41026);
nand U42798 (N_42798,N_40302,N_41285);
nor U42799 (N_42799,N_41184,N_41567);
nand U42800 (N_42800,N_41887,N_41931);
nor U42801 (N_42801,N_40283,N_40178);
or U42802 (N_42802,N_40789,N_41080);
nor U42803 (N_42803,N_41689,N_40995);
nor U42804 (N_42804,N_41381,N_41223);
nand U42805 (N_42805,N_40774,N_40447);
and U42806 (N_42806,N_41108,N_40115);
nand U42807 (N_42807,N_41770,N_41437);
or U42808 (N_42808,N_41281,N_40082);
and U42809 (N_42809,N_41955,N_41216);
or U42810 (N_42810,N_40274,N_41298);
nor U42811 (N_42811,N_41025,N_40017);
and U42812 (N_42812,N_41796,N_41047);
and U42813 (N_42813,N_41845,N_41236);
and U42814 (N_42814,N_41622,N_41867);
nor U42815 (N_42815,N_40940,N_40877);
nor U42816 (N_42816,N_40014,N_40445);
xor U42817 (N_42817,N_40227,N_41819);
nand U42818 (N_42818,N_41200,N_40152);
and U42819 (N_42819,N_40365,N_41140);
xnor U42820 (N_42820,N_41484,N_41721);
xnor U42821 (N_42821,N_41919,N_41112);
and U42822 (N_42822,N_40580,N_41990);
nor U42823 (N_42823,N_40241,N_41734);
xor U42824 (N_42824,N_41720,N_40101);
xnor U42825 (N_42825,N_41478,N_40716);
xnor U42826 (N_42826,N_40506,N_41167);
xnor U42827 (N_42827,N_41169,N_40621);
nor U42828 (N_42828,N_41325,N_41790);
xnor U42829 (N_42829,N_41485,N_40160);
or U42830 (N_42830,N_41711,N_41139);
nor U42831 (N_42831,N_40801,N_41758);
nor U42832 (N_42832,N_40817,N_40203);
and U42833 (N_42833,N_40508,N_41783);
or U42834 (N_42834,N_40437,N_40359);
or U42835 (N_42835,N_40193,N_40547);
xor U42836 (N_42836,N_40153,N_40086);
nor U42837 (N_42837,N_41769,N_41117);
or U42838 (N_42838,N_41969,N_40311);
nor U42839 (N_42839,N_41705,N_40229);
nand U42840 (N_42840,N_41651,N_40732);
and U42841 (N_42841,N_40124,N_41057);
nand U42842 (N_42842,N_40488,N_41598);
nand U42843 (N_42843,N_40439,N_41487);
nor U42844 (N_42844,N_41425,N_40509);
nor U42845 (N_42845,N_40148,N_41500);
xor U42846 (N_42846,N_41469,N_41896);
nor U42847 (N_42847,N_41453,N_40131);
nand U42848 (N_42848,N_40874,N_40291);
and U42849 (N_42849,N_41331,N_41055);
nor U42850 (N_42850,N_40871,N_40562);
nor U42851 (N_42851,N_40652,N_41360);
and U42852 (N_42852,N_40731,N_41174);
nand U42853 (N_42853,N_40459,N_40264);
and U42854 (N_42854,N_41094,N_41901);
xnor U42855 (N_42855,N_40751,N_40828);
xnor U42856 (N_42856,N_40754,N_40592);
and U42857 (N_42857,N_41313,N_41940);
xor U42858 (N_42858,N_41274,N_41647);
or U42859 (N_42859,N_40963,N_41273);
nand U42860 (N_42860,N_41010,N_41600);
nor U42861 (N_42861,N_40566,N_41894);
nand U42862 (N_42862,N_41002,N_40584);
nand U42863 (N_42863,N_41468,N_40173);
and U42864 (N_42864,N_40208,N_40761);
or U42865 (N_42865,N_40905,N_40904);
nor U42866 (N_42866,N_41086,N_40932);
or U42867 (N_42867,N_41359,N_40278);
nor U42868 (N_42868,N_41987,N_40338);
xnor U42869 (N_42869,N_41729,N_40656);
nor U42870 (N_42870,N_41084,N_41153);
nand U42871 (N_42871,N_41638,N_41707);
nand U42872 (N_42872,N_41417,N_40670);
nand U42873 (N_42873,N_40887,N_40471);
nor U42874 (N_42874,N_40038,N_41390);
nor U42875 (N_42875,N_40833,N_41886);
or U42876 (N_42876,N_40782,N_40499);
xor U42877 (N_42877,N_40702,N_41621);
or U42878 (N_42878,N_40523,N_40418);
and U42879 (N_42879,N_41054,N_41226);
and U42880 (N_42880,N_40219,N_40690);
xor U42881 (N_42881,N_41161,N_41259);
xnor U42882 (N_42882,N_40258,N_41740);
xor U42883 (N_42883,N_41791,N_40165);
and U42884 (N_42884,N_40622,N_41155);
or U42885 (N_42885,N_41846,N_41890);
nand U42886 (N_42886,N_40950,N_41091);
nand U42887 (N_42887,N_40910,N_40998);
nand U42888 (N_42888,N_40736,N_41170);
nor U42889 (N_42889,N_41565,N_40129);
xnor U42890 (N_42890,N_41536,N_41544);
nor U42891 (N_42891,N_41296,N_40677);
nand U42892 (N_42892,N_40810,N_41430);
nand U42893 (N_42893,N_40438,N_41753);
nand U42894 (N_42894,N_41512,N_41318);
xnor U42895 (N_42895,N_41173,N_40992);
xor U42896 (N_42896,N_40183,N_41580);
xor U42897 (N_42897,N_40465,N_41039);
or U42898 (N_42898,N_41932,N_40710);
xnor U42899 (N_42899,N_41467,N_40414);
and U42900 (N_42900,N_41426,N_41214);
nor U42901 (N_42901,N_40510,N_40202);
or U42902 (N_42902,N_41083,N_40999);
xnor U42903 (N_42903,N_41443,N_40200);
nand U42904 (N_42904,N_41736,N_40307);
or U42905 (N_42905,N_40976,N_41704);
nand U42906 (N_42906,N_40369,N_41268);
or U42907 (N_42907,N_40723,N_40860);
nand U42908 (N_42908,N_41982,N_40002);
xnor U42909 (N_42909,N_41836,N_40689);
xnor U42910 (N_42910,N_41569,N_41579);
and U42911 (N_42911,N_40357,N_40397);
or U42912 (N_42912,N_41715,N_41667);
and U42913 (N_42913,N_40901,N_40469);
or U42914 (N_42914,N_41311,N_41085);
or U42915 (N_42915,N_40684,N_41961);
nand U42916 (N_42916,N_41833,N_41219);
nor U42917 (N_42917,N_40386,N_40339);
and U42918 (N_42918,N_41043,N_41860);
nor U42919 (N_42919,N_41349,N_40748);
or U42920 (N_42920,N_41065,N_41461);
and U42921 (N_42921,N_40540,N_40886);
nand U42922 (N_42922,N_41000,N_40713);
nor U42923 (N_42923,N_40489,N_41432);
or U42924 (N_42924,N_40889,N_41636);
xnor U42925 (N_42925,N_41450,N_40705);
or U42926 (N_42926,N_41632,N_40925);
and U42927 (N_42927,N_40996,N_40955);
and U42928 (N_42928,N_40557,N_41851);
xor U42929 (N_42929,N_40306,N_41596);
nor U42930 (N_42930,N_41133,N_41022);
and U42931 (N_42931,N_41692,N_41725);
or U42932 (N_42932,N_41792,N_41664);
xnor U42933 (N_42933,N_40862,N_41547);
nand U42934 (N_42934,N_40842,N_41344);
nor U42935 (N_42935,N_40947,N_41723);
or U42936 (N_42936,N_40811,N_40704);
xnor U42937 (N_42937,N_41966,N_41946);
and U42938 (N_42938,N_40783,N_41364);
and U42939 (N_42939,N_40037,N_41674);
nand U42940 (N_42940,N_41046,N_40415);
and U42941 (N_42941,N_40117,N_40374);
and U42942 (N_42942,N_41189,N_41951);
xnor U42943 (N_42943,N_40559,N_40938);
nor U42944 (N_42944,N_40408,N_40728);
or U42945 (N_42945,N_40305,N_40417);
and U42946 (N_42946,N_41442,N_40475);
xor U42947 (N_42947,N_40893,N_40126);
nor U42948 (N_42948,N_40988,N_41830);
and U42949 (N_42949,N_40209,N_40261);
nand U42950 (N_42950,N_40013,N_40141);
nor U42951 (N_42951,N_40367,N_41581);
and U42952 (N_42952,N_40342,N_41745);
xnor U42953 (N_42953,N_40042,N_41918);
or U42954 (N_42954,N_40001,N_40272);
xnor U42955 (N_42955,N_40144,N_40595);
nand U42956 (N_42956,N_40560,N_41300);
xnor U42957 (N_42957,N_41436,N_40009);
nand U42958 (N_42958,N_40003,N_41070);
or U42959 (N_42959,N_40260,N_41889);
or U42960 (N_42960,N_41677,N_40157);
nor U42961 (N_42961,N_40861,N_41532);
nand U42962 (N_42962,N_40337,N_41922);
and U42963 (N_42963,N_41471,N_41508);
or U42964 (N_42964,N_40519,N_40926);
nor U42965 (N_42965,N_41272,N_40680);
xor U42966 (N_42966,N_40330,N_40617);
or U42967 (N_42967,N_40796,N_40204);
xnor U42968 (N_42968,N_41557,N_40820);
and U42969 (N_42969,N_40083,N_41767);
nand U42970 (N_42970,N_41611,N_40936);
xor U42971 (N_42971,N_40777,N_41759);
nor U42972 (N_42972,N_41190,N_41089);
nor U42973 (N_42973,N_40583,N_40185);
nor U42974 (N_42974,N_40982,N_41681);
or U42975 (N_42975,N_41548,N_40391);
xnor U42976 (N_42976,N_40577,N_41828);
xnor U42977 (N_42977,N_41713,N_40502);
nand U42978 (N_42978,N_40079,N_40589);
xor U42979 (N_42979,N_41763,N_40217);
nor U42980 (N_42980,N_41292,N_40741);
nand U42981 (N_42981,N_40244,N_41253);
or U42982 (N_42982,N_40211,N_41949);
and U42983 (N_42983,N_41857,N_41844);
and U42984 (N_42984,N_40591,N_41826);
and U42985 (N_42985,N_40807,N_40775);
xnor U42986 (N_42986,N_41655,N_41802);
nor U42987 (N_42987,N_41203,N_41307);
nand U42988 (N_42988,N_40423,N_41115);
nor U42989 (N_42989,N_40627,N_40740);
nor U42990 (N_42990,N_40100,N_40929);
nor U42991 (N_42991,N_40221,N_40243);
nand U42992 (N_42992,N_41428,N_40637);
and U42993 (N_42993,N_41212,N_41553);
nor U42994 (N_42994,N_41334,N_40454);
nor U42995 (N_42995,N_41158,N_41370);
nand U42996 (N_42996,N_40065,N_40952);
or U42997 (N_42997,N_41097,N_41348);
or U42998 (N_42998,N_41654,N_40123);
xor U42999 (N_42999,N_40697,N_41424);
nand U43000 (N_43000,N_41199,N_41924);
or U43001 (N_43001,N_40529,N_41297);
nor U43002 (N_43002,N_41136,N_41509);
or U43003 (N_43003,N_40827,N_40879);
or U43004 (N_43004,N_41652,N_41963);
xnor U43005 (N_43005,N_40089,N_40777);
and U43006 (N_43006,N_40474,N_41026);
or U43007 (N_43007,N_40785,N_41106);
nor U43008 (N_43008,N_41121,N_40459);
xnor U43009 (N_43009,N_41863,N_41338);
or U43010 (N_43010,N_41032,N_40395);
nor U43011 (N_43011,N_41358,N_40197);
nor U43012 (N_43012,N_40329,N_40191);
nor U43013 (N_43013,N_41175,N_41336);
and U43014 (N_43014,N_41591,N_41359);
nor U43015 (N_43015,N_40862,N_41788);
or U43016 (N_43016,N_41280,N_40185);
or U43017 (N_43017,N_41838,N_41680);
or U43018 (N_43018,N_41909,N_41851);
xnor U43019 (N_43019,N_41315,N_41090);
xnor U43020 (N_43020,N_40061,N_40736);
and U43021 (N_43021,N_40465,N_41088);
xor U43022 (N_43022,N_41525,N_40775);
nor U43023 (N_43023,N_40592,N_41645);
or U43024 (N_43024,N_41986,N_40812);
or U43025 (N_43025,N_41289,N_40882);
xnor U43026 (N_43026,N_40965,N_41596);
xnor U43027 (N_43027,N_41622,N_40467);
and U43028 (N_43028,N_41261,N_40618);
and U43029 (N_43029,N_40544,N_41314);
and U43030 (N_43030,N_40848,N_41461);
and U43031 (N_43031,N_41247,N_40260);
or U43032 (N_43032,N_40635,N_41186);
nand U43033 (N_43033,N_40165,N_40174);
nand U43034 (N_43034,N_41322,N_41536);
xor U43035 (N_43035,N_40613,N_40331);
or U43036 (N_43036,N_40560,N_40259);
nand U43037 (N_43037,N_41306,N_41922);
xnor U43038 (N_43038,N_41378,N_41688);
and U43039 (N_43039,N_40373,N_41227);
nand U43040 (N_43040,N_41748,N_41601);
xor U43041 (N_43041,N_40647,N_41267);
nand U43042 (N_43042,N_41228,N_40887);
or U43043 (N_43043,N_41464,N_40723);
nor U43044 (N_43044,N_40530,N_40697);
xor U43045 (N_43045,N_40425,N_41156);
nand U43046 (N_43046,N_40807,N_40383);
and U43047 (N_43047,N_41929,N_41300);
xor U43048 (N_43048,N_41122,N_41825);
or U43049 (N_43049,N_41773,N_40592);
or U43050 (N_43050,N_40753,N_41226);
and U43051 (N_43051,N_41918,N_40969);
or U43052 (N_43052,N_40777,N_41499);
and U43053 (N_43053,N_40901,N_41237);
nor U43054 (N_43054,N_41934,N_40006);
xnor U43055 (N_43055,N_41312,N_40753);
and U43056 (N_43056,N_40068,N_41904);
nor U43057 (N_43057,N_40914,N_40725);
nand U43058 (N_43058,N_41615,N_41351);
xnor U43059 (N_43059,N_40710,N_41412);
or U43060 (N_43060,N_40095,N_41203);
nand U43061 (N_43061,N_41622,N_41422);
nor U43062 (N_43062,N_40446,N_41957);
nor U43063 (N_43063,N_41095,N_41528);
and U43064 (N_43064,N_40590,N_41465);
and U43065 (N_43065,N_40900,N_40892);
or U43066 (N_43066,N_40597,N_40432);
nand U43067 (N_43067,N_40584,N_40702);
xor U43068 (N_43068,N_41552,N_41607);
nand U43069 (N_43069,N_40056,N_40852);
nand U43070 (N_43070,N_40552,N_40380);
and U43071 (N_43071,N_41057,N_41294);
and U43072 (N_43072,N_40481,N_41955);
nand U43073 (N_43073,N_41671,N_40434);
nor U43074 (N_43074,N_41702,N_40416);
xor U43075 (N_43075,N_40839,N_41148);
nand U43076 (N_43076,N_41054,N_40185);
or U43077 (N_43077,N_40633,N_41364);
or U43078 (N_43078,N_41970,N_41137);
or U43079 (N_43079,N_40669,N_41126);
nor U43080 (N_43080,N_41381,N_40314);
xor U43081 (N_43081,N_40069,N_40828);
or U43082 (N_43082,N_40571,N_41151);
nand U43083 (N_43083,N_40919,N_40579);
or U43084 (N_43084,N_41247,N_41353);
xor U43085 (N_43085,N_41441,N_41140);
or U43086 (N_43086,N_41275,N_41520);
and U43087 (N_43087,N_40445,N_40313);
and U43088 (N_43088,N_41997,N_41931);
nor U43089 (N_43089,N_41753,N_41298);
xor U43090 (N_43090,N_40123,N_41145);
nand U43091 (N_43091,N_40940,N_41756);
xor U43092 (N_43092,N_41630,N_40778);
or U43093 (N_43093,N_40793,N_41350);
or U43094 (N_43094,N_41070,N_41754);
nand U43095 (N_43095,N_40194,N_40472);
and U43096 (N_43096,N_40934,N_41258);
and U43097 (N_43097,N_40833,N_40447);
or U43098 (N_43098,N_41969,N_40701);
xnor U43099 (N_43099,N_41005,N_40344);
and U43100 (N_43100,N_41412,N_40959);
or U43101 (N_43101,N_40478,N_41770);
or U43102 (N_43102,N_40516,N_41431);
nor U43103 (N_43103,N_40655,N_41510);
or U43104 (N_43104,N_41562,N_41133);
nor U43105 (N_43105,N_40744,N_40644);
or U43106 (N_43106,N_40049,N_41317);
xnor U43107 (N_43107,N_41666,N_40231);
nand U43108 (N_43108,N_41815,N_41087);
and U43109 (N_43109,N_40537,N_40163);
nand U43110 (N_43110,N_40296,N_40447);
nor U43111 (N_43111,N_41027,N_40366);
or U43112 (N_43112,N_41834,N_40360);
xnor U43113 (N_43113,N_41499,N_40236);
or U43114 (N_43114,N_41344,N_41164);
xor U43115 (N_43115,N_40570,N_40095);
nor U43116 (N_43116,N_41619,N_41816);
nor U43117 (N_43117,N_41773,N_40199);
xnor U43118 (N_43118,N_41084,N_40042);
nand U43119 (N_43119,N_41515,N_41227);
or U43120 (N_43120,N_41955,N_41217);
or U43121 (N_43121,N_41230,N_40650);
or U43122 (N_43122,N_41108,N_40986);
nand U43123 (N_43123,N_40011,N_40802);
nand U43124 (N_43124,N_41804,N_40775);
or U43125 (N_43125,N_41080,N_40704);
nand U43126 (N_43126,N_40260,N_40063);
and U43127 (N_43127,N_40155,N_41561);
and U43128 (N_43128,N_41661,N_41710);
or U43129 (N_43129,N_41968,N_41236);
nand U43130 (N_43130,N_41061,N_40440);
or U43131 (N_43131,N_40959,N_41004);
nand U43132 (N_43132,N_40099,N_41803);
nand U43133 (N_43133,N_41801,N_41151);
or U43134 (N_43134,N_41083,N_41260);
nor U43135 (N_43135,N_41614,N_41606);
nand U43136 (N_43136,N_41073,N_41226);
nor U43137 (N_43137,N_41312,N_40774);
nor U43138 (N_43138,N_40154,N_41183);
xor U43139 (N_43139,N_40415,N_40703);
nor U43140 (N_43140,N_40483,N_40322);
nand U43141 (N_43141,N_40001,N_41610);
nor U43142 (N_43142,N_41633,N_41364);
nand U43143 (N_43143,N_40192,N_41616);
or U43144 (N_43144,N_40052,N_40130);
nor U43145 (N_43145,N_40602,N_40689);
nor U43146 (N_43146,N_41840,N_41520);
nand U43147 (N_43147,N_41668,N_41375);
nor U43148 (N_43148,N_41882,N_41250);
or U43149 (N_43149,N_41909,N_40949);
nor U43150 (N_43150,N_40266,N_41147);
nor U43151 (N_43151,N_40235,N_41260);
or U43152 (N_43152,N_41521,N_40888);
or U43153 (N_43153,N_40880,N_40955);
xnor U43154 (N_43154,N_40878,N_41500);
or U43155 (N_43155,N_41591,N_40711);
and U43156 (N_43156,N_40762,N_41999);
and U43157 (N_43157,N_40426,N_40897);
nor U43158 (N_43158,N_40305,N_40937);
nor U43159 (N_43159,N_40478,N_40313);
nor U43160 (N_43160,N_41090,N_40029);
xor U43161 (N_43161,N_40014,N_41104);
nand U43162 (N_43162,N_41820,N_41265);
nand U43163 (N_43163,N_41571,N_40387);
nand U43164 (N_43164,N_41932,N_41248);
nor U43165 (N_43165,N_41305,N_41316);
nand U43166 (N_43166,N_40717,N_41991);
and U43167 (N_43167,N_40133,N_40074);
and U43168 (N_43168,N_40188,N_40901);
nand U43169 (N_43169,N_40728,N_40168);
nand U43170 (N_43170,N_41621,N_41066);
or U43171 (N_43171,N_41050,N_41244);
nand U43172 (N_43172,N_41616,N_41965);
and U43173 (N_43173,N_41221,N_40909);
nor U43174 (N_43174,N_40421,N_40572);
or U43175 (N_43175,N_40633,N_40989);
nor U43176 (N_43176,N_40351,N_40484);
nor U43177 (N_43177,N_40755,N_40319);
and U43178 (N_43178,N_40751,N_40786);
and U43179 (N_43179,N_41994,N_40853);
nand U43180 (N_43180,N_40679,N_41091);
and U43181 (N_43181,N_40243,N_41838);
xnor U43182 (N_43182,N_41218,N_41576);
nand U43183 (N_43183,N_40037,N_40697);
and U43184 (N_43184,N_40082,N_41598);
xnor U43185 (N_43185,N_41940,N_40212);
nand U43186 (N_43186,N_40051,N_40448);
nand U43187 (N_43187,N_40430,N_41765);
or U43188 (N_43188,N_40255,N_40260);
nand U43189 (N_43189,N_40662,N_40248);
xnor U43190 (N_43190,N_40531,N_40847);
nor U43191 (N_43191,N_41774,N_40294);
and U43192 (N_43192,N_41773,N_41679);
and U43193 (N_43193,N_40191,N_41378);
xor U43194 (N_43194,N_41020,N_41976);
nand U43195 (N_43195,N_40205,N_41131);
nand U43196 (N_43196,N_41945,N_40112);
xor U43197 (N_43197,N_40202,N_41634);
nor U43198 (N_43198,N_41048,N_41748);
or U43199 (N_43199,N_40240,N_40057);
nor U43200 (N_43200,N_40902,N_40853);
nand U43201 (N_43201,N_41038,N_41677);
nand U43202 (N_43202,N_41551,N_41079);
and U43203 (N_43203,N_40203,N_41745);
or U43204 (N_43204,N_40273,N_40514);
or U43205 (N_43205,N_40246,N_40569);
xor U43206 (N_43206,N_41080,N_41226);
xor U43207 (N_43207,N_40017,N_41186);
or U43208 (N_43208,N_40810,N_40561);
nand U43209 (N_43209,N_41559,N_41609);
xor U43210 (N_43210,N_40382,N_40901);
and U43211 (N_43211,N_41039,N_40385);
nand U43212 (N_43212,N_41136,N_40570);
nand U43213 (N_43213,N_40576,N_41282);
or U43214 (N_43214,N_40861,N_40540);
nand U43215 (N_43215,N_41168,N_41178);
xor U43216 (N_43216,N_40039,N_41606);
or U43217 (N_43217,N_40348,N_41425);
and U43218 (N_43218,N_40710,N_40003);
xnor U43219 (N_43219,N_40877,N_40171);
nand U43220 (N_43220,N_40599,N_40778);
nor U43221 (N_43221,N_40969,N_41023);
nor U43222 (N_43222,N_41025,N_41163);
and U43223 (N_43223,N_40982,N_40428);
xor U43224 (N_43224,N_41256,N_40716);
nand U43225 (N_43225,N_40458,N_41996);
and U43226 (N_43226,N_40903,N_40106);
or U43227 (N_43227,N_40140,N_41018);
and U43228 (N_43228,N_41154,N_41895);
xor U43229 (N_43229,N_40741,N_41944);
xor U43230 (N_43230,N_41029,N_41803);
and U43231 (N_43231,N_41564,N_40226);
xor U43232 (N_43232,N_41466,N_41227);
xor U43233 (N_43233,N_40682,N_40995);
or U43234 (N_43234,N_41986,N_41593);
or U43235 (N_43235,N_40712,N_40177);
nand U43236 (N_43236,N_40852,N_40132);
and U43237 (N_43237,N_41283,N_40380);
and U43238 (N_43238,N_41038,N_40938);
nand U43239 (N_43239,N_41974,N_40604);
nand U43240 (N_43240,N_40343,N_41219);
nand U43241 (N_43241,N_40578,N_40819);
or U43242 (N_43242,N_41273,N_41781);
and U43243 (N_43243,N_41779,N_41026);
and U43244 (N_43244,N_41042,N_40774);
nor U43245 (N_43245,N_41717,N_40272);
xnor U43246 (N_43246,N_41187,N_41827);
xor U43247 (N_43247,N_40169,N_41069);
nor U43248 (N_43248,N_40199,N_40344);
xnor U43249 (N_43249,N_40642,N_41035);
and U43250 (N_43250,N_40739,N_40268);
nor U43251 (N_43251,N_40148,N_41683);
xnor U43252 (N_43252,N_41315,N_41993);
xor U43253 (N_43253,N_41242,N_41956);
and U43254 (N_43254,N_41921,N_41501);
xnor U43255 (N_43255,N_41744,N_40965);
nor U43256 (N_43256,N_41882,N_40063);
xnor U43257 (N_43257,N_40781,N_41151);
nand U43258 (N_43258,N_41306,N_40749);
nor U43259 (N_43259,N_40736,N_40859);
xor U43260 (N_43260,N_41316,N_41885);
nand U43261 (N_43261,N_40577,N_41532);
nand U43262 (N_43262,N_40107,N_41565);
or U43263 (N_43263,N_41534,N_41684);
nand U43264 (N_43264,N_41421,N_40569);
or U43265 (N_43265,N_40551,N_41781);
or U43266 (N_43266,N_41797,N_41127);
nand U43267 (N_43267,N_41630,N_40022);
xnor U43268 (N_43268,N_40003,N_40070);
nand U43269 (N_43269,N_41564,N_41918);
nand U43270 (N_43270,N_41765,N_40731);
and U43271 (N_43271,N_41615,N_41943);
nor U43272 (N_43272,N_40756,N_40855);
or U43273 (N_43273,N_41716,N_41126);
nand U43274 (N_43274,N_40408,N_40268);
nor U43275 (N_43275,N_41562,N_41613);
and U43276 (N_43276,N_41902,N_40191);
or U43277 (N_43277,N_41330,N_40245);
nand U43278 (N_43278,N_41704,N_40133);
and U43279 (N_43279,N_40412,N_40523);
or U43280 (N_43280,N_41656,N_41596);
nor U43281 (N_43281,N_40876,N_40907);
or U43282 (N_43282,N_40890,N_41850);
and U43283 (N_43283,N_40962,N_40050);
or U43284 (N_43284,N_40102,N_40216);
or U43285 (N_43285,N_41555,N_41161);
nand U43286 (N_43286,N_40734,N_41287);
nand U43287 (N_43287,N_40244,N_41125);
xor U43288 (N_43288,N_41729,N_40827);
nor U43289 (N_43289,N_41090,N_41696);
and U43290 (N_43290,N_41158,N_40737);
and U43291 (N_43291,N_41027,N_41677);
nand U43292 (N_43292,N_41037,N_41969);
xor U43293 (N_43293,N_40150,N_41651);
and U43294 (N_43294,N_40439,N_41439);
xor U43295 (N_43295,N_41684,N_41342);
xnor U43296 (N_43296,N_41073,N_41658);
xor U43297 (N_43297,N_40342,N_40549);
and U43298 (N_43298,N_41501,N_40030);
nand U43299 (N_43299,N_41980,N_41651);
xnor U43300 (N_43300,N_41226,N_40618);
and U43301 (N_43301,N_40635,N_40819);
or U43302 (N_43302,N_40638,N_40236);
nor U43303 (N_43303,N_41862,N_40597);
nand U43304 (N_43304,N_41860,N_40472);
or U43305 (N_43305,N_40066,N_41568);
or U43306 (N_43306,N_40299,N_40374);
nand U43307 (N_43307,N_40211,N_41005);
nand U43308 (N_43308,N_40081,N_41700);
and U43309 (N_43309,N_41106,N_41407);
nor U43310 (N_43310,N_41487,N_40372);
xnor U43311 (N_43311,N_40779,N_40966);
or U43312 (N_43312,N_40238,N_40389);
nand U43313 (N_43313,N_41200,N_40690);
nor U43314 (N_43314,N_41792,N_40945);
or U43315 (N_43315,N_41312,N_40883);
nand U43316 (N_43316,N_41528,N_41447);
xor U43317 (N_43317,N_41989,N_41948);
nand U43318 (N_43318,N_41495,N_40819);
xnor U43319 (N_43319,N_40900,N_41121);
nand U43320 (N_43320,N_41589,N_41504);
nor U43321 (N_43321,N_41381,N_41138);
nor U43322 (N_43322,N_41130,N_41604);
nor U43323 (N_43323,N_40057,N_41541);
xor U43324 (N_43324,N_41016,N_41224);
and U43325 (N_43325,N_40480,N_41946);
nand U43326 (N_43326,N_40739,N_41303);
and U43327 (N_43327,N_40763,N_41176);
nand U43328 (N_43328,N_41498,N_41478);
nor U43329 (N_43329,N_41383,N_40008);
or U43330 (N_43330,N_40607,N_41971);
nor U43331 (N_43331,N_40724,N_40560);
xnor U43332 (N_43332,N_41176,N_40868);
nor U43333 (N_43333,N_41096,N_40500);
and U43334 (N_43334,N_40551,N_41754);
nor U43335 (N_43335,N_40202,N_40658);
nand U43336 (N_43336,N_41533,N_40400);
and U43337 (N_43337,N_40294,N_41479);
xor U43338 (N_43338,N_40468,N_41982);
nand U43339 (N_43339,N_41958,N_41380);
or U43340 (N_43340,N_41090,N_41405);
or U43341 (N_43341,N_40204,N_40764);
or U43342 (N_43342,N_40773,N_40388);
or U43343 (N_43343,N_40896,N_41435);
or U43344 (N_43344,N_41241,N_40258);
or U43345 (N_43345,N_40681,N_40147);
nor U43346 (N_43346,N_41805,N_41799);
xnor U43347 (N_43347,N_40229,N_41816);
nor U43348 (N_43348,N_40929,N_41449);
and U43349 (N_43349,N_40444,N_41276);
and U43350 (N_43350,N_41019,N_40403);
nor U43351 (N_43351,N_41475,N_40025);
and U43352 (N_43352,N_41818,N_41895);
and U43353 (N_43353,N_41867,N_40949);
and U43354 (N_43354,N_41897,N_40898);
nand U43355 (N_43355,N_41717,N_41737);
nor U43356 (N_43356,N_40895,N_41135);
and U43357 (N_43357,N_41657,N_40424);
or U43358 (N_43358,N_40470,N_40225);
and U43359 (N_43359,N_41081,N_40984);
nand U43360 (N_43360,N_41600,N_41647);
xnor U43361 (N_43361,N_41229,N_41682);
xor U43362 (N_43362,N_40889,N_40416);
nor U43363 (N_43363,N_40813,N_40260);
nand U43364 (N_43364,N_41683,N_40822);
nor U43365 (N_43365,N_41641,N_41962);
or U43366 (N_43366,N_41521,N_40850);
nand U43367 (N_43367,N_41791,N_40512);
nand U43368 (N_43368,N_40378,N_41542);
and U43369 (N_43369,N_41068,N_41998);
nand U43370 (N_43370,N_40993,N_40345);
nand U43371 (N_43371,N_41437,N_40151);
or U43372 (N_43372,N_40959,N_40404);
and U43373 (N_43373,N_41099,N_41742);
or U43374 (N_43374,N_40408,N_41301);
xor U43375 (N_43375,N_40118,N_40201);
nand U43376 (N_43376,N_41755,N_40001);
and U43377 (N_43377,N_41270,N_40534);
nand U43378 (N_43378,N_41547,N_41141);
and U43379 (N_43379,N_40225,N_40342);
nor U43380 (N_43380,N_41550,N_41345);
or U43381 (N_43381,N_40645,N_41083);
xnor U43382 (N_43382,N_41293,N_40784);
xnor U43383 (N_43383,N_40322,N_41797);
and U43384 (N_43384,N_41266,N_41524);
nand U43385 (N_43385,N_41783,N_41378);
xor U43386 (N_43386,N_40176,N_41055);
and U43387 (N_43387,N_40963,N_41897);
or U43388 (N_43388,N_41693,N_40466);
nor U43389 (N_43389,N_41469,N_40538);
nand U43390 (N_43390,N_41922,N_41688);
xnor U43391 (N_43391,N_40867,N_41290);
and U43392 (N_43392,N_41353,N_40741);
and U43393 (N_43393,N_40340,N_41166);
or U43394 (N_43394,N_41390,N_41067);
xnor U43395 (N_43395,N_41618,N_40717);
nor U43396 (N_43396,N_40398,N_41541);
and U43397 (N_43397,N_40533,N_40136);
or U43398 (N_43398,N_41857,N_41632);
and U43399 (N_43399,N_40844,N_40443);
or U43400 (N_43400,N_41863,N_40470);
nor U43401 (N_43401,N_40200,N_40781);
and U43402 (N_43402,N_40835,N_40805);
nand U43403 (N_43403,N_40191,N_40576);
and U43404 (N_43404,N_41487,N_40930);
or U43405 (N_43405,N_41090,N_41957);
and U43406 (N_43406,N_41055,N_40875);
nand U43407 (N_43407,N_40083,N_41086);
or U43408 (N_43408,N_41507,N_40092);
nand U43409 (N_43409,N_41604,N_40412);
nand U43410 (N_43410,N_41828,N_40695);
nand U43411 (N_43411,N_40506,N_40309);
xor U43412 (N_43412,N_41420,N_40924);
nor U43413 (N_43413,N_41230,N_41250);
nand U43414 (N_43414,N_41596,N_40913);
or U43415 (N_43415,N_40549,N_40511);
and U43416 (N_43416,N_41083,N_41559);
and U43417 (N_43417,N_40453,N_40018);
nand U43418 (N_43418,N_41865,N_41841);
xor U43419 (N_43419,N_40604,N_41368);
nand U43420 (N_43420,N_41475,N_40856);
nor U43421 (N_43421,N_40869,N_41916);
nand U43422 (N_43422,N_41275,N_41610);
xnor U43423 (N_43423,N_41022,N_41369);
or U43424 (N_43424,N_40311,N_40659);
and U43425 (N_43425,N_40736,N_40166);
xor U43426 (N_43426,N_41045,N_41948);
nor U43427 (N_43427,N_40172,N_40950);
and U43428 (N_43428,N_41610,N_41488);
nand U43429 (N_43429,N_41544,N_41492);
nand U43430 (N_43430,N_40334,N_41963);
nor U43431 (N_43431,N_41692,N_41657);
or U43432 (N_43432,N_40306,N_40745);
nand U43433 (N_43433,N_41965,N_41909);
or U43434 (N_43434,N_40241,N_40221);
nor U43435 (N_43435,N_40120,N_41918);
nor U43436 (N_43436,N_41612,N_41843);
and U43437 (N_43437,N_40638,N_40095);
or U43438 (N_43438,N_41019,N_40127);
or U43439 (N_43439,N_40788,N_40383);
nor U43440 (N_43440,N_40008,N_40432);
nor U43441 (N_43441,N_40837,N_40716);
xor U43442 (N_43442,N_40901,N_41182);
and U43443 (N_43443,N_41842,N_40617);
nor U43444 (N_43444,N_41259,N_41181);
nand U43445 (N_43445,N_41704,N_41828);
and U43446 (N_43446,N_40156,N_40204);
or U43447 (N_43447,N_40751,N_41107);
nor U43448 (N_43448,N_40588,N_41674);
nor U43449 (N_43449,N_41993,N_41491);
or U43450 (N_43450,N_40834,N_41646);
or U43451 (N_43451,N_40166,N_41834);
or U43452 (N_43452,N_40480,N_40555);
nor U43453 (N_43453,N_40825,N_40930);
nand U43454 (N_43454,N_40622,N_41045);
nor U43455 (N_43455,N_41311,N_40636);
and U43456 (N_43456,N_40425,N_41264);
nor U43457 (N_43457,N_41988,N_40446);
xnor U43458 (N_43458,N_41686,N_40727);
and U43459 (N_43459,N_41875,N_41426);
or U43460 (N_43460,N_40416,N_41271);
nor U43461 (N_43461,N_41597,N_40268);
or U43462 (N_43462,N_41852,N_40033);
nor U43463 (N_43463,N_40509,N_40104);
and U43464 (N_43464,N_40912,N_40955);
xnor U43465 (N_43465,N_41185,N_41468);
and U43466 (N_43466,N_41681,N_41061);
and U43467 (N_43467,N_41100,N_41705);
xor U43468 (N_43468,N_41369,N_41558);
xnor U43469 (N_43469,N_41889,N_41022);
nand U43470 (N_43470,N_40940,N_41373);
nand U43471 (N_43471,N_40334,N_41696);
nand U43472 (N_43472,N_40409,N_41955);
xnor U43473 (N_43473,N_41130,N_41690);
or U43474 (N_43474,N_41091,N_40590);
nand U43475 (N_43475,N_40021,N_41555);
xor U43476 (N_43476,N_40100,N_40897);
and U43477 (N_43477,N_41355,N_41397);
xor U43478 (N_43478,N_41282,N_41983);
nand U43479 (N_43479,N_41178,N_41291);
or U43480 (N_43480,N_40785,N_40819);
or U43481 (N_43481,N_40979,N_41815);
or U43482 (N_43482,N_41277,N_41455);
and U43483 (N_43483,N_40108,N_40708);
nor U43484 (N_43484,N_41701,N_40885);
nor U43485 (N_43485,N_40157,N_41790);
nand U43486 (N_43486,N_40238,N_40563);
or U43487 (N_43487,N_40728,N_41781);
nor U43488 (N_43488,N_41858,N_40012);
xnor U43489 (N_43489,N_41463,N_40209);
and U43490 (N_43490,N_41584,N_41505);
and U43491 (N_43491,N_41946,N_41138);
nand U43492 (N_43492,N_40876,N_40979);
nor U43493 (N_43493,N_41331,N_41487);
xor U43494 (N_43494,N_40124,N_40265);
and U43495 (N_43495,N_40545,N_41932);
nand U43496 (N_43496,N_40575,N_41236);
xor U43497 (N_43497,N_40289,N_41612);
nand U43498 (N_43498,N_41685,N_40764);
and U43499 (N_43499,N_40265,N_41367);
or U43500 (N_43500,N_40480,N_41771);
nand U43501 (N_43501,N_40119,N_41975);
or U43502 (N_43502,N_41387,N_41717);
nand U43503 (N_43503,N_40193,N_41237);
or U43504 (N_43504,N_41683,N_40998);
nor U43505 (N_43505,N_41486,N_41367);
xor U43506 (N_43506,N_40335,N_40774);
and U43507 (N_43507,N_41196,N_40734);
nor U43508 (N_43508,N_40275,N_41986);
nand U43509 (N_43509,N_41852,N_40054);
or U43510 (N_43510,N_40237,N_41495);
xor U43511 (N_43511,N_40090,N_40862);
or U43512 (N_43512,N_41620,N_41961);
xnor U43513 (N_43513,N_40762,N_41177);
and U43514 (N_43514,N_40820,N_41896);
nand U43515 (N_43515,N_41026,N_41339);
and U43516 (N_43516,N_40804,N_40447);
or U43517 (N_43517,N_40279,N_40588);
nor U43518 (N_43518,N_41498,N_41042);
and U43519 (N_43519,N_41490,N_40606);
nand U43520 (N_43520,N_40948,N_40994);
and U43521 (N_43521,N_41878,N_40797);
or U43522 (N_43522,N_41779,N_41154);
and U43523 (N_43523,N_41800,N_40396);
nand U43524 (N_43524,N_41577,N_40409);
and U43525 (N_43525,N_40112,N_41556);
and U43526 (N_43526,N_40916,N_41836);
and U43527 (N_43527,N_41641,N_41984);
or U43528 (N_43528,N_41387,N_40600);
xor U43529 (N_43529,N_41342,N_40211);
xor U43530 (N_43530,N_41188,N_40349);
nand U43531 (N_43531,N_41534,N_40021);
or U43532 (N_43532,N_41396,N_40355);
nor U43533 (N_43533,N_41847,N_40413);
and U43534 (N_43534,N_41868,N_40315);
and U43535 (N_43535,N_41762,N_40226);
nand U43536 (N_43536,N_40678,N_40459);
nand U43537 (N_43537,N_40799,N_41689);
and U43538 (N_43538,N_41802,N_40921);
or U43539 (N_43539,N_41322,N_40648);
xor U43540 (N_43540,N_41293,N_40879);
nor U43541 (N_43541,N_41656,N_40134);
and U43542 (N_43542,N_40473,N_41788);
xor U43543 (N_43543,N_40760,N_40555);
nor U43544 (N_43544,N_41510,N_41530);
or U43545 (N_43545,N_41915,N_41231);
or U43546 (N_43546,N_40007,N_40047);
nand U43547 (N_43547,N_40494,N_40474);
nor U43548 (N_43548,N_41945,N_41501);
nor U43549 (N_43549,N_40405,N_41895);
or U43550 (N_43550,N_40459,N_40451);
or U43551 (N_43551,N_40371,N_41490);
nand U43552 (N_43552,N_41231,N_40394);
nand U43553 (N_43553,N_41409,N_41081);
nand U43554 (N_43554,N_41653,N_41363);
nor U43555 (N_43555,N_40957,N_40761);
and U43556 (N_43556,N_40999,N_40792);
nand U43557 (N_43557,N_41141,N_40865);
nand U43558 (N_43558,N_41121,N_40092);
xnor U43559 (N_43559,N_40376,N_41929);
xor U43560 (N_43560,N_41290,N_40699);
or U43561 (N_43561,N_40177,N_41675);
nand U43562 (N_43562,N_41421,N_40865);
or U43563 (N_43563,N_41482,N_41489);
xor U43564 (N_43564,N_40069,N_40755);
nand U43565 (N_43565,N_41452,N_40409);
and U43566 (N_43566,N_40627,N_41074);
xor U43567 (N_43567,N_40365,N_41032);
or U43568 (N_43568,N_41618,N_40058);
xor U43569 (N_43569,N_40658,N_40315);
or U43570 (N_43570,N_41022,N_41801);
nand U43571 (N_43571,N_40535,N_40113);
and U43572 (N_43572,N_40414,N_40545);
or U43573 (N_43573,N_41619,N_40219);
nand U43574 (N_43574,N_41195,N_41773);
nor U43575 (N_43575,N_40600,N_41424);
or U43576 (N_43576,N_41073,N_41405);
or U43577 (N_43577,N_41918,N_40503);
xnor U43578 (N_43578,N_41600,N_41369);
nor U43579 (N_43579,N_40474,N_41621);
xnor U43580 (N_43580,N_40882,N_40144);
xor U43581 (N_43581,N_41153,N_41591);
and U43582 (N_43582,N_41740,N_41128);
and U43583 (N_43583,N_40676,N_41401);
xor U43584 (N_43584,N_41636,N_40930);
and U43585 (N_43585,N_41396,N_41991);
nand U43586 (N_43586,N_40338,N_41524);
nor U43587 (N_43587,N_40826,N_41889);
or U43588 (N_43588,N_40745,N_40451);
and U43589 (N_43589,N_40614,N_41306);
and U43590 (N_43590,N_40049,N_41290);
nand U43591 (N_43591,N_40127,N_40875);
nand U43592 (N_43592,N_40676,N_41263);
nor U43593 (N_43593,N_41008,N_40231);
or U43594 (N_43594,N_41183,N_41522);
and U43595 (N_43595,N_40717,N_40899);
xnor U43596 (N_43596,N_41388,N_40154);
nor U43597 (N_43597,N_40817,N_40773);
and U43598 (N_43598,N_40061,N_40263);
xor U43599 (N_43599,N_41790,N_40476);
xnor U43600 (N_43600,N_40684,N_40040);
and U43601 (N_43601,N_40491,N_41522);
or U43602 (N_43602,N_40750,N_41013);
nor U43603 (N_43603,N_40290,N_40461);
xnor U43604 (N_43604,N_41132,N_40317);
nand U43605 (N_43605,N_41909,N_41035);
xnor U43606 (N_43606,N_41091,N_41605);
nor U43607 (N_43607,N_40422,N_41382);
xor U43608 (N_43608,N_41833,N_41394);
nor U43609 (N_43609,N_41267,N_41336);
or U43610 (N_43610,N_40056,N_40386);
nand U43611 (N_43611,N_41349,N_40471);
nor U43612 (N_43612,N_40748,N_40219);
nor U43613 (N_43613,N_41447,N_41115);
xnor U43614 (N_43614,N_41800,N_41827);
and U43615 (N_43615,N_41478,N_40668);
nor U43616 (N_43616,N_41240,N_41004);
nor U43617 (N_43617,N_41536,N_40355);
nand U43618 (N_43618,N_41034,N_40219);
or U43619 (N_43619,N_41224,N_41060);
and U43620 (N_43620,N_40866,N_41041);
nand U43621 (N_43621,N_41204,N_40226);
or U43622 (N_43622,N_40219,N_41347);
nand U43623 (N_43623,N_40635,N_40672);
xor U43624 (N_43624,N_41667,N_40780);
and U43625 (N_43625,N_40616,N_40048);
or U43626 (N_43626,N_41129,N_41284);
or U43627 (N_43627,N_41991,N_41569);
nand U43628 (N_43628,N_41387,N_40923);
xnor U43629 (N_43629,N_40007,N_41290);
or U43630 (N_43630,N_40123,N_41038);
xnor U43631 (N_43631,N_40960,N_41221);
and U43632 (N_43632,N_41585,N_41425);
xnor U43633 (N_43633,N_41719,N_40235);
xnor U43634 (N_43634,N_40191,N_40677);
or U43635 (N_43635,N_41505,N_41515);
xnor U43636 (N_43636,N_40277,N_41659);
xnor U43637 (N_43637,N_41618,N_40359);
and U43638 (N_43638,N_41025,N_40369);
xnor U43639 (N_43639,N_41355,N_40352);
or U43640 (N_43640,N_41401,N_40367);
xor U43641 (N_43641,N_40024,N_41161);
xor U43642 (N_43642,N_41666,N_40275);
and U43643 (N_43643,N_40251,N_40093);
or U43644 (N_43644,N_41387,N_40231);
or U43645 (N_43645,N_40856,N_40422);
nor U43646 (N_43646,N_40570,N_40446);
and U43647 (N_43647,N_40124,N_40442);
nand U43648 (N_43648,N_40804,N_41786);
or U43649 (N_43649,N_40463,N_40061);
xor U43650 (N_43650,N_41270,N_40418);
xor U43651 (N_43651,N_40342,N_41654);
or U43652 (N_43652,N_41899,N_40139);
and U43653 (N_43653,N_41980,N_41455);
nor U43654 (N_43654,N_40040,N_41814);
or U43655 (N_43655,N_41284,N_41558);
nor U43656 (N_43656,N_41996,N_41288);
nor U43657 (N_43657,N_40033,N_41046);
and U43658 (N_43658,N_40347,N_40797);
nand U43659 (N_43659,N_41797,N_41920);
nor U43660 (N_43660,N_40359,N_41779);
or U43661 (N_43661,N_40991,N_40408);
or U43662 (N_43662,N_41766,N_41276);
xor U43663 (N_43663,N_40404,N_40517);
nand U43664 (N_43664,N_41359,N_40290);
or U43665 (N_43665,N_41120,N_41543);
and U43666 (N_43666,N_40308,N_41841);
or U43667 (N_43667,N_41037,N_40161);
or U43668 (N_43668,N_40887,N_40518);
nor U43669 (N_43669,N_40777,N_41567);
nor U43670 (N_43670,N_41723,N_41014);
nor U43671 (N_43671,N_41349,N_40369);
nand U43672 (N_43672,N_40695,N_41026);
or U43673 (N_43673,N_40555,N_41672);
xor U43674 (N_43674,N_41044,N_41971);
nor U43675 (N_43675,N_41355,N_40817);
xor U43676 (N_43676,N_40340,N_41794);
and U43677 (N_43677,N_40486,N_40090);
xor U43678 (N_43678,N_41154,N_40868);
and U43679 (N_43679,N_41876,N_41835);
nor U43680 (N_43680,N_40689,N_41415);
nand U43681 (N_43681,N_40187,N_41799);
nand U43682 (N_43682,N_41016,N_41968);
and U43683 (N_43683,N_40877,N_41089);
or U43684 (N_43684,N_40725,N_40932);
and U43685 (N_43685,N_40454,N_41804);
and U43686 (N_43686,N_40377,N_41649);
nor U43687 (N_43687,N_41865,N_40513);
nor U43688 (N_43688,N_40703,N_41048);
xnor U43689 (N_43689,N_40835,N_40237);
or U43690 (N_43690,N_41431,N_40999);
nand U43691 (N_43691,N_40446,N_40556);
nand U43692 (N_43692,N_41980,N_41754);
nand U43693 (N_43693,N_41249,N_41660);
or U43694 (N_43694,N_40841,N_40004);
and U43695 (N_43695,N_41410,N_41920);
or U43696 (N_43696,N_41571,N_41333);
nor U43697 (N_43697,N_41066,N_41960);
nor U43698 (N_43698,N_40417,N_41928);
or U43699 (N_43699,N_41712,N_40747);
nor U43700 (N_43700,N_41579,N_41429);
nor U43701 (N_43701,N_41043,N_41017);
nor U43702 (N_43702,N_41704,N_40990);
or U43703 (N_43703,N_41847,N_40658);
or U43704 (N_43704,N_41457,N_40885);
and U43705 (N_43705,N_41304,N_40073);
and U43706 (N_43706,N_41040,N_40726);
or U43707 (N_43707,N_40276,N_41888);
nor U43708 (N_43708,N_40633,N_41932);
xor U43709 (N_43709,N_40578,N_40629);
and U43710 (N_43710,N_41944,N_40018);
or U43711 (N_43711,N_40082,N_41237);
or U43712 (N_43712,N_40571,N_41861);
or U43713 (N_43713,N_41048,N_40708);
nor U43714 (N_43714,N_41147,N_41871);
or U43715 (N_43715,N_41195,N_40236);
nor U43716 (N_43716,N_40931,N_41152);
nand U43717 (N_43717,N_41254,N_41482);
xnor U43718 (N_43718,N_41732,N_40239);
xor U43719 (N_43719,N_41481,N_40098);
nand U43720 (N_43720,N_40216,N_40917);
or U43721 (N_43721,N_40597,N_40068);
or U43722 (N_43722,N_40223,N_40244);
xor U43723 (N_43723,N_41031,N_41419);
xor U43724 (N_43724,N_41803,N_40185);
and U43725 (N_43725,N_41353,N_40162);
and U43726 (N_43726,N_40681,N_41839);
or U43727 (N_43727,N_41551,N_41629);
or U43728 (N_43728,N_40852,N_41810);
nor U43729 (N_43729,N_41698,N_40569);
xor U43730 (N_43730,N_41030,N_40603);
and U43731 (N_43731,N_41491,N_41740);
nand U43732 (N_43732,N_41219,N_41114);
and U43733 (N_43733,N_41489,N_41816);
and U43734 (N_43734,N_40238,N_41125);
or U43735 (N_43735,N_40581,N_40388);
nor U43736 (N_43736,N_41546,N_40954);
xnor U43737 (N_43737,N_40583,N_40135);
and U43738 (N_43738,N_41832,N_40564);
xor U43739 (N_43739,N_41591,N_41102);
nor U43740 (N_43740,N_40111,N_40299);
and U43741 (N_43741,N_41101,N_40684);
or U43742 (N_43742,N_40862,N_40551);
xnor U43743 (N_43743,N_41480,N_41545);
nand U43744 (N_43744,N_41475,N_40815);
nor U43745 (N_43745,N_40648,N_41235);
xor U43746 (N_43746,N_40314,N_41479);
xnor U43747 (N_43747,N_40754,N_40839);
or U43748 (N_43748,N_41112,N_40302);
and U43749 (N_43749,N_41218,N_40664);
or U43750 (N_43750,N_40060,N_41530);
nor U43751 (N_43751,N_41071,N_41415);
xnor U43752 (N_43752,N_40437,N_41722);
nor U43753 (N_43753,N_41681,N_41516);
xnor U43754 (N_43754,N_40153,N_41917);
xor U43755 (N_43755,N_40136,N_40243);
and U43756 (N_43756,N_41019,N_40123);
xnor U43757 (N_43757,N_41285,N_40633);
and U43758 (N_43758,N_41453,N_41110);
nor U43759 (N_43759,N_41620,N_41307);
xnor U43760 (N_43760,N_41383,N_40389);
or U43761 (N_43761,N_41366,N_41569);
and U43762 (N_43762,N_40510,N_40584);
and U43763 (N_43763,N_41243,N_41659);
or U43764 (N_43764,N_41107,N_40546);
and U43765 (N_43765,N_40993,N_41768);
and U43766 (N_43766,N_40163,N_41236);
xor U43767 (N_43767,N_40930,N_40617);
xnor U43768 (N_43768,N_40290,N_40281);
xnor U43769 (N_43769,N_40839,N_40406);
or U43770 (N_43770,N_41420,N_41272);
xor U43771 (N_43771,N_41409,N_41934);
or U43772 (N_43772,N_41946,N_41867);
nand U43773 (N_43773,N_40758,N_41993);
nand U43774 (N_43774,N_40695,N_41122);
and U43775 (N_43775,N_41802,N_40455);
or U43776 (N_43776,N_40858,N_41054);
xor U43777 (N_43777,N_40981,N_41053);
or U43778 (N_43778,N_40278,N_40997);
and U43779 (N_43779,N_40043,N_40463);
nor U43780 (N_43780,N_40331,N_40545);
nand U43781 (N_43781,N_40727,N_40383);
nand U43782 (N_43782,N_41642,N_41573);
xnor U43783 (N_43783,N_40212,N_40912);
xnor U43784 (N_43784,N_40620,N_41803);
and U43785 (N_43785,N_41656,N_41263);
nand U43786 (N_43786,N_40197,N_40729);
nand U43787 (N_43787,N_41124,N_41538);
and U43788 (N_43788,N_40444,N_40002);
nand U43789 (N_43789,N_40804,N_41822);
or U43790 (N_43790,N_41992,N_40943);
nand U43791 (N_43791,N_40814,N_40366);
xor U43792 (N_43792,N_41095,N_41635);
or U43793 (N_43793,N_40995,N_40902);
nor U43794 (N_43794,N_41332,N_40153);
nand U43795 (N_43795,N_41197,N_41259);
nand U43796 (N_43796,N_40987,N_40070);
and U43797 (N_43797,N_41833,N_40916);
or U43798 (N_43798,N_41698,N_41036);
and U43799 (N_43799,N_40351,N_40128);
and U43800 (N_43800,N_40582,N_40790);
nand U43801 (N_43801,N_40952,N_40170);
nand U43802 (N_43802,N_40674,N_41788);
xor U43803 (N_43803,N_40650,N_41599);
nand U43804 (N_43804,N_41746,N_41876);
and U43805 (N_43805,N_40128,N_40191);
nor U43806 (N_43806,N_41866,N_41555);
or U43807 (N_43807,N_41292,N_41991);
nor U43808 (N_43808,N_41237,N_41973);
nor U43809 (N_43809,N_40381,N_40031);
nand U43810 (N_43810,N_41283,N_40112);
xnor U43811 (N_43811,N_40162,N_41872);
nand U43812 (N_43812,N_41885,N_40881);
or U43813 (N_43813,N_40530,N_41790);
and U43814 (N_43814,N_41752,N_40826);
and U43815 (N_43815,N_40298,N_41999);
nor U43816 (N_43816,N_40165,N_41646);
nand U43817 (N_43817,N_41018,N_41935);
nand U43818 (N_43818,N_40067,N_41442);
or U43819 (N_43819,N_41543,N_41168);
xor U43820 (N_43820,N_41426,N_40647);
nor U43821 (N_43821,N_40769,N_40298);
xnor U43822 (N_43822,N_41499,N_40109);
or U43823 (N_43823,N_41703,N_40939);
nand U43824 (N_43824,N_41245,N_40106);
nand U43825 (N_43825,N_40682,N_41905);
xnor U43826 (N_43826,N_40306,N_40696);
nor U43827 (N_43827,N_40245,N_40166);
xnor U43828 (N_43828,N_40356,N_40135);
nand U43829 (N_43829,N_41930,N_40348);
xor U43830 (N_43830,N_40105,N_41487);
or U43831 (N_43831,N_40786,N_40531);
nand U43832 (N_43832,N_40141,N_40618);
nor U43833 (N_43833,N_40271,N_41736);
or U43834 (N_43834,N_41004,N_41405);
xor U43835 (N_43835,N_41166,N_41862);
nand U43836 (N_43836,N_40119,N_41421);
and U43837 (N_43837,N_40820,N_40107);
xnor U43838 (N_43838,N_40415,N_40043);
nor U43839 (N_43839,N_40940,N_40319);
and U43840 (N_43840,N_40983,N_40272);
xnor U43841 (N_43841,N_40083,N_40500);
and U43842 (N_43842,N_41044,N_41806);
or U43843 (N_43843,N_40047,N_41818);
nor U43844 (N_43844,N_41507,N_40186);
or U43845 (N_43845,N_40780,N_41485);
or U43846 (N_43846,N_40491,N_40151);
or U43847 (N_43847,N_40265,N_41846);
or U43848 (N_43848,N_41356,N_40409);
and U43849 (N_43849,N_40490,N_41659);
xor U43850 (N_43850,N_40535,N_41550);
nand U43851 (N_43851,N_41165,N_41761);
or U43852 (N_43852,N_41095,N_40767);
and U43853 (N_43853,N_41239,N_40643);
nor U43854 (N_43854,N_41062,N_41824);
nand U43855 (N_43855,N_40027,N_41016);
nor U43856 (N_43856,N_40906,N_41165);
nor U43857 (N_43857,N_40864,N_40081);
and U43858 (N_43858,N_41711,N_41586);
nand U43859 (N_43859,N_41104,N_41633);
or U43860 (N_43860,N_40335,N_40172);
or U43861 (N_43861,N_40632,N_41315);
or U43862 (N_43862,N_41447,N_40055);
or U43863 (N_43863,N_40659,N_40663);
xor U43864 (N_43864,N_40412,N_40209);
and U43865 (N_43865,N_41441,N_41705);
nor U43866 (N_43866,N_40319,N_41810);
nand U43867 (N_43867,N_40281,N_41281);
nand U43868 (N_43868,N_40960,N_41095);
and U43869 (N_43869,N_41044,N_41079);
nor U43870 (N_43870,N_40085,N_41746);
xnor U43871 (N_43871,N_41521,N_40778);
nand U43872 (N_43872,N_41796,N_41817);
and U43873 (N_43873,N_41072,N_41400);
nor U43874 (N_43874,N_41168,N_40241);
xor U43875 (N_43875,N_41301,N_40502);
nand U43876 (N_43876,N_40727,N_40533);
nor U43877 (N_43877,N_40206,N_41058);
and U43878 (N_43878,N_41322,N_41116);
xnor U43879 (N_43879,N_41055,N_41559);
and U43880 (N_43880,N_40232,N_41347);
xor U43881 (N_43881,N_40617,N_40730);
or U43882 (N_43882,N_41212,N_40062);
nand U43883 (N_43883,N_40509,N_41633);
nor U43884 (N_43884,N_41026,N_40740);
nand U43885 (N_43885,N_40727,N_40877);
or U43886 (N_43886,N_41235,N_41911);
nor U43887 (N_43887,N_41500,N_41626);
and U43888 (N_43888,N_41209,N_41153);
and U43889 (N_43889,N_41507,N_40448);
and U43890 (N_43890,N_41454,N_41374);
nor U43891 (N_43891,N_40667,N_40240);
nor U43892 (N_43892,N_41792,N_41752);
and U43893 (N_43893,N_41421,N_40416);
nand U43894 (N_43894,N_40055,N_41877);
xor U43895 (N_43895,N_40226,N_41435);
nand U43896 (N_43896,N_40453,N_41621);
xor U43897 (N_43897,N_40056,N_41133);
nand U43898 (N_43898,N_41118,N_40241);
and U43899 (N_43899,N_41922,N_40951);
nor U43900 (N_43900,N_40325,N_41048);
nor U43901 (N_43901,N_41843,N_40723);
xor U43902 (N_43902,N_41770,N_41981);
or U43903 (N_43903,N_40046,N_41746);
xor U43904 (N_43904,N_40171,N_41243);
xnor U43905 (N_43905,N_40656,N_41262);
xnor U43906 (N_43906,N_40745,N_41936);
xnor U43907 (N_43907,N_40362,N_40806);
and U43908 (N_43908,N_41357,N_41260);
or U43909 (N_43909,N_40172,N_41967);
and U43910 (N_43910,N_41215,N_41920);
xnor U43911 (N_43911,N_41445,N_40426);
nor U43912 (N_43912,N_40407,N_41261);
nor U43913 (N_43913,N_40681,N_40354);
xor U43914 (N_43914,N_41973,N_40869);
and U43915 (N_43915,N_41956,N_41766);
or U43916 (N_43916,N_41251,N_41990);
nand U43917 (N_43917,N_40371,N_40169);
and U43918 (N_43918,N_40521,N_41470);
nand U43919 (N_43919,N_41921,N_40470);
nor U43920 (N_43920,N_41539,N_41548);
nor U43921 (N_43921,N_41004,N_40014);
nand U43922 (N_43922,N_41204,N_40718);
or U43923 (N_43923,N_41965,N_40962);
nor U43924 (N_43924,N_41509,N_41949);
nand U43925 (N_43925,N_40573,N_40734);
nand U43926 (N_43926,N_40643,N_40011);
nor U43927 (N_43927,N_40573,N_41488);
or U43928 (N_43928,N_40923,N_40187);
nor U43929 (N_43929,N_40730,N_40178);
nor U43930 (N_43930,N_41028,N_40669);
nand U43931 (N_43931,N_41659,N_41551);
nor U43932 (N_43932,N_41035,N_41547);
nor U43933 (N_43933,N_40007,N_40140);
or U43934 (N_43934,N_40991,N_40653);
nand U43935 (N_43935,N_40854,N_41519);
nand U43936 (N_43936,N_40015,N_41650);
and U43937 (N_43937,N_41018,N_40595);
nand U43938 (N_43938,N_41819,N_40271);
or U43939 (N_43939,N_40940,N_41693);
or U43940 (N_43940,N_41398,N_41528);
nor U43941 (N_43941,N_41836,N_40318);
or U43942 (N_43942,N_41138,N_40312);
xor U43943 (N_43943,N_40288,N_40492);
or U43944 (N_43944,N_41141,N_41041);
nand U43945 (N_43945,N_41862,N_40279);
nand U43946 (N_43946,N_41533,N_40315);
nand U43947 (N_43947,N_40747,N_40262);
xor U43948 (N_43948,N_40144,N_41857);
or U43949 (N_43949,N_40382,N_41855);
xor U43950 (N_43950,N_40547,N_40211);
or U43951 (N_43951,N_40257,N_41119);
nand U43952 (N_43952,N_41742,N_41802);
or U43953 (N_43953,N_40839,N_40813);
nand U43954 (N_43954,N_40452,N_41102);
or U43955 (N_43955,N_40071,N_41885);
nor U43956 (N_43956,N_40607,N_40464);
nor U43957 (N_43957,N_41436,N_40555);
nor U43958 (N_43958,N_40047,N_40506);
xnor U43959 (N_43959,N_40098,N_41982);
or U43960 (N_43960,N_40121,N_41203);
or U43961 (N_43961,N_40963,N_41268);
nor U43962 (N_43962,N_41578,N_40260);
xnor U43963 (N_43963,N_41968,N_40009);
xnor U43964 (N_43964,N_41194,N_41661);
nand U43965 (N_43965,N_40397,N_40003);
or U43966 (N_43966,N_41249,N_40710);
nor U43967 (N_43967,N_40484,N_40249);
or U43968 (N_43968,N_41500,N_40515);
xor U43969 (N_43969,N_40824,N_41570);
nand U43970 (N_43970,N_40355,N_41103);
and U43971 (N_43971,N_41638,N_41240);
xnor U43972 (N_43972,N_40349,N_40819);
nand U43973 (N_43973,N_40579,N_41330);
xnor U43974 (N_43974,N_41622,N_40799);
nor U43975 (N_43975,N_41573,N_40120);
and U43976 (N_43976,N_41219,N_41242);
xor U43977 (N_43977,N_40412,N_41691);
xor U43978 (N_43978,N_40500,N_40391);
or U43979 (N_43979,N_41689,N_40976);
or U43980 (N_43980,N_40435,N_40636);
and U43981 (N_43981,N_41076,N_41642);
nor U43982 (N_43982,N_41425,N_40025);
or U43983 (N_43983,N_40550,N_41590);
nand U43984 (N_43984,N_41033,N_41615);
or U43985 (N_43985,N_40091,N_40412);
xor U43986 (N_43986,N_40725,N_41864);
and U43987 (N_43987,N_40064,N_41627);
or U43988 (N_43988,N_41166,N_41810);
nand U43989 (N_43989,N_40901,N_41003);
nor U43990 (N_43990,N_41633,N_40723);
and U43991 (N_43991,N_40539,N_41369);
or U43992 (N_43992,N_41400,N_41046);
nand U43993 (N_43993,N_41605,N_40431);
nor U43994 (N_43994,N_41526,N_41759);
and U43995 (N_43995,N_41306,N_40491);
xnor U43996 (N_43996,N_41003,N_41432);
nand U43997 (N_43997,N_41604,N_40674);
and U43998 (N_43998,N_41197,N_40670);
and U43999 (N_43999,N_40711,N_41858);
xnor U44000 (N_44000,N_43063,N_42335);
and U44001 (N_44001,N_43347,N_42490);
and U44002 (N_44002,N_43760,N_42113);
and U44003 (N_44003,N_43505,N_43822);
or U44004 (N_44004,N_42909,N_42189);
xor U44005 (N_44005,N_43386,N_43232);
or U44006 (N_44006,N_42617,N_43754);
xnor U44007 (N_44007,N_42213,N_43591);
xor U44008 (N_44008,N_43617,N_43324);
or U44009 (N_44009,N_42595,N_42583);
nor U44010 (N_44010,N_43940,N_42683);
and U44011 (N_44011,N_43047,N_42770);
nand U44012 (N_44012,N_42358,N_42936);
and U44013 (N_44013,N_43529,N_42160);
xnor U44014 (N_44014,N_42257,N_43878);
or U44015 (N_44015,N_42647,N_42179);
xnor U44016 (N_44016,N_43424,N_43629);
or U44017 (N_44017,N_42688,N_42435);
nor U44018 (N_44018,N_42570,N_42137);
nand U44019 (N_44019,N_43301,N_43259);
or U44020 (N_44020,N_42550,N_43042);
and U44021 (N_44021,N_43903,N_43191);
xor U44022 (N_44022,N_43968,N_42785);
and U44023 (N_44023,N_43094,N_43739);
nor U44024 (N_44024,N_43525,N_42916);
and U44025 (N_44025,N_42798,N_43491);
or U44026 (N_44026,N_43279,N_42328);
or U44027 (N_44027,N_42873,N_42065);
nor U44028 (N_44028,N_43138,N_43181);
xor U44029 (N_44029,N_42912,N_43574);
or U44030 (N_44030,N_42453,N_43183);
and U44031 (N_44031,N_42981,N_43784);
and U44032 (N_44032,N_43111,N_43829);
or U44033 (N_44033,N_42043,N_42634);
or U44034 (N_44034,N_43560,N_43960);
xor U44035 (N_44035,N_43241,N_43297);
and U44036 (N_44036,N_42158,N_43925);
nor U44037 (N_44037,N_42661,N_43680);
nand U44038 (N_44038,N_42007,N_43412);
nand U44039 (N_44039,N_42140,N_42467);
or U44040 (N_44040,N_43351,N_42170);
nand U44041 (N_44041,N_43665,N_42760);
nor U44042 (N_44042,N_43821,N_42466);
and U44043 (N_44043,N_42939,N_42388);
or U44044 (N_44044,N_42008,N_42559);
nor U44045 (N_44045,N_42613,N_42588);
nand U44046 (N_44046,N_43485,N_42988);
and U44047 (N_44047,N_42247,N_43467);
xnor U44048 (N_44048,N_43220,N_42290);
or U44049 (N_44049,N_42071,N_42494);
xnor U44050 (N_44050,N_43995,N_43189);
nor U44051 (N_44051,N_43300,N_42356);
nand U44052 (N_44052,N_42864,N_43742);
xnor U44053 (N_44053,N_42394,N_43603);
or U44054 (N_44054,N_42793,N_43270);
xor U44055 (N_44055,N_43834,N_43783);
xor U44056 (N_44056,N_42042,N_42064);
nor U44057 (N_44057,N_42221,N_42716);
nor U44058 (N_44058,N_42668,N_43846);
nand U44059 (N_44059,N_43098,N_42723);
nor U44060 (N_44060,N_43576,N_43964);
and U44061 (N_44061,N_43712,N_42692);
nand U44062 (N_44062,N_43379,N_43371);
nand U44063 (N_44063,N_42802,N_42927);
nor U44064 (N_44064,N_42609,N_42139);
xnor U44065 (N_44065,N_42000,N_43420);
nor U44066 (N_44066,N_42407,N_43332);
nor U44067 (N_44067,N_43985,N_42225);
nor U44068 (N_44068,N_43905,N_42294);
or U44069 (N_44069,N_42729,N_43253);
xnor U44070 (N_44070,N_42994,N_43668);
nor U44071 (N_44071,N_42787,N_42266);
and U44072 (N_44072,N_43280,N_43557);
and U44073 (N_44073,N_43669,N_42258);
nor U44074 (N_44074,N_43409,N_42307);
nand U44075 (N_44075,N_43996,N_42788);
nand U44076 (N_44076,N_42431,N_42100);
or U44077 (N_44077,N_42244,N_42302);
nand U44078 (N_44078,N_42357,N_43274);
and U44079 (N_44079,N_43951,N_43394);
and U44080 (N_44080,N_43173,N_42301);
nor U44081 (N_44081,N_43879,N_42995);
xnor U44082 (N_44082,N_43919,N_42519);
and U44083 (N_44083,N_43166,N_42974);
nor U44084 (N_44084,N_43040,N_43992);
nor U44085 (N_44085,N_43918,N_42932);
xnor U44086 (N_44086,N_42708,N_43334);
nand U44087 (N_44087,N_43585,N_43015);
or U44088 (N_44088,N_43848,N_42085);
nor U44089 (N_44089,N_42272,N_42555);
or U44090 (N_44090,N_43343,N_43462);
or U44091 (N_44091,N_43683,N_42251);
xnor U44092 (N_44092,N_43400,N_42281);
nor U44093 (N_44093,N_43598,N_43445);
nand U44094 (N_44094,N_42843,N_43008);
xor U44095 (N_44095,N_42949,N_42567);
xnor U44096 (N_44096,N_42432,N_43152);
nor U44097 (N_44097,N_42915,N_43179);
nor U44098 (N_44098,N_42649,N_42155);
nor U44099 (N_44099,N_42102,N_42740);
nand U44100 (N_44100,N_43647,N_42738);
and U44101 (N_44101,N_43229,N_43818);
or U44102 (N_44102,N_43894,N_42090);
nor U44103 (N_44103,N_43490,N_42709);
xnor U44104 (N_44104,N_43054,N_43134);
and U44105 (N_44105,N_43933,N_42376);
and U44106 (N_44106,N_42292,N_43973);
nor U44107 (N_44107,N_43091,N_43026);
and U44108 (N_44108,N_42077,N_43767);
or U44109 (N_44109,N_43844,N_43611);
nor U44110 (N_44110,N_43965,N_42954);
or U44111 (N_44111,N_43478,N_42083);
or U44112 (N_44112,N_43066,N_42947);
nor U44113 (N_44113,N_43573,N_42908);
and U44114 (N_44114,N_42461,N_42628);
nand U44115 (N_44115,N_42030,N_42766);
xor U44116 (N_44116,N_42642,N_43750);
xnor U44117 (N_44117,N_43261,N_42854);
xnor U44118 (N_44118,N_43877,N_42196);
nand U44119 (N_44119,N_42901,N_42999);
nor U44120 (N_44120,N_43667,N_42874);
or U44121 (N_44121,N_43791,N_43129);
nor U44122 (N_44122,N_43582,N_42353);
and U44123 (N_44123,N_42586,N_42492);
or U44124 (N_44124,N_43081,N_42713);
nand U44125 (N_44125,N_43793,N_42336);
nand U44126 (N_44126,N_42054,N_43616);
or U44127 (N_44127,N_42327,N_42419);
and U44128 (N_44128,N_43044,N_42914);
or U44129 (N_44129,N_42626,N_42049);
nand U44130 (N_44130,N_42003,N_43049);
nor U44131 (N_44131,N_42868,N_43644);
or U44132 (N_44132,N_42533,N_43219);
or U44133 (N_44133,N_42010,N_42438);
xor U44134 (N_44134,N_43163,N_42429);
xor U44135 (N_44135,N_43169,N_43530);
xor U44136 (N_44136,N_42293,N_43789);
nand U44137 (N_44137,N_42451,N_42141);
nand U44138 (N_44138,N_42767,N_43645);
or U44139 (N_44139,N_43920,N_43836);
xnor U44140 (N_44140,N_43359,N_42022);
nand U44141 (N_44141,N_43774,N_43869);
xnor U44142 (N_44142,N_43177,N_42020);
and U44143 (N_44143,N_42488,N_43917);
nand U44144 (N_44144,N_43795,N_43514);
nor U44145 (N_44145,N_43811,N_42544);
or U44146 (N_44146,N_43225,N_43859);
nand U44147 (N_44147,N_42062,N_42489);
and U44148 (N_44148,N_43234,N_42958);
nor U44149 (N_44149,N_42314,N_43841);
nor U44150 (N_44150,N_42430,N_42774);
xor U44151 (N_44151,N_42200,N_43757);
nand U44152 (N_44152,N_43715,N_43271);
xnor U44153 (N_44153,N_42512,N_43392);
or U44154 (N_44154,N_43747,N_42153);
xnor U44155 (N_44155,N_43753,N_42863);
nand U44156 (N_44156,N_42930,N_42816);
or U44157 (N_44157,N_42922,N_43308);
nor U44158 (N_44158,N_43387,N_42361);
nand U44159 (N_44159,N_42066,N_43151);
xnor U44160 (N_44160,N_42470,N_42571);
or U44161 (N_44161,N_43638,N_43200);
nor U44162 (N_44162,N_43425,N_42385);
or U44163 (N_44163,N_43547,N_43099);
or U44164 (N_44164,N_43938,N_43655);
nor U44165 (N_44165,N_42581,N_43405);
nor U44166 (N_44166,N_42562,N_42056);
nor U44167 (N_44167,N_43036,N_42233);
and U44168 (N_44168,N_42693,N_42454);
nand U44169 (N_44169,N_42354,N_43499);
xnor U44170 (N_44170,N_42822,N_43536);
and U44171 (N_44171,N_42082,N_43595);
or U44172 (N_44172,N_42261,N_42029);
xnor U44173 (N_44173,N_42190,N_43814);
xnor U44174 (N_44174,N_43150,N_43549);
xnor U44175 (N_44175,N_43796,N_43454);
and U44176 (N_44176,N_42607,N_43475);
or U44177 (N_44177,N_42526,N_42323);
nand U44178 (N_44178,N_43546,N_43051);
and U44179 (N_44179,N_43362,N_43931);
and U44180 (N_44180,N_43993,N_43289);
xnor U44181 (N_44181,N_42289,N_42117);
and U44182 (N_44182,N_43205,N_42277);
nand U44183 (N_44183,N_43787,N_42724);
nor U44184 (N_44184,N_42406,N_43780);
xor U44185 (N_44185,N_42841,N_42624);
nand U44186 (N_44186,N_43306,N_43866);
or U44187 (N_44187,N_43902,N_43493);
or U44188 (N_44188,N_43315,N_42993);
and U44189 (N_44189,N_43843,N_42161);
or U44190 (N_44190,N_42875,N_42836);
nand U44191 (N_44191,N_42097,N_43874);
or U44192 (N_44192,N_42989,N_42659);
nand U44193 (N_44193,N_42831,N_43430);
or U44194 (N_44194,N_43587,N_43688);
or U44195 (N_44195,N_42918,N_43093);
nor U44196 (N_44196,N_42871,N_42757);
and U44197 (N_44197,N_43446,N_43907);
nor U44198 (N_44198,N_42449,N_43358);
or U44199 (N_44199,N_43268,N_43620);
xnor U44200 (N_44200,N_42346,N_42001);
or U44201 (N_44201,N_42011,N_43311);
nor U44202 (N_44202,N_42185,N_43293);
nor U44203 (N_44203,N_43687,N_42395);
xor U44204 (N_44204,N_42515,N_43520);
and U44205 (N_44205,N_42920,N_43666);
nand U44206 (N_44206,N_42675,N_43136);
and U44207 (N_44207,N_42574,N_43501);
xnor U44208 (N_44208,N_42402,N_42373);
and U44209 (N_44209,N_42173,N_43000);
nand U44210 (N_44210,N_43033,N_42664);
xnor U44211 (N_44211,N_42762,N_42149);
xor U44212 (N_44212,N_42685,N_42603);
nor U44213 (N_44213,N_42534,N_42735);
and U44214 (N_44214,N_42471,N_43427);
nor U44215 (N_44215,N_42672,N_43007);
nor U44216 (N_44216,N_42138,N_43982);
nor U44217 (N_44217,N_42789,N_42241);
or U44218 (N_44218,N_42697,N_43231);
or U44219 (N_44219,N_42681,N_43159);
xnor U44220 (N_44220,N_43075,N_43762);
nand U44221 (N_44221,N_43414,N_42345);
nand U44222 (N_44222,N_42630,N_43707);
nand U44223 (N_44223,N_43722,N_42950);
xor U44224 (N_44224,N_42881,N_42265);
or U44225 (N_44225,N_42483,N_43615);
nand U44226 (N_44226,N_43786,N_43608);
or U44227 (N_44227,N_42464,N_43227);
nor U44228 (N_44228,N_42622,N_43823);
and U44229 (N_44229,N_42084,N_42690);
nand U44230 (N_44230,N_42542,N_42876);
nand U44231 (N_44231,N_42764,N_43524);
nand U44232 (N_44232,N_43221,N_42771);
and U44233 (N_44233,N_42734,N_42312);
nor U44234 (N_44234,N_43552,N_42144);
nor U44235 (N_44235,N_43817,N_42703);
xnor U44236 (N_44236,N_42387,N_42931);
or U44237 (N_44237,N_43987,N_43165);
nor U44238 (N_44238,N_42486,N_43978);
nor U44239 (N_44239,N_43888,N_42645);
nand U44240 (N_44240,N_43005,N_43941);
nand U44241 (N_44241,N_43277,N_42543);
xor U44242 (N_44242,N_43592,N_43802);
xnor U44243 (N_44243,N_43676,N_42990);
nor U44244 (N_44244,N_42132,N_42790);
or U44245 (N_44245,N_43816,N_42652);
nor U44246 (N_44246,N_42456,N_42380);
nor U44247 (N_44247,N_43117,N_43368);
nor U44248 (N_44248,N_43391,N_42725);
nor U44249 (N_44249,N_43443,N_43050);
xnor U44250 (N_44250,N_42428,N_42627);
nor U44251 (N_44251,N_42107,N_42520);
or U44252 (N_44252,N_42638,N_43135);
nand U44253 (N_44253,N_42168,N_42363);
and U44254 (N_44254,N_43466,N_43519);
xor U44255 (N_44255,N_42338,N_43022);
nor U44256 (N_44256,N_43635,N_43590);
nor U44257 (N_44257,N_42946,N_42375);
and U44258 (N_44258,N_42135,N_43407);
and U44259 (N_44259,N_42699,N_42210);
xor U44260 (N_44260,N_42513,N_42215);
nand U44261 (N_44261,N_43428,N_42459);
nand U44262 (N_44262,N_42014,N_43704);
xor U44263 (N_44263,N_43484,N_43577);
xor U44264 (N_44264,N_43981,N_43373);
xnor U44265 (N_44265,N_43532,N_43447);
xor U44266 (N_44266,N_42303,N_43527);
nand U44267 (N_44267,N_42598,N_42339);
and U44268 (N_44268,N_43618,N_43521);
and U44269 (N_44269,N_43523,N_42287);
and U44270 (N_44270,N_43876,N_42805);
nand U44271 (N_44271,N_42463,N_42905);
nand U44272 (N_44272,N_43959,N_42465);
nand U44273 (N_44273,N_42860,N_43141);
xor U44274 (N_44274,N_42561,N_43310);
and U44275 (N_44275,N_42839,N_43526);
nand U44276 (N_44276,N_43323,N_42678);
xor U44277 (N_44277,N_43926,N_43283);
xnor U44278 (N_44278,N_43423,N_42126);
and U44279 (N_44279,N_43991,N_42565);
or U44280 (N_44280,N_42316,N_42156);
and U44281 (N_44281,N_42481,N_42031);
xor U44282 (N_44282,N_43276,N_43284);
nand U44283 (N_44283,N_42013,N_43132);
nand U44284 (N_44284,N_43282,N_43867);
and U44285 (N_44285,N_43360,N_42367);
xor U44286 (N_44286,N_42986,N_43448);
nor U44287 (N_44287,N_42162,N_42879);
or U44288 (N_44288,N_43773,N_43353);
or U44289 (N_44289,N_43746,N_43732);
or U44290 (N_44290,N_43201,N_43735);
and U44291 (N_44291,N_42423,N_42830);
nand U44292 (N_44292,N_42101,N_42671);
and U44293 (N_44293,N_42195,N_42743);
nor U44294 (N_44294,N_43439,N_42252);
nand U44295 (N_44295,N_43537,N_43316);
and U44296 (N_44296,N_42779,N_43455);
or U44297 (N_44297,N_43893,N_43014);
xor U44298 (N_44298,N_42103,N_42827);
xnor U44299 (N_44299,N_42374,N_42178);
and U44300 (N_44300,N_43193,N_42892);
and U44301 (N_44301,N_42411,N_42476);
or U44302 (N_44302,N_43733,N_43575);
and U44303 (N_44303,N_43952,N_42517);
or U44304 (N_44304,N_42991,N_43634);
and U44305 (N_44305,N_42953,N_42450);
nand U44306 (N_44306,N_43511,N_43325);
xor U44307 (N_44307,N_43660,N_43375);
and U44308 (N_44308,N_42291,N_43679);
xnor U44309 (N_44309,N_42035,N_43236);
and U44310 (N_44310,N_42823,N_42590);
or U44311 (N_44311,N_42006,N_43623);
and U44312 (N_44312,N_43745,N_42019);
xor U44313 (N_44313,N_43436,N_42305);
nand U44314 (N_44314,N_42768,N_43857);
and U44315 (N_44315,N_42255,N_43035);
xnor U44316 (N_44316,N_42756,N_42984);
nor U44317 (N_44317,N_42485,N_43174);
and U44318 (N_44318,N_43649,N_42352);
and U44319 (N_44319,N_43184,N_42612);
nor U44320 (N_44320,N_42899,N_43724);
nor U44321 (N_44321,N_43365,N_42573);
nand U44322 (N_44322,N_43759,N_43604);
and U44323 (N_44323,N_43095,N_42437);
nor U44324 (N_44324,N_42941,N_43309);
nor U44325 (N_44325,N_43614,N_42903);
nand U44326 (N_44326,N_42315,N_43214);
and U44327 (N_44327,N_43019,N_43432);
nor U44328 (N_44328,N_42318,N_42209);
nand U44329 (N_44329,N_43442,N_43492);
nor U44330 (N_44330,N_42795,N_43143);
or U44331 (N_44331,N_43705,N_42580);
xor U44332 (N_44332,N_42585,N_43648);
nand U44333 (N_44333,N_42017,N_43674);
nand U44334 (N_44334,N_42528,N_43197);
or U44335 (N_44335,N_42938,N_42749);
nor U44336 (N_44336,N_43998,N_43067);
xor U44337 (N_44337,N_43643,N_43216);
nor U44338 (N_44338,N_43589,N_43522);
nor U44339 (N_44339,N_42809,N_43226);
and U44340 (N_44340,N_42641,N_42263);
nand U44341 (N_44341,N_42973,N_42321);
nor U44342 (N_44342,N_43207,N_42553);
nor U44343 (N_44343,N_42782,N_43642);
nand U44344 (N_44344,N_43901,N_42803);
xor U44345 (N_44345,N_43772,N_42186);
nor U44346 (N_44346,N_42143,N_42217);
nand U44347 (N_44347,N_43507,N_43775);
and U44348 (N_44348,N_43555,N_42504);
nor U44349 (N_44349,N_42781,N_43078);
and U44350 (N_44350,N_43686,N_42184);
and U44351 (N_44351,N_43534,N_42442);
nand U44352 (N_44352,N_42473,N_43662);
nand U44353 (N_44353,N_43041,N_43781);
nor U44354 (N_44354,N_42880,N_42424);
xor U44355 (N_44355,N_42378,N_42028);
xor U44356 (N_44356,N_42259,N_43376);
nand U44357 (N_44357,N_43971,N_43853);
nor U44358 (N_44358,N_43550,N_43923);
and U44359 (N_44359,N_42531,N_42837);
nor U44360 (N_44360,N_43806,N_43065);
xor U44361 (N_44361,N_42667,N_43073);
and U44362 (N_44362,N_42413,N_43977);
xnor U44363 (N_44363,N_42507,N_42971);
xnor U44364 (N_44364,N_42576,N_43950);
or U44365 (N_44365,N_43140,N_42655);
nand U44366 (N_44366,N_43060,N_42208);
nor U44367 (N_44367,N_43266,N_43090);
xnor U44368 (N_44368,N_42698,N_42500);
nor U44369 (N_44369,N_43936,N_42582);
xnor U44370 (N_44370,N_43771,N_43086);
and U44371 (N_44371,N_42382,N_43883);
nor U44372 (N_44372,N_42276,N_43383);
nor U44373 (N_44373,N_43922,N_42957);
nand U44374 (N_44374,N_42288,N_42324);
or U44375 (N_44375,N_43468,N_43429);
nor U44376 (N_44376,N_42333,N_43769);
nand U44377 (N_44377,N_43855,N_43770);
xnor U44378 (N_44378,N_42439,N_42418);
and U44379 (N_44379,N_43963,N_43625);
and U44380 (N_44380,N_42797,N_43540);
or U44381 (N_44381,N_43654,N_43109);
or U44382 (N_44382,N_42639,N_42980);
nor U44383 (N_44383,N_43006,N_43994);
nor U44384 (N_44384,N_42817,N_43498);
nand U44385 (N_44385,N_42621,N_43048);
xor U44386 (N_44386,N_42845,N_42521);
and U44387 (N_44387,N_43886,N_43417);
nor U44388 (N_44388,N_43438,N_42337);
nand U44389 (N_44389,N_43533,N_43377);
or U44390 (N_44390,N_43218,N_42237);
nor U44391 (N_44391,N_42778,N_42744);
nor U44392 (N_44392,N_43228,N_42012);
and U44393 (N_44393,N_43967,N_42942);
nand U44394 (N_44394,N_43194,N_43633);
and U44395 (N_44395,N_43502,N_43082);
nor U44396 (N_44396,N_42249,N_42351);
or U44397 (N_44397,N_42036,N_43906);
xor U44398 (N_44398,N_43720,N_43570);
xnor U44399 (N_44399,N_43858,N_43449);
or U44400 (N_44400,N_43864,N_43947);
nand U44401 (N_44401,N_43327,N_42821);
nor U44402 (N_44402,N_43800,N_43128);
nand U44403 (N_44403,N_43110,N_43397);
and U44404 (N_44404,N_43291,N_42911);
or U44405 (N_44405,N_43390,N_43700);
or U44406 (N_44406,N_43808,N_42427);
and U44407 (N_44407,N_42242,N_43304);
nand U44408 (N_44408,N_42154,N_43356);
or U44409 (N_44409,N_42283,N_42086);
and U44410 (N_44410,N_42720,N_42355);
nand U44411 (N_44411,N_43743,N_43085);
nand U44412 (N_44412,N_42308,N_43809);
nor U44413 (N_44413,N_42963,N_42207);
or U44414 (N_44414,N_42886,N_43190);
xnor U44415 (N_44415,N_42384,N_42150);
xor U44416 (N_44416,N_43659,N_42243);
nor U44417 (N_44417,N_43021,N_42917);
nor U44418 (N_44418,N_42273,N_43029);
nand U44419 (N_44419,N_43398,N_42956);
xnor U44420 (N_44420,N_43278,N_43096);
or U44421 (N_44421,N_42940,N_43698);
nand U44422 (N_44422,N_42660,N_42523);
nor U44423 (N_44423,N_42152,N_43953);
xor U44424 (N_44424,N_42885,N_42393);
or U44425 (N_44425,N_42887,N_43804);
nand U44426 (N_44426,N_42067,N_42890);
xnor U44427 (N_44427,N_43758,N_43341);
nand U44428 (N_44428,N_42578,N_42371);
xor U44429 (N_44429,N_43556,N_43212);
nor U44430 (N_44430,N_43559,N_42410);
nand U44431 (N_44431,N_43170,N_43037);
nor U44432 (N_44432,N_42165,N_43144);
xnor U44433 (N_44433,N_42965,N_42616);
or U44434 (N_44434,N_42631,N_43374);
or U44435 (N_44435,N_43908,N_43119);
and U44436 (N_44436,N_42342,N_42188);
and U44437 (N_44437,N_43752,N_43097);
and U44438 (N_44438,N_43785,N_42964);
nor U44439 (N_44439,N_42902,N_42349);
xnor U44440 (N_44440,N_43406,N_42623);
and U44441 (N_44441,N_43388,N_43500);
nor U44442 (N_44442,N_43849,N_42810);
nand U44443 (N_44443,N_43223,N_42643);
and U44444 (N_44444,N_43012,N_42566);
xor U44445 (N_44445,N_43419,N_42389);
nand U44446 (N_44446,N_42426,N_43069);
or U44447 (N_44447,N_43675,N_42040);
nor U44448 (N_44448,N_42594,N_42304);
nor U44449 (N_44449,N_43980,N_42775);
nand U44450 (N_44450,N_42896,N_42441);
and U44451 (N_44451,N_42646,N_42813);
nand U44452 (N_44452,N_42219,N_43719);
nor U44453 (N_44453,N_43562,N_42945);
nand U44454 (N_44454,N_43003,N_43120);
nor U44455 (N_44455,N_43815,N_43267);
xnor U44456 (N_44456,N_43303,N_43621);
nand U44457 (N_44457,N_42112,N_43820);
and U44458 (N_44458,N_42166,N_42446);
and U44459 (N_44459,N_43255,N_42721);
or U44460 (N_44460,N_42861,N_42472);
xor U44461 (N_44461,N_43929,N_43433);
nand U44462 (N_44462,N_42808,N_42601);
nand U44463 (N_44463,N_42034,N_42877);
and U44464 (N_44464,N_43142,N_43799);
xor U44465 (N_44465,N_43435,N_43102);
or U44466 (N_44466,N_43508,N_43413);
or U44467 (N_44467,N_42919,N_42344);
nor U44468 (N_44468,N_42651,N_42811);
and U44469 (N_44469,N_43865,N_43250);
and U44470 (N_44470,N_42087,N_43717);
and U44471 (N_44471,N_42759,N_42267);
and U44472 (N_44472,N_43213,N_43870);
or U44473 (N_44473,N_43763,N_42282);
nor U44474 (N_44474,N_42812,N_43074);
and U44475 (N_44475,N_43175,N_43630);
nand U44476 (N_44476,N_42791,N_42985);
nand U44477 (N_44477,N_43613,N_43935);
nand U44478 (N_44478,N_43456,N_42761);
and U44479 (N_44479,N_42405,N_43211);
xnor U44480 (N_44480,N_43337,N_43314);
or U44481 (N_44481,N_43622,N_42203);
nor U44482 (N_44482,N_42487,N_43710);
nor U44483 (N_44483,N_42894,N_42669);
nor U44484 (N_44484,N_42474,N_43914);
xnor U44485 (N_44485,N_42694,N_43909);
and U44486 (N_44486,N_42167,N_42633);
and U44487 (N_44487,N_42460,N_43131);
nor U44488 (N_44488,N_43990,N_42701);
or U44489 (N_44489,N_43565,N_42514);
nand U44490 (N_44490,N_42091,N_42620);
or U44491 (N_44491,N_42882,N_42921);
nand U44492 (N_44492,N_42181,N_42271);
nand U44493 (N_44493,N_43064,N_42972);
nor U44494 (N_44494,N_43457,N_43404);
xor U44495 (N_44495,N_42852,N_42700);
nand U44496 (N_44496,N_43782,N_43727);
xnor U44497 (N_44497,N_42401,N_42127);
and U44498 (N_44498,N_42814,N_43708);
or U44499 (N_44499,N_42458,N_43681);
nor U44500 (N_44500,N_42391,N_43488);
nand U44501 (N_44501,N_42250,N_42635);
xor U44502 (N_44502,N_43224,N_43954);
xnor U44503 (N_44503,N_43639,N_42379);
xnor U44504 (N_44504,N_42392,N_43510);
or U44505 (N_44505,N_42975,N_43709);
or U44506 (N_44506,N_43663,N_42591);
and U44507 (N_44507,N_42510,N_43600);
nor U44508 (N_44508,N_43104,N_43807);
nand U44509 (N_44509,N_42502,N_42080);
xnor U44510 (N_44510,N_42420,N_43528);
nand U44511 (N_44511,N_42230,N_43154);
xnor U44512 (N_44512,N_42278,N_43084);
and U44513 (N_44513,N_43972,N_43024);
xnor U44514 (N_44514,N_43512,N_43930);
nor U44515 (N_44515,N_42926,N_42849);
or U44516 (N_44516,N_43338,N_42479);
or U44517 (N_44517,N_43336,N_43805);
or U44518 (N_44518,N_43330,N_42900);
or U44519 (N_44519,N_43363,N_43450);
and U44520 (N_44520,N_42201,N_43402);
nor U44521 (N_44521,N_42298,N_43581);
nor U44522 (N_44522,N_43531,N_42850);
xor U44523 (N_44523,N_42889,N_42577);
or U44524 (N_44524,N_42996,N_42403);
nor U44525 (N_44525,N_42268,N_42935);
and U44526 (N_44526,N_42895,N_42637);
and U44527 (N_44527,N_42977,N_43602);
nand U44528 (N_44528,N_43023,N_42075);
or U44529 (N_44529,N_43452,N_43538);
and U44530 (N_44530,N_42239,N_43369);
nand U44531 (N_44531,N_42151,N_43477);
nor U44532 (N_44532,N_42296,N_42755);
and U44533 (N_44533,N_43637,N_42717);
nand U44534 (N_44534,N_43695,N_43105);
xor U44535 (N_44535,N_42320,N_42199);
and U44536 (N_44536,N_43056,N_42044);
or U44537 (N_44537,N_43032,N_42695);
nor U44538 (N_44538,N_42377,N_42673);
and U44539 (N_44539,N_43852,N_43464);
xnor U44540 (N_44540,N_43344,N_43946);
xnor U44541 (N_44541,N_42119,N_42684);
nand U44542 (N_44542,N_43837,N_42269);
nand U44543 (N_44543,N_43320,N_43803);
or U44544 (N_44544,N_43607,N_42592);
or U44545 (N_44545,N_43596,N_42129);
nand U44546 (N_44546,N_42038,N_42632);
and U44547 (N_44547,N_43087,N_42840);
xor U44548 (N_44548,N_43403,N_42300);
and U44549 (N_44549,N_43955,N_42969);
nor U44550 (N_44550,N_43480,N_42477);
nand U44551 (N_44551,N_43340,N_42711);
and U44552 (N_44552,N_42792,N_43350);
and U44553 (N_44553,N_43880,N_43898);
or U44554 (N_44554,N_43010,N_43509);
xnor U44555 (N_44555,N_42493,N_42214);
nor U44556 (N_44556,N_43670,N_42176);
nand U44557 (N_44557,N_42096,N_42383);
xor U44558 (N_44558,N_42496,N_43009);
xnor U44559 (N_44559,N_43856,N_43765);
nor U44560 (N_44560,N_42884,N_43691);
xnor U44561 (N_44561,N_43958,N_42913);
xor U44562 (N_44562,N_43101,N_42747);
and U44563 (N_44563,N_43899,N_43355);
xor U44564 (N_44564,N_42865,N_43285);
and U44565 (N_44565,N_43335,N_42110);
xor U44566 (N_44566,N_42898,N_43764);
nor U44567 (N_44567,N_43415,N_42122);
and U44568 (N_44568,N_43126,N_43797);
nand U44569 (N_44569,N_43418,N_42216);
xor U44570 (N_44570,N_42937,N_43943);
and U44571 (N_44571,N_42722,N_43384);
nand U44572 (N_44572,N_42340,N_42187);
nor U44573 (N_44573,N_43263,N_42706);
nand U44574 (N_44574,N_42686,N_43871);
xnor U44575 (N_44575,N_43734,N_43543);
nand U44576 (N_44576,N_43706,N_42560);
nor U44577 (N_44577,N_42360,N_43610);
or U44578 (N_44578,N_43957,N_43755);
nand U44579 (N_44579,N_43677,N_42815);
nand U44580 (N_44580,N_43932,N_43058);
or U44581 (N_44581,N_43281,N_43192);
nor U44582 (N_44582,N_43671,N_42260);
nand U44583 (N_44583,N_43632,N_42869);
xor U44584 (N_44584,N_43437,N_42444);
xnor U44585 (N_44585,N_43875,N_43966);
nor U44586 (N_44586,N_43245,N_43792);
or U44587 (N_44587,N_43470,N_43487);
or U44588 (N_44588,N_43233,N_43046);
and U44589 (N_44589,N_43020,N_42906);
nor U44590 (N_44590,N_42677,N_42579);
nor U44591 (N_44591,N_43378,N_43106);
xnor U44592 (N_44592,N_42857,N_42741);
or U44593 (N_44593,N_42099,N_43586);
nor U44594 (N_44594,N_43328,N_42820);
nor U44595 (N_44595,N_42398,N_43850);
xnor U44596 (N_44596,N_43061,N_42226);
or U44597 (N_44597,N_42171,N_43609);
xor U44598 (N_44598,N_43260,N_42362);
and U44599 (N_44599,N_43626,N_43256);
nand U44600 (N_44600,N_43504,N_42524);
and U44601 (N_44601,N_43290,N_42491);
or U44602 (N_44602,N_43729,N_42396);
nor U44603 (N_44603,N_42564,N_42676);
nor U44604 (N_44604,N_42910,N_43070);
or U44605 (N_44605,N_42754,N_43593);
and U44606 (N_44606,N_43605,N_43657);
and U44607 (N_44607,N_42838,N_43381);
xor U44608 (N_44608,N_42615,N_42847);
nor U44609 (N_44609,N_42348,N_42499);
nor U44610 (N_44610,N_42967,N_43396);
and U44611 (N_44611,N_42452,N_43701);
nand U44612 (N_44612,N_43030,N_43286);
nor U44613 (N_44613,N_43928,N_43385);
and U44614 (N_44614,N_42800,N_42835);
nor U44615 (N_44615,N_42046,N_43518);
nand U44616 (N_44616,N_42048,N_42807);
nor U44617 (N_44617,N_43217,N_43318);
xor U44618 (N_44618,N_43884,N_42386);
or U44619 (N_44619,N_42962,N_42705);
and U44620 (N_44620,N_42842,N_43089);
nand U44621 (N_44621,N_42506,N_43039);
xnor U44622 (N_44622,N_43215,N_42397);
and U44623 (N_44623,N_43833,N_43599);
nand U44624 (N_44624,N_42848,N_42682);
nor U44625 (N_44625,N_43243,N_42205);
nand U44626 (N_44626,N_43411,N_42872);
nand U44627 (N_44627,N_42979,N_43295);
xor U44628 (N_44628,N_42177,N_43882);
or U44629 (N_44629,N_43364,N_42331);
and U44630 (N_44630,N_43945,N_43298);
nor U44631 (N_44631,N_43116,N_43842);
xor U44632 (N_44632,N_43566,N_43986);
nand U44633 (N_44633,N_43548,N_43399);
nand U44634 (N_44634,N_42944,N_43690);
nor U44635 (N_44635,N_43458,N_42240);
nor U44636 (N_44636,N_42462,N_43516);
xor U44637 (N_44637,N_43651,N_42404);
nand U44638 (N_44638,N_43597,N_43969);
and U44639 (N_44639,N_43862,N_42753);
nand U44640 (N_44640,N_42055,N_42309);
xor U44641 (N_44641,N_42796,N_42326);
nor U44642 (N_44642,N_43984,N_42859);
xor U44643 (N_44643,N_42399,N_42737);
nand U44644 (N_44644,N_42704,N_42742);
and U44645 (N_44645,N_43696,N_42604);
nand U44646 (N_44646,N_42952,N_42522);
nand U44647 (N_44647,N_42169,N_43125);
or U44648 (N_44648,N_43956,N_43471);
and U44649 (N_44649,N_43851,N_42883);
and U44650 (N_44650,N_43421,N_43744);
nor U44651 (N_44651,N_42846,N_42718);
or U44652 (N_44652,N_43172,N_42365);
nand U44653 (N_44653,N_42540,N_43723);
and U44654 (N_44654,N_42033,N_42134);
nor U44655 (N_44655,N_42878,N_43975);
and U44656 (N_44656,N_42072,N_42317);
and U44657 (N_44657,N_43265,N_43002);
and U44658 (N_44658,N_43294,N_42417);
xnor U44659 (N_44659,N_42366,N_42076);
or U44660 (N_44660,N_42416,N_42834);
and U44661 (N_44661,N_42587,N_43673);
and U44662 (N_44662,N_42095,N_42763);
xnor U44663 (N_44663,N_43601,N_43580);
xnor U44664 (N_44664,N_42425,N_43222);
nor U44665 (N_44665,N_43198,N_43028);
nor U44666 (N_44666,N_43474,N_43713);
or U44667 (N_44667,N_42804,N_42050);
nand U44668 (N_44668,N_43252,N_43017);
or U44669 (N_44669,N_42018,N_43472);
nor U44670 (N_44670,N_42211,N_42248);
and U44671 (N_44671,N_42231,N_43636);
xor U44672 (N_44672,N_42608,N_43176);
and U44673 (N_44673,N_42133,N_42262);
or U44674 (N_44674,N_42801,N_43513);
nor U44675 (N_44675,N_43962,N_43461);
and U44676 (N_44676,N_42254,N_42182);
xnor U44677 (N_44677,N_42866,N_43057);
or U44678 (N_44678,N_42313,N_42961);
or U44679 (N_44679,N_42223,N_43465);
xor U44680 (N_44680,N_42147,N_42016);
and U44681 (N_44681,N_43702,N_42640);
nor U44682 (N_44682,N_42750,N_42537);
xnor U44683 (N_44683,N_43887,N_43761);
or U44684 (N_44684,N_43756,N_42710);
nor U44685 (N_44685,N_42128,N_43890);
or U44686 (N_44686,N_43199,N_43410);
or U44687 (N_44687,N_43408,N_43678);
nand U44688 (N_44688,N_42114,N_43921);
and U44689 (N_44689,N_43441,N_42088);
xor U44690 (N_44690,N_42270,N_43168);
nand U44691 (N_44691,N_42194,N_42657);
xor U44692 (N_44692,N_42978,N_43483);
nand U44693 (N_44693,N_42589,N_42501);
or U44694 (N_44694,N_42867,N_42306);
and U44695 (N_44695,N_42712,N_43563);
nand U44696 (N_44696,N_42334,N_42746);
xor U44697 (N_44697,N_42228,N_42319);
xnor U44698 (N_44698,N_42907,N_43195);
or U44699 (N_44699,N_42976,N_43845);
xnor U44700 (N_44700,N_43551,N_43370);
or U44701 (N_44701,N_42575,N_43187);
xnor U44702 (N_44702,N_43571,N_43299);
or U44703 (N_44703,N_42172,N_43317);
or U44704 (N_44704,N_43203,N_43481);
and U44705 (N_44705,N_42436,N_43357);
nor U44706 (N_44706,N_43121,N_42893);
nand U44707 (N_44707,N_43269,N_42123);
xor U44708 (N_44708,N_43812,N_43367);
or U44709 (N_44709,N_43656,N_42731);
xnor U44710 (N_44710,N_43970,N_43497);
and U44711 (N_44711,N_42274,N_43204);
or U44712 (N_44712,N_43631,N_43319);
nand U44713 (N_44713,N_43149,N_43572);
xor U44714 (N_44714,N_42739,N_42853);
xnor U44715 (N_44715,N_43153,N_43584);
or U44716 (N_44716,N_42605,N_42212);
xor U44717 (N_44717,N_42527,N_42924);
nor U44718 (N_44718,N_43292,N_43794);
and U44719 (N_44719,N_42057,N_43788);
nand U44720 (N_44720,N_43145,N_42109);
xor U44721 (N_44721,N_43322,N_43249);
xnor U44722 (N_44722,N_43148,N_42124);
nand U44723 (N_44723,N_42058,N_42535);
and U44724 (N_44724,N_42434,N_43868);
nor U44725 (N_44725,N_42532,N_42142);
and U44726 (N_44726,N_43694,N_42037);
or U44727 (N_44727,N_43476,N_43372);
and U44728 (N_44728,N_43242,N_43459);
xor U44729 (N_44729,N_43164,N_42060);
nand U44730 (N_44730,N_42484,N_42563);
and U44731 (N_44731,N_42025,N_43779);
nand U44732 (N_44732,N_43913,N_43053);
nor U44733 (N_44733,N_43544,N_43088);
xor U44734 (N_44734,N_42833,N_43473);
or U44735 (N_44735,N_43431,N_43366);
xnor U44736 (N_44736,N_43916,N_42870);
or U44737 (N_44737,N_42381,N_42079);
nor U44738 (N_44738,N_42204,N_43881);
xor U44739 (N_44739,N_42414,N_43389);
and U44740 (N_44740,N_43251,N_43254);
xor U44741 (N_44741,N_43004,N_42163);
nand U44742 (N_44742,N_43157,N_42665);
or U44743 (N_44743,N_43703,N_43983);
nor U44744 (N_44744,N_42844,N_42600);
nand U44745 (N_44745,N_43778,N_43167);
nand U44746 (N_44746,N_43068,N_43275);
and U44747 (N_44747,N_43999,N_43737);
and U44748 (N_44748,N_42511,N_42440);
and U44749 (N_44749,N_42131,N_42730);
nand U44750 (N_44750,N_42529,N_43974);
and U44751 (N_44751,N_43264,N_42482);
or U44752 (N_44752,N_43891,N_42636);
nand U44753 (N_44753,N_42120,N_43451);
and U44754 (N_44754,N_43989,N_42777);
nand U44755 (N_44755,N_43684,N_42275);
xor U44756 (N_44756,N_43942,N_42238);
nor U44757 (N_44757,N_42246,N_43819);
nor U44758 (N_44758,N_42554,N_42541);
or U44759 (N_44759,N_42136,N_43331);
xor U44760 (N_44760,N_42125,N_42359);
or U44761 (N_44761,N_43124,N_43100);
nor U44762 (N_44762,N_42063,N_43685);
or U44763 (N_44763,N_43258,N_42116);
xnor U44764 (N_44764,N_42610,N_43349);
xor U44765 (N_44765,N_43161,N_42059);
xor U44766 (N_44766,N_42002,N_42745);
and U44767 (N_44767,N_42925,N_42332);
nor U44768 (N_44768,N_43640,N_42732);
nand U44769 (N_44769,N_43352,N_43348);
nor U44770 (N_44770,N_43517,N_42551);
xor U44771 (N_44771,N_43469,N_43801);
nand U44772 (N_44772,N_43077,N_42475);
and U44773 (N_44773,N_43826,N_42232);
nor U44774 (N_44774,N_42457,N_43641);
or U44775 (N_44775,N_43001,N_43146);
nor U44776 (N_44776,N_43139,N_43749);
and U44777 (N_44777,N_42193,N_42078);
xnor U44778 (N_44778,N_42015,N_43725);
nor U44779 (N_44779,N_42047,N_42236);
nand U44780 (N_44780,N_42498,N_42118);
and U44781 (N_44781,N_42409,N_43692);
xor U44782 (N_44782,N_43937,N_43071);
nor U44783 (N_44783,N_42648,N_42503);
or U44784 (N_44784,N_43988,N_42943);
xnor U44785 (N_44785,N_42696,N_42786);
nand U44786 (N_44786,N_43976,N_42422);
nor U44787 (N_44787,N_43579,N_42897);
or U44788 (N_44788,N_42776,N_43594);
nand U44789 (N_44789,N_42297,N_43156);
and U44790 (N_44790,N_43401,N_42180);
or U44791 (N_44791,N_42372,N_43736);
nor U44792 (N_44792,N_42279,N_42347);
nand U44793 (N_44793,N_43897,N_43247);
or U44794 (N_44794,N_42081,N_42468);
xor U44795 (N_44795,N_42068,N_43558);
xnor U44796 (N_44796,N_43896,N_43835);
nand U44797 (N_44797,N_42829,N_42235);
nor U44798 (N_44798,N_43776,N_43262);
nor U44799 (N_44799,N_43944,N_42549);
nand U44800 (N_44800,N_43354,N_43202);
nor U44801 (N_44801,N_43011,N_42558);
and U44802 (N_44802,N_43103,N_42370);
xnor U44803 (N_44803,N_42736,N_42322);
and U44804 (N_44804,N_43380,N_43716);
or U44805 (N_44805,N_42552,N_43578);
nor U44806 (N_44806,N_42691,N_43130);
nor U44807 (N_44807,N_43904,N_43257);
or U44808 (N_44808,N_42733,N_42784);
nor U44809 (N_44809,N_43731,N_43672);
and U44810 (N_44810,N_42093,N_43721);
nor U44811 (N_44811,N_42662,N_43016);
nor U44812 (N_44812,N_43209,N_42175);
xor U44813 (N_44813,N_43313,N_42928);
or U44814 (N_44814,N_42041,N_42518);
and U44815 (N_44815,N_42773,N_43515);
nor U44816 (N_44816,N_42658,N_43463);
and U44817 (N_44817,N_43112,N_43180);
nand U44818 (N_44818,N_42614,N_43568);
nor U44819 (N_44819,N_42987,N_42227);
xnor U44820 (N_44820,N_42783,N_43158);
or U44821 (N_44821,N_43237,N_42412);
and U44822 (N_44822,N_42619,N_43711);
nand U44823 (N_44823,N_42045,N_42593);
nand U44824 (N_44824,N_42443,N_42005);
xnor U44825 (N_44825,N_43186,N_43506);
or U44826 (N_44826,N_43045,N_42997);
nor U44827 (N_44827,N_43137,N_43395);
or U44828 (N_44828,N_42004,N_42546);
nand U44829 (N_44829,N_43503,N_43915);
xor U44830 (N_44830,N_43460,N_43554);
or U44831 (N_44831,N_42955,N_43133);
and U44832 (N_44832,N_42727,N_43079);
nor U44833 (N_44833,N_43889,N_42670);
xnor U44834 (N_44834,N_43627,N_42825);
nor U44835 (N_44835,N_43885,N_43346);
or U44836 (N_44836,N_43948,N_42024);
xor U44837 (N_44837,N_43479,N_42284);
nor U44838 (N_44838,N_43393,N_42888);
nand U44839 (N_44839,N_42923,N_42959);
xnor U44840 (N_44840,N_43208,N_43382);
nand U44841 (N_44841,N_43055,N_42421);
or U44842 (N_44842,N_42824,N_42569);
or U44843 (N_44843,N_42148,N_42769);
or U44844 (N_44844,N_43730,N_42934);
and U44845 (N_44845,N_43123,N_42548);
xnor U44846 (N_44846,N_42159,N_42311);
xnor U44847 (N_44847,N_42400,N_42183);
or U44848 (N_44848,N_43624,N_42832);
and U44849 (N_44849,N_42089,N_43569);
xor U44850 (N_44850,N_42108,N_43444);
nor U44851 (N_44851,N_42726,N_43939);
nor U44852 (N_44852,N_43273,N_42329);
xor U44853 (N_44853,N_42547,N_42584);
and U44854 (N_44854,N_43798,N_42644);
and U44855 (N_44855,N_42415,N_42325);
xor U44856 (N_44856,N_42679,N_42433);
or U44857 (N_44857,N_43766,N_42951);
xor U44858 (N_44858,N_43542,N_42061);
xor U44859 (N_44859,N_43307,N_43873);
xor U44860 (N_44860,N_42618,N_43838);
nor U44861 (N_44861,N_43628,N_43567);
and U44862 (N_44862,N_42794,N_42663);
nor U44863 (N_44863,N_42966,N_43718);
nor U44864 (N_44864,N_43080,N_43312);
xor U44865 (N_44865,N_42929,N_42751);
nor U44866 (N_44866,N_42105,N_43027);
nor U44867 (N_44867,N_42023,N_43561);
nor U44868 (N_44868,N_42202,N_42299);
and U44869 (N_44869,N_43541,N_42983);
or U44870 (N_44870,N_42280,N_42752);
and U44871 (N_44871,N_42220,N_42497);
nor U44872 (N_44872,N_43927,N_42508);
nand U44873 (N_44873,N_43013,N_43997);
xor U44874 (N_44874,N_43248,N_42960);
xnor U44875 (N_44875,N_43900,N_42819);
and U44876 (N_44876,N_42599,N_42027);
nand U44877 (N_44877,N_43246,N_43434);
or U44878 (N_44878,N_42256,N_43038);
nand U44879 (N_44879,N_43288,N_43892);
xor U44880 (N_44880,N_43287,N_42039);
nand U44881 (N_44881,N_42596,N_42557);
nor U44882 (N_44882,N_42772,N_43949);
xnor U44883 (N_44883,N_43321,N_43813);
nand U44884 (N_44884,N_42052,N_43059);
nor U44885 (N_44885,N_43188,N_43495);
nor U44886 (N_44886,N_42341,N_43895);
or U44887 (N_44887,N_43751,N_42728);
nand U44888 (N_44888,N_42369,N_43612);
xnor U44889 (N_44889,N_42653,N_42495);
or U44890 (N_44890,N_42364,N_42689);
or U44891 (N_44891,N_42806,N_43025);
nor U44892 (N_44892,N_43453,N_42094);
and U44893 (N_44893,N_43539,N_43790);
nand U44894 (N_44894,N_42597,N_42715);
nor U44895 (N_44895,N_43076,N_42343);
nor U44896 (N_44896,N_42765,N_43244);
and U44897 (N_44897,N_43034,N_42674);
or U44898 (N_44898,N_43697,N_42536);
nand U44899 (N_44899,N_42408,N_42509);
and U44900 (N_44900,N_42191,N_42115);
xor U44901 (N_44901,N_42350,N_43108);
nand U44902 (N_44902,N_42998,N_42111);
nor U44903 (N_44903,N_43178,N_42074);
and U44904 (N_44904,N_43825,N_43496);
and U44905 (N_44905,N_42568,N_43535);
nor U44906 (N_44906,N_42625,N_43230);
xnor U44907 (N_44907,N_43162,N_42445);
nand U44908 (N_44908,N_43768,N_43031);
nand U44909 (N_44909,N_43910,N_42968);
or U44910 (N_44910,N_42719,N_42070);
or U44911 (N_44911,N_42799,N_43486);
xor U44912 (N_44912,N_43714,N_43361);
or U44913 (N_44913,N_42862,N_42245);
xnor U44914 (N_44914,N_43738,N_42606);
or U44915 (N_44915,N_43564,N_43118);
xnor U44916 (N_44916,N_42106,N_42455);
xor U44917 (N_44917,N_43107,N_43832);
nor U44918 (N_44918,N_43588,N_42629);
or U44919 (N_44919,N_42145,N_42602);
nor U44920 (N_44920,N_43682,N_42146);
xnor U44921 (N_44921,N_42224,N_43861);
nor U44922 (N_44922,N_43122,N_43147);
nor U44923 (N_44923,N_43018,N_43911);
nor U44924 (N_44924,N_43863,N_42538);
and U44925 (N_44925,N_43777,N_42157);
and U44926 (N_44926,N_42758,N_42654);
xor U44927 (N_44927,N_42666,N_42818);
and U44928 (N_44928,N_43545,N_42858);
nor U44929 (N_44929,N_43824,N_43127);
and U44930 (N_44930,N_43726,N_42891);
and U44931 (N_44931,N_43553,N_43238);
and U44932 (N_44932,N_43339,N_43482);
xor U44933 (N_44933,N_42130,N_42197);
nand U44934 (N_44934,N_43196,N_42447);
nand U44935 (N_44935,N_43210,N_42121);
or U44936 (N_44936,N_43740,N_42539);
xor U44937 (N_44937,N_42714,N_42748);
nand U44938 (N_44938,N_42702,N_43489);
nand U44939 (N_44939,N_43342,N_42982);
nor U44940 (N_44940,N_43839,N_43240);
nor U44941 (N_44941,N_43854,N_42707);
nand U44942 (N_44942,N_43741,N_42206);
and U44943 (N_44943,N_42992,N_43830);
nor U44944 (N_44944,N_42572,N_43155);
or U44945 (N_44945,N_43699,N_43422);
nor U44946 (N_44946,N_42948,N_43171);
nor U44947 (N_44947,N_42556,N_42828);
and U44948 (N_44948,N_43583,N_43693);
nand U44949 (N_44949,N_42053,N_42164);
xnor U44950 (N_44950,N_43661,N_43305);
xor U44951 (N_44951,N_42680,N_42904);
and U44952 (N_44952,N_43426,N_43827);
or U44953 (N_44953,N_43646,N_43182);
nor U44954 (N_44954,N_43653,N_43912);
nor U44955 (N_44955,N_42687,N_42192);
and U44956 (N_44956,N_42480,N_42469);
and U44957 (N_44957,N_42826,N_43924);
nand U44958 (N_44958,N_42970,N_43831);
xor U44959 (N_44959,N_43619,N_43689);
nand U44960 (N_44960,N_42780,N_42253);
nor U44961 (N_44961,N_42545,N_43115);
nand U44962 (N_44962,N_43302,N_43043);
and U44963 (N_44963,N_42478,N_42611);
xnor U44964 (N_44964,N_43658,N_42032);
nor U44965 (N_44965,N_43272,N_42009);
nor U44966 (N_44966,N_42021,N_43160);
nor U44967 (N_44967,N_42026,N_42656);
xnor U44968 (N_44968,N_42285,N_43345);
or U44969 (N_44969,N_43652,N_43606);
or U44970 (N_44970,N_43872,N_43934);
and U44971 (N_44971,N_43092,N_42448);
xnor U44972 (N_44972,N_42092,N_42530);
and U44973 (N_44973,N_42650,N_42234);
nor U44974 (N_44974,N_43860,N_42855);
xnor U44975 (N_44975,N_42104,N_42073);
or U44976 (N_44976,N_43296,N_42851);
nand U44977 (N_44977,N_43748,N_43664);
and U44978 (N_44978,N_42174,N_42933);
nand U44979 (N_44979,N_42390,N_43728);
or U44980 (N_44980,N_43114,N_42222);
nand U44981 (N_44981,N_42310,N_42198);
xnor U44982 (N_44982,N_43052,N_42505);
or U44983 (N_44983,N_43062,N_43650);
and U44984 (N_44984,N_42218,N_43961);
nor U44985 (N_44985,N_42856,N_43416);
xor U44986 (N_44986,N_42516,N_43072);
or U44987 (N_44987,N_43979,N_43329);
xnor U44988 (N_44988,N_42229,N_42295);
xor U44989 (N_44989,N_42525,N_43840);
nor U44990 (N_44990,N_43083,N_42069);
nand U44991 (N_44991,N_42264,N_43326);
xnor U44992 (N_44992,N_43239,N_43494);
or U44993 (N_44993,N_42051,N_42368);
and U44994 (N_44994,N_42098,N_43440);
and U44995 (N_44995,N_43828,N_43847);
and U44996 (N_44996,N_43810,N_42330);
or U44997 (N_44997,N_43206,N_43235);
nand U44998 (N_44998,N_42286,N_43333);
and U44999 (N_44999,N_43185,N_43113);
nor U45000 (N_45000,N_42441,N_42606);
or U45001 (N_45001,N_42731,N_43051);
nor U45002 (N_45002,N_42812,N_42595);
nor U45003 (N_45003,N_42199,N_43036);
nor U45004 (N_45004,N_43356,N_42225);
nand U45005 (N_45005,N_43668,N_42473);
or U45006 (N_45006,N_42618,N_42550);
nor U45007 (N_45007,N_42388,N_42264);
nor U45008 (N_45008,N_42724,N_42301);
xnor U45009 (N_45009,N_43915,N_43352);
nor U45010 (N_45010,N_42266,N_42906);
nor U45011 (N_45011,N_42818,N_42690);
or U45012 (N_45012,N_42830,N_43820);
nand U45013 (N_45013,N_43047,N_43201);
and U45014 (N_45014,N_42172,N_42596);
or U45015 (N_45015,N_42767,N_43345);
xor U45016 (N_45016,N_42695,N_42275);
and U45017 (N_45017,N_43722,N_42214);
xor U45018 (N_45018,N_43933,N_43662);
and U45019 (N_45019,N_42266,N_42160);
and U45020 (N_45020,N_42238,N_43328);
or U45021 (N_45021,N_42534,N_42795);
or U45022 (N_45022,N_43373,N_43259);
xor U45023 (N_45023,N_43749,N_42047);
and U45024 (N_45024,N_42319,N_42715);
or U45025 (N_45025,N_43633,N_43688);
nor U45026 (N_45026,N_42290,N_42401);
or U45027 (N_45027,N_42837,N_42854);
xor U45028 (N_45028,N_42894,N_42638);
and U45029 (N_45029,N_43958,N_43658);
xnor U45030 (N_45030,N_43296,N_43440);
and U45031 (N_45031,N_42612,N_43858);
and U45032 (N_45032,N_42086,N_42764);
or U45033 (N_45033,N_43905,N_43644);
nor U45034 (N_45034,N_42118,N_42910);
nand U45035 (N_45035,N_42488,N_43136);
nand U45036 (N_45036,N_42171,N_42153);
nand U45037 (N_45037,N_42644,N_43055);
and U45038 (N_45038,N_43271,N_43640);
and U45039 (N_45039,N_42877,N_42461);
or U45040 (N_45040,N_42390,N_42517);
and U45041 (N_45041,N_42126,N_42381);
or U45042 (N_45042,N_42554,N_43574);
xnor U45043 (N_45043,N_42589,N_43541);
nor U45044 (N_45044,N_43567,N_42886);
nor U45045 (N_45045,N_43957,N_43772);
and U45046 (N_45046,N_42211,N_42285);
and U45047 (N_45047,N_42695,N_42838);
nand U45048 (N_45048,N_42820,N_43081);
xor U45049 (N_45049,N_42945,N_42879);
xor U45050 (N_45050,N_42152,N_42145);
or U45051 (N_45051,N_43815,N_42992);
or U45052 (N_45052,N_43945,N_43632);
nor U45053 (N_45053,N_43696,N_43681);
nor U45054 (N_45054,N_42158,N_43782);
nand U45055 (N_45055,N_43903,N_42304);
and U45056 (N_45056,N_42304,N_43817);
or U45057 (N_45057,N_42814,N_42571);
and U45058 (N_45058,N_42994,N_43879);
nor U45059 (N_45059,N_42682,N_43850);
and U45060 (N_45060,N_43145,N_42983);
and U45061 (N_45061,N_43154,N_43723);
nor U45062 (N_45062,N_42767,N_43649);
nor U45063 (N_45063,N_42933,N_43370);
nor U45064 (N_45064,N_42258,N_42904);
or U45065 (N_45065,N_43320,N_43665);
or U45066 (N_45066,N_42233,N_42333);
and U45067 (N_45067,N_43942,N_42554);
xnor U45068 (N_45068,N_42715,N_43789);
xnor U45069 (N_45069,N_43638,N_43728);
and U45070 (N_45070,N_42144,N_43565);
nand U45071 (N_45071,N_43750,N_42653);
nand U45072 (N_45072,N_43401,N_42099);
or U45073 (N_45073,N_42904,N_43169);
nor U45074 (N_45074,N_43628,N_42036);
nor U45075 (N_45075,N_42904,N_42438);
nand U45076 (N_45076,N_42297,N_42132);
nand U45077 (N_45077,N_42465,N_42503);
and U45078 (N_45078,N_43609,N_43865);
and U45079 (N_45079,N_43739,N_43720);
and U45080 (N_45080,N_42733,N_42020);
and U45081 (N_45081,N_43169,N_43957);
and U45082 (N_45082,N_42887,N_43494);
or U45083 (N_45083,N_42107,N_42037);
and U45084 (N_45084,N_42322,N_42220);
nor U45085 (N_45085,N_43456,N_42427);
nor U45086 (N_45086,N_43081,N_43120);
and U45087 (N_45087,N_43345,N_43766);
nand U45088 (N_45088,N_43931,N_43402);
nand U45089 (N_45089,N_43420,N_42608);
or U45090 (N_45090,N_42573,N_43088);
nand U45091 (N_45091,N_42634,N_42535);
nor U45092 (N_45092,N_43252,N_42492);
nor U45093 (N_45093,N_42442,N_43435);
nand U45094 (N_45094,N_42051,N_43310);
nor U45095 (N_45095,N_42256,N_42119);
and U45096 (N_45096,N_42889,N_43650);
or U45097 (N_45097,N_43810,N_43509);
nand U45098 (N_45098,N_43037,N_43722);
xor U45099 (N_45099,N_43268,N_42905);
nor U45100 (N_45100,N_42646,N_43626);
xnor U45101 (N_45101,N_43990,N_42846);
nor U45102 (N_45102,N_42180,N_43485);
nand U45103 (N_45103,N_42969,N_43786);
xor U45104 (N_45104,N_42132,N_43539);
nand U45105 (N_45105,N_42176,N_43801);
or U45106 (N_45106,N_43377,N_43973);
or U45107 (N_45107,N_42393,N_43444);
xnor U45108 (N_45108,N_43032,N_43706);
and U45109 (N_45109,N_43162,N_42756);
nor U45110 (N_45110,N_43410,N_42690);
nand U45111 (N_45111,N_43194,N_42562);
and U45112 (N_45112,N_43263,N_42621);
nand U45113 (N_45113,N_42204,N_42477);
or U45114 (N_45114,N_43915,N_43220);
nor U45115 (N_45115,N_43001,N_42467);
xor U45116 (N_45116,N_42918,N_43695);
xnor U45117 (N_45117,N_42424,N_43453);
and U45118 (N_45118,N_43300,N_42361);
xnor U45119 (N_45119,N_43495,N_43398);
or U45120 (N_45120,N_43951,N_43877);
and U45121 (N_45121,N_43007,N_42130);
nor U45122 (N_45122,N_42345,N_42383);
nand U45123 (N_45123,N_43790,N_42902);
or U45124 (N_45124,N_42985,N_43297);
xor U45125 (N_45125,N_42721,N_43503);
nand U45126 (N_45126,N_42000,N_42193);
and U45127 (N_45127,N_43937,N_43975);
and U45128 (N_45128,N_43963,N_42675);
xor U45129 (N_45129,N_43326,N_42887);
xnor U45130 (N_45130,N_43700,N_43509);
nand U45131 (N_45131,N_42519,N_42810);
nand U45132 (N_45132,N_42708,N_43102);
nor U45133 (N_45133,N_42009,N_43554);
nand U45134 (N_45134,N_42939,N_43123);
and U45135 (N_45135,N_43643,N_42264);
or U45136 (N_45136,N_42088,N_43063);
nand U45137 (N_45137,N_42872,N_42102);
or U45138 (N_45138,N_43911,N_42691);
nand U45139 (N_45139,N_43686,N_43736);
nor U45140 (N_45140,N_43492,N_43688);
nand U45141 (N_45141,N_42433,N_43823);
nor U45142 (N_45142,N_42681,N_42743);
nand U45143 (N_45143,N_43385,N_43968);
nand U45144 (N_45144,N_42439,N_42277);
xor U45145 (N_45145,N_42694,N_43569);
or U45146 (N_45146,N_42534,N_43413);
nor U45147 (N_45147,N_43330,N_43961);
and U45148 (N_45148,N_42847,N_42652);
nand U45149 (N_45149,N_42390,N_42453);
nand U45150 (N_45150,N_43538,N_42443);
nor U45151 (N_45151,N_42421,N_42142);
nor U45152 (N_45152,N_42160,N_43727);
nand U45153 (N_45153,N_42494,N_42412);
nand U45154 (N_45154,N_43339,N_43547);
and U45155 (N_45155,N_42870,N_42152);
nand U45156 (N_45156,N_42909,N_43985);
or U45157 (N_45157,N_43936,N_43799);
nand U45158 (N_45158,N_43791,N_42209);
nand U45159 (N_45159,N_42439,N_43882);
or U45160 (N_45160,N_42242,N_42663);
nand U45161 (N_45161,N_43910,N_42138);
and U45162 (N_45162,N_42137,N_42202);
nor U45163 (N_45163,N_43263,N_43463);
xnor U45164 (N_45164,N_43587,N_43220);
or U45165 (N_45165,N_43783,N_42434);
nand U45166 (N_45166,N_43032,N_42574);
nor U45167 (N_45167,N_43593,N_43466);
and U45168 (N_45168,N_42141,N_43255);
and U45169 (N_45169,N_43313,N_43733);
nand U45170 (N_45170,N_42776,N_42685);
or U45171 (N_45171,N_43042,N_42073);
and U45172 (N_45172,N_43867,N_42143);
nand U45173 (N_45173,N_43854,N_43029);
or U45174 (N_45174,N_43331,N_42697);
nor U45175 (N_45175,N_42246,N_43719);
nand U45176 (N_45176,N_42447,N_42036);
nand U45177 (N_45177,N_43892,N_43838);
or U45178 (N_45178,N_42711,N_43599);
or U45179 (N_45179,N_43546,N_43068);
and U45180 (N_45180,N_43929,N_43171);
and U45181 (N_45181,N_43680,N_43172);
xnor U45182 (N_45182,N_42211,N_42442);
and U45183 (N_45183,N_42435,N_43184);
xnor U45184 (N_45184,N_42007,N_42642);
nand U45185 (N_45185,N_42688,N_43840);
xnor U45186 (N_45186,N_43492,N_43778);
nand U45187 (N_45187,N_42797,N_42815);
xor U45188 (N_45188,N_42973,N_42767);
and U45189 (N_45189,N_42118,N_42636);
or U45190 (N_45190,N_43628,N_42563);
nor U45191 (N_45191,N_42266,N_43133);
and U45192 (N_45192,N_43206,N_42490);
nor U45193 (N_45193,N_43308,N_42112);
or U45194 (N_45194,N_42328,N_42749);
xnor U45195 (N_45195,N_43062,N_43689);
xnor U45196 (N_45196,N_43274,N_42407);
and U45197 (N_45197,N_42455,N_43504);
nand U45198 (N_45198,N_42019,N_43537);
and U45199 (N_45199,N_43292,N_43051);
nor U45200 (N_45200,N_42513,N_42740);
nand U45201 (N_45201,N_42253,N_43526);
nor U45202 (N_45202,N_42275,N_43335);
and U45203 (N_45203,N_43255,N_43600);
xor U45204 (N_45204,N_43613,N_42392);
nand U45205 (N_45205,N_42650,N_42757);
and U45206 (N_45206,N_42383,N_42001);
or U45207 (N_45207,N_42573,N_43874);
and U45208 (N_45208,N_43121,N_43947);
xnor U45209 (N_45209,N_43977,N_42087);
nand U45210 (N_45210,N_42800,N_42822);
and U45211 (N_45211,N_43790,N_42705);
xnor U45212 (N_45212,N_43823,N_42452);
nor U45213 (N_45213,N_42957,N_43049);
xnor U45214 (N_45214,N_42890,N_42247);
nor U45215 (N_45215,N_42319,N_43299);
or U45216 (N_45216,N_43394,N_42631);
and U45217 (N_45217,N_43618,N_43598);
or U45218 (N_45218,N_42497,N_42964);
nand U45219 (N_45219,N_43912,N_42608);
and U45220 (N_45220,N_43547,N_43450);
nand U45221 (N_45221,N_42295,N_43514);
and U45222 (N_45222,N_43973,N_42823);
xor U45223 (N_45223,N_42126,N_43477);
nand U45224 (N_45224,N_43831,N_42016);
nand U45225 (N_45225,N_43378,N_42385);
or U45226 (N_45226,N_42977,N_43563);
xnor U45227 (N_45227,N_42954,N_43520);
or U45228 (N_45228,N_42666,N_42711);
nor U45229 (N_45229,N_43974,N_43561);
xnor U45230 (N_45230,N_42135,N_43966);
xor U45231 (N_45231,N_43657,N_42671);
xnor U45232 (N_45232,N_43442,N_43181);
nor U45233 (N_45233,N_43087,N_42905);
and U45234 (N_45234,N_43252,N_43452);
nor U45235 (N_45235,N_43815,N_42557);
or U45236 (N_45236,N_42261,N_43898);
xor U45237 (N_45237,N_43094,N_43664);
nand U45238 (N_45238,N_42926,N_43061);
and U45239 (N_45239,N_42221,N_43193);
nand U45240 (N_45240,N_43381,N_43788);
xnor U45241 (N_45241,N_42129,N_43178);
and U45242 (N_45242,N_43832,N_43294);
and U45243 (N_45243,N_42239,N_42718);
nor U45244 (N_45244,N_42800,N_42904);
nand U45245 (N_45245,N_42555,N_43878);
and U45246 (N_45246,N_42689,N_43673);
nand U45247 (N_45247,N_42684,N_42403);
and U45248 (N_45248,N_42944,N_42886);
xnor U45249 (N_45249,N_42443,N_42888);
nand U45250 (N_45250,N_42650,N_42009);
nor U45251 (N_45251,N_42594,N_42421);
nor U45252 (N_45252,N_43271,N_42386);
or U45253 (N_45253,N_43111,N_42116);
xor U45254 (N_45254,N_42324,N_43596);
nand U45255 (N_45255,N_42761,N_42506);
nand U45256 (N_45256,N_42705,N_43853);
xnor U45257 (N_45257,N_43783,N_42271);
nor U45258 (N_45258,N_43513,N_43016);
nand U45259 (N_45259,N_42713,N_43278);
nor U45260 (N_45260,N_42904,N_42933);
or U45261 (N_45261,N_43091,N_43932);
nor U45262 (N_45262,N_43648,N_43005);
or U45263 (N_45263,N_43188,N_42769);
xor U45264 (N_45264,N_43621,N_43264);
nand U45265 (N_45265,N_42098,N_42564);
nand U45266 (N_45266,N_43716,N_43890);
nand U45267 (N_45267,N_42502,N_43807);
xor U45268 (N_45268,N_43354,N_42174);
nor U45269 (N_45269,N_43957,N_42070);
xnor U45270 (N_45270,N_43082,N_42032);
or U45271 (N_45271,N_43307,N_43351);
and U45272 (N_45272,N_42131,N_43215);
nor U45273 (N_45273,N_43576,N_43604);
nand U45274 (N_45274,N_43465,N_43754);
and U45275 (N_45275,N_43224,N_42855);
or U45276 (N_45276,N_43374,N_43059);
xnor U45277 (N_45277,N_42459,N_42331);
nand U45278 (N_45278,N_43459,N_43412);
xor U45279 (N_45279,N_42260,N_42660);
and U45280 (N_45280,N_43246,N_42889);
xnor U45281 (N_45281,N_43269,N_43715);
nor U45282 (N_45282,N_43976,N_43614);
nor U45283 (N_45283,N_43439,N_42894);
nor U45284 (N_45284,N_42347,N_43558);
nor U45285 (N_45285,N_43754,N_42212);
or U45286 (N_45286,N_43280,N_42244);
nor U45287 (N_45287,N_42107,N_42064);
or U45288 (N_45288,N_43366,N_42491);
nor U45289 (N_45289,N_42668,N_43353);
xnor U45290 (N_45290,N_42138,N_42579);
nand U45291 (N_45291,N_43810,N_42476);
and U45292 (N_45292,N_43637,N_42299);
xnor U45293 (N_45293,N_42679,N_43986);
or U45294 (N_45294,N_43809,N_43480);
or U45295 (N_45295,N_42898,N_42952);
or U45296 (N_45296,N_42583,N_42694);
xor U45297 (N_45297,N_43444,N_42428);
or U45298 (N_45298,N_43423,N_43851);
and U45299 (N_45299,N_43714,N_43884);
xnor U45300 (N_45300,N_43321,N_42816);
or U45301 (N_45301,N_43892,N_42719);
or U45302 (N_45302,N_43183,N_42125);
nand U45303 (N_45303,N_43052,N_42956);
or U45304 (N_45304,N_43407,N_42803);
xor U45305 (N_45305,N_42344,N_43395);
nor U45306 (N_45306,N_43863,N_42748);
and U45307 (N_45307,N_42753,N_43294);
and U45308 (N_45308,N_43904,N_43996);
and U45309 (N_45309,N_43354,N_43595);
nand U45310 (N_45310,N_43981,N_42644);
xnor U45311 (N_45311,N_43770,N_42878);
xnor U45312 (N_45312,N_42597,N_43943);
or U45313 (N_45313,N_42227,N_42443);
or U45314 (N_45314,N_42914,N_43990);
and U45315 (N_45315,N_43100,N_43596);
xnor U45316 (N_45316,N_43920,N_42126);
or U45317 (N_45317,N_43429,N_43735);
xor U45318 (N_45318,N_42501,N_42708);
xnor U45319 (N_45319,N_43120,N_43734);
xor U45320 (N_45320,N_42757,N_42474);
or U45321 (N_45321,N_43104,N_42386);
nand U45322 (N_45322,N_42978,N_42268);
nand U45323 (N_45323,N_42071,N_42678);
xnor U45324 (N_45324,N_42790,N_43180);
xnor U45325 (N_45325,N_42331,N_42416);
nor U45326 (N_45326,N_42517,N_42004);
and U45327 (N_45327,N_42491,N_43805);
nor U45328 (N_45328,N_42382,N_43090);
nand U45329 (N_45329,N_43772,N_43131);
or U45330 (N_45330,N_43745,N_42233);
nor U45331 (N_45331,N_43984,N_42293);
or U45332 (N_45332,N_43007,N_43651);
and U45333 (N_45333,N_42304,N_43713);
nor U45334 (N_45334,N_42876,N_43697);
and U45335 (N_45335,N_42636,N_43980);
xor U45336 (N_45336,N_43152,N_42396);
or U45337 (N_45337,N_43660,N_43842);
nand U45338 (N_45338,N_43336,N_43290);
and U45339 (N_45339,N_43799,N_42086);
or U45340 (N_45340,N_43141,N_43717);
or U45341 (N_45341,N_42498,N_42881);
nand U45342 (N_45342,N_42550,N_43305);
nor U45343 (N_45343,N_43206,N_42474);
nand U45344 (N_45344,N_42756,N_42544);
or U45345 (N_45345,N_42037,N_43366);
nand U45346 (N_45346,N_43615,N_43108);
or U45347 (N_45347,N_43553,N_43738);
or U45348 (N_45348,N_43428,N_43304);
nand U45349 (N_45349,N_43783,N_43226);
or U45350 (N_45350,N_42997,N_42989);
xnor U45351 (N_45351,N_43418,N_42972);
or U45352 (N_45352,N_43480,N_43160);
nand U45353 (N_45353,N_42251,N_43306);
or U45354 (N_45354,N_43657,N_42071);
nand U45355 (N_45355,N_42937,N_42004);
xor U45356 (N_45356,N_42813,N_42381);
xor U45357 (N_45357,N_42657,N_42827);
and U45358 (N_45358,N_42693,N_43793);
nand U45359 (N_45359,N_43705,N_43191);
xnor U45360 (N_45360,N_43469,N_43374);
nor U45361 (N_45361,N_42112,N_43137);
or U45362 (N_45362,N_42693,N_42780);
nor U45363 (N_45363,N_43545,N_42266);
or U45364 (N_45364,N_42575,N_42229);
or U45365 (N_45365,N_42921,N_43104);
nor U45366 (N_45366,N_43782,N_43807);
nor U45367 (N_45367,N_42784,N_43781);
and U45368 (N_45368,N_43194,N_42201);
xnor U45369 (N_45369,N_42625,N_42777);
or U45370 (N_45370,N_42658,N_43433);
nand U45371 (N_45371,N_43062,N_42430);
xor U45372 (N_45372,N_42151,N_42697);
xor U45373 (N_45373,N_42408,N_42785);
nand U45374 (N_45374,N_42306,N_42272);
and U45375 (N_45375,N_43711,N_42665);
or U45376 (N_45376,N_43816,N_42579);
nor U45377 (N_45377,N_42649,N_43305);
nor U45378 (N_45378,N_43256,N_42055);
nand U45379 (N_45379,N_43103,N_43749);
or U45380 (N_45380,N_42232,N_42907);
and U45381 (N_45381,N_42847,N_43244);
nor U45382 (N_45382,N_42915,N_43649);
nor U45383 (N_45383,N_43518,N_42071);
nand U45384 (N_45384,N_42542,N_42393);
xor U45385 (N_45385,N_42822,N_43939);
xor U45386 (N_45386,N_42833,N_42030);
nand U45387 (N_45387,N_42289,N_42880);
or U45388 (N_45388,N_43319,N_42283);
and U45389 (N_45389,N_42819,N_43166);
nand U45390 (N_45390,N_42510,N_43058);
or U45391 (N_45391,N_43530,N_42404);
xnor U45392 (N_45392,N_42191,N_42936);
nor U45393 (N_45393,N_43967,N_42728);
and U45394 (N_45394,N_43243,N_42361);
nand U45395 (N_45395,N_42425,N_43744);
xor U45396 (N_45396,N_42895,N_42603);
xor U45397 (N_45397,N_42118,N_42209);
xnor U45398 (N_45398,N_43477,N_42623);
nor U45399 (N_45399,N_42539,N_43315);
xor U45400 (N_45400,N_42818,N_43914);
nand U45401 (N_45401,N_43205,N_43136);
and U45402 (N_45402,N_43859,N_43360);
nand U45403 (N_45403,N_42367,N_42251);
xnor U45404 (N_45404,N_43844,N_42107);
nand U45405 (N_45405,N_43213,N_42959);
or U45406 (N_45406,N_43538,N_42580);
and U45407 (N_45407,N_43296,N_42748);
or U45408 (N_45408,N_42828,N_43054);
xnor U45409 (N_45409,N_43888,N_43720);
or U45410 (N_45410,N_43266,N_42016);
xnor U45411 (N_45411,N_42535,N_43717);
and U45412 (N_45412,N_43020,N_42157);
and U45413 (N_45413,N_43206,N_42702);
and U45414 (N_45414,N_42564,N_43431);
or U45415 (N_45415,N_43383,N_43437);
or U45416 (N_45416,N_42286,N_43313);
nor U45417 (N_45417,N_43830,N_42499);
xnor U45418 (N_45418,N_43242,N_43553);
and U45419 (N_45419,N_42239,N_43393);
nand U45420 (N_45420,N_43797,N_43013);
or U45421 (N_45421,N_42494,N_43385);
nor U45422 (N_45422,N_43982,N_43797);
and U45423 (N_45423,N_43553,N_42030);
xnor U45424 (N_45424,N_42211,N_42580);
and U45425 (N_45425,N_43982,N_43131);
nand U45426 (N_45426,N_43082,N_42191);
xnor U45427 (N_45427,N_42832,N_42072);
xnor U45428 (N_45428,N_42450,N_43904);
nand U45429 (N_45429,N_43156,N_43437);
or U45430 (N_45430,N_43468,N_42310);
nor U45431 (N_45431,N_43607,N_43771);
and U45432 (N_45432,N_43122,N_43600);
xnor U45433 (N_45433,N_43970,N_42328);
xnor U45434 (N_45434,N_42549,N_42846);
and U45435 (N_45435,N_42923,N_43748);
nor U45436 (N_45436,N_43885,N_43385);
or U45437 (N_45437,N_43108,N_42383);
and U45438 (N_45438,N_42179,N_43677);
nor U45439 (N_45439,N_42767,N_43076);
xnor U45440 (N_45440,N_42503,N_42221);
nand U45441 (N_45441,N_43267,N_43183);
and U45442 (N_45442,N_42959,N_42972);
xnor U45443 (N_45443,N_42661,N_42411);
or U45444 (N_45444,N_43220,N_42088);
nor U45445 (N_45445,N_43909,N_42802);
nand U45446 (N_45446,N_42970,N_43701);
or U45447 (N_45447,N_42339,N_43060);
xnor U45448 (N_45448,N_43370,N_43044);
xnor U45449 (N_45449,N_42404,N_43882);
or U45450 (N_45450,N_42389,N_43068);
and U45451 (N_45451,N_43361,N_43764);
nor U45452 (N_45452,N_42794,N_42034);
nor U45453 (N_45453,N_43892,N_42853);
nor U45454 (N_45454,N_43347,N_43044);
nand U45455 (N_45455,N_43664,N_42389);
xnor U45456 (N_45456,N_43857,N_43930);
nor U45457 (N_45457,N_43525,N_42651);
and U45458 (N_45458,N_43212,N_43016);
nand U45459 (N_45459,N_42835,N_42981);
and U45460 (N_45460,N_42809,N_43198);
and U45461 (N_45461,N_42036,N_42817);
nor U45462 (N_45462,N_42602,N_42635);
nor U45463 (N_45463,N_42073,N_42425);
nor U45464 (N_45464,N_43243,N_42238);
and U45465 (N_45465,N_43569,N_43007);
nor U45466 (N_45466,N_42392,N_43147);
nand U45467 (N_45467,N_43985,N_42877);
nor U45468 (N_45468,N_42355,N_42447);
and U45469 (N_45469,N_42025,N_42525);
or U45470 (N_45470,N_42945,N_43957);
and U45471 (N_45471,N_43385,N_43539);
nor U45472 (N_45472,N_43007,N_43632);
or U45473 (N_45473,N_43331,N_42268);
or U45474 (N_45474,N_42959,N_42230);
xor U45475 (N_45475,N_43398,N_43385);
nor U45476 (N_45476,N_42811,N_43259);
or U45477 (N_45477,N_42800,N_42868);
xor U45478 (N_45478,N_42413,N_42941);
and U45479 (N_45479,N_42879,N_42342);
nand U45480 (N_45480,N_42721,N_42377);
and U45481 (N_45481,N_42327,N_43113);
nor U45482 (N_45482,N_43904,N_43187);
nand U45483 (N_45483,N_43605,N_43213);
nand U45484 (N_45484,N_43217,N_42789);
nand U45485 (N_45485,N_43332,N_43739);
or U45486 (N_45486,N_42965,N_42352);
and U45487 (N_45487,N_43767,N_43458);
nand U45488 (N_45488,N_43176,N_42207);
nand U45489 (N_45489,N_42722,N_43152);
nand U45490 (N_45490,N_43211,N_43223);
xor U45491 (N_45491,N_42049,N_43931);
or U45492 (N_45492,N_43663,N_43402);
xor U45493 (N_45493,N_42240,N_42923);
nand U45494 (N_45494,N_42882,N_42972);
xnor U45495 (N_45495,N_42629,N_43265);
or U45496 (N_45496,N_42191,N_42924);
xnor U45497 (N_45497,N_43934,N_43426);
nand U45498 (N_45498,N_43192,N_43308);
nor U45499 (N_45499,N_43217,N_43292);
nand U45500 (N_45500,N_42725,N_43590);
nand U45501 (N_45501,N_42683,N_43360);
and U45502 (N_45502,N_43508,N_43963);
xnor U45503 (N_45503,N_42972,N_43037);
or U45504 (N_45504,N_42376,N_43335);
or U45505 (N_45505,N_43740,N_43375);
xnor U45506 (N_45506,N_42073,N_42776);
and U45507 (N_45507,N_43282,N_42243);
nand U45508 (N_45508,N_42554,N_43250);
xor U45509 (N_45509,N_43986,N_42464);
xnor U45510 (N_45510,N_42242,N_42459);
and U45511 (N_45511,N_42975,N_43863);
and U45512 (N_45512,N_42555,N_43785);
nand U45513 (N_45513,N_42111,N_42729);
xor U45514 (N_45514,N_43876,N_42277);
or U45515 (N_45515,N_42455,N_43947);
or U45516 (N_45516,N_42432,N_43489);
nand U45517 (N_45517,N_42601,N_43935);
and U45518 (N_45518,N_43803,N_42345);
nand U45519 (N_45519,N_43844,N_42290);
and U45520 (N_45520,N_42210,N_43585);
or U45521 (N_45521,N_42561,N_43272);
xnor U45522 (N_45522,N_42153,N_42572);
and U45523 (N_45523,N_42731,N_42621);
nand U45524 (N_45524,N_43532,N_43317);
xor U45525 (N_45525,N_42103,N_43821);
nor U45526 (N_45526,N_42125,N_43827);
or U45527 (N_45527,N_43465,N_42210);
nand U45528 (N_45528,N_43789,N_42849);
xor U45529 (N_45529,N_42472,N_43742);
nand U45530 (N_45530,N_43929,N_42683);
or U45531 (N_45531,N_42858,N_42098);
and U45532 (N_45532,N_42542,N_42666);
or U45533 (N_45533,N_42431,N_42126);
or U45534 (N_45534,N_42865,N_43244);
nor U45535 (N_45535,N_43704,N_43290);
xor U45536 (N_45536,N_42031,N_43409);
or U45537 (N_45537,N_42813,N_42246);
and U45538 (N_45538,N_43735,N_43150);
or U45539 (N_45539,N_42996,N_43322);
and U45540 (N_45540,N_42037,N_42058);
or U45541 (N_45541,N_43236,N_43453);
or U45542 (N_45542,N_43910,N_42020);
nor U45543 (N_45543,N_43899,N_43166);
xor U45544 (N_45544,N_43035,N_42380);
nand U45545 (N_45545,N_42836,N_43879);
xnor U45546 (N_45546,N_43973,N_42860);
and U45547 (N_45547,N_43842,N_42741);
nand U45548 (N_45548,N_43925,N_43103);
nand U45549 (N_45549,N_43077,N_43074);
xnor U45550 (N_45550,N_43963,N_43064);
nand U45551 (N_45551,N_43073,N_42795);
or U45552 (N_45552,N_43670,N_43477);
nor U45553 (N_45553,N_43030,N_42424);
nor U45554 (N_45554,N_43124,N_43342);
nand U45555 (N_45555,N_43212,N_43509);
nor U45556 (N_45556,N_42079,N_43178);
and U45557 (N_45557,N_42064,N_43919);
nor U45558 (N_45558,N_43732,N_42960);
nand U45559 (N_45559,N_43396,N_43607);
nor U45560 (N_45560,N_42628,N_42360);
nand U45561 (N_45561,N_42069,N_43496);
and U45562 (N_45562,N_43533,N_42656);
xor U45563 (N_45563,N_43676,N_43733);
nand U45564 (N_45564,N_42163,N_43187);
and U45565 (N_45565,N_43460,N_43396);
or U45566 (N_45566,N_43109,N_43730);
or U45567 (N_45567,N_43522,N_43287);
xor U45568 (N_45568,N_42880,N_42907);
xnor U45569 (N_45569,N_42886,N_43518);
or U45570 (N_45570,N_43356,N_42910);
and U45571 (N_45571,N_42147,N_42435);
nand U45572 (N_45572,N_43598,N_43850);
or U45573 (N_45573,N_43849,N_43332);
nor U45574 (N_45574,N_43477,N_42564);
and U45575 (N_45575,N_43594,N_43496);
nand U45576 (N_45576,N_42360,N_42137);
nand U45577 (N_45577,N_42012,N_43807);
or U45578 (N_45578,N_43143,N_43872);
nand U45579 (N_45579,N_42144,N_42658);
nor U45580 (N_45580,N_43649,N_43288);
xor U45581 (N_45581,N_43780,N_42393);
and U45582 (N_45582,N_43806,N_43662);
and U45583 (N_45583,N_43658,N_42773);
nand U45584 (N_45584,N_43461,N_43467);
or U45585 (N_45585,N_42294,N_43373);
nor U45586 (N_45586,N_43957,N_43205);
nor U45587 (N_45587,N_43949,N_42186);
or U45588 (N_45588,N_43930,N_42999);
xor U45589 (N_45589,N_43793,N_43232);
nor U45590 (N_45590,N_42087,N_42673);
or U45591 (N_45591,N_43440,N_43805);
nand U45592 (N_45592,N_42918,N_42859);
or U45593 (N_45593,N_42400,N_43666);
nor U45594 (N_45594,N_43693,N_42464);
nand U45595 (N_45595,N_42371,N_42041);
nand U45596 (N_45596,N_43139,N_42007);
xor U45597 (N_45597,N_43536,N_43246);
or U45598 (N_45598,N_42046,N_43484);
and U45599 (N_45599,N_42841,N_43758);
nor U45600 (N_45600,N_42253,N_42955);
nor U45601 (N_45601,N_43436,N_42037);
and U45602 (N_45602,N_43635,N_42667);
nand U45603 (N_45603,N_42602,N_42960);
and U45604 (N_45604,N_43519,N_42011);
or U45605 (N_45605,N_42383,N_42118);
nand U45606 (N_45606,N_42050,N_43162);
or U45607 (N_45607,N_43028,N_42772);
nand U45608 (N_45608,N_42692,N_43412);
nand U45609 (N_45609,N_43582,N_43557);
and U45610 (N_45610,N_42698,N_42899);
or U45611 (N_45611,N_43166,N_43114);
nand U45612 (N_45612,N_43365,N_42226);
xor U45613 (N_45613,N_42891,N_43596);
nor U45614 (N_45614,N_43728,N_43865);
nand U45615 (N_45615,N_42572,N_43411);
xnor U45616 (N_45616,N_43432,N_42622);
nand U45617 (N_45617,N_42629,N_42104);
and U45618 (N_45618,N_43859,N_43523);
nor U45619 (N_45619,N_42342,N_43399);
or U45620 (N_45620,N_43180,N_42635);
nor U45621 (N_45621,N_43416,N_43360);
xnor U45622 (N_45622,N_43937,N_42342);
nor U45623 (N_45623,N_43293,N_43660);
xor U45624 (N_45624,N_42992,N_43548);
xor U45625 (N_45625,N_42840,N_42113);
nand U45626 (N_45626,N_42999,N_42796);
and U45627 (N_45627,N_43809,N_43339);
nand U45628 (N_45628,N_43026,N_43709);
and U45629 (N_45629,N_42575,N_42233);
nand U45630 (N_45630,N_42253,N_43424);
nor U45631 (N_45631,N_42983,N_43051);
xor U45632 (N_45632,N_43411,N_42152);
nand U45633 (N_45633,N_43405,N_43794);
nand U45634 (N_45634,N_43178,N_42072);
xnor U45635 (N_45635,N_42914,N_43168);
nand U45636 (N_45636,N_42935,N_42629);
nor U45637 (N_45637,N_42856,N_43713);
nor U45638 (N_45638,N_42844,N_42028);
nand U45639 (N_45639,N_42703,N_42255);
nor U45640 (N_45640,N_42921,N_42015);
nor U45641 (N_45641,N_43338,N_43633);
or U45642 (N_45642,N_42382,N_43461);
nor U45643 (N_45643,N_42412,N_43775);
nor U45644 (N_45644,N_43879,N_42397);
nand U45645 (N_45645,N_42599,N_43683);
xnor U45646 (N_45646,N_42988,N_42889);
nor U45647 (N_45647,N_43743,N_43521);
and U45648 (N_45648,N_42820,N_43583);
and U45649 (N_45649,N_42843,N_43882);
or U45650 (N_45650,N_43976,N_42317);
xor U45651 (N_45651,N_42521,N_43405);
nand U45652 (N_45652,N_43637,N_42927);
and U45653 (N_45653,N_42257,N_43498);
or U45654 (N_45654,N_43679,N_43958);
and U45655 (N_45655,N_42709,N_42608);
nor U45656 (N_45656,N_42140,N_42958);
or U45657 (N_45657,N_42454,N_43897);
and U45658 (N_45658,N_42808,N_42648);
xnor U45659 (N_45659,N_43283,N_43911);
nand U45660 (N_45660,N_43631,N_42388);
and U45661 (N_45661,N_43757,N_42340);
nor U45662 (N_45662,N_42200,N_43148);
xor U45663 (N_45663,N_43259,N_43683);
nor U45664 (N_45664,N_42077,N_43427);
nand U45665 (N_45665,N_42677,N_43821);
and U45666 (N_45666,N_42720,N_42357);
nor U45667 (N_45667,N_43260,N_42668);
and U45668 (N_45668,N_42823,N_43632);
nor U45669 (N_45669,N_42010,N_42642);
nor U45670 (N_45670,N_43387,N_42023);
and U45671 (N_45671,N_42906,N_43177);
nand U45672 (N_45672,N_43201,N_43193);
or U45673 (N_45673,N_43861,N_43677);
or U45674 (N_45674,N_43197,N_43482);
nand U45675 (N_45675,N_42085,N_43041);
nor U45676 (N_45676,N_42107,N_43778);
and U45677 (N_45677,N_43992,N_42063);
xor U45678 (N_45678,N_43645,N_42786);
and U45679 (N_45679,N_43128,N_42435);
and U45680 (N_45680,N_42387,N_42294);
nand U45681 (N_45681,N_42318,N_42249);
xor U45682 (N_45682,N_42711,N_43074);
and U45683 (N_45683,N_42267,N_43783);
or U45684 (N_45684,N_42960,N_43371);
and U45685 (N_45685,N_43625,N_42625);
nand U45686 (N_45686,N_43856,N_42666);
nand U45687 (N_45687,N_43634,N_42438);
and U45688 (N_45688,N_43680,N_43900);
nand U45689 (N_45689,N_43328,N_42935);
xnor U45690 (N_45690,N_42507,N_42950);
and U45691 (N_45691,N_42079,N_42713);
or U45692 (N_45692,N_42782,N_42770);
nand U45693 (N_45693,N_42858,N_43478);
nand U45694 (N_45694,N_43416,N_42589);
nand U45695 (N_45695,N_42525,N_42202);
xnor U45696 (N_45696,N_43954,N_43806);
or U45697 (N_45697,N_42719,N_42681);
or U45698 (N_45698,N_43037,N_43684);
and U45699 (N_45699,N_42529,N_43521);
or U45700 (N_45700,N_42403,N_43344);
xor U45701 (N_45701,N_43168,N_43291);
or U45702 (N_45702,N_42753,N_42519);
nor U45703 (N_45703,N_43426,N_42818);
xnor U45704 (N_45704,N_43531,N_43103);
and U45705 (N_45705,N_42139,N_42274);
and U45706 (N_45706,N_43395,N_42119);
and U45707 (N_45707,N_42966,N_42582);
nand U45708 (N_45708,N_42330,N_43964);
nor U45709 (N_45709,N_43010,N_43821);
xor U45710 (N_45710,N_42516,N_42192);
nor U45711 (N_45711,N_42908,N_43053);
or U45712 (N_45712,N_43869,N_43795);
nand U45713 (N_45713,N_43027,N_42577);
xnor U45714 (N_45714,N_42112,N_42279);
xnor U45715 (N_45715,N_43469,N_43174);
nand U45716 (N_45716,N_42369,N_43910);
and U45717 (N_45717,N_43957,N_42240);
nor U45718 (N_45718,N_42265,N_43337);
nor U45719 (N_45719,N_42870,N_43243);
xnor U45720 (N_45720,N_43937,N_42497);
and U45721 (N_45721,N_43805,N_42323);
nor U45722 (N_45722,N_43967,N_43840);
xnor U45723 (N_45723,N_42999,N_43656);
and U45724 (N_45724,N_42602,N_42146);
and U45725 (N_45725,N_43593,N_43699);
nor U45726 (N_45726,N_43395,N_42979);
nand U45727 (N_45727,N_43562,N_43725);
or U45728 (N_45728,N_43472,N_43295);
or U45729 (N_45729,N_43149,N_42299);
nand U45730 (N_45730,N_42497,N_43901);
and U45731 (N_45731,N_43978,N_42782);
nand U45732 (N_45732,N_42348,N_42439);
nand U45733 (N_45733,N_42660,N_42464);
or U45734 (N_45734,N_43775,N_42301);
and U45735 (N_45735,N_43517,N_43748);
nand U45736 (N_45736,N_43967,N_43762);
nand U45737 (N_45737,N_42593,N_43143);
nor U45738 (N_45738,N_42895,N_42229);
xnor U45739 (N_45739,N_42966,N_42328);
or U45740 (N_45740,N_42039,N_42955);
xor U45741 (N_45741,N_43875,N_43376);
and U45742 (N_45742,N_43790,N_42427);
nor U45743 (N_45743,N_42736,N_43828);
nand U45744 (N_45744,N_43317,N_43005);
or U45745 (N_45745,N_43886,N_43842);
and U45746 (N_45746,N_43507,N_43527);
xor U45747 (N_45747,N_42283,N_43287);
or U45748 (N_45748,N_43356,N_42728);
nand U45749 (N_45749,N_42386,N_42085);
xnor U45750 (N_45750,N_42473,N_42764);
and U45751 (N_45751,N_43642,N_42278);
nand U45752 (N_45752,N_43255,N_42917);
or U45753 (N_45753,N_43180,N_43394);
xor U45754 (N_45754,N_42240,N_42780);
xor U45755 (N_45755,N_42304,N_43715);
xor U45756 (N_45756,N_42676,N_42643);
xnor U45757 (N_45757,N_43594,N_42228);
nand U45758 (N_45758,N_43847,N_42759);
nand U45759 (N_45759,N_42715,N_42994);
and U45760 (N_45760,N_42148,N_43146);
or U45761 (N_45761,N_43298,N_42926);
nand U45762 (N_45762,N_43190,N_43457);
nor U45763 (N_45763,N_43869,N_42511);
nor U45764 (N_45764,N_42514,N_43607);
nor U45765 (N_45765,N_42984,N_43915);
and U45766 (N_45766,N_43701,N_42957);
and U45767 (N_45767,N_43577,N_43166);
or U45768 (N_45768,N_42084,N_42936);
nor U45769 (N_45769,N_43031,N_43483);
and U45770 (N_45770,N_42745,N_43662);
and U45771 (N_45771,N_43256,N_43577);
and U45772 (N_45772,N_43956,N_43172);
xnor U45773 (N_45773,N_42404,N_43664);
and U45774 (N_45774,N_42564,N_42379);
nand U45775 (N_45775,N_43524,N_43984);
or U45776 (N_45776,N_43907,N_43506);
and U45777 (N_45777,N_42240,N_42499);
or U45778 (N_45778,N_42384,N_42812);
and U45779 (N_45779,N_43770,N_42717);
xnor U45780 (N_45780,N_42817,N_43378);
or U45781 (N_45781,N_43041,N_42050);
nand U45782 (N_45782,N_42346,N_42636);
nor U45783 (N_45783,N_43115,N_43359);
and U45784 (N_45784,N_42560,N_43721);
nor U45785 (N_45785,N_43365,N_43649);
and U45786 (N_45786,N_42535,N_42200);
or U45787 (N_45787,N_42834,N_43115);
nand U45788 (N_45788,N_42498,N_42855);
xor U45789 (N_45789,N_42011,N_43424);
or U45790 (N_45790,N_43800,N_42833);
nor U45791 (N_45791,N_42412,N_42838);
xor U45792 (N_45792,N_43226,N_43236);
nand U45793 (N_45793,N_42456,N_43806);
xnor U45794 (N_45794,N_43866,N_43587);
or U45795 (N_45795,N_42135,N_43660);
nand U45796 (N_45796,N_42082,N_43546);
nand U45797 (N_45797,N_42374,N_43864);
and U45798 (N_45798,N_43162,N_42394);
or U45799 (N_45799,N_42551,N_43479);
nor U45800 (N_45800,N_42736,N_43481);
and U45801 (N_45801,N_43499,N_42020);
nor U45802 (N_45802,N_43118,N_42460);
or U45803 (N_45803,N_43785,N_43166);
nor U45804 (N_45804,N_42011,N_42641);
nand U45805 (N_45805,N_42523,N_43490);
nor U45806 (N_45806,N_42631,N_43305);
and U45807 (N_45807,N_42938,N_43495);
nand U45808 (N_45808,N_43768,N_42600);
or U45809 (N_45809,N_42512,N_42528);
nand U45810 (N_45810,N_43054,N_43413);
xnor U45811 (N_45811,N_42660,N_43714);
or U45812 (N_45812,N_43581,N_42255);
nand U45813 (N_45813,N_42037,N_42158);
nor U45814 (N_45814,N_43176,N_43483);
nand U45815 (N_45815,N_42675,N_42492);
or U45816 (N_45816,N_43342,N_43277);
nand U45817 (N_45817,N_43194,N_43036);
nor U45818 (N_45818,N_42233,N_42120);
nor U45819 (N_45819,N_42982,N_42594);
and U45820 (N_45820,N_42402,N_42952);
xnor U45821 (N_45821,N_42290,N_42559);
or U45822 (N_45822,N_43795,N_43116);
nor U45823 (N_45823,N_42544,N_42350);
nor U45824 (N_45824,N_43063,N_42338);
or U45825 (N_45825,N_42202,N_42228);
and U45826 (N_45826,N_43145,N_42475);
and U45827 (N_45827,N_43287,N_43141);
or U45828 (N_45828,N_43941,N_42627);
nor U45829 (N_45829,N_43050,N_43340);
xnor U45830 (N_45830,N_42996,N_43457);
xnor U45831 (N_45831,N_43897,N_42152);
and U45832 (N_45832,N_43048,N_43788);
xor U45833 (N_45833,N_42542,N_43685);
and U45834 (N_45834,N_43351,N_43322);
nand U45835 (N_45835,N_43753,N_43438);
nor U45836 (N_45836,N_43282,N_43355);
nand U45837 (N_45837,N_43514,N_42766);
nor U45838 (N_45838,N_42282,N_42700);
nand U45839 (N_45839,N_43322,N_43817);
nor U45840 (N_45840,N_43418,N_43575);
xor U45841 (N_45841,N_42269,N_43980);
and U45842 (N_45842,N_43014,N_42572);
xor U45843 (N_45843,N_42332,N_42023);
nand U45844 (N_45844,N_43105,N_42135);
xnor U45845 (N_45845,N_42348,N_42509);
xnor U45846 (N_45846,N_43373,N_42343);
or U45847 (N_45847,N_42683,N_42388);
or U45848 (N_45848,N_42925,N_43115);
nor U45849 (N_45849,N_43263,N_42339);
xnor U45850 (N_45850,N_43096,N_42834);
xor U45851 (N_45851,N_43166,N_42220);
nor U45852 (N_45852,N_42988,N_42921);
xor U45853 (N_45853,N_42641,N_43128);
xor U45854 (N_45854,N_42720,N_43610);
or U45855 (N_45855,N_42415,N_43140);
nand U45856 (N_45856,N_43120,N_42207);
or U45857 (N_45857,N_42897,N_43710);
or U45858 (N_45858,N_43652,N_43581);
or U45859 (N_45859,N_43140,N_42503);
and U45860 (N_45860,N_43760,N_42235);
xnor U45861 (N_45861,N_43076,N_42830);
nand U45862 (N_45862,N_42181,N_42247);
or U45863 (N_45863,N_42972,N_42332);
xor U45864 (N_45864,N_42054,N_43419);
and U45865 (N_45865,N_43299,N_43541);
and U45866 (N_45866,N_42689,N_43910);
xnor U45867 (N_45867,N_42909,N_42593);
or U45868 (N_45868,N_42017,N_42985);
xnor U45869 (N_45869,N_42081,N_42819);
nand U45870 (N_45870,N_42637,N_43669);
nand U45871 (N_45871,N_42299,N_42394);
or U45872 (N_45872,N_43929,N_43856);
xnor U45873 (N_45873,N_42415,N_43963);
nand U45874 (N_45874,N_42267,N_42838);
nor U45875 (N_45875,N_42044,N_42406);
and U45876 (N_45876,N_42637,N_42266);
or U45877 (N_45877,N_43356,N_43968);
nand U45878 (N_45878,N_42596,N_42062);
and U45879 (N_45879,N_43554,N_42855);
nand U45880 (N_45880,N_43755,N_43143);
or U45881 (N_45881,N_43889,N_42269);
nand U45882 (N_45882,N_43497,N_42711);
or U45883 (N_45883,N_42797,N_42825);
and U45884 (N_45884,N_42237,N_43756);
and U45885 (N_45885,N_43321,N_42120);
xnor U45886 (N_45886,N_42293,N_43619);
nor U45887 (N_45887,N_43283,N_42405);
xor U45888 (N_45888,N_42221,N_42786);
and U45889 (N_45889,N_43213,N_43422);
nor U45890 (N_45890,N_43907,N_43803);
nand U45891 (N_45891,N_42848,N_43283);
xnor U45892 (N_45892,N_42453,N_43219);
or U45893 (N_45893,N_42590,N_42739);
nand U45894 (N_45894,N_43602,N_42275);
xnor U45895 (N_45895,N_42460,N_43629);
xnor U45896 (N_45896,N_42933,N_42052);
nor U45897 (N_45897,N_42678,N_42792);
nor U45898 (N_45898,N_43407,N_43134);
xor U45899 (N_45899,N_43573,N_42864);
xnor U45900 (N_45900,N_42262,N_43755);
or U45901 (N_45901,N_43085,N_43773);
or U45902 (N_45902,N_43786,N_42817);
or U45903 (N_45903,N_42820,N_43538);
nand U45904 (N_45904,N_43797,N_43568);
or U45905 (N_45905,N_43555,N_42104);
nand U45906 (N_45906,N_42134,N_43045);
or U45907 (N_45907,N_42428,N_42142);
nand U45908 (N_45908,N_43397,N_43465);
nor U45909 (N_45909,N_42329,N_43743);
and U45910 (N_45910,N_42934,N_43373);
or U45911 (N_45911,N_42295,N_42782);
and U45912 (N_45912,N_42854,N_42663);
nand U45913 (N_45913,N_42145,N_43472);
or U45914 (N_45914,N_42972,N_43149);
and U45915 (N_45915,N_42232,N_43447);
xnor U45916 (N_45916,N_43893,N_42631);
and U45917 (N_45917,N_43830,N_43699);
or U45918 (N_45918,N_43561,N_42055);
nand U45919 (N_45919,N_43428,N_43402);
nand U45920 (N_45920,N_42737,N_42631);
nand U45921 (N_45921,N_43809,N_42902);
xor U45922 (N_45922,N_42144,N_43534);
nand U45923 (N_45923,N_42784,N_43313);
or U45924 (N_45924,N_43668,N_43118);
and U45925 (N_45925,N_42917,N_43368);
and U45926 (N_45926,N_42704,N_42117);
and U45927 (N_45927,N_43416,N_42042);
xor U45928 (N_45928,N_42149,N_42650);
nand U45929 (N_45929,N_42914,N_42758);
xnor U45930 (N_45930,N_43370,N_42913);
nand U45931 (N_45931,N_42465,N_42800);
and U45932 (N_45932,N_43667,N_42399);
and U45933 (N_45933,N_42070,N_43717);
xnor U45934 (N_45934,N_43575,N_43025);
or U45935 (N_45935,N_42286,N_43286);
nand U45936 (N_45936,N_43310,N_42116);
and U45937 (N_45937,N_43217,N_42668);
and U45938 (N_45938,N_42004,N_43374);
xnor U45939 (N_45939,N_43551,N_42526);
xnor U45940 (N_45940,N_42389,N_42084);
nor U45941 (N_45941,N_42474,N_43667);
nor U45942 (N_45942,N_42034,N_43397);
nor U45943 (N_45943,N_42202,N_43553);
xor U45944 (N_45944,N_42582,N_42198);
and U45945 (N_45945,N_43380,N_43234);
nor U45946 (N_45946,N_43390,N_42327);
and U45947 (N_45947,N_42158,N_43251);
nand U45948 (N_45948,N_42071,N_42301);
nor U45949 (N_45949,N_43571,N_42618);
nand U45950 (N_45950,N_42246,N_42226);
and U45951 (N_45951,N_42019,N_42231);
nor U45952 (N_45952,N_42576,N_43457);
nor U45953 (N_45953,N_43525,N_43087);
and U45954 (N_45954,N_43676,N_43639);
or U45955 (N_45955,N_42863,N_42929);
nand U45956 (N_45956,N_43122,N_43579);
or U45957 (N_45957,N_43212,N_43083);
and U45958 (N_45958,N_42423,N_43989);
xnor U45959 (N_45959,N_42929,N_43998);
nor U45960 (N_45960,N_43021,N_42157);
or U45961 (N_45961,N_42330,N_43976);
nand U45962 (N_45962,N_43773,N_43562);
and U45963 (N_45963,N_42747,N_43890);
and U45964 (N_45964,N_42665,N_42909);
xnor U45965 (N_45965,N_42592,N_42971);
nor U45966 (N_45966,N_42807,N_43551);
nand U45967 (N_45967,N_42965,N_43703);
nor U45968 (N_45968,N_43018,N_42285);
and U45969 (N_45969,N_43455,N_42718);
nor U45970 (N_45970,N_42094,N_43673);
and U45971 (N_45971,N_43069,N_43431);
nand U45972 (N_45972,N_43749,N_42064);
nor U45973 (N_45973,N_43163,N_43664);
nand U45974 (N_45974,N_43011,N_43492);
or U45975 (N_45975,N_42315,N_43187);
and U45976 (N_45976,N_42858,N_42356);
and U45977 (N_45977,N_43902,N_42182);
or U45978 (N_45978,N_43909,N_43486);
or U45979 (N_45979,N_43208,N_42374);
and U45980 (N_45980,N_43723,N_43559);
nor U45981 (N_45981,N_43731,N_43452);
nand U45982 (N_45982,N_43232,N_43196);
or U45983 (N_45983,N_43138,N_43597);
nand U45984 (N_45984,N_43002,N_43597);
nor U45985 (N_45985,N_43528,N_42693);
xor U45986 (N_45986,N_43931,N_42737);
and U45987 (N_45987,N_43860,N_42863);
nand U45988 (N_45988,N_42455,N_42485);
nand U45989 (N_45989,N_42009,N_43992);
nor U45990 (N_45990,N_43082,N_42060);
or U45991 (N_45991,N_42040,N_43311);
and U45992 (N_45992,N_43268,N_42843);
or U45993 (N_45993,N_43180,N_42893);
nand U45994 (N_45994,N_42047,N_43571);
or U45995 (N_45995,N_43232,N_43298);
xnor U45996 (N_45996,N_42123,N_43576);
or U45997 (N_45997,N_43418,N_42892);
nand U45998 (N_45998,N_43033,N_43808);
and U45999 (N_45999,N_42024,N_43859);
xnor U46000 (N_46000,N_44946,N_45573);
and U46001 (N_46001,N_44428,N_44338);
or U46002 (N_46002,N_44918,N_44206);
or U46003 (N_46003,N_45729,N_45687);
and U46004 (N_46004,N_45000,N_44583);
nor U46005 (N_46005,N_45787,N_45739);
xor U46006 (N_46006,N_44689,N_44216);
and U46007 (N_46007,N_45992,N_45018);
or U46008 (N_46008,N_44587,N_44022);
nand U46009 (N_46009,N_44287,N_45988);
xnor U46010 (N_46010,N_44616,N_45067);
nor U46011 (N_46011,N_45124,N_45637);
nor U46012 (N_46012,N_44808,N_44292);
nand U46013 (N_46013,N_44248,N_45071);
and U46014 (N_46014,N_45888,N_45492);
or U46015 (N_46015,N_44602,N_45732);
or U46016 (N_46016,N_45140,N_44974);
or U46017 (N_46017,N_44351,N_44896);
and U46018 (N_46018,N_44840,N_45223);
nor U46019 (N_46019,N_44620,N_44515);
xnor U46020 (N_46020,N_45106,N_44607);
nand U46021 (N_46021,N_44357,N_45551);
xnor U46022 (N_46022,N_45785,N_44847);
nand U46023 (N_46023,N_45279,N_44824);
and U46024 (N_46024,N_44508,N_44105);
nor U46025 (N_46025,N_44766,N_45376);
xor U46026 (N_46026,N_45144,N_44276);
and U46027 (N_46027,N_44716,N_45002);
nor U46028 (N_46028,N_45201,N_44399);
nand U46029 (N_46029,N_45126,N_44679);
or U46030 (N_46030,N_44736,N_44113);
or U46031 (N_46031,N_44042,N_45504);
or U46032 (N_46032,N_44463,N_44036);
or U46033 (N_46033,N_45819,N_44321);
or U46034 (N_46034,N_45475,N_45967);
nor U46035 (N_46035,N_44584,N_44656);
or U46036 (N_46036,N_44640,N_45483);
and U46037 (N_46037,N_45565,N_44412);
nor U46038 (N_46038,N_44898,N_44062);
or U46039 (N_46039,N_45286,N_45911);
xor U46040 (N_46040,N_44245,N_45516);
xnor U46041 (N_46041,N_45069,N_45085);
and U46042 (N_46042,N_45287,N_45994);
xnor U46043 (N_46043,N_45448,N_44140);
or U46044 (N_46044,N_45354,N_44746);
xor U46045 (N_46045,N_45908,N_45547);
nand U46046 (N_46046,N_44127,N_44851);
and U46047 (N_46047,N_45629,N_44384);
nor U46048 (N_46048,N_45428,N_45304);
nand U46049 (N_46049,N_44010,N_44073);
or U46050 (N_46050,N_45865,N_45133);
xnor U46051 (N_46051,N_44516,N_45394);
nor U46052 (N_46052,N_45808,N_45505);
xor U46053 (N_46053,N_45156,N_45659);
or U46054 (N_46054,N_44241,N_44458);
xor U46055 (N_46055,N_44183,N_44492);
nand U46056 (N_46056,N_45767,N_45612);
and U46057 (N_46057,N_45571,N_44854);
nor U46058 (N_46058,N_45523,N_45939);
nand U46059 (N_46059,N_45555,N_45771);
and U46060 (N_46060,N_44398,N_44953);
or U46061 (N_46061,N_45519,N_44538);
nand U46062 (N_46062,N_44955,N_45609);
or U46063 (N_46063,N_45185,N_44517);
nor U46064 (N_46064,N_44718,N_45564);
xor U46065 (N_46065,N_44522,N_45957);
nand U46066 (N_46066,N_45820,N_45353);
nand U46067 (N_46067,N_44792,N_45092);
or U46068 (N_46068,N_44368,N_44800);
nor U46069 (N_46069,N_45860,N_45466);
nand U46070 (N_46070,N_44141,N_45081);
and U46071 (N_46071,N_44876,N_44580);
nand U46072 (N_46072,N_45363,N_44992);
nor U46073 (N_46073,N_45235,N_45530);
or U46074 (N_46074,N_44775,N_44197);
nand U46075 (N_46075,N_45907,N_45230);
and U46076 (N_46076,N_44260,N_45097);
xnor U46077 (N_46077,N_44919,N_45618);
or U46078 (N_46078,N_45675,N_45923);
and U46079 (N_46079,N_44664,N_44661);
and U46080 (N_46080,N_45434,N_45150);
nand U46081 (N_46081,N_45281,N_45242);
and U46082 (N_46082,N_44378,N_45259);
and U46083 (N_46083,N_45449,N_44281);
xor U46084 (N_46084,N_44817,N_45722);
xnor U46085 (N_46085,N_45545,N_45111);
xnor U46086 (N_46086,N_45674,N_44171);
nand U46087 (N_46087,N_44383,N_45415);
nor U46088 (N_46088,N_45750,N_45568);
or U46089 (N_46089,N_45958,N_44158);
xor U46090 (N_46090,N_45080,N_45747);
and U46091 (N_46091,N_44329,N_44560);
xor U46092 (N_46092,N_44026,N_44971);
nor U46093 (N_46093,N_45697,N_45973);
nor U46094 (N_46094,N_44174,N_45768);
or U46095 (N_46095,N_45815,N_45567);
nand U46096 (N_46096,N_45987,N_45333);
or U46097 (N_46097,N_44308,N_45758);
or U46098 (N_46098,N_44404,N_45636);
nand U46099 (N_46099,N_44966,N_45340);
nor U46100 (N_46100,N_45798,N_44456);
or U46101 (N_46101,N_44816,N_44262);
or U46102 (N_46102,N_45137,N_44848);
nor U46103 (N_46103,N_45847,N_44430);
nand U46104 (N_46104,N_45773,N_45754);
and U46105 (N_46105,N_44938,N_44674);
xor U46106 (N_46106,N_44393,N_44423);
nor U46107 (N_46107,N_44944,N_44299);
xor U46108 (N_46108,N_44549,N_45107);
nor U46109 (N_46109,N_44509,N_44998);
or U46110 (N_46110,N_45876,N_44787);
nor U46111 (N_46111,N_45859,N_45948);
nand U46112 (N_46112,N_44180,N_44985);
nand U46113 (N_46113,N_44785,N_44364);
nand U46114 (N_46114,N_44796,N_45592);
nand U46115 (N_46115,N_45816,N_44238);
and U46116 (N_46116,N_44909,N_44728);
xor U46117 (N_46117,N_45227,N_45460);
xnor U46118 (N_46118,N_44436,N_45195);
and U46119 (N_46119,N_44185,N_45702);
nand U46120 (N_46120,N_44879,N_45190);
nand U46121 (N_46121,N_45375,N_44625);
or U46122 (N_46122,N_44326,N_45465);
or U46123 (N_46123,N_45200,N_45942);
nand U46124 (N_46124,N_45009,N_45109);
nand U46125 (N_46125,N_44566,N_45469);
xor U46126 (N_46126,N_45061,N_45826);
or U46127 (N_46127,N_45797,N_44646);
and U46128 (N_46128,N_45209,N_45393);
nor U46129 (N_46129,N_45057,N_45828);
nor U46130 (N_46130,N_44480,N_45639);
and U46131 (N_46131,N_45944,N_45507);
nor U46132 (N_46132,N_44426,N_44878);
nor U46133 (N_46133,N_45409,N_45361);
nand U46134 (N_46134,N_44934,N_44561);
or U46135 (N_46135,N_44343,N_45709);
and U46136 (N_46136,N_44818,N_44341);
nand U46137 (N_46137,N_45053,N_44781);
and U46138 (N_46138,N_44272,N_45197);
nor U46139 (N_46139,N_45662,N_45162);
and U46140 (N_46140,N_44608,N_44937);
xor U46141 (N_46141,N_45803,N_44478);
nor U46142 (N_46142,N_44332,N_45924);
or U46143 (N_46143,N_44350,N_45717);
and U46144 (N_46144,N_44900,N_45093);
nand U46145 (N_46145,N_44941,N_45897);
nand U46146 (N_46146,N_45921,N_44410);
nor U46147 (N_46147,N_45779,N_44578);
xnor U46148 (N_46148,N_44672,N_44565);
or U46149 (N_46149,N_44479,N_44903);
and U46150 (N_46150,N_44634,N_45682);
or U46151 (N_46151,N_44089,N_44988);
nand U46152 (N_46152,N_44852,N_45514);
nor U46153 (N_46153,N_45213,N_45003);
nand U46154 (N_46154,N_45496,N_44451);
xnor U46155 (N_46155,N_45270,N_45313);
and U46156 (N_46156,N_44550,N_44576);
and U46157 (N_46157,N_45892,N_44837);
and U46158 (N_46158,N_44211,N_44239);
or U46159 (N_46159,N_44474,N_44846);
nor U46160 (N_46160,N_45367,N_45362);
or U46161 (N_46161,N_44629,N_44845);
and U46162 (N_46162,N_44986,N_45290);
xnor U46163 (N_46163,N_44473,N_45142);
nand U46164 (N_46164,N_45622,N_44527);
or U46165 (N_46165,N_44790,N_44496);
xor U46166 (N_46166,N_44717,N_44791);
nand U46167 (N_46167,N_45688,N_45045);
nand U46168 (N_46168,N_44405,N_44635);
or U46169 (N_46169,N_44553,N_44370);
xor U46170 (N_46170,N_44149,N_45341);
xnor U46171 (N_46171,N_44096,N_45438);
nand U46172 (N_46172,N_44546,N_45116);
or U46173 (N_46173,N_45904,N_44659);
nor U46174 (N_46174,N_45872,N_44881);
and U46175 (N_46175,N_44415,N_44493);
or U46176 (N_46176,N_44855,N_44588);
or U46177 (N_46177,N_44614,N_44555);
nand U46178 (N_46178,N_44932,N_44631);
or U46179 (N_46179,N_44325,N_45595);
and U46180 (N_46180,N_44853,N_44313);
xnor U46181 (N_46181,N_45184,N_44075);
xnor U46182 (N_46182,N_44880,N_45342);
xor U46183 (N_46183,N_45205,N_44653);
and U46184 (N_46184,N_45015,N_44155);
and U46185 (N_46185,N_45864,N_44088);
nor U46186 (N_46186,N_44673,N_44598);
nand U46187 (N_46187,N_45099,N_45079);
nand U46188 (N_46188,N_44891,N_44641);
nand U46189 (N_46189,N_44314,N_45463);
or U46190 (N_46190,N_44406,N_45539);
nand U46191 (N_46191,N_44340,N_44890);
nor U46192 (N_46192,N_44109,N_45563);
nand U46193 (N_46193,N_44452,N_45578);
xnor U46194 (N_46194,N_44825,N_44031);
xnor U46195 (N_46195,N_45305,N_44693);
xnor U46196 (N_46196,N_44166,N_44633);
and U46197 (N_46197,N_45764,N_44823);
nor U46198 (N_46198,N_44860,N_45701);
xnor U46199 (N_46199,N_44161,N_45405);
nor U46200 (N_46200,N_45384,N_45078);
or U46201 (N_46201,N_45387,N_45010);
nand U46202 (N_46202,N_44121,N_45154);
and U46203 (N_46203,N_45218,N_44004);
and U46204 (N_46204,N_45168,N_45536);
or U46205 (N_46205,N_44250,N_44061);
xor U46206 (N_46206,N_44135,N_45733);
nand U46207 (N_46207,N_45382,N_45268);
and U46208 (N_46208,N_44793,N_44665);
nand U46209 (N_46209,N_44472,N_45901);
and U46210 (N_46210,N_44571,N_45303);
nor U46211 (N_46211,N_44084,N_45765);
nand U46212 (N_46212,N_44295,N_45147);
and U46213 (N_46213,N_44815,N_45026);
nand U46214 (N_46214,N_44839,N_44297);
nand U46215 (N_46215,N_44142,N_45331);
xor U46216 (N_46216,N_45343,N_45174);
nand U46217 (N_46217,N_45856,N_45143);
nand U46218 (N_46218,N_45931,N_44687);
nor U46219 (N_46219,N_45572,N_45373);
and U46220 (N_46220,N_45456,N_45068);
nor U46221 (N_46221,N_45446,N_45721);
nor U46222 (N_46222,N_44386,N_45339);
nor U46223 (N_46223,N_44371,N_44290);
or U46224 (N_46224,N_44895,N_44417);
nor U46225 (N_46225,N_45755,N_44117);
nor U46226 (N_46226,N_45678,N_45014);
nand U46227 (N_46227,N_44301,N_45048);
nor U46228 (N_46228,N_45544,N_45976);
or U46229 (N_46229,N_44735,N_44585);
nand U46230 (N_46230,N_44726,N_44702);
nor U46231 (N_46231,N_45207,N_44365);
or U46232 (N_46232,N_44367,N_45730);
xnor U46233 (N_46233,N_44320,N_44048);
nor U46234 (N_46234,N_45294,N_45800);
nand U46235 (N_46235,N_44432,N_45677);
and U46236 (N_46236,N_44756,N_45600);
nand U46237 (N_46237,N_45685,N_44226);
xor U46238 (N_46238,N_45635,N_45710);
or U46239 (N_46239,N_44168,N_44810);
xnor U46240 (N_46240,N_45704,N_45882);
and U46241 (N_46241,N_44202,N_45051);
or U46242 (N_46242,N_45262,N_45017);
xor U46243 (N_46243,N_44025,N_45982);
nor U46244 (N_46244,N_44794,N_44685);
or U46245 (N_46245,N_44425,N_45113);
xor U46246 (N_46246,N_44220,N_44738);
nand U46247 (N_46247,N_44867,N_44795);
xnor U46248 (N_46248,N_45086,N_45176);
or U46249 (N_46249,N_45309,N_45711);
or U46250 (N_46250,N_45756,N_44044);
nor U46251 (N_46251,N_45273,N_45953);
nor U46252 (N_46252,N_44092,N_45358);
or U46253 (N_46253,N_45866,N_45699);
and U46254 (N_46254,N_45408,N_44982);
xnor U46255 (N_46255,N_45810,N_45254);
and U46256 (N_46256,N_44058,N_44445);
nor U46257 (N_46257,N_44481,N_45625);
xnor U46258 (N_46258,N_45788,N_44275);
xnor U46259 (N_46259,N_45941,N_44139);
nand U46260 (N_46260,N_45412,N_45100);
nor U46261 (N_46261,N_45591,N_45245);
or U46262 (N_46262,N_44129,N_44060);
nand U46263 (N_46263,N_45736,N_44501);
nor U46264 (N_46264,N_44812,N_44242);
nor U46265 (N_46265,N_45135,N_44112);
nand U46266 (N_46266,N_44041,N_44352);
and U46267 (N_46267,N_45666,N_45321);
nand U46268 (N_46268,N_44051,N_44028);
and U46269 (N_46269,N_45902,N_45575);
nand U46270 (N_46270,N_45115,N_45265);
and U46271 (N_46271,N_45216,N_44596);
or U46272 (N_46272,N_45500,N_45984);
and U46273 (N_46273,N_44768,N_45593);
nor U46274 (N_46274,N_44045,N_45929);
nor U46275 (N_46275,N_45224,N_45282);
and U46276 (N_46276,N_44539,N_44310);
or U46277 (N_46277,N_45577,N_44594);
xnor U46278 (N_46278,N_44654,N_45590);
or U46279 (N_46279,N_45997,N_44874);
nand U46280 (N_46280,N_44579,N_45686);
and U46281 (N_46281,N_45665,N_45096);
nand U46282 (N_46282,N_44940,N_45933);
nor U46283 (N_46283,N_44122,N_45183);
nor U46284 (N_46284,N_44151,N_44957);
or U46285 (N_46285,N_45647,N_45851);
nand U46286 (N_46286,N_45608,N_45926);
xor U46287 (N_46287,N_45813,N_44928);
or U46288 (N_46288,N_44315,N_44021);
nor U46289 (N_46289,N_45420,N_45878);
nor U46290 (N_46290,N_44069,N_45762);
or U46291 (N_46291,N_45237,N_44134);
nor U46292 (N_46292,N_45966,N_45356);
xnor U46293 (N_46293,N_45980,N_44385);
nor U46294 (N_46294,N_45292,N_44111);
nor U46295 (N_46295,N_45127,N_44462);
or U46296 (N_46296,N_44963,N_44873);
and U46297 (N_46297,N_45936,N_44930);
nand U46298 (N_46298,N_45386,N_45171);
nor U46299 (N_46299,N_45199,N_45658);
and U46300 (N_46300,N_44869,N_45350);
nor U46301 (N_46301,N_44783,N_44468);
and U46302 (N_46302,N_45841,N_44666);
and U46303 (N_46303,N_45244,N_44413);
nor U46304 (N_46304,N_45794,N_45410);
xor U46305 (N_46305,N_44434,N_44083);
nand U46306 (N_46306,N_44628,N_45239);
or U46307 (N_46307,N_45617,N_45377);
nand U46308 (N_46308,N_45480,N_45403);
nand U46309 (N_46309,N_44347,N_44150);
nor U46310 (N_46310,N_45570,N_45352);
and U46311 (N_46311,N_45164,N_45473);
or U46312 (N_46312,N_45510,N_45975);
or U46313 (N_46313,N_44017,N_44369);
xor U46314 (N_46314,N_45916,N_45034);
nand U46315 (N_46315,N_45013,N_44005);
xnor U46316 (N_46316,N_45186,N_45046);
or U46317 (N_46317,N_44914,N_44229);
or U46318 (N_46318,N_44175,N_44771);
or U46319 (N_46319,N_45249,N_45182);
nand U46320 (N_46320,N_44905,N_44249);
xnor U46321 (N_46321,N_45493,N_45338);
xor U46322 (N_46322,N_45024,N_45839);
nor U46323 (N_46323,N_45430,N_44006);
xor U46324 (N_46324,N_44188,N_45712);
or U46325 (N_46325,N_45596,N_45757);
xnor U46326 (N_46326,N_44801,N_44520);
and U46327 (N_46327,N_45495,N_44186);
xor U46328 (N_46328,N_45760,N_45920);
xor U46329 (N_46329,N_45349,N_44231);
nand U46330 (N_46330,N_44870,N_45720);
or U46331 (N_46331,N_45324,N_44037);
nor U46332 (N_46332,N_44376,N_44849);
nor U46333 (N_46333,N_45491,N_44683);
and U46334 (N_46334,N_45807,N_45020);
xor U46335 (N_46335,N_44038,N_45646);
or U46336 (N_46336,N_44304,N_44573);
or U46337 (N_46337,N_44605,N_44176);
and U46338 (N_46338,N_44729,N_44564);
xnor U46339 (N_46339,N_45474,N_45940);
xor U46340 (N_46340,N_44850,N_45970);
nand U46341 (N_46341,N_45744,N_45044);
and U46342 (N_46342,N_44001,N_45334);
nand U46343 (N_46343,N_44471,N_45642);
xor U46344 (N_46344,N_44780,N_44951);
nand U46345 (N_46345,N_45795,N_45588);
and U46346 (N_46346,N_44532,N_44972);
nor U46347 (N_46347,N_44644,N_44433);
nand U46348 (N_46348,N_44563,N_44733);
and U46349 (N_46349,N_45753,N_44234);
nor U46350 (N_46350,N_45777,N_45319);
nor U46351 (N_46351,N_44582,N_45241);
and U46352 (N_46352,N_44671,N_45643);
nand U46353 (N_46353,N_44429,N_44328);
or U46354 (N_46354,N_44612,N_45512);
nor U46355 (N_46355,N_45713,N_45553);
nor U46356 (N_46356,N_45977,N_44007);
or U46357 (N_46357,N_45731,N_45909);
xnor U46358 (N_46358,N_45995,N_44136);
xor U46359 (N_46359,N_44411,N_44894);
xnor U46360 (N_46360,N_44125,N_45243);
nor U46361 (N_46361,N_45478,N_44630);
xor U46362 (N_46362,N_45968,N_45439);
and U46363 (N_46363,N_44146,N_44306);
or U46364 (N_46364,N_44543,N_44029);
nand U46365 (N_46365,N_44106,N_44396);
nand U46366 (N_46366,N_45132,N_44259);
xnor U46367 (N_46367,N_44487,N_45814);
nor U46368 (N_46368,N_45613,N_44513);
xor U46369 (N_46369,N_44252,N_45895);
nor U46370 (N_46370,N_45255,N_45293);
or U46371 (N_46371,N_45032,N_44018);
xnor U46372 (N_46372,N_44567,N_45834);
xor U46373 (N_46373,N_45741,N_45885);
and U46374 (N_46374,N_44877,N_44609);
and U46375 (N_46375,N_44266,N_45670);
and U46376 (N_46376,N_44907,N_44160);
xnor U46377 (N_46377,N_45634,N_45260);
and U46378 (N_46378,N_44862,N_44901);
xor U46379 (N_46379,N_44777,N_45138);
xnor U46380 (N_46380,N_45442,N_45891);
or U46381 (N_46381,N_44484,N_45311);
nor U46382 (N_46382,N_44642,N_45318);
nand U46383 (N_46383,N_45153,N_44556);
or U46384 (N_46384,N_45915,N_45027);
nand U46385 (N_46385,N_44558,N_44236);
nand U46386 (N_46386,N_45327,N_45212);
nor U46387 (N_46387,N_44931,N_45307);
nand U46388 (N_46388,N_45535,N_44032);
xor U46389 (N_46389,N_44143,N_45627);
and U46390 (N_46390,N_44819,N_45922);
xnor U46391 (N_46391,N_45468,N_45030);
or U46392 (N_46392,N_44568,N_45886);
xor U46393 (N_46393,N_44622,N_44030);
and U46394 (N_46394,N_45599,N_44443);
or U46395 (N_46395,N_44882,N_45167);
nand U46396 (N_46396,N_44649,N_45188);
nor U46397 (N_46397,N_45910,N_45837);
or U46398 (N_46398,N_45210,N_44660);
or U46399 (N_46399,N_45157,N_44886);
and U46400 (N_46400,N_44130,N_44066);
xor U46401 (N_46401,N_44043,N_45831);
and U46402 (N_46402,N_45679,N_44745);
or U46403 (N_46403,N_44589,N_44958);
or U46404 (N_46404,N_45052,N_44913);
and U46405 (N_46405,N_44495,N_45652);
or U46406 (N_46406,N_45776,N_44137);
nor U46407 (N_46407,N_44518,N_45169);
nand U46408 (N_46408,N_44271,N_44834);
xnor U46409 (N_46409,N_44779,N_45371);
and U46410 (N_46410,N_45894,N_44912);
nor U46411 (N_46411,N_45369,N_45951);
or U46412 (N_46412,N_45518,N_45073);
and U46413 (N_46413,N_45134,N_44696);
nor U46414 (N_46414,N_44805,N_45914);
nand U46415 (N_46415,N_45511,N_44826);
and U46416 (N_46416,N_44773,N_45850);
or U46417 (N_46417,N_44163,N_45074);
xor U46418 (N_46418,N_44449,N_44720);
nand U46419 (N_46419,N_45288,N_44739);
xor U46420 (N_46420,N_44713,N_45938);
nand U46421 (N_46421,N_45125,N_45986);
nand U46422 (N_46422,N_45784,N_44214);
or U46423 (N_46423,N_45348,N_44521);
nor U46424 (N_46424,N_45484,N_44939);
nor U46425 (N_46425,N_44500,N_45005);
or U46426 (N_46426,N_44806,N_44540);
xnor U46427 (N_46427,N_44157,N_44514);
nor U46428 (N_46428,N_44994,N_44755);
or U46429 (N_46429,N_45253,N_45330);
or U46430 (N_46430,N_45738,N_44270);
nand U46431 (N_46431,N_44204,N_45094);
or U46432 (N_46432,N_45857,N_44668);
nand U46433 (N_46433,N_45566,N_44942);
and U46434 (N_46434,N_45221,N_44014);
nor U46435 (N_46435,N_45487,N_45846);
or U46436 (N_46436,N_45214,N_45783);
or U46437 (N_46437,N_44593,N_44722);
nor U46438 (N_46438,N_44191,N_44688);
and U46439 (N_46439,N_44759,N_44925);
or U46440 (N_46440,N_45441,N_45335);
nand U46441 (N_46441,N_45192,N_45683);
and U46442 (N_46442,N_44747,N_45267);
nand U46443 (N_46443,N_45606,N_44537);
nor U46444 (N_46444,N_45715,N_45737);
or U46445 (N_46445,N_44483,N_45998);
nor U46446 (N_46446,N_44694,N_44068);
xnor U46447 (N_46447,N_45039,N_44858);
or U46448 (N_46448,N_44770,N_45752);
xnor U46449 (N_46449,N_45781,N_44557);
nor U46450 (N_46450,N_45574,N_44335);
xor U46451 (N_46451,N_45694,N_45641);
nor U46452 (N_46452,N_45378,N_44316);
or U46453 (N_46453,N_44647,N_44488);
or U46454 (N_46454,N_45440,N_45996);
or U46455 (N_46455,N_45896,N_44402);
or U46456 (N_46456,N_45211,N_44435);
nor U46457 (N_46457,N_44305,N_45619);
xnor U46458 (N_46458,N_44504,N_45047);
xnor U46459 (N_46459,N_45962,N_44650);
and U46460 (N_46460,N_44119,N_45978);
xnor U46461 (N_46461,N_45379,N_45041);
nand U46462 (N_46462,N_44945,N_44662);
or U46463 (N_46463,N_44677,N_44570);
or U46464 (N_46464,N_44167,N_44727);
and U46465 (N_46465,N_45277,N_45433);
or U46466 (N_46466,N_45170,N_44243);
or U46467 (N_46467,N_44450,N_44969);
and U46468 (N_46468,N_44764,N_44948);
and U46469 (N_46469,N_45871,N_44172);
or U46470 (N_46470,N_45424,N_44381);
or U46471 (N_46471,N_45389,N_45672);
and U46472 (N_46472,N_44120,N_44349);
and U46473 (N_46473,N_45422,N_44389);
nand U46474 (N_46474,N_44192,N_45064);
and U46475 (N_46475,N_45453,N_44392);
and U46476 (N_46476,N_45118,N_44279);
or U46477 (N_46477,N_44623,N_45299);
nor U46478 (N_46478,N_44822,N_45222);
and U46479 (N_46479,N_45825,N_44908);
xnor U46480 (N_46480,N_44959,N_44064);
and U46481 (N_46481,N_45040,N_45822);
or U46482 (N_46482,N_44431,N_45918);
nor U46483 (N_46483,N_45950,N_44205);
or U46484 (N_46484,N_45528,N_44933);
nand U46485 (N_46485,N_44523,N_44170);
xor U46486 (N_46486,N_45421,N_44104);
nand U46487 (N_46487,N_45368,N_44379);
xor U46488 (N_46488,N_44973,N_44189);
nand U46489 (N_46489,N_45217,N_44547);
xnor U46490 (N_46490,N_44758,N_44078);
xnor U46491 (N_46491,N_45661,N_45947);
and U46492 (N_46492,N_45129,N_45793);
and U46493 (N_46493,N_45202,N_44701);
and U46494 (N_46494,N_45189,N_45275);
xor U46495 (N_46495,N_44144,N_44789);
nor U46496 (N_46496,N_45228,N_45700);
xor U46497 (N_46497,N_44511,N_45809);
nand U46498 (N_46498,N_44725,N_44485);
and U46499 (N_46499,N_45937,N_45559);
nand U46500 (N_46500,N_44678,N_45435);
xnor U46501 (N_46501,N_45411,N_45072);
and U46502 (N_46502,N_45862,N_45043);
xnor U46503 (N_46503,N_44228,N_45136);
or U46504 (N_46504,N_44618,N_44444);
or U46505 (N_46505,N_44591,N_45443);
nand U46506 (N_46506,N_44173,N_44981);
xor U46507 (N_46507,N_44154,N_44600);
nor U46508 (N_46508,N_44915,N_45139);
and U46509 (N_46509,N_44437,N_45796);
nor U46510 (N_46510,N_45471,N_45925);
and U46511 (N_46511,N_44871,N_45062);
or U46512 (N_46512,N_45959,N_45905);
nand U46513 (N_46513,N_44505,N_45402);
xnor U46514 (N_46514,N_44264,N_45927);
and U46515 (N_46515,N_45522,N_44535);
nand U46516 (N_46516,N_44606,N_45821);
xnor U46517 (N_46517,N_45160,N_44544);
nor U46518 (N_46518,N_44207,N_45488);
or U46519 (N_46519,N_44237,N_45684);
nand U46520 (N_46520,N_44541,N_44980);
xnor U46521 (N_46521,N_44804,N_45623);
xor U46522 (N_46522,N_44681,N_45280);
nand U46523 (N_46523,N_45316,N_45166);
nor U46524 (N_46524,N_45397,N_45749);
xor U46525 (N_46525,N_45499,N_45001);
or U46526 (N_46526,N_45123,N_44712);
and U46527 (N_46527,N_44960,N_44454);
nor U46528 (N_46528,N_44637,N_44531);
or U46529 (N_46529,N_45858,N_44507);
nor U46530 (N_46530,N_44813,N_45705);
nand U46531 (N_46531,N_44708,N_44447);
xnor U46532 (N_46532,N_45102,N_45965);
nand U46533 (N_46533,N_45250,N_44082);
nand U46534 (N_46534,N_45130,N_45734);
and U46535 (N_46535,N_44752,N_45095);
and U46536 (N_46536,N_45019,N_45594);
and U46537 (N_46537,N_45525,N_45893);
or U46538 (N_46538,N_44698,N_44979);
nor U46539 (N_46539,N_45532,N_45314);
nor U46540 (N_46540,N_45240,N_45742);
nor U46541 (N_46541,N_44838,N_45289);
or U46542 (N_46542,N_44265,N_45695);
nand U46543 (N_46543,N_45543,N_44285);
nor U46544 (N_46544,N_44181,N_44461);
xor U46545 (N_46545,N_45521,N_44296);
or U46546 (N_46546,N_44274,N_44224);
and U46547 (N_46547,N_44107,N_45817);
xor U46548 (N_46548,N_45101,N_44990);
and U46549 (N_46549,N_44706,N_44273);
nand U46550 (N_46550,N_44528,N_44097);
xnor U46551 (N_46551,N_44311,N_45383);
nand U46552 (N_46552,N_45954,N_45301);
nor U46553 (N_46553,N_45601,N_44569);
nand U46554 (N_46554,N_44697,N_44828);
and U46555 (N_46555,N_45725,N_45119);
and U46556 (N_46556,N_45935,N_44318);
or U46557 (N_46557,N_45236,N_45829);
xnor U46558 (N_46558,N_45297,N_44344);
nor U46559 (N_46559,N_45981,N_45066);
and U46560 (N_46560,N_45991,N_45450);
nor U46561 (N_46561,N_45486,N_44529);
xnor U46562 (N_46562,N_45506,N_44949);
and U46563 (N_46563,N_44603,N_44639);
or U46564 (N_46564,N_44519,N_44247);
xnor U46565 (N_46565,N_45006,N_44235);
or U46566 (N_46566,N_44682,N_44750);
xnor U46567 (N_46567,N_44178,N_44184);
nand U46568 (N_46568,N_44977,N_44502);
xor U46569 (N_46569,N_44498,N_45698);
nand U46570 (N_46570,N_45597,N_45323);
xor U46571 (N_46571,N_45903,N_44741);
nand U46572 (N_46572,N_45252,N_45204);
xor U46573 (N_46573,N_44095,N_44049);
xnor U46574 (N_46574,N_44162,N_45630);
nand U46575 (N_46575,N_44291,N_44391);
or U46576 (N_46576,N_44684,N_44407);
and U46577 (N_46577,N_45537,N_45302);
nand U46578 (N_46578,N_44020,N_45861);
nand U46579 (N_46579,N_44744,N_44841);
or U46580 (N_46580,N_45558,N_44888);
or U46581 (N_46581,N_44740,N_45481);
xor U46582 (N_46582,N_44293,N_44551);
and U46583 (N_46583,N_44926,N_45110);
xnor U46584 (N_46584,N_45426,N_44289);
nand U46585 (N_46585,N_45763,N_44968);
nor U46586 (N_46586,N_44667,N_45663);
xor U46587 (N_46587,N_45569,N_45088);
or U46588 (N_46588,N_44268,N_44455);
xnor U46589 (N_46589,N_45880,N_45624);
nand U46590 (N_46590,N_45727,N_44597);
nor U46591 (N_46591,N_45502,N_45489);
and U46592 (N_46592,N_45317,N_45952);
nor U46593 (N_46593,N_45413,N_44169);
nor U46594 (N_46594,N_44778,N_45120);
nor U46595 (N_46595,N_45759,N_44053);
or U46596 (N_46596,N_45431,N_44464);
and U46597 (N_46597,N_45638,N_44730);
or U46598 (N_46598,N_44772,N_45964);
and U46599 (N_46599,N_45900,N_44892);
nand U46600 (N_46600,N_45655,N_45883);
nor U46601 (N_46601,N_45983,N_44947);
and U46602 (N_46602,N_45141,N_44586);
and U46603 (N_46603,N_44387,N_45726);
xor U46604 (N_46604,N_44924,N_45065);
and U46605 (N_46605,N_45653,N_44643);
and U46606 (N_46606,N_44193,N_45989);
xnor U46607 (N_46607,N_45640,N_44194);
or U46608 (N_46608,N_45075,N_45312);
nand U46609 (N_46609,N_45370,N_44574);
and U46610 (N_46610,N_44156,N_44989);
or U46611 (N_46611,N_45503,N_44427);
and U46612 (N_46612,N_45208,N_45560);
xor U46613 (N_46613,N_44382,N_45960);
nand U46614 (N_46614,N_44476,N_44148);
xnor U46615 (N_46615,N_44615,N_45836);
and U46616 (N_46616,N_44309,N_45761);
nand U46617 (N_46617,N_44337,N_45668);
nor U46618 (N_46618,N_44669,N_45056);
and U46619 (N_46619,N_44754,N_45789);
xor U46620 (N_46620,N_44534,N_45689);
and U46621 (N_46621,N_44590,N_44027);
and U46622 (N_46622,N_44927,N_44999);
nor U46623 (N_46623,N_45283,N_44145);
or U46624 (N_46624,N_45346,N_45451);
or U46625 (N_46625,N_45692,N_45219);
xnor U46626 (N_46626,N_44658,N_44330);
or U46627 (N_46627,N_45644,N_44916);
and U46628 (N_46628,N_44645,N_44763);
and U46629 (N_46629,N_44562,N_44284);
nand U46630 (N_46630,N_45278,N_44835);
and U46631 (N_46631,N_44008,N_45416);
and U46632 (N_46632,N_44056,N_45517);
or U46633 (N_46633,N_45586,N_45971);
nor U46634 (N_46634,N_44533,N_45028);
nor U46635 (N_46635,N_44497,N_44814);
xor U46636 (N_46636,N_44035,N_44422);
and U46637 (N_46637,N_44700,N_44294);
nand U46638 (N_46638,N_44355,N_44525);
and U46639 (N_46639,N_45091,N_44278);
nand U46640 (N_46640,N_44012,N_44221);
nor U46641 (N_46641,N_45868,N_44374);
nand U46642 (N_46642,N_45117,N_45146);
nand U46643 (N_46643,N_44039,N_44288);
nor U46644 (N_46644,N_45562,N_45472);
nand U46645 (N_46645,N_45775,N_44680);
xnor U46646 (N_46646,N_44737,N_44530);
xor U46647 (N_46647,N_45181,N_44690);
nor U46648 (N_46648,N_45054,N_45552);
and U46649 (N_46649,N_44961,N_45614);
nor U46650 (N_46650,N_44240,N_45844);
xnor U46651 (N_46651,N_44705,N_45520);
or U46652 (N_46652,N_44510,N_45291);
nor U46653 (N_46653,N_44448,N_44910);
and U46654 (N_46654,N_45226,N_44993);
nand U46655 (N_46655,N_44124,N_44359);
and U46656 (N_46656,N_45231,N_45791);
and U46657 (N_46657,N_45012,N_45112);
and U46658 (N_46658,N_44453,N_44843);
or U46659 (N_46659,N_44071,N_45380);
nand U46660 (N_46660,N_45329,N_45746);
nand U46661 (N_46661,N_44719,N_45031);
xnor U46662 (N_46662,N_45890,N_45234);
nor U46663 (N_46663,N_45158,N_45248);
nand U46664 (N_46664,N_45229,N_44377);
or U46665 (N_46665,N_45664,N_44552);
and U46666 (N_46666,N_45529,N_44128);
or U46667 (N_46667,N_44195,N_44346);
nand U46668 (N_46668,N_44223,N_45145);
or U46669 (N_46669,N_44280,N_44929);
or U46670 (N_46670,N_45276,N_44198);
or U46671 (N_46671,N_44131,N_44003);
nor U46672 (N_46672,N_44177,N_45203);
and U46673 (N_46673,N_44094,N_45187);
nor U46674 (N_46674,N_44187,N_44592);
nand U46675 (N_46675,N_45628,N_45285);
or U46676 (N_46676,N_44863,N_44984);
nor U46677 (N_46677,N_45385,N_45611);
and U46678 (N_46678,N_44132,N_45059);
and U46679 (N_46679,N_45633,N_45527);
nor U46680 (N_46680,N_45840,N_44554);
xor U46681 (N_46681,N_44657,N_45999);
xnor U46682 (N_46682,N_45812,N_45554);
and U46683 (N_46683,N_44408,N_45853);
xnor U46684 (N_46684,N_45108,N_45546);
and U46685 (N_46685,N_45930,N_44967);
or U46686 (N_46686,N_45152,N_44324);
xnor U46687 (N_46687,N_45598,N_45357);
xor U46688 (N_46688,N_44126,N_45549);
and U46689 (N_46689,N_44821,N_45246);
xor U46690 (N_46690,N_44506,N_44074);
nor U46691 (N_46691,N_44477,N_44286);
and U46692 (N_46692,N_45206,N_45557);
or U46693 (N_46693,N_45306,N_44710);
nor U46694 (N_46694,N_45427,N_44334);
and U46695 (N_46695,N_45025,N_45476);
nor U46696 (N_46696,N_44317,N_44965);
xor U46697 (N_46697,N_45906,N_45770);
and U46698 (N_46698,N_44100,N_45513);
xor U46699 (N_46699,N_44651,N_44753);
nor U46700 (N_46700,N_44373,N_45610);
xor U46701 (N_46701,N_45708,N_45121);
xnor U46702 (N_46702,N_44906,N_45786);
and U46703 (N_46703,N_44152,N_44923);
nand U46704 (N_46704,N_44442,N_44219);
and U46705 (N_46705,N_45723,N_44889);
nor U46706 (N_46706,N_44695,N_45155);
and U46707 (N_46707,N_44486,N_45220);
xnor U46708 (N_46708,N_44872,N_45508);
or U46709 (N_46709,N_44638,N_45974);
nand U46710 (N_46710,N_44624,N_44784);
nor U46711 (N_46711,N_44232,N_44063);
nand U46712 (N_46712,N_45359,N_45580);
nand U46713 (N_46713,N_45718,N_45772);
nor U46714 (N_46714,N_44034,N_44209);
and U46715 (N_46715,N_45748,N_45148);
xor U46716 (N_46716,N_45407,N_45042);
or U46717 (N_46717,N_44251,N_45414);
nand U46718 (N_46718,N_44950,N_45404);
or U46719 (N_46719,N_45912,N_44077);
xnor U46720 (N_46720,N_45849,N_44200);
or U46721 (N_46721,N_44619,N_45029);
or U46722 (N_46722,N_45194,N_44358);
nor U46723 (N_46723,N_45023,N_44190);
or U46724 (N_46724,N_44499,N_44460);
nand U46725 (N_46725,N_45780,N_45485);
xnor U46726 (N_46726,N_45366,N_44256);
nor U46727 (N_46727,N_44081,N_45792);
and U46728 (N_46728,N_45833,N_44099);
xor U46729 (N_46729,N_44976,N_44116);
nand U46730 (N_46730,N_44323,N_45706);
and U46731 (N_46731,N_44090,N_44997);
nor U46732 (N_46732,N_44648,N_44830);
xnor U46733 (N_46733,N_44675,N_45855);
nor U46734 (N_46734,N_44482,N_45541);
nand U46735 (N_46735,N_44842,N_44512);
nor U46736 (N_46736,N_45175,N_45300);
xor U46737 (N_46737,N_44611,N_45782);
nor U46738 (N_46738,N_44093,N_44617);
nor U46739 (N_46739,N_45298,N_44199);
nand U46740 (N_46740,N_44345,N_44621);
and U46741 (N_46741,N_44857,N_44595);
and U46742 (N_46742,N_44962,N_44749);
nor U46743 (N_46743,N_45870,N_45272);
nand U46744 (N_46744,N_44331,N_44401);
xnor U46745 (N_46745,N_44388,N_44394);
nor U46746 (N_46746,N_45161,N_45256);
xnor U46747 (N_46747,N_45806,N_44255);
and U46748 (N_46748,N_44743,N_44788);
or U46749 (N_46749,N_44055,N_44098);
nor U46750 (N_46750,N_44864,N_44164);
nand U46751 (N_46751,N_45919,N_44964);
or U46752 (N_46752,N_44802,N_45524);
xnor U46753 (N_46753,N_44277,N_44459);
xnor U46754 (N_46754,N_44230,N_45585);
xor U46755 (N_46755,N_44859,N_45667);
xnor U46756 (N_46756,N_44298,N_45751);
xnor U46757 (N_46757,N_45049,N_45271);
xor U46758 (N_46758,N_45322,N_45645);
and U46759 (N_46759,N_45258,N_45284);
xor U46760 (N_46760,N_45607,N_44936);
and U46761 (N_46761,N_45461,N_44921);
or U46762 (N_46762,N_45452,N_45945);
xor U46763 (N_46763,N_44983,N_44312);
xor U46764 (N_46764,N_44715,N_44632);
nand U46765 (N_46765,N_45766,N_44087);
nand U46766 (N_46766,N_45036,N_44467);
xnor U46767 (N_46767,N_44920,N_44952);
nor U46768 (N_46768,N_45419,N_44196);
nand U46769 (N_46769,N_44663,N_44079);
and U46770 (N_46770,N_44076,N_45103);
nand U46771 (N_46771,N_44059,N_45673);
nor U46772 (N_46772,N_45477,N_45955);
nand U46773 (N_46773,N_44375,N_44721);
nor U46774 (N_46774,N_45716,N_45728);
xor U46775 (N_46775,N_45191,N_44734);
and U46776 (N_46776,N_44601,N_44363);
nand U46777 (N_46777,N_44820,N_44760);
xor U46778 (N_46778,N_45863,N_45626);
or U46779 (N_46779,N_44809,N_45037);
and U46780 (N_46780,N_45582,N_45531);
and U46781 (N_46781,N_45320,N_44503);
xor U46782 (N_46782,N_44153,N_44421);
or U46783 (N_46783,N_44302,N_45347);
nor U46784 (N_46784,N_44897,N_45845);
and U46785 (N_46785,N_45889,N_45774);
or U46786 (N_46786,N_44307,N_45374);
xor U46787 (N_46787,N_44009,N_44218);
xor U46788 (N_46788,N_45251,N_45266);
nor U46789 (N_46789,N_44267,N_45899);
or U46790 (N_46790,N_44856,N_45724);
or U46791 (N_46791,N_44676,N_44023);
nor U46792 (N_46792,N_45464,N_45033);
xor U46793 (N_46793,N_44282,N_45696);
and U46794 (N_46794,N_45310,N_45388);
or U46795 (N_46795,N_45215,N_44975);
nor U46796 (N_46796,N_45396,N_45400);
or U46797 (N_46797,N_44762,N_45615);
xnor U46798 (N_46798,N_45799,N_45447);
xnor U46799 (N_46799,N_45360,N_45501);
nand U46800 (N_46800,N_45867,N_44996);
xor U46801 (N_46801,N_44258,N_45778);
xor U46802 (N_46802,N_45055,N_44875);
xor U46803 (N_46803,N_44711,N_44201);
and U46804 (N_46804,N_45177,N_44692);
or U46805 (N_46805,N_45707,N_45007);
xor U46806 (N_46806,N_45657,N_45390);
or U46807 (N_46807,N_44782,N_45490);
nor U46808 (N_46808,N_45651,N_44626);
and U46809 (N_46809,N_44709,N_44811);
or U46810 (N_46810,N_45497,N_44091);
nand U46811 (N_46811,N_45875,N_45325);
and U46812 (N_46812,N_45848,N_45913);
nand U46813 (N_46813,N_44118,N_45969);
nand U46814 (N_46814,N_44110,N_44536);
xnor U46815 (N_46815,N_44339,N_45315);
nor U46816 (N_46816,N_44604,N_44222);
nor U46817 (N_46817,N_45060,N_45445);
and U46818 (N_46818,N_45621,N_44865);
nor U46819 (N_46819,N_44133,N_45579);
or U46820 (N_46820,N_44115,N_45196);
nand U46821 (N_46821,N_44572,N_45467);
xor U46822 (N_46822,N_45538,N_45620);
and U46823 (N_46823,N_45395,N_45928);
nand U46824 (N_46824,N_44465,N_44526);
nor U46825 (N_46825,N_45365,N_44360);
xor U46826 (N_46826,N_44147,N_45589);
and U46827 (N_46827,N_45401,N_44559);
or U46828 (N_46828,N_45676,N_45128);
or U46829 (N_46829,N_45961,N_44362);
or U46830 (N_46830,N_44475,N_45854);
and U46831 (N_46831,N_44182,N_44440);
or U46832 (N_46832,N_45151,N_44446);
nor U46833 (N_46833,N_45459,N_44943);
or U46834 (N_46834,N_45180,N_44832);
or U46835 (N_46835,N_45104,N_45542);
xnor U46836 (N_46836,N_45990,N_45515);
and U46837 (N_46837,N_44065,N_44080);
nor U46838 (N_46838,N_45076,N_45090);
or U46839 (N_46839,N_44040,N_44319);
xnor U46840 (N_46840,N_45671,N_44019);
xor U46841 (N_46841,N_45550,N_44731);
or U46842 (N_46842,N_44599,N_44610);
nor U46843 (N_46843,N_44263,N_44085);
nand U46844 (N_46844,N_45877,N_45344);
xnor U46845 (N_46845,N_44466,N_45351);
xnor U46846 (N_46846,N_44704,N_44054);
nand U46847 (N_46847,N_44336,N_45830);
xor U46848 (N_46848,N_45693,N_44469);
or U46849 (N_46849,N_45233,N_45131);
xor U46850 (N_46850,N_45719,N_45238);
or U46851 (N_46851,N_44652,N_44046);
xor U46852 (N_46852,N_45406,N_45035);
and U46853 (N_46853,N_44108,N_45398);
nor U46854 (N_46854,N_44416,N_45082);
or U46855 (N_46855,N_45509,N_45884);
or U46856 (N_46856,N_45616,N_45691);
or U46857 (N_46857,N_45455,N_44524);
nand U46858 (N_46858,N_45308,N_44577);
and U46859 (N_46859,N_44899,N_44769);
and U46860 (N_46860,N_45232,N_44887);
and U46861 (N_46861,N_44917,N_44861);
or U46862 (N_46862,N_44724,N_44655);
or U46863 (N_46863,N_45603,N_44883);
nand U46864 (N_46864,N_45063,N_44732);
nor U46865 (N_46865,N_45083,N_45963);
and U46866 (N_46866,N_44123,N_44798);
xnor U46867 (N_46867,N_45583,N_44356);
or U46868 (N_46868,N_44893,N_45381);
xnor U46869 (N_46869,N_45261,N_45004);
xnor U46870 (N_46870,N_44470,N_45326);
and U46871 (N_46871,N_45956,N_44203);
and U46872 (N_46872,N_45985,N_44414);
nor U46873 (N_46873,N_45869,N_45423);
or U46874 (N_46874,N_44774,N_45898);
xnor U46875 (N_46875,N_45735,N_45745);
nand U46876 (N_46876,N_44627,N_45656);
nand U46877 (N_46877,N_45008,N_45077);
or U46878 (N_46878,N_44165,N_44767);
or U46879 (N_46879,N_45835,N_45050);
xnor U46880 (N_46880,N_45587,N_44424);
nor U46881 (N_46881,N_45457,N_45852);
xnor U46882 (N_46882,N_44420,N_45089);
or U46883 (N_46883,N_45418,N_44269);
or U46884 (N_46884,N_44011,N_44807);
nand U46885 (N_46885,N_44581,N_44366);
nor U46886 (N_46886,N_44419,N_45556);
xnor U46887 (N_46887,N_44836,N_44757);
xor U46888 (N_46888,N_45149,N_45364);
nor U46889 (N_46889,N_45949,N_45172);
nand U46890 (N_46890,N_45650,N_44253);
or U46891 (N_46891,N_44776,N_45494);
nor U46892 (N_46892,N_44390,N_44327);
or U46893 (N_46893,N_45818,N_45432);
nor U46894 (N_46894,N_44016,N_45540);
nand U46895 (N_46895,N_44545,N_44354);
nor U46896 (N_46896,N_45887,N_44057);
xnor U46897 (N_46897,N_45163,N_45669);
xor U46898 (N_46898,N_45648,N_44699);
nand U46899 (N_46899,N_44254,N_45804);
xnor U46900 (N_46900,N_44244,N_44833);
or U46901 (N_46901,N_45801,N_45979);
or U46902 (N_46902,N_44844,N_44691);
xor U46903 (N_46903,N_44761,N_44457);
nand U46904 (N_46904,N_44322,N_45295);
nand U46905 (N_46905,N_45429,N_44179);
nand U46906 (N_46906,N_44707,N_44490);
nand U46907 (N_46907,N_44885,N_45274);
and U46908 (N_46908,N_44575,N_44866);
and U46909 (N_46909,N_44246,N_44439);
xor U46910 (N_46910,N_45703,N_45392);
and U46911 (N_46911,N_45740,N_44353);
or U46912 (N_46912,N_44159,N_45874);
or U46913 (N_46913,N_45832,N_45827);
or U46914 (N_46914,N_45355,N_44904);
nand U46915 (N_46915,N_45479,N_45165);
or U46916 (N_46916,N_45372,N_45605);
nor U46917 (N_46917,N_44372,N_45179);
and U46918 (N_46918,N_44995,N_45917);
nor U46919 (N_46919,N_44548,N_45681);
and U46920 (N_46920,N_44786,N_45823);
nor U46921 (N_46921,N_45934,N_44225);
nand U46922 (N_46922,N_44257,N_45257);
or U46923 (N_46923,N_44613,N_44922);
nand U46924 (N_46924,N_45533,N_45016);
or U46925 (N_46925,N_44827,N_44072);
xnor U46926 (N_46926,N_45561,N_45399);
or U46927 (N_46927,N_44024,N_45824);
nor U46928 (N_46928,N_45454,N_45437);
xnor U46929 (N_46929,N_44542,N_44212);
nor U46930 (N_46930,N_45842,N_44261);
nand U46931 (N_46931,N_45470,N_44342);
or U46932 (N_46932,N_44911,N_44361);
or U46933 (N_46933,N_45946,N_45087);
and U46934 (N_46934,N_44070,N_45581);
or U46935 (N_46935,N_45790,N_45345);
nor U46936 (N_46936,N_45993,N_44987);
and U46937 (N_46937,N_44491,N_44348);
nand U46938 (N_46938,N_44333,N_44395);
and U46939 (N_46939,N_44884,N_45482);
nand U46940 (N_46940,N_45873,N_45943);
and U46941 (N_46941,N_44283,N_44400);
and U46942 (N_46942,N_44751,N_44397);
nand U46943 (N_46943,N_45604,N_44000);
and U46944 (N_46944,N_44636,N_44380);
nand U46945 (N_46945,N_45838,N_44102);
and U46946 (N_46946,N_44686,N_45337);
nand U46947 (N_46947,N_44868,N_45011);
and U46948 (N_46948,N_44829,N_44101);
nor U46949 (N_46949,N_44799,N_45247);
or U46950 (N_46950,N_44703,N_45021);
xor U46951 (N_46951,N_44138,N_45632);
xor U46952 (N_46952,N_44956,N_45173);
or U46953 (N_46953,N_44067,N_44409);
nand U46954 (N_46954,N_45743,N_44978);
xnor U46955 (N_46955,N_45584,N_45198);
nand U46956 (N_46956,N_44002,N_45714);
or U46957 (N_46957,N_45084,N_45332);
and U46958 (N_46958,N_45498,N_45680);
nand U46959 (N_46959,N_45114,N_44015);
or U46960 (N_46960,N_45631,N_45534);
xnor U46961 (N_46961,N_44047,N_44797);
or U46962 (N_46962,N_45805,N_45881);
or U46963 (N_46963,N_45690,N_44217);
nor U46964 (N_46964,N_45444,N_45225);
and U46965 (N_46965,N_44210,N_45296);
xnor U46966 (N_46966,N_44742,N_45328);
and U46967 (N_46967,N_44418,N_44489);
nor U46968 (N_46968,N_44714,N_44670);
nor U46969 (N_46969,N_45193,N_45098);
nor U46970 (N_46970,N_44831,N_45417);
xnor U46971 (N_46971,N_44403,N_45458);
or U46972 (N_46972,N_44114,N_44765);
or U46973 (N_46973,N_45336,N_44300);
nor U46974 (N_46974,N_44033,N_44050);
or U46975 (N_46975,N_45879,N_45122);
nand U46976 (N_46976,N_44213,N_45070);
nor U46977 (N_46977,N_44215,N_45548);
nand U46978 (N_46978,N_44935,N_44233);
nor U46979 (N_46979,N_45660,N_45038);
nand U46980 (N_46980,N_45178,N_45602);
xor U46981 (N_46981,N_45425,N_44052);
or U46982 (N_46982,N_45769,N_45391);
nor U46983 (N_46983,N_44103,N_45462);
nor U46984 (N_46984,N_44227,N_45263);
and U46985 (N_46985,N_44441,N_44902);
or U46986 (N_46986,N_44954,N_44013);
xnor U46987 (N_46987,N_44748,N_45264);
nor U46988 (N_46988,N_44494,N_44086);
xor U46989 (N_46989,N_45972,N_45654);
and U46990 (N_46990,N_44803,N_44208);
xor U46991 (N_46991,N_44303,N_45022);
nor U46992 (N_46992,N_44723,N_45159);
nor U46993 (N_46993,N_44991,N_45811);
or U46994 (N_46994,N_45436,N_45269);
or U46995 (N_46995,N_45058,N_45802);
or U46996 (N_46996,N_45843,N_45105);
and U46997 (N_46997,N_45526,N_45649);
nand U46998 (N_46998,N_45932,N_45576);
nand U46999 (N_46999,N_44438,N_44970);
nor U47000 (N_47000,N_44369,N_44876);
and U47001 (N_47001,N_44893,N_44745);
or U47002 (N_47002,N_45181,N_44504);
nand U47003 (N_47003,N_45978,N_44156);
nor U47004 (N_47004,N_45336,N_45937);
nor U47005 (N_47005,N_44207,N_45290);
xnor U47006 (N_47006,N_45569,N_45222);
nand U47007 (N_47007,N_45531,N_45071);
or U47008 (N_47008,N_45639,N_44460);
and U47009 (N_47009,N_45547,N_45440);
or U47010 (N_47010,N_44254,N_45122);
and U47011 (N_47011,N_44703,N_44817);
and U47012 (N_47012,N_45016,N_45255);
xor U47013 (N_47013,N_44467,N_45396);
xor U47014 (N_47014,N_44661,N_44105);
nand U47015 (N_47015,N_44099,N_45788);
and U47016 (N_47016,N_44379,N_44117);
xnor U47017 (N_47017,N_45898,N_45527);
nand U47018 (N_47018,N_45526,N_45867);
nand U47019 (N_47019,N_44668,N_45087);
nand U47020 (N_47020,N_44831,N_45964);
nor U47021 (N_47021,N_44404,N_44989);
nor U47022 (N_47022,N_45854,N_45479);
and U47023 (N_47023,N_44164,N_44978);
and U47024 (N_47024,N_44641,N_44186);
xnor U47025 (N_47025,N_45370,N_44570);
nor U47026 (N_47026,N_44104,N_45988);
xnor U47027 (N_47027,N_45375,N_45422);
or U47028 (N_47028,N_44694,N_45808);
nor U47029 (N_47029,N_45000,N_45690);
or U47030 (N_47030,N_44202,N_44035);
or U47031 (N_47031,N_45767,N_45439);
or U47032 (N_47032,N_44315,N_44895);
and U47033 (N_47033,N_44647,N_45734);
nand U47034 (N_47034,N_45099,N_44455);
xnor U47035 (N_47035,N_44810,N_45362);
nand U47036 (N_47036,N_44558,N_45086);
or U47037 (N_47037,N_45286,N_44358);
and U47038 (N_47038,N_45937,N_45717);
and U47039 (N_47039,N_44128,N_45080);
nor U47040 (N_47040,N_44489,N_45976);
nor U47041 (N_47041,N_44152,N_44321);
or U47042 (N_47042,N_44996,N_44415);
nor U47043 (N_47043,N_44029,N_45734);
xnor U47044 (N_47044,N_44493,N_45607);
or U47045 (N_47045,N_44892,N_45710);
and U47046 (N_47046,N_45978,N_44077);
or U47047 (N_47047,N_45448,N_44758);
or U47048 (N_47048,N_45164,N_45938);
nand U47049 (N_47049,N_44394,N_44365);
nand U47050 (N_47050,N_45098,N_45827);
and U47051 (N_47051,N_45851,N_44667);
and U47052 (N_47052,N_44962,N_45474);
nand U47053 (N_47053,N_44618,N_44704);
xor U47054 (N_47054,N_44224,N_45633);
or U47055 (N_47055,N_44161,N_45969);
xor U47056 (N_47056,N_45710,N_45385);
xor U47057 (N_47057,N_44539,N_45367);
and U47058 (N_47058,N_44453,N_45437);
nand U47059 (N_47059,N_44014,N_45762);
nor U47060 (N_47060,N_45428,N_44203);
or U47061 (N_47061,N_44931,N_45954);
or U47062 (N_47062,N_44609,N_44701);
and U47063 (N_47063,N_45570,N_45907);
or U47064 (N_47064,N_44119,N_44095);
nand U47065 (N_47065,N_44948,N_45272);
and U47066 (N_47066,N_45693,N_45955);
and U47067 (N_47067,N_45339,N_44184);
or U47068 (N_47068,N_44637,N_45932);
nand U47069 (N_47069,N_44874,N_44612);
and U47070 (N_47070,N_45941,N_44246);
nand U47071 (N_47071,N_45793,N_45960);
and U47072 (N_47072,N_44903,N_44818);
nand U47073 (N_47073,N_44658,N_45595);
or U47074 (N_47074,N_44367,N_45599);
or U47075 (N_47075,N_44288,N_45352);
or U47076 (N_47076,N_44703,N_45979);
nor U47077 (N_47077,N_45404,N_44905);
or U47078 (N_47078,N_45000,N_45873);
or U47079 (N_47079,N_44608,N_44841);
nor U47080 (N_47080,N_45703,N_44487);
nand U47081 (N_47081,N_45258,N_44620);
and U47082 (N_47082,N_45701,N_45024);
xor U47083 (N_47083,N_44899,N_44977);
xnor U47084 (N_47084,N_44931,N_45327);
xnor U47085 (N_47085,N_44568,N_45603);
nor U47086 (N_47086,N_44403,N_44272);
nor U47087 (N_47087,N_45606,N_44145);
nand U47088 (N_47088,N_44522,N_44725);
nand U47089 (N_47089,N_44862,N_45149);
nand U47090 (N_47090,N_44596,N_44372);
or U47091 (N_47091,N_45632,N_45742);
nand U47092 (N_47092,N_45465,N_45975);
and U47093 (N_47093,N_44482,N_44067);
nor U47094 (N_47094,N_44243,N_45393);
nor U47095 (N_47095,N_44056,N_44974);
xor U47096 (N_47096,N_44862,N_44524);
nor U47097 (N_47097,N_45133,N_44153);
nand U47098 (N_47098,N_44695,N_44863);
and U47099 (N_47099,N_45037,N_45776);
nor U47100 (N_47100,N_45773,N_44821);
nand U47101 (N_47101,N_45577,N_44669);
and U47102 (N_47102,N_45404,N_45662);
and U47103 (N_47103,N_44996,N_44662);
nor U47104 (N_47104,N_45022,N_45567);
and U47105 (N_47105,N_44480,N_44608);
or U47106 (N_47106,N_44582,N_44804);
and U47107 (N_47107,N_45656,N_44335);
or U47108 (N_47108,N_45754,N_44651);
nor U47109 (N_47109,N_44409,N_45215);
nor U47110 (N_47110,N_45871,N_44829);
xnor U47111 (N_47111,N_45157,N_45556);
nand U47112 (N_47112,N_45110,N_45149);
nor U47113 (N_47113,N_44454,N_45197);
xor U47114 (N_47114,N_44680,N_44102);
or U47115 (N_47115,N_44745,N_44597);
or U47116 (N_47116,N_44012,N_44944);
xnor U47117 (N_47117,N_44924,N_44754);
nor U47118 (N_47118,N_45471,N_44549);
xnor U47119 (N_47119,N_45762,N_44165);
xor U47120 (N_47120,N_44155,N_44695);
or U47121 (N_47121,N_44603,N_44362);
nor U47122 (N_47122,N_45092,N_44449);
xnor U47123 (N_47123,N_44154,N_44800);
or U47124 (N_47124,N_45969,N_44206);
nor U47125 (N_47125,N_45892,N_44494);
nand U47126 (N_47126,N_45261,N_44400);
nand U47127 (N_47127,N_44263,N_44885);
nand U47128 (N_47128,N_44206,N_45760);
and U47129 (N_47129,N_45114,N_45491);
nand U47130 (N_47130,N_45781,N_44705);
or U47131 (N_47131,N_45276,N_45531);
nor U47132 (N_47132,N_44628,N_44924);
nor U47133 (N_47133,N_44710,N_44527);
nand U47134 (N_47134,N_45790,N_45244);
and U47135 (N_47135,N_45200,N_44853);
and U47136 (N_47136,N_45203,N_45880);
xnor U47137 (N_47137,N_45674,N_45596);
nand U47138 (N_47138,N_44792,N_45488);
nor U47139 (N_47139,N_45166,N_44635);
nor U47140 (N_47140,N_44556,N_45948);
or U47141 (N_47141,N_45080,N_44949);
nor U47142 (N_47142,N_45997,N_45446);
and U47143 (N_47143,N_45082,N_45621);
and U47144 (N_47144,N_45857,N_45497);
xor U47145 (N_47145,N_44483,N_44235);
nand U47146 (N_47146,N_44445,N_44459);
nor U47147 (N_47147,N_44823,N_45537);
nand U47148 (N_47148,N_44039,N_44276);
xor U47149 (N_47149,N_45529,N_45022);
nand U47150 (N_47150,N_44089,N_45944);
xnor U47151 (N_47151,N_44387,N_44584);
xor U47152 (N_47152,N_44452,N_45531);
and U47153 (N_47153,N_44917,N_44737);
or U47154 (N_47154,N_44485,N_44889);
or U47155 (N_47155,N_45098,N_44725);
or U47156 (N_47156,N_44299,N_45263);
xnor U47157 (N_47157,N_45829,N_44916);
xnor U47158 (N_47158,N_45338,N_45179);
or U47159 (N_47159,N_45574,N_44666);
nand U47160 (N_47160,N_44349,N_45071);
nand U47161 (N_47161,N_44275,N_45611);
nor U47162 (N_47162,N_44172,N_45113);
or U47163 (N_47163,N_45637,N_45045);
nand U47164 (N_47164,N_45854,N_45090);
or U47165 (N_47165,N_45887,N_44542);
and U47166 (N_47166,N_45550,N_44259);
and U47167 (N_47167,N_44299,N_44449);
xnor U47168 (N_47168,N_44457,N_44916);
and U47169 (N_47169,N_44641,N_45624);
nand U47170 (N_47170,N_45239,N_45376);
nor U47171 (N_47171,N_44442,N_44670);
or U47172 (N_47172,N_45710,N_45897);
nand U47173 (N_47173,N_44127,N_45672);
or U47174 (N_47174,N_44342,N_44790);
or U47175 (N_47175,N_44888,N_45136);
xor U47176 (N_47176,N_44897,N_44442);
or U47177 (N_47177,N_45134,N_44421);
and U47178 (N_47178,N_45856,N_45617);
nor U47179 (N_47179,N_45597,N_45021);
and U47180 (N_47180,N_45260,N_44494);
xor U47181 (N_47181,N_44988,N_44338);
nor U47182 (N_47182,N_45752,N_44442);
or U47183 (N_47183,N_44447,N_44744);
or U47184 (N_47184,N_44811,N_45958);
xor U47185 (N_47185,N_44137,N_44314);
nand U47186 (N_47186,N_44567,N_45840);
nor U47187 (N_47187,N_44126,N_45655);
xor U47188 (N_47188,N_44206,N_45909);
and U47189 (N_47189,N_45843,N_44587);
or U47190 (N_47190,N_44154,N_44899);
and U47191 (N_47191,N_44158,N_45234);
nand U47192 (N_47192,N_44705,N_45307);
or U47193 (N_47193,N_44456,N_45120);
or U47194 (N_47194,N_45653,N_44360);
nand U47195 (N_47195,N_44868,N_45472);
nor U47196 (N_47196,N_45798,N_45897);
xnor U47197 (N_47197,N_45534,N_45929);
nand U47198 (N_47198,N_44352,N_44485);
and U47199 (N_47199,N_45242,N_44981);
nand U47200 (N_47200,N_44174,N_45014);
and U47201 (N_47201,N_45169,N_45478);
or U47202 (N_47202,N_44465,N_45067);
nor U47203 (N_47203,N_45544,N_44210);
nor U47204 (N_47204,N_44171,N_45494);
nand U47205 (N_47205,N_44542,N_44722);
xor U47206 (N_47206,N_45984,N_45258);
xor U47207 (N_47207,N_44009,N_45544);
and U47208 (N_47208,N_44063,N_44412);
nor U47209 (N_47209,N_45598,N_45630);
xnor U47210 (N_47210,N_45128,N_44446);
and U47211 (N_47211,N_44492,N_45832);
xnor U47212 (N_47212,N_45431,N_44687);
nand U47213 (N_47213,N_45757,N_44545);
nand U47214 (N_47214,N_44151,N_45258);
xor U47215 (N_47215,N_45760,N_44000);
or U47216 (N_47216,N_45745,N_44028);
xnor U47217 (N_47217,N_45168,N_45948);
nand U47218 (N_47218,N_44532,N_44214);
or U47219 (N_47219,N_44253,N_45851);
nor U47220 (N_47220,N_44308,N_45649);
nor U47221 (N_47221,N_45728,N_44534);
nor U47222 (N_47222,N_44786,N_45699);
nand U47223 (N_47223,N_45790,N_44950);
nor U47224 (N_47224,N_45276,N_45613);
xnor U47225 (N_47225,N_45618,N_45723);
or U47226 (N_47226,N_44389,N_45714);
or U47227 (N_47227,N_45111,N_45346);
nor U47228 (N_47228,N_45020,N_45472);
and U47229 (N_47229,N_44082,N_45455);
nand U47230 (N_47230,N_45063,N_44851);
or U47231 (N_47231,N_45351,N_45804);
xnor U47232 (N_47232,N_45056,N_45720);
nor U47233 (N_47233,N_45108,N_44527);
xnor U47234 (N_47234,N_45951,N_44809);
nand U47235 (N_47235,N_45179,N_45143);
nor U47236 (N_47236,N_44235,N_45586);
xor U47237 (N_47237,N_44009,N_44611);
nor U47238 (N_47238,N_45428,N_44231);
nor U47239 (N_47239,N_44850,N_44220);
or U47240 (N_47240,N_44305,N_44252);
xor U47241 (N_47241,N_45217,N_45040);
and U47242 (N_47242,N_44648,N_44876);
or U47243 (N_47243,N_45321,N_45291);
nand U47244 (N_47244,N_45496,N_45309);
and U47245 (N_47245,N_44086,N_45089);
and U47246 (N_47246,N_44840,N_45411);
nor U47247 (N_47247,N_44717,N_45510);
and U47248 (N_47248,N_44123,N_45940);
nand U47249 (N_47249,N_44954,N_44565);
xnor U47250 (N_47250,N_44096,N_45533);
or U47251 (N_47251,N_44221,N_44112);
xnor U47252 (N_47252,N_44264,N_44649);
nor U47253 (N_47253,N_45150,N_44869);
and U47254 (N_47254,N_45375,N_45921);
xnor U47255 (N_47255,N_44013,N_45496);
xor U47256 (N_47256,N_45161,N_45499);
nor U47257 (N_47257,N_44155,N_45400);
nand U47258 (N_47258,N_44233,N_44162);
xor U47259 (N_47259,N_45353,N_45230);
nand U47260 (N_47260,N_45025,N_44445);
xor U47261 (N_47261,N_45008,N_45759);
nor U47262 (N_47262,N_44813,N_44530);
xnor U47263 (N_47263,N_44405,N_44488);
and U47264 (N_47264,N_44025,N_44384);
xnor U47265 (N_47265,N_44145,N_44749);
nor U47266 (N_47266,N_45386,N_45704);
and U47267 (N_47267,N_44902,N_45596);
and U47268 (N_47268,N_44395,N_45786);
nand U47269 (N_47269,N_44000,N_44411);
or U47270 (N_47270,N_44353,N_44623);
and U47271 (N_47271,N_44405,N_45524);
nand U47272 (N_47272,N_44662,N_45660);
and U47273 (N_47273,N_45411,N_45653);
or U47274 (N_47274,N_44644,N_44999);
or U47275 (N_47275,N_44229,N_44472);
xor U47276 (N_47276,N_45338,N_45272);
and U47277 (N_47277,N_45972,N_44014);
nor U47278 (N_47278,N_45780,N_44403);
nand U47279 (N_47279,N_45185,N_44808);
xnor U47280 (N_47280,N_44728,N_45113);
nor U47281 (N_47281,N_44726,N_44009);
xnor U47282 (N_47282,N_45335,N_44469);
and U47283 (N_47283,N_44797,N_44462);
and U47284 (N_47284,N_45193,N_45568);
and U47285 (N_47285,N_44690,N_45666);
xor U47286 (N_47286,N_45637,N_44323);
or U47287 (N_47287,N_44694,N_45675);
nor U47288 (N_47288,N_44441,N_45159);
nand U47289 (N_47289,N_44925,N_44427);
xnor U47290 (N_47290,N_44648,N_45173);
or U47291 (N_47291,N_45678,N_45451);
xnor U47292 (N_47292,N_45444,N_45971);
nor U47293 (N_47293,N_44813,N_44341);
xor U47294 (N_47294,N_44514,N_45665);
nor U47295 (N_47295,N_44778,N_45023);
nand U47296 (N_47296,N_45728,N_45668);
nand U47297 (N_47297,N_45260,N_45932);
or U47298 (N_47298,N_44515,N_44529);
and U47299 (N_47299,N_44342,N_44579);
or U47300 (N_47300,N_45729,N_45535);
or U47301 (N_47301,N_44773,N_44367);
or U47302 (N_47302,N_45132,N_45685);
nand U47303 (N_47303,N_44862,N_45396);
nor U47304 (N_47304,N_44722,N_44994);
nand U47305 (N_47305,N_45640,N_45383);
or U47306 (N_47306,N_45193,N_45003);
or U47307 (N_47307,N_44690,N_44754);
nand U47308 (N_47308,N_44761,N_44348);
or U47309 (N_47309,N_45860,N_45563);
nor U47310 (N_47310,N_44249,N_44638);
xnor U47311 (N_47311,N_44614,N_45887);
and U47312 (N_47312,N_44669,N_44498);
nand U47313 (N_47313,N_44015,N_44004);
or U47314 (N_47314,N_44847,N_45433);
nand U47315 (N_47315,N_44551,N_45982);
nand U47316 (N_47316,N_45714,N_44483);
nor U47317 (N_47317,N_44154,N_45695);
nand U47318 (N_47318,N_45970,N_45467);
nor U47319 (N_47319,N_45840,N_45029);
nand U47320 (N_47320,N_45815,N_44774);
nor U47321 (N_47321,N_44585,N_45766);
or U47322 (N_47322,N_45517,N_45821);
nor U47323 (N_47323,N_44229,N_44606);
xnor U47324 (N_47324,N_44264,N_44833);
xnor U47325 (N_47325,N_44922,N_45666);
nor U47326 (N_47326,N_44850,N_45917);
nor U47327 (N_47327,N_44147,N_44123);
or U47328 (N_47328,N_45557,N_44088);
nand U47329 (N_47329,N_44185,N_44873);
nor U47330 (N_47330,N_44685,N_44337);
nand U47331 (N_47331,N_45589,N_44095);
and U47332 (N_47332,N_45503,N_45650);
and U47333 (N_47333,N_44592,N_44521);
xnor U47334 (N_47334,N_44848,N_45663);
and U47335 (N_47335,N_45323,N_44196);
or U47336 (N_47336,N_45639,N_44438);
and U47337 (N_47337,N_45583,N_45723);
and U47338 (N_47338,N_44993,N_45473);
nand U47339 (N_47339,N_45678,N_44965);
xor U47340 (N_47340,N_45439,N_45761);
nand U47341 (N_47341,N_44652,N_44248);
nand U47342 (N_47342,N_44204,N_45227);
nand U47343 (N_47343,N_44762,N_45724);
and U47344 (N_47344,N_45814,N_45678);
nor U47345 (N_47345,N_44793,N_45075);
xor U47346 (N_47346,N_44720,N_44867);
nand U47347 (N_47347,N_44554,N_45206);
nand U47348 (N_47348,N_45135,N_44735);
and U47349 (N_47349,N_44343,N_45541);
and U47350 (N_47350,N_44831,N_44701);
xnor U47351 (N_47351,N_44347,N_44760);
and U47352 (N_47352,N_45681,N_44501);
and U47353 (N_47353,N_44354,N_44004);
and U47354 (N_47354,N_44207,N_45892);
or U47355 (N_47355,N_45560,N_44350);
or U47356 (N_47356,N_45859,N_45869);
xor U47357 (N_47357,N_45451,N_45943);
xor U47358 (N_47358,N_45892,N_44849);
and U47359 (N_47359,N_44244,N_44595);
and U47360 (N_47360,N_44123,N_45289);
xnor U47361 (N_47361,N_45875,N_45006);
nand U47362 (N_47362,N_45064,N_45343);
nand U47363 (N_47363,N_45848,N_45807);
or U47364 (N_47364,N_44791,N_45955);
xnor U47365 (N_47365,N_44908,N_44886);
nor U47366 (N_47366,N_45502,N_45684);
xnor U47367 (N_47367,N_44973,N_44640);
nor U47368 (N_47368,N_44453,N_44173);
or U47369 (N_47369,N_44440,N_44865);
nor U47370 (N_47370,N_44593,N_45605);
nand U47371 (N_47371,N_45604,N_44026);
xor U47372 (N_47372,N_45561,N_45704);
and U47373 (N_47373,N_44955,N_45978);
and U47374 (N_47374,N_45059,N_44631);
and U47375 (N_47375,N_44202,N_44443);
nand U47376 (N_47376,N_45939,N_44901);
or U47377 (N_47377,N_44997,N_44353);
nand U47378 (N_47378,N_44580,N_44820);
and U47379 (N_47379,N_45533,N_45682);
nor U47380 (N_47380,N_45063,N_45585);
and U47381 (N_47381,N_44326,N_45189);
or U47382 (N_47382,N_45189,N_45524);
nand U47383 (N_47383,N_45497,N_45453);
nor U47384 (N_47384,N_45742,N_45416);
nor U47385 (N_47385,N_45739,N_44647);
nand U47386 (N_47386,N_45325,N_45742);
and U47387 (N_47387,N_44357,N_44602);
nand U47388 (N_47388,N_45842,N_44541);
nand U47389 (N_47389,N_44967,N_45177);
nand U47390 (N_47390,N_44761,N_45044);
and U47391 (N_47391,N_45049,N_44582);
nor U47392 (N_47392,N_44314,N_44752);
or U47393 (N_47393,N_44175,N_45731);
nor U47394 (N_47394,N_45404,N_44376);
xor U47395 (N_47395,N_45075,N_45179);
or U47396 (N_47396,N_45905,N_44822);
and U47397 (N_47397,N_44633,N_44395);
nand U47398 (N_47398,N_45146,N_44367);
nor U47399 (N_47399,N_45638,N_45342);
or U47400 (N_47400,N_45242,N_44796);
nand U47401 (N_47401,N_44084,N_45484);
nand U47402 (N_47402,N_44503,N_45545);
and U47403 (N_47403,N_44391,N_45766);
and U47404 (N_47404,N_45440,N_45962);
xor U47405 (N_47405,N_45264,N_44006);
or U47406 (N_47406,N_44616,N_44169);
nand U47407 (N_47407,N_44713,N_44633);
xnor U47408 (N_47408,N_44961,N_45475);
and U47409 (N_47409,N_44843,N_45501);
and U47410 (N_47410,N_45537,N_44934);
and U47411 (N_47411,N_45384,N_45723);
xor U47412 (N_47412,N_44248,N_45961);
or U47413 (N_47413,N_45395,N_44969);
xnor U47414 (N_47414,N_44404,N_44211);
nor U47415 (N_47415,N_44590,N_45483);
and U47416 (N_47416,N_45016,N_44342);
nand U47417 (N_47417,N_45487,N_45963);
or U47418 (N_47418,N_45923,N_45478);
and U47419 (N_47419,N_44800,N_44127);
or U47420 (N_47420,N_44900,N_44243);
and U47421 (N_47421,N_45515,N_45570);
or U47422 (N_47422,N_45539,N_45685);
xor U47423 (N_47423,N_45509,N_45874);
nor U47424 (N_47424,N_45995,N_45150);
nand U47425 (N_47425,N_44984,N_45814);
nand U47426 (N_47426,N_45761,N_44992);
xnor U47427 (N_47427,N_44710,N_44746);
nand U47428 (N_47428,N_45024,N_45767);
and U47429 (N_47429,N_45034,N_45933);
nor U47430 (N_47430,N_44969,N_45345);
nor U47431 (N_47431,N_45826,N_44822);
nor U47432 (N_47432,N_45157,N_44802);
and U47433 (N_47433,N_44660,N_45248);
or U47434 (N_47434,N_45184,N_44895);
or U47435 (N_47435,N_45346,N_44021);
nor U47436 (N_47436,N_44361,N_45658);
xor U47437 (N_47437,N_45320,N_44550);
xnor U47438 (N_47438,N_45076,N_44108);
or U47439 (N_47439,N_44216,N_45849);
nand U47440 (N_47440,N_45203,N_45047);
and U47441 (N_47441,N_45396,N_44185);
and U47442 (N_47442,N_45001,N_44554);
or U47443 (N_47443,N_45136,N_44924);
xnor U47444 (N_47444,N_45808,N_44898);
nand U47445 (N_47445,N_44970,N_44114);
nand U47446 (N_47446,N_45599,N_44862);
and U47447 (N_47447,N_44039,N_44169);
xnor U47448 (N_47448,N_44334,N_45034);
nor U47449 (N_47449,N_44234,N_44215);
nand U47450 (N_47450,N_45502,N_44438);
and U47451 (N_47451,N_44883,N_45480);
xnor U47452 (N_47452,N_45061,N_45878);
nand U47453 (N_47453,N_44135,N_44629);
xor U47454 (N_47454,N_44055,N_44566);
nand U47455 (N_47455,N_45885,N_45956);
xor U47456 (N_47456,N_44222,N_44493);
nor U47457 (N_47457,N_45792,N_45406);
nand U47458 (N_47458,N_45178,N_45825);
and U47459 (N_47459,N_44551,N_45279);
xnor U47460 (N_47460,N_44793,N_44052);
or U47461 (N_47461,N_45049,N_45637);
nor U47462 (N_47462,N_44632,N_44664);
nand U47463 (N_47463,N_44165,N_45280);
or U47464 (N_47464,N_44170,N_45965);
or U47465 (N_47465,N_45545,N_45722);
nand U47466 (N_47466,N_45718,N_45604);
or U47467 (N_47467,N_45696,N_45410);
xor U47468 (N_47468,N_45774,N_44193);
nor U47469 (N_47469,N_44940,N_44625);
nor U47470 (N_47470,N_44772,N_45653);
xnor U47471 (N_47471,N_45900,N_45501);
or U47472 (N_47472,N_44449,N_45022);
and U47473 (N_47473,N_44727,N_44619);
nand U47474 (N_47474,N_44043,N_45195);
and U47475 (N_47475,N_44571,N_44353);
nor U47476 (N_47476,N_45448,N_45236);
xnor U47477 (N_47477,N_45328,N_45281);
and U47478 (N_47478,N_44495,N_45838);
nor U47479 (N_47479,N_45362,N_44670);
and U47480 (N_47480,N_44271,N_44652);
and U47481 (N_47481,N_44911,N_44309);
nand U47482 (N_47482,N_45740,N_44246);
nand U47483 (N_47483,N_44660,N_45123);
nor U47484 (N_47484,N_45225,N_45592);
nor U47485 (N_47485,N_45917,N_44649);
nor U47486 (N_47486,N_45077,N_45599);
xor U47487 (N_47487,N_45222,N_44592);
and U47488 (N_47488,N_44974,N_44186);
nor U47489 (N_47489,N_45958,N_44704);
nor U47490 (N_47490,N_45600,N_45681);
or U47491 (N_47491,N_45336,N_45775);
and U47492 (N_47492,N_44714,N_45459);
nand U47493 (N_47493,N_45266,N_45838);
xnor U47494 (N_47494,N_44388,N_45599);
and U47495 (N_47495,N_45500,N_44706);
nor U47496 (N_47496,N_44821,N_44068);
and U47497 (N_47497,N_45123,N_45174);
nor U47498 (N_47498,N_45939,N_44214);
or U47499 (N_47499,N_45673,N_44155);
nand U47500 (N_47500,N_44306,N_45633);
nand U47501 (N_47501,N_45750,N_44651);
xnor U47502 (N_47502,N_44724,N_44059);
nand U47503 (N_47503,N_44674,N_44442);
nor U47504 (N_47504,N_44137,N_45618);
nor U47505 (N_47505,N_45098,N_45401);
xnor U47506 (N_47506,N_45522,N_44649);
and U47507 (N_47507,N_45616,N_44772);
nand U47508 (N_47508,N_45643,N_44604);
and U47509 (N_47509,N_44085,N_45608);
xor U47510 (N_47510,N_44738,N_44558);
nor U47511 (N_47511,N_45834,N_45451);
nor U47512 (N_47512,N_45794,N_44648);
or U47513 (N_47513,N_45526,N_45784);
nor U47514 (N_47514,N_44441,N_44131);
xor U47515 (N_47515,N_45566,N_45202);
xor U47516 (N_47516,N_45749,N_45507);
nand U47517 (N_47517,N_45999,N_44846);
and U47518 (N_47518,N_45978,N_44293);
or U47519 (N_47519,N_44728,N_44054);
nor U47520 (N_47520,N_44404,N_44813);
or U47521 (N_47521,N_44864,N_45606);
and U47522 (N_47522,N_44298,N_44349);
nand U47523 (N_47523,N_45294,N_44020);
or U47524 (N_47524,N_45161,N_45397);
nor U47525 (N_47525,N_45857,N_45938);
xnor U47526 (N_47526,N_45928,N_44236);
xor U47527 (N_47527,N_45406,N_44169);
nand U47528 (N_47528,N_44699,N_45571);
nor U47529 (N_47529,N_44587,N_44233);
and U47530 (N_47530,N_45836,N_45517);
xnor U47531 (N_47531,N_44861,N_45217);
and U47532 (N_47532,N_45892,N_45139);
and U47533 (N_47533,N_44844,N_45852);
or U47534 (N_47534,N_45787,N_44818);
nor U47535 (N_47535,N_45804,N_44416);
nand U47536 (N_47536,N_45638,N_45919);
nor U47537 (N_47537,N_45992,N_44453);
or U47538 (N_47538,N_44639,N_45751);
xor U47539 (N_47539,N_45363,N_45019);
nand U47540 (N_47540,N_44357,N_44861);
nand U47541 (N_47541,N_44797,N_44865);
xor U47542 (N_47542,N_44959,N_45293);
nand U47543 (N_47543,N_45974,N_44792);
and U47544 (N_47544,N_45105,N_44298);
and U47545 (N_47545,N_45952,N_44063);
xnor U47546 (N_47546,N_44143,N_44614);
or U47547 (N_47547,N_44776,N_44191);
xnor U47548 (N_47548,N_45242,N_44363);
nand U47549 (N_47549,N_44120,N_45456);
nand U47550 (N_47550,N_45172,N_44210);
and U47551 (N_47551,N_45097,N_45110);
xor U47552 (N_47552,N_45013,N_44302);
nor U47553 (N_47553,N_44849,N_45985);
and U47554 (N_47554,N_44803,N_45933);
xnor U47555 (N_47555,N_45245,N_45785);
nand U47556 (N_47556,N_45337,N_44494);
nand U47557 (N_47557,N_45734,N_45515);
xor U47558 (N_47558,N_44454,N_44274);
xor U47559 (N_47559,N_45637,N_45883);
nor U47560 (N_47560,N_45588,N_44342);
xor U47561 (N_47561,N_44079,N_44377);
nand U47562 (N_47562,N_45250,N_44905);
and U47563 (N_47563,N_44008,N_45886);
nor U47564 (N_47564,N_45987,N_44550);
xor U47565 (N_47565,N_44501,N_45325);
nor U47566 (N_47566,N_44191,N_44936);
and U47567 (N_47567,N_44335,N_44358);
or U47568 (N_47568,N_45259,N_44222);
and U47569 (N_47569,N_44378,N_45863);
nand U47570 (N_47570,N_44796,N_44841);
xor U47571 (N_47571,N_44696,N_45916);
nor U47572 (N_47572,N_44019,N_45832);
or U47573 (N_47573,N_45540,N_44017);
and U47574 (N_47574,N_45620,N_45717);
and U47575 (N_47575,N_45808,N_44932);
nand U47576 (N_47576,N_44720,N_44415);
xor U47577 (N_47577,N_45125,N_45394);
xnor U47578 (N_47578,N_44402,N_44629);
xor U47579 (N_47579,N_45615,N_45185);
xor U47580 (N_47580,N_45843,N_45854);
xnor U47581 (N_47581,N_45092,N_45383);
nand U47582 (N_47582,N_44607,N_45847);
nand U47583 (N_47583,N_44677,N_45657);
nor U47584 (N_47584,N_45015,N_44527);
xor U47585 (N_47585,N_45557,N_45817);
and U47586 (N_47586,N_45991,N_44315);
nand U47587 (N_47587,N_45983,N_44168);
nand U47588 (N_47588,N_45199,N_45927);
and U47589 (N_47589,N_44289,N_45002);
or U47590 (N_47590,N_45241,N_44599);
nand U47591 (N_47591,N_44821,N_45253);
and U47592 (N_47592,N_45966,N_44969);
xnor U47593 (N_47593,N_44890,N_45669);
nor U47594 (N_47594,N_44970,N_44145);
or U47595 (N_47595,N_44289,N_44377);
nor U47596 (N_47596,N_45395,N_45042);
xor U47597 (N_47597,N_44349,N_44807);
nor U47598 (N_47598,N_44476,N_44158);
xnor U47599 (N_47599,N_44444,N_44710);
or U47600 (N_47600,N_45902,N_44325);
xnor U47601 (N_47601,N_45133,N_45588);
and U47602 (N_47602,N_44775,N_44568);
nand U47603 (N_47603,N_44945,N_44638);
and U47604 (N_47604,N_44846,N_44624);
nor U47605 (N_47605,N_45582,N_45487);
or U47606 (N_47606,N_45959,N_44581);
xor U47607 (N_47607,N_45709,N_44511);
nand U47608 (N_47608,N_45578,N_44346);
or U47609 (N_47609,N_44816,N_44711);
nor U47610 (N_47610,N_45850,N_45799);
or U47611 (N_47611,N_45615,N_45144);
xor U47612 (N_47612,N_44979,N_45387);
xnor U47613 (N_47613,N_44576,N_45518);
nor U47614 (N_47614,N_44542,N_45840);
or U47615 (N_47615,N_45701,N_45679);
nand U47616 (N_47616,N_44275,N_45363);
xor U47617 (N_47617,N_44598,N_45668);
xnor U47618 (N_47618,N_44607,N_44904);
nand U47619 (N_47619,N_44966,N_44834);
or U47620 (N_47620,N_44166,N_44053);
or U47621 (N_47621,N_45987,N_45590);
or U47622 (N_47622,N_44874,N_44977);
nor U47623 (N_47623,N_44284,N_44436);
nor U47624 (N_47624,N_44434,N_45760);
and U47625 (N_47625,N_45503,N_44279);
and U47626 (N_47626,N_44790,N_44490);
nand U47627 (N_47627,N_45303,N_45438);
or U47628 (N_47628,N_45475,N_44327);
or U47629 (N_47629,N_45623,N_44137);
and U47630 (N_47630,N_45812,N_44306);
and U47631 (N_47631,N_44541,N_44002);
xnor U47632 (N_47632,N_45745,N_45148);
nor U47633 (N_47633,N_44179,N_44983);
xnor U47634 (N_47634,N_45043,N_45996);
nand U47635 (N_47635,N_44158,N_45872);
or U47636 (N_47636,N_45603,N_44744);
or U47637 (N_47637,N_45601,N_44741);
or U47638 (N_47638,N_45341,N_45408);
or U47639 (N_47639,N_44191,N_44746);
or U47640 (N_47640,N_45709,N_44815);
nor U47641 (N_47641,N_44194,N_44602);
xor U47642 (N_47642,N_45941,N_45093);
or U47643 (N_47643,N_45845,N_45252);
nor U47644 (N_47644,N_44566,N_45211);
and U47645 (N_47645,N_45939,N_45903);
nand U47646 (N_47646,N_44828,N_44169);
nand U47647 (N_47647,N_44619,N_44307);
nand U47648 (N_47648,N_45571,N_44416);
and U47649 (N_47649,N_44574,N_45548);
nor U47650 (N_47650,N_45220,N_44342);
and U47651 (N_47651,N_44228,N_45648);
xor U47652 (N_47652,N_45814,N_44820);
xnor U47653 (N_47653,N_44834,N_45744);
xor U47654 (N_47654,N_44490,N_45762);
xor U47655 (N_47655,N_44766,N_45308);
or U47656 (N_47656,N_45232,N_45978);
nand U47657 (N_47657,N_44293,N_45285);
and U47658 (N_47658,N_44224,N_45995);
and U47659 (N_47659,N_44745,N_45973);
nand U47660 (N_47660,N_44992,N_45269);
nor U47661 (N_47661,N_44543,N_45034);
or U47662 (N_47662,N_44127,N_44420);
or U47663 (N_47663,N_45270,N_45950);
nand U47664 (N_47664,N_45628,N_44647);
xnor U47665 (N_47665,N_44931,N_45142);
xor U47666 (N_47666,N_45120,N_44733);
nor U47667 (N_47667,N_45626,N_45167);
and U47668 (N_47668,N_44307,N_45615);
nor U47669 (N_47669,N_45822,N_45944);
or U47670 (N_47670,N_45263,N_44147);
nor U47671 (N_47671,N_45038,N_44296);
xnor U47672 (N_47672,N_44311,N_45637);
nand U47673 (N_47673,N_45432,N_44505);
nand U47674 (N_47674,N_44151,N_44719);
nor U47675 (N_47675,N_44762,N_44021);
nand U47676 (N_47676,N_44585,N_44817);
and U47677 (N_47677,N_45277,N_44087);
and U47678 (N_47678,N_45999,N_44590);
nor U47679 (N_47679,N_45780,N_44269);
and U47680 (N_47680,N_44822,N_45054);
and U47681 (N_47681,N_45179,N_45679);
nand U47682 (N_47682,N_44233,N_45497);
or U47683 (N_47683,N_44743,N_45134);
or U47684 (N_47684,N_44141,N_45078);
or U47685 (N_47685,N_45256,N_44555);
or U47686 (N_47686,N_45522,N_44606);
and U47687 (N_47687,N_45867,N_44283);
and U47688 (N_47688,N_44342,N_45155);
xor U47689 (N_47689,N_45544,N_44308);
nor U47690 (N_47690,N_45640,N_45135);
and U47691 (N_47691,N_45577,N_44177);
nand U47692 (N_47692,N_44034,N_45153);
nor U47693 (N_47693,N_44238,N_44339);
nand U47694 (N_47694,N_45352,N_45721);
nand U47695 (N_47695,N_45303,N_44867);
nor U47696 (N_47696,N_44374,N_44935);
xnor U47697 (N_47697,N_44089,N_44276);
nand U47698 (N_47698,N_45060,N_44958);
or U47699 (N_47699,N_45410,N_44333);
and U47700 (N_47700,N_45963,N_44335);
nor U47701 (N_47701,N_45478,N_44878);
or U47702 (N_47702,N_44753,N_45448);
and U47703 (N_47703,N_45430,N_45622);
or U47704 (N_47704,N_44986,N_45655);
and U47705 (N_47705,N_44733,N_45593);
nand U47706 (N_47706,N_44972,N_44301);
or U47707 (N_47707,N_44810,N_44697);
nor U47708 (N_47708,N_45272,N_45399);
or U47709 (N_47709,N_44389,N_44815);
nand U47710 (N_47710,N_45883,N_44394);
xor U47711 (N_47711,N_45353,N_45793);
nand U47712 (N_47712,N_44964,N_44615);
nand U47713 (N_47713,N_45525,N_45819);
nand U47714 (N_47714,N_45756,N_44595);
xor U47715 (N_47715,N_45526,N_45739);
and U47716 (N_47716,N_45458,N_45447);
xor U47717 (N_47717,N_44309,N_44977);
nor U47718 (N_47718,N_44733,N_45708);
nor U47719 (N_47719,N_44861,N_44228);
nor U47720 (N_47720,N_44660,N_44254);
nor U47721 (N_47721,N_45018,N_45436);
xor U47722 (N_47722,N_44244,N_44280);
nor U47723 (N_47723,N_44605,N_45933);
and U47724 (N_47724,N_44247,N_44922);
nand U47725 (N_47725,N_44940,N_45258);
or U47726 (N_47726,N_45242,N_44453);
or U47727 (N_47727,N_45928,N_44173);
nor U47728 (N_47728,N_44215,N_44603);
or U47729 (N_47729,N_45349,N_44755);
nand U47730 (N_47730,N_44976,N_44210);
nor U47731 (N_47731,N_44918,N_45173);
nor U47732 (N_47732,N_44448,N_44583);
nor U47733 (N_47733,N_45807,N_45990);
xor U47734 (N_47734,N_45793,N_44511);
or U47735 (N_47735,N_44190,N_45393);
and U47736 (N_47736,N_44952,N_45450);
xnor U47737 (N_47737,N_44208,N_44025);
nand U47738 (N_47738,N_44009,N_45166);
and U47739 (N_47739,N_45310,N_44753);
nor U47740 (N_47740,N_44288,N_44370);
or U47741 (N_47741,N_45621,N_44382);
or U47742 (N_47742,N_45494,N_45431);
and U47743 (N_47743,N_45023,N_44126);
nor U47744 (N_47744,N_44614,N_45453);
nand U47745 (N_47745,N_44430,N_44495);
nor U47746 (N_47746,N_44641,N_45448);
xor U47747 (N_47747,N_45287,N_45856);
nor U47748 (N_47748,N_45656,N_45441);
nand U47749 (N_47749,N_44951,N_45862);
xor U47750 (N_47750,N_45580,N_44730);
and U47751 (N_47751,N_45377,N_44618);
or U47752 (N_47752,N_44139,N_44601);
nand U47753 (N_47753,N_45931,N_44540);
xor U47754 (N_47754,N_44474,N_44664);
xor U47755 (N_47755,N_44632,N_44565);
or U47756 (N_47756,N_45823,N_45043);
and U47757 (N_47757,N_44214,N_44869);
nand U47758 (N_47758,N_45505,N_45661);
nor U47759 (N_47759,N_45759,N_44264);
nor U47760 (N_47760,N_44408,N_45064);
xor U47761 (N_47761,N_44207,N_45552);
nor U47762 (N_47762,N_44805,N_44123);
or U47763 (N_47763,N_44503,N_45096);
xor U47764 (N_47764,N_44045,N_44620);
nor U47765 (N_47765,N_45920,N_44142);
and U47766 (N_47766,N_44055,N_45576);
nand U47767 (N_47767,N_44195,N_45053);
or U47768 (N_47768,N_45912,N_44128);
or U47769 (N_47769,N_44137,N_44714);
nor U47770 (N_47770,N_45844,N_45201);
or U47771 (N_47771,N_44150,N_44902);
nor U47772 (N_47772,N_45586,N_45200);
xnor U47773 (N_47773,N_44216,N_45347);
nand U47774 (N_47774,N_45177,N_45804);
xor U47775 (N_47775,N_44879,N_44765);
or U47776 (N_47776,N_45926,N_45715);
or U47777 (N_47777,N_45035,N_45606);
nor U47778 (N_47778,N_45470,N_45655);
xnor U47779 (N_47779,N_45174,N_44448);
and U47780 (N_47780,N_45943,N_44189);
xor U47781 (N_47781,N_44129,N_45145);
or U47782 (N_47782,N_45049,N_44260);
nor U47783 (N_47783,N_45348,N_44847);
and U47784 (N_47784,N_45474,N_45480);
nor U47785 (N_47785,N_45832,N_45600);
xnor U47786 (N_47786,N_44125,N_44604);
nor U47787 (N_47787,N_44501,N_45939);
nand U47788 (N_47788,N_44967,N_45050);
or U47789 (N_47789,N_45741,N_44740);
xor U47790 (N_47790,N_44159,N_44535);
and U47791 (N_47791,N_45651,N_45288);
or U47792 (N_47792,N_45088,N_45111);
or U47793 (N_47793,N_44247,N_45370);
and U47794 (N_47794,N_44764,N_45367);
and U47795 (N_47795,N_45052,N_45740);
or U47796 (N_47796,N_44821,N_44289);
nor U47797 (N_47797,N_45747,N_45392);
nand U47798 (N_47798,N_44429,N_45505);
and U47799 (N_47799,N_45305,N_44806);
nand U47800 (N_47800,N_45617,N_45644);
and U47801 (N_47801,N_44890,N_44604);
nor U47802 (N_47802,N_45214,N_44169);
and U47803 (N_47803,N_45541,N_44175);
nand U47804 (N_47804,N_44840,N_45701);
nor U47805 (N_47805,N_44550,N_45729);
nor U47806 (N_47806,N_45287,N_45076);
or U47807 (N_47807,N_45642,N_44663);
nand U47808 (N_47808,N_44083,N_44947);
xnor U47809 (N_47809,N_45061,N_44944);
nor U47810 (N_47810,N_44743,N_45462);
and U47811 (N_47811,N_44764,N_44886);
and U47812 (N_47812,N_45755,N_44224);
nand U47813 (N_47813,N_45356,N_45321);
nor U47814 (N_47814,N_44235,N_45591);
nand U47815 (N_47815,N_44869,N_45156);
and U47816 (N_47816,N_45032,N_45343);
nand U47817 (N_47817,N_44612,N_45541);
or U47818 (N_47818,N_44115,N_44416);
xnor U47819 (N_47819,N_45565,N_44691);
nand U47820 (N_47820,N_45170,N_45761);
nand U47821 (N_47821,N_44516,N_45721);
and U47822 (N_47822,N_44046,N_45488);
and U47823 (N_47823,N_45018,N_44945);
or U47824 (N_47824,N_45091,N_44044);
and U47825 (N_47825,N_45583,N_44042);
nor U47826 (N_47826,N_44978,N_45927);
nand U47827 (N_47827,N_45166,N_44655);
nand U47828 (N_47828,N_44901,N_44725);
nor U47829 (N_47829,N_45513,N_45170);
or U47830 (N_47830,N_44824,N_44776);
or U47831 (N_47831,N_44392,N_45218);
xor U47832 (N_47832,N_45392,N_44588);
nand U47833 (N_47833,N_45542,N_44478);
xor U47834 (N_47834,N_44547,N_45125);
and U47835 (N_47835,N_45434,N_44939);
and U47836 (N_47836,N_44792,N_44096);
nor U47837 (N_47837,N_44379,N_44760);
nand U47838 (N_47838,N_44460,N_45469);
nor U47839 (N_47839,N_45676,N_44656);
and U47840 (N_47840,N_45310,N_45295);
xnor U47841 (N_47841,N_44337,N_45254);
nand U47842 (N_47842,N_45584,N_45312);
nand U47843 (N_47843,N_45820,N_44918);
and U47844 (N_47844,N_45046,N_44304);
xnor U47845 (N_47845,N_44270,N_45640);
nor U47846 (N_47846,N_44687,N_44414);
and U47847 (N_47847,N_45972,N_44328);
or U47848 (N_47848,N_45158,N_45869);
xnor U47849 (N_47849,N_45118,N_44050);
and U47850 (N_47850,N_45290,N_45442);
or U47851 (N_47851,N_45502,N_45180);
and U47852 (N_47852,N_45284,N_45514);
nor U47853 (N_47853,N_44237,N_44555);
nor U47854 (N_47854,N_45732,N_45580);
xor U47855 (N_47855,N_44886,N_44871);
nand U47856 (N_47856,N_45167,N_44242);
nand U47857 (N_47857,N_44236,N_45143);
nand U47858 (N_47858,N_45185,N_44000);
or U47859 (N_47859,N_44043,N_44412);
and U47860 (N_47860,N_45302,N_45642);
xor U47861 (N_47861,N_45844,N_45100);
xnor U47862 (N_47862,N_44111,N_44409);
or U47863 (N_47863,N_44992,N_44430);
nor U47864 (N_47864,N_45969,N_44381);
xor U47865 (N_47865,N_45749,N_44613);
nor U47866 (N_47866,N_44386,N_45314);
nand U47867 (N_47867,N_44520,N_44763);
xor U47868 (N_47868,N_45712,N_44680);
xnor U47869 (N_47869,N_44486,N_44833);
and U47870 (N_47870,N_44075,N_44682);
or U47871 (N_47871,N_45121,N_45103);
nor U47872 (N_47872,N_44704,N_45847);
nand U47873 (N_47873,N_45857,N_44443);
or U47874 (N_47874,N_45628,N_45350);
and U47875 (N_47875,N_45839,N_44732);
and U47876 (N_47876,N_44047,N_44117);
and U47877 (N_47877,N_45423,N_45258);
nor U47878 (N_47878,N_44962,N_45869);
and U47879 (N_47879,N_44221,N_44288);
and U47880 (N_47880,N_44398,N_45037);
and U47881 (N_47881,N_44154,N_44196);
or U47882 (N_47882,N_44301,N_45025);
and U47883 (N_47883,N_44756,N_44654);
or U47884 (N_47884,N_45979,N_45665);
nor U47885 (N_47885,N_44635,N_44064);
xor U47886 (N_47886,N_45085,N_45916);
or U47887 (N_47887,N_44517,N_44359);
and U47888 (N_47888,N_44064,N_45150);
or U47889 (N_47889,N_45994,N_44362);
and U47890 (N_47890,N_44481,N_44122);
or U47891 (N_47891,N_44824,N_45654);
nor U47892 (N_47892,N_45956,N_44075);
nand U47893 (N_47893,N_45651,N_45106);
xnor U47894 (N_47894,N_45436,N_45875);
xnor U47895 (N_47895,N_45153,N_44305);
nand U47896 (N_47896,N_45128,N_44681);
xor U47897 (N_47897,N_45788,N_44473);
and U47898 (N_47898,N_45246,N_44820);
and U47899 (N_47899,N_44973,N_44797);
and U47900 (N_47900,N_44972,N_45211);
nor U47901 (N_47901,N_45391,N_44818);
or U47902 (N_47902,N_45962,N_45920);
nor U47903 (N_47903,N_44784,N_45496);
nand U47904 (N_47904,N_44738,N_44112);
or U47905 (N_47905,N_44875,N_45342);
and U47906 (N_47906,N_44266,N_44552);
nand U47907 (N_47907,N_45986,N_44283);
or U47908 (N_47908,N_44032,N_44726);
or U47909 (N_47909,N_45121,N_44412);
or U47910 (N_47910,N_45925,N_44348);
or U47911 (N_47911,N_44293,N_44939);
nor U47912 (N_47912,N_45810,N_45107);
xor U47913 (N_47913,N_45288,N_45116);
nand U47914 (N_47914,N_44218,N_45659);
nor U47915 (N_47915,N_45607,N_45154);
and U47916 (N_47916,N_45731,N_45694);
xor U47917 (N_47917,N_45633,N_45052);
xor U47918 (N_47918,N_45704,N_44279);
nand U47919 (N_47919,N_44655,N_45102);
nor U47920 (N_47920,N_44868,N_44817);
nor U47921 (N_47921,N_44032,N_45369);
nand U47922 (N_47922,N_45154,N_44635);
xor U47923 (N_47923,N_45736,N_44220);
or U47924 (N_47924,N_45499,N_44511);
nor U47925 (N_47925,N_44195,N_45279);
nor U47926 (N_47926,N_45297,N_44540);
or U47927 (N_47927,N_44111,N_44065);
or U47928 (N_47928,N_44427,N_45536);
or U47929 (N_47929,N_44268,N_45626);
and U47930 (N_47930,N_45041,N_45696);
or U47931 (N_47931,N_44306,N_45640);
and U47932 (N_47932,N_44467,N_45972);
nor U47933 (N_47933,N_44140,N_45152);
or U47934 (N_47934,N_44386,N_44792);
xor U47935 (N_47935,N_45611,N_44805);
xnor U47936 (N_47936,N_44191,N_45268);
or U47937 (N_47937,N_45757,N_44915);
and U47938 (N_47938,N_44778,N_45295);
and U47939 (N_47939,N_44278,N_44105);
nor U47940 (N_47940,N_44459,N_45614);
xor U47941 (N_47941,N_45769,N_44360);
or U47942 (N_47942,N_44230,N_44363);
and U47943 (N_47943,N_44532,N_44192);
nand U47944 (N_47944,N_45534,N_44731);
xor U47945 (N_47945,N_44472,N_44648);
nor U47946 (N_47946,N_45926,N_45160);
nor U47947 (N_47947,N_44511,N_45601);
nor U47948 (N_47948,N_45132,N_45834);
xnor U47949 (N_47949,N_44541,N_44275);
nor U47950 (N_47950,N_44835,N_44323);
and U47951 (N_47951,N_44673,N_45215);
xnor U47952 (N_47952,N_44178,N_45811);
nand U47953 (N_47953,N_45085,N_45785);
or U47954 (N_47954,N_45812,N_45485);
nor U47955 (N_47955,N_45366,N_45477);
or U47956 (N_47956,N_44972,N_45476);
xnor U47957 (N_47957,N_45602,N_45114);
nor U47958 (N_47958,N_45856,N_44535);
xor U47959 (N_47959,N_45842,N_45105);
xor U47960 (N_47960,N_44407,N_44630);
nor U47961 (N_47961,N_44479,N_45603);
or U47962 (N_47962,N_44619,N_44412);
or U47963 (N_47963,N_45090,N_45680);
or U47964 (N_47964,N_45828,N_44110);
or U47965 (N_47965,N_44458,N_45684);
and U47966 (N_47966,N_45106,N_44434);
xnor U47967 (N_47967,N_44019,N_45742);
or U47968 (N_47968,N_44846,N_45274);
xnor U47969 (N_47969,N_44294,N_45228);
and U47970 (N_47970,N_45237,N_45417);
nand U47971 (N_47971,N_44555,N_44841);
and U47972 (N_47972,N_44478,N_45689);
and U47973 (N_47973,N_45860,N_44702);
nand U47974 (N_47974,N_44423,N_44244);
nor U47975 (N_47975,N_44024,N_44740);
nor U47976 (N_47976,N_45441,N_44749);
xnor U47977 (N_47977,N_45900,N_44895);
nor U47978 (N_47978,N_45214,N_44899);
nand U47979 (N_47979,N_44236,N_45347);
nor U47980 (N_47980,N_45827,N_44728);
nand U47981 (N_47981,N_45734,N_45200);
nand U47982 (N_47982,N_44933,N_44132);
and U47983 (N_47983,N_45030,N_44402);
nand U47984 (N_47984,N_44146,N_44958);
nand U47985 (N_47985,N_45202,N_45192);
nand U47986 (N_47986,N_44075,N_44892);
or U47987 (N_47987,N_44487,N_45393);
nand U47988 (N_47988,N_45157,N_44209);
or U47989 (N_47989,N_44519,N_44559);
nand U47990 (N_47990,N_45862,N_45290);
or U47991 (N_47991,N_44165,N_45049);
and U47992 (N_47992,N_44236,N_45951);
xor U47993 (N_47993,N_44123,N_44702);
nand U47994 (N_47994,N_45253,N_45939);
or U47995 (N_47995,N_44204,N_45814);
xor U47996 (N_47996,N_44168,N_45584);
or U47997 (N_47997,N_45398,N_44576);
or U47998 (N_47998,N_44118,N_45660);
or U47999 (N_47999,N_44163,N_44562);
xor U48000 (N_48000,N_46149,N_47317);
nand U48001 (N_48001,N_47533,N_47682);
and U48002 (N_48002,N_47426,N_46958);
or U48003 (N_48003,N_47824,N_47852);
and U48004 (N_48004,N_47540,N_46131);
or U48005 (N_48005,N_47982,N_46936);
and U48006 (N_48006,N_46431,N_47470);
nand U48007 (N_48007,N_46946,N_46109);
nand U48008 (N_48008,N_46278,N_46274);
nor U48009 (N_48009,N_46897,N_46286);
xnor U48010 (N_48010,N_46712,N_46486);
or U48011 (N_48011,N_46208,N_47198);
and U48012 (N_48012,N_46056,N_46942);
nand U48013 (N_48013,N_47603,N_46061);
xor U48014 (N_48014,N_46226,N_46156);
and U48015 (N_48015,N_47397,N_47525);
or U48016 (N_48016,N_46643,N_47559);
nand U48017 (N_48017,N_47891,N_47574);
nor U48018 (N_48018,N_47339,N_46285);
nor U48019 (N_48019,N_47671,N_47674);
and U48020 (N_48020,N_47965,N_46784);
and U48021 (N_48021,N_47335,N_46080);
nor U48022 (N_48022,N_47362,N_46279);
xor U48023 (N_48023,N_46573,N_46235);
nor U48024 (N_48024,N_47940,N_46395);
xor U48025 (N_48025,N_46619,N_46141);
and U48026 (N_48026,N_46657,N_47732);
or U48027 (N_48027,N_47528,N_46821);
or U48028 (N_48028,N_46336,N_47399);
or U48029 (N_48029,N_46353,N_47132);
nor U48030 (N_48030,N_47589,N_46242);
xor U48031 (N_48031,N_46847,N_46763);
xor U48032 (N_48032,N_47214,N_47297);
nor U48033 (N_48033,N_47127,N_47762);
nand U48034 (N_48034,N_47223,N_46802);
xnor U48035 (N_48035,N_47555,N_46114);
or U48036 (N_48036,N_47867,N_46315);
or U48037 (N_48037,N_46751,N_47471);
nor U48038 (N_48038,N_47462,N_47913);
and U48039 (N_48039,N_46685,N_46715);
nand U48040 (N_48040,N_46995,N_47429);
xnor U48041 (N_48041,N_47286,N_46369);
and U48042 (N_48042,N_47902,N_46649);
xnor U48043 (N_48043,N_46566,N_46009);
nand U48044 (N_48044,N_46373,N_46873);
and U48045 (N_48045,N_46005,N_47669);
xor U48046 (N_48046,N_47253,N_46391);
xor U48047 (N_48047,N_46684,N_46010);
or U48048 (N_48048,N_47222,N_47738);
and U48049 (N_48049,N_47787,N_46406);
nor U48050 (N_48050,N_47615,N_47323);
xnor U48051 (N_48051,N_47013,N_47600);
nor U48052 (N_48052,N_47308,N_47990);
nor U48053 (N_48053,N_47404,N_47702);
and U48054 (N_48054,N_46551,N_47206);
xnor U48055 (N_48055,N_46927,N_47376);
nor U48056 (N_48056,N_47654,N_46179);
and U48057 (N_48057,N_47751,N_46600);
xnor U48058 (N_48058,N_47455,N_46744);
and U48059 (N_48059,N_46256,N_47623);
nor U48060 (N_48060,N_47507,N_46337);
or U48061 (N_48061,N_47854,N_47861);
nand U48062 (N_48062,N_47766,N_47349);
nand U48063 (N_48063,N_46941,N_46667);
nor U48064 (N_48064,N_47184,N_47529);
xnor U48065 (N_48065,N_46713,N_47642);
xnor U48066 (N_48066,N_46289,N_47120);
xor U48067 (N_48067,N_46961,N_47084);
xor U48068 (N_48068,N_46819,N_47964);
or U48069 (N_48069,N_47065,N_47107);
xor U48070 (N_48070,N_46525,N_46546);
xor U48071 (N_48071,N_47128,N_47703);
and U48072 (N_48072,N_46025,N_47234);
and U48073 (N_48073,N_46326,N_46816);
or U48074 (N_48074,N_46264,N_47432);
nand U48075 (N_48075,N_46970,N_47450);
and U48076 (N_48076,N_47488,N_47826);
and U48077 (N_48077,N_47262,N_47465);
and U48078 (N_48078,N_46664,N_46119);
nand U48079 (N_48079,N_47845,N_47409);
nor U48080 (N_48080,N_46872,N_46000);
or U48081 (N_48081,N_46298,N_47447);
xor U48082 (N_48082,N_46929,N_46008);
nor U48083 (N_48083,N_47009,N_46268);
and U48084 (N_48084,N_47320,N_47698);
and U48085 (N_48085,N_47236,N_47496);
nand U48086 (N_48086,N_47866,N_46940);
and U48087 (N_48087,N_46676,N_46645);
xor U48088 (N_48088,N_47730,N_46169);
xnor U48089 (N_48089,N_47140,N_47176);
nand U48090 (N_48090,N_47242,N_47341);
xor U48091 (N_48091,N_46201,N_47967);
and U48092 (N_48092,N_46239,N_47293);
and U48093 (N_48093,N_46213,N_46878);
or U48094 (N_48094,N_46794,N_47494);
nand U48095 (N_48095,N_47984,N_47799);
nor U48096 (N_48096,N_47464,N_47553);
nand U48097 (N_48097,N_46560,N_47241);
and U48098 (N_48098,N_46194,N_47933);
nand U48099 (N_48099,N_47680,N_46624);
and U48100 (N_48100,N_46252,N_47343);
xnor U48101 (N_48101,N_47576,N_46734);
or U48102 (N_48102,N_46209,N_46185);
nor U48103 (N_48103,N_47405,N_47472);
xor U48104 (N_48104,N_47060,N_46582);
nand U48105 (N_48105,N_47029,N_46233);
nor U48106 (N_48106,N_46294,N_47749);
nand U48107 (N_48107,N_46426,N_47452);
and U48108 (N_48108,N_47484,N_47015);
nor U48109 (N_48109,N_47584,N_46276);
xnor U48110 (N_48110,N_46089,N_47103);
nand U48111 (N_48111,N_47192,N_47633);
nand U48112 (N_48112,N_46133,N_46272);
and U48113 (N_48113,N_47023,N_46764);
or U48114 (N_48114,N_47769,N_47461);
xor U48115 (N_48115,N_47081,N_46104);
and U48116 (N_48116,N_46701,N_47147);
and U48117 (N_48117,N_47263,N_47713);
nor U48118 (N_48118,N_47044,N_47071);
and U48119 (N_48119,N_46693,N_47728);
or U48120 (N_48120,N_47768,N_46898);
or U48121 (N_48121,N_47003,N_46521);
and U48122 (N_48122,N_47827,N_46586);
or U48123 (N_48123,N_47934,N_47284);
and U48124 (N_48124,N_46911,N_46733);
nand U48125 (N_48125,N_47275,N_46505);
nand U48126 (N_48126,N_47058,N_47538);
nand U48127 (N_48127,N_47955,N_46162);
or U48128 (N_48128,N_46524,N_47704);
or U48129 (N_48129,N_46792,N_46931);
nor U48130 (N_48130,N_47304,N_47428);
nor U48131 (N_48131,N_46223,N_47947);
nand U48132 (N_48132,N_46519,N_47066);
nand U48133 (N_48133,N_47314,N_46504);
nor U48134 (N_48134,N_47620,N_47853);
or U48135 (N_48135,N_47252,N_47425);
xnor U48136 (N_48136,N_47739,N_47996);
nor U48137 (N_48137,N_47594,N_47387);
and U48138 (N_48138,N_46583,N_46771);
nor U48139 (N_48139,N_47232,N_47788);
or U48140 (N_48140,N_46402,N_46983);
nor U48141 (N_48141,N_47067,N_47267);
and U48142 (N_48142,N_46992,N_47761);
nand U48143 (N_48143,N_46532,N_46158);
nand U48144 (N_48144,N_47613,N_46774);
xnor U48145 (N_48145,N_47268,N_46606);
nor U48146 (N_48146,N_47477,N_47005);
and U48147 (N_48147,N_46815,N_46448);
nand U48148 (N_48148,N_47256,N_46623);
xnor U48149 (N_48149,N_47634,N_47040);
xnor U48150 (N_48150,N_47298,N_47229);
xnor U48151 (N_48151,N_46168,N_46167);
or U48152 (N_48152,N_47294,N_47281);
nand U48153 (N_48153,N_46053,N_47356);
nor U48154 (N_48154,N_47032,N_46066);
or U48155 (N_48155,N_47554,N_47161);
nand U48156 (N_48156,N_46218,N_47331);
nand U48157 (N_48157,N_47312,N_47403);
nand U48158 (N_48158,N_46430,N_46500);
nand U48159 (N_48159,N_47817,N_46030);
xnor U48160 (N_48160,N_46248,N_46175);
xor U48161 (N_48161,N_46522,N_46882);
nand U48162 (N_48162,N_46097,N_46446);
xor U48163 (N_48163,N_47953,N_47687);
nor U48164 (N_48164,N_46984,N_46379);
and U48165 (N_48165,N_47750,N_47959);
and U48166 (N_48166,N_47802,N_46189);
nor U48167 (N_48167,N_47441,N_47686);
nand U48168 (N_48168,N_47381,N_47001);
and U48169 (N_48169,N_46367,N_46830);
and U48170 (N_48170,N_46536,N_47338);
nor U48171 (N_48171,N_47099,N_46967);
xnor U48172 (N_48172,N_47608,N_46644);
xor U48173 (N_48173,N_47460,N_47763);
or U48174 (N_48174,N_46765,N_46266);
nor U48175 (N_48175,N_46717,N_47083);
xor U48176 (N_48176,N_47150,N_47621);
nor U48177 (N_48177,N_47135,N_47487);
xnor U48178 (N_48178,N_47021,N_46745);
xnor U48179 (N_48179,N_47875,N_47547);
nor U48180 (N_48180,N_46543,N_47243);
and U48181 (N_48181,N_47193,N_47577);
or U48182 (N_48182,N_47927,N_47166);
xnor U48183 (N_48183,N_46043,N_47882);
nand U48184 (N_48184,N_47438,N_46981);
and U48185 (N_48185,N_46442,N_47264);
xnor U48186 (N_48186,N_46051,N_47718);
nand U48187 (N_48187,N_46420,N_47524);
nand U48188 (N_48188,N_47442,N_47870);
nand U48189 (N_48189,N_46232,N_47998);
or U48190 (N_48190,N_47857,N_46605);
and U48191 (N_48191,N_46885,N_46640);
nand U48192 (N_48192,N_46956,N_47911);
nor U48193 (N_48193,N_47435,N_46265);
xnor U48194 (N_48194,N_46799,N_47086);
xor U48195 (N_48195,N_46952,N_46359);
or U48196 (N_48196,N_47725,N_46325);
and U48197 (N_48197,N_47693,N_46258);
and U48198 (N_48198,N_47110,N_46107);
xnor U48199 (N_48199,N_47808,N_46128);
nand U48200 (N_48200,N_47195,N_46140);
and U48201 (N_48201,N_47138,N_47564);
nand U48202 (N_48202,N_47624,N_46318);
nand U48203 (N_48203,N_46028,N_46464);
nor U48204 (N_48204,N_46953,N_46074);
nor U48205 (N_48205,N_47890,N_47893);
and U48206 (N_48206,N_47042,N_46598);
nor U48207 (N_48207,N_47119,N_47977);
and U48208 (N_48208,N_46165,N_47935);
and U48209 (N_48209,N_47586,N_46388);
or U48210 (N_48210,N_47420,N_46916);
and U48211 (N_48211,N_47770,N_47760);
nor U48212 (N_48212,N_47720,N_47638);
nor U48213 (N_48213,N_47944,N_47324);
nand U48214 (N_48214,N_47115,N_47412);
xor U48215 (N_48215,N_47434,N_47892);
xor U48216 (N_48216,N_46636,N_47492);
nor U48217 (N_48217,N_46578,N_46806);
nor U48218 (N_48218,N_46839,N_47809);
nand U48219 (N_48219,N_46782,N_47345);
or U48220 (N_48220,N_46033,N_46793);
and U48221 (N_48221,N_46204,N_46400);
xnor U48222 (N_48222,N_46416,N_47661);
nand U48223 (N_48223,N_46835,N_46300);
xor U48224 (N_48224,N_47024,N_47048);
nor U48225 (N_48225,N_47102,N_47868);
xnor U48226 (N_48226,N_46572,N_47677);
or U48227 (N_48227,N_47748,N_47351);
and U48228 (N_48228,N_47203,N_47796);
nand U48229 (N_48229,N_47658,N_47532);
or U48230 (N_48230,N_47869,N_47105);
and U48231 (N_48231,N_46018,N_47018);
nor U48232 (N_48232,N_47392,N_46236);
nor U48233 (N_48233,N_46454,N_46186);
nand U48234 (N_48234,N_46243,N_47148);
and U48235 (N_48235,N_46432,N_46562);
xnor U48236 (N_48236,N_47122,N_47061);
nand U48237 (N_48237,N_46284,N_46498);
nand U48238 (N_48238,N_47276,N_46377);
or U48239 (N_48239,N_47963,N_47273);
xor U48240 (N_48240,N_47966,N_47475);
and U48241 (N_48241,N_46100,N_47563);
nand U48242 (N_48242,N_46917,N_47847);
and U48243 (N_48243,N_47142,N_46758);
nor U48244 (N_48244,N_47172,N_46251);
nor U48245 (N_48245,N_46328,N_46138);
and U48246 (N_48246,N_47567,N_46621);
and U48247 (N_48247,N_46852,N_47446);
nand U48248 (N_48248,N_46081,N_47958);
xnor U48249 (N_48249,N_47792,N_47517);
or U48250 (N_48250,N_46125,N_46151);
or U48251 (N_48251,N_47910,N_46260);
nor U48252 (N_48252,N_46220,N_46665);
nand U48253 (N_48253,N_47520,N_46646);
or U48254 (N_48254,N_46057,N_47419);
nand U48255 (N_48255,N_47188,N_47579);
nor U48256 (N_48256,N_47781,N_47043);
nor U48257 (N_48257,N_46212,N_47280);
nor U48258 (N_48258,N_46293,N_46727);
nand U48259 (N_48259,N_47975,N_47137);
nor U48260 (N_48260,N_46322,N_47437);
and U48261 (N_48261,N_47512,N_46688);
nand U48262 (N_48262,N_47016,N_46316);
and U48263 (N_48263,N_46569,N_46820);
nand U48264 (N_48264,N_47415,N_46738);
xnor U48265 (N_48265,N_46216,N_46062);
or U48266 (N_48266,N_46357,N_46973);
xor U48267 (N_48267,N_47812,N_47290);
xor U48268 (N_48268,N_46867,N_46964);
and U48269 (N_48269,N_46237,N_47622);
and U48270 (N_48270,N_46622,N_46153);
nor U48271 (N_48271,N_46085,N_47591);
nor U48272 (N_48272,N_46540,N_47053);
xnor U48273 (N_48273,N_47519,N_47939);
nor U48274 (N_48274,N_46050,N_46036);
nand U48275 (N_48275,N_46451,N_47816);
or U48276 (N_48276,N_47443,N_47948);
nand U48277 (N_48277,N_47557,N_47696);
xnor U48278 (N_48278,N_46843,N_46585);
nor U48279 (N_48279,N_47932,N_47235);
and U48280 (N_48280,N_46881,N_47736);
nand U48281 (N_48281,N_46960,N_47509);
xor U48282 (N_48282,N_46122,N_47803);
and U48283 (N_48283,N_46689,N_47333);
or U48284 (N_48284,N_47480,N_47052);
nor U48285 (N_48285,N_47466,N_46205);
and U48286 (N_48286,N_46732,N_46393);
or U48287 (N_48287,N_46283,N_47375);
nor U48288 (N_48288,N_46642,N_47012);
nor U48289 (N_48289,N_46273,N_47271);
or U48290 (N_48290,N_46674,N_47406);
xnor U48291 (N_48291,N_46512,N_46360);
nand U48292 (N_48292,N_46550,N_46297);
or U48293 (N_48293,N_46335,N_46989);
nor U48294 (N_48294,N_46575,N_47772);
nor U48295 (N_48295,N_46980,N_46307);
and U48296 (N_48296,N_47237,N_47900);
nor U48297 (N_48297,N_46726,N_46737);
nor U48298 (N_48298,N_47800,N_46375);
xor U48299 (N_48299,N_47095,N_46113);
and U48300 (N_48300,N_46945,N_46574);
xnor U48301 (N_48301,N_47082,N_47248);
and U48302 (N_48302,N_46392,N_47898);
nor U48303 (N_48303,N_47660,N_46925);
and U48304 (N_48304,N_47597,N_47031);
xor U48305 (N_48305,N_46757,N_46708);
xnor U48306 (N_48306,N_46846,N_47240);
nor U48307 (N_48307,N_46382,N_47499);
and U48308 (N_48308,N_47549,N_46553);
and U48309 (N_48309,N_47636,N_47478);
xor U48310 (N_48310,N_47265,N_46954);
nor U48311 (N_48311,N_47929,N_47169);
nor U48312 (N_48312,N_47836,N_47778);
nand U48313 (N_48313,N_47108,N_47578);
nand U48314 (N_48314,N_47740,N_47617);
nand U48315 (N_48315,N_46506,N_46091);
xnor U48316 (N_48316,N_47605,N_46760);
nor U48317 (N_48317,N_47019,N_46513);
nand U48318 (N_48318,N_46035,N_46919);
xor U48319 (N_48319,N_47296,N_46245);
nor U48320 (N_48320,N_46673,N_47684);
nor U48321 (N_48321,N_47651,N_47077);
nor U48322 (N_48322,N_46417,N_47261);
nor U48323 (N_48323,N_46497,N_47628);
and U48324 (N_48324,N_46652,N_46714);
or U48325 (N_48325,N_47092,N_46705);
and U48326 (N_48326,N_46761,N_47350);
or U48327 (N_48327,N_47346,N_47491);
nor U48328 (N_48328,N_46786,N_46287);
nor U48329 (N_48329,N_46604,N_47228);
or U48330 (N_48330,N_47552,N_47080);
nor U48331 (N_48331,N_47655,N_46282);
xor U48332 (N_48332,N_46001,N_46059);
nor U48333 (N_48333,N_47175,N_46955);
or U48334 (N_48334,N_47546,N_46127);
xor U48335 (N_48335,N_46824,N_46399);
and U48336 (N_48336,N_46440,N_47136);
xnor U48337 (N_48337,N_47220,N_46317);
and U48338 (N_48338,N_46034,N_46154);
nor U48339 (N_48339,N_47199,N_47954);
or U48340 (N_48340,N_46538,N_46148);
nor U48341 (N_48341,N_46889,N_47451);
xnor U48342 (N_48342,N_47377,N_46858);
and U48343 (N_48343,N_47151,N_46221);
nand U48344 (N_48344,N_47683,N_46988);
and U48345 (N_48345,N_47771,N_46343);
nand U48346 (N_48346,N_46719,N_46002);
xor U48347 (N_48347,N_47970,N_46787);
and U48348 (N_48348,N_47697,N_47074);
or U48349 (N_48349,N_46421,N_47431);
nor U48350 (N_48350,N_46775,N_47689);
xnor U48351 (N_48351,N_47146,N_46129);
xor U48352 (N_48352,N_47112,N_47194);
nor U48353 (N_48353,N_46290,N_46742);
xnor U48354 (N_48354,N_46135,N_47316);
or U48355 (N_48355,N_47530,N_46249);
and U48356 (N_48356,N_47908,N_47598);
nand U48357 (N_48357,N_46770,N_46837);
and U48358 (N_48358,N_46172,N_47968);
xnor U48359 (N_48359,N_46704,N_47340);
xor U48360 (N_48360,N_46874,N_46374);
nor U48361 (N_48361,N_47522,N_46038);
nor U48362 (N_48362,N_47389,N_47145);
nand U48363 (N_48363,N_47550,N_46994);
nor U48364 (N_48364,N_47291,N_46262);
and U48365 (N_48365,N_46990,N_46703);
nor U48366 (N_48366,N_47513,N_47495);
xnor U48367 (N_48367,N_46511,N_47486);
nor U48368 (N_48368,N_47079,N_47879);
nor U48369 (N_48369,N_47498,N_47794);
and U48370 (N_48370,N_46996,N_46174);
or U48371 (N_48371,N_46594,N_46354);
and U48372 (N_48372,N_47611,N_46414);
nor U48373 (N_48373,N_47418,N_47154);
and U48374 (N_48374,N_46428,N_47274);
nor U48375 (N_48375,N_46422,N_46031);
nand U48376 (N_48376,N_46870,N_46480);
xor U48377 (N_48377,N_46492,N_47855);
xor U48378 (N_48378,N_46338,N_46581);
or U48379 (N_48379,N_47444,N_47640);
xnor U48380 (N_48380,N_46344,N_47657);
nor U48381 (N_48381,N_46052,N_46230);
nand U48382 (N_48382,N_46444,N_46320);
nand U48383 (N_48383,N_46231,N_47037);
nand U48384 (N_48384,N_46020,N_47733);
xnor U48385 (N_48385,N_47159,N_47117);
and U48386 (N_48386,N_47871,N_47779);
and U48387 (N_48387,N_46831,N_46333);
or U48388 (N_48388,N_46781,N_47695);
and U48389 (N_48389,N_47832,N_47485);
nor U48390 (N_48390,N_47279,N_47489);
nor U48391 (N_48391,N_47822,N_46501);
nand U48392 (N_48392,N_47059,N_47459);
and U48393 (N_48393,N_47991,N_47363);
and U48394 (N_48394,N_46396,N_47215);
or U48395 (N_48395,N_47997,N_46634);
or U48396 (N_48396,N_47601,N_47407);
xor U48397 (N_48397,N_47886,N_47722);
or U48398 (N_48398,N_47413,N_47301);
or U48399 (N_48399,N_47219,N_46670);
nand U48400 (N_48400,N_47244,N_47789);
nand U48401 (N_48401,N_46556,N_47197);
nor U48402 (N_48402,N_47925,N_47260);
nor U48403 (N_48403,N_47508,N_46804);
nand U48404 (N_48404,N_46969,N_46707);
and U48405 (N_48405,N_46101,N_47731);
and U48406 (N_48406,N_47978,N_47098);
nor U48407 (N_48407,N_47878,N_47500);
or U48408 (N_48408,N_47008,N_46656);
and U48409 (N_48409,N_47208,N_46507);
and U48410 (N_48410,N_47224,N_47833);
nor U48411 (N_48411,N_47510,N_46669);
nand U48412 (N_48412,N_46329,N_47726);
xnor U48413 (N_48413,N_47211,N_47795);
nor U48414 (N_48414,N_47034,N_46476);
or U48415 (N_48415,N_46084,N_46601);
xor U48416 (N_48416,N_47473,N_46099);
and U48417 (N_48417,N_46384,N_47665);
nand U48418 (N_48418,N_46588,N_47957);
and U48419 (N_48419,N_46222,N_47479);
nand U48420 (N_48420,N_47300,N_47742);
nand U48421 (N_48421,N_47004,N_47883);
and U48422 (N_48422,N_47468,N_46876);
nor U48423 (N_48423,N_46437,N_47850);
or U48424 (N_48424,N_46895,N_46219);
xor U48425 (N_48425,N_47337,N_46177);
nand U48426 (N_48426,N_46527,N_47179);
and U48427 (N_48427,N_46675,N_47398);
nand U48428 (N_48428,N_46557,N_47659);
and U48429 (N_48429,N_46938,N_46609);
and U48430 (N_48430,N_46016,N_47126);
or U48431 (N_48431,N_46880,N_46901);
nor U48432 (N_48432,N_47889,N_46577);
xnor U48433 (N_48433,N_46853,N_47164);
nand U48434 (N_48434,N_47656,N_47181);
or U48435 (N_48435,N_47097,N_46661);
or U48436 (N_48436,N_46072,N_47952);
xnor U48437 (N_48437,N_47503,N_47070);
or U48438 (N_48438,N_46635,N_47125);
and U48439 (N_48439,N_46592,N_46612);
xor U48440 (N_48440,N_47445,N_47851);
and U48441 (N_48441,N_46436,N_46241);
and U48442 (N_48442,N_46533,N_47129);
nor U48443 (N_48443,N_47453,N_46544);
nand U48444 (N_48444,N_47033,N_47299);
or U48445 (N_48445,N_46397,N_46514);
nor U48446 (N_48446,N_47028,N_47254);
and U48447 (N_48447,N_47049,N_46461);
nand U48448 (N_48448,N_47705,N_46568);
and U48449 (N_48449,N_46349,N_47675);
xor U48450 (N_48450,N_47226,N_47999);
xnor U48451 (N_48451,N_47385,N_46425);
xor U48452 (N_48452,N_46735,N_47329);
or U48453 (N_48453,N_47873,N_46494);
nor U48454 (N_48454,N_47165,N_46968);
nand U48455 (N_48455,N_46766,N_47541);
and U48456 (N_48456,N_47629,N_46370);
or U48457 (N_48457,N_46173,N_46007);
nor U48458 (N_48458,N_47950,N_47745);
nor U48459 (N_48459,N_47956,N_46342);
nand U48460 (N_48460,N_46229,N_47050);
and U48461 (N_48461,N_46918,N_47637);
xnor U48462 (N_48462,N_46462,N_46844);
nand U48463 (N_48463,N_47690,N_46796);
nand U48464 (N_48464,N_46810,N_46313);
xnor U48465 (N_48465,N_46608,N_47765);
xnor U48466 (N_48466,N_47251,N_46126);
xor U48467 (N_48467,N_46227,N_46848);
and U48468 (N_48468,N_46418,N_47414);
or U48469 (N_48469,N_47724,N_47257);
or U48470 (N_48470,N_47653,N_46679);
xor U48471 (N_48471,N_47209,N_47283);
xor U48472 (N_48472,N_47884,N_47325);
or U48473 (N_48473,N_46206,N_46197);
nor U48474 (N_48474,N_47402,N_47839);
and U48475 (N_48475,N_47992,N_47318);
and U48476 (N_48476,N_47152,N_47831);
xnor U48477 (N_48477,N_46065,N_47862);
nor U48478 (N_48478,N_47834,N_46552);
or U48479 (N_48479,N_47786,N_46275);
nor U48480 (N_48480,N_46438,N_47588);
xnor U48481 (N_48481,N_47006,N_46681);
or U48482 (N_48482,N_47667,N_46121);
nor U48483 (N_48483,N_47109,N_46517);
nor U48484 (N_48484,N_47764,N_46170);
or U48485 (N_48485,N_47632,N_47924);
or U48486 (N_48486,N_46356,N_46306);
nand U48487 (N_48487,N_46999,N_46615);
nor U48488 (N_48488,N_47727,N_46654);
nor U48489 (N_48489,N_47210,N_46749);
xnor U48490 (N_48490,N_47828,N_47729);
and U48491 (N_48491,N_46523,N_46270);
and U48492 (N_48492,N_46372,N_47743);
nand U48493 (N_48493,N_47707,N_47545);
xnor U48494 (N_48494,N_46860,N_47838);
and U48495 (N_48495,N_47616,N_47051);
xor U48496 (N_48496,N_47526,N_47056);
or U48497 (N_48497,N_46259,N_46617);
nor U48498 (N_48498,N_47951,N_46628);
or U48499 (N_48499,N_47185,N_47604);
and U48500 (N_48500,N_46147,N_46934);
nand U48501 (N_48501,N_47319,N_46884);
and U48502 (N_48502,N_47481,N_47895);
and U48503 (N_48503,N_46027,N_46826);
nor U48504 (N_48504,N_46145,N_47100);
and U48505 (N_48505,N_46403,N_46817);
nor U48506 (N_48506,N_46639,N_46489);
and U48507 (N_48507,N_47981,N_46347);
and U48508 (N_48508,N_46415,N_47618);
nor U48509 (N_48509,N_47570,N_46026);
or U48510 (N_48510,N_47178,N_47189);
or U48511 (N_48511,N_47309,N_46836);
xnor U48512 (N_48512,N_46724,N_46073);
and U48513 (N_48513,N_47941,N_46312);
and U48514 (N_48514,N_46003,N_47183);
nor U48515 (N_48515,N_47785,N_46641);
and U48516 (N_48516,N_47609,N_46529);
nand U48517 (N_48517,N_46161,N_47639);
xnor U48518 (N_48518,N_46962,N_46214);
or U48519 (N_48519,N_46902,N_47942);
xnor U48520 (N_48520,N_47818,N_47711);
nand U48521 (N_48521,N_46750,N_46659);
xor U48522 (N_48522,N_46632,N_47245);
and U48523 (N_48523,N_46045,N_47133);
and U48524 (N_48524,N_46965,N_46467);
nor U48525 (N_48525,N_47502,N_47841);
nand U48526 (N_48526,N_46797,N_47646);
nor U48527 (N_48527,N_46134,N_46769);
and U48528 (N_48528,N_47780,N_46683);
xnor U48529 (N_48529,N_47233,N_46192);
and U48530 (N_48530,N_47390,N_47899);
nor U48531 (N_48531,N_46075,N_47672);
or U48532 (N_48532,N_46183,N_46244);
or U48533 (N_48533,N_47515,N_47255);
and U48534 (N_48534,N_47928,N_47272);
and U48535 (N_48535,N_47068,N_46160);
and U48536 (N_48536,N_47569,N_47170);
and U48537 (N_48537,N_46723,N_46380);
xor U48538 (N_48538,N_47162,N_46217);
nand U48539 (N_48539,N_47815,N_46651);
or U48540 (N_48540,N_47200,N_46845);
or U48541 (N_48541,N_47433,N_46710);
nand U48542 (N_48542,N_47221,N_46827);
or U48543 (N_48543,N_46697,N_47864);
and U48544 (N_48544,N_46638,N_46869);
nor U48545 (N_48545,N_47041,N_46663);
nor U48546 (N_48546,N_47747,N_46637);
and U48547 (N_48547,N_47355,N_47776);
nor U48548 (N_48548,N_46424,N_46103);
or U48549 (N_48549,N_46453,N_46579);
nand U48550 (N_48550,N_47000,N_46466);
xor U48551 (N_48551,N_46404,N_46120);
nor U48552 (N_48552,N_47313,N_47374);
or U48553 (N_48553,N_47790,N_46610);
nor U48554 (N_48554,N_46324,N_47302);
or U48555 (N_48555,N_46363,N_46894);
nand U48556 (N_48556,N_46423,N_47369);
xor U48557 (N_48557,N_47980,N_46408);
xnor U48558 (N_48558,N_46224,N_47535);
xnor U48559 (N_48559,N_47773,N_47055);
and U48560 (N_48560,N_47582,N_47571);
and U48561 (N_48561,N_47091,N_47880);
nand U48562 (N_48562,N_47627,N_46971);
or U48563 (N_48563,N_46042,N_46299);
nor U48564 (N_48564,N_46047,N_47993);
and U48565 (N_48565,N_46024,N_47840);
nand U48566 (N_48566,N_47511,N_47022);
nand U48567 (N_48567,N_47315,N_47612);
xnor U48568 (N_48568,N_47177,N_47038);
or U48569 (N_48569,N_46136,N_46439);
or U48570 (N_48570,N_46779,N_47946);
nand U48571 (N_48571,N_47664,N_46620);
nand U48572 (N_48572,N_46443,N_47116);
or U48573 (N_48573,N_47755,N_46875);
and U48574 (N_48574,N_47919,N_46459);
nor U48575 (N_48575,N_46152,N_46143);
or U48576 (N_48576,N_46288,N_46484);
xnor U48577 (N_48577,N_46250,N_46593);
or U48578 (N_48578,N_46441,N_47388);
xnor U48579 (N_48579,N_46032,N_47805);
nor U48580 (N_48580,N_46825,N_47625);
and U48581 (N_48581,N_46923,N_46090);
nand U48582 (N_48582,N_47463,N_47396);
or U48583 (N_48583,N_46914,N_46803);
nand U48584 (N_48584,N_47877,N_46851);
xor U48585 (N_48585,N_46111,N_46309);
xnor U48586 (N_48586,N_47843,N_47774);
nand U48587 (N_48587,N_47380,N_46920);
nor U48588 (N_48588,N_46747,N_47367);
nand U48589 (N_48589,N_47784,N_47506);
nand U48590 (N_48590,N_46928,N_46350);
nor U48591 (N_48591,N_46548,N_47187);
nor U48592 (N_48592,N_46469,N_46215);
or U48593 (N_48593,N_46362,N_47134);
xor U48594 (N_48594,N_46280,N_46974);
nand U48595 (N_48595,N_46132,N_46558);
or U48596 (N_48596,N_47130,N_46785);
nor U48597 (N_48597,N_46427,N_47849);
nor U48598 (N_48598,N_47332,N_46470);
nand U48599 (N_48599,N_47482,N_47157);
nand U48600 (N_48600,N_47035,N_47971);
or U48601 (N_48601,N_46716,N_46071);
nor U48602 (N_48602,N_47825,N_46691);
nand U48603 (N_48603,N_46741,N_46864);
or U48604 (N_48604,N_46323,N_47923);
nand U48605 (N_48605,N_47424,N_47906);
or U48606 (N_48606,N_46472,N_47876);
or U48607 (N_48607,N_46068,N_46531);
or U48608 (N_48608,N_46899,N_47094);
or U48609 (N_48609,N_46130,N_46800);
and U48610 (N_48610,N_47230,N_46096);
nand U48611 (N_48611,N_47912,N_47917);
nand U48612 (N_48612,N_47327,N_47701);
and U48613 (N_48613,N_46926,N_46662);
xnor U48614 (N_48614,N_47514,N_47218);
and U48615 (N_48615,N_46892,N_46181);
xor U48616 (N_48616,N_46891,N_46935);
nand U48617 (N_48617,N_46570,N_47057);
nor U48618 (N_48618,N_46626,N_46871);
or U48619 (N_48619,N_47539,N_46199);
or U48620 (N_48620,N_47737,N_46411);
or U48621 (N_48621,N_47078,N_46754);
and U48622 (N_48622,N_47644,N_46381);
xor U48623 (N_48623,N_46580,N_46371);
nor U48624 (N_48624,N_46255,N_46567);
xnor U48625 (N_48625,N_46238,N_46972);
xor U48626 (N_48626,N_46004,N_46813);
and U48627 (N_48627,N_46339,N_47562);
xnor U48628 (N_48628,N_47668,N_47681);
and U48629 (N_48629,N_47201,N_46576);
or U48630 (N_48630,N_46368,N_46178);
nor U48631 (N_48631,N_46093,N_47096);
xnor U48632 (N_48632,N_46904,N_47926);
or U48633 (N_48633,N_46296,N_47813);
or U48634 (N_48634,N_47143,N_46694);
nor U48635 (N_48635,N_47983,N_47174);
nand U48636 (N_48636,N_47101,N_47907);
nand U48637 (N_48637,N_46748,N_47587);
and U48638 (N_48638,N_46950,N_47692);
nand U48639 (N_48639,N_46412,N_47417);
nand U48640 (N_48640,N_46849,N_46937);
xor U48641 (N_48641,N_47814,N_46110);
xnor U48642 (N_48642,N_47217,N_46385);
or U48643 (N_48643,N_46908,N_46776);
nand U48644 (N_48644,N_47797,N_47026);
nand U48645 (N_48645,N_46355,N_47069);
nand U48646 (N_48646,N_47558,N_47989);
and U48647 (N_48647,N_47842,N_47699);
and U48648 (N_48648,N_46171,N_46795);
nor U48649 (N_48649,N_46678,N_46361);
nand U48650 (N_48650,N_47670,N_46040);
and U48651 (N_48651,N_46456,N_47918);
and U48652 (N_48652,N_47721,N_46660);
nand U48653 (N_48653,N_47897,N_47909);
or U48654 (N_48654,N_46041,N_47856);
or U48655 (N_48655,N_46473,N_46254);
xnor U48656 (N_48656,N_46458,N_47469);
and U48657 (N_48657,N_47328,N_47819);
nor U48658 (N_48658,N_47285,N_46449);
nor U48659 (N_48659,N_46759,N_46933);
or U48660 (N_48660,N_47716,N_46808);
xnor U48661 (N_48661,N_46893,N_46389);
nand U48662 (N_48662,N_46069,N_46301);
and U48663 (N_48663,N_46124,N_47619);
xnor U48664 (N_48664,N_47278,N_46228);
or U48665 (N_48665,N_47292,N_47076);
or U48666 (N_48666,N_47225,N_47449);
nor U48667 (N_48667,N_47820,N_46063);
nor U48668 (N_48668,N_46234,N_46711);
xor U48669 (N_48669,N_47830,N_46006);
and U48670 (N_48670,N_46526,N_46777);
nand U48671 (N_48671,N_47401,N_46752);
xor U48672 (N_48672,N_46888,N_47227);
or U48673 (N_48673,N_46144,N_47650);
nand U48674 (N_48674,N_46520,N_47490);
nor U48675 (N_48675,N_47807,N_46979);
xor U48676 (N_48676,N_47804,N_47121);
and U48677 (N_48677,N_47581,N_46014);
nand U48678 (N_48678,N_47734,N_47504);
nor U48679 (N_48679,N_47551,N_47123);
and U48680 (N_48680,N_46490,N_46319);
xnor U48681 (N_48681,N_47379,N_47282);
nor U48682 (N_48682,N_46611,N_46471);
and U48683 (N_48683,N_47518,N_46584);
nor U48684 (N_48684,N_47708,N_46783);
or U48685 (N_48685,N_46773,N_46613);
nand U48686 (N_48686,N_46861,N_47342);
nor U48687 (N_48687,N_46502,N_47937);
and U48688 (N_48688,N_47806,N_47783);
nor U48689 (N_48689,N_47846,N_47167);
nand U48690 (N_48690,N_47754,N_47714);
nor U48691 (N_48691,N_47543,N_46450);
and U48692 (N_48692,N_47207,N_46549);
or U48693 (N_48693,N_46398,N_46944);
nor U48694 (N_48694,N_47717,N_46887);
or U48695 (N_48695,N_47190,N_47631);
and U48696 (N_48696,N_47583,N_47585);
and U48697 (N_48697,N_47063,N_46092);
nor U48698 (N_48698,N_47039,N_46801);
xor U48699 (N_48699,N_46508,N_47168);
and U48700 (N_48700,N_47089,N_46877);
xor U48701 (N_48701,N_47393,N_46696);
xnor U48702 (N_48702,N_46195,N_47767);
xnor U48703 (N_48703,N_46921,N_46332);
nor U48704 (N_48704,N_47483,N_47649);
or U48705 (N_48705,N_46479,N_46413);
xor U48706 (N_48706,N_47360,N_46188);
xnor U48707 (N_48707,N_47679,N_46516);
xor U48708 (N_48708,N_47239,N_46807);
or U48709 (N_48709,N_47614,N_46011);
nor U48710 (N_48710,N_46341,N_46535);
nor U48711 (N_48711,N_46477,N_46023);
nand U48712 (N_48712,N_46303,N_46327);
or U48713 (N_48713,N_47894,N_46730);
nor U48714 (N_48714,N_46478,N_46842);
or U48715 (N_48715,N_47905,N_46079);
or U48716 (N_48716,N_46348,N_46267);
xor U48717 (N_48717,N_46597,N_46633);
xor U48718 (N_48718,N_46865,N_46591);
nor U48719 (N_48719,N_47972,N_46166);
or U48720 (N_48720,N_46991,N_47709);
nor U48721 (N_48721,N_46736,N_46563);
or U48722 (N_48722,N_46647,N_47973);
or U48723 (N_48723,N_46859,N_46352);
nor U48724 (N_48724,N_47382,N_46155);
nand U48725 (N_48725,N_47476,N_46509);
nor U48726 (N_48726,N_47394,N_46346);
nor U48727 (N_48727,N_46729,N_47759);
nand U48728 (N_48728,N_47844,N_46044);
and U48729 (N_48729,N_47011,N_46070);
nor U48730 (N_48730,N_46650,N_47020);
nor U48731 (N_48731,N_46975,N_46302);
or U48732 (N_48732,N_46924,N_47930);
nor U48733 (N_48733,N_46022,N_46115);
nor U48734 (N_48734,N_47186,N_46184);
or U48735 (N_48735,N_47410,N_46029);
nor U48736 (N_48736,N_47408,N_47921);
nor U48737 (N_48737,N_46078,N_46077);
nor U48738 (N_48738,N_46225,N_46554);
xor U48739 (N_48739,N_46487,N_46912);
or U48740 (N_48740,N_46559,N_47798);
xor U48741 (N_48741,N_46949,N_46746);
nand U48742 (N_48742,N_47896,N_47663);
and U48743 (N_48743,N_46616,N_47372);
or U48744 (N_48744,N_47865,N_46753);
or U48745 (N_48745,N_46672,N_47986);
nand U48746 (N_48746,N_46957,N_47439);
nand U48747 (N_48747,N_46862,N_47361);
nand U48748 (N_48748,N_46037,N_47216);
nor U48749 (N_48749,N_46137,N_46058);
and U48750 (N_48750,N_47536,N_46982);
or U48751 (N_48751,N_47922,N_46429);
nand U48752 (N_48752,N_47793,N_46150);
nor U48753 (N_48753,N_47860,N_46087);
nand U48754 (N_48754,N_46834,N_47238);
xor U48755 (N_48755,N_46863,N_47352);
nor U48756 (N_48756,N_46019,N_46474);
xor U48757 (N_48757,N_46269,N_46376);
and U48758 (N_48758,N_47090,N_46985);
nor U48759 (N_48759,N_47710,N_46823);
nand U48760 (N_48760,N_47270,N_46364);
nor U48761 (N_48761,N_46409,N_47474);
nand U48762 (N_48762,N_46291,N_47920);
or U48763 (N_48763,N_47212,N_47606);
xnor U48764 (N_48764,N_47118,N_46655);
nand U48765 (N_48765,N_47544,N_46879);
xor U48766 (N_48766,N_46561,N_46419);
nand U48767 (N_48767,N_46618,N_47881);
nand U48768 (N_48768,N_46157,N_46690);
nor U48769 (N_48769,N_46648,N_46518);
nand U48770 (N_48770,N_47887,N_47448);
nand U48771 (N_48771,N_47289,N_47810);
xnor U48772 (N_48772,N_47277,N_47287);
and U48773 (N_48773,N_47647,N_47305);
nor U48774 (N_48774,N_46725,N_47685);
or U48775 (N_48775,N_46146,N_47073);
xor U48776 (N_48776,N_47590,N_47635);
nor U48777 (N_48777,N_46587,N_46589);
and U48778 (N_48778,N_47602,N_46903);
nor U48779 (N_48779,N_46314,N_46700);
and U48780 (N_48780,N_46571,N_46321);
and U48781 (N_48781,N_47566,N_46039);
nor U48782 (N_48782,N_46866,N_46142);
xnor U48783 (N_48783,N_47962,N_46829);
and U48784 (N_48784,N_47269,N_46198);
nand U48785 (N_48785,N_47593,N_46123);
xnor U48786 (N_48786,N_46539,N_46909);
and U48787 (N_48787,N_46811,N_46541);
nand U48788 (N_48788,N_46485,N_46993);
or U48789 (N_48789,N_47673,N_47371);
xor U48790 (N_48790,N_46706,N_47149);
nor U48791 (N_48791,N_47821,N_47630);
and U48792 (N_48792,N_46798,N_47088);
nand U48793 (N_48793,N_47691,N_46791);
nor U48794 (N_48794,N_46207,N_46728);
nor U48795 (N_48795,N_47648,N_46310);
nand U48796 (N_48796,N_47915,N_47572);
nand U48797 (N_48797,N_47662,N_46828);
nand U48798 (N_48798,N_47756,N_46564);
nor U48799 (N_48799,N_46176,N_47111);
and U48800 (N_48800,N_46094,N_46182);
and U48801 (N_48801,N_46271,N_47386);
or U48802 (N_48802,N_46943,N_47777);
nor U48803 (N_48803,N_47131,N_46699);
nand U48804 (N_48804,N_46963,N_46064);
nand U48805 (N_48805,N_47811,N_46702);
nand U48806 (N_48806,N_46822,N_46789);
nor U48807 (N_48807,N_47113,N_46200);
or U48808 (N_48808,N_46261,N_47062);
nor U48809 (N_48809,N_47580,N_47961);
nor U48810 (N_48810,N_46345,N_47358);
xnor U48811 (N_48811,N_46590,N_47144);
and U48812 (N_48812,N_47497,N_47916);
and U48813 (N_48813,N_47106,N_46106);
and U48814 (N_48814,N_47758,N_46159);
nor U48815 (N_48815,N_46812,N_46939);
or U48816 (N_48816,N_47365,N_46387);
nor U48817 (N_48817,N_47694,N_46932);
nor U48818 (N_48818,N_46658,N_47936);
nand U48819 (N_48819,N_46854,N_47370);
xnor U48820 (N_48820,N_47231,N_46460);
or U48821 (N_48821,N_47007,N_47775);
nand U48822 (N_48822,N_46088,N_47030);
and U48823 (N_48823,N_47560,N_46102);
nor U48824 (N_48824,N_47054,N_46528);
xnor U48825 (N_48825,N_46163,N_46756);
and U48826 (N_48826,N_47311,N_47568);
xor U48827 (N_48827,N_46407,N_46190);
or U48828 (N_48828,N_47139,N_46457);
nand U48829 (N_48829,N_47523,N_47440);
or U48830 (N_48830,N_47537,N_46809);
nand U48831 (N_48831,N_47171,N_47307);
and U48832 (N_48832,N_46906,N_46365);
nand U48833 (N_48833,N_47688,N_46814);
nor U48834 (N_48834,N_46790,N_47156);
xor U48835 (N_48835,N_47974,N_47025);
or U48836 (N_48836,N_46203,N_47715);
and U48837 (N_48837,N_46832,N_47247);
or U48838 (N_48838,N_47326,N_46977);
nand U48839 (N_48839,N_47931,N_47180);
or U48840 (N_48840,N_46978,N_47596);
nand U48841 (N_48841,N_47565,N_46740);
nor U48842 (N_48842,N_47249,N_47163);
and U48843 (N_48843,N_46666,N_47676);
or U48844 (N_48844,N_46046,N_47336);
nand U48845 (N_48845,N_46435,N_46193);
and U48846 (N_48846,N_46305,N_47573);
xor U48847 (N_48847,N_47322,N_47949);
xor U48848 (N_48848,N_47561,N_47903);
nand U48849 (N_48849,N_46067,N_47347);
or U48850 (N_48850,N_46083,N_46139);
nand U48851 (N_48851,N_47017,N_46281);
nor U48852 (N_48852,N_47607,N_47741);
nor U48853 (N_48853,N_46915,N_46997);
and U48854 (N_48854,N_46805,N_47104);
and U48855 (N_48855,N_46687,N_47303);
xor U48856 (N_48856,N_46386,N_46247);
xor U48857 (N_48857,N_47173,N_47595);
xor U48858 (N_48858,N_46595,N_46698);
nand U48859 (N_48859,N_47045,N_46445);
xor U48860 (N_48860,N_46116,N_46488);
and U48861 (N_48861,N_46017,N_46211);
xor U48862 (N_48862,N_47458,N_47047);
nand U48863 (N_48863,N_46340,N_47885);
and U48864 (N_48864,N_46599,N_47782);
and U48865 (N_48865,N_46631,N_47114);
nor U48866 (N_48866,N_46959,N_47521);
and U48867 (N_48867,N_46434,N_46021);
xnor U48868 (N_48868,N_46607,N_46295);
or U48869 (N_48869,N_47712,N_47266);
nor U48870 (N_48870,N_47542,N_47976);
or U48871 (N_48871,N_46475,N_47592);
or U48872 (N_48872,N_46614,N_46653);
nor U48873 (N_48873,N_46277,N_47250);
xnor U48874 (N_48874,N_46491,N_47357);
or U48875 (N_48875,N_47960,N_47010);
xnor U48876 (N_48876,N_46482,N_47400);
nor U48877 (N_48877,N_47383,N_46055);
or U48878 (N_48878,N_47288,N_47757);
xnor U48879 (N_48879,N_46433,N_47155);
and U48880 (N_48880,N_46922,N_46850);
xnor U48881 (N_48881,N_46263,N_47191);
nand U48882 (N_48882,N_46731,N_47723);
nor U48883 (N_48883,N_47202,N_46060);
and U48884 (N_48884,N_46627,N_47411);
nand U48885 (N_48885,N_46692,N_47837);
or U48886 (N_48886,N_47421,N_46191);
nand U48887 (N_48887,N_47205,N_47610);
or U48888 (N_48888,N_47354,N_46680);
or U48889 (N_48889,N_46481,N_47599);
and U48890 (N_48890,N_46890,N_47430);
or U48891 (N_48891,N_47454,N_46686);
and U48892 (N_48892,N_47259,N_47075);
or U48893 (N_48893,N_46463,N_46447);
nor U48894 (N_48894,N_47456,N_47874);
nor U48895 (N_48895,N_46483,N_47652);
nand U48896 (N_48896,N_47306,N_46257);
and U48897 (N_48897,N_46330,N_46410);
xnor U48898 (N_48898,N_47330,N_46530);
or U48899 (N_48899,N_46390,N_46840);
and U48900 (N_48900,N_47422,N_46868);
or U48901 (N_48901,N_47995,N_46086);
xnor U48902 (N_48902,N_46394,N_47423);
nand U48903 (N_48903,N_46117,N_46625);
nand U48904 (N_48904,N_47321,N_47516);
xor U48905 (N_48905,N_47196,N_46966);
xor U48906 (N_48906,N_46721,N_46196);
xnor U48907 (N_48907,N_46838,N_46767);
xnor U48908 (N_48908,N_47829,N_47085);
nand U48909 (N_48909,N_46596,N_46468);
and U48910 (N_48910,N_46998,N_46082);
nor U48911 (N_48911,N_47985,N_47002);
nor U48912 (N_48912,N_46105,N_46401);
xnor U48913 (N_48913,N_47863,N_46331);
xor U48914 (N_48914,N_47204,N_47416);
nand U48915 (N_48915,N_47213,N_46076);
xnor U48916 (N_48916,N_47888,N_47368);
or U48917 (N_48917,N_47384,N_47823);
and U48918 (N_48918,N_46668,N_47641);
or U48919 (N_48919,N_47706,N_46383);
xor U48920 (N_48920,N_47719,N_47501);
nor U48921 (N_48921,N_46948,N_46054);
and U48922 (N_48922,N_46164,N_46112);
nor U48923 (N_48923,N_47348,N_46951);
nand U48924 (N_48924,N_47969,N_46907);
or U48925 (N_48925,N_47872,N_46709);
xnor U48926 (N_48926,N_46841,N_47945);
and U48927 (N_48927,N_46405,N_47158);
nor U48928 (N_48928,N_46334,N_47678);
xnor U48929 (N_48929,N_47835,N_47643);
or U48930 (N_48930,N_47391,N_46253);
nand U48931 (N_48931,N_46015,N_46603);
nand U48932 (N_48932,N_47994,N_46510);
nand U48933 (N_48933,N_46930,N_47359);
nor U48934 (N_48934,N_47505,N_46905);
nand U48935 (N_48935,N_46095,N_47548);
xor U48936 (N_48936,N_46743,N_47072);
nand U48937 (N_48937,N_47859,N_46722);
xor U48938 (N_48938,N_46913,N_46896);
or U48939 (N_48939,N_46883,N_46818);
nor U48940 (N_48940,N_46292,N_47427);
xnor U48941 (N_48941,N_47373,N_46187);
or U48942 (N_48942,N_46630,N_47791);
xor U48943 (N_48943,N_47378,N_46246);
or U48944 (N_48944,N_47467,N_46778);
and U48945 (N_48945,N_46210,N_47014);
nand U48946 (N_48946,N_47527,N_47848);
nand U48947 (N_48947,N_46496,N_46515);
nor U48948 (N_48948,N_46987,N_46240);
xor U48949 (N_48949,N_46772,N_46542);
nor U48950 (N_48950,N_47753,N_47027);
nand U48951 (N_48951,N_47141,N_47979);
nor U48952 (N_48952,N_46537,N_47752);
nand U48953 (N_48953,N_47436,N_47987);
or U48954 (N_48954,N_47914,N_46555);
or U48955 (N_48955,N_46788,N_47457);
or U48956 (N_48956,N_47746,N_46049);
or U48957 (N_48957,N_47093,N_47938);
nand U48958 (N_48958,N_46768,N_46012);
nor U48959 (N_48959,N_47246,N_47124);
nand U48960 (N_48960,N_47988,N_47493);
and U48961 (N_48961,N_46695,N_47087);
nor U48962 (N_48962,N_47534,N_46986);
nand U48963 (N_48963,N_47901,N_46499);
nand U48964 (N_48964,N_46602,N_46311);
xnor U48965 (N_48965,N_46857,N_47353);
nor U48966 (N_48966,N_46720,N_46202);
or U48967 (N_48967,N_47666,N_46098);
and U48968 (N_48968,N_46503,N_46304);
nor U48969 (N_48969,N_46351,N_47310);
nor U48970 (N_48970,N_46629,N_47645);
xnor U48971 (N_48971,N_46180,N_47182);
nor U48972 (N_48972,N_46378,N_46366);
xnor U48973 (N_48973,N_46108,N_46718);
nor U48974 (N_48974,N_46755,N_47531);
nor U48975 (N_48975,N_47064,N_46910);
xnor U48976 (N_48976,N_46976,N_46013);
nor U48977 (N_48977,N_47858,N_46900);
nand U48978 (N_48978,N_46855,N_47046);
xnor U48979 (N_48979,N_46493,N_47334);
xnor U48980 (N_48980,N_46780,N_47364);
and U48981 (N_48981,N_47258,N_47575);
xor U48982 (N_48982,N_46565,N_46452);
nor U48983 (N_48983,N_46677,N_47801);
xor U48984 (N_48984,N_46358,N_47626);
and U48985 (N_48985,N_46308,N_46947);
nor U48986 (N_48986,N_46118,N_46739);
and U48987 (N_48987,N_46886,N_47295);
and U48988 (N_48988,N_46762,N_47395);
nor U48989 (N_48989,N_47744,N_46856);
xor U48990 (N_48990,N_47943,N_46534);
nor U48991 (N_48991,N_46048,N_47904);
nor U48992 (N_48992,N_46455,N_46495);
xnor U48993 (N_48993,N_46545,N_46671);
and U48994 (N_48994,N_47700,N_47344);
and U48995 (N_48995,N_46833,N_47735);
nor U48996 (N_48996,N_47556,N_46465);
nor U48997 (N_48997,N_47153,N_47036);
nor U48998 (N_48998,N_46682,N_47366);
xor U48999 (N_48999,N_47160,N_46547);
nor U49000 (N_49000,N_47260,N_47215);
nor U49001 (N_49001,N_46123,N_47015);
nand U49002 (N_49002,N_47347,N_46916);
and U49003 (N_49003,N_46881,N_46352);
nand U49004 (N_49004,N_47308,N_46958);
xnor U49005 (N_49005,N_47935,N_46961);
nor U49006 (N_49006,N_46742,N_47268);
nand U49007 (N_49007,N_46490,N_46360);
and U49008 (N_49008,N_47798,N_46161);
or U49009 (N_49009,N_47943,N_47379);
nor U49010 (N_49010,N_46165,N_47292);
nand U49011 (N_49011,N_46142,N_46553);
nand U49012 (N_49012,N_47427,N_47472);
and U49013 (N_49013,N_46607,N_46292);
and U49014 (N_49014,N_46853,N_46485);
nor U49015 (N_49015,N_47587,N_46678);
xor U49016 (N_49016,N_47642,N_46985);
nand U49017 (N_49017,N_46815,N_47021);
nor U49018 (N_49018,N_47782,N_47124);
nand U49019 (N_49019,N_46529,N_47525);
xnor U49020 (N_49020,N_46081,N_46203);
xor U49021 (N_49021,N_47959,N_46959);
nand U49022 (N_49022,N_46800,N_46544);
and U49023 (N_49023,N_46832,N_46297);
and U49024 (N_49024,N_46708,N_47917);
xor U49025 (N_49025,N_47506,N_47607);
xor U49026 (N_49026,N_46587,N_46405);
nor U49027 (N_49027,N_46312,N_46604);
nor U49028 (N_49028,N_47952,N_46396);
nor U49029 (N_49029,N_46186,N_47889);
nand U49030 (N_49030,N_46856,N_47852);
nand U49031 (N_49031,N_47495,N_47359);
nand U49032 (N_49032,N_46786,N_46919);
or U49033 (N_49033,N_46064,N_47595);
nand U49034 (N_49034,N_47982,N_46847);
or U49035 (N_49035,N_46750,N_46568);
xor U49036 (N_49036,N_46846,N_46581);
nand U49037 (N_49037,N_47262,N_47757);
nand U49038 (N_49038,N_46215,N_46808);
and U49039 (N_49039,N_46446,N_46997);
nand U49040 (N_49040,N_46989,N_47968);
xnor U49041 (N_49041,N_46996,N_47650);
nand U49042 (N_49042,N_46604,N_46893);
or U49043 (N_49043,N_46556,N_46292);
nand U49044 (N_49044,N_46606,N_47090);
nor U49045 (N_49045,N_47209,N_46406);
nor U49046 (N_49046,N_47133,N_47021);
nor U49047 (N_49047,N_47769,N_47968);
or U49048 (N_49048,N_47129,N_46315);
nor U49049 (N_49049,N_46993,N_46404);
nor U49050 (N_49050,N_47717,N_46164);
nand U49051 (N_49051,N_47580,N_47510);
and U49052 (N_49052,N_47308,N_47939);
and U49053 (N_49053,N_47283,N_46681);
or U49054 (N_49054,N_46511,N_46003);
nand U49055 (N_49055,N_46346,N_46545);
and U49056 (N_49056,N_47897,N_47394);
and U49057 (N_49057,N_47689,N_47022);
and U49058 (N_49058,N_47949,N_47586);
or U49059 (N_49059,N_47564,N_46673);
or U49060 (N_49060,N_47640,N_46649);
nor U49061 (N_49061,N_46039,N_46638);
nor U49062 (N_49062,N_46160,N_46263);
nor U49063 (N_49063,N_47990,N_47716);
and U49064 (N_49064,N_46100,N_46735);
and U49065 (N_49065,N_47652,N_46230);
and U49066 (N_49066,N_47702,N_46658);
nor U49067 (N_49067,N_47523,N_47631);
nor U49068 (N_49068,N_47168,N_47450);
nand U49069 (N_49069,N_46044,N_46879);
nand U49070 (N_49070,N_47877,N_46545);
and U49071 (N_49071,N_47277,N_46410);
and U49072 (N_49072,N_47676,N_46876);
or U49073 (N_49073,N_46697,N_47014);
or U49074 (N_49074,N_46506,N_46818);
or U49075 (N_49075,N_46621,N_46670);
nor U49076 (N_49076,N_47204,N_46266);
or U49077 (N_49077,N_47134,N_47306);
nor U49078 (N_49078,N_47294,N_46148);
xnor U49079 (N_49079,N_47317,N_47704);
nand U49080 (N_49080,N_47627,N_46782);
or U49081 (N_49081,N_47189,N_47608);
xnor U49082 (N_49082,N_46402,N_47031);
nand U49083 (N_49083,N_46895,N_47809);
nand U49084 (N_49084,N_47064,N_47608);
xnor U49085 (N_49085,N_46900,N_47612);
or U49086 (N_49086,N_46825,N_47623);
and U49087 (N_49087,N_46831,N_47312);
nor U49088 (N_49088,N_46647,N_47834);
and U49089 (N_49089,N_47316,N_47590);
and U49090 (N_49090,N_46770,N_47826);
or U49091 (N_49091,N_46431,N_47713);
and U49092 (N_49092,N_47767,N_46636);
or U49093 (N_49093,N_47460,N_47241);
xnor U49094 (N_49094,N_47258,N_46642);
nand U49095 (N_49095,N_46816,N_46932);
nor U49096 (N_49096,N_46893,N_47721);
nand U49097 (N_49097,N_47673,N_47938);
nand U49098 (N_49098,N_47473,N_46760);
nand U49099 (N_49099,N_46174,N_46514);
nor U49100 (N_49100,N_47064,N_47449);
and U49101 (N_49101,N_47258,N_46347);
and U49102 (N_49102,N_47089,N_46058);
nand U49103 (N_49103,N_46090,N_46920);
xnor U49104 (N_49104,N_47886,N_47980);
or U49105 (N_49105,N_47746,N_47362);
nand U49106 (N_49106,N_47267,N_47999);
xnor U49107 (N_49107,N_47389,N_47369);
or U49108 (N_49108,N_47927,N_46775);
and U49109 (N_49109,N_46780,N_47370);
and U49110 (N_49110,N_47161,N_47066);
xor U49111 (N_49111,N_46463,N_46386);
xnor U49112 (N_49112,N_47062,N_46431);
xor U49113 (N_49113,N_46533,N_46433);
xnor U49114 (N_49114,N_46632,N_46075);
and U49115 (N_49115,N_47885,N_47535);
nand U49116 (N_49116,N_46141,N_47147);
and U49117 (N_49117,N_46065,N_47633);
and U49118 (N_49118,N_47304,N_46125);
nor U49119 (N_49119,N_46643,N_46701);
or U49120 (N_49120,N_46391,N_46099);
or U49121 (N_49121,N_47094,N_46308);
or U49122 (N_49122,N_47761,N_46443);
and U49123 (N_49123,N_46945,N_46034);
or U49124 (N_49124,N_47535,N_46725);
or U49125 (N_49125,N_47877,N_47495);
nor U49126 (N_49126,N_46171,N_47503);
xor U49127 (N_49127,N_47409,N_46046);
nand U49128 (N_49128,N_46346,N_47118);
nor U49129 (N_49129,N_47354,N_47532);
and U49130 (N_49130,N_47692,N_47142);
nor U49131 (N_49131,N_47971,N_46735);
or U49132 (N_49132,N_46713,N_46826);
or U49133 (N_49133,N_47997,N_46063);
nand U49134 (N_49134,N_46426,N_46211);
or U49135 (N_49135,N_46636,N_47761);
or U49136 (N_49136,N_46069,N_47403);
nand U49137 (N_49137,N_47283,N_46703);
or U49138 (N_49138,N_46717,N_47705);
or U49139 (N_49139,N_47684,N_46752);
xor U49140 (N_49140,N_47690,N_46974);
xor U49141 (N_49141,N_46478,N_47226);
or U49142 (N_49142,N_46326,N_47611);
and U49143 (N_49143,N_46637,N_46170);
xnor U49144 (N_49144,N_47998,N_46695);
or U49145 (N_49145,N_47804,N_47505);
or U49146 (N_49146,N_46515,N_47059);
and U49147 (N_49147,N_47605,N_46710);
nand U49148 (N_49148,N_47275,N_46621);
nand U49149 (N_49149,N_47776,N_46310);
nand U49150 (N_49150,N_47302,N_47667);
and U49151 (N_49151,N_46092,N_46293);
and U49152 (N_49152,N_46382,N_47127);
and U49153 (N_49153,N_47786,N_46591);
nand U49154 (N_49154,N_47721,N_46616);
nand U49155 (N_49155,N_46696,N_46481);
nor U49156 (N_49156,N_47062,N_47380);
nand U49157 (N_49157,N_46732,N_47362);
xor U49158 (N_49158,N_47985,N_46438);
nor U49159 (N_49159,N_46891,N_46493);
or U49160 (N_49160,N_47677,N_46067);
xnor U49161 (N_49161,N_47604,N_47353);
nor U49162 (N_49162,N_46654,N_47769);
or U49163 (N_49163,N_47960,N_46115);
and U49164 (N_49164,N_47048,N_47621);
nand U49165 (N_49165,N_46554,N_46572);
nor U49166 (N_49166,N_47946,N_46198);
nor U49167 (N_49167,N_46926,N_47741);
nor U49168 (N_49168,N_47182,N_47833);
nand U49169 (N_49169,N_46037,N_47447);
and U49170 (N_49170,N_47116,N_46896);
xor U49171 (N_49171,N_46572,N_47441);
nand U49172 (N_49172,N_47959,N_47890);
or U49173 (N_49173,N_47637,N_47569);
or U49174 (N_49174,N_46991,N_46695);
and U49175 (N_49175,N_47220,N_46287);
nor U49176 (N_49176,N_47138,N_47950);
nor U49177 (N_49177,N_46182,N_46125);
or U49178 (N_49178,N_47447,N_47967);
xor U49179 (N_49179,N_46271,N_47653);
or U49180 (N_49180,N_47301,N_47877);
nor U49181 (N_49181,N_47437,N_47556);
nand U49182 (N_49182,N_46302,N_46331);
or U49183 (N_49183,N_46946,N_46859);
nor U49184 (N_49184,N_46490,N_47390);
nand U49185 (N_49185,N_46720,N_46618);
xnor U49186 (N_49186,N_47156,N_46322);
nand U49187 (N_49187,N_47520,N_46182);
xor U49188 (N_49188,N_47012,N_46345);
or U49189 (N_49189,N_46308,N_47886);
or U49190 (N_49190,N_47523,N_46092);
nand U49191 (N_49191,N_47212,N_47005);
nor U49192 (N_49192,N_46010,N_46258);
or U49193 (N_49193,N_47409,N_47011);
or U49194 (N_49194,N_47479,N_47322);
or U49195 (N_49195,N_47922,N_46400);
nand U49196 (N_49196,N_47927,N_46709);
nor U49197 (N_49197,N_47157,N_46810);
and U49198 (N_49198,N_46427,N_46394);
or U49199 (N_49199,N_46807,N_47558);
nor U49200 (N_49200,N_47013,N_46782);
and U49201 (N_49201,N_47040,N_47155);
xor U49202 (N_49202,N_47074,N_47715);
nand U49203 (N_49203,N_46088,N_47490);
nand U49204 (N_49204,N_46417,N_46953);
nor U49205 (N_49205,N_46088,N_46633);
nor U49206 (N_49206,N_46578,N_47286);
and U49207 (N_49207,N_47435,N_46154);
nor U49208 (N_49208,N_46247,N_46165);
or U49209 (N_49209,N_47869,N_46797);
xor U49210 (N_49210,N_46411,N_46812);
xor U49211 (N_49211,N_47072,N_46142);
xor U49212 (N_49212,N_47401,N_47169);
nor U49213 (N_49213,N_46741,N_47657);
nor U49214 (N_49214,N_47806,N_46744);
nor U49215 (N_49215,N_47964,N_46964);
and U49216 (N_49216,N_46996,N_47337);
xnor U49217 (N_49217,N_46181,N_47147);
or U49218 (N_49218,N_46817,N_46366);
nand U49219 (N_49219,N_47372,N_47183);
nand U49220 (N_49220,N_46463,N_46169);
or U49221 (N_49221,N_47018,N_46454);
xnor U49222 (N_49222,N_47517,N_46057);
nor U49223 (N_49223,N_46517,N_47948);
nor U49224 (N_49224,N_46221,N_46016);
and U49225 (N_49225,N_46034,N_47803);
or U49226 (N_49226,N_47441,N_46117);
xor U49227 (N_49227,N_46796,N_46281);
and U49228 (N_49228,N_47976,N_47030);
nand U49229 (N_49229,N_47624,N_46927);
nor U49230 (N_49230,N_46438,N_46762);
and U49231 (N_49231,N_47083,N_46726);
or U49232 (N_49232,N_46605,N_46371);
or U49233 (N_49233,N_47931,N_46250);
nor U49234 (N_49234,N_46299,N_47895);
nand U49235 (N_49235,N_47164,N_47295);
and U49236 (N_49236,N_46105,N_47332);
xor U49237 (N_49237,N_46614,N_46120);
xor U49238 (N_49238,N_47729,N_46987);
or U49239 (N_49239,N_47950,N_46169);
xor U49240 (N_49240,N_46573,N_46982);
nor U49241 (N_49241,N_46189,N_47407);
or U49242 (N_49242,N_46313,N_46934);
and U49243 (N_49243,N_47265,N_47248);
or U49244 (N_49244,N_46788,N_47654);
nand U49245 (N_49245,N_47488,N_47852);
or U49246 (N_49246,N_47068,N_46888);
xor U49247 (N_49247,N_46475,N_46554);
nand U49248 (N_49248,N_47195,N_47154);
and U49249 (N_49249,N_47845,N_47997);
and U49250 (N_49250,N_46807,N_47449);
xor U49251 (N_49251,N_46455,N_47678);
nand U49252 (N_49252,N_46694,N_46471);
nand U49253 (N_49253,N_46442,N_46645);
or U49254 (N_49254,N_46113,N_47914);
xnor U49255 (N_49255,N_47427,N_47553);
or U49256 (N_49256,N_46348,N_47584);
and U49257 (N_49257,N_47034,N_47511);
nand U49258 (N_49258,N_46888,N_46856);
nand U49259 (N_49259,N_46138,N_46769);
and U49260 (N_49260,N_46216,N_46813);
nand U49261 (N_49261,N_46198,N_46088);
nor U49262 (N_49262,N_46359,N_46209);
or U49263 (N_49263,N_47479,N_46119);
nor U49264 (N_49264,N_46495,N_46380);
or U49265 (N_49265,N_46751,N_46504);
or U49266 (N_49266,N_46611,N_47367);
or U49267 (N_49267,N_46316,N_46992);
or U49268 (N_49268,N_47529,N_46460);
xnor U49269 (N_49269,N_46784,N_46292);
xor U49270 (N_49270,N_47873,N_47839);
xnor U49271 (N_49271,N_47140,N_46362);
xor U49272 (N_49272,N_46855,N_46579);
nand U49273 (N_49273,N_46645,N_46539);
or U49274 (N_49274,N_47922,N_46818);
or U49275 (N_49275,N_47400,N_47278);
nor U49276 (N_49276,N_47012,N_47198);
nand U49277 (N_49277,N_46372,N_47426);
nor U49278 (N_49278,N_47590,N_46687);
or U49279 (N_49279,N_47257,N_47239);
and U49280 (N_49280,N_46445,N_46728);
and U49281 (N_49281,N_46082,N_47906);
and U49282 (N_49282,N_47224,N_46970);
nor U49283 (N_49283,N_47212,N_46689);
nand U49284 (N_49284,N_47920,N_47279);
nand U49285 (N_49285,N_47404,N_46855);
and U49286 (N_49286,N_47178,N_46036);
or U49287 (N_49287,N_46778,N_46992);
nor U49288 (N_49288,N_47202,N_47711);
or U49289 (N_49289,N_46419,N_47197);
xnor U49290 (N_49290,N_47042,N_46757);
or U49291 (N_49291,N_46414,N_47835);
xnor U49292 (N_49292,N_47635,N_46168);
and U49293 (N_49293,N_47597,N_46791);
nor U49294 (N_49294,N_47196,N_46622);
and U49295 (N_49295,N_46674,N_46060);
xnor U49296 (N_49296,N_46097,N_46279);
nand U49297 (N_49297,N_47479,N_47218);
or U49298 (N_49298,N_46797,N_46183);
nor U49299 (N_49299,N_46824,N_46696);
xnor U49300 (N_49300,N_46395,N_47956);
nor U49301 (N_49301,N_47670,N_47009);
and U49302 (N_49302,N_46697,N_47456);
or U49303 (N_49303,N_46973,N_47842);
nand U49304 (N_49304,N_46820,N_46238);
or U49305 (N_49305,N_46429,N_47037);
nand U49306 (N_49306,N_47632,N_46800);
nor U49307 (N_49307,N_47903,N_47309);
nand U49308 (N_49308,N_47842,N_46597);
nor U49309 (N_49309,N_46594,N_47348);
xnor U49310 (N_49310,N_46376,N_47430);
and U49311 (N_49311,N_47772,N_47414);
or U49312 (N_49312,N_47629,N_46891);
or U49313 (N_49313,N_47948,N_47596);
nand U49314 (N_49314,N_46204,N_46745);
nor U49315 (N_49315,N_47739,N_47801);
xnor U49316 (N_49316,N_46679,N_47086);
or U49317 (N_49317,N_47711,N_47298);
xor U49318 (N_49318,N_46066,N_47078);
and U49319 (N_49319,N_46957,N_46804);
nor U49320 (N_49320,N_46144,N_47738);
nor U49321 (N_49321,N_46153,N_46243);
or U49322 (N_49322,N_47005,N_46395);
xor U49323 (N_49323,N_46553,N_47785);
nand U49324 (N_49324,N_47588,N_47266);
nor U49325 (N_49325,N_47161,N_46872);
nand U49326 (N_49326,N_46449,N_46548);
nor U49327 (N_49327,N_47860,N_47176);
and U49328 (N_49328,N_46158,N_47270);
or U49329 (N_49329,N_46348,N_47840);
nor U49330 (N_49330,N_46618,N_46844);
and U49331 (N_49331,N_47958,N_47428);
nand U49332 (N_49332,N_47409,N_47809);
nor U49333 (N_49333,N_46098,N_47581);
and U49334 (N_49334,N_47893,N_46390);
nand U49335 (N_49335,N_47893,N_47860);
xor U49336 (N_49336,N_46242,N_47361);
nor U49337 (N_49337,N_46909,N_46089);
nor U49338 (N_49338,N_46680,N_47969);
nor U49339 (N_49339,N_46006,N_46866);
or U49340 (N_49340,N_46020,N_46797);
and U49341 (N_49341,N_47673,N_47748);
xnor U49342 (N_49342,N_46140,N_47364);
or U49343 (N_49343,N_47003,N_46511);
or U49344 (N_49344,N_47038,N_46116);
xnor U49345 (N_49345,N_46156,N_47334);
or U49346 (N_49346,N_47179,N_47861);
or U49347 (N_49347,N_47737,N_47861);
or U49348 (N_49348,N_46439,N_46285);
xnor U49349 (N_49349,N_46608,N_46225);
and U49350 (N_49350,N_47338,N_47379);
xnor U49351 (N_49351,N_46785,N_46636);
nor U49352 (N_49352,N_46304,N_46781);
nor U49353 (N_49353,N_46158,N_47912);
and U49354 (N_49354,N_47807,N_46717);
xnor U49355 (N_49355,N_46326,N_46338);
and U49356 (N_49356,N_47019,N_47968);
nor U49357 (N_49357,N_46311,N_47824);
nor U49358 (N_49358,N_46147,N_47694);
or U49359 (N_49359,N_46136,N_46497);
or U49360 (N_49360,N_47636,N_47901);
or U49361 (N_49361,N_46194,N_47447);
xor U49362 (N_49362,N_47559,N_47314);
nand U49363 (N_49363,N_46616,N_46124);
and U49364 (N_49364,N_46080,N_46931);
xnor U49365 (N_49365,N_47019,N_46345);
and U49366 (N_49366,N_47267,N_46940);
and U49367 (N_49367,N_46074,N_46580);
or U49368 (N_49368,N_47477,N_46270);
nand U49369 (N_49369,N_46135,N_46205);
and U49370 (N_49370,N_47923,N_46225);
nand U49371 (N_49371,N_46408,N_46113);
or U49372 (N_49372,N_46106,N_47138);
xnor U49373 (N_49373,N_46154,N_47810);
and U49374 (N_49374,N_46591,N_47588);
nor U49375 (N_49375,N_46910,N_46300);
or U49376 (N_49376,N_47923,N_46928);
nand U49377 (N_49377,N_47857,N_47000);
xnor U49378 (N_49378,N_47551,N_47308);
xnor U49379 (N_49379,N_46479,N_47120);
or U49380 (N_49380,N_46872,N_47888);
xor U49381 (N_49381,N_46068,N_46554);
xor U49382 (N_49382,N_47476,N_47873);
nand U49383 (N_49383,N_47785,N_46058);
xnor U49384 (N_49384,N_46711,N_47656);
and U49385 (N_49385,N_46069,N_46319);
nor U49386 (N_49386,N_47212,N_46805);
nor U49387 (N_49387,N_46839,N_46358);
or U49388 (N_49388,N_46395,N_46814);
nand U49389 (N_49389,N_46105,N_46580);
nand U49390 (N_49390,N_46275,N_47239);
or U49391 (N_49391,N_46408,N_46146);
and U49392 (N_49392,N_46404,N_47789);
nor U49393 (N_49393,N_46468,N_46608);
and U49394 (N_49394,N_47920,N_47016);
xor U49395 (N_49395,N_47534,N_46490);
and U49396 (N_49396,N_46265,N_47195);
nor U49397 (N_49397,N_47257,N_46540);
nand U49398 (N_49398,N_47742,N_46271);
nand U49399 (N_49399,N_47565,N_47476);
xnor U49400 (N_49400,N_47070,N_46537);
and U49401 (N_49401,N_47476,N_47691);
nand U49402 (N_49402,N_46003,N_46863);
and U49403 (N_49403,N_46606,N_46545);
nor U49404 (N_49404,N_46239,N_47397);
nand U49405 (N_49405,N_47833,N_47868);
nand U49406 (N_49406,N_46249,N_47956);
or U49407 (N_49407,N_47762,N_46767);
and U49408 (N_49408,N_46455,N_46158);
xnor U49409 (N_49409,N_46424,N_46610);
nor U49410 (N_49410,N_46286,N_47358);
nand U49411 (N_49411,N_46150,N_47424);
and U49412 (N_49412,N_47442,N_46418);
xnor U49413 (N_49413,N_47247,N_46069);
and U49414 (N_49414,N_46345,N_47899);
xor U49415 (N_49415,N_46257,N_46202);
xnor U49416 (N_49416,N_47306,N_46177);
nor U49417 (N_49417,N_47637,N_47620);
xnor U49418 (N_49418,N_46855,N_46658);
nor U49419 (N_49419,N_46187,N_46852);
nand U49420 (N_49420,N_47556,N_46709);
xor U49421 (N_49421,N_46469,N_46692);
and U49422 (N_49422,N_46814,N_46551);
nand U49423 (N_49423,N_47358,N_47728);
and U49424 (N_49424,N_46961,N_47594);
nor U49425 (N_49425,N_46555,N_47853);
nand U49426 (N_49426,N_47846,N_47129);
nand U49427 (N_49427,N_47439,N_47368);
and U49428 (N_49428,N_46598,N_46468);
nor U49429 (N_49429,N_46821,N_47368);
and U49430 (N_49430,N_46643,N_47763);
nand U49431 (N_49431,N_47004,N_47958);
nand U49432 (N_49432,N_46122,N_47485);
nand U49433 (N_49433,N_47801,N_47319);
nor U49434 (N_49434,N_47470,N_47647);
and U49435 (N_49435,N_47005,N_47103);
nor U49436 (N_49436,N_47164,N_46725);
xnor U49437 (N_49437,N_47249,N_47688);
nor U49438 (N_49438,N_46102,N_46528);
nor U49439 (N_49439,N_47386,N_46032);
and U49440 (N_49440,N_47988,N_47610);
nor U49441 (N_49441,N_47535,N_46470);
nand U49442 (N_49442,N_47330,N_47046);
nor U49443 (N_49443,N_47709,N_47572);
xnor U49444 (N_49444,N_47117,N_47101);
and U49445 (N_49445,N_47245,N_46126);
xor U49446 (N_49446,N_47990,N_47543);
and U49447 (N_49447,N_46637,N_46755);
and U49448 (N_49448,N_47241,N_47473);
nand U49449 (N_49449,N_47485,N_46339);
nand U49450 (N_49450,N_47814,N_46918);
or U49451 (N_49451,N_47763,N_46500);
and U49452 (N_49452,N_47200,N_47449);
nand U49453 (N_49453,N_47611,N_46250);
or U49454 (N_49454,N_46556,N_46062);
and U49455 (N_49455,N_46219,N_47695);
or U49456 (N_49456,N_46367,N_47741);
nor U49457 (N_49457,N_46456,N_47419);
xor U49458 (N_49458,N_47266,N_46452);
xor U49459 (N_49459,N_47590,N_47565);
xnor U49460 (N_49460,N_46799,N_46849);
nor U49461 (N_49461,N_47922,N_46044);
or U49462 (N_49462,N_47102,N_46708);
nor U49463 (N_49463,N_47977,N_47646);
nor U49464 (N_49464,N_47687,N_47350);
and U49465 (N_49465,N_47482,N_47917);
nor U49466 (N_49466,N_47138,N_47054);
xor U49467 (N_49467,N_46121,N_47543);
nand U49468 (N_49468,N_46219,N_46015);
nor U49469 (N_49469,N_47988,N_47355);
and U49470 (N_49470,N_47763,N_46604);
nand U49471 (N_49471,N_46182,N_46454);
nand U49472 (N_49472,N_46289,N_47741);
nand U49473 (N_49473,N_47987,N_46380);
and U49474 (N_49474,N_46013,N_46131);
or U49475 (N_49475,N_47017,N_47513);
nand U49476 (N_49476,N_46725,N_46060);
nand U49477 (N_49477,N_47178,N_47445);
xnor U49478 (N_49478,N_46379,N_46594);
nand U49479 (N_49479,N_47069,N_46981);
nand U49480 (N_49480,N_46099,N_46648);
and U49481 (N_49481,N_47356,N_46314);
xor U49482 (N_49482,N_47175,N_46042);
or U49483 (N_49483,N_47333,N_46639);
nand U49484 (N_49484,N_46025,N_47297);
nor U49485 (N_49485,N_47515,N_46479);
xor U49486 (N_49486,N_47142,N_47933);
xor U49487 (N_49487,N_47553,N_47740);
xnor U49488 (N_49488,N_47989,N_46240);
nand U49489 (N_49489,N_46494,N_47990);
or U49490 (N_49490,N_47995,N_46285);
nor U49491 (N_49491,N_47376,N_47182);
nor U49492 (N_49492,N_46644,N_46204);
nor U49493 (N_49493,N_47525,N_47740);
nor U49494 (N_49494,N_47588,N_46699);
xor U49495 (N_49495,N_46539,N_46827);
or U49496 (N_49496,N_46344,N_46820);
and U49497 (N_49497,N_47449,N_47945);
or U49498 (N_49498,N_46855,N_47922);
nand U49499 (N_49499,N_47785,N_47442);
xor U49500 (N_49500,N_47631,N_46403);
xor U49501 (N_49501,N_46931,N_47043);
xor U49502 (N_49502,N_47637,N_47545);
nor U49503 (N_49503,N_46332,N_47174);
or U49504 (N_49504,N_46433,N_46482);
and U49505 (N_49505,N_47298,N_46967);
and U49506 (N_49506,N_47158,N_47862);
nand U49507 (N_49507,N_47675,N_47136);
nand U49508 (N_49508,N_46155,N_47010);
nor U49509 (N_49509,N_47682,N_47101);
xor U49510 (N_49510,N_46381,N_46747);
or U49511 (N_49511,N_47897,N_46322);
nand U49512 (N_49512,N_46562,N_47016);
or U49513 (N_49513,N_47977,N_46519);
nor U49514 (N_49514,N_46828,N_46150);
and U49515 (N_49515,N_47267,N_46047);
or U49516 (N_49516,N_47312,N_47468);
xor U49517 (N_49517,N_46103,N_47400);
or U49518 (N_49518,N_47241,N_47662);
or U49519 (N_49519,N_46758,N_47819);
nor U49520 (N_49520,N_47270,N_47007);
or U49521 (N_49521,N_47104,N_46496);
nand U49522 (N_49522,N_46777,N_47322);
and U49523 (N_49523,N_47036,N_47979);
nand U49524 (N_49524,N_46072,N_46076);
nor U49525 (N_49525,N_46283,N_46313);
and U49526 (N_49526,N_46315,N_47173);
and U49527 (N_49527,N_47058,N_47956);
xor U49528 (N_49528,N_46469,N_47238);
xnor U49529 (N_49529,N_47756,N_46291);
or U49530 (N_49530,N_46861,N_46952);
nand U49531 (N_49531,N_46287,N_46671);
and U49532 (N_49532,N_46929,N_46941);
nor U49533 (N_49533,N_46119,N_47979);
and U49534 (N_49534,N_46856,N_47767);
and U49535 (N_49535,N_47434,N_47205);
and U49536 (N_49536,N_47141,N_46920);
and U49537 (N_49537,N_46537,N_47015);
and U49538 (N_49538,N_46354,N_46613);
xnor U49539 (N_49539,N_47954,N_47554);
nor U49540 (N_49540,N_47541,N_47670);
nand U49541 (N_49541,N_47019,N_46182);
nand U49542 (N_49542,N_46485,N_46544);
or U49543 (N_49543,N_46176,N_47683);
xnor U49544 (N_49544,N_47594,N_47198);
nor U49545 (N_49545,N_47111,N_46605);
or U49546 (N_49546,N_47351,N_47485);
xnor U49547 (N_49547,N_46010,N_47880);
nor U49548 (N_49548,N_46706,N_46328);
xor U49549 (N_49549,N_47818,N_46429);
and U49550 (N_49550,N_46482,N_47152);
nand U49551 (N_49551,N_46033,N_47880);
xor U49552 (N_49552,N_46298,N_46045);
nand U49553 (N_49553,N_46198,N_46766);
xnor U49554 (N_49554,N_47063,N_46673);
nand U49555 (N_49555,N_47931,N_47829);
xor U49556 (N_49556,N_47974,N_47692);
or U49557 (N_49557,N_47628,N_47869);
and U49558 (N_49558,N_46990,N_46939);
or U49559 (N_49559,N_46686,N_47754);
or U49560 (N_49560,N_47927,N_46792);
nor U49561 (N_49561,N_46049,N_47184);
xnor U49562 (N_49562,N_46077,N_46684);
nand U49563 (N_49563,N_47458,N_46167);
and U49564 (N_49564,N_47793,N_47679);
nor U49565 (N_49565,N_46859,N_46683);
nand U49566 (N_49566,N_47246,N_47212);
or U49567 (N_49567,N_46123,N_47085);
nand U49568 (N_49568,N_46949,N_47898);
or U49569 (N_49569,N_47790,N_47138);
and U49570 (N_49570,N_47018,N_47738);
or U49571 (N_49571,N_46802,N_47936);
xnor U49572 (N_49572,N_46630,N_47554);
nand U49573 (N_49573,N_47510,N_46847);
nand U49574 (N_49574,N_47295,N_47375);
or U49575 (N_49575,N_47917,N_46219);
xnor U49576 (N_49576,N_47837,N_47476);
nand U49577 (N_49577,N_47629,N_47719);
and U49578 (N_49578,N_47623,N_47490);
and U49579 (N_49579,N_46514,N_47144);
xor U49580 (N_49580,N_46908,N_47785);
nand U49581 (N_49581,N_47678,N_46414);
nor U49582 (N_49582,N_47634,N_46120);
xnor U49583 (N_49583,N_47462,N_46884);
or U49584 (N_49584,N_47293,N_47466);
nand U49585 (N_49585,N_46463,N_46888);
nor U49586 (N_49586,N_46351,N_47058);
nand U49587 (N_49587,N_46499,N_47462);
xnor U49588 (N_49588,N_46256,N_47584);
or U49589 (N_49589,N_46950,N_47171);
and U49590 (N_49590,N_46453,N_46204);
and U49591 (N_49591,N_47930,N_47087);
xnor U49592 (N_49592,N_46891,N_46396);
xor U49593 (N_49593,N_46010,N_47315);
and U49594 (N_49594,N_46878,N_46938);
and U49595 (N_49595,N_47935,N_46945);
xnor U49596 (N_49596,N_47907,N_46063);
or U49597 (N_49597,N_46273,N_46053);
and U49598 (N_49598,N_47332,N_47503);
xnor U49599 (N_49599,N_47648,N_46780);
nand U49600 (N_49600,N_47860,N_47199);
or U49601 (N_49601,N_46769,N_47479);
nand U49602 (N_49602,N_46790,N_46663);
xnor U49603 (N_49603,N_47548,N_47678);
or U49604 (N_49604,N_47177,N_47042);
nand U49605 (N_49605,N_46115,N_47104);
and U49606 (N_49606,N_47198,N_47547);
and U49607 (N_49607,N_46423,N_46952);
nand U49608 (N_49608,N_47269,N_47669);
xnor U49609 (N_49609,N_46829,N_46677);
or U49610 (N_49610,N_46724,N_47612);
and U49611 (N_49611,N_47839,N_47634);
or U49612 (N_49612,N_47922,N_47194);
nand U49613 (N_49613,N_47566,N_46963);
nor U49614 (N_49614,N_47655,N_47887);
or U49615 (N_49615,N_47395,N_47652);
xnor U49616 (N_49616,N_46885,N_46162);
xnor U49617 (N_49617,N_47562,N_46846);
nand U49618 (N_49618,N_46701,N_47523);
nand U49619 (N_49619,N_47816,N_47693);
xnor U49620 (N_49620,N_47601,N_46121);
or U49621 (N_49621,N_47302,N_46977);
xor U49622 (N_49622,N_47343,N_46559);
or U49623 (N_49623,N_46940,N_47712);
xnor U49624 (N_49624,N_47107,N_47112);
and U49625 (N_49625,N_46064,N_46825);
nor U49626 (N_49626,N_46838,N_47286);
nand U49627 (N_49627,N_47112,N_46183);
nor U49628 (N_49628,N_47643,N_47195);
nor U49629 (N_49629,N_47603,N_46482);
nand U49630 (N_49630,N_47862,N_46222);
nand U49631 (N_49631,N_47405,N_46497);
nor U49632 (N_49632,N_47966,N_47516);
nand U49633 (N_49633,N_46515,N_47959);
xor U49634 (N_49634,N_47157,N_47080);
or U49635 (N_49635,N_46455,N_47952);
nor U49636 (N_49636,N_46098,N_47445);
and U49637 (N_49637,N_46192,N_46333);
xor U49638 (N_49638,N_47913,N_46402);
nand U49639 (N_49639,N_47950,N_46090);
nand U49640 (N_49640,N_46936,N_46416);
nand U49641 (N_49641,N_46589,N_47997);
or U49642 (N_49642,N_47371,N_46209);
or U49643 (N_49643,N_46446,N_47765);
xor U49644 (N_49644,N_47379,N_46298);
nor U49645 (N_49645,N_47263,N_46189);
nor U49646 (N_49646,N_46840,N_47516);
xor U49647 (N_49647,N_46874,N_47294);
xor U49648 (N_49648,N_47673,N_47292);
xnor U49649 (N_49649,N_47050,N_46210);
or U49650 (N_49650,N_47237,N_46937);
xnor U49651 (N_49651,N_47203,N_46702);
nor U49652 (N_49652,N_47391,N_47372);
xor U49653 (N_49653,N_47772,N_47390);
xor U49654 (N_49654,N_46221,N_47771);
nand U49655 (N_49655,N_46928,N_46654);
xnor U49656 (N_49656,N_46209,N_47584);
and U49657 (N_49657,N_47664,N_47599);
and U49658 (N_49658,N_46662,N_46200);
and U49659 (N_49659,N_47203,N_47910);
nor U49660 (N_49660,N_46907,N_47348);
or U49661 (N_49661,N_47597,N_47972);
nand U49662 (N_49662,N_47447,N_47075);
nand U49663 (N_49663,N_47874,N_47423);
nand U49664 (N_49664,N_46555,N_47205);
xnor U49665 (N_49665,N_47662,N_46951);
xor U49666 (N_49666,N_46025,N_46081);
nand U49667 (N_49667,N_47721,N_47062);
xnor U49668 (N_49668,N_47980,N_46303);
nor U49669 (N_49669,N_46474,N_46355);
nand U49670 (N_49670,N_46402,N_46615);
nor U49671 (N_49671,N_47034,N_46627);
nor U49672 (N_49672,N_47752,N_46722);
nand U49673 (N_49673,N_47707,N_47223);
nor U49674 (N_49674,N_46556,N_47840);
and U49675 (N_49675,N_47992,N_47071);
xnor U49676 (N_49676,N_46927,N_47145);
xor U49677 (N_49677,N_47823,N_46169);
xnor U49678 (N_49678,N_46907,N_47520);
and U49679 (N_49679,N_47848,N_46657);
xnor U49680 (N_49680,N_46573,N_47797);
or U49681 (N_49681,N_47422,N_46583);
nor U49682 (N_49682,N_46848,N_46510);
or U49683 (N_49683,N_46343,N_46430);
xnor U49684 (N_49684,N_46148,N_46942);
xnor U49685 (N_49685,N_46837,N_46880);
or U49686 (N_49686,N_46808,N_46340);
nand U49687 (N_49687,N_46198,N_47521);
and U49688 (N_49688,N_46547,N_47708);
or U49689 (N_49689,N_47695,N_46076);
nand U49690 (N_49690,N_46734,N_47798);
nor U49691 (N_49691,N_47757,N_46074);
or U49692 (N_49692,N_47954,N_46956);
nor U49693 (N_49693,N_46213,N_46299);
xnor U49694 (N_49694,N_47053,N_47423);
nor U49695 (N_49695,N_46075,N_47782);
and U49696 (N_49696,N_47735,N_46944);
and U49697 (N_49697,N_47424,N_46125);
or U49698 (N_49698,N_46555,N_47551);
nand U49699 (N_49699,N_47425,N_47854);
and U49700 (N_49700,N_46738,N_47749);
nor U49701 (N_49701,N_46233,N_47373);
or U49702 (N_49702,N_47171,N_47624);
or U49703 (N_49703,N_47488,N_46298);
xnor U49704 (N_49704,N_47902,N_47289);
xor U49705 (N_49705,N_47116,N_46058);
xor U49706 (N_49706,N_47640,N_46344);
nor U49707 (N_49707,N_46513,N_47451);
nand U49708 (N_49708,N_47561,N_46841);
or U49709 (N_49709,N_47845,N_47793);
and U49710 (N_49710,N_47273,N_46331);
xor U49711 (N_49711,N_47682,N_47138);
xnor U49712 (N_49712,N_47178,N_47171);
xor U49713 (N_49713,N_47767,N_47033);
nor U49714 (N_49714,N_46248,N_46827);
nor U49715 (N_49715,N_47711,N_46894);
and U49716 (N_49716,N_46676,N_46273);
nand U49717 (N_49717,N_46125,N_46638);
xnor U49718 (N_49718,N_46029,N_46270);
and U49719 (N_49719,N_47739,N_47247);
nand U49720 (N_49720,N_47186,N_46991);
nand U49721 (N_49721,N_46443,N_47373);
nor U49722 (N_49722,N_46571,N_46072);
or U49723 (N_49723,N_46094,N_47023);
nand U49724 (N_49724,N_47642,N_46907);
and U49725 (N_49725,N_47727,N_47941);
and U49726 (N_49726,N_47093,N_46422);
nor U49727 (N_49727,N_46253,N_46010);
xor U49728 (N_49728,N_46801,N_46787);
or U49729 (N_49729,N_47257,N_47856);
nor U49730 (N_49730,N_46840,N_46330);
nor U49731 (N_49731,N_46325,N_47174);
nor U49732 (N_49732,N_47068,N_47664);
or U49733 (N_49733,N_46701,N_46386);
or U49734 (N_49734,N_46303,N_47348);
xor U49735 (N_49735,N_46452,N_47761);
xnor U49736 (N_49736,N_47406,N_46550);
or U49737 (N_49737,N_46491,N_47886);
xor U49738 (N_49738,N_47781,N_47638);
nor U49739 (N_49739,N_46253,N_46050);
nand U49740 (N_49740,N_46079,N_46320);
or U49741 (N_49741,N_47813,N_47426);
xor U49742 (N_49742,N_47641,N_47453);
or U49743 (N_49743,N_46413,N_46246);
nor U49744 (N_49744,N_47258,N_46245);
or U49745 (N_49745,N_46284,N_46894);
nor U49746 (N_49746,N_46530,N_46655);
nand U49747 (N_49747,N_46855,N_47294);
and U49748 (N_49748,N_47384,N_46712);
or U49749 (N_49749,N_46375,N_47382);
and U49750 (N_49750,N_47049,N_47750);
and U49751 (N_49751,N_46234,N_46958);
or U49752 (N_49752,N_47333,N_46924);
nand U49753 (N_49753,N_46368,N_46485);
nand U49754 (N_49754,N_46649,N_46847);
xnor U49755 (N_49755,N_46580,N_46867);
and U49756 (N_49756,N_46729,N_46547);
xnor U49757 (N_49757,N_47180,N_47692);
nand U49758 (N_49758,N_47490,N_46754);
or U49759 (N_49759,N_47300,N_47071);
or U49760 (N_49760,N_46968,N_47166);
xnor U49761 (N_49761,N_47029,N_47515);
or U49762 (N_49762,N_47364,N_47070);
or U49763 (N_49763,N_47783,N_47724);
xnor U49764 (N_49764,N_46555,N_47519);
and U49765 (N_49765,N_47777,N_47953);
and U49766 (N_49766,N_47479,N_46922);
or U49767 (N_49767,N_47757,N_46956);
nand U49768 (N_49768,N_46578,N_46975);
or U49769 (N_49769,N_47473,N_47629);
and U49770 (N_49770,N_46124,N_46576);
xnor U49771 (N_49771,N_46624,N_46962);
nor U49772 (N_49772,N_47713,N_46315);
xor U49773 (N_49773,N_47818,N_47696);
nand U49774 (N_49774,N_47879,N_47601);
or U49775 (N_49775,N_47369,N_47715);
and U49776 (N_49776,N_47511,N_47137);
nor U49777 (N_49777,N_46882,N_46428);
or U49778 (N_49778,N_47851,N_46619);
or U49779 (N_49779,N_47909,N_46342);
nor U49780 (N_49780,N_47854,N_46099);
nand U49781 (N_49781,N_46971,N_46532);
nor U49782 (N_49782,N_47294,N_46366);
and U49783 (N_49783,N_46752,N_46893);
nand U49784 (N_49784,N_47649,N_46259);
nor U49785 (N_49785,N_47706,N_46773);
nand U49786 (N_49786,N_47789,N_46011);
nand U49787 (N_49787,N_47545,N_47590);
nor U49788 (N_49788,N_47122,N_47588);
and U49789 (N_49789,N_46157,N_47578);
or U49790 (N_49790,N_46276,N_46268);
or U49791 (N_49791,N_46600,N_47869);
nand U49792 (N_49792,N_46630,N_47694);
and U49793 (N_49793,N_46514,N_46212);
nor U49794 (N_49794,N_47512,N_46069);
and U49795 (N_49795,N_47976,N_46872);
or U49796 (N_49796,N_46296,N_46512);
or U49797 (N_49797,N_46737,N_47173);
nand U49798 (N_49798,N_46111,N_46480);
or U49799 (N_49799,N_46278,N_47050);
and U49800 (N_49800,N_47398,N_47278);
or U49801 (N_49801,N_47681,N_47364);
nand U49802 (N_49802,N_46636,N_46331);
xnor U49803 (N_49803,N_47416,N_46472);
xnor U49804 (N_49804,N_46281,N_46844);
or U49805 (N_49805,N_47193,N_47422);
nand U49806 (N_49806,N_46061,N_46645);
xnor U49807 (N_49807,N_47950,N_46214);
or U49808 (N_49808,N_46455,N_47762);
xor U49809 (N_49809,N_46580,N_47002);
and U49810 (N_49810,N_46180,N_46605);
nor U49811 (N_49811,N_47035,N_46913);
nand U49812 (N_49812,N_47249,N_47474);
nand U49813 (N_49813,N_47987,N_47428);
nand U49814 (N_49814,N_47372,N_47030);
and U49815 (N_49815,N_47513,N_46576);
xnor U49816 (N_49816,N_46815,N_47050);
nor U49817 (N_49817,N_46101,N_47440);
and U49818 (N_49818,N_46472,N_46671);
and U49819 (N_49819,N_46740,N_46447);
and U49820 (N_49820,N_46545,N_47080);
or U49821 (N_49821,N_47191,N_46707);
nand U49822 (N_49822,N_47005,N_47533);
nor U49823 (N_49823,N_47194,N_46266);
or U49824 (N_49824,N_47683,N_46021);
nor U49825 (N_49825,N_47200,N_47524);
nor U49826 (N_49826,N_46468,N_46342);
nand U49827 (N_49827,N_46590,N_47316);
xor U49828 (N_49828,N_47787,N_46732);
nand U49829 (N_49829,N_46637,N_47926);
xnor U49830 (N_49830,N_47679,N_47079);
or U49831 (N_49831,N_46549,N_46005);
or U49832 (N_49832,N_47347,N_47287);
and U49833 (N_49833,N_47645,N_46756);
xnor U49834 (N_49834,N_47845,N_46561);
xnor U49835 (N_49835,N_47551,N_47437);
nor U49836 (N_49836,N_46099,N_46072);
or U49837 (N_49837,N_47731,N_47573);
nand U49838 (N_49838,N_47359,N_47431);
nor U49839 (N_49839,N_47150,N_47343);
or U49840 (N_49840,N_46170,N_47040);
nor U49841 (N_49841,N_47906,N_46148);
xnor U49842 (N_49842,N_47376,N_46359);
xor U49843 (N_49843,N_46277,N_47142);
nor U49844 (N_49844,N_47359,N_46924);
nor U49845 (N_49845,N_46247,N_46563);
xor U49846 (N_49846,N_46955,N_46972);
nand U49847 (N_49847,N_47843,N_46680);
or U49848 (N_49848,N_46487,N_47658);
nand U49849 (N_49849,N_46322,N_46728);
nor U49850 (N_49850,N_46218,N_46501);
and U49851 (N_49851,N_46539,N_47646);
xor U49852 (N_49852,N_46014,N_47198);
nand U49853 (N_49853,N_46414,N_46237);
nand U49854 (N_49854,N_46395,N_47199);
or U49855 (N_49855,N_46755,N_46942);
and U49856 (N_49856,N_47731,N_47779);
nor U49857 (N_49857,N_47769,N_47636);
nor U49858 (N_49858,N_46844,N_46541);
xnor U49859 (N_49859,N_46607,N_47908);
nand U49860 (N_49860,N_47105,N_46031);
xnor U49861 (N_49861,N_46718,N_47127);
or U49862 (N_49862,N_47278,N_46784);
xnor U49863 (N_49863,N_47468,N_47908);
nor U49864 (N_49864,N_46190,N_47133);
nor U49865 (N_49865,N_46178,N_46561);
nand U49866 (N_49866,N_46604,N_46053);
xnor U49867 (N_49867,N_46315,N_46005);
xnor U49868 (N_49868,N_47759,N_46652);
xnor U49869 (N_49869,N_46353,N_46276);
nand U49870 (N_49870,N_47200,N_47724);
nor U49871 (N_49871,N_46495,N_47914);
xnor U49872 (N_49872,N_46860,N_47705);
xor U49873 (N_49873,N_47859,N_46841);
nand U49874 (N_49874,N_46285,N_46905);
and U49875 (N_49875,N_46957,N_47711);
nand U49876 (N_49876,N_47179,N_47347);
or U49877 (N_49877,N_47275,N_46821);
nor U49878 (N_49878,N_47350,N_47309);
xnor U49879 (N_49879,N_47886,N_47541);
nor U49880 (N_49880,N_47612,N_46681);
nand U49881 (N_49881,N_47481,N_46501);
nor U49882 (N_49882,N_46128,N_47376);
and U49883 (N_49883,N_46101,N_46356);
nor U49884 (N_49884,N_46390,N_47881);
nor U49885 (N_49885,N_46342,N_46329);
nand U49886 (N_49886,N_47800,N_46665);
or U49887 (N_49887,N_47133,N_47094);
nand U49888 (N_49888,N_47961,N_47245);
or U49889 (N_49889,N_47291,N_47959);
nor U49890 (N_49890,N_46973,N_47032);
or U49891 (N_49891,N_47520,N_47869);
nand U49892 (N_49892,N_46980,N_47127);
or U49893 (N_49893,N_47382,N_47280);
nand U49894 (N_49894,N_47829,N_46626);
and U49895 (N_49895,N_46105,N_47941);
nand U49896 (N_49896,N_46536,N_46177);
nor U49897 (N_49897,N_46858,N_47106);
and U49898 (N_49898,N_47111,N_47171);
and U49899 (N_49899,N_46160,N_47863);
and U49900 (N_49900,N_46074,N_46832);
nand U49901 (N_49901,N_46914,N_47767);
or U49902 (N_49902,N_47916,N_46986);
nor U49903 (N_49903,N_46677,N_47286);
nor U49904 (N_49904,N_47317,N_46653);
and U49905 (N_49905,N_47093,N_46700);
nand U49906 (N_49906,N_46771,N_46689);
nor U49907 (N_49907,N_47528,N_47901);
and U49908 (N_49908,N_47717,N_46930);
xnor U49909 (N_49909,N_46272,N_46930);
and U49910 (N_49910,N_46945,N_46333);
or U49911 (N_49911,N_47001,N_46825);
or U49912 (N_49912,N_46676,N_47489);
nand U49913 (N_49913,N_46076,N_47603);
xnor U49914 (N_49914,N_46546,N_46534);
nand U49915 (N_49915,N_47670,N_46331);
nand U49916 (N_49916,N_46186,N_46974);
or U49917 (N_49917,N_46295,N_47344);
or U49918 (N_49918,N_47759,N_46206);
nand U49919 (N_49919,N_46107,N_47132);
nor U49920 (N_49920,N_46438,N_47139);
or U49921 (N_49921,N_46225,N_47438);
and U49922 (N_49922,N_46059,N_47529);
or U49923 (N_49923,N_47045,N_47901);
and U49924 (N_49924,N_46680,N_46436);
nor U49925 (N_49925,N_47174,N_46303);
nor U49926 (N_49926,N_47398,N_46012);
nand U49927 (N_49927,N_47365,N_47768);
xor U49928 (N_49928,N_47439,N_47423);
xnor U49929 (N_49929,N_47753,N_47848);
xnor U49930 (N_49930,N_47535,N_47279);
or U49931 (N_49931,N_46125,N_47764);
nand U49932 (N_49932,N_46796,N_46641);
or U49933 (N_49933,N_46784,N_46431);
xor U49934 (N_49934,N_47877,N_46413);
nand U49935 (N_49935,N_47575,N_46481);
nand U49936 (N_49936,N_46762,N_47338);
xnor U49937 (N_49937,N_46282,N_46363);
or U49938 (N_49938,N_46184,N_47984);
nand U49939 (N_49939,N_47491,N_46773);
and U49940 (N_49940,N_46023,N_46674);
and U49941 (N_49941,N_46374,N_47850);
nand U49942 (N_49942,N_46950,N_46621);
and U49943 (N_49943,N_47406,N_47959);
and U49944 (N_49944,N_47301,N_47134);
and U49945 (N_49945,N_46341,N_46815);
nand U49946 (N_49946,N_46958,N_46138);
and U49947 (N_49947,N_46828,N_47039);
and U49948 (N_49948,N_47102,N_47289);
or U49949 (N_49949,N_46489,N_47632);
or U49950 (N_49950,N_46373,N_46425);
xnor U49951 (N_49951,N_46443,N_47312);
and U49952 (N_49952,N_46301,N_47094);
nand U49953 (N_49953,N_47551,N_47029);
xnor U49954 (N_49954,N_46309,N_47164);
and U49955 (N_49955,N_46422,N_46160);
xor U49956 (N_49956,N_46643,N_47958);
xnor U49957 (N_49957,N_47640,N_47596);
nand U49958 (N_49958,N_47971,N_47836);
nand U49959 (N_49959,N_46616,N_46130);
and U49960 (N_49960,N_46955,N_46591);
and U49961 (N_49961,N_47222,N_47064);
nand U49962 (N_49962,N_46241,N_46274);
nand U49963 (N_49963,N_47639,N_47297);
nor U49964 (N_49964,N_47895,N_46403);
or U49965 (N_49965,N_46553,N_47178);
xor U49966 (N_49966,N_47136,N_46752);
nor U49967 (N_49967,N_47840,N_46925);
or U49968 (N_49968,N_47200,N_47511);
xnor U49969 (N_49969,N_47439,N_47553);
nand U49970 (N_49970,N_47492,N_46349);
or U49971 (N_49971,N_46131,N_46069);
or U49972 (N_49972,N_46837,N_47876);
nor U49973 (N_49973,N_46044,N_46815);
nand U49974 (N_49974,N_47268,N_46669);
nor U49975 (N_49975,N_46949,N_46234);
nor U49976 (N_49976,N_47880,N_47504);
or U49977 (N_49977,N_47383,N_47424);
nor U49978 (N_49978,N_47902,N_47612);
nor U49979 (N_49979,N_46436,N_46627);
nor U49980 (N_49980,N_46357,N_47721);
nand U49981 (N_49981,N_46571,N_47301);
xnor U49982 (N_49982,N_46886,N_46680);
and U49983 (N_49983,N_47829,N_47595);
xor U49984 (N_49984,N_46078,N_46823);
xnor U49985 (N_49985,N_46149,N_47246);
and U49986 (N_49986,N_47927,N_46669);
nand U49987 (N_49987,N_46404,N_46790);
nor U49988 (N_49988,N_46710,N_46867);
and U49989 (N_49989,N_47167,N_47170);
or U49990 (N_49990,N_46764,N_46282);
or U49991 (N_49991,N_47394,N_46125);
nor U49992 (N_49992,N_46889,N_46713);
xor U49993 (N_49993,N_47304,N_46559);
xor U49994 (N_49994,N_47835,N_47913);
xnor U49995 (N_49995,N_47143,N_46817);
and U49996 (N_49996,N_46885,N_46666);
nor U49997 (N_49997,N_46384,N_47212);
nor U49998 (N_49998,N_47789,N_46531);
and U49999 (N_49999,N_47707,N_46573);
or UO_0 (O_0,N_48184,N_49763);
or UO_1 (O_1,N_48925,N_49550);
xnor UO_2 (O_2,N_48927,N_49357);
and UO_3 (O_3,N_48391,N_49923);
and UO_4 (O_4,N_49999,N_48257);
nor UO_5 (O_5,N_48756,N_49842);
xor UO_6 (O_6,N_49782,N_48906);
or UO_7 (O_7,N_49257,N_49616);
and UO_8 (O_8,N_48804,N_48339);
or UO_9 (O_9,N_48643,N_48626);
or UO_10 (O_10,N_48381,N_49491);
nor UO_11 (O_11,N_49530,N_49803);
nand UO_12 (O_12,N_49986,N_49844);
and UO_13 (O_13,N_48870,N_48053);
and UO_14 (O_14,N_49266,N_48664);
or UO_15 (O_15,N_49663,N_48075);
xnor UO_16 (O_16,N_49374,N_49811);
or UO_17 (O_17,N_48665,N_49454);
nor UO_18 (O_18,N_49768,N_48002);
and UO_19 (O_19,N_48742,N_49890);
xnor UO_20 (O_20,N_48315,N_49035);
and UO_21 (O_21,N_49958,N_49916);
or UO_22 (O_22,N_48644,N_48486);
nor UO_23 (O_23,N_49444,N_48966);
nor UO_24 (O_24,N_49242,N_49697);
nand UO_25 (O_25,N_48316,N_49073);
xor UO_26 (O_26,N_48885,N_49928);
nand UO_27 (O_27,N_48780,N_49812);
nor UO_28 (O_28,N_49148,N_49282);
or UO_29 (O_29,N_49941,N_48960);
xor UO_30 (O_30,N_49533,N_48671);
and UO_31 (O_31,N_49887,N_48303);
nor UO_32 (O_32,N_49818,N_48089);
or UO_33 (O_33,N_49336,N_49070);
and UO_34 (O_34,N_48628,N_48731);
nor UO_35 (O_35,N_49370,N_49171);
nand UO_36 (O_36,N_48956,N_49784);
nor UO_37 (O_37,N_49541,N_48692);
xor UO_38 (O_38,N_49447,N_48313);
xor UO_39 (O_39,N_48173,N_49824);
nor UO_40 (O_40,N_49553,N_49211);
nor UO_41 (O_41,N_49959,N_48368);
xnor UO_42 (O_42,N_48565,N_48761);
nor UO_43 (O_43,N_49639,N_48524);
or UO_44 (O_44,N_49421,N_49854);
nand UO_45 (O_45,N_49201,N_49097);
nor UO_46 (O_46,N_48485,N_48588);
nor UO_47 (O_47,N_49267,N_49919);
xor UO_48 (O_48,N_49861,N_49415);
and UO_49 (O_49,N_49482,N_48146);
and UO_50 (O_50,N_49858,N_49046);
nor UO_51 (O_51,N_49290,N_49284);
xnor UO_52 (O_52,N_49412,N_49004);
or UO_53 (O_53,N_48504,N_49310);
xor UO_54 (O_54,N_49321,N_48129);
xor UO_55 (O_55,N_49126,N_49566);
xor UO_56 (O_56,N_49124,N_49892);
or UO_57 (O_57,N_48225,N_49876);
xnor UO_58 (O_58,N_49921,N_48206);
and UO_59 (O_59,N_49857,N_48943);
nand UO_60 (O_60,N_48387,N_49484);
or UO_61 (O_61,N_49413,N_48957);
xor UO_62 (O_62,N_49728,N_49625);
nor UO_63 (O_63,N_49390,N_49689);
nor UO_64 (O_64,N_48685,N_49723);
and UO_65 (O_65,N_49260,N_48564);
or UO_66 (O_66,N_49508,N_48152);
xnor UO_67 (O_67,N_48690,N_49925);
nand UO_68 (O_68,N_48520,N_49078);
xnor UO_69 (O_69,N_49951,N_48868);
nor UO_70 (O_70,N_49236,N_49081);
xor UO_71 (O_71,N_49462,N_48069);
and UO_72 (O_72,N_49702,N_48730);
nor UO_73 (O_73,N_49871,N_49957);
nor UO_74 (O_74,N_49044,N_49250);
and UO_75 (O_75,N_48041,N_48077);
or UO_76 (O_76,N_49439,N_49608);
nand UO_77 (O_77,N_48662,N_49855);
and UO_78 (O_78,N_49375,N_48229);
and UO_79 (O_79,N_49518,N_48603);
nand UO_80 (O_80,N_48784,N_49688);
nand UO_81 (O_81,N_49934,N_48170);
or UO_82 (O_82,N_48047,N_48156);
or UO_83 (O_83,N_48113,N_48670);
nor UO_84 (O_84,N_48490,N_48590);
and UO_85 (O_85,N_48970,N_49547);
xor UO_86 (O_86,N_49975,N_49036);
and UO_87 (O_87,N_48085,N_48620);
and UO_88 (O_88,N_48306,N_48634);
and UO_89 (O_89,N_49781,N_49752);
nand UO_90 (O_90,N_48031,N_48509);
nor UO_91 (O_91,N_48890,N_49993);
or UO_92 (O_92,N_49299,N_48540);
xor UO_93 (O_93,N_48648,N_49833);
nor UO_94 (O_94,N_48572,N_49516);
xor UO_95 (O_95,N_48379,N_49886);
xnor UO_96 (O_96,N_48724,N_48618);
nor UO_97 (O_97,N_48500,N_49604);
xnor UO_98 (O_98,N_48232,N_49438);
or UO_99 (O_99,N_49806,N_49182);
nor UO_100 (O_100,N_48439,N_48120);
and UO_101 (O_101,N_48076,N_48808);
xnor UO_102 (O_102,N_48998,N_48298);
nand UO_103 (O_103,N_49234,N_49636);
or UO_104 (O_104,N_49387,N_49634);
nor UO_105 (O_105,N_48897,N_48760);
nor UO_106 (O_106,N_49903,N_48332);
nand UO_107 (O_107,N_48973,N_49402);
nor UO_108 (O_108,N_49393,N_48932);
nand UO_109 (O_109,N_48445,N_48281);
or UO_110 (O_110,N_48096,N_48362);
or UO_111 (O_111,N_49762,N_49346);
or UO_112 (O_112,N_48062,N_49076);
nor UO_113 (O_113,N_49621,N_49622);
xor UO_114 (O_114,N_49092,N_48452);
or UO_115 (O_115,N_49796,N_49511);
or UO_116 (O_116,N_49361,N_48659);
nand UO_117 (O_117,N_48043,N_49667);
and UO_118 (O_118,N_48848,N_48050);
or UO_119 (O_119,N_48242,N_49713);
nand UO_120 (O_120,N_48811,N_49584);
or UO_121 (O_121,N_48916,N_49388);
or UO_122 (O_122,N_49660,N_49365);
nor UO_123 (O_123,N_48460,N_48866);
nor UO_124 (O_124,N_48834,N_48978);
nand UO_125 (O_125,N_48674,N_48488);
xor UO_126 (O_126,N_48483,N_49990);
or UO_127 (O_127,N_49258,N_48678);
or UO_128 (O_128,N_48243,N_49397);
nand UO_129 (O_129,N_49896,N_49265);
nor UO_130 (O_130,N_49938,N_49263);
or UO_131 (O_131,N_48398,N_48657);
and UO_132 (O_132,N_49683,N_48934);
nor UO_133 (O_133,N_48975,N_49061);
nor UO_134 (O_134,N_49253,N_48860);
or UO_135 (O_135,N_48449,N_48568);
nor UO_136 (O_136,N_49481,N_48142);
and UO_137 (O_137,N_49411,N_49316);
nor UO_138 (O_138,N_48376,N_48613);
xor UO_139 (O_139,N_49955,N_48884);
or UO_140 (O_140,N_48974,N_48616);
nor UO_141 (O_141,N_48933,N_49731);
nand UO_142 (O_142,N_48841,N_48244);
nand UO_143 (O_143,N_48738,N_48091);
or UO_144 (O_144,N_48570,N_48723);
nor UO_145 (O_145,N_49757,N_49449);
nand UO_146 (O_146,N_49554,N_49488);
nor UO_147 (O_147,N_49870,N_49213);
nor UO_148 (O_148,N_49074,N_49527);
nand UO_149 (O_149,N_48030,N_48915);
nand UO_150 (O_150,N_48382,N_48319);
nor UO_151 (O_151,N_49270,N_49297);
or UO_152 (O_152,N_48487,N_49730);
nand UO_153 (O_153,N_48755,N_49973);
nor UO_154 (O_154,N_49602,N_48917);
and UO_155 (O_155,N_49807,N_49232);
nor UO_156 (O_156,N_49269,N_48873);
nand UO_157 (O_157,N_49948,N_49820);
xor UO_158 (O_158,N_49256,N_49565);
nand UO_159 (O_159,N_48631,N_49804);
and UO_160 (O_160,N_48469,N_48880);
xor UO_161 (O_161,N_48743,N_48965);
and UO_162 (O_162,N_48849,N_49588);
xor UO_163 (O_163,N_49669,N_49308);
and UO_164 (O_164,N_48431,N_48250);
or UO_165 (O_165,N_49909,N_49254);
or UO_166 (O_166,N_48102,N_49718);
nor UO_167 (O_167,N_49240,N_48337);
or UO_168 (O_168,N_49889,N_48856);
nor UO_169 (O_169,N_48324,N_49027);
nand UO_170 (O_170,N_48872,N_49740);
xor UO_171 (O_171,N_49430,N_48370);
xnor UO_172 (O_172,N_49012,N_48832);
xnor UO_173 (O_173,N_49332,N_48419);
nor UO_174 (O_174,N_48611,N_49726);
nor UO_175 (O_175,N_48165,N_49897);
or UO_176 (O_176,N_48167,N_48058);
or UO_177 (O_177,N_49272,N_48991);
xor UO_178 (O_178,N_49817,N_49335);
nand UO_179 (O_179,N_48428,N_48843);
nand UO_180 (O_180,N_48412,N_49091);
and UO_181 (O_181,N_49274,N_49991);
xnor UO_182 (O_182,N_49230,N_48175);
or UO_183 (O_183,N_49144,N_48942);
nor UO_184 (O_184,N_49868,N_49159);
nor UO_185 (O_185,N_48435,N_48100);
nor UO_186 (O_186,N_48793,N_49408);
and UO_187 (O_187,N_49156,N_48852);
xnor UO_188 (O_188,N_48189,N_48846);
and UO_189 (O_189,N_49347,N_49245);
or UO_190 (O_190,N_48208,N_48740);
nand UO_191 (O_191,N_49984,N_48327);
and UO_192 (O_192,N_48171,N_49377);
or UO_193 (O_193,N_49798,N_48499);
and UO_194 (O_194,N_48360,N_49135);
or UO_195 (O_195,N_49102,N_48065);
xor UO_196 (O_196,N_48317,N_49138);
and UO_197 (O_197,N_48702,N_48335);
nor UO_198 (O_198,N_48402,N_49312);
nor UO_199 (O_199,N_49536,N_48624);
or UO_200 (O_200,N_49523,N_48747);
xnor UO_201 (O_201,N_49017,N_48087);
or UO_202 (O_202,N_48253,N_48106);
nor UO_203 (O_203,N_48677,N_48092);
nand UO_204 (O_204,N_48645,N_49205);
xor UO_205 (O_205,N_48931,N_48116);
xnor UO_206 (O_206,N_49195,N_48254);
and UO_207 (O_207,N_49400,N_48221);
nor UO_208 (O_208,N_48961,N_48114);
nor UO_209 (O_209,N_49980,N_48049);
or UO_210 (O_210,N_48413,N_49594);
nand UO_211 (O_211,N_48821,N_48256);
and UO_212 (O_212,N_48967,N_49985);
nor UO_213 (O_213,N_49560,N_49732);
and UO_214 (O_214,N_48018,N_49895);
xor UO_215 (O_215,N_48223,N_48894);
or UO_216 (O_216,N_49741,N_48700);
and UO_217 (O_217,N_48004,N_48022);
xor UO_218 (O_218,N_48105,N_49907);
nand UO_219 (O_219,N_48132,N_49847);
xnor UO_220 (O_220,N_48727,N_48517);
and UO_221 (O_221,N_49943,N_48796);
nor UO_222 (O_222,N_48433,N_49598);
nor UO_223 (O_223,N_49268,N_48667);
and UO_224 (O_224,N_49545,N_48656);
nand UO_225 (O_225,N_49194,N_49303);
nor UO_226 (O_226,N_49829,N_48660);
xnor UO_227 (O_227,N_48212,N_48734);
nand UO_228 (O_228,N_48981,N_48163);
xnor UO_229 (O_229,N_49600,N_48078);
or UO_230 (O_230,N_49132,N_48086);
xnor UO_231 (O_231,N_49926,N_48371);
and UO_232 (O_232,N_48014,N_49341);
and UO_233 (O_233,N_48591,N_49678);
xor UO_234 (O_234,N_48573,N_48307);
and UO_235 (O_235,N_48814,N_48627);
xor UO_236 (O_236,N_48513,N_48533);
nor UO_237 (O_237,N_48385,N_48501);
xnor UO_238 (O_238,N_48125,N_48815);
nand UO_239 (O_239,N_48145,N_48782);
and UO_240 (O_240,N_48394,N_49040);
nor UO_241 (O_241,N_48080,N_49404);
xnor UO_242 (O_242,N_48340,N_49152);
nand UO_243 (O_243,N_48987,N_48825);
and UO_244 (O_244,N_49662,N_48265);
nor UO_245 (O_245,N_48448,N_48422);
and UO_246 (O_246,N_49932,N_49627);
nand UO_247 (O_247,N_48630,N_49682);
xnor UO_248 (O_248,N_48952,N_49771);
xnor UO_249 (O_249,N_48023,N_49499);
and UO_250 (O_250,N_49154,N_48876);
nor UO_251 (O_251,N_49434,N_49472);
xnor UO_252 (O_252,N_48800,N_49995);
xnor UO_253 (O_253,N_48118,N_48141);
or UO_254 (O_254,N_49416,N_49770);
nor UO_255 (O_255,N_48705,N_48709);
or UO_256 (O_256,N_49106,N_48123);
xor UO_257 (O_257,N_48473,N_48838);
or UO_258 (O_258,N_48712,N_49134);
or UO_259 (O_259,N_48928,N_49637);
nand UO_260 (O_260,N_49789,N_48126);
xnor UO_261 (O_261,N_49239,N_49930);
or UO_262 (O_262,N_48465,N_49165);
or UO_263 (O_263,N_48632,N_48638);
and UO_264 (O_264,N_49203,N_49657);
nor UO_265 (O_265,N_48836,N_48230);
xnor UO_266 (O_266,N_48548,N_48110);
or UO_267 (O_267,N_49304,N_49425);
xnor UO_268 (O_268,N_49087,N_49243);
xnor UO_269 (O_269,N_49317,N_48680);
xnor UO_270 (O_270,N_48929,N_48331);
or UO_271 (O_271,N_49799,N_48607);
nor UO_272 (O_272,N_49210,N_48646);
nor UO_273 (O_273,N_48482,N_48720);
nor UO_274 (O_274,N_49215,N_48012);
and UO_275 (O_275,N_49681,N_48149);
xnor UO_276 (O_276,N_48356,N_49075);
nand UO_277 (O_277,N_48877,N_49071);
nand UO_278 (O_278,N_48429,N_49121);
nand UO_279 (O_279,N_49917,N_49822);
nand UO_280 (O_280,N_48071,N_49721);
and UO_281 (O_281,N_48283,N_48423);
or UO_282 (O_282,N_49456,N_49575);
xor UO_283 (O_283,N_48322,N_49675);
nand UO_284 (O_284,N_48357,N_48920);
nor UO_285 (O_285,N_48308,N_49451);
or UO_286 (O_286,N_48652,N_49694);
nor UO_287 (O_287,N_49352,N_48042);
nor UO_288 (O_288,N_49275,N_49733);
nor UO_289 (O_289,N_48336,N_48693);
or UO_290 (O_290,N_49028,N_49853);
or UO_291 (O_291,N_49661,N_48701);
nand UO_292 (O_292,N_49725,N_48893);
nor UO_293 (O_293,N_49107,N_49793);
nand UO_294 (O_294,N_49248,N_49504);
nor UO_295 (O_295,N_48179,N_49389);
nand UO_296 (O_296,N_49922,N_48910);
nand UO_297 (O_297,N_49836,N_48599);
xor UO_298 (O_298,N_49231,N_49698);
xnor UO_299 (O_299,N_48434,N_49173);
and UO_300 (O_300,N_48426,N_49734);
and UO_301 (O_301,N_49291,N_49947);
nand UO_302 (O_302,N_49143,N_48831);
or UO_303 (O_303,N_49997,N_49176);
nor UO_304 (O_304,N_49724,N_48268);
nor UO_305 (O_305,N_49739,N_49477);
xor UO_306 (O_306,N_49116,N_48299);
nor UO_307 (O_307,N_49761,N_49368);
or UO_308 (O_308,N_48468,N_48200);
nand UO_309 (O_309,N_48919,N_49181);
and UO_310 (O_310,N_48397,N_49615);
xor UO_311 (O_311,N_48502,N_49406);
nor UO_312 (O_312,N_48844,N_48380);
xor UO_313 (O_313,N_48081,N_49571);
xor UO_314 (O_314,N_49348,N_49618);
xor UO_315 (O_315,N_48577,N_49470);
and UO_316 (O_316,N_48177,N_48421);
nor UO_317 (O_317,N_48668,N_49570);
and UO_318 (O_318,N_48217,N_49431);
and UO_319 (O_319,N_48914,N_48054);
nor UO_320 (O_320,N_49160,N_48450);
or UO_321 (O_321,N_48204,N_48569);
nand UO_322 (O_322,N_48290,N_48036);
xor UO_323 (O_323,N_49830,N_49577);
or UO_324 (O_324,N_49561,N_49048);
or UO_325 (O_325,N_49340,N_49020);
and UO_326 (O_326,N_49880,N_49183);
nand UO_327 (O_327,N_49384,N_49506);
or UO_328 (O_328,N_49302,N_48990);
or UO_329 (O_329,N_49300,N_49515);
or UO_330 (O_330,N_49283,N_48545);
or UO_331 (O_331,N_49791,N_49151);
nor UO_332 (O_332,N_49949,N_48222);
xor UO_333 (O_333,N_48555,N_49816);
nand UO_334 (O_334,N_49095,N_49502);
xor UO_335 (O_335,N_48194,N_48608);
or UO_336 (O_336,N_48311,N_49202);
xnor UO_337 (O_337,N_48072,N_49041);
or UO_338 (O_338,N_48378,N_49053);
nand UO_339 (O_339,N_48561,N_49869);
nor UO_340 (O_340,N_48689,N_49845);
nand UO_341 (O_341,N_49631,N_48532);
nor UO_342 (O_342,N_48822,N_48805);
nand UO_343 (O_343,N_48140,N_49133);
nand UO_344 (O_344,N_49542,N_48629);
and UO_345 (O_345,N_49950,N_49100);
nor UO_346 (O_346,N_48048,N_49805);
or UO_347 (O_347,N_49420,N_49819);
or UO_348 (O_348,N_49517,N_49326);
or UO_349 (O_349,N_48348,N_49687);
and UO_350 (O_350,N_48249,N_48586);
or UO_351 (O_351,N_49096,N_49380);
or UO_352 (O_352,N_49077,N_48017);
and UO_353 (O_353,N_48228,N_49422);
and UO_354 (O_354,N_49360,N_49356);
xor UO_355 (O_355,N_49426,N_48637);
nor UO_356 (O_356,N_48640,N_48850);
and UO_357 (O_357,N_48959,N_49177);
nand UO_358 (O_358,N_48539,N_48136);
nor UO_359 (O_359,N_48526,N_48489);
nor UO_360 (O_360,N_48898,N_48737);
and UO_361 (O_361,N_49052,N_49480);
or UO_362 (O_362,N_49666,N_48055);
nand UO_363 (O_363,N_48409,N_49318);
or UO_364 (O_364,N_49686,N_49611);
nor UO_365 (O_365,N_48079,N_49395);
xnor UO_366 (O_366,N_49136,N_49503);
or UO_367 (O_367,N_49277,N_49204);
nor UO_368 (O_368,N_48016,N_49825);
xor UO_369 (O_369,N_48295,N_49872);
xor UO_370 (O_370,N_48158,N_48766);
and UO_371 (O_371,N_48205,N_49748);
nand UO_372 (O_372,N_48006,N_48277);
and UO_373 (O_373,N_49742,N_48716);
and UO_374 (O_374,N_49787,N_49716);
nor UO_375 (O_375,N_48459,N_49437);
and UO_376 (O_376,N_48466,N_48013);
or UO_377 (O_377,N_48736,N_48606);
and UO_378 (O_378,N_48993,N_49963);
or UO_379 (O_379,N_48111,N_48550);
nand UO_380 (O_380,N_49163,N_48771);
nand UO_381 (O_381,N_49717,N_49207);
nor UO_382 (O_382,N_49864,N_49605);
nor UO_383 (O_383,N_48183,N_48563);
xor UO_384 (O_384,N_48270,N_49241);
nand UO_385 (O_385,N_48726,N_49585);
and UO_386 (O_386,N_48134,N_48829);
xnor UO_387 (O_387,N_48887,N_48444);
xnor UO_388 (O_388,N_49228,N_48349);
and UO_389 (O_389,N_49233,N_49802);
and UO_390 (O_390,N_49122,N_49493);
xor UO_391 (O_391,N_48647,N_49601);
nor UO_392 (O_392,N_48447,N_48262);
or UO_393 (O_393,N_48571,N_48024);
or UO_394 (O_394,N_48816,N_48739);
and UO_395 (O_395,N_48554,N_48455);
nand UO_396 (O_396,N_49089,N_49051);
nor UO_397 (O_397,N_48227,N_48128);
and UO_398 (O_398,N_48478,N_49131);
nand UO_399 (O_399,N_48777,N_48625);
nor UO_400 (O_400,N_48273,N_49305);
and UO_401 (O_401,N_48681,N_48301);
or UO_402 (O_402,N_48330,N_48699);
and UO_403 (O_403,N_48538,N_48430);
and UO_404 (O_404,N_49823,N_49767);
and UO_405 (O_405,N_49330,N_48708);
and UO_406 (O_406,N_48003,N_49405);
nand UO_407 (O_407,N_48574,N_48279);
or UO_408 (O_408,N_48992,N_48264);
xor UO_409 (O_409,N_48878,N_48786);
xor UO_410 (O_410,N_48009,N_49010);
and UO_411 (O_411,N_49313,N_49252);
xnor UO_412 (O_412,N_49821,N_49946);
or UO_413 (O_413,N_49883,N_49744);
nor UO_414 (O_414,N_48521,N_48365);
and UO_415 (O_415,N_48476,N_49129);
nand UO_416 (O_416,N_49125,N_48903);
xnor UO_417 (O_417,N_49031,N_49019);
or UO_418 (O_418,N_48187,N_48542);
nand UO_419 (O_419,N_49727,N_49063);
and UO_420 (O_420,N_49196,N_49496);
xnor UO_421 (O_421,N_49647,N_48735);
or UO_422 (O_422,N_48781,N_49485);
or UO_423 (O_423,N_49358,N_48663);
nand UO_424 (O_424,N_49712,N_48988);
nand UO_425 (O_425,N_48040,N_49200);
and UO_426 (O_426,N_48060,N_48185);
xnor UO_427 (O_427,N_49677,N_49746);
xor UO_428 (O_428,N_48896,N_49766);
xor UO_429 (O_429,N_49112,N_48669);
and UO_430 (O_430,N_48168,N_48425);
nand UO_431 (O_431,N_48010,N_49756);
nor UO_432 (O_432,N_49902,N_49068);
nor UO_433 (O_433,N_48122,N_48345);
xor UO_434 (O_434,N_48581,N_49815);
or UO_435 (O_435,N_48790,N_48220);
nand UO_436 (O_436,N_49906,N_48686);
and UO_437 (O_437,N_48839,N_49015);
nand UO_438 (O_438,N_48984,N_49064);
nor UO_439 (O_439,N_48810,N_48964);
nor UO_440 (O_440,N_48911,N_49996);
or UO_441 (O_441,N_49994,N_48101);
and UO_442 (O_442,N_48936,N_49952);
xnor UO_443 (O_443,N_49033,N_49414);
nand UO_444 (O_444,N_49054,N_48779);
and UO_445 (O_445,N_49977,N_49128);
or UO_446 (O_446,N_48722,N_49140);
nand UO_447 (O_447,N_48698,N_48395);
xnor UO_448 (O_448,N_48234,N_48057);
or UO_449 (O_449,N_49337,N_49497);
xnor UO_450 (O_450,N_49987,N_49433);
nand UO_451 (O_451,N_48121,N_49610);
and UO_452 (O_452,N_48666,N_48763);
nor UO_453 (O_453,N_48713,N_48366);
xnor UO_454 (O_454,N_48178,N_48696);
xor UO_455 (O_455,N_48600,N_48117);
xor UO_456 (O_456,N_48405,N_48192);
and UO_457 (O_457,N_49684,N_48480);
nand UO_458 (O_458,N_49954,N_49057);
xor UO_459 (O_459,N_49953,N_49262);
or UO_460 (O_460,N_48037,N_48494);
nand UO_461 (O_461,N_48715,N_48704);
nor UO_462 (O_462,N_49008,N_49372);
nor UO_463 (O_463,N_49664,N_48551);
nor UO_464 (O_464,N_48847,N_48442);
nand UO_465 (O_465,N_49379,N_48237);
nand UO_466 (O_466,N_49198,N_48462);
xnor UO_467 (O_467,N_48605,N_49220);
nor UO_468 (O_468,N_49016,N_48641);
nand UO_469 (O_469,N_49155,N_49624);
xor UO_470 (O_470,N_48310,N_49632);
nand UO_471 (O_471,N_48567,N_49164);
nand UO_472 (O_472,N_49882,N_48056);
nor UO_473 (O_473,N_48963,N_48246);
xnor UO_474 (O_474,N_49924,N_49557);
and UO_475 (O_475,N_49099,N_49276);
or UO_476 (O_476,N_48675,N_48828);
xor UO_477 (O_477,N_49696,N_49371);
or UO_478 (O_478,N_48694,N_49369);
or UO_479 (O_479,N_48383,N_48437);
or UO_480 (O_480,N_48744,N_49311);
nor UO_481 (O_481,N_48097,N_49510);
xnor UO_482 (O_482,N_49777,N_49080);
and UO_483 (O_483,N_48131,N_48995);
and UO_484 (O_484,N_48809,N_48417);
and UO_485 (O_485,N_48388,N_48706);
xor UO_486 (O_486,N_49877,N_49025);
nor UO_487 (O_487,N_49323,N_48214);
nor UO_488 (O_488,N_49178,N_49736);
or UO_489 (O_489,N_48239,N_48635);
nand UO_490 (O_490,N_48374,N_49069);
xor UO_491 (O_491,N_48610,N_49193);
nor UO_492 (O_492,N_49797,N_48944);
nor UO_493 (O_493,N_48070,N_49778);
and UO_494 (O_494,N_49592,N_49349);
nor UO_495 (O_495,N_49559,N_48682);
xor UO_496 (O_496,N_49676,N_49385);
nor UO_497 (O_497,N_49441,N_48748);
nor UO_498 (O_498,N_48045,N_49966);
xor UO_499 (O_499,N_49982,N_49759);
xor UO_500 (O_500,N_48935,N_49586);
nor UO_501 (O_501,N_49720,N_49013);
or UO_502 (O_502,N_48438,N_48358);
nand UO_503 (O_503,N_48350,N_49968);
nand UO_504 (O_504,N_49247,N_48410);
xnor UO_505 (O_505,N_48019,N_49794);
or UO_506 (O_506,N_48725,N_49514);
xnor UO_507 (O_507,N_49229,N_49988);
xor UO_508 (O_508,N_49264,N_48552);
xnor UO_509 (O_509,N_49613,N_49001);
nand UO_510 (O_510,N_49603,N_48046);
and UO_511 (O_511,N_49281,N_49185);
nor UO_512 (O_512,N_48464,N_48575);
xor UO_513 (O_513,N_48457,N_48549);
xnor UO_514 (O_514,N_48719,N_48874);
or UO_515 (O_515,N_49538,N_48946);
and UO_516 (O_516,N_48553,N_49137);
or UO_517 (O_517,N_48593,N_48688);
and UO_518 (O_518,N_48446,N_48636);
nor UO_519 (O_519,N_48424,N_49322);
nor UO_520 (O_520,N_49319,N_49735);
nand UO_521 (O_521,N_48389,N_49094);
xnor UO_522 (O_522,N_49353,N_48066);
xor UO_523 (O_523,N_48236,N_49307);
and UO_524 (O_524,N_49226,N_49293);
nand UO_525 (O_525,N_49055,N_49118);
and UO_526 (O_526,N_48139,N_48980);
or UO_527 (O_527,N_48443,N_48661);
or UO_528 (O_528,N_48164,N_49117);
or UO_529 (O_529,N_48093,N_49826);
or UO_530 (O_530,N_48812,N_49428);
or UO_531 (O_531,N_48939,N_49900);
and UO_532 (O_532,N_48979,N_48757);
or UO_533 (O_533,N_48354,N_48458);
nand UO_534 (O_534,N_48359,N_48255);
nand UO_535 (O_535,N_49446,N_48619);
nand UO_536 (O_536,N_49644,N_48393);
or UO_537 (O_537,N_49249,N_49309);
and UO_538 (O_538,N_48304,N_49544);
xor UO_539 (O_539,N_49929,N_49668);
xnor UO_540 (O_540,N_48456,N_49674);
nand UO_541 (O_541,N_49672,N_48785);
xor UO_542 (O_542,N_48404,N_49945);
and UO_543 (O_543,N_48147,N_48601);
nand UO_544 (O_544,N_48203,N_48717);
nor UO_545 (O_545,N_49933,N_49255);
or UO_546 (O_546,N_48986,N_48506);
nor UO_547 (O_547,N_49227,N_48400);
and UO_548 (O_548,N_48733,N_49655);
nor UO_549 (O_549,N_49525,N_49329);
nor UO_550 (O_550,N_48515,N_48186);
nand UO_551 (O_551,N_49715,N_48518);
xor UO_552 (O_552,N_49620,N_49813);
nor UO_553 (O_553,N_49537,N_49745);
nor UO_554 (O_554,N_49753,N_48598);
xor UO_555 (O_555,N_49120,N_49827);
nand UO_556 (O_556,N_48021,N_49920);
xor UO_557 (O_557,N_49992,N_49429);
nor UO_558 (O_558,N_48094,N_48000);
nor UO_559 (O_559,N_48044,N_48157);
or UO_560 (O_560,N_48921,N_48369);
nand UO_561 (O_561,N_49168,N_48653);
or UO_562 (O_562,N_49614,N_49520);
or UO_563 (O_563,N_48495,N_49567);
nor UO_564 (O_564,N_48259,N_48767);
nor UO_565 (O_565,N_48913,N_48769);
and UO_566 (O_566,N_49795,N_49381);
nand UO_567 (O_567,N_48875,N_48213);
or UO_568 (O_568,N_49695,N_48231);
xor UO_569 (O_569,N_48900,N_49539);
and UO_570 (O_570,N_49528,N_48818);
xnor UO_571 (O_571,N_49574,N_48248);
xnor UO_572 (O_572,N_49366,N_48454);
xnor UO_573 (O_573,N_48557,N_49692);
nor UO_574 (O_574,N_48436,N_48193);
nor UO_575 (O_575,N_49750,N_49640);
nand UO_576 (O_576,N_49259,N_48714);
or UO_577 (O_577,N_49800,N_48161);
xor UO_578 (O_578,N_49314,N_48902);
nand UO_579 (O_579,N_49908,N_48516);
and UO_580 (O_580,N_48883,N_48758);
nand UO_581 (O_581,N_48827,N_49500);
nor UO_582 (O_582,N_48160,N_48399);
nor UO_583 (O_583,N_48280,N_48741);
and UO_584 (O_584,N_48658,N_49860);
xnor UO_585 (O_585,N_49765,N_48059);
xnor UO_586 (O_586,N_49540,N_49841);
and UO_587 (O_587,N_49467,N_49532);
nor UO_588 (O_588,N_48621,N_49912);
nor UO_589 (O_589,N_48418,N_49214);
and UO_590 (O_590,N_48289,N_48302);
xor UO_591 (O_591,N_49056,N_49442);
xor UO_592 (O_592,N_49543,N_49161);
nor UO_593 (O_593,N_48288,N_49364);
or UO_594 (O_594,N_49261,N_48240);
xnor UO_595 (O_595,N_48088,N_48034);
or UO_596 (O_596,N_49331,N_48245);
nand UO_597 (O_597,N_48005,N_48924);
nor UO_598 (O_598,N_49505,N_49840);
and UO_599 (O_599,N_49376,N_49749);
nand UO_600 (O_600,N_48612,N_48067);
nand UO_601 (O_601,N_48833,N_48511);
nand UO_602 (O_602,N_49737,N_49453);
and UO_603 (O_603,N_49223,N_49478);
nor UO_604 (O_604,N_48566,N_48342);
xor UO_605 (O_605,N_49788,N_49396);
or UO_606 (O_606,N_49866,N_49979);
nor UO_607 (O_607,N_48174,N_49172);
nor UO_608 (O_608,N_49961,N_49835);
xor UO_609 (O_609,N_49382,N_49848);
or UO_610 (O_610,N_49865,N_49832);
nand UO_611 (O_611,N_48218,N_49058);
xnor UO_612 (O_612,N_49572,N_49246);
nand UO_613 (O_613,N_49179,N_48226);
nand UO_614 (O_614,N_49351,N_48353);
and UO_615 (O_615,N_48527,N_48084);
or UO_616 (O_616,N_48823,N_49512);
nor UO_617 (O_617,N_48474,N_48143);
nand UO_618 (O_618,N_48795,N_49549);
nand UO_619 (O_619,N_49021,N_49555);
nor UO_620 (O_620,N_48751,N_49489);
and UO_621 (O_621,N_48461,N_48895);
and UO_622 (O_622,N_48558,N_49427);
or UO_623 (O_623,N_48416,N_48746);
nand UO_624 (O_624,N_48127,N_49479);
and UO_625 (O_625,N_49563,N_49710);
xor UO_626 (O_626,N_48938,N_49189);
nor UO_627 (O_627,N_49251,N_49108);
and UO_628 (O_628,N_48510,N_48453);
or UO_629 (O_629,N_48528,N_48219);
or UO_630 (O_630,N_48503,N_48854);
nor UO_631 (O_631,N_49005,N_49967);
or UO_632 (O_632,N_48862,N_48820);
nor UO_633 (O_633,N_49894,N_49911);
xnor UO_634 (O_634,N_48655,N_48241);
nand UO_635 (O_635,N_49838,N_48074);
nor UO_636 (O_636,N_49939,N_49568);
xor UO_637 (O_637,N_48364,N_48772);
nor UO_638 (O_638,N_48144,N_49315);
and UO_639 (O_639,N_49589,N_49719);
or UO_640 (O_640,N_48562,N_48377);
or UO_641 (O_641,N_49130,N_48901);
and UO_642 (O_642,N_49964,N_49045);
xnor UO_643 (O_643,N_49111,N_49881);
nor UO_644 (O_644,N_48801,N_49700);
and UO_645 (O_645,N_49670,N_48314);
nand UO_646 (O_646,N_49591,N_49551);
xnor UO_647 (O_647,N_49628,N_48033);
or UO_648 (O_648,N_48420,N_48291);
and UO_649 (O_649,N_48276,N_49150);
nor UO_650 (O_650,N_49754,N_48320);
or UO_651 (O_651,N_49651,N_48971);
nand UO_652 (O_652,N_48806,N_49237);
nand UO_653 (O_653,N_48972,N_48803);
and UO_654 (O_654,N_48032,N_48765);
or UO_655 (O_655,N_49018,N_49363);
nand UO_656 (O_656,N_48325,N_49654);
xor UO_657 (O_657,N_48064,N_48813);
and UO_658 (O_658,N_49652,N_48355);
nand UO_659 (O_659,N_49507,N_48198);
nand UO_660 (O_660,N_49956,N_49050);
xnor UO_661 (O_661,N_49535,N_48347);
and UO_662 (O_662,N_48926,N_49587);
and UO_663 (O_663,N_48863,N_49286);
nand UO_664 (O_664,N_48718,N_49901);
nor UO_665 (O_665,N_48587,N_48266);
nor UO_666 (O_666,N_48729,N_48026);
nand UO_667 (O_667,N_48284,N_49110);
and UO_668 (O_668,N_49524,N_49184);
xor UO_669 (O_669,N_49162,N_48776);
nor UO_670 (O_670,N_49888,N_49435);
nand UO_671 (O_671,N_49709,N_49287);
and UO_672 (O_672,N_48798,N_48797);
or UO_673 (O_673,N_48305,N_48817);
nor UO_674 (O_674,N_48497,N_48543);
nand UO_675 (O_675,N_49659,N_49597);
nand UO_676 (O_676,N_49146,N_49022);
nand UO_677 (O_677,N_48498,N_49473);
or UO_678 (O_678,N_49219,N_48985);
and UO_679 (O_679,N_49452,N_48775);
or UO_680 (O_680,N_49474,N_48753);
and UO_681 (O_681,N_48233,N_49086);
nor UO_682 (O_682,N_49007,N_48650);
and UO_683 (O_683,N_49606,N_48799);
and UO_684 (O_684,N_49609,N_49301);
or UO_685 (O_685,N_49190,N_48602);
and UO_686 (O_686,N_49612,N_48432);
or UO_687 (O_687,N_49115,N_48861);
nor UO_688 (O_688,N_49918,N_48754);
xnor UO_689 (O_689,N_48989,N_48169);
nor UO_690 (O_690,N_48061,N_48479);
or UO_691 (O_691,N_49775,N_49082);
or UO_692 (O_692,N_48930,N_49169);
and UO_693 (O_693,N_48341,N_48541);
and UO_694 (O_694,N_48247,N_49101);
and UO_695 (O_695,N_49373,N_48773);
nand UO_696 (O_696,N_49852,N_49225);
and UO_697 (O_697,N_48293,N_48215);
or UO_698 (O_698,N_49023,N_49216);
and UO_699 (O_699,N_48099,N_49448);
nor UO_700 (O_700,N_48386,N_49362);
nand UO_701 (O_701,N_49738,N_49450);
or UO_702 (O_702,N_48275,N_49898);
nor UO_703 (O_703,N_48840,N_48063);
nor UO_704 (O_704,N_49685,N_49417);
nor UO_705 (O_705,N_48585,N_48615);
and UO_706 (O_706,N_49690,N_49656);
and UO_707 (O_707,N_48326,N_49079);
nand UO_708 (O_708,N_48560,N_49529);
nand UO_709 (O_709,N_48869,N_48762);
nand UO_710 (O_710,N_49208,N_49521);
and UO_711 (O_711,N_48683,N_49774);
nor UO_712 (O_712,N_49810,N_48372);
nor UO_713 (O_713,N_48507,N_49940);
or UO_714 (O_714,N_49047,N_49893);
nand UO_715 (O_715,N_48951,N_49471);
and UO_716 (O_716,N_49333,N_49937);
xnor UO_717 (O_717,N_48604,N_49339);
xnor UO_718 (O_718,N_48020,N_48352);
or UO_719 (O_719,N_48830,N_49199);
and UO_720 (O_720,N_48403,N_49649);
xnor UO_721 (O_721,N_49648,N_48082);
or UO_722 (O_722,N_49714,N_48576);
nand UO_723 (O_723,N_48115,N_48982);
and UO_724 (O_724,N_49552,N_48904);
nand UO_725 (O_725,N_49147,N_49187);
or UO_726 (O_726,N_48802,N_49546);
and UO_727 (O_727,N_49722,N_49843);
xnor UO_728 (O_728,N_48344,N_49065);
and UO_729 (O_729,N_49424,N_48710);
xnor UO_730 (O_730,N_49180,N_48864);
and UO_731 (O_731,N_48949,N_48296);
nor UO_732 (O_732,N_48039,N_48285);
nor UO_733 (O_733,N_49418,N_49809);
and UO_734 (O_734,N_49875,N_49706);
or UO_735 (O_735,N_49490,N_48819);
nand UO_736 (O_736,N_49878,N_48211);
xor UO_737 (O_737,N_49145,N_49186);
nor UO_738 (O_738,N_48791,N_48589);
nor UO_739 (O_739,N_49032,N_48639);
nand UO_740 (O_740,N_49109,N_48038);
or UO_741 (O_741,N_49786,N_48977);
nor UO_742 (O_742,N_48475,N_49392);
xor UO_743 (O_743,N_48768,N_49910);
or UO_744 (O_744,N_49519,N_48764);
xnor UO_745 (O_745,N_48789,N_49465);
nor UO_746 (O_746,N_48098,N_49776);
or UO_747 (O_747,N_48871,N_48287);
and UO_748 (O_748,N_48544,N_48835);
xor UO_749 (O_749,N_48937,N_49167);
or UO_750 (O_750,N_49222,N_49289);
nor UO_751 (O_751,N_49142,N_49935);
nand UO_752 (O_752,N_48559,N_49711);
or UO_753 (O_753,N_48375,N_49970);
and UO_754 (O_754,N_49969,N_48649);
and UO_755 (O_755,N_48535,N_48414);
and UO_756 (O_756,N_48300,N_49494);
and UO_757 (O_757,N_49378,N_49244);
and UO_758 (O_758,N_49679,N_48642);
nand UO_759 (O_759,N_48531,N_48492);
xor UO_760 (O_760,N_49285,N_48962);
and UO_761 (O_761,N_49629,N_48857);
and UO_762 (O_762,N_48481,N_48969);
or UO_763 (O_763,N_49891,N_49067);
or UO_764 (O_764,N_48137,N_48401);
and UO_765 (O_765,N_48051,N_48108);
nand UO_766 (O_766,N_49403,N_49899);
nand UO_767 (O_767,N_49399,N_49801);
and UO_768 (O_768,N_48886,N_49849);
or UO_769 (O_769,N_48623,N_49083);
and UO_770 (O_770,N_49665,N_48338);
nor UO_771 (O_771,N_48679,N_48858);
nand UO_772 (O_772,N_48373,N_49296);
nand UO_773 (O_773,N_49831,N_49562);
and UO_774 (O_774,N_49011,N_49394);
and UO_775 (O_775,N_49905,N_49641);
nand UO_776 (O_776,N_48519,N_49170);
and UO_777 (O_777,N_49703,N_48888);
xnor UO_778 (O_778,N_48155,N_49599);
nand UO_779 (O_779,N_49037,N_48274);
xor UO_780 (O_780,N_49976,N_48787);
and UO_781 (O_781,N_48191,N_49139);
nand UO_782 (O_782,N_49873,N_49014);
and UO_783 (O_783,N_49278,N_48508);
or UO_784 (O_784,N_49009,N_49105);
or UO_785 (O_785,N_49582,N_49059);
and UO_786 (O_786,N_48721,N_48728);
nor UO_787 (O_787,N_48103,N_48073);
xnor UO_788 (O_788,N_49209,N_49217);
nand UO_789 (O_789,N_48826,N_49461);
nor UO_790 (O_790,N_48750,N_49534);
xor UO_791 (O_791,N_49850,N_49280);
nand UO_792 (O_792,N_48684,N_49743);
xor UO_793 (O_793,N_48711,N_48238);
nor UO_794 (O_794,N_49084,N_49295);
nor UO_795 (O_795,N_49062,N_48090);
xnor UO_796 (O_796,N_48530,N_48529);
nand UO_797 (O_797,N_48367,N_49680);
or UO_798 (O_798,N_49558,N_48028);
or UO_799 (O_799,N_48783,N_48609);
or UO_800 (O_800,N_49328,N_49464);
xor UO_801 (O_801,N_48505,N_48008);
nor UO_802 (O_802,N_49114,N_48950);
and UO_803 (O_803,N_48881,N_49707);
and UO_804 (O_804,N_49191,N_49034);
xnor UO_805 (O_805,N_49492,N_48584);
xor UO_806 (O_806,N_49407,N_48891);
or UO_807 (O_807,N_48011,N_49792);
nor UO_808 (O_808,N_48889,N_49635);
nor UO_809 (O_809,N_48968,N_48536);
nand UO_810 (O_810,N_48522,N_48778);
nor UO_811 (O_811,N_48133,N_49344);
or UO_812 (O_812,N_49814,N_48029);
and UO_813 (O_813,N_49221,N_48472);
and UO_814 (O_814,N_49699,N_48384);
nor UO_815 (O_815,N_48899,N_49174);
nand UO_816 (O_816,N_49391,N_48035);
nand UO_817 (O_817,N_49457,N_49779);
xnor UO_818 (O_818,N_49638,N_48470);
xor UO_819 (O_819,N_48001,N_49175);
or UO_820 (O_820,N_48788,N_48673);
and UO_821 (O_821,N_49513,N_48958);
xor UO_822 (O_822,N_48210,N_48484);
or UO_823 (O_823,N_49595,N_48135);
xor UO_824 (O_824,N_48580,N_49747);
nor UO_825 (O_825,N_48537,N_49000);
xor UO_826 (O_826,N_48297,N_49483);
nor UO_827 (O_827,N_49874,N_49780);
nor UO_828 (O_828,N_48216,N_48622);
nand UO_829 (O_829,N_49410,N_48390);
nor UO_830 (O_830,N_49522,N_49026);
and UO_831 (O_831,N_49642,N_49188);
nand UO_832 (O_832,N_48309,N_48351);
nor UO_833 (O_833,N_48408,N_48851);
xnor UO_834 (O_834,N_49630,N_49834);
xor UO_835 (O_835,N_49701,N_49072);
nor UO_836 (O_836,N_48909,N_49856);
nand UO_837 (O_837,N_49808,N_49235);
xnor UO_838 (O_838,N_48329,N_49650);
or UO_839 (O_839,N_48853,N_48427);
nor UO_840 (O_840,N_49783,N_48148);
and UO_841 (O_841,N_49583,N_49192);
nor UO_842 (O_842,N_49760,N_49944);
nor UO_843 (O_843,N_48282,N_48271);
nand UO_844 (O_844,N_49419,N_48286);
or UO_845 (O_845,N_48124,N_49927);
or UO_846 (O_846,N_48119,N_48321);
nor UO_847 (O_847,N_49342,N_49093);
nand UO_848 (O_848,N_48947,N_48007);
nor UO_849 (O_849,N_49633,N_48415);
nor UO_850 (O_850,N_48107,N_48837);
nor UO_851 (O_851,N_49367,N_49158);
xnor UO_852 (O_852,N_48263,N_49043);
nor UO_853 (O_853,N_49960,N_49607);
xnor UO_854 (O_854,N_48199,N_48441);
or UO_855 (O_855,N_48583,N_49623);
nand UO_856 (O_856,N_48770,N_48083);
and UO_857 (O_857,N_48252,N_48278);
nand UO_858 (O_858,N_49501,N_49460);
xor UO_859 (O_859,N_48467,N_48407);
nor UO_860 (O_860,N_49576,N_49693);
or UO_861 (O_861,N_49306,N_49383);
and UO_862 (O_862,N_48859,N_49863);
nand UO_863 (O_863,N_49002,N_49708);
xnor UO_864 (O_864,N_49981,N_48406);
xnor UO_865 (O_865,N_49088,N_49153);
and UO_866 (O_866,N_49673,N_48151);
nand UO_867 (O_867,N_49704,N_48202);
or UO_868 (O_868,N_48251,N_48922);
and UO_869 (O_869,N_49617,N_48824);
nor UO_870 (O_870,N_48312,N_48188);
and UO_871 (O_871,N_49024,N_48676);
nand UO_872 (O_872,N_49113,N_48579);
nand UO_873 (O_873,N_49913,N_48556);
nand UO_874 (O_874,N_48687,N_49166);
nand UO_875 (O_875,N_49790,N_48451);
nor UO_876 (O_876,N_49334,N_48794);
or UO_877 (O_877,N_49978,N_48945);
nand UO_878 (O_878,N_48343,N_48166);
or UO_879 (O_879,N_48130,N_48491);
nor UO_880 (O_880,N_49455,N_48855);
nand UO_881 (O_881,N_49458,N_48842);
xor UO_882 (O_882,N_48918,N_48865);
xor UO_883 (O_883,N_48015,N_49619);
nand UO_884 (O_884,N_48845,N_49355);
or UO_885 (O_885,N_49936,N_49974);
nor UO_886 (O_886,N_48333,N_49409);
xor UO_887 (O_887,N_49596,N_49038);
xor UO_888 (O_888,N_48109,N_49556);
nor UO_889 (O_889,N_49862,N_49066);
nand UO_890 (O_890,N_49548,N_48633);
nand UO_891 (O_891,N_48209,N_49729);
or UO_892 (O_892,N_49915,N_49646);
xnor UO_893 (O_893,N_49769,N_49049);
and UO_894 (O_894,N_48534,N_49751);
nand UO_895 (O_895,N_48905,N_49580);
or UO_896 (O_896,N_48578,N_48912);
nand UO_897 (O_897,N_48954,N_48703);
and UO_898 (O_898,N_48154,N_48594);
or UO_899 (O_899,N_49931,N_49298);
nand UO_900 (O_900,N_48392,N_48292);
or UO_901 (O_901,N_49867,N_49495);
or UO_902 (O_902,N_48867,N_48159);
xnor UO_903 (O_903,N_49772,N_49294);
nand UO_904 (O_904,N_48272,N_49962);
nor UO_905 (O_905,N_48260,N_48190);
nor UO_906 (O_906,N_48651,N_49042);
nand UO_907 (O_907,N_49119,N_49324);
nor UO_908 (O_908,N_49658,N_48411);
xnor UO_909 (O_909,N_48025,N_48150);
or UO_910 (O_910,N_48294,N_49060);
nand UO_911 (O_911,N_48672,N_48752);
nand UO_912 (O_912,N_48176,N_49773);
or UO_913 (O_913,N_49320,N_49197);
xor UO_914 (O_914,N_49645,N_49104);
xnor UO_915 (O_915,N_48172,N_49581);
or UO_916 (O_916,N_48471,N_49764);
xor UO_917 (O_917,N_49983,N_48983);
xor UO_918 (O_918,N_49029,N_48807);
xnor UO_919 (O_919,N_48224,N_48095);
nor UO_920 (O_920,N_49498,N_49879);
nor UO_921 (O_921,N_48104,N_49218);
nand UO_922 (O_922,N_48953,N_49443);
or UO_923 (O_923,N_49030,N_49423);
xnor UO_924 (O_924,N_49755,N_49965);
and UO_925 (O_925,N_49475,N_49564);
nor UO_926 (O_926,N_48361,N_48201);
and UO_927 (O_927,N_48614,N_49149);
xnor UO_928 (O_928,N_48976,N_49238);
or UO_929 (O_929,N_49003,N_48523);
and UO_930 (O_930,N_48695,N_48879);
nor UO_931 (O_931,N_48597,N_49359);
nor UO_932 (O_932,N_48948,N_48749);
nand UO_933 (O_933,N_48617,N_48180);
xnor UO_934 (O_934,N_48182,N_48907);
or UO_935 (O_935,N_49141,N_48068);
and UO_936 (O_936,N_48496,N_49123);
and UO_937 (O_937,N_49466,N_49338);
nand UO_938 (O_938,N_48654,N_48052);
nor UO_939 (O_939,N_49469,N_48745);
nand UO_940 (O_940,N_49224,N_48514);
or UO_941 (O_941,N_48196,N_48346);
nor UO_942 (O_942,N_48892,N_49098);
and UO_943 (O_943,N_48908,N_48112);
nor UO_944 (O_944,N_49445,N_49885);
and UO_945 (O_945,N_49345,N_49705);
xnor UO_946 (O_946,N_48162,N_48195);
and UO_947 (O_947,N_48396,N_49593);
nor UO_948 (O_948,N_49271,N_48547);
nand UO_949 (O_949,N_48267,N_49487);
nor UO_950 (O_950,N_49526,N_48546);
nand UO_951 (O_951,N_48996,N_49432);
xnor UO_952 (O_952,N_48440,N_48269);
xor UO_953 (O_953,N_49859,N_48235);
xnor UO_954 (O_954,N_49989,N_49343);
xnor UO_955 (O_955,N_48595,N_48334);
or UO_956 (O_956,N_48940,N_49006);
or UO_957 (O_957,N_49085,N_49292);
nor UO_958 (O_958,N_49998,N_49386);
or UO_959 (O_959,N_48955,N_48697);
nand UO_960 (O_960,N_48323,N_49884);
nor UO_961 (O_961,N_49350,N_48318);
xnor UO_962 (O_962,N_48363,N_49288);
nand UO_963 (O_963,N_48512,N_49643);
nor UO_964 (O_964,N_49914,N_48882);
and UO_965 (O_965,N_49436,N_48261);
nand UO_966 (O_966,N_48463,N_49463);
and UO_967 (O_967,N_49157,N_48759);
xor UO_968 (O_968,N_49785,N_49828);
nand UO_969 (O_969,N_49354,N_49401);
and UO_970 (O_970,N_48596,N_49206);
or UO_971 (O_971,N_49578,N_48027);
xnor UO_972 (O_972,N_49839,N_49579);
nand UO_973 (O_973,N_49626,N_48582);
and UO_974 (O_974,N_49590,N_48941);
and UO_975 (O_975,N_48732,N_48207);
xnor UO_976 (O_976,N_48997,N_48493);
nand UO_977 (O_977,N_48707,N_49971);
nor UO_978 (O_978,N_49212,N_48153);
and UO_979 (O_979,N_48592,N_49327);
or UO_980 (O_980,N_48994,N_48923);
nor UO_981 (O_981,N_49531,N_49573);
and UO_982 (O_982,N_49846,N_49090);
nand UO_983 (O_983,N_49837,N_49671);
and UO_984 (O_984,N_49273,N_49509);
nor UO_985 (O_985,N_49476,N_48477);
and UO_986 (O_986,N_49103,N_49972);
nand UO_987 (O_987,N_48691,N_49459);
xor UO_988 (O_988,N_49904,N_48138);
and UO_989 (O_989,N_48525,N_49758);
and UO_990 (O_990,N_49486,N_49127);
nor UO_991 (O_991,N_49440,N_49398);
or UO_992 (O_992,N_49851,N_49325);
or UO_993 (O_993,N_49468,N_48792);
xor UO_994 (O_994,N_48999,N_49942);
nor UO_995 (O_995,N_49279,N_49691);
nor UO_996 (O_996,N_48774,N_48197);
nand UO_997 (O_997,N_49039,N_48181);
or UO_998 (O_998,N_48328,N_49653);
nor UO_999 (O_999,N_49569,N_48258);
nor UO_1000 (O_1000,N_48455,N_49280);
xor UO_1001 (O_1001,N_49003,N_48755);
xnor UO_1002 (O_1002,N_49606,N_49674);
and UO_1003 (O_1003,N_49350,N_49903);
and UO_1004 (O_1004,N_49274,N_49682);
and UO_1005 (O_1005,N_48388,N_49146);
or UO_1006 (O_1006,N_48779,N_49486);
and UO_1007 (O_1007,N_48499,N_48036);
and UO_1008 (O_1008,N_49065,N_49550);
nor UO_1009 (O_1009,N_48089,N_49399);
nor UO_1010 (O_1010,N_48089,N_48750);
xnor UO_1011 (O_1011,N_48521,N_49652);
nor UO_1012 (O_1012,N_48141,N_49759);
and UO_1013 (O_1013,N_49976,N_49028);
xnor UO_1014 (O_1014,N_49318,N_49818);
or UO_1015 (O_1015,N_49252,N_48918);
and UO_1016 (O_1016,N_48236,N_49573);
nand UO_1017 (O_1017,N_49270,N_49462);
and UO_1018 (O_1018,N_48733,N_49661);
or UO_1019 (O_1019,N_48079,N_49546);
or UO_1020 (O_1020,N_48834,N_48095);
nor UO_1021 (O_1021,N_49140,N_49469);
nand UO_1022 (O_1022,N_49049,N_48013);
and UO_1023 (O_1023,N_48316,N_48591);
xnor UO_1024 (O_1024,N_49169,N_49705);
xor UO_1025 (O_1025,N_49658,N_49142);
nor UO_1026 (O_1026,N_48368,N_49888);
and UO_1027 (O_1027,N_49904,N_48069);
xnor UO_1028 (O_1028,N_48384,N_48253);
nand UO_1029 (O_1029,N_49870,N_49295);
xnor UO_1030 (O_1030,N_48064,N_49660);
nand UO_1031 (O_1031,N_49028,N_48037);
or UO_1032 (O_1032,N_49099,N_49952);
xnor UO_1033 (O_1033,N_48868,N_49263);
or UO_1034 (O_1034,N_48551,N_48052);
and UO_1035 (O_1035,N_48571,N_48237);
and UO_1036 (O_1036,N_48883,N_49122);
nor UO_1037 (O_1037,N_48867,N_49346);
nor UO_1038 (O_1038,N_49014,N_49641);
xor UO_1039 (O_1039,N_48984,N_48777);
and UO_1040 (O_1040,N_49855,N_48760);
nand UO_1041 (O_1041,N_49289,N_48449);
xnor UO_1042 (O_1042,N_48878,N_49030);
or UO_1043 (O_1043,N_48921,N_48031);
nand UO_1044 (O_1044,N_48348,N_49597);
nand UO_1045 (O_1045,N_49462,N_48650);
or UO_1046 (O_1046,N_48363,N_48243);
or UO_1047 (O_1047,N_48424,N_48170);
or UO_1048 (O_1048,N_48678,N_49083);
nor UO_1049 (O_1049,N_49164,N_49678);
or UO_1050 (O_1050,N_48670,N_49477);
and UO_1051 (O_1051,N_49628,N_48546);
xnor UO_1052 (O_1052,N_48188,N_48195);
nand UO_1053 (O_1053,N_48057,N_49665);
and UO_1054 (O_1054,N_48348,N_48693);
nor UO_1055 (O_1055,N_49643,N_49895);
xnor UO_1056 (O_1056,N_49566,N_48743);
xor UO_1057 (O_1057,N_49064,N_48491);
nand UO_1058 (O_1058,N_48571,N_48360);
nor UO_1059 (O_1059,N_49089,N_48133);
or UO_1060 (O_1060,N_49050,N_48770);
nand UO_1061 (O_1061,N_49143,N_49295);
nand UO_1062 (O_1062,N_48254,N_49738);
and UO_1063 (O_1063,N_49931,N_48987);
and UO_1064 (O_1064,N_48852,N_48464);
nand UO_1065 (O_1065,N_48109,N_48567);
nor UO_1066 (O_1066,N_48550,N_49159);
nor UO_1067 (O_1067,N_48013,N_49283);
or UO_1068 (O_1068,N_48417,N_49941);
and UO_1069 (O_1069,N_49518,N_49790);
nor UO_1070 (O_1070,N_49474,N_49591);
and UO_1071 (O_1071,N_48727,N_49734);
nor UO_1072 (O_1072,N_49302,N_48491);
nand UO_1073 (O_1073,N_49900,N_48733);
nor UO_1074 (O_1074,N_48248,N_48883);
and UO_1075 (O_1075,N_49541,N_49180);
or UO_1076 (O_1076,N_49580,N_48546);
xnor UO_1077 (O_1077,N_48105,N_49678);
and UO_1078 (O_1078,N_48975,N_49900);
nor UO_1079 (O_1079,N_49314,N_49394);
nor UO_1080 (O_1080,N_49104,N_49718);
or UO_1081 (O_1081,N_49370,N_49132);
or UO_1082 (O_1082,N_48460,N_48858);
xor UO_1083 (O_1083,N_48572,N_49384);
xor UO_1084 (O_1084,N_49399,N_48601);
xnor UO_1085 (O_1085,N_49703,N_49932);
nor UO_1086 (O_1086,N_49891,N_49992);
nand UO_1087 (O_1087,N_49696,N_49421);
or UO_1088 (O_1088,N_48100,N_49433);
nor UO_1089 (O_1089,N_49056,N_48217);
and UO_1090 (O_1090,N_49422,N_49995);
nor UO_1091 (O_1091,N_48937,N_49876);
nand UO_1092 (O_1092,N_48267,N_49560);
nor UO_1093 (O_1093,N_48678,N_49519);
nand UO_1094 (O_1094,N_48432,N_49593);
and UO_1095 (O_1095,N_48476,N_49397);
nor UO_1096 (O_1096,N_48792,N_48869);
or UO_1097 (O_1097,N_48569,N_48991);
nand UO_1098 (O_1098,N_49339,N_49903);
and UO_1099 (O_1099,N_49077,N_49788);
nor UO_1100 (O_1100,N_49712,N_48010);
nand UO_1101 (O_1101,N_49193,N_48489);
xor UO_1102 (O_1102,N_49691,N_48350);
nor UO_1103 (O_1103,N_48942,N_48672);
or UO_1104 (O_1104,N_48317,N_48228);
or UO_1105 (O_1105,N_48131,N_49786);
nor UO_1106 (O_1106,N_48962,N_48035);
nand UO_1107 (O_1107,N_49895,N_48731);
and UO_1108 (O_1108,N_49249,N_49401);
nor UO_1109 (O_1109,N_48029,N_49220);
or UO_1110 (O_1110,N_49801,N_49326);
nor UO_1111 (O_1111,N_49041,N_48280);
or UO_1112 (O_1112,N_49956,N_49965);
xnor UO_1113 (O_1113,N_49266,N_48268);
nand UO_1114 (O_1114,N_48271,N_49065);
xor UO_1115 (O_1115,N_49755,N_49597);
and UO_1116 (O_1116,N_49324,N_49798);
nor UO_1117 (O_1117,N_48349,N_48566);
nand UO_1118 (O_1118,N_48942,N_49515);
nor UO_1119 (O_1119,N_49397,N_48669);
xnor UO_1120 (O_1120,N_48630,N_48743);
xor UO_1121 (O_1121,N_49704,N_49150);
or UO_1122 (O_1122,N_48005,N_48300);
or UO_1123 (O_1123,N_48207,N_49813);
xor UO_1124 (O_1124,N_49506,N_49441);
and UO_1125 (O_1125,N_49498,N_49258);
nand UO_1126 (O_1126,N_48114,N_48031);
and UO_1127 (O_1127,N_49996,N_48353);
nand UO_1128 (O_1128,N_49242,N_49033);
or UO_1129 (O_1129,N_49178,N_48873);
nand UO_1130 (O_1130,N_49506,N_49931);
nand UO_1131 (O_1131,N_48918,N_48522);
nor UO_1132 (O_1132,N_49963,N_48039);
nor UO_1133 (O_1133,N_48511,N_48405);
and UO_1134 (O_1134,N_48813,N_49802);
and UO_1135 (O_1135,N_48947,N_48989);
and UO_1136 (O_1136,N_49919,N_49177);
or UO_1137 (O_1137,N_49136,N_48822);
nand UO_1138 (O_1138,N_48812,N_48493);
nand UO_1139 (O_1139,N_48608,N_48289);
nor UO_1140 (O_1140,N_48493,N_48749);
and UO_1141 (O_1141,N_48262,N_48716);
and UO_1142 (O_1142,N_49082,N_49003);
or UO_1143 (O_1143,N_49324,N_48812);
nand UO_1144 (O_1144,N_48364,N_49599);
xor UO_1145 (O_1145,N_49299,N_49264);
xnor UO_1146 (O_1146,N_48616,N_48576);
and UO_1147 (O_1147,N_49174,N_48399);
xor UO_1148 (O_1148,N_49791,N_48756);
or UO_1149 (O_1149,N_49615,N_49446);
xnor UO_1150 (O_1150,N_48400,N_49642);
or UO_1151 (O_1151,N_48488,N_48234);
nor UO_1152 (O_1152,N_49967,N_48548);
nor UO_1153 (O_1153,N_49198,N_49197);
xor UO_1154 (O_1154,N_49389,N_49717);
or UO_1155 (O_1155,N_49658,N_49581);
nor UO_1156 (O_1156,N_48352,N_48131);
and UO_1157 (O_1157,N_49388,N_49851);
and UO_1158 (O_1158,N_48943,N_49394);
and UO_1159 (O_1159,N_49462,N_49001);
xor UO_1160 (O_1160,N_49429,N_49088);
xor UO_1161 (O_1161,N_49146,N_49502);
or UO_1162 (O_1162,N_49508,N_49243);
nand UO_1163 (O_1163,N_48677,N_49209);
and UO_1164 (O_1164,N_49035,N_49813);
xor UO_1165 (O_1165,N_49508,N_49937);
or UO_1166 (O_1166,N_48979,N_49873);
and UO_1167 (O_1167,N_48953,N_49746);
nor UO_1168 (O_1168,N_48401,N_48381);
or UO_1169 (O_1169,N_48285,N_48913);
nand UO_1170 (O_1170,N_48275,N_49667);
or UO_1171 (O_1171,N_48657,N_49560);
xor UO_1172 (O_1172,N_48493,N_48418);
and UO_1173 (O_1173,N_49978,N_49346);
and UO_1174 (O_1174,N_48356,N_48042);
and UO_1175 (O_1175,N_48927,N_48323);
and UO_1176 (O_1176,N_48469,N_48781);
nor UO_1177 (O_1177,N_49173,N_49400);
xnor UO_1178 (O_1178,N_48792,N_49333);
or UO_1179 (O_1179,N_49258,N_49678);
nor UO_1180 (O_1180,N_49279,N_48519);
xor UO_1181 (O_1181,N_48741,N_49102);
and UO_1182 (O_1182,N_48280,N_49810);
and UO_1183 (O_1183,N_49090,N_49988);
or UO_1184 (O_1184,N_49787,N_49767);
or UO_1185 (O_1185,N_49489,N_48469);
or UO_1186 (O_1186,N_49339,N_48897);
or UO_1187 (O_1187,N_49385,N_49640);
and UO_1188 (O_1188,N_48707,N_48465);
nor UO_1189 (O_1189,N_49195,N_49217);
nor UO_1190 (O_1190,N_48568,N_49690);
nor UO_1191 (O_1191,N_48970,N_48798);
and UO_1192 (O_1192,N_49524,N_48430);
nand UO_1193 (O_1193,N_49644,N_49676);
xor UO_1194 (O_1194,N_48525,N_49419);
xor UO_1195 (O_1195,N_49730,N_48636);
nor UO_1196 (O_1196,N_49844,N_48590);
nor UO_1197 (O_1197,N_49821,N_49492);
and UO_1198 (O_1198,N_48054,N_48909);
or UO_1199 (O_1199,N_48059,N_48984);
and UO_1200 (O_1200,N_49564,N_48813);
nor UO_1201 (O_1201,N_48139,N_48147);
or UO_1202 (O_1202,N_48386,N_48382);
xnor UO_1203 (O_1203,N_49645,N_49682);
nand UO_1204 (O_1204,N_48629,N_48719);
nor UO_1205 (O_1205,N_48944,N_49748);
nor UO_1206 (O_1206,N_49774,N_49491);
or UO_1207 (O_1207,N_49729,N_48985);
xor UO_1208 (O_1208,N_48585,N_48673);
or UO_1209 (O_1209,N_49038,N_49345);
or UO_1210 (O_1210,N_48663,N_49366);
or UO_1211 (O_1211,N_49693,N_48409);
nand UO_1212 (O_1212,N_49668,N_49688);
nand UO_1213 (O_1213,N_48416,N_48268);
nand UO_1214 (O_1214,N_48772,N_49171);
xor UO_1215 (O_1215,N_49923,N_48770);
nor UO_1216 (O_1216,N_48042,N_48194);
nor UO_1217 (O_1217,N_49530,N_49296);
and UO_1218 (O_1218,N_48980,N_49379);
or UO_1219 (O_1219,N_48604,N_49634);
or UO_1220 (O_1220,N_48996,N_48688);
and UO_1221 (O_1221,N_49126,N_48463);
nor UO_1222 (O_1222,N_48787,N_48790);
nor UO_1223 (O_1223,N_49508,N_48317);
xor UO_1224 (O_1224,N_49839,N_49266);
nand UO_1225 (O_1225,N_48665,N_48140);
and UO_1226 (O_1226,N_48573,N_49574);
nor UO_1227 (O_1227,N_49473,N_48223);
nor UO_1228 (O_1228,N_48686,N_48709);
nand UO_1229 (O_1229,N_48140,N_49688);
and UO_1230 (O_1230,N_49954,N_49307);
nor UO_1231 (O_1231,N_49170,N_48038);
nand UO_1232 (O_1232,N_49866,N_49307);
nor UO_1233 (O_1233,N_48706,N_49263);
or UO_1234 (O_1234,N_49601,N_49178);
and UO_1235 (O_1235,N_49820,N_49094);
nor UO_1236 (O_1236,N_48771,N_48339);
and UO_1237 (O_1237,N_49627,N_48211);
nor UO_1238 (O_1238,N_49012,N_48116);
xnor UO_1239 (O_1239,N_49802,N_49753);
nor UO_1240 (O_1240,N_48119,N_48620);
nand UO_1241 (O_1241,N_49683,N_49987);
nor UO_1242 (O_1242,N_49037,N_48855);
xnor UO_1243 (O_1243,N_49710,N_49879);
or UO_1244 (O_1244,N_49332,N_49242);
and UO_1245 (O_1245,N_49417,N_49759);
xor UO_1246 (O_1246,N_48284,N_49854);
or UO_1247 (O_1247,N_48461,N_49554);
xnor UO_1248 (O_1248,N_49091,N_48889);
xnor UO_1249 (O_1249,N_48097,N_48221);
and UO_1250 (O_1250,N_48463,N_49859);
xor UO_1251 (O_1251,N_48238,N_48926);
nor UO_1252 (O_1252,N_49388,N_48738);
and UO_1253 (O_1253,N_48262,N_49996);
or UO_1254 (O_1254,N_48455,N_48968);
or UO_1255 (O_1255,N_49967,N_49046);
xnor UO_1256 (O_1256,N_49350,N_49879);
or UO_1257 (O_1257,N_49080,N_48795);
xnor UO_1258 (O_1258,N_48626,N_49471);
or UO_1259 (O_1259,N_49314,N_49940);
xnor UO_1260 (O_1260,N_49255,N_48670);
xnor UO_1261 (O_1261,N_48695,N_49775);
or UO_1262 (O_1262,N_48172,N_49870);
and UO_1263 (O_1263,N_48466,N_48689);
xnor UO_1264 (O_1264,N_48331,N_48531);
and UO_1265 (O_1265,N_49854,N_49221);
nand UO_1266 (O_1266,N_48947,N_48488);
nor UO_1267 (O_1267,N_49074,N_48675);
nand UO_1268 (O_1268,N_48226,N_48536);
nor UO_1269 (O_1269,N_48731,N_49799);
or UO_1270 (O_1270,N_49370,N_49228);
nand UO_1271 (O_1271,N_48226,N_49440);
and UO_1272 (O_1272,N_49536,N_49435);
and UO_1273 (O_1273,N_48754,N_48984);
or UO_1274 (O_1274,N_49672,N_49435);
nand UO_1275 (O_1275,N_49641,N_49503);
or UO_1276 (O_1276,N_49746,N_49290);
or UO_1277 (O_1277,N_49897,N_48781);
and UO_1278 (O_1278,N_48243,N_49027);
nor UO_1279 (O_1279,N_49247,N_48104);
nor UO_1280 (O_1280,N_49770,N_48385);
or UO_1281 (O_1281,N_48975,N_48656);
and UO_1282 (O_1282,N_49657,N_49062);
nor UO_1283 (O_1283,N_48330,N_49630);
and UO_1284 (O_1284,N_49286,N_49022);
and UO_1285 (O_1285,N_48789,N_48000);
nand UO_1286 (O_1286,N_48050,N_49028);
nor UO_1287 (O_1287,N_48442,N_49479);
xnor UO_1288 (O_1288,N_48269,N_48529);
nor UO_1289 (O_1289,N_49401,N_48812);
xor UO_1290 (O_1290,N_48372,N_49064);
xnor UO_1291 (O_1291,N_48003,N_49649);
nor UO_1292 (O_1292,N_48476,N_48357);
nor UO_1293 (O_1293,N_48006,N_48302);
xnor UO_1294 (O_1294,N_48507,N_49993);
xor UO_1295 (O_1295,N_48663,N_48260);
nand UO_1296 (O_1296,N_48099,N_48567);
or UO_1297 (O_1297,N_48310,N_48013);
or UO_1298 (O_1298,N_48184,N_49187);
xnor UO_1299 (O_1299,N_49910,N_48980);
xor UO_1300 (O_1300,N_49257,N_48242);
nor UO_1301 (O_1301,N_49968,N_48686);
and UO_1302 (O_1302,N_48181,N_48318);
and UO_1303 (O_1303,N_49051,N_49909);
xor UO_1304 (O_1304,N_49098,N_49127);
nand UO_1305 (O_1305,N_48955,N_48432);
or UO_1306 (O_1306,N_48429,N_49863);
and UO_1307 (O_1307,N_49240,N_49285);
and UO_1308 (O_1308,N_48185,N_49286);
xnor UO_1309 (O_1309,N_48810,N_48174);
xor UO_1310 (O_1310,N_48370,N_48193);
nand UO_1311 (O_1311,N_48567,N_48354);
nor UO_1312 (O_1312,N_49756,N_48225);
nand UO_1313 (O_1313,N_49426,N_49262);
and UO_1314 (O_1314,N_48006,N_49512);
nor UO_1315 (O_1315,N_48387,N_49160);
nor UO_1316 (O_1316,N_48184,N_48319);
xnor UO_1317 (O_1317,N_48458,N_49634);
and UO_1318 (O_1318,N_49519,N_49621);
or UO_1319 (O_1319,N_49415,N_48699);
nor UO_1320 (O_1320,N_48717,N_48055);
or UO_1321 (O_1321,N_48148,N_49588);
nor UO_1322 (O_1322,N_49295,N_49208);
or UO_1323 (O_1323,N_48624,N_49108);
or UO_1324 (O_1324,N_49199,N_49809);
and UO_1325 (O_1325,N_49295,N_48939);
and UO_1326 (O_1326,N_49186,N_48494);
or UO_1327 (O_1327,N_48578,N_48452);
xor UO_1328 (O_1328,N_48175,N_49354);
and UO_1329 (O_1329,N_48978,N_49694);
and UO_1330 (O_1330,N_48079,N_49296);
nor UO_1331 (O_1331,N_48193,N_49462);
nor UO_1332 (O_1332,N_48550,N_49038);
and UO_1333 (O_1333,N_49190,N_49230);
nor UO_1334 (O_1334,N_49375,N_48982);
xnor UO_1335 (O_1335,N_48917,N_48190);
xnor UO_1336 (O_1336,N_49071,N_49803);
nor UO_1337 (O_1337,N_49343,N_49629);
or UO_1338 (O_1338,N_49902,N_49489);
xnor UO_1339 (O_1339,N_48187,N_49550);
nand UO_1340 (O_1340,N_49236,N_49038);
or UO_1341 (O_1341,N_49757,N_49174);
xor UO_1342 (O_1342,N_48008,N_49411);
and UO_1343 (O_1343,N_48100,N_48119);
nand UO_1344 (O_1344,N_49058,N_48096);
and UO_1345 (O_1345,N_49393,N_48028);
nor UO_1346 (O_1346,N_49696,N_49608);
nand UO_1347 (O_1347,N_49629,N_49442);
nor UO_1348 (O_1348,N_48899,N_48941);
and UO_1349 (O_1349,N_48117,N_49158);
nand UO_1350 (O_1350,N_49763,N_49272);
nand UO_1351 (O_1351,N_48516,N_49398);
nand UO_1352 (O_1352,N_48347,N_49617);
nand UO_1353 (O_1353,N_48026,N_49833);
and UO_1354 (O_1354,N_48388,N_49666);
and UO_1355 (O_1355,N_49703,N_49568);
and UO_1356 (O_1356,N_48785,N_48401);
xnor UO_1357 (O_1357,N_49969,N_49743);
and UO_1358 (O_1358,N_49156,N_49887);
nand UO_1359 (O_1359,N_48176,N_49341);
nor UO_1360 (O_1360,N_49500,N_49172);
or UO_1361 (O_1361,N_49169,N_48016);
xnor UO_1362 (O_1362,N_48227,N_48889);
or UO_1363 (O_1363,N_48220,N_49821);
or UO_1364 (O_1364,N_48266,N_48089);
xor UO_1365 (O_1365,N_48738,N_49123);
nand UO_1366 (O_1366,N_49321,N_48285);
nor UO_1367 (O_1367,N_49049,N_49450);
or UO_1368 (O_1368,N_49198,N_48183);
nand UO_1369 (O_1369,N_49977,N_49984);
and UO_1370 (O_1370,N_48661,N_48376);
nor UO_1371 (O_1371,N_49226,N_48180);
nand UO_1372 (O_1372,N_48643,N_48722);
nor UO_1373 (O_1373,N_49382,N_49238);
and UO_1374 (O_1374,N_49750,N_49502);
nor UO_1375 (O_1375,N_49542,N_49275);
xnor UO_1376 (O_1376,N_48965,N_49887);
and UO_1377 (O_1377,N_48600,N_48306);
nor UO_1378 (O_1378,N_48404,N_48112);
and UO_1379 (O_1379,N_49693,N_49864);
xor UO_1380 (O_1380,N_48936,N_49529);
xnor UO_1381 (O_1381,N_48703,N_49730);
nand UO_1382 (O_1382,N_48407,N_49437);
xor UO_1383 (O_1383,N_49764,N_49357);
nor UO_1384 (O_1384,N_49417,N_48851);
xnor UO_1385 (O_1385,N_48339,N_48604);
nor UO_1386 (O_1386,N_48284,N_49552);
nor UO_1387 (O_1387,N_49802,N_48445);
xnor UO_1388 (O_1388,N_49829,N_49627);
nand UO_1389 (O_1389,N_49363,N_49738);
nor UO_1390 (O_1390,N_49973,N_48039);
xor UO_1391 (O_1391,N_48528,N_48672);
nor UO_1392 (O_1392,N_49037,N_49525);
nand UO_1393 (O_1393,N_48014,N_49058);
or UO_1394 (O_1394,N_48080,N_48140);
nor UO_1395 (O_1395,N_49344,N_49976);
nor UO_1396 (O_1396,N_49724,N_49417);
or UO_1397 (O_1397,N_49305,N_48299);
or UO_1398 (O_1398,N_49451,N_48509);
xnor UO_1399 (O_1399,N_49694,N_48898);
xnor UO_1400 (O_1400,N_49373,N_49254);
xnor UO_1401 (O_1401,N_48865,N_48388);
xor UO_1402 (O_1402,N_48284,N_49691);
nor UO_1403 (O_1403,N_49910,N_48078);
nand UO_1404 (O_1404,N_49710,N_49374);
xor UO_1405 (O_1405,N_49374,N_49016);
or UO_1406 (O_1406,N_49830,N_49679);
nor UO_1407 (O_1407,N_49815,N_49246);
nor UO_1408 (O_1408,N_48842,N_48278);
or UO_1409 (O_1409,N_48203,N_49020);
nor UO_1410 (O_1410,N_48835,N_48497);
or UO_1411 (O_1411,N_48485,N_48630);
xnor UO_1412 (O_1412,N_49374,N_49161);
and UO_1413 (O_1413,N_49575,N_49664);
or UO_1414 (O_1414,N_49378,N_48294);
nand UO_1415 (O_1415,N_48038,N_48402);
nor UO_1416 (O_1416,N_49721,N_49027);
and UO_1417 (O_1417,N_49667,N_49956);
nand UO_1418 (O_1418,N_48389,N_49807);
nor UO_1419 (O_1419,N_48573,N_49595);
and UO_1420 (O_1420,N_49721,N_48471);
xnor UO_1421 (O_1421,N_48701,N_49708);
nor UO_1422 (O_1422,N_49389,N_49027);
or UO_1423 (O_1423,N_48815,N_48322);
nor UO_1424 (O_1424,N_49315,N_48776);
and UO_1425 (O_1425,N_48011,N_48003);
xor UO_1426 (O_1426,N_49698,N_48165);
xnor UO_1427 (O_1427,N_48406,N_48063);
or UO_1428 (O_1428,N_48487,N_49934);
nand UO_1429 (O_1429,N_48142,N_48215);
xnor UO_1430 (O_1430,N_49633,N_48468);
nor UO_1431 (O_1431,N_49887,N_49607);
and UO_1432 (O_1432,N_48409,N_48175);
or UO_1433 (O_1433,N_48980,N_48764);
nor UO_1434 (O_1434,N_49896,N_49971);
and UO_1435 (O_1435,N_48889,N_49734);
or UO_1436 (O_1436,N_49618,N_48824);
xnor UO_1437 (O_1437,N_48837,N_49459);
xor UO_1438 (O_1438,N_49672,N_48610);
nand UO_1439 (O_1439,N_48949,N_49552);
xor UO_1440 (O_1440,N_48722,N_49174);
and UO_1441 (O_1441,N_48026,N_48048);
nor UO_1442 (O_1442,N_48380,N_48552);
nand UO_1443 (O_1443,N_49786,N_48756);
and UO_1444 (O_1444,N_49367,N_48810);
xor UO_1445 (O_1445,N_48698,N_49600);
nor UO_1446 (O_1446,N_49645,N_49179);
nor UO_1447 (O_1447,N_49783,N_48779);
xor UO_1448 (O_1448,N_48964,N_49841);
and UO_1449 (O_1449,N_48805,N_49589);
xor UO_1450 (O_1450,N_48282,N_49195);
xnor UO_1451 (O_1451,N_49494,N_49011);
nand UO_1452 (O_1452,N_49063,N_48037);
xor UO_1453 (O_1453,N_49972,N_48282);
or UO_1454 (O_1454,N_49032,N_48903);
or UO_1455 (O_1455,N_49553,N_48434);
or UO_1456 (O_1456,N_49054,N_49198);
and UO_1457 (O_1457,N_48958,N_48663);
and UO_1458 (O_1458,N_49490,N_49871);
and UO_1459 (O_1459,N_49001,N_48682);
or UO_1460 (O_1460,N_48851,N_49577);
nor UO_1461 (O_1461,N_49572,N_48832);
nand UO_1462 (O_1462,N_48907,N_48126);
and UO_1463 (O_1463,N_48422,N_48328);
or UO_1464 (O_1464,N_48847,N_49017);
or UO_1465 (O_1465,N_48823,N_48643);
and UO_1466 (O_1466,N_48220,N_48007);
or UO_1467 (O_1467,N_49806,N_48281);
xor UO_1468 (O_1468,N_49700,N_49757);
nor UO_1469 (O_1469,N_49318,N_48458);
nor UO_1470 (O_1470,N_48346,N_48591);
and UO_1471 (O_1471,N_49201,N_48814);
or UO_1472 (O_1472,N_48081,N_48860);
xor UO_1473 (O_1473,N_48102,N_49583);
nand UO_1474 (O_1474,N_48211,N_49377);
xor UO_1475 (O_1475,N_48419,N_49350);
nor UO_1476 (O_1476,N_49805,N_48190);
or UO_1477 (O_1477,N_49706,N_48358);
nand UO_1478 (O_1478,N_48889,N_49111);
nor UO_1479 (O_1479,N_48066,N_49669);
and UO_1480 (O_1480,N_49062,N_48385);
and UO_1481 (O_1481,N_48061,N_49132);
nor UO_1482 (O_1482,N_48273,N_49906);
and UO_1483 (O_1483,N_49369,N_48486);
nand UO_1484 (O_1484,N_48251,N_48478);
and UO_1485 (O_1485,N_48047,N_48840);
and UO_1486 (O_1486,N_49582,N_49007);
nand UO_1487 (O_1487,N_49792,N_48646);
and UO_1488 (O_1488,N_48177,N_48668);
nor UO_1489 (O_1489,N_49960,N_48391);
and UO_1490 (O_1490,N_48211,N_48988);
nand UO_1491 (O_1491,N_48193,N_48822);
nand UO_1492 (O_1492,N_49508,N_49357);
or UO_1493 (O_1493,N_49412,N_48714);
xnor UO_1494 (O_1494,N_48920,N_49858);
or UO_1495 (O_1495,N_49087,N_49671);
and UO_1496 (O_1496,N_48897,N_49080);
nor UO_1497 (O_1497,N_48013,N_48214);
or UO_1498 (O_1498,N_49253,N_48145);
and UO_1499 (O_1499,N_48150,N_49331);
nand UO_1500 (O_1500,N_48359,N_49512);
or UO_1501 (O_1501,N_48566,N_48783);
xnor UO_1502 (O_1502,N_49896,N_48566);
and UO_1503 (O_1503,N_48695,N_48039);
xnor UO_1504 (O_1504,N_48598,N_49343);
nand UO_1505 (O_1505,N_48285,N_48278);
xnor UO_1506 (O_1506,N_49180,N_48910);
nor UO_1507 (O_1507,N_48622,N_49127);
nor UO_1508 (O_1508,N_49371,N_48888);
xor UO_1509 (O_1509,N_48843,N_49675);
nand UO_1510 (O_1510,N_49604,N_49224);
nand UO_1511 (O_1511,N_49419,N_48919);
nor UO_1512 (O_1512,N_49595,N_48268);
xnor UO_1513 (O_1513,N_49041,N_48875);
and UO_1514 (O_1514,N_49211,N_49735);
nor UO_1515 (O_1515,N_49165,N_49222);
xnor UO_1516 (O_1516,N_49806,N_48715);
xor UO_1517 (O_1517,N_49078,N_49616);
xnor UO_1518 (O_1518,N_48886,N_48617);
and UO_1519 (O_1519,N_48450,N_49543);
or UO_1520 (O_1520,N_49902,N_48570);
nand UO_1521 (O_1521,N_49544,N_49036);
nand UO_1522 (O_1522,N_48794,N_48253);
xor UO_1523 (O_1523,N_48563,N_49315);
and UO_1524 (O_1524,N_48763,N_48866);
nor UO_1525 (O_1525,N_49591,N_49935);
or UO_1526 (O_1526,N_49571,N_49691);
nand UO_1527 (O_1527,N_49551,N_49359);
and UO_1528 (O_1528,N_49820,N_49413);
and UO_1529 (O_1529,N_48008,N_49741);
nor UO_1530 (O_1530,N_48664,N_49323);
or UO_1531 (O_1531,N_49020,N_48548);
xnor UO_1532 (O_1532,N_49195,N_48399);
or UO_1533 (O_1533,N_48077,N_48546);
nand UO_1534 (O_1534,N_49506,N_48098);
xor UO_1535 (O_1535,N_48971,N_49529);
nor UO_1536 (O_1536,N_49368,N_48212);
or UO_1537 (O_1537,N_49831,N_48561);
nor UO_1538 (O_1538,N_49419,N_48322);
nor UO_1539 (O_1539,N_49787,N_48798);
or UO_1540 (O_1540,N_48925,N_49760);
nor UO_1541 (O_1541,N_48400,N_48718);
nand UO_1542 (O_1542,N_49752,N_48031);
xnor UO_1543 (O_1543,N_49929,N_48267);
xor UO_1544 (O_1544,N_48890,N_48278);
and UO_1545 (O_1545,N_48034,N_48551);
and UO_1546 (O_1546,N_48672,N_49509);
xor UO_1547 (O_1547,N_49960,N_48680);
xor UO_1548 (O_1548,N_48104,N_49035);
and UO_1549 (O_1549,N_48668,N_48101);
nor UO_1550 (O_1550,N_48568,N_48323);
nand UO_1551 (O_1551,N_48773,N_48255);
and UO_1552 (O_1552,N_49212,N_48335);
or UO_1553 (O_1553,N_48975,N_48523);
nor UO_1554 (O_1554,N_48830,N_48321);
xnor UO_1555 (O_1555,N_48006,N_48790);
and UO_1556 (O_1556,N_49548,N_49219);
and UO_1557 (O_1557,N_48337,N_49968);
nor UO_1558 (O_1558,N_49517,N_49998);
or UO_1559 (O_1559,N_49351,N_48147);
and UO_1560 (O_1560,N_48162,N_49383);
or UO_1561 (O_1561,N_49726,N_48413);
nor UO_1562 (O_1562,N_48410,N_48558);
or UO_1563 (O_1563,N_49932,N_49111);
nor UO_1564 (O_1564,N_48663,N_48017);
nand UO_1565 (O_1565,N_48411,N_48002);
and UO_1566 (O_1566,N_48277,N_49401);
or UO_1567 (O_1567,N_49225,N_48567);
nor UO_1568 (O_1568,N_48876,N_48300);
nor UO_1569 (O_1569,N_49017,N_48487);
xnor UO_1570 (O_1570,N_48858,N_49519);
xnor UO_1571 (O_1571,N_48184,N_49613);
nor UO_1572 (O_1572,N_49483,N_48656);
or UO_1573 (O_1573,N_49474,N_49733);
xor UO_1574 (O_1574,N_48443,N_48821);
or UO_1575 (O_1575,N_48786,N_48664);
xnor UO_1576 (O_1576,N_48045,N_48190);
and UO_1577 (O_1577,N_49445,N_49261);
and UO_1578 (O_1578,N_49180,N_49421);
and UO_1579 (O_1579,N_49700,N_49075);
and UO_1580 (O_1580,N_48619,N_48021);
nor UO_1581 (O_1581,N_48723,N_49540);
nor UO_1582 (O_1582,N_48577,N_48239);
and UO_1583 (O_1583,N_49820,N_48237);
and UO_1584 (O_1584,N_48007,N_49681);
nand UO_1585 (O_1585,N_48793,N_48158);
or UO_1586 (O_1586,N_49864,N_49757);
and UO_1587 (O_1587,N_49303,N_49439);
nand UO_1588 (O_1588,N_48733,N_49223);
nor UO_1589 (O_1589,N_49674,N_49291);
nor UO_1590 (O_1590,N_49343,N_49872);
xor UO_1591 (O_1591,N_49904,N_48357);
xor UO_1592 (O_1592,N_48994,N_49630);
nand UO_1593 (O_1593,N_49567,N_48228);
nand UO_1594 (O_1594,N_48281,N_48558);
and UO_1595 (O_1595,N_48832,N_49092);
and UO_1596 (O_1596,N_48725,N_49325);
nand UO_1597 (O_1597,N_49422,N_48780);
xor UO_1598 (O_1598,N_49973,N_49457);
and UO_1599 (O_1599,N_49166,N_49713);
xnor UO_1600 (O_1600,N_48531,N_48702);
xnor UO_1601 (O_1601,N_49514,N_49788);
nand UO_1602 (O_1602,N_48137,N_48606);
nand UO_1603 (O_1603,N_49881,N_48800);
nor UO_1604 (O_1604,N_49458,N_49842);
or UO_1605 (O_1605,N_48506,N_49397);
nor UO_1606 (O_1606,N_48397,N_49121);
nand UO_1607 (O_1607,N_49821,N_49453);
xor UO_1608 (O_1608,N_48155,N_49028);
and UO_1609 (O_1609,N_48910,N_49636);
or UO_1610 (O_1610,N_49146,N_48077);
nor UO_1611 (O_1611,N_49981,N_48827);
nand UO_1612 (O_1612,N_49239,N_48832);
or UO_1613 (O_1613,N_48168,N_49657);
nor UO_1614 (O_1614,N_48210,N_49903);
or UO_1615 (O_1615,N_49978,N_48149);
nor UO_1616 (O_1616,N_49028,N_49612);
nor UO_1617 (O_1617,N_49942,N_49015);
nor UO_1618 (O_1618,N_48406,N_48239);
nand UO_1619 (O_1619,N_49033,N_49631);
nand UO_1620 (O_1620,N_49080,N_48686);
nand UO_1621 (O_1621,N_49905,N_48603);
nor UO_1622 (O_1622,N_49121,N_48463);
xor UO_1623 (O_1623,N_49253,N_48471);
nor UO_1624 (O_1624,N_48992,N_49848);
and UO_1625 (O_1625,N_48455,N_48948);
and UO_1626 (O_1626,N_48071,N_48289);
nor UO_1627 (O_1627,N_49690,N_48742);
nor UO_1628 (O_1628,N_49514,N_49171);
nor UO_1629 (O_1629,N_48566,N_48570);
and UO_1630 (O_1630,N_49149,N_49973);
or UO_1631 (O_1631,N_48480,N_48196);
nand UO_1632 (O_1632,N_49456,N_48532);
and UO_1633 (O_1633,N_48016,N_49085);
or UO_1634 (O_1634,N_49064,N_48101);
or UO_1635 (O_1635,N_48693,N_48330);
nor UO_1636 (O_1636,N_49870,N_48243);
nand UO_1637 (O_1637,N_48156,N_49776);
xor UO_1638 (O_1638,N_49889,N_48910);
and UO_1639 (O_1639,N_48602,N_48958);
xor UO_1640 (O_1640,N_49778,N_49309);
and UO_1641 (O_1641,N_48385,N_49386);
or UO_1642 (O_1642,N_48497,N_49662);
and UO_1643 (O_1643,N_49142,N_49126);
nor UO_1644 (O_1644,N_49488,N_49892);
and UO_1645 (O_1645,N_48065,N_48086);
xor UO_1646 (O_1646,N_49395,N_48566);
xor UO_1647 (O_1647,N_49245,N_49537);
and UO_1648 (O_1648,N_48496,N_48407);
or UO_1649 (O_1649,N_49131,N_48158);
nand UO_1650 (O_1650,N_49355,N_49348);
or UO_1651 (O_1651,N_49842,N_49883);
nor UO_1652 (O_1652,N_48065,N_48968);
or UO_1653 (O_1653,N_49699,N_48454);
xnor UO_1654 (O_1654,N_49800,N_49593);
or UO_1655 (O_1655,N_48924,N_49116);
and UO_1656 (O_1656,N_48398,N_48994);
and UO_1657 (O_1657,N_48804,N_49355);
nand UO_1658 (O_1658,N_49730,N_49506);
or UO_1659 (O_1659,N_49604,N_48000);
and UO_1660 (O_1660,N_49668,N_48971);
xor UO_1661 (O_1661,N_48363,N_49526);
xor UO_1662 (O_1662,N_49924,N_48125);
nand UO_1663 (O_1663,N_49597,N_49434);
xnor UO_1664 (O_1664,N_49050,N_48843);
and UO_1665 (O_1665,N_48270,N_48708);
nand UO_1666 (O_1666,N_49727,N_49242);
and UO_1667 (O_1667,N_49042,N_49381);
or UO_1668 (O_1668,N_48178,N_49877);
and UO_1669 (O_1669,N_49646,N_48235);
nor UO_1670 (O_1670,N_49761,N_48380);
xor UO_1671 (O_1671,N_48706,N_49298);
and UO_1672 (O_1672,N_48566,N_49132);
and UO_1673 (O_1673,N_48888,N_48119);
or UO_1674 (O_1674,N_48114,N_49993);
xnor UO_1675 (O_1675,N_48144,N_48043);
or UO_1676 (O_1676,N_49327,N_49523);
nand UO_1677 (O_1677,N_49032,N_48132);
nor UO_1678 (O_1678,N_49527,N_48790);
nor UO_1679 (O_1679,N_49586,N_49531);
or UO_1680 (O_1680,N_48405,N_48921);
nor UO_1681 (O_1681,N_48232,N_48768);
nand UO_1682 (O_1682,N_48624,N_48463);
and UO_1683 (O_1683,N_49932,N_48115);
nand UO_1684 (O_1684,N_48878,N_48009);
and UO_1685 (O_1685,N_48153,N_49603);
and UO_1686 (O_1686,N_48807,N_48477);
nand UO_1687 (O_1687,N_49699,N_48922);
nor UO_1688 (O_1688,N_48400,N_48656);
nor UO_1689 (O_1689,N_49605,N_48239);
xor UO_1690 (O_1690,N_48817,N_49778);
or UO_1691 (O_1691,N_48620,N_48943);
or UO_1692 (O_1692,N_48852,N_48510);
and UO_1693 (O_1693,N_49302,N_49531);
and UO_1694 (O_1694,N_48736,N_48560);
nor UO_1695 (O_1695,N_48836,N_49876);
and UO_1696 (O_1696,N_49516,N_49786);
and UO_1697 (O_1697,N_49950,N_49415);
nand UO_1698 (O_1698,N_49968,N_48844);
nand UO_1699 (O_1699,N_48645,N_48370);
or UO_1700 (O_1700,N_49125,N_49914);
xor UO_1701 (O_1701,N_48537,N_48666);
xnor UO_1702 (O_1702,N_49131,N_49014);
or UO_1703 (O_1703,N_48975,N_48775);
or UO_1704 (O_1704,N_49849,N_49452);
and UO_1705 (O_1705,N_48308,N_48424);
and UO_1706 (O_1706,N_48223,N_49345);
nand UO_1707 (O_1707,N_49110,N_48544);
nor UO_1708 (O_1708,N_48132,N_49737);
and UO_1709 (O_1709,N_49516,N_49090);
nor UO_1710 (O_1710,N_49901,N_49578);
nor UO_1711 (O_1711,N_49664,N_49548);
and UO_1712 (O_1712,N_49827,N_48072);
nor UO_1713 (O_1713,N_49216,N_48253);
nand UO_1714 (O_1714,N_48331,N_48428);
xor UO_1715 (O_1715,N_49269,N_49498);
xor UO_1716 (O_1716,N_48821,N_48307);
xor UO_1717 (O_1717,N_48154,N_48033);
or UO_1718 (O_1718,N_48036,N_49293);
or UO_1719 (O_1719,N_48635,N_48567);
nor UO_1720 (O_1720,N_48225,N_49031);
nor UO_1721 (O_1721,N_49925,N_49880);
nand UO_1722 (O_1722,N_48341,N_48792);
or UO_1723 (O_1723,N_49917,N_48064);
or UO_1724 (O_1724,N_48309,N_49214);
xor UO_1725 (O_1725,N_48260,N_48011);
nor UO_1726 (O_1726,N_49951,N_49495);
and UO_1727 (O_1727,N_48865,N_48854);
or UO_1728 (O_1728,N_49344,N_49660);
and UO_1729 (O_1729,N_48754,N_49107);
and UO_1730 (O_1730,N_48155,N_48779);
xor UO_1731 (O_1731,N_48471,N_48761);
nand UO_1732 (O_1732,N_49224,N_49087);
and UO_1733 (O_1733,N_49030,N_49738);
nor UO_1734 (O_1734,N_49039,N_49087);
or UO_1735 (O_1735,N_49776,N_49174);
nor UO_1736 (O_1736,N_49245,N_48578);
nor UO_1737 (O_1737,N_49823,N_49085);
and UO_1738 (O_1738,N_48493,N_49134);
and UO_1739 (O_1739,N_48182,N_48099);
and UO_1740 (O_1740,N_48820,N_48182);
nor UO_1741 (O_1741,N_48488,N_48395);
xor UO_1742 (O_1742,N_49542,N_48369);
and UO_1743 (O_1743,N_49955,N_49745);
or UO_1744 (O_1744,N_49509,N_49791);
nand UO_1745 (O_1745,N_48579,N_49352);
nand UO_1746 (O_1746,N_49004,N_48179);
and UO_1747 (O_1747,N_49468,N_49447);
xor UO_1748 (O_1748,N_48144,N_49823);
nor UO_1749 (O_1749,N_49652,N_49596);
or UO_1750 (O_1750,N_49230,N_48731);
nand UO_1751 (O_1751,N_49232,N_49501);
and UO_1752 (O_1752,N_49731,N_49837);
and UO_1753 (O_1753,N_48702,N_48718);
xor UO_1754 (O_1754,N_48221,N_49162);
xnor UO_1755 (O_1755,N_49306,N_48893);
nor UO_1756 (O_1756,N_48082,N_49354);
nor UO_1757 (O_1757,N_48534,N_49025);
or UO_1758 (O_1758,N_49002,N_49819);
nor UO_1759 (O_1759,N_48327,N_49102);
xor UO_1760 (O_1760,N_49413,N_48192);
xnor UO_1761 (O_1761,N_49694,N_48550);
and UO_1762 (O_1762,N_48245,N_49644);
xnor UO_1763 (O_1763,N_49254,N_49506);
and UO_1764 (O_1764,N_48767,N_48384);
and UO_1765 (O_1765,N_49634,N_48193);
xor UO_1766 (O_1766,N_49357,N_48911);
or UO_1767 (O_1767,N_49385,N_48510);
nand UO_1768 (O_1768,N_49306,N_49497);
or UO_1769 (O_1769,N_48959,N_48702);
nand UO_1770 (O_1770,N_48578,N_48522);
nor UO_1771 (O_1771,N_48031,N_48582);
and UO_1772 (O_1772,N_48809,N_49481);
xnor UO_1773 (O_1773,N_49622,N_48050);
nor UO_1774 (O_1774,N_48473,N_49562);
xor UO_1775 (O_1775,N_48834,N_49719);
and UO_1776 (O_1776,N_49242,N_48519);
nand UO_1777 (O_1777,N_48362,N_49277);
or UO_1778 (O_1778,N_49126,N_48915);
nor UO_1779 (O_1779,N_49711,N_49853);
nor UO_1780 (O_1780,N_48951,N_48985);
or UO_1781 (O_1781,N_48819,N_48822);
nor UO_1782 (O_1782,N_49130,N_48567);
and UO_1783 (O_1783,N_48753,N_49449);
xnor UO_1784 (O_1784,N_48736,N_48868);
and UO_1785 (O_1785,N_49271,N_49506);
nand UO_1786 (O_1786,N_48319,N_48662);
and UO_1787 (O_1787,N_48439,N_49449);
xor UO_1788 (O_1788,N_48472,N_48601);
nand UO_1789 (O_1789,N_48084,N_48233);
nor UO_1790 (O_1790,N_49183,N_49574);
or UO_1791 (O_1791,N_48922,N_48264);
or UO_1792 (O_1792,N_48623,N_48190);
nor UO_1793 (O_1793,N_49577,N_49892);
nand UO_1794 (O_1794,N_49071,N_49343);
nor UO_1795 (O_1795,N_49891,N_49740);
and UO_1796 (O_1796,N_48210,N_49839);
nor UO_1797 (O_1797,N_49330,N_48309);
or UO_1798 (O_1798,N_49933,N_49528);
xor UO_1799 (O_1799,N_48933,N_49449);
nor UO_1800 (O_1800,N_49255,N_49137);
nor UO_1801 (O_1801,N_48878,N_49708);
nand UO_1802 (O_1802,N_49690,N_48613);
and UO_1803 (O_1803,N_49707,N_48614);
nor UO_1804 (O_1804,N_48208,N_48297);
nor UO_1805 (O_1805,N_49592,N_49002);
nor UO_1806 (O_1806,N_49160,N_49667);
or UO_1807 (O_1807,N_48015,N_49070);
or UO_1808 (O_1808,N_49853,N_49394);
nor UO_1809 (O_1809,N_49326,N_49448);
and UO_1810 (O_1810,N_49908,N_49553);
nor UO_1811 (O_1811,N_48183,N_49528);
xor UO_1812 (O_1812,N_49878,N_48728);
or UO_1813 (O_1813,N_49788,N_49376);
and UO_1814 (O_1814,N_49760,N_48388);
and UO_1815 (O_1815,N_48036,N_49040);
nand UO_1816 (O_1816,N_49595,N_48821);
and UO_1817 (O_1817,N_48299,N_48425);
and UO_1818 (O_1818,N_48753,N_48155);
nand UO_1819 (O_1819,N_48989,N_49450);
nor UO_1820 (O_1820,N_49974,N_49618);
nor UO_1821 (O_1821,N_48913,N_48917);
or UO_1822 (O_1822,N_49864,N_48020);
xor UO_1823 (O_1823,N_48107,N_48069);
xnor UO_1824 (O_1824,N_48606,N_48098);
xor UO_1825 (O_1825,N_48609,N_48202);
nor UO_1826 (O_1826,N_48425,N_48470);
xor UO_1827 (O_1827,N_49708,N_48824);
nand UO_1828 (O_1828,N_49734,N_49372);
and UO_1829 (O_1829,N_48755,N_48237);
or UO_1830 (O_1830,N_48674,N_48357);
or UO_1831 (O_1831,N_48107,N_49076);
or UO_1832 (O_1832,N_49497,N_49002);
or UO_1833 (O_1833,N_49773,N_48742);
nor UO_1834 (O_1834,N_48821,N_49423);
and UO_1835 (O_1835,N_48261,N_49292);
nand UO_1836 (O_1836,N_49155,N_49237);
nor UO_1837 (O_1837,N_49406,N_48000);
nor UO_1838 (O_1838,N_49012,N_49939);
or UO_1839 (O_1839,N_49182,N_48092);
and UO_1840 (O_1840,N_49723,N_49064);
nand UO_1841 (O_1841,N_49490,N_48123);
nand UO_1842 (O_1842,N_48015,N_48105);
nor UO_1843 (O_1843,N_48506,N_49187);
nand UO_1844 (O_1844,N_48040,N_48503);
nand UO_1845 (O_1845,N_48372,N_49754);
or UO_1846 (O_1846,N_48296,N_49055);
nor UO_1847 (O_1847,N_49662,N_48252);
or UO_1848 (O_1848,N_49246,N_49547);
nand UO_1849 (O_1849,N_48357,N_49575);
nor UO_1850 (O_1850,N_49664,N_49313);
or UO_1851 (O_1851,N_48076,N_48474);
nand UO_1852 (O_1852,N_49658,N_48095);
xor UO_1853 (O_1853,N_48105,N_49021);
nor UO_1854 (O_1854,N_48386,N_48133);
or UO_1855 (O_1855,N_49120,N_48848);
xor UO_1856 (O_1856,N_49394,N_49520);
xor UO_1857 (O_1857,N_48513,N_48866);
nand UO_1858 (O_1858,N_49536,N_49503);
nand UO_1859 (O_1859,N_48038,N_49049);
nand UO_1860 (O_1860,N_49350,N_48094);
nor UO_1861 (O_1861,N_48656,N_49444);
xor UO_1862 (O_1862,N_48968,N_49168);
and UO_1863 (O_1863,N_48319,N_49730);
nor UO_1864 (O_1864,N_48048,N_49701);
and UO_1865 (O_1865,N_48103,N_49063);
nand UO_1866 (O_1866,N_49434,N_49116);
or UO_1867 (O_1867,N_48431,N_48083);
nand UO_1868 (O_1868,N_48845,N_48644);
and UO_1869 (O_1869,N_49717,N_49169);
and UO_1870 (O_1870,N_48244,N_48916);
nand UO_1871 (O_1871,N_49250,N_49709);
xnor UO_1872 (O_1872,N_48508,N_49833);
or UO_1873 (O_1873,N_49922,N_48568);
and UO_1874 (O_1874,N_49987,N_48365);
nor UO_1875 (O_1875,N_49856,N_49851);
or UO_1876 (O_1876,N_48791,N_49658);
nand UO_1877 (O_1877,N_49477,N_49097);
or UO_1878 (O_1878,N_48645,N_48386);
nor UO_1879 (O_1879,N_49219,N_49947);
nand UO_1880 (O_1880,N_49486,N_48466);
or UO_1881 (O_1881,N_49944,N_49064);
nand UO_1882 (O_1882,N_48334,N_49377);
nor UO_1883 (O_1883,N_49673,N_49631);
nand UO_1884 (O_1884,N_48750,N_49593);
or UO_1885 (O_1885,N_49077,N_48711);
and UO_1886 (O_1886,N_49616,N_48990);
and UO_1887 (O_1887,N_48939,N_49269);
nand UO_1888 (O_1888,N_49644,N_48280);
and UO_1889 (O_1889,N_49371,N_48964);
xor UO_1890 (O_1890,N_49885,N_49807);
or UO_1891 (O_1891,N_49036,N_48102);
or UO_1892 (O_1892,N_48111,N_48562);
xor UO_1893 (O_1893,N_48979,N_48010);
nor UO_1894 (O_1894,N_49313,N_49028);
nand UO_1895 (O_1895,N_48509,N_49996);
nor UO_1896 (O_1896,N_49988,N_49921);
nand UO_1897 (O_1897,N_49952,N_48031);
xor UO_1898 (O_1898,N_49024,N_48154);
nand UO_1899 (O_1899,N_49197,N_49069);
or UO_1900 (O_1900,N_48091,N_49600);
or UO_1901 (O_1901,N_48692,N_48650);
nand UO_1902 (O_1902,N_48895,N_49264);
nor UO_1903 (O_1903,N_48658,N_48754);
nor UO_1904 (O_1904,N_48653,N_49923);
nand UO_1905 (O_1905,N_49969,N_49482);
and UO_1906 (O_1906,N_48510,N_49947);
nor UO_1907 (O_1907,N_49461,N_48797);
or UO_1908 (O_1908,N_49765,N_48191);
or UO_1909 (O_1909,N_48360,N_48844);
nand UO_1910 (O_1910,N_49095,N_48708);
nor UO_1911 (O_1911,N_48886,N_48786);
xnor UO_1912 (O_1912,N_48475,N_49771);
or UO_1913 (O_1913,N_48047,N_48577);
nor UO_1914 (O_1914,N_48575,N_49496);
xor UO_1915 (O_1915,N_48816,N_48244);
nand UO_1916 (O_1916,N_48019,N_49420);
nor UO_1917 (O_1917,N_49866,N_48160);
or UO_1918 (O_1918,N_48369,N_49792);
and UO_1919 (O_1919,N_49833,N_48487);
nor UO_1920 (O_1920,N_48437,N_49972);
and UO_1921 (O_1921,N_49099,N_48540);
or UO_1922 (O_1922,N_49624,N_48587);
nand UO_1923 (O_1923,N_49095,N_49421);
or UO_1924 (O_1924,N_48573,N_48457);
and UO_1925 (O_1925,N_49821,N_48205);
and UO_1926 (O_1926,N_49458,N_48258);
xor UO_1927 (O_1927,N_48471,N_49619);
and UO_1928 (O_1928,N_49421,N_49428);
and UO_1929 (O_1929,N_48077,N_48247);
or UO_1930 (O_1930,N_48108,N_48129);
xor UO_1931 (O_1931,N_48906,N_48915);
or UO_1932 (O_1932,N_48303,N_48168);
or UO_1933 (O_1933,N_49036,N_48488);
nor UO_1934 (O_1934,N_49829,N_49445);
nand UO_1935 (O_1935,N_49654,N_49853);
and UO_1936 (O_1936,N_49239,N_49492);
nor UO_1937 (O_1937,N_49051,N_48480);
nor UO_1938 (O_1938,N_48321,N_49146);
nand UO_1939 (O_1939,N_48380,N_49916);
or UO_1940 (O_1940,N_49216,N_48516);
and UO_1941 (O_1941,N_48793,N_49620);
nor UO_1942 (O_1942,N_48500,N_48591);
or UO_1943 (O_1943,N_49369,N_49979);
and UO_1944 (O_1944,N_48831,N_49595);
xor UO_1945 (O_1945,N_49702,N_49455);
xor UO_1946 (O_1946,N_48777,N_48258);
nor UO_1947 (O_1947,N_49137,N_49918);
nor UO_1948 (O_1948,N_48349,N_49143);
and UO_1949 (O_1949,N_48908,N_48499);
nor UO_1950 (O_1950,N_48508,N_49000);
nand UO_1951 (O_1951,N_49743,N_48825);
xor UO_1952 (O_1952,N_49999,N_48246);
and UO_1953 (O_1953,N_49685,N_49222);
nor UO_1954 (O_1954,N_49483,N_49634);
and UO_1955 (O_1955,N_49024,N_48235);
nor UO_1956 (O_1956,N_49345,N_48141);
nand UO_1957 (O_1957,N_49133,N_49499);
and UO_1958 (O_1958,N_49960,N_48453);
or UO_1959 (O_1959,N_48802,N_48126);
and UO_1960 (O_1960,N_49201,N_48410);
or UO_1961 (O_1961,N_48883,N_49903);
nor UO_1962 (O_1962,N_49504,N_49948);
or UO_1963 (O_1963,N_49681,N_48961);
or UO_1964 (O_1964,N_48164,N_48891);
nand UO_1965 (O_1965,N_48646,N_48367);
xnor UO_1966 (O_1966,N_49027,N_49962);
nand UO_1967 (O_1967,N_49158,N_48177);
or UO_1968 (O_1968,N_49227,N_48114);
and UO_1969 (O_1969,N_48260,N_48079);
nor UO_1970 (O_1970,N_49664,N_49031);
or UO_1971 (O_1971,N_49775,N_49505);
xor UO_1972 (O_1972,N_48653,N_49511);
nand UO_1973 (O_1973,N_48238,N_48934);
nand UO_1974 (O_1974,N_48303,N_49524);
nor UO_1975 (O_1975,N_49670,N_49896);
xnor UO_1976 (O_1976,N_48099,N_49149);
nor UO_1977 (O_1977,N_48445,N_48293);
nand UO_1978 (O_1978,N_49108,N_48915);
or UO_1979 (O_1979,N_49571,N_48710);
nor UO_1980 (O_1980,N_48514,N_48790);
and UO_1981 (O_1981,N_49100,N_48228);
or UO_1982 (O_1982,N_49832,N_48509);
nor UO_1983 (O_1983,N_49015,N_49722);
and UO_1984 (O_1984,N_49598,N_48353);
or UO_1985 (O_1985,N_49701,N_49742);
nor UO_1986 (O_1986,N_49938,N_49396);
xnor UO_1987 (O_1987,N_48068,N_49422);
or UO_1988 (O_1988,N_49304,N_48022);
xnor UO_1989 (O_1989,N_49255,N_49478);
and UO_1990 (O_1990,N_49170,N_49709);
xor UO_1991 (O_1991,N_48771,N_48184);
and UO_1992 (O_1992,N_48098,N_48569);
or UO_1993 (O_1993,N_49842,N_48123);
nand UO_1994 (O_1994,N_48890,N_48817);
or UO_1995 (O_1995,N_49777,N_49470);
nor UO_1996 (O_1996,N_48014,N_49165);
xnor UO_1997 (O_1997,N_48261,N_49646);
xor UO_1998 (O_1998,N_48594,N_49704);
nor UO_1999 (O_1999,N_48921,N_48212);
nor UO_2000 (O_2000,N_48481,N_49771);
nor UO_2001 (O_2001,N_49299,N_49084);
xnor UO_2002 (O_2002,N_48022,N_49564);
nand UO_2003 (O_2003,N_49229,N_48288);
and UO_2004 (O_2004,N_49062,N_48664);
xnor UO_2005 (O_2005,N_48766,N_49280);
or UO_2006 (O_2006,N_48023,N_48820);
nand UO_2007 (O_2007,N_49411,N_48063);
or UO_2008 (O_2008,N_48563,N_48055);
and UO_2009 (O_2009,N_48521,N_48621);
and UO_2010 (O_2010,N_49954,N_49369);
nand UO_2011 (O_2011,N_49074,N_48768);
nor UO_2012 (O_2012,N_49096,N_49660);
nand UO_2013 (O_2013,N_48635,N_48184);
or UO_2014 (O_2014,N_49207,N_49404);
and UO_2015 (O_2015,N_49083,N_49772);
or UO_2016 (O_2016,N_49597,N_48376);
and UO_2017 (O_2017,N_49466,N_48355);
or UO_2018 (O_2018,N_48663,N_49107);
nor UO_2019 (O_2019,N_49470,N_49875);
nor UO_2020 (O_2020,N_49383,N_49114);
and UO_2021 (O_2021,N_48171,N_48734);
nand UO_2022 (O_2022,N_49650,N_49767);
nand UO_2023 (O_2023,N_48842,N_49894);
nand UO_2024 (O_2024,N_48365,N_49957);
xnor UO_2025 (O_2025,N_48309,N_48260);
xor UO_2026 (O_2026,N_49104,N_48745);
xnor UO_2027 (O_2027,N_49863,N_48608);
and UO_2028 (O_2028,N_49602,N_48189);
nand UO_2029 (O_2029,N_49847,N_48447);
and UO_2030 (O_2030,N_48799,N_49604);
and UO_2031 (O_2031,N_48364,N_48587);
and UO_2032 (O_2032,N_48203,N_49224);
nor UO_2033 (O_2033,N_49542,N_48257);
xor UO_2034 (O_2034,N_49579,N_49367);
and UO_2035 (O_2035,N_48217,N_49386);
xnor UO_2036 (O_2036,N_48140,N_48022);
or UO_2037 (O_2037,N_48357,N_48083);
nor UO_2038 (O_2038,N_49879,N_49492);
xor UO_2039 (O_2039,N_49652,N_48144);
or UO_2040 (O_2040,N_48935,N_48267);
xnor UO_2041 (O_2041,N_49779,N_49370);
xor UO_2042 (O_2042,N_48613,N_48866);
and UO_2043 (O_2043,N_49715,N_48192);
nand UO_2044 (O_2044,N_49987,N_48172);
and UO_2045 (O_2045,N_49451,N_49930);
xor UO_2046 (O_2046,N_49306,N_48044);
nand UO_2047 (O_2047,N_49987,N_49734);
nand UO_2048 (O_2048,N_48256,N_48517);
nor UO_2049 (O_2049,N_49577,N_49022);
nor UO_2050 (O_2050,N_49230,N_49539);
nand UO_2051 (O_2051,N_49078,N_48324);
and UO_2052 (O_2052,N_49685,N_48666);
nor UO_2053 (O_2053,N_48496,N_48059);
or UO_2054 (O_2054,N_48968,N_49912);
or UO_2055 (O_2055,N_49528,N_48540);
nand UO_2056 (O_2056,N_48561,N_48165);
and UO_2057 (O_2057,N_48412,N_48034);
nor UO_2058 (O_2058,N_48957,N_48010);
nand UO_2059 (O_2059,N_49812,N_49113);
nor UO_2060 (O_2060,N_49410,N_48196);
nor UO_2061 (O_2061,N_48418,N_49064);
xnor UO_2062 (O_2062,N_48446,N_48919);
or UO_2063 (O_2063,N_49939,N_48833);
xor UO_2064 (O_2064,N_49305,N_48657);
or UO_2065 (O_2065,N_49926,N_48686);
and UO_2066 (O_2066,N_49786,N_48719);
nand UO_2067 (O_2067,N_49882,N_49640);
xor UO_2068 (O_2068,N_48778,N_48442);
nor UO_2069 (O_2069,N_49197,N_48406);
or UO_2070 (O_2070,N_48143,N_48287);
nor UO_2071 (O_2071,N_48314,N_48195);
nor UO_2072 (O_2072,N_49706,N_48437);
xnor UO_2073 (O_2073,N_49419,N_49879);
nand UO_2074 (O_2074,N_48028,N_49043);
or UO_2075 (O_2075,N_49016,N_49199);
or UO_2076 (O_2076,N_48523,N_49908);
nor UO_2077 (O_2077,N_49603,N_49886);
nand UO_2078 (O_2078,N_49780,N_48284);
or UO_2079 (O_2079,N_48708,N_48595);
xnor UO_2080 (O_2080,N_48466,N_48878);
or UO_2081 (O_2081,N_49025,N_48987);
nand UO_2082 (O_2082,N_49251,N_49990);
and UO_2083 (O_2083,N_49808,N_48263);
xor UO_2084 (O_2084,N_48163,N_49784);
nor UO_2085 (O_2085,N_48055,N_48405);
xor UO_2086 (O_2086,N_49138,N_48481);
xor UO_2087 (O_2087,N_48441,N_48968);
nor UO_2088 (O_2088,N_48256,N_48074);
nand UO_2089 (O_2089,N_48883,N_48906);
or UO_2090 (O_2090,N_48107,N_49824);
xnor UO_2091 (O_2091,N_49076,N_49463);
nand UO_2092 (O_2092,N_48071,N_49125);
nand UO_2093 (O_2093,N_48307,N_49310);
nand UO_2094 (O_2094,N_48111,N_48344);
xnor UO_2095 (O_2095,N_49648,N_49904);
or UO_2096 (O_2096,N_48232,N_48774);
xor UO_2097 (O_2097,N_49657,N_48100);
or UO_2098 (O_2098,N_49311,N_49662);
xnor UO_2099 (O_2099,N_48792,N_48359);
nand UO_2100 (O_2100,N_48050,N_49922);
nor UO_2101 (O_2101,N_48324,N_49348);
nor UO_2102 (O_2102,N_49711,N_48937);
nand UO_2103 (O_2103,N_49917,N_49570);
xor UO_2104 (O_2104,N_48607,N_49552);
xnor UO_2105 (O_2105,N_48903,N_49225);
or UO_2106 (O_2106,N_49022,N_49980);
and UO_2107 (O_2107,N_48624,N_49116);
and UO_2108 (O_2108,N_48347,N_48943);
and UO_2109 (O_2109,N_48717,N_49685);
nand UO_2110 (O_2110,N_48269,N_48178);
nand UO_2111 (O_2111,N_48608,N_48101);
and UO_2112 (O_2112,N_49043,N_49319);
xnor UO_2113 (O_2113,N_48891,N_48076);
or UO_2114 (O_2114,N_48159,N_48010);
nand UO_2115 (O_2115,N_48051,N_48325);
xnor UO_2116 (O_2116,N_48704,N_49481);
and UO_2117 (O_2117,N_49167,N_49176);
and UO_2118 (O_2118,N_48737,N_48310);
and UO_2119 (O_2119,N_49193,N_48224);
nor UO_2120 (O_2120,N_49062,N_49612);
nor UO_2121 (O_2121,N_49118,N_48429);
nor UO_2122 (O_2122,N_49430,N_48705);
xor UO_2123 (O_2123,N_48671,N_49203);
and UO_2124 (O_2124,N_48165,N_49458);
nor UO_2125 (O_2125,N_48675,N_49212);
or UO_2126 (O_2126,N_49682,N_48652);
xnor UO_2127 (O_2127,N_48086,N_48803);
xnor UO_2128 (O_2128,N_48873,N_49563);
xnor UO_2129 (O_2129,N_49547,N_48175);
or UO_2130 (O_2130,N_48383,N_48920);
xnor UO_2131 (O_2131,N_49773,N_48662);
and UO_2132 (O_2132,N_49392,N_48895);
nand UO_2133 (O_2133,N_49663,N_48160);
nand UO_2134 (O_2134,N_48935,N_48126);
nor UO_2135 (O_2135,N_49554,N_49364);
nand UO_2136 (O_2136,N_49009,N_49593);
nor UO_2137 (O_2137,N_49639,N_48121);
or UO_2138 (O_2138,N_48824,N_48243);
nor UO_2139 (O_2139,N_48102,N_49049);
nor UO_2140 (O_2140,N_49856,N_49296);
nand UO_2141 (O_2141,N_48548,N_48182);
nand UO_2142 (O_2142,N_48241,N_49866);
or UO_2143 (O_2143,N_49145,N_49595);
nor UO_2144 (O_2144,N_49556,N_49244);
nand UO_2145 (O_2145,N_48260,N_48406);
xnor UO_2146 (O_2146,N_49937,N_49294);
nor UO_2147 (O_2147,N_49174,N_49126);
nand UO_2148 (O_2148,N_49554,N_48983);
nand UO_2149 (O_2149,N_48968,N_48063);
and UO_2150 (O_2150,N_48628,N_48179);
and UO_2151 (O_2151,N_48111,N_49106);
nand UO_2152 (O_2152,N_48928,N_49152);
nor UO_2153 (O_2153,N_49555,N_49620);
and UO_2154 (O_2154,N_48208,N_49000);
or UO_2155 (O_2155,N_48768,N_49335);
nand UO_2156 (O_2156,N_48878,N_49206);
or UO_2157 (O_2157,N_48425,N_49689);
and UO_2158 (O_2158,N_49578,N_49265);
or UO_2159 (O_2159,N_49460,N_49219);
and UO_2160 (O_2160,N_49279,N_49303);
and UO_2161 (O_2161,N_48044,N_49729);
xor UO_2162 (O_2162,N_48690,N_48716);
and UO_2163 (O_2163,N_49875,N_49651);
or UO_2164 (O_2164,N_48645,N_48604);
nor UO_2165 (O_2165,N_49834,N_49946);
or UO_2166 (O_2166,N_48727,N_48394);
and UO_2167 (O_2167,N_48272,N_49279);
nand UO_2168 (O_2168,N_48411,N_49876);
xnor UO_2169 (O_2169,N_49914,N_48281);
or UO_2170 (O_2170,N_48968,N_48792);
and UO_2171 (O_2171,N_49166,N_48603);
or UO_2172 (O_2172,N_49310,N_49839);
xnor UO_2173 (O_2173,N_48304,N_49825);
or UO_2174 (O_2174,N_49156,N_49229);
and UO_2175 (O_2175,N_49696,N_48552);
or UO_2176 (O_2176,N_49929,N_49836);
nand UO_2177 (O_2177,N_49789,N_49709);
xnor UO_2178 (O_2178,N_49849,N_49650);
or UO_2179 (O_2179,N_48247,N_48280);
xnor UO_2180 (O_2180,N_48691,N_48320);
xor UO_2181 (O_2181,N_48438,N_49108);
nor UO_2182 (O_2182,N_48227,N_49868);
and UO_2183 (O_2183,N_49135,N_48355);
nor UO_2184 (O_2184,N_49723,N_48941);
xor UO_2185 (O_2185,N_48233,N_48311);
xnor UO_2186 (O_2186,N_49385,N_49568);
nand UO_2187 (O_2187,N_48291,N_48571);
and UO_2188 (O_2188,N_49865,N_49321);
xnor UO_2189 (O_2189,N_48590,N_49900);
and UO_2190 (O_2190,N_48044,N_49399);
xnor UO_2191 (O_2191,N_49374,N_49666);
nor UO_2192 (O_2192,N_48797,N_48643);
or UO_2193 (O_2193,N_49272,N_48662);
nor UO_2194 (O_2194,N_48013,N_49670);
nand UO_2195 (O_2195,N_48987,N_48210);
nor UO_2196 (O_2196,N_49970,N_48419);
and UO_2197 (O_2197,N_49945,N_49854);
nor UO_2198 (O_2198,N_48605,N_48957);
and UO_2199 (O_2199,N_49158,N_49563);
nor UO_2200 (O_2200,N_49091,N_49033);
or UO_2201 (O_2201,N_49698,N_49564);
and UO_2202 (O_2202,N_49545,N_49718);
nor UO_2203 (O_2203,N_49770,N_49421);
nor UO_2204 (O_2204,N_48818,N_49473);
or UO_2205 (O_2205,N_49018,N_48667);
xnor UO_2206 (O_2206,N_49933,N_48564);
nor UO_2207 (O_2207,N_49829,N_49088);
xor UO_2208 (O_2208,N_49548,N_48087);
nor UO_2209 (O_2209,N_48082,N_48003);
and UO_2210 (O_2210,N_49309,N_48582);
and UO_2211 (O_2211,N_49092,N_48026);
and UO_2212 (O_2212,N_48656,N_49290);
or UO_2213 (O_2213,N_48927,N_49132);
and UO_2214 (O_2214,N_49035,N_48618);
and UO_2215 (O_2215,N_49590,N_49781);
nand UO_2216 (O_2216,N_49158,N_49329);
xor UO_2217 (O_2217,N_48186,N_48038);
nand UO_2218 (O_2218,N_49554,N_49559);
xor UO_2219 (O_2219,N_48343,N_49363);
nand UO_2220 (O_2220,N_48413,N_48434);
nor UO_2221 (O_2221,N_48800,N_49121);
xor UO_2222 (O_2222,N_49304,N_49643);
nor UO_2223 (O_2223,N_48427,N_48576);
xnor UO_2224 (O_2224,N_48113,N_48997);
and UO_2225 (O_2225,N_48641,N_49194);
nand UO_2226 (O_2226,N_48155,N_48295);
nor UO_2227 (O_2227,N_48491,N_49709);
nand UO_2228 (O_2228,N_48071,N_49867);
nand UO_2229 (O_2229,N_49872,N_48890);
nand UO_2230 (O_2230,N_49326,N_49623);
nand UO_2231 (O_2231,N_49659,N_48004);
nand UO_2232 (O_2232,N_49005,N_48386);
xor UO_2233 (O_2233,N_48853,N_49203);
or UO_2234 (O_2234,N_49710,N_49820);
or UO_2235 (O_2235,N_49951,N_49593);
nor UO_2236 (O_2236,N_49507,N_48877);
nand UO_2237 (O_2237,N_49924,N_48339);
nor UO_2238 (O_2238,N_49361,N_48734);
xor UO_2239 (O_2239,N_48153,N_48131);
nand UO_2240 (O_2240,N_49916,N_49510);
and UO_2241 (O_2241,N_48505,N_48408);
and UO_2242 (O_2242,N_48337,N_48215);
nor UO_2243 (O_2243,N_48131,N_48175);
xnor UO_2244 (O_2244,N_48055,N_48892);
nand UO_2245 (O_2245,N_48355,N_48472);
and UO_2246 (O_2246,N_48713,N_48735);
or UO_2247 (O_2247,N_48327,N_49868);
nand UO_2248 (O_2248,N_49979,N_49863);
nor UO_2249 (O_2249,N_48760,N_48560);
and UO_2250 (O_2250,N_48247,N_48576);
xor UO_2251 (O_2251,N_49050,N_48802);
nor UO_2252 (O_2252,N_49938,N_49696);
nand UO_2253 (O_2253,N_49859,N_48080);
xor UO_2254 (O_2254,N_48776,N_48706);
nor UO_2255 (O_2255,N_48310,N_49933);
and UO_2256 (O_2256,N_49039,N_49120);
and UO_2257 (O_2257,N_49964,N_48008);
nand UO_2258 (O_2258,N_49042,N_49403);
nor UO_2259 (O_2259,N_49753,N_48385);
nor UO_2260 (O_2260,N_48164,N_48163);
nor UO_2261 (O_2261,N_48230,N_48808);
and UO_2262 (O_2262,N_48196,N_48358);
nor UO_2263 (O_2263,N_48479,N_48348);
or UO_2264 (O_2264,N_48792,N_48394);
xnor UO_2265 (O_2265,N_48387,N_49888);
xnor UO_2266 (O_2266,N_48968,N_48867);
xnor UO_2267 (O_2267,N_49901,N_49317);
or UO_2268 (O_2268,N_48013,N_49813);
or UO_2269 (O_2269,N_48106,N_49216);
or UO_2270 (O_2270,N_48099,N_48502);
or UO_2271 (O_2271,N_49226,N_49352);
xnor UO_2272 (O_2272,N_49834,N_48792);
nand UO_2273 (O_2273,N_48165,N_49816);
nand UO_2274 (O_2274,N_49889,N_49462);
nor UO_2275 (O_2275,N_49789,N_48843);
or UO_2276 (O_2276,N_48697,N_48526);
or UO_2277 (O_2277,N_49224,N_49818);
xor UO_2278 (O_2278,N_48686,N_48638);
nor UO_2279 (O_2279,N_48245,N_48412);
or UO_2280 (O_2280,N_49196,N_49222);
and UO_2281 (O_2281,N_49666,N_49982);
and UO_2282 (O_2282,N_48650,N_49748);
and UO_2283 (O_2283,N_48354,N_49868);
nand UO_2284 (O_2284,N_48035,N_49505);
and UO_2285 (O_2285,N_49767,N_49264);
or UO_2286 (O_2286,N_49584,N_48531);
and UO_2287 (O_2287,N_49652,N_48027);
nor UO_2288 (O_2288,N_48880,N_49990);
and UO_2289 (O_2289,N_49798,N_49660);
and UO_2290 (O_2290,N_49392,N_48564);
or UO_2291 (O_2291,N_49719,N_48913);
nand UO_2292 (O_2292,N_49397,N_48173);
and UO_2293 (O_2293,N_49571,N_48767);
nand UO_2294 (O_2294,N_48486,N_49861);
or UO_2295 (O_2295,N_48730,N_48477);
nand UO_2296 (O_2296,N_49397,N_49299);
xor UO_2297 (O_2297,N_48305,N_48487);
nor UO_2298 (O_2298,N_49325,N_48746);
and UO_2299 (O_2299,N_49354,N_48999);
nand UO_2300 (O_2300,N_49792,N_48714);
xnor UO_2301 (O_2301,N_49458,N_48306);
xor UO_2302 (O_2302,N_49647,N_48340);
nand UO_2303 (O_2303,N_48474,N_48327);
or UO_2304 (O_2304,N_49731,N_49730);
xnor UO_2305 (O_2305,N_48236,N_49731);
or UO_2306 (O_2306,N_48147,N_49970);
xor UO_2307 (O_2307,N_49813,N_48618);
or UO_2308 (O_2308,N_49545,N_48918);
nor UO_2309 (O_2309,N_48201,N_48786);
xnor UO_2310 (O_2310,N_49177,N_49711);
nand UO_2311 (O_2311,N_49369,N_48953);
or UO_2312 (O_2312,N_48460,N_48518);
or UO_2313 (O_2313,N_48405,N_49718);
nor UO_2314 (O_2314,N_48562,N_49905);
nor UO_2315 (O_2315,N_48723,N_49215);
nor UO_2316 (O_2316,N_49563,N_48719);
or UO_2317 (O_2317,N_49222,N_49400);
xor UO_2318 (O_2318,N_48161,N_49506);
or UO_2319 (O_2319,N_48429,N_48523);
xnor UO_2320 (O_2320,N_49013,N_48793);
and UO_2321 (O_2321,N_48647,N_49272);
nor UO_2322 (O_2322,N_49743,N_48629);
and UO_2323 (O_2323,N_48386,N_49732);
and UO_2324 (O_2324,N_48066,N_49307);
and UO_2325 (O_2325,N_49599,N_48522);
xnor UO_2326 (O_2326,N_49022,N_49065);
nor UO_2327 (O_2327,N_49809,N_48026);
nand UO_2328 (O_2328,N_49062,N_48940);
nor UO_2329 (O_2329,N_49087,N_49150);
xnor UO_2330 (O_2330,N_49013,N_48226);
nand UO_2331 (O_2331,N_48014,N_49972);
nor UO_2332 (O_2332,N_49931,N_49718);
and UO_2333 (O_2333,N_49125,N_49337);
or UO_2334 (O_2334,N_48756,N_49020);
nand UO_2335 (O_2335,N_49618,N_48593);
and UO_2336 (O_2336,N_48758,N_48847);
nor UO_2337 (O_2337,N_49654,N_48182);
xor UO_2338 (O_2338,N_49908,N_48414);
nand UO_2339 (O_2339,N_48961,N_49631);
nor UO_2340 (O_2340,N_48078,N_49397);
xor UO_2341 (O_2341,N_48981,N_49983);
and UO_2342 (O_2342,N_48532,N_48531);
nor UO_2343 (O_2343,N_48223,N_48819);
and UO_2344 (O_2344,N_48100,N_48751);
nor UO_2345 (O_2345,N_48760,N_49090);
xor UO_2346 (O_2346,N_49212,N_48952);
xnor UO_2347 (O_2347,N_49176,N_49199);
nand UO_2348 (O_2348,N_49563,N_48026);
or UO_2349 (O_2349,N_48090,N_48955);
and UO_2350 (O_2350,N_49117,N_48618);
xnor UO_2351 (O_2351,N_48576,N_48993);
and UO_2352 (O_2352,N_48942,N_49148);
or UO_2353 (O_2353,N_48591,N_49692);
or UO_2354 (O_2354,N_49728,N_49986);
or UO_2355 (O_2355,N_48744,N_49104);
xnor UO_2356 (O_2356,N_49511,N_48547);
or UO_2357 (O_2357,N_48189,N_48493);
nor UO_2358 (O_2358,N_49442,N_48430);
xor UO_2359 (O_2359,N_48110,N_48964);
or UO_2360 (O_2360,N_49670,N_49594);
or UO_2361 (O_2361,N_48921,N_48639);
and UO_2362 (O_2362,N_49260,N_48208);
nand UO_2363 (O_2363,N_49897,N_48524);
or UO_2364 (O_2364,N_48130,N_49660);
and UO_2365 (O_2365,N_49253,N_48783);
or UO_2366 (O_2366,N_48676,N_49166);
xor UO_2367 (O_2367,N_48054,N_49893);
nand UO_2368 (O_2368,N_48204,N_49735);
xor UO_2369 (O_2369,N_49110,N_49211);
and UO_2370 (O_2370,N_49746,N_49293);
and UO_2371 (O_2371,N_49735,N_48871);
nand UO_2372 (O_2372,N_48563,N_48732);
xnor UO_2373 (O_2373,N_49090,N_48177);
xor UO_2374 (O_2374,N_49152,N_48952);
nand UO_2375 (O_2375,N_49370,N_48885);
nand UO_2376 (O_2376,N_48869,N_48540);
nand UO_2377 (O_2377,N_48365,N_48011);
and UO_2378 (O_2378,N_48669,N_49492);
and UO_2379 (O_2379,N_49706,N_48096);
nand UO_2380 (O_2380,N_49910,N_48597);
xnor UO_2381 (O_2381,N_48279,N_49219);
nand UO_2382 (O_2382,N_48381,N_49000);
xor UO_2383 (O_2383,N_49553,N_49488);
xnor UO_2384 (O_2384,N_48697,N_49863);
nand UO_2385 (O_2385,N_48707,N_48187);
nor UO_2386 (O_2386,N_48726,N_49186);
or UO_2387 (O_2387,N_48641,N_48415);
nand UO_2388 (O_2388,N_48433,N_49329);
and UO_2389 (O_2389,N_48736,N_49327);
nor UO_2390 (O_2390,N_48076,N_49881);
nand UO_2391 (O_2391,N_48424,N_48351);
and UO_2392 (O_2392,N_49307,N_49209);
or UO_2393 (O_2393,N_48409,N_49724);
xor UO_2394 (O_2394,N_48584,N_48047);
nand UO_2395 (O_2395,N_49943,N_48269);
and UO_2396 (O_2396,N_48617,N_48107);
or UO_2397 (O_2397,N_48789,N_49456);
or UO_2398 (O_2398,N_49588,N_48663);
xor UO_2399 (O_2399,N_48584,N_49543);
and UO_2400 (O_2400,N_49936,N_49983);
or UO_2401 (O_2401,N_48270,N_49550);
and UO_2402 (O_2402,N_48287,N_48742);
nor UO_2403 (O_2403,N_49701,N_48262);
nor UO_2404 (O_2404,N_48668,N_48641);
nand UO_2405 (O_2405,N_48634,N_48104);
nor UO_2406 (O_2406,N_48740,N_49188);
and UO_2407 (O_2407,N_49124,N_49004);
and UO_2408 (O_2408,N_49085,N_48333);
or UO_2409 (O_2409,N_49538,N_48402);
nor UO_2410 (O_2410,N_48609,N_49704);
xor UO_2411 (O_2411,N_48205,N_49391);
nand UO_2412 (O_2412,N_49685,N_49131);
or UO_2413 (O_2413,N_48454,N_49629);
nor UO_2414 (O_2414,N_49724,N_49003);
xor UO_2415 (O_2415,N_49771,N_48013);
nand UO_2416 (O_2416,N_49568,N_48798);
nand UO_2417 (O_2417,N_49571,N_48265);
nand UO_2418 (O_2418,N_48905,N_49112);
xor UO_2419 (O_2419,N_48000,N_49532);
and UO_2420 (O_2420,N_49178,N_49290);
nor UO_2421 (O_2421,N_48468,N_49133);
xnor UO_2422 (O_2422,N_49011,N_48604);
nand UO_2423 (O_2423,N_48954,N_48786);
nand UO_2424 (O_2424,N_48236,N_49503);
nand UO_2425 (O_2425,N_49797,N_49447);
or UO_2426 (O_2426,N_48669,N_49858);
nor UO_2427 (O_2427,N_49808,N_48450);
or UO_2428 (O_2428,N_48064,N_49400);
nor UO_2429 (O_2429,N_48949,N_49941);
xor UO_2430 (O_2430,N_48773,N_48774);
nand UO_2431 (O_2431,N_48394,N_48420);
and UO_2432 (O_2432,N_49878,N_48998);
nor UO_2433 (O_2433,N_49009,N_49486);
or UO_2434 (O_2434,N_49647,N_49898);
or UO_2435 (O_2435,N_48235,N_48422);
nor UO_2436 (O_2436,N_49679,N_49312);
xor UO_2437 (O_2437,N_49815,N_49894);
xor UO_2438 (O_2438,N_48942,N_48099);
nand UO_2439 (O_2439,N_49722,N_48425);
nor UO_2440 (O_2440,N_49814,N_48265);
nand UO_2441 (O_2441,N_48143,N_48832);
xnor UO_2442 (O_2442,N_48191,N_49552);
nor UO_2443 (O_2443,N_49086,N_49645);
xor UO_2444 (O_2444,N_48513,N_48049);
or UO_2445 (O_2445,N_48754,N_49116);
and UO_2446 (O_2446,N_48276,N_49395);
and UO_2447 (O_2447,N_48148,N_49683);
and UO_2448 (O_2448,N_48905,N_48171);
nor UO_2449 (O_2449,N_49888,N_48972);
or UO_2450 (O_2450,N_49702,N_48205);
or UO_2451 (O_2451,N_48551,N_49909);
or UO_2452 (O_2452,N_48114,N_49565);
or UO_2453 (O_2453,N_48669,N_49473);
and UO_2454 (O_2454,N_49974,N_49193);
and UO_2455 (O_2455,N_48791,N_49739);
xnor UO_2456 (O_2456,N_48406,N_49464);
and UO_2457 (O_2457,N_49149,N_48071);
xor UO_2458 (O_2458,N_49574,N_48626);
or UO_2459 (O_2459,N_49772,N_49891);
nand UO_2460 (O_2460,N_49667,N_48573);
or UO_2461 (O_2461,N_49992,N_49545);
or UO_2462 (O_2462,N_49637,N_48075);
and UO_2463 (O_2463,N_49811,N_48471);
or UO_2464 (O_2464,N_48865,N_48538);
nor UO_2465 (O_2465,N_48259,N_49296);
nand UO_2466 (O_2466,N_49228,N_49138);
xor UO_2467 (O_2467,N_48656,N_49375);
nand UO_2468 (O_2468,N_49184,N_48143);
xor UO_2469 (O_2469,N_48043,N_48618);
or UO_2470 (O_2470,N_49481,N_48733);
and UO_2471 (O_2471,N_48486,N_49557);
xnor UO_2472 (O_2472,N_49966,N_49825);
xnor UO_2473 (O_2473,N_49554,N_48247);
nand UO_2474 (O_2474,N_48110,N_49305);
xnor UO_2475 (O_2475,N_48191,N_48101);
or UO_2476 (O_2476,N_49289,N_49822);
and UO_2477 (O_2477,N_49978,N_48946);
and UO_2478 (O_2478,N_48569,N_48665);
or UO_2479 (O_2479,N_49832,N_48952);
nor UO_2480 (O_2480,N_48924,N_49025);
nor UO_2481 (O_2481,N_48794,N_48280);
and UO_2482 (O_2482,N_48992,N_48813);
nor UO_2483 (O_2483,N_49238,N_49752);
nor UO_2484 (O_2484,N_48059,N_49582);
xnor UO_2485 (O_2485,N_49212,N_48264);
or UO_2486 (O_2486,N_48430,N_48061);
nor UO_2487 (O_2487,N_48999,N_49265);
or UO_2488 (O_2488,N_48288,N_49523);
nor UO_2489 (O_2489,N_48015,N_48266);
nor UO_2490 (O_2490,N_48463,N_49712);
or UO_2491 (O_2491,N_48878,N_49889);
nand UO_2492 (O_2492,N_49165,N_48357);
xor UO_2493 (O_2493,N_48461,N_49509);
nand UO_2494 (O_2494,N_49523,N_48041);
or UO_2495 (O_2495,N_49833,N_48052);
nand UO_2496 (O_2496,N_49979,N_49727);
or UO_2497 (O_2497,N_48610,N_48469);
nor UO_2498 (O_2498,N_48372,N_49732);
or UO_2499 (O_2499,N_48544,N_49575);
and UO_2500 (O_2500,N_49009,N_49989);
or UO_2501 (O_2501,N_48077,N_49830);
xor UO_2502 (O_2502,N_49429,N_49549);
nor UO_2503 (O_2503,N_48664,N_48345);
nand UO_2504 (O_2504,N_49689,N_48970);
xor UO_2505 (O_2505,N_48357,N_49227);
and UO_2506 (O_2506,N_48064,N_48571);
nand UO_2507 (O_2507,N_48456,N_48469);
nor UO_2508 (O_2508,N_48731,N_49427);
and UO_2509 (O_2509,N_49952,N_49199);
xnor UO_2510 (O_2510,N_48131,N_49772);
nor UO_2511 (O_2511,N_49014,N_48692);
or UO_2512 (O_2512,N_49320,N_49822);
nand UO_2513 (O_2513,N_48829,N_48155);
nor UO_2514 (O_2514,N_49554,N_48924);
nand UO_2515 (O_2515,N_48382,N_49923);
nand UO_2516 (O_2516,N_48640,N_48685);
nor UO_2517 (O_2517,N_48065,N_49445);
or UO_2518 (O_2518,N_48763,N_49668);
nor UO_2519 (O_2519,N_49346,N_48111);
or UO_2520 (O_2520,N_48293,N_48200);
or UO_2521 (O_2521,N_49807,N_49773);
nand UO_2522 (O_2522,N_49158,N_49273);
nand UO_2523 (O_2523,N_48514,N_48307);
nand UO_2524 (O_2524,N_48309,N_49779);
nor UO_2525 (O_2525,N_49530,N_49223);
xnor UO_2526 (O_2526,N_48083,N_49925);
xnor UO_2527 (O_2527,N_48754,N_48234);
or UO_2528 (O_2528,N_48168,N_49153);
xnor UO_2529 (O_2529,N_49554,N_49166);
nor UO_2530 (O_2530,N_49257,N_49404);
xor UO_2531 (O_2531,N_48887,N_49317);
or UO_2532 (O_2532,N_48752,N_48501);
or UO_2533 (O_2533,N_48982,N_48639);
or UO_2534 (O_2534,N_49059,N_48990);
or UO_2535 (O_2535,N_48643,N_49524);
or UO_2536 (O_2536,N_48522,N_48902);
xnor UO_2537 (O_2537,N_48621,N_48195);
nand UO_2538 (O_2538,N_48882,N_49118);
or UO_2539 (O_2539,N_48984,N_49711);
and UO_2540 (O_2540,N_49860,N_48612);
nor UO_2541 (O_2541,N_49710,N_49587);
xnor UO_2542 (O_2542,N_49255,N_48102);
or UO_2543 (O_2543,N_48671,N_49830);
or UO_2544 (O_2544,N_48847,N_49319);
nor UO_2545 (O_2545,N_48246,N_49309);
or UO_2546 (O_2546,N_48086,N_49222);
xnor UO_2547 (O_2547,N_48134,N_49282);
or UO_2548 (O_2548,N_48695,N_49902);
xor UO_2549 (O_2549,N_48694,N_49747);
nand UO_2550 (O_2550,N_48416,N_48812);
and UO_2551 (O_2551,N_48234,N_48766);
or UO_2552 (O_2552,N_48256,N_48956);
nand UO_2553 (O_2553,N_49886,N_48402);
xnor UO_2554 (O_2554,N_48259,N_48963);
and UO_2555 (O_2555,N_48559,N_48620);
and UO_2556 (O_2556,N_49745,N_49236);
xnor UO_2557 (O_2557,N_48468,N_48282);
and UO_2558 (O_2558,N_49101,N_48803);
and UO_2559 (O_2559,N_49992,N_49179);
or UO_2560 (O_2560,N_49226,N_48785);
nand UO_2561 (O_2561,N_49171,N_48709);
nand UO_2562 (O_2562,N_48228,N_48769);
nand UO_2563 (O_2563,N_48448,N_48187);
xor UO_2564 (O_2564,N_49871,N_49301);
nand UO_2565 (O_2565,N_49649,N_49259);
and UO_2566 (O_2566,N_49927,N_49940);
and UO_2567 (O_2567,N_49498,N_48597);
nor UO_2568 (O_2568,N_48184,N_49350);
nand UO_2569 (O_2569,N_49371,N_48757);
nor UO_2570 (O_2570,N_49848,N_49836);
or UO_2571 (O_2571,N_48653,N_49541);
or UO_2572 (O_2572,N_48673,N_48313);
and UO_2573 (O_2573,N_49375,N_49665);
and UO_2574 (O_2574,N_49978,N_49267);
nand UO_2575 (O_2575,N_49854,N_48257);
xor UO_2576 (O_2576,N_49972,N_49220);
and UO_2577 (O_2577,N_48872,N_48694);
or UO_2578 (O_2578,N_49060,N_48722);
nand UO_2579 (O_2579,N_48811,N_49600);
xor UO_2580 (O_2580,N_48483,N_49451);
nand UO_2581 (O_2581,N_48952,N_48356);
or UO_2582 (O_2582,N_49549,N_49050);
or UO_2583 (O_2583,N_49969,N_48690);
or UO_2584 (O_2584,N_48126,N_49604);
xnor UO_2585 (O_2585,N_49671,N_49597);
nor UO_2586 (O_2586,N_48436,N_48746);
xor UO_2587 (O_2587,N_49231,N_49600);
xnor UO_2588 (O_2588,N_49932,N_48276);
or UO_2589 (O_2589,N_48524,N_49128);
xor UO_2590 (O_2590,N_49788,N_48246);
nor UO_2591 (O_2591,N_48116,N_49505);
nand UO_2592 (O_2592,N_48094,N_48426);
and UO_2593 (O_2593,N_49952,N_48875);
nand UO_2594 (O_2594,N_48723,N_48935);
or UO_2595 (O_2595,N_49711,N_48442);
xor UO_2596 (O_2596,N_49141,N_48737);
nand UO_2597 (O_2597,N_48953,N_48982);
and UO_2598 (O_2598,N_49635,N_49041);
xnor UO_2599 (O_2599,N_49207,N_49377);
and UO_2600 (O_2600,N_49411,N_48417);
and UO_2601 (O_2601,N_48264,N_49035);
nor UO_2602 (O_2602,N_48324,N_48484);
and UO_2603 (O_2603,N_48538,N_49887);
xor UO_2604 (O_2604,N_49129,N_48313);
nand UO_2605 (O_2605,N_48400,N_49902);
nor UO_2606 (O_2606,N_49495,N_48364);
xnor UO_2607 (O_2607,N_49937,N_48660);
nand UO_2608 (O_2608,N_48847,N_49967);
xnor UO_2609 (O_2609,N_49267,N_49083);
xor UO_2610 (O_2610,N_48604,N_48622);
nand UO_2611 (O_2611,N_49223,N_49488);
and UO_2612 (O_2612,N_48299,N_49704);
nand UO_2613 (O_2613,N_49852,N_49636);
and UO_2614 (O_2614,N_48590,N_48599);
or UO_2615 (O_2615,N_49443,N_48216);
nand UO_2616 (O_2616,N_48363,N_48162);
and UO_2617 (O_2617,N_48434,N_49719);
nand UO_2618 (O_2618,N_49500,N_48810);
or UO_2619 (O_2619,N_49002,N_49690);
nor UO_2620 (O_2620,N_48251,N_49178);
nand UO_2621 (O_2621,N_48760,N_48532);
and UO_2622 (O_2622,N_49011,N_48391);
nor UO_2623 (O_2623,N_48406,N_48184);
xnor UO_2624 (O_2624,N_48440,N_48707);
xor UO_2625 (O_2625,N_48120,N_48052);
nand UO_2626 (O_2626,N_49645,N_49508);
and UO_2627 (O_2627,N_49188,N_49361);
nand UO_2628 (O_2628,N_48179,N_48283);
or UO_2629 (O_2629,N_48095,N_48759);
and UO_2630 (O_2630,N_48586,N_48130);
and UO_2631 (O_2631,N_49872,N_48792);
and UO_2632 (O_2632,N_49997,N_48053);
nand UO_2633 (O_2633,N_48254,N_48867);
xor UO_2634 (O_2634,N_49314,N_48227);
nor UO_2635 (O_2635,N_49882,N_49067);
or UO_2636 (O_2636,N_48217,N_48413);
nor UO_2637 (O_2637,N_49708,N_49198);
and UO_2638 (O_2638,N_49693,N_49779);
nand UO_2639 (O_2639,N_48177,N_49095);
nand UO_2640 (O_2640,N_49389,N_48775);
xor UO_2641 (O_2641,N_48123,N_48415);
and UO_2642 (O_2642,N_48974,N_48043);
or UO_2643 (O_2643,N_49601,N_49599);
and UO_2644 (O_2644,N_49698,N_49935);
nand UO_2645 (O_2645,N_49330,N_48687);
xnor UO_2646 (O_2646,N_48392,N_49142);
or UO_2647 (O_2647,N_49761,N_49183);
or UO_2648 (O_2648,N_48729,N_48144);
or UO_2649 (O_2649,N_48612,N_48657);
nand UO_2650 (O_2650,N_48910,N_49505);
and UO_2651 (O_2651,N_49220,N_49278);
nor UO_2652 (O_2652,N_49022,N_48013);
nor UO_2653 (O_2653,N_49523,N_49941);
or UO_2654 (O_2654,N_48062,N_49914);
or UO_2655 (O_2655,N_48962,N_48616);
nor UO_2656 (O_2656,N_48746,N_48215);
and UO_2657 (O_2657,N_48661,N_49909);
or UO_2658 (O_2658,N_49548,N_49181);
and UO_2659 (O_2659,N_48120,N_48339);
nand UO_2660 (O_2660,N_49609,N_48939);
nor UO_2661 (O_2661,N_49103,N_49738);
nor UO_2662 (O_2662,N_48163,N_48663);
xor UO_2663 (O_2663,N_49461,N_48385);
and UO_2664 (O_2664,N_48835,N_49284);
nor UO_2665 (O_2665,N_48646,N_48053);
xnor UO_2666 (O_2666,N_48652,N_49047);
and UO_2667 (O_2667,N_48052,N_48557);
and UO_2668 (O_2668,N_48779,N_49463);
xnor UO_2669 (O_2669,N_49109,N_49330);
nand UO_2670 (O_2670,N_49821,N_48622);
nand UO_2671 (O_2671,N_49585,N_48330);
nor UO_2672 (O_2672,N_49592,N_48059);
or UO_2673 (O_2673,N_49435,N_49575);
or UO_2674 (O_2674,N_48329,N_49305);
nand UO_2675 (O_2675,N_48096,N_48775);
xnor UO_2676 (O_2676,N_48654,N_48234);
or UO_2677 (O_2677,N_49766,N_49591);
nor UO_2678 (O_2678,N_48063,N_48926);
xor UO_2679 (O_2679,N_49932,N_49179);
xnor UO_2680 (O_2680,N_49353,N_49953);
nor UO_2681 (O_2681,N_49003,N_48285);
nor UO_2682 (O_2682,N_49781,N_48585);
and UO_2683 (O_2683,N_49166,N_49644);
or UO_2684 (O_2684,N_49784,N_49278);
and UO_2685 (O_2685,N_49289,N_49148);
and UO_2686 (O_2686,N_49653,N_49541);
or UO_2687 (O_2687,N_48214,N_49314);
or UO_2688 (O_2688,N_49002,N_49134);
or UO_2689 (O_2689,N_49254,N_48073);
or UO_2690 (O_2690,N_48282,N_48089);
nor UO_2691 (O_2691,N_49070,N_48764);
nor UO_2692 (O_2692,N_48398,N_49736);
xor UO_2693 (O_2693,N_49503,N_48704);
nor UO_2694 (O_2694,N_48166,N_48212);
and UO_2695 (O_2695,N_48555,N_48468);
nand UO_2696 (O_2696,N_48102,N_49033);
and UO_2697 (O_2697,N_48582,N_48329);
nor UO_2698 (O_2698,N_48813,N_48961);
xor UO_2699 (O_2699,N_49001,N_48595);
nand UO_2700 (O_2700,N_49495,N_49711);
and UO_2701 (O_2701,N_48964,N_49208);
xnor UO_2702 (O_2702,N_49223,N_48586);
and UO_2703 (O_2703,N_49710,N_48143);
nor UO_2704 (O_2704,N_49347,N_49392);
and UO_2705 (O_2705,N_48235,N_48153);
nand UO_2706 (O_2706,N_48492,N_48276);
nand UO_2707 (O_2707,N_48990,N_48512);
and UO_2708 (O_2708,N_49696,N_49601);
xnor UO_2709 (O_2709,N_48571,N_49133);
nand UO_2710 (O_2710,N_48210,N_48919);
or UO_2711 (O_2711,N_49786,N_49799);
xor UO_2712 (O_2712,N_49495,N_49905);
nor UO_2713 (O_2713,N_49414,N_49013);
xor UO_2714 (O_2714,N_48688,N_48718);
or UO_2715 (O_2715,N_49924,N_48375);
and UO_2716 (O_2716,N_48881,N_48481);
xor UO_2717 (O_2717,N_48217,N_49649);
nand UO_2718 (O_2718,N_48259,N_48101);
and UO_2719 (O_2719,N_48643,N_49068);
or UO_2720 (O_2720,N_48933,N_48546);
and UO_2721 (O_2721,N_48789,N_49430);
or UO_2722 (O_2722,N_49256,N_48514);
or UO_2723 (O_2723,N_48544,N_49765);
nand UO_2724 (O_2724,N_48165,N_48245);
nand UO_2725 (O_2725,N_49156,N_48362);
nor UO_2726 (O_2726,N_48156,N_48165);
or UO_2727 (O_2727,N_49754,N_49809);
and UO_2728 (O_2728,N_48892,N_48108);
xnor UO_2729 (O_2729,N_48247,N_49195);
nor UO_2730 (O_2730,N_49143,N_49074);
or UO_2731 (O_2731,N_49093,N_49145);
or UO_2732 (O_2732,N_49856,N_49641);
and UO_2733 (O_2733,N_48183,N_48864);
nand UO_2734 (O_2734,N_48488,N_49855);
nor UO_2735 (O_2735,N_49503,N_49751);
nand UO_2736 (O_2736,N_49769,N_49468);
nand UO_2737 (O_2737,N_48661,N_49232);
and UO_2738 (O_2738,N_48245,N_48520);
nand UO_2739 (O_2739,N_49340,N_49393);
nand UO_2740 (O_2740,N_49593,N_48745);
xnor UO_2741 (O_2741,N_48051,N_49187);
nor UO_2742 (O_2742,N_48650,N_49640);
xnor UO_2743 (O_2743,N_48975,N_48415);
or UO_2744 (O_2744,N_49996,N_49163);
or UO_2745 (O_2745,N_49831,N_49198);
or UO_2746 (O_2746,N_48117,N_49850);
xor UO_2747 (O_2747,N_49901,N_48769);
nand UO_2748 (O_2748,N_49566,N_48050);
xor UO_2749 (O_2749,N_49168,N_49611);
xnor UO_2750 (O_2750,N_49397,N_49885);
nand UO_2751 (O_2751,N_48846,N_49013);
and UO_2752 (O_2752,N_48408,N_49927);
nand UO_2753 (O_2753,N_49157,N_48779);
or UO_2754 (O_2754,N_48532,N_48860);
and UO_2755 (O_2755,N_49656,N_48965);
and UO_2756 (O_2756,N_49890,N_48707);
xor UO_2757 (O_2757,N_48079,N_49173);
or UO_2758 (O_2758,N_49187,N_48356);
or UO_2759 (O_2759,N_49564,N_48557);
and UO_2760 (O_2760,N_48599,N_49458);
or UO_2761 (O_2761,N_49539,N_49564);
or UO_2762 (O_2762,N_49213,N_49326);
and UO_2763 (O_2763,N_49715,N_48225);
or UO_2764 (O_2764,N_49252,N_48330);
and UO_2765 (O_2765,N_49590,N_48290);
nor UO_2766 (O_2766,N_49944,N_48036);
and UO_2767 (O_2767,N_48511,N_48645);
nand UO_2768 (O_2768,N_48952,N_49998);
nand UO_2769 (O_2769,N_49692,N_48701);
or UO_2770 (O_2770,N_49508,N_48165);
nand UO_2771 (O_2771,N_48203,N_49737);
and UO_2772 (O_2772,N_49411,N_49505);
xnor UO_2773 (O_2773,N_49453,N_49783);
or UO_2774 (O_2774,N_49424,N_48598);
or UO_2775 (O_2775,N_49828,N_48988);
xnor UO_2776 (O_2776,N_49976,N_49486);
or UO_2777 (O_2777,N_49772,N_49423);
or UO_2778 (O_2778,N_48809,N_48863);
xor UO_2779 (O_2779,N_48312,N_48724);
nand UO_2780 (O_2780,N_49318,N_48053);
xor UO_2781 (O_2781,N_49228,N_49253);
and UO_2782 (O_2782,N_48639,N_49687);
or UO_2783 (O_2783,N_48917,N_49215);
xnor UO_2784 (O_2784,N_49524,N_48101);
xor UO_2785 (O_2785,N_48456,N_48685);
xor UO_2786 (O_2786,N_49828,N_49456);
xnor UO_2787 (O_2787,N_48267,N_49831);
nand UO_2788 (O_2788,N_48113,N_49751);
and UO_2789 (O_2789,N_48121,N_49704);
and UO_2790 (O_2790,N_49475,N_49260);
and UO_2791 (O_2791,N_48585,N_48453);
nand UO_2792 (O_2792,N_49074,N_48658);
or UO_2793 (O_2793,N_49956,N_48371);
xnor UO_2794 (O_2794,N_49088,N_49849);
xor UO_2795 (O_2795,N_48964,N_49823);
or UO_2796 (O_2796,N_48440,N_48766);
xor UO_2797 (O_2797,N_48366,N_48065);
and UO_2798 (O_2798,N_48193,N_49846);
nor UO_2799 (O_2799,N_49037,N_49731);
nand UO_2800 (O_2800,N_48304,N_49775);
xor UO_2801 (O_2801,N_49525,N_49585);
nand UO_2802 (O_2802,N_49581,N_48721);
nand UO_2803 (O_2803,N_49703,N_48572);
and UO_2804 (O_2804,N_49866,N_49750);
or UO_2805 (O_2805,N_48070,N_49455);
and UO_2806 (O_2806,N_48613,N_48269);
or UO_2807 (O_2807,N_49448,N_49060);
nand UO_2808 (O_2808,N_49385,N_48101);
xor UO_2809 (O_2809,N_49153,N_48496);
xnor UO_2810 (O_2810,N_49494,N_48562);
nor UO_2811 (O_2811,N_48345,N_49278);
nand UO_2812 (O_2812,N_48851,N_48830);
xnor UO_2813 (O_2813,N_49438,N_48919);
or UO_2814 (O_2814,N_49749,N_48897);
nor UO_2815 (O_2815,N_48227,N_48455);
and UO_2816 (O_2816,N_48587,N_49169);
and UO_2817 (O_2817,N_48841,N_48329);
nand UO_2818 (O_2818,N_49547,N_48987);
and UO_2819 (O_2819,N_49017,N_49165);
or UO_2820 (O_2820,N_48374,N_49797);
nand UO_2821 (O_2821,N_48749,N_49138);
nand UO_2822 (O_2822,N_49117,N_48150);
or UO_2823 (O_2823,N_49237,N_49660);
nor UO_2824 (O_2824,N_48801,N_48266);
nand UO_2825 (O_2825,N_48170,N_48305);
nand UO_2826 (O_2826,N_49375,N_49817);
or UO_2827 (O_2827,N_48767,N_49951);
and UO_2828 (O_2828,N_49562,N_48004);
or UO_2829 (O_2829,N_49009,N_48970);
xor UO_2830 (O_2830,N_49259,N_49755);
or UO_2831 (O_2831,N_49257,N_49475);
nand UO_2832 (O_2832,N_48798,N_49004);
or UO_2833 (O_2833,N_49035,N_49150);
nor UO_2834 (O_2834,N_49512,N_49006);
nand UO_2835 (O_2835,N_49246,N_48779);
nand UO_2836 (O_2836,N_48068,N_49757);
and UO_2837 (O_2837,N_49370,N_49402);
or UO_2838 (O_2838,N_48154,N_49141);
nand UO_2839 (O_2839,N_49744,N_49901);
nor UO_2840 (O_2840,N_49375,N_48265);
or UO_2841 (O_2841,N_49141,N_49608);
nand UO_2842 (O_2842,N_48170,N_48825);
and UO_2843 (O_2843,N_48572,N_48770);
xor UO_2844 (O_2844,N_49794,N_49248);
xor UO_2845 (O_2845,N_49205,N_49357);
nand UO_2846 (O_2846,N_48848,N_49278);
nor UO_2847 (O_2847,N_49370,N_49231);
nor UO_2848 (O_2848,N_48077,N_49233);
and UO_2849 (O_2849,N_49782,N_49356);
and UO_2850 (O_2850,N_49439,N_49442);
xnor UO_2851 (O_2851,N_49885,N_49860);
nand UO_2852 (O_2852,N_49503,N_49723);
xnor UO_2853 (O_2853,N_48064,N_48828);
nor UO_2854 (O_2854,N_49877,N_48948);
nor UO_2855 (O_2855,N_49757,N_49176);
nand UO_2856 (O_2856,N_48208,N_48094);
nand UO_2857 (O_2857,N_48708,N_48415);
or UO_2858 (O_2858,N_49192,N_48307);
nor UO_2859 (O_2859,N_48328,N_48222);
or UO_2860 (O_2860,N_49358,N_49567);
xnor UO_2861 (O_2861,N_48690,N_49194);
nand UO_2862 (O_2862,N_49489,N_49318);
and UO_2863 (O_2863,N_48707,N_48973);
nor UO_2864 (O_2864,N_48741,N_49286);
nand UO_2865 (O_2865,N_48414,N_48609);
nand UO_2866 (O_2866,N_48676,N_49209);
nand UO_2867 (O_2867,N_49430,N_49492);
xnor UO_2868 (O_2868,N_48971,N_48002);
or UO_2869 (O_2869,N_49627,N_49135);
xor UO_2870 (O_2870,N_48438,N_49228);
or UO_2871 (O_2871,N_48257,N_49700);
or UO_2872 (O_2872,N_49199,N_49779);
xnor UO_2873 (O_2873,N_48069,N_48409);
nand UO_2874 (O_2874,N_48657,N_48621);
or UO_2875 (O_2875,N_48953,N_49545);
nand UO_2876 (O_2876,N_48569,N_49124);
nand UO_2877 (O_2877,N_49663,N_49615);
xnor UO_2878 (O_2878,N_49400,N_48693);
nor UO_2879 (O_2879,N_48381,N_48408);
nor UO_2880 (O_2880,N_48720,N_49081);
nand UO_2881 (O_2881,N_48587,N_48602);
and UO_2882 (O_2882,N_49352,N_48197);
xnor UO_2883 (O_2883,N_48426,N_49221);
or UO_2884 (O_2884,N_48875,N_48508);
and UO_2885 (O_2885,N_48226,N_48083);
and UO_2886 (O_2886,N_48522,N_49788);
xor UO_2887 (O_2887,N_49322,N_48719);
and UO_2888 (O_2888,N_48993,N_48920);
and UO_2889 (O_2889,N_49338,N_48327);
nand UO_2890 (O_2890,N_48811,N_49131);
and UO_2891 (O_2891,N_48665,N_48315);
or UO_2892 (O_2892,N_49169,N_49290);
and UO_2893 (O_2893,N_48378,N_49484);
nand UO_2894 (O_2894,N_49582,N_49096);
and UO_2895 (O_2895,N_48803,N_49075);
nor UO_2896 (O_2896,N_48770,N_49136);
and UO_2897 (O_2897,N_48555,N_48294);
nand UO_2898 (O_2898,N_49166,N_49494);
xor UO_2899 (O_2899,N_49362,N_48682);
nor UO_2900 (O_2900,N_49289,N_48224);
nand UO_2901 (O_2901,N_48990,N_49208);
nand UO_2902 (O_2902,N_49590,N_48826);
xor UO_2903 (O_2903,N_49675,N_48157);
nand UO_2904 (O_2904,N_48214,N_48395);
nand UO_2905 (O_2905,N_48644,N_48327);
nor UO_2906 (O_2906,N_49597,N_48901);
xor UO_2907 (O_2907,N_49374,N_49091);
or UO_2908 (O_2908,N_49688,N_49298);
xor UO_2909 (O_2909,N_48721,N_48694);
and UO_2910 (O_2910,N_48223,N_49326);
nand UO_2911 (O_2911,N_48370,N_49016);
nand UO_2912 (O_2912,N_49808,N_49224);
nand UO_2913 (O_2913,N_48293,N_48984);
nand UO_2914 (O_2914,N_49084,N_48466);
xnor UO_2915 (O_2915,N_48385,N_49602);
nand UO_2916 (O_2916,N_48730,N_48520);
xnor UO_2917 (O_2917,N_48901,N_49242);
xnor UO_2918 (O_2918,N_49450,N_48666);
nor UO_2919 (O_2919,N_49164,N_49156);
nand UO_2920 (O_2920,N_48182,N_49440);
xnor UO_2921 (O_2921,N_48360,N_48874);
nand UO_2922 (O_2922,N_48220,N_49598);
and UO_2923 (O_2923,N_49196,N_49390);
nand UO_2924 (O_2924,N_49519,N_49088);
and UO_2925 (O_2925,N_49111,N_48646);
nor UO_2926 (O_2926,N_48403,N_48671);
nand UO_2927 (O_2927,N_48598,N_48225);
nand UO_2928 (O_2928,N_49793,N_48678);
nand UO_2929 (O_2929,N_49267,N_48317);
nor UO_2930 (O_2930,N_48003,N_49674);
xor UO_2931 (O_2931,N_48729,N_49283);
nor UO_2932 (O_2932,N_49873,N_49228);
nand UO_2933 (O_2933,N_49448,N_48253);
and UO_2934 (O_2934,N_48281,N_49202);
nand UO_2935 (O_2935,N_49895,N_49378);
xor UO_2936 (O_2936,N_48712,N_49761);
and UO_2937 (O_2937,N_48523,N_48670);
or UO_2938 (O_2938,N_49998,N_48511);
xor UO_2939 (O_2939,N_48256,N_48556);
and UO_2940 (O_2940,N_48685,N_49444);
nor UO_2941 (O_2941,N_49163,N_49188);
xnor UO_2942 (O_2942,N_49946,N_48431);
xor UO_2943 (O_2943,N_48962,N_48965);
xor UO_2944 (O_2944,N_49686,N_48949);
nor UO_2945 (O_2945,N_48182,N_49064);
xnor UO_2946 (O_2946,N_48634,N_48601);
nor UO_2947 (O_2947,N_49136,N_49773);
xnor UO_2948 (O_2948,N_48162,N_49472);
and UO_2949 (O_2949,N_48181,N_48189);
nand UO_2950 (O_2950,N_48721,N_48606);
or UO_2951 (O_2951,N_48703,N_48809);
nor UO_2952 (O_2952,N_48618,N_48492);
nand UO_2953 (O_2953,N_48780,N_49294);
or UO_2954 (O_2954,N_48423,N_48206);
nor UO_2955 (O_2955,N_48558,N_49700);
nand UO_2956 (O_2956,N_49259,N_49408);
and UO_2957 (O_2957,N_49591,N_48731);
nor UO_2958 (O_2958,N_48378,N_48450);
and UO_2959 (O_2959,N_49239,N_48961);
xnor UO_2960 (O_2960,N_48982,N_48022);
and UO_2961 (O_2961,N_48301,N_49435);
and UO_2962 (O_2962,N_49891,N_49031);
nor UO_2963 (O_2963,N_49212,N_48655);
and UO_2964 (O_2964,N_49880,N_49588);
nor UO_2965 (O_2965,N_48359,N_49714);
xor UO_2966 (O_2966,N_49416,N_48960);
xor UO_2967 (O_2967,N_49751,N_49276);
xnor UO_2968 (O_2968,N_49630,N_48997);
and UO_2969 (O_2969,N_48842,N_48275);
nor UO_2970 (O_2970,N_49608,N_49514);
nor UO_2971 (O_2971,N_49172,N_49364);
and UO_2972 (O_2972,N_49247,N_48545);
nor UO_2973 (O_2973,N_48210,N_48476);
nand UO_2974 (O_2974,N_48167,N_49165);
nor UO_2975 (O_2975,N_49981,N_48509);
xnor UO_2976 (O_2976,N_49020,N_48125);
nor UO_2977 (O_2977,N_49144,N_48938);
xor UO_2978 (O_2978,N_49763,N_48935);
nand UO_2979 (O_2979,N_49578,N_49864);
and UO_2980 (O_2980,N_49839,N_49444);
nand UO_2981 (O_2981,N_49847,N_48377);
nand UO_2982 (O_2982,N_48179,N_48305);
nand UO_2983 (O_2983,N_48220,N_48811);
xor UO_2984 (O_2984,N_48754,N_48575);
nor UO_2985 (O_2985,N_49462,N_48774);
xor UO_2986 (O_2986,N_49521,N_49800);
or UO_2987 (O_2987,N_49175,N_49430);
and UO_2988 (O_2988,N_49008,N_49989);
xor UO_2989 (O_2989,N_48922,N_49238);
nor UO_2990 (O_2990,N_48009,N_49977);
and UO_2991 (O_2991,N_49897,N_48527);
nand UO_2992 (O_2992,N_49125,N_49847);
nand UO_2993 (O_2993,N_48296,N_49893);
xor UO_2994 (O_2994,N_49245,N_49270);
xor UO_2995 (O_2995,N_49232,N_48682);
xnor UO_2996 (O_2996,N_48205,N_48257);
or UO_2997 (O_2997,N_49216,N_48503);
xnor UO_2998 (O_2998,N_48776,N_48578);
xnor UO_2999 (O_2999,N_48506,N_49449);
or UO_3000 (O_3000,N_48982,N_49499);
nor UO_3001 (O_3001,N_49072,N_48260);
xor UO_3002 (O_3002,N_48843,N_48338);
nor UO_3003 (O_3003,N_49235,N_49609);
and UO_3004 (O_3004,N_48173,N_48983);
xnor UO_3005 (O_3005,N_49197,N_48101);
and UO_3006 (O_3006,N_48166,N_48261);
nor UO_3007 (O_3007,N_49648,N_49762);
nand UO_3008 (O_3008,N_48864,N_48480);
and UO_3009 (O_3009,N_48446,N_49615);
nand UO_3010 (O_3010,N_48363,N_48842);
nor UO_3011 (O_3011,N_49644,N_49756);
or UO_3012 (O_3012,N_49297,N_49618);
and UO_3013 (O_3013,N_48425,N_48204);
nand UO_3014 (O_3014,N_49244,N_49631);
xnor UO_3015 (O_3015,N_49465,N_48381);
or UO_3016 (O_3016,N_48412,N_49821);
nor UO_3017 (O_3017,N_49465,N_48602);
xnor UO_3018 (O_3018,N_49720,N_49831);
nor UO_3019 (O_3019,N_48391,N_48295);
nand UO_3020 (O_3020,N_48525,N_49954);
and UO_3021 (O_3021,N_48175,N_48000);
nand UO_3022 (O_3022,N_48720,N_48378);
nor UO_3023 (O_3023,N_49826,N_49140);
nor UO_3024 (O_3024,N_48279,N_49203);
nor UO_3025 (O_3025,N_48585,N_48224);
or UO_3026 (O_3026,N_49423,N_49928);
xnor UO_3027 (O_3027,N_49230,N_49171);
nand UO_3028 (O_3028,N_48104,N_49696);
nand UO_3029 (O_3029,N_48839,N_49387);
nand UO_3030 (O_3030,N_48528,N_49813);
and UO_3031 (O_3031,N_48994,N_49938);
nand UO_3032 (O_3032,N_48222,N_49546);
nor UO_3033 (O_3033,N_48412,N_49399);
and UO_3034 (O_3034,N_48672,N_48489);
nand UO_3035 (O_3035,N_49887,N_49778);
xnor UO_3036 (O_3036,N_49916,N_49321);
nor UO_3037 (O_3037,N_49856,N_48303);
and UO_3038 (O_3038,N_48254,N_48628);
xnor UO_3039 (O_3039,N_49779,N_48691);
nand UO_3040 (O_3040,N_48070,N_48094);
or UO_3041 (O_3041,N_49405,N_48908);
nor UO_3042 (O_3042,N_49035,N_49325);
nor UO_3043 (O_3043,N_49659,N_49460);
or UO_3044 (O_3044,N_49114,N_49951);
and UO_3045 (O_3045,N_49242,N_48657);
or UO_3046 (O_3046,N_48341,N_49766);
nor UO_3047 (O_3047,N_48593,N_48770);
or UO_3048 (O_3048,N_48689,N_49653);
nand UO_3049 (O_3049,N_49167,N_48225);
nand UO_3050 (O_3050,N_49131,N_48488);
nand UO_3051 (O_3051,N_48205,N_48747);
or UO_3052 (O_3052,N_49156,N_49073);
and UO_3053 (O_3053,N_49123,N_48631);
and UO_3054 (O_3054,N_49346,N_49392);
nor UO_3055 (O_3055,N_48530,N_48707);
or UO_3056 (O_3056,N_48561,N_49799);
or UO_3057 (O_3057,N_48536,N_48503);
or UO_3058 (O_3058,N_48534,N_48976);
xnor UO_3059 (O_3059,N_48782,N_49352);
xnor UO_3060 (O_3060,N_48895,N_48687);
and UO_3061 (O_3061,N_49190,N_49669);
nand UO_3062 (O_3062,N_48697,N_49505);
xor UO_3063 (O_3063,N_49723,N_48815);
or UO_3064 (O_3064,N_49687,N_49187);
or UO_3065 (O_3065,N_48879,N_48886);
and UO_3066 (O_3066,N_48112,N_48928);
and UO_3067 (O_3067,N_48717,N_49885);
nand UO_3068 (O_3068,N_48839,N_49964);
nand UO_3069 (O_3069,N_49040,N_48442);
or UO_3070 (O_3070,N_49054,N_49938);
xor UO_3071 (O_3071,N_48915,N_48649);
nand UO_3072 (O_3072,N_49318,N_49897);
and UO_3073 (O_3073,N_49792,N_49461);
and UO_3074 (O_3074,N_49769,N_49881);
and UO_3075 (O_3075,N_48055,N_48900);
nand UO_3076 (O_3076,N_48730,N_49550);
nor UO_3077 (O_3077,N_48801,N_49732);
nand UO_3078 (O_3078,N_48977,N_49237);
nand UO_3079 (O_3079,N_48447,N_48842);
nor UO_3080 (O_3080,N_48432,N_49940);
and UO_3081 (O_3081,N_48290,N_49424);
nor UO_3082 (O_3082,N_49668,N_48305);
and UO_3083 (O_3083,N_48595,N_48326);
and UO_3084 (O_3084,N_49940,N_49419);
nor UO_3085 (O_3085,N_49433,N_49242);
and UO_3086 (O_3086,N_48323,N_49542);
nor UO_3087 (O_3087,N_48669,N_49255);
and UO_3088 (O_3088,N_49718,N_49879);
and UO_3089 (O_3089,N_49237,N_49373);
nand UO_3090 (O_3090,N_48076,N_49595);
nand UO_3091 (O_3091,N_49176,N_49241);
nor UO_3092 (O_3092,N_48869,N_48864);
or UO_3093 (O_3093,N_48018,N_48689);
xnor UO_3094 (O_3094,N_49292,N_48669);
or UO_3095 (O_3095,N_48225,N_49863);
nor UO_3096 (O_3096,N_48591,N_49283);
or UO_3097 (O_3097,N_48222,N_49996);
or UO_3098 (O_3098,N_49033,N_48254);
xnor UO_3099 (O_3099,N_48923,N_49938);
or UO_3100 (O_3100,N_49464,N_49776);
or UO_3101 (O_3101,N_49343,N_48532);
nand UO_3102 (O_3102,N_49665,N_49179);
and UO_3103 (O_3103,N_48709,N_49669);
nand UO_3104 (O_3104,N_48011,N_48051);
nand UO_3105 (O_3105,N_49351,N_49563);
and UO_3106 (O_3106,N_49539,N_49094);
nand UO_3107 (O_3107,N_49301,N_48005);
xor UO_3108 (O_3108,N_49416,N_49327);
nand UO_3109 (O_3109,N_49171,N_48973);
nor UO_3110 (O_3110,N_48321,N_49585);
or UO_3111 (O_3111,N_48226,N_49860);
and UO_3112 (O_3112,N_49827,N_49253);
nor UO_3113 (O_3113,N_49753,N_48539);
xnor UO_3114 (O_3114,N_48174,N_49014);
xor UO_3115 (O_3115,N_49039,N_48169);
xnor UO_3116 (O_3116,N_49354,N_49618);
nor UO_3117 (O_3117,N_48287,N_48660);
nand UO_3118 (O_3118,N_49032,N_48902);
xnor UO_3119 (O_3119,N_48290,N_48424);
and UO_3120 (O_3120,N_49309,N_48271);
nand UO_3121 (O_3121,N_49813,N_49009);
nor UO_3122 (O_3122,N_48980,N_49512);
xor UO_3123 (O_3123,N_48152,N_48768);
or UO_3124 (O_3124,N_49260,N_49468);
nor UO_3125 (O_3125,N_48338,N_48540);
nor UO_3126 (O_3126,N_49277,N_49309);
xor UO_3127 (O_3127,N_48216,N_49709);
and UO_3128 (O_3128,N_49546,N_49243);
nand UO_3129 (O_3129,N_48860,N_49287);
or UO_3130 (O_3130,N_48256,N_48985);
nand UO_3131 (O_3131,N_49911,N_48231);
nor UO_3132 (O_3132,N_48822,N_48390);
or UO_3133 (O_3133,N_49581,N_49679);
nor UO_3134 (O_3134,N_49102,N_48593);
and UO_3135 (O_3135,N_49376,N_48909);
nand UO_3136 (O_3136,N_48835,N_49025);
nor UO_3137 (O_3137,N_49391,N_48460);
and UO_3138 (O_3138,N_48041,N_49935);
or UO_3139 (O_3139,N_49164,N_49653);
nand UO_3140 (O_3140,N_48038,N_49141);
and UO_3141 (O_3141,N_49418,N_49036);
nor UO_3142 (O_3142,N_49545,N_49517);
nor UO_3143 (O_3143,N_49300,N_49157);
or UO_3144 (O_3144,N_48989,N_49014);
or UO_3145 (O_3145,N_48428,N_49531);
xnor UO_3146 (O_3146,N_48820,N_49783);
nand UO_3147 (O_3147,N_49911,N_49857);
xnor UO_3148 (O_3148,N_49026,N_48608);
or UO_3149 (O_3149,N_49621,N_49995);
nor UO_3150 (O_3150,N_48968,N_48076);
nand UO_3151 (O_3151,N_49024,N_48170);
or UO_3152 (O_3152,N_49135,N_49923);
nand UO_3153 (O_3153,N_48034,N_49474);
nor UO_3154 (O_3154,N_49617,N_48493);
xnor UO_3155 (O_3155,N_49767,N_48528);
xor UO_3156 (O_3156,N_49997,N_49424);
nand UO_3157 (O_3157,N_48685,N_49142);
and UO_3158 (O_3158,N_49964,N_48132);
or UO_3159 (O_3159,N_49725,N_49163);
xnor UO_3160 (O_3160,N_49147,N_48158);
nor UO_3161 (O_3161,N_49387,N_49229);
and UO_3162 (O_3162,N_49469,N_48085);
and UO_3163 (O_3163,N_48662,N_49892);
or UO_3164 (O_3164,N_48284,N_48073);
and UO_3165 (O_3165,N_49796,N_49601);
nor UO_3166 (O_3166,N_48182,N_49449);
nor UO_3167 (O_3167,N_48207,N_49444);
xor UO_3168 (O_3168,N_48543,N_49457);
or UO_3169 (O_3169,N_49353,N_49986);
or UO_3170 (O_3170,N_49037,N_48261);
and UO_3171 (O_3171,N_49717,N_48873);
nand UO_3172 (O_3172,N_48303,N_49649);
and UO_3173 (O_3173,N_49289,N_49472);
and UO_3174 (O_3174,N_48868,N_48904);
nand UO_3175 (O_3175,N_48394,N_49116);
nor UO_3176 (O_3176,N_48482,N_49551);
and UO_3177 (O_3177,N_49091,N_49625);
xor UO_3178 (O_3178,N_48358,N_49378);
nand UO_3179 (O_3179,N_49774,N_48378);
or UO_3180 (O_3180,N_48867,N_48707);
xor UO_3181 (O_3181,N_48918,N_49657);
nor UO_3182 (O_3182,N_48738,N_48525);
and UO_3183 (O_3183,N_49549,N_48501);
xor UO_3184 (O_3184,N_49451,N_49103);
and UO_3185 (O_3185,N_49588,N_49057);
nor UO_3186 (O_3186,N_49865,N_48149);
xor UO_3187 (O_3187,N_48197,N_49714);
or UO_3188 (O_3188,N_48123,N_48668);
nand UO_3189 (O_3189,N_48116,N_48728);
nor UO_3190 (O_3190,N_49901,N_48380);
xor UO_3191 (O_3191,N_48059,N_48336);
nor UO_3192 (O_3192,N_49494,N_48125);
nand UO_3193 (O_3193,N_48234,N_49721);
nor UO_3194 (O_3194,N_48744,N_49883);
xor UO_3195 (O_3195,N_49517,N_49543);
and UO_3196 (O_3196,N_49839,N_48700);
or UO_3197 (O_3197,N_49698,N_48776);
and UO_3198 (O_3198,N_48934,N_49658);
nand UO_3199 (O_3199,N_49849,N_49901);
nand UO_3200 (O_3200,N_48141,N_48424);
nor UO_3201 (O_3201,N_48357,N_48270);
and UO_3202 (O_3202,N_49833,N_48307);
and UO_3203 (O_3203,N_49288,N_49826);
or UO_3204 (O_3204,N_48087,N_48417);
nor UO_3205 (O_3205,N_49521,N_49915);
and UO_3206 (O_3206,N_48173,N_48220);
or UO_3207 (O_3207,N_49671,N_49363);
or UO_3208 (O_3208,N_49814,N_48312);
and UO_3209 (O_3209,N_49960,N_49608);
and UO_3210 (O_3210,N_49548,N_49686);
nand UO_3211 (O_3211,N_49008,N_49827);
nand UO_3212 (O_3212,N_49954,N_49461);
nand UO_3213 (O_3213,N_48500,N_48652);
and UO_3214 (O_3214,N_48559,N_49429);
xnor UO_3215 (O_3215,N_49929,N_48197);
nand UO_3216 (O_3216,N_48145,N_48533);
nand UO_3217 (O_3217,N_49529,N_49771);
and UO_3218 (O_3218,N_49738,N_48672);
nor UO_3219 (O_3219,N_48734,N_49864);
and UO_3220 (O_3220,N_49754,N_48868);
or UO_3221 (O_3221,N_49525,N_48928);
or UO_3222 (O_3222,N_48292,N_48314);
and UO_3223 (O_3223,N_49394,N_49182);
nor UO_3224 (O_3224,N_48157,N_49807);
nor UO_3225 (O_3225,N_49109,N_48119);
nor UO_3226 (O_3226,N_48512,N_49321);
nand UO_3227 (O_3227,N_48603,N_49304);
nor UO_3228 (O_3228,N_48033,N_48848);
or UO_3229 (O_3229,N_48563,N_48781);
or UO_3230 (O_3230,N_49911,N_48720);
nor UO_3231 (O_3231,N_49514,N_48421);
xor UO_3232 (O_3232,N_49950,N_48710);
and UO_3233 (O_3233,N_48186,N_49875);
xnor UO_3234 (O_3234,N_48552,N_49813);
nand UO_3235 (O_3235,N_49381,N_49047);
xor UO_3236 (O_3236,N_48225,N_48290);
nor UO_3237 (O_3237,N_49845,N_48827);
nand UO_3238 (O_3238,N_48927,N_49318);
nor UO_3239 (O_3239,N_48020,N_49844);
nand UO_3240 (O_3240,N_48639,N_48989);
and UO_3241 (O_3241,N_48071,N_48628);
nand UO_3242 (O_3242,N_48534,N_48686);
xor UO_3243 (O_3243,N_49454,N_49605);
xnor UO_3244 (O_3244,N_49345,N_48459);
or UO_3245 (O_3245,N_48421,N_48302);
nand UO_3246 (O_3246,N_49438,N_49522);
nor UO_3247 (O_3247,N_48722,N_48606);
nor UO_3248 (O_3248,N_49541,N_49004);
or UO_3249 (O_3249,N_48885,N_48796);
nand UO_3250 (O_3250,N_49478,N_48114);
xnor UO_3251 (O_3251,N_48686,N_49514);
nand UO_3252 (O_3252,N_48598,N_49027);
nand UO_3253 (O_3253,N_49641,N_49976);
nor UO_3254 (O_3254,N_48284,N_48789);
or UO_3255 (O_3255,N_48340,N_49044);
nand UO_3256 (O_3256,N_48618,N_49913);
nand UO_3257 (O_3257,N_49305,N_49830);
nand UO_3258 (O_3258,N_49551,N_48363);
nor UO_3259 (O_3259,N_49222,N_48348);
and UO_3260 (O_3260,N_49686,N_49212);
nand UO_3261 (O_3261,N_49722,N_49715);
xor UO_3262 (O_3262,N_48324,N_48851);
and UO_3263 (O_3263,N_49705,N_48210);
or UO_3264 (O_3264,N_48084,N_48053);
or UO_3265 (O_3265,N_48504,N_48997);
xnor UO_3266 (O_3266,N_49721,N_49436);
and UO_3267 (O_3267,N_48758,N_49429);
nand UO_3268 (O_3268,N_49876,N_49074);
xnor UO_3269 (O_3269,N_48024,N_49889);
nand UO_3270 (O_3270,N_49906,N_49402);
xnor UO_3271 (O_3271,N_49820,N_49306);
nand UO_3272 (O_3272,N_48607,N_48677);
nor UO_3273 (O_3273,N_48788,N_48639);
nor UO_3274 (O_3274,N_49317,N_48031);
xnor UO_3275 (O_3275,N_49612,N_49453);
and UO_3276 (O_3276,N_49863,N_49161);
nand UO_3277 (O_3277,N_49088,N_49468);
or UO_3278 (O_3278,N_49334,N_48077);
and UO_3279 (O_3279,N_49199,N_49473);
nor UO_3280 (O_3280,N_49184,N_48691);
nor UO_3281 (O_3281,N_49609,N_48374);
nand UO_3282 (O_3282,N_48600,N_49742);
or UO_3283 (O_3283,N_48340,N_49239);
and UO_3284 (O_3284,N_48603,N_48150);
and UO_3285 (O_3285,N_48210,N_48069);
nand UO_3286 (O_3286,N_48500,N_49989);
nor UO_3287 (O_3287,N_48099,N_49350);
nor UO_3288 (O_3288,N_49613,N_49660);
nor UO_3289 (O_3289,N_49612,N_49812);
xor UO_3290 (O_3290,N_49364,N_49523);
nand UO_3291 (O_3291,N_48134,N_48962);
nor UO_3292 (O_3292,N_48173,N_48059);
nor UO_3293 (O_3293,N_49413,N_49334);
nor UO_3294 (O_3294,N_48178,N_49958);
xor UO_3295 (O_3295,N_49192,N_49889);
or UO_3296 (O_3296,N_48343,N_48372);
or UO_3297 (O_3297,N_49311,N_48075);
or UO_3298 (O_3298,N_49014,N_48748);
xnor UO_3299 (O_3299,N_49595,N_48983);
and UO_3300 (O_3300,N_49966,N_49463);
xnor UO_3301 (O_3301,N_49275,N_49244);
xnor UO_3302 (O_3302,N_49118,N_49435);
xnor UO_3303 (O_3303,N_49525,N_48337);
nor UO_3304 (O_3304,N_48760,N_48652);
nor UO_3305 (O_3305,N_49764,N_49703);
xnor UO_3306 (O_3306,N_48558,N_49189);
xnor UO_3307 (O_3307,N_49974,N_48361);
xnor UO_3308 (O_3308,N_48488,N_48012);
nor UO_3309 (O_3309,N_48211,N_49279);
xor UO_3310 (O_3310,N_49284,N_49065);
nand UO_3311 (O_3311,N_49267,N_49009);
xnor UO_3312 (O_3312,N_48578,N_49428);
or UO_3313 (O_3313,N_49691,N_49062);
and UO_3314 (O_3314,N_49328,N_49735);
xnor UO_3315 (O_3315,N_49513,N_48605);
xnor UO_3316 (O_3316,N_49586,N_49136);
and UO_3317 (O_3317,N_48034,N_49767);
and UO_3318 (O_3318,N_48051,N_49969);
xor UO_3319 (O_3319,N_49648,N_48943);
nor UO_3320 (O_3320,N_48179,N_48608);
nor UO_3321 (O_3321,N_49834,N_48117);
nor UO_3322 (O_3322,N_49425,N_48801);
and UO_3323 (O_3323,N_49632,N_48125);
nand UO_3324 (O_3324,N_48481,N_49069);
nor UO_3325 (O_3325,N_49732,N_48638);
nand UO_3326 (O_3326,N_48084,N_48989);
nand UO_3327 (O_3327,N_49503,N_48917);
and UO_3328 (O_3328,N_48044,N_49875);
and UO_3329 (O_3329,N_48840,N_48416);
and UO_3330 (O_3330,N_49986,N_49503);
or UO_3331 (O_3331,N_48669,N_48244);
nand UO_3332 (O_3332,N_48590,N_49613);
nor UO_3333 (O_3333,N_49841,N_48117);
xor UO_3334 (O_3334,N_49063,N_48374);
or UO_3335 (O_3335,N_48176,N_49674);
or UO_3336 (O_3336,N_48659,N_48095);
or UO_3337 (O_3337,N_49376,N_48253);
nand UO_3338 (O_3338,N_49436,N_48488);
and UO_3339 (O_3339,N_48975,N_48109);
nand UO_3340 (O_3340,N_48936,N_49563);
nor UO_3341 (O_3341,N_48749,N_49042);
nand UO_3342 (O_3342,N_48489,N_48628);
and UO_3343 (O_3343,N_49655,N_49510);
and UO_3344 (O_3344,N_49543,N_48237);
nor UO_3345 (O_3345,N_49853,N_49964);
and UO_3346 (O_3346,N_49352,N_48677);
and UO_3347 (O_3347,N_49439,N_48538);
nor UO_3348 (O_3348,N_48487,N_49781);
xnor UO_3349 (O_3349,N_48690,N_48479);
or UO_3350 (O_3350,N_49266,N_48048);
or UO_3351 (O_3351,N_48302,N_49336);
nor UO_3352 (O_3352,N_48563,N_49112);
or UO_3353 (O_3353,N_49720,N_48600);
and UO_3354 (O_3354,N_49608,N_48866);
and UO_3355 (O_3355,N_48571,N_49139);
and UO_3356 (O_3356,N_48710,N_49601);
nand UO_3357 (O_3357,N_48320,N_49545);
or UO_3358 (O_3358,N_48833,N_48394);
and UO_3359 (O_3359,N_48000,N_48627);
nand UO_3360 (O_3360,N_49024,N_49825);
nor UO_3361 (O_3361,N_49222,N_49474);
and UO_3362 (O_3362,N_48346,N_48738);
nand UO_3363 (O_3363,N_48035,N_49800);
and UO_3364 (O_3364,N_48950,N_49050);
and UO_3365 (O_3365,N_49766,N_48058);
nor UO_3366 (O_3366,N_49516,N_49781);
nor UO_3367 (O_3367,N_48780,N_48695);
and UO_3368 (O_3368,N_49117,N_48196);
xor UO_3369 (O_3369,N_49209,N_48943);
nand UO_3370 (O_3370,N_48913,N_49253);
nor UO_3371 (O_3371,N_48253,N_49438);
xnor UO_3372 (O_3372,N_48544,N_49281);
xor UO_3373 (O_3373,N_49268,N_48764);
nand UO_3374 (O_3374,N_48047,N_49109);
xor UO_3375 (O_3375,N_48365,N_48802);
or UO_3376 (O_3376,N_48294,N_49921);
nor UO_3377 (O_3377,N_48581,N_48455);
nor UO_3378 (O_3378,N_48144,N_49848);
xor UO_3379 (O_3379,N_49617,N_49030);
or UO_3380 (O_3380,N_49140,N_48519);
nand UO_3381 (O_3381,N_49989,N_49237);
xor UO_3382 (O_3382,N_48087,N_48103);
and UO_3383 (O_3383,N_48919,N_48682);
nand UO_3384 (O_3384,N_48142,N_49513);
and UO_3385 (O_3385,N_49489,N_48096);
xnor UO_3386 (O_3386,N_49215,N_48319);
or UO_3387 (O_3387,N_49536,N_49605);
nand UO_3388 (O_3388,N_49555,N_49845);
and UO_3389 (O_3389,N_48948,N_49063);
nand UO_3390 (O_3390,N_48419,N_49442);
or UO_3391 (O_3391,N_48515,N_48601);
and UO_3392 (O_3392,N_49430,N_48225);
nor UO_3393 (O_3393,N_48754,N_48140);
xor UO_3394 (O_3394,N_48487,N_49515);
and UO_3395 (O_3395,N_49305,N_48956);
nand UO_3396 (O_3396,N_48381,N_48697);
nor UO_3397 (O_3397,N_48304,N_48358);
xnor UO_3398 (O_3398,N_49951,N_48516);
xor UO_3399 (O_3399,N_48135,N_49531);
or UO_3400 (O_3400,N_48563,N_49570);
or UO_3401 (O_3401,N_48409,N_49392);
or UO_3402 (O_3402,N_48973,N_49030);
nor UO_3403 (O_3403,N_48797,N_48940);
or UO_3404 (O_3404,N_48865,N_49007);
or UO_3405 (O_3405,N_49850,N_48834);
and UO_3406 (O_3406,N_49105,N_49290);
nand UO_3407 (O_3407,N_49068,N_49411);
xnor UO_3408 (O_3408,N_48545,N_48465);
nor UO_3409 (O_3409,N_49062,N_49152);
nand UO_3410 (O_3410,N_49113,N_49953);
nand UO_3411 (O_3411,N_49826,N_48307);
and UO_3412 (O_3412,N_49260,N_48981);
nand UO_3413 (O_3413,N_48845,N_49061);
nand UO_3414 (O_3414,N_49840,N_48175);
and UO_3415 (O_3415,N_49433,N_49623);
or UO_3416 (O_3416,N_49591,N_48123);
xnor UO_3417 (O_3417,N_48325,N_49692);
and UO_3418 (O_3418,N_49546,N_48320);
or UO_3419 (O_3419,N_49408,N_48995);
or UO_3420 (O_3420,N_48231,N_48817);
and UO_3421 (O_3421,N_49487,N_49683);
nor UO_3422 (O_3422,N_49654,N_48355);
and UO_3423 (O_3423,N_49874,N_48631);
or UO_3424 (O_3424,N_48626,N_48192);
or UO_3425 (O_3425,N_48975,N_49347);
xor UO_3426 (O_3426,N_49811,N_48073);
nand UO_3427 (O_3427,N_49064,N_48975);
or UO_3428 (O_3428,N_48058,N_48095);
xnor UO_3429 (O_3429,N_48276,N_49741);
and UO_3430 (O_3430,N_49483,N_48250);
and UO_3431 (O_3431,N_48252,N_48103);
xor UO_3432 (O_3432,N_49954,N_49370);
or UO_3433 (O_3433,N_48428,N_49768);
and UO_3434 (O_3434,N_49710,N_49852);
nor UO_3435 (O_3435,N_49627,N_48134);
nor UO_3436 (O_3436,N_48215,N_48058);
or UO_3437 (O_3437,N_48826,N_49884);
or UO_3438 (O_3438,N_48686,N_48706);
xnor UO_3439 (O_3439,N_49410,N_48057);
nand UO_3440 (O_3440,N_48535,N_48431);
xnor UO_3441 (O_3441,N_48610,N_48938);
nand UO_3442 (O_3442,N_49977,N_49292);
xnor UO_3443 (O_3443,N_48026,N_49848);
nand UO_3444 (O_3444,N_49518,N_48916);
xor UO_3445 (O_3445,N_48978,N_49636);
and UO_3446 (O_3446,N_49442,N_48300);
nand UO_3447 (O_3447,N_48426,N_48527);
and UO_3448 (O_3448,N_49783,N_48084);
xor UO_3449 (O_3449,N_48989,N_48701);
xor UO_3450 (O_3450,N_48781,N_48214);
nor UO_3451 (O_3451,N_48728,N_48758);
nand UO_3452 (O_3452,N_49356,N_48815);
xor UO_3453 (O_3453,N_49421,N_48244);
xnor UO_3454 (O_3454,N_48956,N_48037);
nor UO_3455 (O_3455,N_48897,N_49448);
nand UO_3456 (O_3456,N_48135,N_49132);
nor UO_3457 (O_3457,N_48830,N_48092);
nand UO_3458 (O_3458,N_48256,N_48478);
xnor UO_3459 (O_3459,N_48074,N_49441);
and UO_3460 (O_3460,N_48697,N_49655);
or UO_3461 (O_3461,N_48118,N_49335);
xor UO_3462 (O_3462,N_49174,N_49865);
or UO_3463 (O_3463,N_49547,N_48019);
xor UO_3464 (O_3464,N_48872,N_48010);
or UO_3465 (O_3465,N_48026,N_49740);
nor UO_3466 (O_3466,N_49914,N_49094);
xor UO_3467 (O_3467,N_49587,N_48540);
and UO_3468 (O_3468,N_49846,N_49088);
and UO_3469 (O_3469,N_48186,N_49881);
and UO_3470 (O_3470,N_49108,N_49340);
or UO_3471 (O_3471,N_49834,N_49599);
xnor UO_3472 (O_3472,N_48009,N_48571);
and UO_3473 (O_3473,N_49010,N_48335);
xnor UO_3474 (O_3474,N_48470,N_48418);
xnor UO_3475 (O_3475,N_49218,N_49413);
and UO_3476 (O_3476,N_49427,N_48527);
nor UO_3477 (O_3477,N_49138,N_48548);
nand UO_3478 (O_3478,N_48255,N_49219);
or UO_3479 (O_3479,N_49832,N_48079);
nand UO_3480 (O_3480,N_49871,N_48940);
nor UO_3481 (O_3481,N_49031,N_48176);
nand UO_3482 (O_3482,N_48821,N_49828);
nand UO_3483 (O_3483,N_49879,N_48112);
and UO_3484 (O_3484,N_48954,N_48036);
and UO_3485 (O_3485,N_48238,N_49314);
or UO_3486 (O_3486,N_49845,N_48953);
or UO_3487 (O_3487,N_48213,N_48240);
xnor UO_3488 (O_3488,N_48616,N_48181);
and UO_3489 (O_3489,N_49338,N_48444);
and UO_3490 (O_3490,N_48512,N_48701);
and UO_3491 (O_3491,N_48199,N_49154);
and UO_3492 (O_3492,N_48659,N_49237);
nand UO_3493 (O_3493,N_49478,N_49947);
and UO_3494 (O_3494,N_48573,N_49538);
or UO_3495 (O_3495,N_49791,N_48332);
or UO_3496 (O_3496,N_49295,N_49746);
nand UO_3497 (O_3497,N_49903,N_49012);
nor UO_3498 (O_3498,N_49295,N_49151);
xor UO_3499 (O_3499,N_49277,N_49422);
xnor UO_3500 (O_3500,N_49966,N_49246);
or UO_3501 (O_3501,N_48143,N_48600);
xor UO_3502 (O_3502,N_49070,N_49232);
and UO_3503 (O_3503,N_49118,N_49361);
and UO_3504 (O_3504,N_48517,N_49072);
nor UO_3505 (O_3505,N_49892,N_49046);
xnor UO_3506 (O_3506,N_48894,N_48178);
nand UO_3507 (O_3507,N_48731,N_48802);
nor UO_3508 (O_3508,N_48348,N_49193);
nand UO_3509 (O_3509,N_48889,N_49972);
xor UO_3510 (O_3510,N_48675,N_48993);
xor UO_3511 (O_3511,N_49924,N_48124);
and UO_3512 (O_3512,N_49920,N_49590);
xor UO_3513 (O_3513,N_48569,N_49469);
nand UO_3514 (O_3514,N_48115,N_48997);
or UO_3515 (O_3515,N_48553,N_49684);
and UO_3516 (O_3516,N_49814,N_48701);
xnor UO_3517 (O_3517,N_49311,N_48022);
xor UO_3518 (O_3518,N_48116,N_49454);
nand UO_3519 (O_3519,N_48076,N_48678);
and UO_3520 (O_3520,N_48940,N_49521);
nand UO_3521 (O_3521,N_49556,N_48713);
and UO_3522 (O_3522,N_49533,N_48026);
nand UO_3523 (O_3523,N_48251,N_48678);
nand UO_3524 (O_3524,N_49593,N_49212);
and UO_3525 (O_3525,N_49796,N_48228);
or UO_3526 (O_3526,N_49312,N_49777);
xnor UO_3527 (O_3527,N_49626,N_49941);
or UO_3528 (O_3528,N_49326,N_48440);
xor UO_3529 (O_3529,N_48443,N_48072);
or UO_3530 (O_3530,N_48130,N_49441);
or UO_3531 (O_3531,N_49245,N_49798);
or UO_3532 (O_3532,N_49412,N_49111);
or UO_3533 (O_3533,N_49314,N_49568);
nor UO_3534 (O_3534,N_49219,N_48674);
nand UO_3535 (O_3535,N_48807,N_49630);
nor UO_3536 (O_3536,N_49539,N_48293);
and UO_3537 (O_3537,N_49374,N_49657);
xnor UO_3538 (O_3538,N_48548,N_49060);
nor UO_3539 (O_3539,N_49466,N_48343);
xor UO_3540 (O_3540,N_48865,N_48219);
or UO_3541 (O_3541,N_49040,N_48919);
xor UO_3542 (O_3542,N_48284,N_48775);
and UO_3543 (O_3543,N_49919,N_49748);
or UO_3544 (O_3544,N_48510,N_49364);
or UO_3545 (O_3545,N_49675,N_49047);
nor UO_3546 (O_3546,N_48017,N_49467);
nand UO_3547 (O_3547,N_48200,N_48946);
or UO_3548 (O_3548,N_48251,N_48970);
xnor UO_3549 (O_3549,N_48172,N_49537);
xnor UO_3550 (O_3550,N_48410,N_48728);
nor UO_3551 (O_3551,N_48913,N_48763);
nand UO_3552 (O_3552,N_48453,N_49632);
nor UO_3553 (O_3553,N_48927,N_48699);
or UO_3554 (O_3554,N_49641,N_49305);
or UO_3555 (O_3555,N_48499,N_49491);
nor UO_3556 (O_3556,N_49038,N_48645);
xor UO_3557 (O_3557,N_49890,N_48023);
nor UO_3558 (O_3558,N_49481,N_48169);
nor UO_3559 (O_3559,N_48011,N_49227);
nor UO_3560 (O_3560,N_49335,N_49313);
and UO_3561 (O_3561,N_48041,N_49643);
or UO_3562 (O_3562,N_48414,N_48668);
and UO_3563 (O_3563,N_48766,N_49838);
xor UO_3564 (O_3564,N_49675,N_49684);
and UO_3565 (O_3565,N_48072,N_49740);
nand UO_3566 (O_3566,N_48396,N_49919);
nor UO_3567 (O_3567,N_48363,N_49852);
nor UO_3568 (O_3568,N_48536,N_49870);
xnor UO_3569 (O_3569,N_49520,N_48674);
nor UO_3570 (O_3570,N_48253,N_49944);
nand UO_3571 (O_3571,N_48016,N_49159);
nor UO_3572 (O_3572,N_49003,N_48757);
nor UO_3573 (O_3573,N_49699,N_49830);
nor UO_3574 (O_3574,N_49483,N_48112);
and UO_3575 (O_3575,N_48309,N_49698);
nor UO_3576 (O_3576,N_49701,N_49971);
nand UO_3577 (O_3577,N_49856,N_48736);
and UO_3578 (O_3578,N_48268,N_48392);
nand UO_3579 (O_3579,N_48012,N_48890);
and UO_3580 (O_3580,N_49727,N_49894);
nor UO_3581 (O_3581,N_49955,N_48689);
or UO_3582 (O_3582,N_49194,N_48722);
and UO_3583 (O_3583,N_48317,N_49744);
and UO_3584 (O_3584,N_49090,N_48771);
xor UO_3585 (O_3585,N_48235,N_49862);
and UO_3586 (O_3586,N_48470,N_48520);
xor UO_3587 (O_3587,N_48575,N_48991);
and UO_3588 (O_3588,N_49210,N_48232);
xor UO_3589 (O_3589,N_48041,N_48745);
nor UO_3590 (O_3590,N_49345,N_48063);
or UO_3591 (O_3591,N_48753,N_48734);
nand UO_3592 (O_3592,N_49814,N_48034);
xnor UO_3593 (O_3593,N_48880,N_49769);
nand UO_3594 (O_3594,N_49661,N_49903);
or UO_3595 (O_3595,N_48654,N_48073);
xnor UO_3596 (O_3596,N_49816,N_48029);
and UO_3597 (O_3597,N_49754,N_48141);
xor UO_3598 (O_3598,N_48171,N_48901);
nand UO_3599 (O_3599,N_49858,N_48382);
or UO_3600 (O_3600,N_49293,N_48367);
and UO_3601 (O_3601,N_48741,N_49832);
nand UO_3602 (O_3602,N_48940,N_48280);
nor UO_3603 (O_3603,N_48958,N_48987);
xnor UO_3604 (O_3604,N_49086,N_49868);
and UO_3605 (O_3605,N_48214,N_49901);
and UO_3606 (O_3606,N_48607,N_49239);
xor UO_3607 (O_3607,N_49575,N_49646);
or UO_3608 (O_3608,N_48589,N_49232);
xnor UO_3609 (O_3609,N_48647,N_49685);
xor UO_3610 (O_3610,N_48467,N_49778);
and UO_3611 (O_3611,N_48586,N_48567);
and UO_3612 (O_3612,N_48468,N_49196);
nor UO_3613 (O_3613,N_49357,N_48003);
and UO_3614 (O_3614,N_49851,N_49270);
or UO_3615 (O_3615,N_48753,N_49074);
nand UO_3616 (O_3616,N_48046,N_49717);
nor UO_3617 (O_3617,N_48983,N_48333);
or UO_3618 (O_3618,N_49975,N_49296);
nor UO_3619 (O_3619,N_48565,N_49088);
and UO_3620 (O_3620,N_48768,N_48004);
or UO_3621 (O_3621,N_49629,N_49259);
or UO_3622 (O_3622,N_49867,N_48468);
xnor UO_3623 (O_3623,N_49189,N_49223);
nand UO_3624 (O_3624,N_48453,N_49559);
and UO_3625 (O_3625,N_49586,N_49110);
or UO_3626 (O_3626,N_48712,N_48985);
nor UO_3627 (O_3627,N_48538,N_49742);
and UO_3628 (O_3628,N_49132,N_48601);
nand UO_3629 (O_3629,N_48271,N_48375);
nor UO_3630 (O_3630,N_48759,N_48470);
and UO_3631 (O_3631,N_49202,N_48093);
nand UO_3632 (O_3632,N_48614,N_49836);
and UO_3633 (O_3633,N_49424,N_48520);
nand UO_3634 (O_3634,N_48815,N_48466);
and UO_3635 (O_3635,N_49977,N_48246);
or UO_3636 (O_3636,N_48506,N_48105);
or UO_3637 (O_3637,N_48438,N_49467);
and UO_3638 (O_3638,N_48182,N_48535);
nor UO_3639 (O_3639,N_48395,N_48383);
nor UO_3640 (O_3640,N_49869,N_48475);
and UO_3641 (O_3641,N_49946,N_49509);
nor UO_3642 (O_3642,N_49253,N_49670);
or UO_3643 (O_3643,N_48455,N_48863);
nor UO_3644 (O_3644,N_48992,N_48699);
nor UO_3645 (O_3645,N_49738,N_49595);
or UO_3646 (O_3646,N_48332,N_48185);
or UO_3647 (O_3647,N_48306,N_49433);
and UO_3648 (O_3648,N_48163,N_48640);
nand UO_3649 (O_3649,N_49498,N_48598);
xor UO_3650 (O_3650,N_48349,N_49551);
nand UO_3651 (O_3651,N_49244,N_49957);
or UO_3652 (O_3652,N_49320,N_48716);
xnor UO_3653 (O_3653,N_49198,N_49948);
or UO_3654 (O_3654,N_48328,N_49829);
and UO_3655 (O_3655,N_48315,N_49230);
nand UO_3656 (O_3656,N_48673,N_48293);
and UO_3657 (O_3657,N_48410,N_49877);
nand UO_3658 (O_3658,N_49411,N_49203);
xnor UO_3659 (O_3659,N_49075,N_48426);
or UO_3660 (O_3660,N_48579,N_48324);
nor UO_3661 (O_3661,N_49670,N_49683);
nand UO_3662 (O_3662,N_49802,N_48325);
and UO_3663 (O_3663,N_48632,N_48595);
nor UO_3664 (O_3664,N_49952,N_48930);
or UO_3665 (O_3665,N_48933,N_49598);
or UO_3666 (O_3666,N_48176,N_48404);
and UO_3667 (O_3667,N_48584,N_49164);
and UO_3668 (O_3668,N_48169,N_49530);
nor UO_3669 (O_3669,N_49184,N_49009);
and UO_3670 (O_3670,N_48244,N_49815);
and UO_3671 (O_3671,N_48404,N_48424);
or UO_3672 (O_3672,N_48922,N_48952);
nand UO_3673 (O_3673,N_49368,N_48470);
and UO_3674 (O_3674,N_49042,N_49080);
nand UO_3675 (O_3675,N_49345,N_48402);
nor UO_3676 (O_3676,N_49765,N_48284);
or UO_3677 (O_3677,N_49137,N_48196);
xnor UO_3678 (O_3678,N_48868,N_49948);
nor UO_3679 (O_3679,N_49303,N_48725);
nor UO_3680 (O_3680,N_48480,N_48987);
or UO_3681 (O_3681,N_48105,N_49399);
nand UO_3682 (O_3682,N_49246,N_48448);
and UO_3683 (O_3683,N_48885,N_48439);
and UO_3684 (O_3684,N_49106,N_49960);
nor UO_3685 (O_3685,N_49956,N_49870);
nor UO_3686 (O_3686,N_48953,N_48128);
nand UO_3687 (O_3687,N_48748,N_48585);
nand UO_3688 (O_3688,N_49867,N_48565);
nand UO_3689 (O_3689,N_48591,N_48453);
nor UO_3690 (O_3690,N_48402,N_49498);
or UO_3691 (O_3691,N_48199,N_48261);
or UO_3692 (O_3692,N_49232,N_49694);
nand UO_3693 (O_3693,N_49432,N_48145);
nand UO_3694 (O_3694,N_48954,N_48238);
nand UO_3695 (O_3695,N_49324,N_48970);
and UO_3696 (O_3696,N_49619,N_48333);
nand UO_3697 (O_3697,N_48975,N_48307);
nor UO_3698 (O_3698,N_49076,N_49661);
xnor UO_3699 (O_3699,N_49117,N_48027);
nor UO_3700 (O_3700,N_48934,N_49941);
and UO_3701 (O_3701,N_49244,N_49061);
xnor UO_3702 (O_3702,N_48963,N_48993);
nand UO_3703 (O_3703,N_48326,N_48360);
xor UO_3704 (O_3704,N_48954,N_49657);
xor UO_3705 (O_3705,N_49959,N_49212);
nand UO_3706 (O_3706,N_49829,N_48339);
and UO_3707 (O_3707,N_49410,N_49014);
nand UO_3708 (O_3708,N_49719,N_48753);
nand UO_3709 (O_3709,N_49017,N_48608);
and UO_3710 (O_3710,N_49484,N_48598);
and UO_3711 (O_3711,N_48075,N_48687);
or UO_3712 (O_3712,N_49927,N_49206);
and UO_3713 (O_3713,N_48771,N_48697);
and UO_3714 (O_3714,N_48408,N_49360);
or UO_3715 (O_3715,N_48733,N_48150);
and UO_3716 (O_3716,N_49561,N_49095);
or UO_3717 (O_3717,N_49934,N_48384);
and UO_3718 (O_3718,N_48716,N_49095);
nor UO_3719 (O_3719,N_49664,N_49961);
and UO_3720 (O_3720,N_49154,N_48892);
xnor UO_3721 (O_3721,N_48460,N_49038);
nor UO_3722 (O_3722,N_49725,N_48179);
and UO_3723 (O_3723,N_48943,N_48331);
and UO_3724 (O_3724,N_49738,N_49641);
nor UO_3725 (O_3725,N_49308,N_49950);
xor UO_3726 (O_3726,N_48097,N_48328);
nand UO_3727 (O_3727,N_48893,N_49180);
xnor UO_3728 (O_3728,N_48065,N_48768);
nor UO_3729 (O_3729,N_49525,N_48577);
or UO_3730 (O_3730,N_48748,N_48089);
or UO_3731 (O_3731,N_49470,N_49061);
nand UO_3732 (O_3732,N_48690,N_48261);
and UO_3733 (O_3733,N_49638,N_48708);
nand UO_3734 (O_3734,N_48696,N_49650);
or UO_3735 (O_3735,N_49388,N_49250);
or UO_3736 (O_3736,N_48107,N_49672);
and UO_3737 (O_3737,N_48051,N_48694);
nor UO_3738 (O_3738,N_48481,N_49690);
or UO_3739 (O_3739,N_48149,N_48235);
or UO_3740 (O_3740,N_49847,N_48014);
or UO_3741 (O_3741,N_48646,N_49137);
nand UO_3742 (O_3742,N_48485,N_48058);
and UO_3743 (O_3743,N_49107,N_49083);
nand UO_3744 (O_3744,N_49759,N_49219);
xnor UO_3745 (O_3745,N_48283,N_48035);
xnor UO_3746 (O_3746,N_48210,N_49929);
or UO_3747 (O_3747,N_49684,N_48309);
nand UO_3748 (O_3748,N_48499,N_49490);
xor UO_3749 (O_3749,N_48555,N_49243);
and UO_3750 (O_3750,N_48290,N_48406);
xor UO_3751 (O_3751,N_48259,N_48192);
or UO_3752 (O_3752,N_49239,N_48463);
nand UO_3753 (O_3753,N_49470,N_49576);
xor UO_3754 (O_3754,N_48280,N_48791);
xor UO_3755 (O_3755,N_49847,N_49480);
nand UO_3756 (O_3756,N_48608,N_49514);
xor UO_3757 (O_3757,N_48477,N_48189);
nor UO_3758 (O_3758,N_48456,N_48536);
and UO_3759 (O_3759,N_48394,N_48085);
nor UO_3760 (O_3760,N_49330,N_49411);
xnor UO_3761 (O_3761,N_48608,N_49235);
or UO_3762 (O_3762,N_49240,N_49417);
nand UO_3763 (O_3763,N_49729,N_49552);
and UO_3764 (O_3764,N_49864,N_48622);
nand UO_3765 (O_3765,N_48367,N_49695);
xor UO_3766 (O_3766,N_48033,N_48453);
or UO_3767 (O_3767,N_49707,N_49925);
or UO_3768 (O_3768,N_49010,N_48100);
and UO_3769 (O_3769,N_49364,N_48683);
or UO_3770 (O_3770,N_49225,N_48683);
or UO_3771 (O_3771,N_48110,N_49705);
xor UO_3772 (O_3772,N_49651,N_49739);
xor UO_3773 (O_3773,N_48492,N_48977);
nor UO_3774 (O_3774,N_48016,N_48945);
and UO_3775 (O_3775,N_48176,N_49171);
nor UO_3776 (O_3776,N_48693,N_49580);
and UO_3777 (O_3777,N_48468,N_49549);
and UO_3778 (O_3778,N_49474,N_48449);
nand UO_3779 (O_3779,N_49690,N_49330);
and UO_3780 (O_3780,N_49908,N_48062);
nor UO_3781 (O_3781,N_49813,N_49953);
nor UO_3782 (O_3782,N_49601,N_49759);
nand UO_3783 (O_3783,N_48735,N_49311);
and UO_3784 (O_3784,N_48341,N_49732);
and UO_3785 (O_3785,N_48033,N_49108);
nor UO_3786 (O_3786,N_48153,N_48331);
and UO_3787 (O_3787,N_48411,N_48555);
nor UO_3788 (O_3788,N_48295,N_48590);
or UO_3789 (O_3789,N_48942,N_49857);
and UO_3790 (O_3790,N_48985,N_49493);
and UO_3791 (O_3791,N_49076,N_48605);
nand UO_3792 (O_3792,N_48877,N_49330);
or UO_3793 (O_3793,N_49004,N_48957);
nand UO_3794 (O_3794,N_48710,N_48761);
nand UO_3795 (O_3795,N_48179,N_48708);
nand UO_3796 (O_3796,N_49663,N_49730);
nand UO_3797 (O_3797,N_49770,N_48283);
or UO_3798 (O_3798,N_48196,N_49943);
nor UO_3799 (O_3799,N_49458,N_49892);
nand UO_3800 (O_3800,N_48358,N_48686);
or UO_3801 (O_3801,N_49823,N_49727);
or UO_3802 (O_3802,N_49981,N_48797);
xor UO_3803 (O_3803,N_48762,N_49293);
nor UO_3804 (O_3804,N_49936,N_48069);
and UO_3805 (O_3805,N_48640,N_48121);
xor UO_3806 (O_3806,N_49829,N_48401);
nor UO_3807 (O_3807,N_49766,N_48428);
xor UO_3808 (O_3808,N_49174,N_48435);
nand UO_3809 (O_3809,N_49276,N_48469);
nand UO_3810 (O_3810,N_49470,N_49689);
and UO_3811 (O_3811,N_48097,N_48933);
or UO_3812 (O_3812,N_49296,N_49275);
nand UO_3813 (O_3813,N_49420,N_48363);
or UO_3814 (O_3814,N_48187,N_48052);
or UO_3815 (O_3815,N_49484,N_48261);
nand UO_3816 (O_3816,N_48404,N_49653);
xnor UO_3817 (O_3817,N_48516,N_49814);
xor UO_3818 (O_3818,N_49945,N_48322);
xnor UO_3819 (O_3819,N_48432,N_48441);
or UO_3820 (O_3820,N_48004,N_49294);
and UO_3821 (O_3821,N_49192,N_48380);
or UO_3822 (O_3822,N_48200,N_49002);
nand UO_3823 (O_3823,N_48985,N_48731);
xnor UO_3824 (O_3824,N_48213,N_49395);
and UO_3825 (O_3825,N_49134,N_49398);
nor UO_3826 (O_3826,N_48109,N_49634);
xnor UO_3827 (O_3827,N_48827,N_48987);
or UO_3828 (O_3828,N_48988,N_49036);
or UO_3829 (O_3829,N_48608,N_48084);
nand UO_3830 (O_3830,N_48638,N_48235);
xor UO_3831 (O_3831,N_49851,N_49212);
nand UO_3832 (O_3832,N_48641,N_48311);
nor UO_3833 (O_3833,N_48479,N_48688);
or UO_3834 (O_3834,N_49701,N_49757);
and UO_3835 (O_3835,N_48477,N_49105);
nand UO_3836 (O_3836,N_48594,N_49778);
nor UO_3837 (O_3837,N_48582,N_49794);
and UO_3838 (O_3838,N_48022,N_49453);
or UO_3839 (O_3839,N_49127,N_49213);
or UO_3840 (O_3840,N_49877,N_48652);
nand UO_3841 (O_3841,N_48637,N_49340);
nor UO_3842 (O_3842,N_49227,N_48796);
nand UO_3843 (O_3843,N_49931,N_48669);
xor UO_3844 (O_3844,N_48202,N_49936);
xor UO_3845 (O_3845,N_48324,N_49738);
and UO_3846 (O_3846,N_48314,N_48696);
nand UO_3847 (O_3847,N_49369,N_49722);
or UO_3848 (O_3848,N_48964,N_48562);
and UO_3849 (O_3849,N_49499,N_49338);
nor UO_3850 (O_3850,N_48123,N_49826);
and UO_3851 (O_3851,N_49763,N_49163);
and UO_3852 (O_3852,N_49903,N_48639);
and UO_3853 (O_3853,N_49627,N_48752);
xor UO_3854 (O_3854,N_49070,N_48659);
nand UO_3855 (O_3855,N_48975,N_49273);
or UO_3856 (O_3856,N_49487,N_49883);
xnor UO_3857 (O_3857,N_48777,N_48072);
xnor UO_3858 (O_3858,N_48559,N_48552);
xor UO_3859 (O_3859,N_49634,N_48366);
xor UO_3860 (O_3860,N_49970,N_48695);
nor UO_3861 (O_3861,N_48606,N_49710);
xor UO_3862 (O_3862,N_48730,N_49823);
nand UO_3863 (O_3863,N_48363,N_48422);
or UO_3864 (O_3864,N_48816,N_49344);
nand UO_3865 (O_3865,N_49991,N_49120);
and UO_3866 (O_3866,N_48625,N_49695);
nor UO_3867 (O_3867,N_49763,N_48887);
nor UO_3868 (O_3868,N_48014,N_48302);
nand UO_3869 (O_3869,N_48041,N_48926);
nand UO_3870 (O_3870,N_49358,N_48780);
xor UO_3871 (O_3871,N_49352,N_48386);
nand UO_3872 (O_3872,N_49209,N_49695);
xnor UO_3873 (O_3873,N_48282,N_48939);
xor UO_3874 (O_3874,N_48691,N_48978);
nor UO_3875 (O_3875,N_49350,N_49329);
nand UO_3876 (O_3876,N_49245,N_49081);
xor UO_3877 (O_3877,N_48534,N_49160);
and UO_3878 (O_3878,N_49924,N_48720);
or UO_3879 (O_3879,N_49018,N_49471);
or UO_3880 (O_3880,N_48726,N_48040);
nor UO_3881 (O_3881,N_49214,N_48432);
nand UO_3882 (O_3882,N_48467,N_49457);
and UO_3883 (O_3883,N_48685,N_49091);
and UO_3884 (O_3884,N_48264,N_48185);
and UO_3885 (O_3885,N_49019,N_49098);
xor UO_3886 (O_3886,N_48433,N_49410);
and UO_3887 (O_3887,N_49922,N_48786);
or UO_3888 (O_3888,N_48309,N_49562);
nor UO_3889 (O_3889,N_48084,N_49739);
nor UO_3890 (O_3890,N_49495,N_48874);
or UO_3891 (O_3891,N_48493,N_48953);
nor UO_3892 (O_3892,N_48638,N_48788);
xor UO_3893 (O_3893,N_49251,N_48096);
nand UO_3894 (O_3894,N_49042,N_48922);
nor UO_3895 (O_3895,N_48286,N_49158);
xnor UO_3896 (O_3896,N_48748,N_48816);
nand UO_3897 (O_3897,N_49454,N_48026);
nor UO_3898 (O_3898,N_49540,N_48525);
nand UO_3899 (O_3899,N_49318,N_48309);
and UO_3900 (O_3900,N_48148,N_49434);
or UO_3901 (O_3901,N_49716,N_49825);
and UO_3902 (O_3902,N_49026,N_49744);
or UO_3903 (O_3903,N_49659,N_49571);
or UO_3904 (O_3904,N_49924,N_48882);
xnor UO_3905 (O_3905,N_49096,N_49822);
nor UO_3906 (O_3906,N_49874,N_49572);
xor UO_3907 (O_3907,N_49467,N_48358);
xnor UO_3908 (O_3908,N_48655,N_48488);
and UO_3909 (O_3909,N_49992,N_48538);
and UO_3910 (O_3910,N_48315,N_49969);
xnor UO_3911 (O_3911,N_48223,N_49050);
nor UO_3912 (O_3912,N_48830,N_48332);
nor UO_3913 (O_3913,N_48698,N_48759);
xnor UO_3914 (O_3914,N_48469,N_49949);
xor UO_3915 (O_3915,N_49928,N_48100);
or UO_3916 (O_3916,N_49325,N_48135);
and UO_3917 (O_3917,N_49029,N_48532);
and UO_3918 (O_3918,N_49478,N_48056);
or UO_3919 (O_3919,N_48209,N_49331);
and UO_3920 (O_3920,N_49849,N_48241);
nor UO_3921 (O_3921,N_49475,N_48379);
nor UO_3922 (O_3922,N_49470,N_48926);
xor UO_3923 (O_3923,N_49367,N_49509);
nor UO_3924 (O_3924,N_49725,N_48890);
xnor UO_3925 (O_3925,N_49932,N_48237);
nor UO_3926 (O_3926,N_48214,N_48040);
nor UO_3927 (O_3927,N_48849,N_48794);
xor UO_3928 (O_3928,N_48001,N_48361);
and UO_3929 (O_3929,N_49403,N_49057);
and UO_3930 (O_3930,N_48088,N_48599);
or UO_3931 (O_3931,N_48699,N_49446);
and UO_3932 (O_3932,N_48657,N_48615);
and UO_3933 (O_3933,N_48933,N_49518);
nand UO_3934 (O_3934,N_48564,N_48775);
xor UO_3935 (O_3935,N_48928,N_48471);
nor UO_3936 (O_3936,N_48516,N_49756);
xnor UO_3937 (O_3937,N_49249,N_48260);
nand UO_3938 (O_3938,N_49049,N_48155);
nand UO_3939 (O_3939,N_48485,N_48256);
xnor UO_3940 (O_3940,N_49524,N_48858);
xor UO_3941 (O_3941,N_49466,N_48567);
nand UO_3942 (O_3942,N_49416,N_49467);
nor UO_3943 (O_3943,N_49788,N_49023);
or UO_3944 (O_3944,N_49004,N_48640);
and UO_3945 (O_3945,N_49979,N_48978);
xor UO_3946 (O_3946,N_49941,N_48609);
and UO_3947 (O_3947,N_48021,N_48870);
nand UO_3948 (O_3948,N_49387,N_49772);
nor UO_3949 (O_3949,N_49520,N_48375);
nand UO_3950 (O_3950,N_48427,N_49317);
nor UO_3951 (O_3951,N_48370,N_48889);
or UO_3952 (O_3952,N_49713,N_48175);
xor UO_3953 (O_3953,N_48174,N_49636);
xor UO_3954 (O_3954,N_48836,N_49652);
nand UO_3955 (O_3955,N_49884,N_49890);
or UO_3956 (O_3956,N_48207,N_49451);
xnor UO_3957 (O_3957,N_49795,N_49205);
nand UO_3958 (O_3958,N_49153,N_49155);
nand UO_3959 (O_3959,N_48375,N_48580);
nand UO_3960 (O_3960,N_49515,N_48843);
or UO_3961 (O_3961,N_49891,N_49844);
nor UO_3962 (O_3962,N_49980,N_48329);
nor UO_3963 (O_3963,N_49443,N_49555);
nand UO_3964 (O_3964,N_49677,N_49324);
nor UO_3965 (O_3965,N_49761,N_48939);
or UO_3966 (O_3966,N_48275,N_49022);
xnor UO_3967 (O_3967,N_49700,N_48910);
nand UO_3968 (O_3968,N_48548,N_49746);
nand UO_3969 (O_3969,N_49042,N_48933);
nor UO_3970 (O_3970,N_48153,N_49600);
nand UO_3971 (O_3971,N_49758,N_49479);
or UO_3972 (O_3972,N_49983,N_49692);
nor UO_3973 (O_3973,N_48768,N_49491);
nor UO_3974 (O_3974,N_48657,N_48640);
and UO_3975 (O_3975,N_48652,N_49671);
and UO_3976 (O_3976,N_49280,N_49915);
xor UO_3977 (O_3977,N_49192,N_48511);
nand UO_3978 (O_3978,N_49723,N_48739);
xor UO_3979 (O_3979,N_48624,N_48363);
nand UO_3980 (O_3980,N_48756,N_49551);
and UO_3981 (O_3981,N_48539,N_48392);
and UO_3982 (O_3982,N_48467,N_49914);
xor UO_3983 (O_3983,N_49618,N_48341);
nor UO_3984 (O_3984,N_48608,N_48996);
and UO_3985 (O_3985,N_49320,N_49339);
or UO_3986 (O_3986,N_49621,N_49560);
nor UO_3987 (O_3987,N_49945,N_48729);
and UO_3988 (O_3988,N_49913,N_49626);
xor UO_3989 (O_3989,N_48988,N_49894);
nor UO_3990 (O_3990,N_48792,N_48418);
xor UO_3991 (O_3991,N_48616,N_48852);
or UO_3992 (O_3992,N_48172,N_48047);
nor UO_3993 (O_3993,N_48938,N_49674);
nor UO_3994 (O_3994,N_49891,N_48919);
and UO_3995 (O_3995,N_48529,N_48037);
or UO_3996 (O_3996,N_49214,N_49064);
or UO_3997 (O_3997,N_48032,N_48342);
xnor UO_3998 (O_3998,N_49719,N_48128);
nor UO_3999 (O_3999,N_48431,N_49914);
or UO_4000 (O_4000,N_48552,N_48583);
nor UO_4001 (O_4001,N_49325,N_49436);
nor UO_4002 (O_4002,N_49989,N_48586);
xor UO_4003 (O_4003,N_48812,N_48513);
xor UO_4004 (O_4004,N_49933,N_48595);
nand UO_4005 (O_4005,N_48802,N_49097);
nor UO_4006 (O_4006,N_48553,N_48771);
nor UO_4007 (O_4007,N_49073,N_49022);
nand UO_4008 (O_4008,N_49406,N_49555);
and UO_4009 (O_4009,N_49847,N_48510);
xor UO_4010 (O_4010,N_48083,N_49787);
or UO_4011 (O_4011,N_48266,N_49918);
and UO_4012 (O_4012,N_49254,N_49586);
nor UO_4013 (O_4013,N_48191,N_48546);
nor UO_4014 (O_4014,N_48567,N_48848);
xnor UO_4015 (O_4015,N_49014,N_49717);
xor UO_4016 (O_4016,N_48931,N_48585);
or UO_4017 (O_4017,N_49118,N_49505);
and UO_4018 (O_4018,N_48268,N_49272);
nand UO_4019 (O_4019,N_49223,N_48891);
nand UO_4020 (O_4020,N_48179,N_49583);
xnor UO_4021 (O_4021,N_49561,N_48147);
nand UO_4022 (O_4022,N_48237,N_48234);
and UO_4023 (O_4023,N_48565,N_49611);
or UO_4024 (O_4024,N_48109,N_48987);
nand UO_4025 (O_4025,N_49120,N_48776);
nor UO_4026 (O_4026,N_49068,N_48476);
and UO_4027 (O_4027,N_48690,N_49069);
xor UO_4028 (O_4028,N_48343,N_48559);
and UO_4029 (O_4029,N_48063,N_49014);
and UO_4030 (O_4030,N_49880,N_48021);
nor UO_4031 (O_4031,N_48286,N_49312);
xnor UO_4032 (O_4032,N_48310,N_48431);
and UO_4033 (O_4033,N_49835,N_48038);
nor UO_4034 (O_4034,N_48695,N_49064);
nor UO_4035 (O_4035,N_48839,N_48751);
or UO_4036 (O_4036,N_49688,N_48168);
and UO_4037 (O_4037,N_49698,N_48379);
nand UO_4038 (O_4038,N_49700,N_48083);
and UO_4039 (O_4039,N_49058,N_48688);
and UO_4040 (O_4040,N_49732,N_48721);
nand UO_4041 (O_4041,N_49611,N_48388);
or UO_4042 (O_4042,N_48396,N_48277);
or UO_4043 (O_4043,N_49148,N_49327);
and UO_4044 (O_4044,N_48300,N_48542);
nand UO_4045 (O_4045,N_48968,N_49520);
nand UO_4046 (O_4046,N_48394,N_48988);
nand UO_4047 (O_4047,N_49812,N_49622);
nand UO_4048 (O_4048,N_49837,N_48321);
nor UO_4049 (O_4049,N_49900,N_49329);
and UO_4050 (O_4050,N_49800,N_49339);
nor UO_4051 (O_4051,N_48334,N_49199);
and UO_4052 (O_4052,N_49498,N_48411);
or UO_4053 (O_4053,N_48553,N_49374);
or UO_4054 (O_4054,N_48517,N_49088);
and UO_4055 (O_4055,N_48890,N_48796);
nor UO_4056 (O_4056,N_48093,N_49265);
and UO_4057 (O_4057,N_49001,N_49334);
nand UO_4058 (O_4058,N_48193,N_48305);
xnor UO_4059 (O_4059,N_49073,N_49665);
nor UO_4060 (O_4060,N_49330,N_48810);
and UO_4061 (O_4061,N_49085,N_48729);
nand UO_4062 (O_4062,N_48809,N_48768);
and UO_4063 (O_4063,N_49106,N_49664);
and UO_4064 (O_4064,N_48220,N_49542);
and UO_4065 (O_4065,N_49050,N_48622);
nand UO_4066 (O_4066,N_48984,N_48725);
xor UO_4067 (O_4067,N_48285,N_48356);
nor UO_4068 (O_4068,N_48326,N_49313);
and UO_4069 (O_4069,N_49765,N_48649);
xor UO_4070 (O_4070,N_48849,N_48236);
and UO_4071 (O_4071,N_49207,N_48456);
xnor UO_4072 (O_4072,N_49570,N_48430);
xnor UO_4073 (O_4073,N_48155,N_49580);
nand UO_4074 (O_4074,N_48458,N_49780);
xor UO_4075 (O_4075,N_49772,N_48080);
nand UO_4076 (O_4076,N_49422,N_48444);
nor UO_4077 (O_4077,N_48055,N_48448);
or UO_4078 (O_4078,N_48711,N_48473);
nand UO_4079 (O_4079,N_48862,N_48761);
nor UO_4080 (O_4080,N_49214,N_48158);
or UO_4081 (O_4081,N_48595,N_49552);
or UO_4082 (O_4082,N_49590,N_48914);
nand UO_4083 (O_4083,N_49373,N_49073);
nor UO_4084 (O_4084,N_49177,N_49547);
xnor UO_4085 (O_4085,N_48124,N_49972);
xnor UO_4086 (O_4086,N_48151,N_48761);
xor UO_4087 (O_4087,N_49008,N_48668);
and UO_4088 (O_4088,N_49581,N_48194);
or UO_4089 (O_4089,N_49541,N_49677);
and UO_4090 (O_4090,N_48623,N_48709);
nand UO_4091 (O_4091,N_48647,N_49842);
or UO_4092 (O_4092,N_48656,N_49610);
nand UO_4093 (O_4093,N_49921,N_49077);
or UO_4094 (O_4094,N_48230,N_49113);
xor UO_4095 (O_4095,N_48607,N_49612);
xnor UO_4096 (O_4096,N_48648,N_48109);
nor UO_4097 (O_4097,N_48495,N_48477);
and UO_4098 (O_4098,N_48378,N_48022);
or UO_4099 (O_4099,N_48699,N_49979);
or UO_4100 (O_4100,N_49972,N_49306);
xor UO_4101 (O_4101,N_48302,N_49209);
nand UO_4102 (O_4102,N_49344,N_49275);
and UO_4103 (O_4103,N_49006,N_48979);
or UO_4104 (O_4104,N_48680,N_48021);
nor UO_4105 (O_4105,N_49833,N_49241);
xor UO_4106 (O_4106,N_48687,N_49284);
or UO_4107 (O_4107,N_48111,N_48421);
xor UO_4108 (O_4108,N_48671,N_48742);
or UO_4109 (O_4109,N_49821,N_48463);
or UO_4110 (O_4110,N_48537,N_49251);
or UO_4111 (O_4111,N_48481,N_49867);
nand UO_4112 (O_4112,N_48016,N_48959);
and UO_4113 (O_4113,N_49426,N_48664);
xor UO_4114 (O_4114,N_48969,N_48442);
or UO_4115 (O_4115,N_49247,N_49946);
nand UO_4116 (O_4116,N_48262,N_48258);
and UO_4117 (O_4117,N_49832,N_48534);
or UO_4118 (O_4118,N_49291,N_48849);
and UO_4119 (O_4119,N_49151,N_49222);
nor UO_4120 (O_4120,N_49535,N_49813);
nor UO_4121 (O_4121,N_49421,N_49213);
nand UO_4122 (O_4122,N_48102,N_49557);
nor UO_4123 (O_4123,N_48221,N_48542);
or UO_4124 (O_4124,N_48193,N_48464);
and UO_4125 (O_4125,N_48892,N_48564);
or UO_4126 (O_4126,N_48387,N_48829);
nor UO_4127 (O_4127,N_48443,N_48788);
nor UO_4128 (O_4128,N_49855,N_48405);
xnor UO_4129 (O_4129,N_49977,N_49648);
or UO_4130 (O_4130,N_48700,N_49656);
nor UO_4131 (O_4131,N_48666,N_48846);
nor UO_4132 (O_4132,N_48206,N_49881);
xor UO_4133 (O_4133,N_49225,N_49437);
nor UO_4134 (O_4134,N_48926,N_49246);
or UO_4135 (O_4135,N_48232,N_48674);
or UO_4136 (O_4136,N_48640,N_49934);
or UO_4137 (O_4137,N_48646,N_49899);
xnor UO_4138 (O_4138,N_48169,N_48231);
nor UO_4139 (O_4139,N_48127,N_48037);
nand UO_4140 (O_4140,N_49940,N_48132);
nor UO_4141 (O_4141,N_49369,N_48965);
nand UO_4142 (O_4142,N_48454,N_48601);
nand UO_4143 (O_4143,N_49571,N_49901);
xnor UO_4144 (O_4144,N_48790,N_48547);
nand UO_4145 (O_4145,N_48650,N_48595);
or UO_4146 (O_4146,N_49880,N_48252);
or UO_4147 (O_4147,N_49916,N_48343);
and UO_4148 (O_4148,N_48729,N_48525);
and UO_4149 (O_4149,N_49104,N_48779);
and UO_4150 (O_4150,N_49765,N_49871);
xor UO_4151 (O_4151,N_49382,N_49439);
nor UO_4152 (O_4152,N_49855,N_49971);
and UO_4153 (O_4153,N_49353,N_49970);
and UO_4154 (O_4154,N_48091,N_48171);
and UO_4155 (O_4155,N_49919,N_49960);
nand UO_4156 (O_4156,N_49332,N_48502);
or UO_4157 (O_4157,N_49318,N_48678);
nand UO_4158 (O_4158,N_49705,N_49407);
xor UO_4159 (O_4159,N_48901,N_48942);
nor UO_4160 (O_4160,N_49785,N_48135);
nor UO_4161 (O_4161,N_49671,N_49842);
or UO_4162 (O_4162,N_49633,N_49330);
or UO_4163 (O_4163,N_49785,N_49640);
xnor UO_4164 (O_4164,N_49159,N_49152);
and UO_4165 (O_4165,N_48944,N_49751);
nor UO_4166 (O_4166,N_48870,N_49708);
and UO_4167 (O_4167,N_49625,N_48308);
nor UO_4168 (O_4168,N_49467,N_49423);
nor UO_4169 (O_4169,N_48142,N_48300);
or UO_4170 (O_4170,N_48563,N_48936);
nand UO_4171 (O_4171,N_48016,N_48048);
nand UO_4172 (O_4172,N_49495,N_49532);
or UO_4173 (O_4173,N_49323,N_49256);
nor UO_4174 (O_4174,N_49713,N_49487);
xor UO_4175 (O_4175,N_48791,N_48815);
or UO_4176 (O_4176,N_49066,N_48573);
and UO_4177 (O_4177,N_49096,N_49659);
xnor UO_4178 (O_4178,N_49948,N_49733);
or UO_4179 (O_4179,N_48873,N_48671);
nor UO_4180 (O_4180,N_48236,N_49265);
nand UO_4181 (O_4181,N_48578,N_48860);
xnor UO_4182 (O_4182,N_48840,N_49313);
and UO_4183 (O_4183,N_48234,N_48897);
or UO_4184 (O_4184,N_49502,N_49728);
nor UO_4185 (O_4185,N_48849,N_48603);
xnor UO_4186 (O_4186,N_48056,N_49818);
xor UO_4187 (O_4187,N_48521,N_49338);
nand UO_4188 (O_4188,N_49058,N_49549);
xnor UO_4189 (O_4189,N_49215,N_48790);
or UO_4190 (O_4190,N_49692,N_49764);
and UO_4191 (O_4191,N_48055,N_49486);
or UO_4192 (O_4192,N_49023,N_49035);
nor UO_4193 (O_4193,N_48205,N_48309);
nor UO_4194 (O_4194,N_49215,N_48753);
xor UO_4195 (O_4195,N_49093,N_49675);
and UO_4196 (O_4196,N_49994,N_49538);
and UO_4197 (O_4197,N_48198,N_48976);
xor UO_4198 (O_4198,N_48844,N_48885);
xor UO_4199 (O_4199,N_49907,N_49767);
and UO_4200 (O_4200,N_49826,N_48950);
and UO_4201 (O_4201,N_49286,N_49555);
nand UO_4202 (O_4202,N_48388,N_49969);
xnor UO_4203 (O_4203,N_48684,N_48923);
xnor UO_4204 (O_4204,N_48819,N_49722);
and UO_4205 (O_4205,N_48979,N_49025);
nand UO_4206 (O_4206,N_48826,N_48278);
or UO_4207 (O_4207,N_49840,N_48960);
or UO_4208 (O_4208,N_49030,N_48540);
xor UO_4209 (O_4209,N_48697,N_49496);
and UO_4210 (O_4210,N_49762,N_49592);
xnor UO_4211 (O_4211,N_49089,N_49878);
and UO_4212 (O_4212,N_48066,N_49235);
xor UO_4213 (O_4213,N_48892,N_49570);
and UO_4214 (O_4214,N_48213,N_49216);
and UO_4215 (O_4215,N_49792,N_48829);
nor UO_4216 (O_4216,N_49084,N_49703);
xor UO_4217 (O_4217,N_49739,N_49948);
nand UO_4218 (O_4218,N_49241,N_49484);
nand UO_4219 (O_4219,N_48084,N_49779);
and UO_4220 (O_4220,N_48455,N_48127);
nor UO_4221 (O_4221,N_48795,N_49971);
or UO_4222 (O_4222,N_49587,N_48767);
or UO_4223 (O_4223,N_48574,N_48668);
and UO_4224 (O_4224,N_48268,N_49081);
or UO_4225 (O_4225,N_48230,N_48280);
xnor UO_4226 (O_4226,N_49361,N_48594);
nand UO_4227 (O_4227,N_48242,N_49376);
xor UO_4228 (O_4228,N_49402,N_49799);
or UO_4229 (O_4229,N_49421,N_48673);
nor UO_4230 (O_4230,N_49824,N_49975);
nand UO_4231 (O_4231,N_48539,N_48042);
and UO_4232 (O_4232,N_48835,N_48811);
xor UO_4233 (O_4233,N_48465,N_48041);
nor UO_4234 (O_4234,N_48491,N_49202);
nand UO_4235 (O_4235,N_48461,N_49003);
nand UO_4236 (O_4236,N_48165,N_48961);
and UO_4237 (O_4237,N_48296,N_48836);
nor UO_4238 (O_4238,N_48805,N_48123);
and UO_4239 (O_4239,N_49534,N_49161);
and UO_4240 (O_4240,N_48349,N_48115);
nor UO_4241 (O_4241,N_49645,N_49200);
nand UO_4242 (O_4242,N_49614,N_48282);
and UO_4243 (O_4243,N_49292,N_48699);
or UO_4244 (O_4244,N_48922,N_49366);
xnor UO_4245 (O_4245,N_48714,N_49738);
or UO_4246 (O_4246,N_49818,N_48253);
and UO_4247 (O_4247,N_49619,N_48617);
xor UO_4248 (O_4248,N_49611,N_49170);
nand UO_4249 (O_4249,N_48404,N_49858);
xnor UO_4250 (O_4250,N_48202,N_48878);
or UO_4251 (O_4251,N_49581,N_49257);
nand UO_4252 (O_4252,N_48994,N_49791);
nor UO_4253 (O_4253,N_48886,N_49028);
or UO_4254 (O_4254,N_49197,N_48867);
nor UO_4255 (O_4255,N_48507,N_49083);
and UO_4256 (O_4256,N_48635,N_48201);
xor UO_4257 (O_4257,N_49501,N_48831);
xor UO_4258 (O_4258,N_49741,N_49165);
or UO_4259 (O_4259,N_49061,N_48188);
nand UO_4260 (O_4260,N_49361,N_48562);
xnor UO_4261 (O_4261,N_48733,N_48111);
and UO_4262 (O_4262,N_49725,N_49651);
and UO_4263 (O_4263,N_49810,N_49291);
nand UO_4264 (O_4264,N_49340,N_48894);
nand UO_4265 (O_4265,N_48222,N_48999);
and UO_4266 (O_4266,N_49394,N_49623);
xor UO_4267 (O_4267,N_49857,N_48281);
or UO_4268 (O_4268,N_48010,N_48751);
nand UO_4269 (O_4269,N_48244,N_48005);
nor UO_4270 (O_4270,N_48299,N_48860);
nand UO_4271 (O_4271,N_48941,N_48371);
xnor UO_4272 (O_4272,N_48366,N_48316);
xor UO_4273 (O_4273,N_49344,N_48033);
xor UO_4274 (O_4274,N_48572,N_48446);
xnor UO_4275 (O_4275,N_48462,N_49136);
xnor UO_4276 (O_4276,N_48322,N_48605);
xnor UO_4277 (O_4277,N_49135,N_49324);
nand UO_4278 (O_4278,N_49296,N_48793);
nand UO_4279 (O_4279,N_49756,N_48182);
xor UO_4280 (O_4280,N_49330,N_48601);
nand UO_4281 (O_4281,N_49864,N_48159);
or UO_4282 (O_4282,N_49672,N_48641);
and UO_4283 (O_4283,N_49266,N_48445);
xor UO_4284 (O_4284,N_49966,N_49846);
xor UO_4285 (O_4285,N_48895,N_49226);
and UO_4286 (O_4286,N_49130,N_48221);
nand UO_4287 (O_4287,N_49857,N_48160);
nor UO_4288 (O_4288,N_49363,N_48904);
nor UO_4289 (O_4289,N_48940,N_48781);
nor UO_4290 (O_4290,N_48224,N_49361);
nor UO_4291 (O_4291,N_48574,N_49163);
nand UO_4292 (O_4292,N_49128,N_48157);
and UO_4293 (O_4293,N_48526,N_49220);
nor UO_4294 (O_4294,N_48682,N_49880);
nor UO_4295 (O_4295,N_49697,N_49255);
nand UO_4296 (O_4296,N_49988,N_48327);
xor UO_4297 (O_4297,N_49051,N_49117);
or UO_4298 (O_4298,N_49434,N_49905);
or UO_4299 (O_4299,N_48724,N_49079);
xnor UO_4300 (O_4300,N_48310,N_48368);
xor UO_4301 (O_4301,N_49299,N_49969);
and UO_4302 (O_4302,N_48384,N_48043);
nand UO_4303 (O_4303,N_48770,N_49497);
and UO_4304 (O_4304,N_49037,N_48455);
nand UO_4305 (O_4305,N_48999,N_48504);
or UO_4306 (O_4306,N_49213,N_48921);
nor UO_4307 (O_4307,N_49150,N_49510);
nor UO_4308 (O_4308,N_48476,N_49130);
nor UO_4309 (O_4309,N_48532,N_48792);
or UO_4310 (O_4310,N_49640,N_49118);
nand UO_4311 (O_4311,N_49949,N_48696);
xor UO_4312 (O_4312,N_49256,N_48615);
nand UO_4313 (O_4313,N_49235,N_49349);
or UO_4314 (O_4314,N_49339,N_48683);
nor UO_4315 (O_4315,N_49734,N_49476);
and UO_4316 (O_4316,N_49543,N_48262);
and UO_4317 (O_4317,N_49843,N_48725);
or UO_4318 (O_4318,N_48104,N_49423);
nand UO_4319 (O_4319,N_48098,N_49852);
xnor UO_4320 (O_4320,N_49823,N_48302);
nand UO_4321 (O_4321,N_48382,N_49040);
or UO_4322 (O_4322,N_48116,N_49717);
nor UO_4323 (O_4323,N_48833,N_48609);
xnor UO_4324 (O_4324,N_49030,N_49392);
xor UO_4325 (O_4325,N_49062,N_49293);
nand UO_4326 (O_4326,N_49476,N_48798);
and UO_4327 (O_4327,N_48312,N_48038);
nor UO_4328 (O_4328,N_48181,N_49783);
or UO_4329 (O_4329,N_49970,N_49425);
xor UO_4330 (O_4330,N_49271,N_48069);
and UO_4331 (O_4331,N_48920,N_48824);
nand UO_4332 (O_4332,N_48919,N_49362);
nor UO_4333 (O_4333,N_49422,N_49288);
nand UO_4334 (O_4334,N_49909,N_49960);
xnor UO_4335 (O_4335,N_49593,N_48483);
nand UO_4336 (O_4336,N_48303,N_48817);
nor UO_4337 (O_4337,N_49936,N_48802);
nor UO_4338 (O_4338,N_49505,N_49324);
nor UO_4339 (O_4339,N_49454,N_49427);
or UO_4340 (O_4340,N_49503,N_48137);
nand UO_4341 (O_4341,N_49260,N_49705);
nand UO_4342 (O_4342,N_48901,N_48225);
xor UO_4343 (O_4343,N_49124,N_49199);
and UO_4344 (O_4344,N_49596,N_48910);
or UO_4345 (O_4345,N_48147,N_49710);
and UO_4346 (O_4346,N_48840,N_48771);
nor UO_4347 (O_4347,N_49177,N_48792);
nand UO_4348 (O_4348,N_49681,N_48469);
nand UO_4349 (O_4349,N_49109,N_49231);
and UO_4350 (O_4350,N_49997,N_48780);
xnor UO_4351 (O_4351,N_48500,N_49100);
nor UO_4352 (O_4352,N_48981,N_48004);
or UO_4353 (O_4353,N_48590,N_49949);
xnor UO_4354 (O_4354,N_49161,N_48065);
nand UO_4355 (O_4355,N_48642,N_48797);
and UO_4356 (O_4356,N_48257,N_48114);
and UO_4357 (O_4357,N_49493,N_49406);
nor UO_4358 (O_4358,N_49025,N_49802);
nor UO_4359 (O_4359,N_49995,N_49802);
nand UO_4360 (O_4360,N_49280,N_48663);
nor UO_4361 (O_4361,N_48002,N_49630);
and UO_4362 (O_4362,N_49588,N_48432);
and UO_4363 (O_4363,N_48149,N_49903);
or UO_4364 (O_4364,N_48383,N_49474);
nand UO_4365 (O_4365,N_48615,N_49407);
nand UO_4366 (O_4366,N_49691,N_49657);
and UO_4367 (O_4367,N_48795,N_49162);
nand UO_4368 (O_4368,N_48895,N_48657);
or UO_4369 (O_4369,N_49509,N_49446);
or UO_4370 (O_4370,N_48979,N_49845);
nand UO_4371 (O_4371,N_49731,N_49651);
nand UO_4372 (O_4372,N_48593,N_48740);
xor UO_4373 (O_4373,N_49974,N_49932);
or UO_4374 (O_4374,N_49209,N_48646);
nand UO_4375 (O_4375,N_49895,N_49458);
nand UO_4376 (O_4376,N_49055,N_49602);
nor UO_4377 (O_4377,N_48426,N_48677);
xor UO_4378 (O_4378,N_49070,N_48336);
xor UO_4379 (O_4379,N_49248,N_49676);
or UO_4380 (O_4380,N_49983,N_48138);
and UO_4381 (O_4381,N_48752,N_49219);
xor UO_4382 (O_4382,N_49122,N_48199);
or UO_4383 (O_4383,N_48395,N_49655);
or UO_4384 (O_4384,N_48330,N_49672);
xnor UO_4385 (O_4385,N_49659,N_48766);
nor UO_4386 (O_4386,N_49694,N_48016);
nand UO_4387 (O_4387,N_48800,N_49549);
and UO_4388 (O_4388,N_48147,N_49364);
nor UO_4389 (O_4389,N_49657,N_48183);
and UO_4390 (O_4390,N_48550,N_49254);
or UO_4391 (O_4391,N_48503,N_49181);
and UO_4392 (O_4392,N_48073,N_48623);
nand UO_4393 (O_4393,N_49500,N_48886);
nor UO_4394 (O_4394,N_48545,N_49093);
and UO_4395 (O_4395,N_48915,N_48556);
or UO_4396 (O_4396,N_48171,N_48684);
and UO_4397 (O_4397,N_48179,N_48394);
nand UO_4398 (O_4398,N_49542,N_49624);
and UO_4399 (O_4399,N_49051,N_48587);
or UO_4400 (O_4400,N_48952,N_48324);
and UO_4401 (O_4401,N_48714,N_49986);
or UO_4402 (O_4402,N_49415,N_48754);
nand UO_4403 (O_4403,N_49819,N_49530);
nor UO_4404 (O_4404,N_49019,N_48044);
nand UO_4405 (O_4405,N_49050,N_49833);
and UO_4406 (O_4406,N_49714,N_48198);
nand UO_4407 (O_4407,N_48073,N_49672);
or UO_4408 (O_4408,N_49967,N_48761);
xor UO_4409 (O_4409,N_49625,N_49506);
and UO_4410 (O_4410,N_48337,N_49603);
nor UO_4411 (O_4411,N_48407,N_49654);
and UO_4412 (O_4412,N_48314,N_48993);
xor UO_4413 (O_4413,N_48352,N_48849);
and UO_4414 (O_4414,N_49694,N_48005);
nand UO_4415 (O_4415,N_48238,N_49863);
xnor UO_4416 (O_4416,N_48403,N_49672);
nor UO_4417 (O_4417,N_49966,N_48934);
nand UO_4418 (O_4418,N_49410,N_49790);
nor UO_4419 (O_4419,N_49903,N_48721);
nand UO_4420 (O_4420,N_48458,N_49191);
nand UO_4421 (O_4421,N_48677,N_48273);
and UO_4422 (O_4422,N_49276,N_48432);
and UO_4423 (O_4423,N_48154,N_49665);
nand UO_4424 (O_4424,N_49561,N_48958);
nand UO_4425 (O_4425,N_48727,N_48862);
nor UO_4426 (O_4426,N_49225,N_48055);
nand UO_4427 (O_4427,N_49859,N_48344);
or UO_4428 (O_4428,N_49813,N_48939);
and UO_4429 (O_4429,N_48320,N_48456);
or UO_4430 (O_4430,N_48059,N_48920);
or UO_4431 (O_4431,N_49017,N_49125);
nor UO_4432 (O_4432,N_49697,N_49659);
xnor UO_4433 (O_4433,N_48636,N_49584);
or UO_4434 (O_4434,N_48917,N_48438);
or UO_4435 (O_4435,N_49069,N_48949);
and UO_4436 (O_4436,N_49208,N_48485);
and UO_4437 (O_4437,N_48282,N_48354);
or UO_4438 (O_4438,N_48041,N_48521);
and UO_4439 (O_4439,N_48400,N_48484);
xnor UO_4440 (O_4440,N_49519,N_49791);
xor UO_4441 (O_4441,N_49147,N_49895);
nor UO_4442 (O_4442,N_48965,N_48231);
xnor UO_4443 (O_4443,N_48313,N_49578);
nor UO_4444 (O_4444,N_49378,N_48579);
nand UO_4445 (O_4445,N_48398,N_49944);
and UO_4446 (O_4446,N_49536,N_49064);
and UO_4447 (O_4447,N_49924,N_49496);
nor UO_4448 (O_4448,N_49152,N_49148);
nand UO_4449 (O_4449,N_48649,N_48801);
and UO_4450 (O_4450,N_49536,N_49055);
or UO_4451 (O_4451,N_49515,N_49354);
nand UO_4452 (O_4452,N_49792,N_48229);
and UO_4453 (O_4453,N_49694,N_49413);
nand UO_4454 (O_4454,N_48993,N_48306);
xor UO_4455 (O_4455,N_48195,N_49767);
and UO_4456 (O_4456,N_49131,N_49508);
xnor UO_4457 (O_4457,N_49704,N_49387);
nand UO_4458 (O_4458,N_48781,N_48591);
nand UO_4459 (O_4459,N_48500,N_49243);
nand UO_4460 (O_4460,N_48377,N_49864);
or UO_4461 (O_4461,N_49217,N_49578);
and UO_4462 (O_4462,N_49505,N_48702);
or UO_4463 (O_4463,N_49711,N_48001);
xnor UO_4464 (O_4464,N_48233,N_48905);
and UO_4465 (O_4465,N_48717,N_48447);
or UO_4466 (O_4466,N_48750,N_49490);
and UO_4467 (O_4467,N_48041,N_48164);
and UO_4468 (O_4468,N_49381,N_48459);
nor UO_4469 (O_4469,N_48548,N_48295);
and UO_4470 (O_4470,N_48698,N_49695);
or UO_4471 (O_4471,N_49087,N_49042);
nor UO_4472 (O_4472,N_49396,N_49306);
nand UO_4473 (O_4473,N_49773,N_48269);
nand UO_4474 (O_4474,N_48826,N_48783);
and UO_4475 (O_4475,N_48598,N_49182);
or UO_4476 (O_4476,N_48471,N_48098);
xor UO_4477 (O_4477,N_48514,N_49168);
nand UO_4478 (O_4478,N_48435,N_48243);
xor UO_4479 (O_4479,N_48826,N_48140);
nor UO_4480 (O_4480,N_48738,N_48613);
and UO_4481 (O_4481,N_48876,N_49908);
and UO_4482 (O_4482,N_49528,N_49141);
and UO_4483 (O_4483,N_49035,N_49194);
or UO_4484 (O_4484,N_49384,N_48180);
nor UO_4485 (O_4485,N_49919,N_48992);
and UO_4486 (O_4486,N_48204,N_49360);
nor UO_4487 (O_4487,N_49531,N_49360);
or UO_4488 (O_4488,N_48826,N_48821);
xnor UO_4489 (O_4489,N_48858,N_48288);
xor UO_4490 (O_4490,N_48003,N_48060);
xnor UO_4491 (O_4491,N_49435,N_48191);
xnor UO_4492 (O_4492,N_48460,N_49525);
nand UO_4493 (O_4493,N_48800,N_48524);
and UO_4494 (O_4494,N_48766,N_49348);
and UO_4495 (O_4495,N_48146,N_49440);
nand UO_4496 (O_4496,N_49553,N_48139);
nand UO_4497 (O_4497,N_49642,N_48377);
nor UO_4498 (O_4498,N_49662,N_49401);
or UO_4499 (O_4499,N_48413,N_49906);
or UO_4500 (O_4500,N_48200,N_48224);
nand UO_4501 (O_4501,N_49984,N_48241);
xnor UO_4502 (O_4502,N_49744,N_49798);
xnor UO_4503 (O_4503,N_48127,N_49220);
nor UO_4504 (O_4504,N_48839,N_49717);
xnor UO_4505 (O_4505,N_49669,N_49418);
nand UO_4506 (O_4506,N_49626,N_48086);
nor UO_4507 (O_4507,N_49414,N_48467);
nand UO_4508 (O_4508,N_49843,N_49016);
nor UO_4509 (O_4509,N_49668,N_48966);
or UO_4510 (O_4510,N_48775,N_48814);
xnor UO_4511 (O_4511,N_49591,N_48796);
and UO_4512 (O_4512,N_48136,N_49307);
or UO_4513 (O_4513,N_49536,N_49862);
nor UO_4514 (O_4514,N_48862,N_49222);
xor UO_4515 (O_4515,N_48745,N_48092);
or UO_4516 (O_4516,N_49730,N_48721);
nand UO_4517 (O_4517,N_49643,N_49586);
xnor UO_4518 (O_4518,N_49337,N_48861);
nand UO_4519 (O_4519,N_48864,N_49228);
or UO_4520 (O_4520,N_48089,N_48069);
nor UO_4521 (O_4521,N_49307,N_48497);
or UO_4522 (O_4522,N_48334,N_48944);
or UO_4523 (O_4523,N_49147,N_49923);
nor UO_4524 (O_4524,N_48228,N_48070);
nand UO_4525 (O_4525,N_48428,N_49707);
nand UO_4526 (O_4526,N_48888,N_49360);
or UO_4527 (O_4527,N_48536,N_48262);
or UO_4528 (O_4528,N_48514,N_48097);
and UO_4529 (O_4529,N_48977,N_48262);
nand UO_4530 (O_4530,N_48496,N_49482);
and UO_4531 (O_4531,N_49555,N_49522);
nand UO_4532 (O_4532,N_48905,N_48637);
xor UO_4533 (O_4533,N_49453,N_49938);
or UO_4534 (O_4534,N_49645,N_49790);
or UO_4535 (O_4535,N_49024,N_48827);
xor UO_4536 (O_4536,N_48885,N_48371);
or UO_4537 (O_4537,N_48810,N_48259);
xnor UO_4538 (O_4538,N_49141,N_48351);
and UO_4539 (O_4539,N_48255,N_48384);
xor UO_4540 (O_4540,N_48713,N_49883);
nor UO_4541 (O_4541,N_49484,N_48818);
or UO_4542 (O_4542,N_48821,N_48389);
or UO_4543 (O_4543,N_48367,N_48960);
xnor UO_4544 (O_4544,N_48429,N_48401);
nand UO_4545 (O_4545,N_48369,N_48584);
nor UO_4546 (O_4546,N_49060,N_49981);
nor UO_4547 (O_4547,N_49896,N_49532);
nor UO_4548 (O_4548,N_49886,N_48503);
or UO_4549 (O_4549,N_49101,N_49913);
xnor UO_4550 (O_4550,N_48476,N_49494);
nand UO_4551 (O_4551,N_48171,N_48064);
and UO_4552 (O_4552,N_48728,N_48111);
and UO_4553 (O_4553,N_49576,N_49345);
nand UO_4554 (O_4554,N_48594,N_49645);
nand UO_4555 (O_4555,N_48479,N_48197);
nand UO_4556 (O_4556,N_49577,N_49530);
nor UO_4557 (O_4557,N_48742,N_49122);
or UO_4558 (O_4558,N_48565,N_49540);
or UO_4559 (O_4559,N_49766,N_48154);
nor UO_4560 (O_4560,N_49104,N_48552);
xor UO_4561 (O_4561,N_49188,N_49579);
nand UO_4562 (O_4562,N_48151,N_48476);
or UO_4563 (O_4563,N_48408,N_49343);
xor UO_4564 (O_4564,N_49148,N_48038);
nor UO_4565 (O_4565,N_48662,N_49991);
and UO_4566 (O_4566,N_49055,N_48474);
nand UO_4567 (O_4567,N_48144,N_48620);
or UO_4568 (O_4568,N_49811,N_49813);
xnor UO_4569 (O_4569,N_49776,N_49301);
nor UO_4570 (O_4570,N_48515,N_49374);
and UO_4571 (O_4571,N_48454,N_49053);
nor UO_4572 (O_4572,N_49483,N_48487);
xnor UO_4573 (O_4573,N_49008,N_48763);
or UO_4574 (O_4574,N_48007,N_49536);
nor UO_4575 (O_4575,N_48335,N_48078);
or UO_4576 (O_4576,N_48583,N_48190);
and UO_4577 (O_4577,N_49162,N_49218);
nand UO_4578 (O_4578,N_49391,N_49184);
and UO_4579 (O_4579,N_49224,N_49661);
or UO_4580 (O_4580,N_48747,N_49771);
xor UO_4581 (O_4581,N_48776,N_48156);
nand UO_4582 (O_4582,N_49520,N_48277);
nor UO_4583 (O_4583,N_49647,N_48137);
and UO_4584 (O_4584,N_49257,N_49345);
xor UO_4585 (O_4585,N_48140,N_49645);
xor UO_4586 (O_4586,N_48810,N_49332);
xor UO_4587 (O_4587,N_48905,N_48805);
nand UO_4588 (O_4588,N_48386,N_48679);
and UO_4589 (O_4589,N_49328,N_48946);
nand UO_4590 (O_4590,N_48196,N_48342);
nand UO_4591 (O_4591,N_49847,N_48347);
xor UO_4592 (O_4592,N_48811,N_49224);
and UO_4593 (O_4593,N_48493,N_48563);
nand UO_4594 (O_4594,N_48185,N_49977);
xnor UO_4595 (O_4595,N_49711,N_49779);
nor UO_4596 (O_4596,N_48244,N_48534);
nand UO_4597 (O_4597,N_49463,N_48788);
nor UO_4598 (O_4598,N_48168,N_48781);
or UO_4599 (O_4599,N_48446,N_49153);
and UO_4600 (O_4600,N_49160,N_48860);
xnor UO_4601 (O_4601,N_49918,N_49080);
nand UO_4602 (O_4602,N_48152,N_49078);
or UO_4603 (O_4603,N_48268,N_48780);
or UO_4604 (O_4604,N_48204,N_48096);
or UO_4605 (O_4605,N_49321,N_48675);
nand UO_4606 (O_4606,N_48938,N_48985);
nor UO_4607 (O_4607,N_48306,N_49007);
nor UO_4608 (O_4608,N_48853,N_49707);
or UO_4609 (O_4609,N_48014,N_49746);
nand UO_4610 (O_4610,N_49876,N_48930);
nor UO_4611 (O_4611,N_49401,N_49446);
or UO_4612 (O_4612,N_49888,N_48139);
nand UO_4613 (O_4613,N_49371,N_48215);
nor UO_4614 (O_4614,N_49873,N_48263);
nor UO_4615 (O_4615,N_49337,N_49402);
and UO_4616 (O_4616,N_48050,N_49918);
or UO_4617 (O_4617,N_48208,N_49978);
or UO_4618 (O_4618,N_48049,N_48969);
and UO_4619 (O_4619,N_48757,N_49607);
nand UO_4620 (O_4620,N_48768,N_48691);
xnor UO_4621 (O_4621,N_49447,N_48736);
nand UO_4622 (O_4622,N_49952,N_49066);
and UO_4623 (O_4623,N_49714,N_49909);
xnor UO_4624 (O_4624,N_48051,N_49937);
or UO_4625 (O_4625,N_49564,N_48865);
nand UO_4626 (O_4626,N_48104,N_49897);
or UO_4627 (O_4627,N_48751,N_49732);
or UO_4628 (O_4628,N_49305,N_49213);
xnor UO_4629 (O_4629,N_48930,N_48246);
nor UO_4630 (O_4630,N_49144,N_48834);
nor UO_4631 (O_4631,N_49977,N_48200);
and UO_4632 (O_4632,N_49262,N_49405);
xnor UO_4633 (O_4633,N_48813,N_49060);
nor UO_4634 (O_4634,N_48473,N_48729);
and UO_4635 (O_4635,N_49287,N_49225);
or UO_4636 (O_4636,N_48161,N_48550);
nand UO_4637 (O_4637,N_49642,N_48418);
nand UO_4638 (O_4638,N_48256,N_48117);
nand UO_4639 (O_4639,N_49481,N_48192);
or UO_4640 (O_4640,N_48830,N_49988);
nor UO_4641 (O_4641,N_48805,N_48710);
or UO_4642 (O_4642,N_48936,N_49067);
or UO_4643 (O_4643,N_48376,N_48098);
nand UO_4644 (O_4644,N_49921,N_49685);
xor UO_4645 (O_4645,N_49134,N_49594);
xnor UO_4646 (O_4646,N_49877,N_49180);
or UO_4647 (O_4647,N_49098,N_49932);
nor UO_4648 (O_4648,N_49406,N_49105);
or UO_4649 (O_4649,N_49166,N_49883);
nand UO_4650 (O_4650,N_49171,N_48187);
or UO_4651 (O_4651,N_48373,N_49201);
nand UO_4652 (O_4652,N_48131,N_48305);
xnor UO_4653 (O_4653,N_49053,N_48764);
and UO_4654 (O_4654,N_49465,N_48804);
or UO_4655 (O_4655,N_48754,N_49940);
nor UO_4656 (O_4656,N_48899,N_49418);
nor UO_4657 (O_4657,N_48558,N_48683);
nand UO_4658 (O_4658,N_48464,N_48194);
and UO_4659 (O_4659,N_48422,N_49555);
nand UO_4660 (O_4660,N_48793,N_48176);
and UO_4661 (O_4661,N_48824,N_48333);
nand UO_4662 (O_4662,N_49355,N_48140);
nor UO_4663 (O_4663,N_49328,N_49859);
and UO_4664 (O_4664,N_48996,N_48992);
nand UO_4665 (O_4665,N_48593,N_48314);
and UO_4666 (O_4666,N_49022,N_48981);
nor UO_4667 (O_4667,N_48963,N_48077);
nand UO_4668 (O_4668,N_48928,N_49965);
nor UO_4669 (O_4669,N_49735,N_48997);
nand UO_4670 (O_4670,N_49422,N_48569);
nand UO_4671 (O_4671,N_49514,N_48046);
and UO_4672 (O_4672,N_49643,N_49101);
and UO_4673 (O_4673,N_48094,N_48893);
xor UO_4674 (O_4674,N_48438,N_49287);
and UO_4675 (O_4675,N_49997,N_48236);
and UO_4676 (O_4676,N_48056,N_48040);
nor UO_4677 (O_4677,N_49355,N_48683);
nor UO_4678 (O_4678,N_48366,N_48182);
or UO_4679 (O_4679,N_49974,N_49541);
nor UO_4680 (O_4680,N_49896,N_49290);
and UO_4681 (O_4681,N_49876,N_49588);
nor UO_4682 (O_4682,N_49041,N_49784);
and UO_4683 (O_4683,N_49898,N_49376);
and UO_4684 (O_4684,N_48964,N_49700);
xor UO_4685 (O_4685,N_49227,N_49403);
or UO_4686 (O_4686,N_49354,N_48579);
nor UO_4687 (O_4687,N_48596,N_49012);
or UO_4688 (O_4688,N_48500,N_48527);
or UO_4689 (O_4689,N_48663,N_48151);
nand UO_4690 (O_4690,N_49182,N_48696);
and UO_4691 (O_4691,N_48227,N_48063);
xnor UO_4692 (O_4692,N_48264,N_48852);
nor UO_4693 (O_4693,N_49382,N_49851);
and UO_4694 (O_4694,N_49287,N_49195);
xor UO_4695 (O_4695,N_48460,N_49439);
xnor UO_4696 (O_4696,N_49946,N_49793);
or UO_4697 (O_4697,N_48441,N_48342);
nand UO_4698 (O_4698,N_48449,N_48822);
or UO_4699 (O_4699,N_49716,N_49577);
and UO_4700 (O_4700,N_49453,N_48516);
nand UO_4701 (O_4701,N_49396,N_48656);
or UO_4702 (O_4702,N_48384,N_48272);
nor UO_4703 (O_4703,N_48160,N_48916);
and UO_4704 (O_4704,N_48380,N_48344);
xor UO_4705 (O_4705,N_49427,N_48935);
and UO_4706 (O_4706,N_48748,N_49575);
xnor UO_4707 (O_4707,N_49735,N_48749);
xor UO_4708 (O_4708,N_48868,N_48471);
nor UO_4709 (O_4709,N_49412,N_49917);
nor UO_4710 (O_4710,N_48897,N_49364);
or UO_4711 (O_4711,N_49627,N_48896);
nor UO_4712 (O_4712,N_48427,N_49396);
nor UO_4713 (O_4713,N_49160,N_49905);
xnor UO_4714 (O_4714,N_49200,N_49078);
xor UO_4715 (O_4715,N_48335,N_48511);
nor UO_4716 (O_4716,N_48106,N_49619);
nand UO_4717 (O_4717,N_49340,N_49055);
nand UO_4718 (O_4718,N_49946,N_48863);
or UO_4719 (O_4719,N_48351,N_49730);
or UO_4720 (O_4720,N_48522,N_48131);
xor UO_4721 (O_4721,N_49255,N_48202);
nand UO_4722 (O_4722,N_48402,N_48838);
nand UO_4723 (O_4723,N_48532,N_49431);
and UO_4724 (O_4724,N_49923,N_49718);
xnor UO_4725 (O_4725,N_48498,N_48270);
nor UO_4726 (O_4726,N_49296,N_49253);
xor UO_4727 (O_4727,N_48903,N_48902);
or UO_4728 (O_4728,N_48310,N_48980);
or UO_4729 (O_4729,N_48177,N_49324);
or UO_4730 (O_4730,N_49251,N_48746);
nor UO_4731 (O_4731,N_49477,N_49908);
nand UO_4732 (O_4732,N_48218,N_48334);
xor UO_4733 (O_4733,N_49772,N_48578);
nor UO_4734 (O_4734,N_49544,N_49220);
nor UO_4735 (O_4735,N_48129,N_49480);
nand UO_4736 (O_4736,N_49137,N_49413);
nand UO_4737 (O_4737,N_49805,N_49978);
and UO_4738 (O_4738,N_48404,N_48894);
xor UO_4739 (O_4739,N_48852,N_48822);
nand UO_4740 (O_4740,N_49191,N_48240);
nand UO_4741 (O_4741,N_48380,N_49859);
xor UO_4742 (O_4742,N_49129,N_48608);
nand UO_4743 (O_4743,N_48512,N_48037);
nor UO_4744 (O_4744,N_49047,N_48408);
nor UO_4745 (O_4745,N_49544,N_48096);
or UO_4746 (O_4746,N_49050,N_49217);
xnor UO_4747 (O_4747,N_49088,N_48599);
or UO_4748 (O_4748,N_48546,N_48180);
nand UO_4749 (O_4749,N_48730,N_48217);
or UO_4750 (O_4750,N_49766,N_48075);
nand UO_4751 (O_4751,N_48642,N_49534);
or UO_4752 (O_4752,N_48244,N_48228);
xnor UO_4753 (O_4753,N_49461,N_49782);
nand UO_4754 (O_4754,N_48543,N_48342);
or UO_4755 (O_4755,N_48352,N_48627);
nand UO_4756 (O_4756,N_48477,N_49938);
xnor UO_4757 (O_4757,N_49468,N_49712);
nand UO_4758 (O_4758,N_49335,N_48240);
xor UO_4759 (O_4759,N_48531,N_48105);
nor UO_4760 (O_4760,N_49499,N_48891);
and UO_4761 (O_4761,N_49367,N_48225);
nor UO_4762 (O_4762,N_49491,N_49857);
nor UO_4763 (O_4763,N_49355,N_48244);
xnor UO_4764 (O_4764,N_49221,N_48357);
nand UO_4765 (O_4765,N_48259,N_48784);
xor UO_4766 (O_4766,N_49257,N_48914);
or UO_4767 (O_4767,N_49956,N_48007);
and UO_4768 (O_4768,N_49569,N_49825);
xor UO_4769 (O_4769,N_49470,N_48669);
nand UO_4770 (O_4770,N_48019,N_49025);
or UO_4771 (O_4771,N_48797,N_48799);
and UO_4772 (O_4772,N_49291,N_48090);
xor UO_4773 (O_4773,N_49595,N_48892);
or UO_4774 (O_4774,N_48597,N_48803);
nor UO_4775 (O_4775,N_49744,N_48077);
xor UO_4776 (O_4776,N_48177,N_49200);
nor UO_4777 (O_4777,N_48652,N_48223);
and UO_4778 (O_4778,N_49115,N_49719);
xor UO_4779 (O_4779,N_49879,N_49299);
or UO_4780 (O_4780,N_48720,N_48460);
xnor UO_4781 (O_4781,N_48007,N_48667);
or UO_4782 (O_4782,N_49156,N_48573);
nand UO_4783 (O_4783,N_48753,N_49193);
xnor UO_4784 (O_4784,N_48298,N_48489);
and UO_4785 (O_4785,N_48179,N_48139);
or UO_4786 (O_4786,N_48652,N_49788);
nand UO_4787 (O_4787,N_49060,N_48058);
and UO_4788 (O_4788,N_48616,N_49791);
or UO_4789 (O_4789,N_49213,N_49670);
xnor UO_4790 (O_4790,N_49332,N_49612);
nand UO_4791 (O_4791,N_49037,N_48853);
nor UO_4792 (O_4792,N_49852,N_49363);
and UO_4793 (O_4793,N_48693,N_49830);
nor UO_4794 (O_4794,N_49412,N_48599);
or UO_4795 (O_4795,N_49138,N_48943);
and UO_4796 (O_4796,N_48788,N_49874);
and UO_4797 (O_4797,N_49931,N_48017);
nand UO_4798 (O_4798,N_48372,N_48763);
nor UO_4799 (O_4799,N_48371,N_49461);
or UO_4800 (O_4800,N_48654,N_48669);
nor UO_4801 (O_4801,N_49899,N_49224);
nand UO_4802 (O_4802,N_49417,N_48219);
or UO_4803 (O_4803,N_48744,N_49528);
or UO_4804 (O_4804,N_48819,N_49531);
nor UO_4805 (O_4805,N_48352,N_48233);
nand UO_4806 (O_4806,N_48519,N_48666);
xor UO_4807 (O_4807,N_48519,N_48498);
nand UO_4808 (O_4808,N_48195,N_48023);
and UO_4809 (O_4809,N_49783,N_48942);
nand UO_4810 (O_4810,N_49652,N_49060);
or UO_4811 (O_4811,N_49540,N_49936);
or UO_4812 (O_4812,N_48370,N_48279);
or UO_4813 (O_4813,N_49032,N_48120);
xnor UO_4814 (O_4814,N_49264,N_48264);
and UO_4815 (O_4815,N_48567,N_48943);
and UO_4816 (O_4816,N_48345,N_49910);
nand UO_4817 (O_4817,N_49727,N_48489);
xnor UO_4818 (O_4818,N_48275,N_49030);
or UO_4819 (O_4819,N_48935,N_48399);
nor UO_4820 (O_4820,N_48185,N_48365);
nor UO_4821 (O_4821,N_49799,N_49488);
and UO_4822 (O_4822,N_49875,N_48135);
and UO_4823 (O_4823,N_49692,N_49048);
nor UO_4824 (O_4824,N_48326,N_49974);
xnor UO_4825 (O_4825,N_49040,N_48961);
nor UO_4826 (O_4826,N_49453,N_48402);
nor UO_4827 (O_4827,N_49938,N_49286);
xnor UO_4828 (O_4828,N_49971,N_48102);
nor UO_4829 (O_4829,N_49229,N_49176);
nand UO_4830 (O_4830,N_48566,N_48945);
nor UO_4831 (O_4831,N_48741,N_49134);
or UO_4832 (O_4832,N_49026,N_49831);
nand UO_4833 (O_4833,N_49986,N_49736);
nand UO_4834 (O_4834,N_49727,N_48975);
xor UO_4835 (O_4835,N_48468,N_48488);
or UO_4836 (O_4836,N_48899,N_49762);
nor UO_4837 (O_4837,N_48267,N_48385);
nand UO_4838 (O_4838,N_48520,N_49678);
xor UO_4839 (O_4839,N_48799,N_49551);
nand UO_4840 (O_4840,N_48897,N_49616);
nor UO_4841 (O_4841,N_48077,N_49419);
xor UO_4842 (O_4842,N_49897,N_48946);
and UO_4843 (O_4843,N_49129,N_48990);
xnor UO_4844 (O_4844,N_49244,N_49906);
or UO_4845 (O_4845,N_49929,N_49645);
or UO_4846 (O_4846,N_48506,N_48778);
and UO_4847 (O_4847,N_49318,N_49674);
nand UO_4848 (O_4848,N_48674,N_49621);
nand UO_4849 (O_4849,N_49935,N_49509);
xnor UO_4850 (O_4850,N_49713,N_49044);
or UO_4851 (O_4851,N_48397,N_48848);
xnor UO_4852 (O_4852,N_49905,N_49551);
and UO_4853 (O_4853,N_49926,N_48326);
nor UO_4854 (O_4854,N_49648,N_49143);
or UO_4855 (O_4855,N_49025,N_49112);
or UO_4856 (O_4856,N_49986,N_49700);
and UO_4857 (O_4857,N_48931,N_49957);
or UO_4858 (O_4858,N_48251,N_48509);
or UO_4859 (O_4859,N_49939,N_49929);
xor UO_4860 (O_4860,N_49630,N_48392);
and UO_4861 (O_4861,N_49356,N_49741);
nand UO_4862 (O_4862,N_48986,N_49291);
nand UO_4863 (O_4863,N_49528,N_48270);
nand UO_4864 (O_4864,N_49591,N_48698);
nor UO_4865 (O_4865,N_49030,N_49159);
and UO_4866 (O_4866,N_48293,N_49667);
xnor UO_4867 (O_4867,N_48701,N_49194);
nor UO_4868 (O_4868,N_48342,N_49258);
and UO_4869 (O_4869,N_49608,N_49790);
xor UO_4870 (O_4870,N_49131,N_48266);
xor UO_4871 (O_4871,N_48286,N_48017);
nand UO_4872 (O_4872,N_49993,N_49692);
and UO_4873 (O_4873,N_48993,N_48037);
xnor UO_4874 (O_4874,N_48664,N_49991);
and UO_4875 (O_4875,N_49257,N_48018);
xor UO_4876 (O_4876,N_48815,N_48886);
nor UO_4877 (O_4877,N_49296,N_49996);
or UO_4878 (O_4878,N_48116,N_49322);
and UO_4879 (O_4879,N_49575,N_48069);
nand UO_4880 (O_4880,N_48247,N_48166);
nor UO_4881 (O_4881,N_49298,N_48802);
nor UO_4882 (O_4882,N_48771,N_48704);
and UO_4883 (O_4883,N_48940,N_48979);
and UO_4884 (O_4884,N_48310,N_49540);
and UO_4885 (O_4885,N_49729,N_48645);
nand UO_4886 (O_4886,N_49218,N_48062);
nand UO_4887 (O_4887,N_48281,N_48181);
and UO_4888 (O_4888,N_48024,N_49917);
xor UO_4889 (O_4889,N_48047,N_48808);
and UO_4890 (O_4890,N_48761,N_49806);
nand UO_4891 (O_4891,N_49929,N_49525);
and UO_4892 (O_4892,N_49181,N_48648);
and UO_4893 (O_4893,N_49712,N_49556);
nor UO_4894 (O_4894,N_48216,N_49643);
or UO_4895 (O_4895,N_48616,N_48582);
and UO_4896 (O_4896,N_48836,N_48274);
or UO_4897 (O_4897,N_49647,N_48613);
nor UO_4898 (O_4898,N_48539,N_49884);
nand UO_4899 (O_4899,N_49409,N_48433);
or UO_4900 (O_4900,N_49446,N_49568);
or UO_4901 (O_4901,N_49698,N_49318);
or UO_4902 (O_4902,N_49813,N_49425);
xor UO_4903 (O_4903,N_49383,N_48069);
or UO_4904 (O_4904,N_48085,N_49090);
and UO_4905 (O_4905,N_49066,N_49437);
nor UO_4906 (O_4906,N_49606,N_49536);
and UO_4907 (O_4907,N_49614,N_49527);
and UO_4908 (O_4908,N_48120,N_49708);
nor UO_4909 (O_4909,N_49896,N_48448);
nor UO_4910 (O_4910,N_48131,N_48579);
and UO_4911 (O_4911,N_48553,N_48350);
nand UO_4912 (O_4912,N_49772,N_49343);
and UO_4913 (O_4913,N_48509,N_48352);
xnor UO_4914 (O_4914,N_49185,N_49977);
nand UO_4915 (O_4915,N_48878,N_48497);
nand UO_4916 (O_4916,N_49659,N_49209);
or UO_4917 (O_4917,N_49581,N_49500);
nand UO_4918 (O_4918,N_49990,N_48889);
xor UO_4919 (O_4919,N_49224,N_48647);
xnor UO_4920 (O_4920,N_48565,N_49102);
or UO_4921 (O_4921,N_49589,N_48354);
nor UO_4922 (O_4922,N_49378,N_48429);
nand UO_4923 (O_4923,N_48067,N_49108);
nand UO_4924 (O_4924,N_48094,N_48606);
nand UO_4925 (O_4925,N_48086,N_49477);
nand UO_4926 (O_4926,N_49692,N_48133);
nand UO_4927 (O_4927,N_48581,N_48625);
nand UO_4928 (O_4928,N_48305,N_49743);
nand UO_4929 (O_4929,N_48947,N_49517);
and UO_4930 (O_4930,N_48081,N_49429);
or UO_4931 (O_4931,N_49410,N_49974);
xor UO_4932 (O_4932,N_49335,N_48928);
nand UO_4933 (O_4933,N_49154,N_49789);
nand UO_4934 (O_4934,N_48465,N_49208);
nor UO_4935 (O_4935,N_48802,N_49665);
nor UO_4936 (O_4936,N_49751,N_49194);
xnor UO_4937 (O_4937,N_49135,N_49531);
nand UO_4938 (O_4938,N_48264,N_49904);
xor UO_4939 (O_4939,N_48980,N_49763);
and UO_4940 (O_4940,N_48160,N_49303);
or UO_4941 (O_4941,N_49060,N_48356);
and UO_4942 (O_4942,N_49733,N_48238);
nor UO_4943 (O_4943,N_48844,N_48090);
or UO_4944 (O_4944,N_48641,N_48401);
nor UO_4945 (O_4945,N_48689,N_48626);
or UO_4946 (O_4946,N_48763,N_48428);
or UO_4947 (O_4947,N_48977,N_49814);
or UO_4948 (O_4948,N_49746,N_48559);
nand UO_4949 (O_4949,N_48525,N_48759);
nor UO_4950 (O_4950,N_49856,N_48319);
xor UO_4951 (O_4951,N_48295,N_49757);
nand UO_4952 (O_4952,N_48298,N_49954);
or UO_4953 (O_4953,N_48174,N_49012);
xor UO_4954 (O_4954,N_49720,N_48087);
nor UO_4955 (O_4955,N_48368,N_49510);
nor UO_4956 (O_4956,N_48184,N_48413);
nor UO_4957 (O_4957,N_49949,N_48838);
nor UO_4958 (O_4958,N_48719,N_48402);
or UO_4959 (O_4959,N_48577,N_49357);
nor UO_4960 (O_4960,N_48317,N_49284);
xnor UO_4961 (O_4961,N_49988,N_48062);
xor UO_4962 (O_4962,N_49302,N_48485);
nand UO_4963 (O_4963,N_48772,N_49771);
xor UO_4964 (O_4964,N_49231,N_48054);
nor UO_4965 (O_4965,N_48313,N_48189);
or UO_4966 (O_4966,N_48029,N_48644);
nand UO_4967 (O_4967,N_49729,N_48774);
xnor UO_4968 (O_4968,N_49240,N_48928);
or UO_4969 (O_4969,N_48397,N_48020);
xnor UO_4970 (O_4970,N_48733,N_48981);
or UO_4971 (O_4971,N_48333,N_49245);
or UO_4972 (O_4972,N_49280,N_48722);
nand UO_4973 (O_4973,N_49044,N_48240);
xor UO_4974 (O_4974,N_48789,N_49548);
nor UO_4975 (O_4975,N_49655,N_49585);
and UO_4976 (O_4976,N_48708,N_49046);
and UO_4977 (O_4977,N_49271,N_49607);
nand UO_4978 (O_4978,N_49502,N_48926);
and UO_4979 (O_4979,N_48211,N_48089);
nor UO_4980 (O_4980,N_48262,N_49050);
nand UO_4981 (O_4981,N_48276,N_48516);
xnor UO_4982 (O_4982,N_48303,N_48274);
and UO_4983 (O_4983,N_48179,N_48093);
or UO_4984 (O_4984,N_48329,N_49127);
nand UO_4985 (O_4985,N_49370,N_49661);
nand UO_4986 (O_4986,N_48141,N_49538);
xor UO_4987 (O_4987,N_49571,N_48645);
and UO_4988 (O_4988,N_48961,N_49981);
or UO_4989 (O_4989,N_49776,N_48583);
or UO_4990 (O_4990,N_48653,N_48362);
nand UO_4991 (O_4991,N_49723,N_48291);
or UO_4992 (O_4992,N_48034,N_49001);
nor UO_4993 (O_4993,N_49258,N_49930);
nor UO_4994 (O_4994,N_49934,N_48618);
or UO_4995 (O_4995,N_48715,N_49774);
nand UO_4996 (O_4996,N_48575,N_49896);
xor UO_4997 (O_4997,N_48144,N_48501);
or UO_4998 (O_4998,N_48907,N_49709);
nor UO_4999 (O_4999,N_48256,N_48599);
endmodule