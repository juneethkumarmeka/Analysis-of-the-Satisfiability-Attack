module basic_500_3000_500_40_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xnor U0 (N_0,In_221,In_248);
or U1 (N_1,In_67,In_268);
xnor U2 (N_2,In_132,In_359);
and U3 (N_3,In_179,In_155);
and U4 (N_4,In_214,In_472);
xor U5 (N_5,In_360,In_143);
or U6 (N_6,In_120,In_471);
or U7 (N_7,In_452,In_31);
xnor U8 (N_8,In_401,In_117);
xnor U9 (N_9,In_498,In_178);
or U10 (N_10,In_449,In_261);
and U11 (N_11,In_157,In_84);
or U12 (N_12,In_108,In_48);
or U13 (N_13,In_349,In_144);
and U14 (N_14,In_455,In_38);
nor U15 (N_15,In_304,In_438);
xor U16 (N_16,In_297,In_152);
and U17 (N_17,In_126,In_239);
nor U18 (N_18,In_474,In_350);
xnor U19 (N_19,In_51,In_167);
nor U20 (N_20,In_34,In_54);
nor U21 (N_21,In_101,In_210);
or U22 (N_22,In_430,In_407);
nand U23 (N_23,In_41,In_104);
nand U24 (N_24,In_388,In_435);
xor U25 (N_25,In_122,In_212);
and U26 (N_26,In_436,In_105);
nand U27 (N_27,In_467,In_331);
or U28 (N_28,In_348,In_309);
nand U29 (N_29,In_247,In_137);
nand U30 (N_30,In_495,In_26);
and U31 (N_31,In_312,In_215);
xnor U32 (N_32,In_386,In_240);
and U33 (N_33,In_58,In_321);
nand U34 (N_34,In_202,In_280);
nor U35 (N_35,In_220,In_32);
or U36 (N_36,In_466,In_194);
xnor U37 (N_37,In_363,In_79);
and U38 (N_38,In_374,In_69);
nor U39 (N_39,In_113,In_400);
nor U40 (N_40,In_376,In_378);
nor U41 (N_41,In_302,In_476);
xor U42 (N_42,In_1,In_486);
and U43 (N_43,In_23,In_196);
and U44 (N_44,In_325,In_465);
xor U45 (N_45,In_477,In_170);
nor U46 (N_46,In_319,In_95);
nor U47 (N_47,In_237,In_209);
nand U48 (N_48,In_433,In_387);
or U49 (N_49,In_227,In_322);
xor U50 (N_50,In_50,In_255);
or U51 (N_51,In_3,In_372);
or U52 (N_52,In_90,In_2);
xor U53 (N_53,In_225,In_276);
or U54 (N_54,In_390,In_65);
nor U55 (N_55,In_417,In_480);
nand U56 (N_56,In_439,In_174);
nand U57 (N_57,In_217,In_173);
or U58 (N_58,In_56,In_269);
xor U59 (N_59,In_145,In_18);
and U60 (N_60,In_427,In_43);
nand U61 (N_61,In_238,In_94);
and U62 (N_62,In_182,In_263);
and U63 (N_63,In_442,In_409);
nor U64 (N_64,In_16,In_298);
or U65 (N_65,In_128,In_275);
nor U66 (N_66,In_460,In_421);
nand U67 (N_67,In_489,In_265);
or U68 (N_68,In_320,In_138);
xor U69 (N_69,In_245,In_20);
xnor U70 (N_70,In_149,In_30);
and U71 (N_71,In_335,In_246);
xnor U72 (N_72,In_166,In_469);
and U73 (N_73,In_461,In_334);
nor U74 (N_74,In_175,In_299);
xor U75 (N_75,In_326,In_395);
and U76 (N_76,N_22,In_192);
and U77 (N_77,In_499,N_55);
and U78 (N_78,In_42,In_340);
nand U79 (N_79,N_68,In_242);
nand U80 (N_80,In_211,N_52);
xnor U81 (N_81,In_154,In_483);
and U82 (N_82,In_347,In_102);
or U83 (N_83,In_267,In_140);
nor U84 (N_84,In_422,In_80);
or U85 (N_85,In_446,In_55);
xor U86 (N_86,In_141,In_163);
nor U87 (N_87,In_453,In_296);
nand U88 (N_88,In_100,In_381);
xnor U89 (N_89,In_253,In_291);
nand U90 (N_90,In_324,In_33);
xnor U91 (N_91,In_307,In_450);
xor U92 (N_92,N_50,In_169);
and U93 (N_93,In_234,In_270);
nand U94 (N_94,N_27,N_30);
nand U95 (N_95,In_497,In_463);
and U96 (N_96,In_345,In_44);
and U97 (N_97,N_18,In_464);
nand U98 (N_98,In_251,In_411);
or U99 (N_99,In_106,In_37);
and U100 (N_100,N_34,In_130);
nor U101 (N_101,In_156,In_481);
nand U102 (N_102,In_213,In_384);
or U103 (N_103,In_158,In_81);
nor U104 (N_104,In_15,In_29);
and U105 (N_105,In_431,N_40);
nor U106 (N_106,In_404,In_188);
nor U107 (N_107,In_236,In_279);
xnor U108 (N_108,In_164,N_45);
or U109 (N_109,In_17,In_457);
or U110 (N_110,In_468,In_162);
xor U111 (N_111,N_28,In_256);
nor U112 (N_112,In_456,In_496);
xnor U113 (N_113,In_60,In_216);
or U114 (N_114,N_6,In_235);
nand U115 (N_115,In_7,In_332);
and U116 (N_116,In_375,In_59);
and U117 (N_117,In_292,In_424);
and U118 (N_118,In_186,In_478);
nand U119 (N_119,In_73,In_273);
xnor U120 (N_120,In_159,In_147);
or U121 (N_121,N_62,In_11);
or U122 (N_122,In_412,In_189);
and U123 (N_123,In_208,In_77);
xnor U124 (N_124,In_254,In_379);
xnor U125 (N_125,In_370,In_98);
nand U126 (N_126,In_362,In_333);
nor U127 (N_127,N_33,In_46);
xor U128 (N_128,In_303,In_165);
xor U129 (N_129,N_41,In_306);
or U130 (N_130,In_364,In_9);
nor U131 (N_131,N_9,In_198);
xnor U132 (N_132,In_85,N_17);
nor U133 (N_133,In_328,In_64);
xnor U134 (N_134,In_199,In_89);
xor U135 (N_135,In_382,N_26);
nand U136 (N_136,In_207,In_408);
nor U137 (N_137,N_66,In_317);
and U138 (N_138,In_353,In_168);
or U139 (N_139,In_103,N_42);
nand U140 (N_140,In_301,In_160);
xnor U141 (N_141,In_419,N_70);
nor U142 (N_142,In_373,In_415);
and U143 (N_143,N_36,N_51);
nand U144 (N_144,N_67,In_330);
nor U145 (N_145,In_244,N_2);
nand U146 (N_146,In_288,N_29);
nand U147 (N_147,In_249,In_92);
or U148 (N_148,In_488,In_27);
or U149 (N_149,N_69,In_286);
xnor U150 (N_150,In_487,N_3);
xor U151 (N_151,In_62,N_112);
nand U152 (N_152,In_300,In_107);
nor U153 (N_153,N_104,N_4);
nand U154 (N_154,N_125,N_19);
nand U155 (N_155,N_138,In_368);
nand U156 (N_156,N_149,In_365);
and U157 (N_157,In_8,N_64);
and U158 (N_158,In_282,In_57);
and U159 (N_159,In_250,N_87);
and U160 (N_160,In_131,N_1);
nand U161 (N_161,In_39,N_72);
or U162 (N_162,N_61,In_318);
nor U163 (N_163,N_47,In_355);
nor U164 (N_164,In_351,In_204);
nor U165 (N_165,In_473,In_440);
xnor U166 (N_166,In_121,N_76);
xor U167 (N_167,In_284,N_113);
or U168 (N_168,N_148,In_96);
nand U169 (N_169,In_63,N_80);
and U170 (N_170,In_281,In_428);
nand U171 (N_171,In_124,In_337);
nor U172 (N_172,In_123,In_183);
nor U173 (N_173,N_59,In_99);
xnor U174 (N_174,In_125,In_490);
or U175 (N_175,In_70,In_136);
xor U176 (N_176,In_203,In_153);
nor U177 (N_177,N_38,N_8);
nand U178 (N_178,In_405,In_134);
nand U179 (N_179,In_393,In_294);
and U180 (N_180,In_0,N_100);
and U181 (N_181,In_201,N_108);
and U182 (N_182,In_341,N_53);
nor U183 (N_183,In_338,N_39);
xnor U184 (N_184,In_479,In_327);
and U185 (N_185,N_24,In_231);
nand U186 (N_186,N_141,N_94);
nand U187 (N_187,In_49,In_40);
and U188 (N_188,In_190,N_93);
nor U189 (N_189,In_403,N_135);
nand U190 (N_190,N_75,In_380);
nand U191 (N_191,In_206,In_287);
nand U192 (N_192,In_323,N_143);
nand U193 (N_193,N_109,In_222);
and U194 (N_194,In_434,N_92);
and U195 (N_195,In_493,In_109);
and U196 (N_196,In_311,In_181);
or U197 (N_197,In_197,N_65);
and U198 (N_198,In_358,In_5);
nor U199 (N_199,N_146,N_101);
and U200 (N_200,In_35,In_52);
nor U201 (N_201,N_78,In_71);
and U202 (N_202,N_107,In_371);
xnor U203 (N_203,In_271,In_83);
xor U204 (N_204,N_60,N_82);
nand U205 (N_205,N_31,In_391);
nor U206 (N_206,In_260,In_462);
nand U207 (N_207,In_361,N_0);
xor U208 (N_208,In_6,In_458);
nand U209 (N_209,In_115,In_447);
nand U210 (N_210,N_43,In_414);
nor U211 (N_211,N_105,In_470);
and U212 (N_212,In_233,N_5);
nor U213 (N_213,In_416,In_343);
xnor U214 (N_214,In_316,In_285);
or U215 (N_215,N_96,N_136);
or U216 (N_216,In_218,N_129);
nand U217 (N_217,In_354,In_290);
or U218 (N_218,In_151,In_315);
xor U219 (N_219,N_118,In_385);
or U220 (N_220,In_184,In_389);
nor U221 (N_221,In_224,N_79);
and U222 (N_222,In_257,N_7);
nand U223 (N_223,N_103,In_226);
or U224 (N_224,N_20,In_392);
xnor U225 (N_225,N_218,In_36);
xor U226 (N_226,N_172,N_144);
nand U227 (N_227,In_13,In_305);
nor U228 (N_228,In_432,In_274);
nand U229 (N_229,N_202,In_171);
and U230 (N_230,N_188,In_283);
nand U231 (N_231,In_277,N_95);
nor U232 (N_232,N_74,In_313);
or U233 (N_233,In_72,N_142);
and U234 (N_234,N_183,N_187);
and U235 (N_235,In_19,N_199);
nor U236 (N_236,In_423,N_114);
nor U237 (N_237,In_437,N_157);
nand U238 (N_238,N_215,N_174);
nor U239 (N_239,In_413,N_123);
nor U240 (N_240,N_81,N_154);
nor U241 (N_241,N_84,N_132);
or U242 (N_242,N_71,N_195);
xnor U243 (N_243,N_89,N_152);
and U244 (N_244,In_356,N_73);
and U245 (N_245,In_10,In_310);
nor U246 (N_246,N_219,In_150);
nand U247 (N_247,In_266,In_53);
nand U248 (N_248,In_91,In_259);
nor U249 (N_249,In_187,In_420);
nand U250 (N_250,N_46,N_37);
nand U251 (N_251,N_15,In_223);
xor U252 (N_252,In_74,N_221);
xnor U253 (N_253,In_76,N_116);
xor U254 (N_254,In_180,In_195);
or U255 (N_255,In_369,In_289);
xor U256 (N_256,In_112,In_406);
and U257 (N_257,In_127,In_142);
or U258 (N_258,N_192,N_160);
nor U259 (N_259,N_49,In_397);
xor U260 (N_260,N_201,N_189);
xnor U261 (N_261,N_159,N_167);
or U262 (N_262,N_171,In_418);
nor U263 (N_263,N_176,N_115);
and U264 (N_264,N_137,In_177);
or U265 (N_265,In_342,N_217);
nor U266 (N_266,N_170,N_168);
nor U267 (N_267,N_97,N_147);
nand U268 (N_268,In_161,In_116);
nand U269 (N_269,In_346,In_228);
xor U270 (N_270,N_163,N_13);
nand U271 (N_271,In_425,In_426);
xor U272 (N_272,N_98,In_482);
or U273 (N_273,In_75,N_166);
nor U274 (N_274,N_182,In_24);
or U275 (N_275,N_208,In_377);
and U276 (N_276,N_151,N_169);
xor U277 (N_277,In_344,N_198);
and U278 (N_278,In_402,N_178);
nand U279 (N_279,N_220,N_161);
nor U280 (N_280,N_99,In_111);
or U281 (N_281,In_14,In_148);
or U282 (N_282,N_158,In_258);
and U283 (N_283,In_475,N_130);
and U284 (N_284,N_126,N_145);
nand U285 (N_285,N_77,N_204);
or U286 (N_286,N_85,In_118);
xor U287 (N_287,In_229,N_139);
nand U288 (N_288,N_121,N_16);
and U289 (N_289,In_494,N_124);
or U290 (N_290,In_264,In_88);
and U291 (N_291,N_140,N_102);
xor U292 (N_292,N_197,In_336);
xnor U293 (N_293,N_191,N_214);
or U294 (N_294,In_119,In_146);
xnor U295 (N_295,In_68,N_200);
and U296 (N_296,In_314,N_23);
xnor U297 (N_297,N_153,In_399);
xnor U298 (N_298,N_131,In_21);
or U299 (N_299,In_176,N_155);
nor U300 (N_300,N_117,N_273);
nor U301 (N_301,N_284,In_443);
nand U302 (N_302,N_241,N_88);
nand U303 (N_303,N_186,In_61);
nor U304 (N_304,N_229,N_275);
nand U305 (N_305,N_83,N_235);
xnor U306 (N_306,N_180,In_12);
nor U307 (N_307,In_394,N_287);
nand U308 (N_308,N_207,In_262);
or U309 (N_309,N_211,N_213);
xor U310 (N_310,In_357,N_110);
or U311 (N_311,N_280,N_133);
and U312 (N_312,In_97,N_251);
nor U313 (N_313,In_295,N_128);
nor U314 (N_314,In_367,In_243);
nor U315 (N_315,In_4,In_398);
and U316 (N_316,N_291,N_203);
nand U317 (N_317,N_249,N_278);
or U318 (N_318,N_156,N_240);
nor U319 (N_319,N_58,N_272);
nor U320 (N_320,In_459,N_266);
nor U321 (N_321,In_47,N_106);
or U322 (N_322,In_329,N_21);
xor U323 (N_323,N_245,N_276);
nor U324 (N_324,In_139,N_283);
nor U325 (N_325,N_234,N_57);
xnor U326 (N_326,N_120,N_233);
or U327 (N_327,N_242,N_270);
and U328 (N_328,In_93,N_122);
xor U329 (N_329,N_288,In_272);
nor U330 (N_330,N_193,N_205);
or U331 (N_331,In_448,N_209);
or U332 (N_332,In_110,In_383);
nand U333 (N_333,N_250,N_63);
xor U334 (N_334,In_396,N_232);
nor U335 (N_335,In_492,N_90);
or U336 (N_336,N_150,In_185);
nor U337 (N_337,N_225,N_184);
xnor U338 (N_338,N_299,In_219);
nor U339 (N_339,In_308,N_293);
nand U340 (N_340,In_129,N_262);
and U341 (N_341,N_12,In_66);
xnor U342 (N_342,N_54,N_44);
or U343 (N_343,In_454,N_263);
nand U344 (N_344,In_366,N_259);
and U345 (N_345,In_241,In_352);
nor U346 (N_346,N_274,In_28);
xor U347 (N_347,N_292,In_172);
nor U348 (N_348,N_164,In_114);
nor U349 (N_349,In_200,In_86);
nor U350 (N_350,In_441,N_285);
xnor U351 (N_351,In_491,In_451);
and U352 (N_352,N_224,N_212);
and U353 (N_353,N_134,In_232);
nand U354 (N_354,N_223,In_45);
and U355 (N_355,In_193,N_228);
nor U356 (N_356,N_260,N_279);
nor U357 (N_357,N_295,N_289);
nand U358 (N_358,N_25,N_237);
nand U359 (N_359,N_255,N_296);
or U360 (N_360,In_444,N_286);
xor U361 (N_361,N_254,N_35);
or U362 (N_362,In_293,In_25);
or U363 (N_363,N_256,N_206);
or U364 (N_364,In_429,N_294);
and U365 (N_365,N_32,N_222);
and U366 (N_366,N_111,N_227);
xnor U367 (N_367,In_22,In_191);
xor U368 (N_368,In_135,In_78);
nand U369 (N_369,N_190,N_210);
and U370 (N_370,N_265,N_179);
xnor U371 (N_371,N_86,N_162);
or U372 (N_372,N_257,N_196);
or U373 (N_373,In_82,N_91);
nor U374 (N_374,N_127,In_133);
xor U375 (N_375,N_247,N_177);
xnor U376 (N_376,N_119,N_309);
and U377 (N_377,N_366,N_243);
and U378 (N_378,N_267,N_352);
xor U379 (N_379,N_48,N_301);
or U380 (N_380,N_324,N_304);
or U381 (N_381,N_353,N_239);
or U382 (N_382,N_216,N_349);
xnor U383 (N_383,N_315,N_335);
or U384 (N_384,N_328,N_277);
nor U385 (N_385,N_230,N_369);
and U386 (N_386,N_361,N_264);
and U387 (N_387,N_319,N_317);
nand U388 (N_388,N_314,N_175);
xor U389 (N_389,N_181,N_11);
nor U390 (N_390,N_350,N_246);
or U391 (N_391,N_370,N_318);
nor U392 (N_392,N_332,N_261);
xnor U393 (N_393,N_358,N_357);
or U394 (N_394,In_445,N_185);
or U395 (N_395,N_343,In_87);
nor U396 (N_396,In_485,N_252);
or U397 (N_397,N_320,N_316);
nand U398 (N_398,N_321,N_347);
or U399 (N_399,N_281,In_484);
nand U400 (N_400,N_322,N_297);
nor U401 (N_401,N_248,N_342);
nand U402 (N_402,In_278,N_329);
and U403 (N_403,N_194,N_268);
or U404 (N_404,N_330,N_308);
xor U405 (N_405,N_345,In_205);
nand U406 (N_406,N_298,N_373);
or U407 (N_407,N_368,N_338);
or U408 (N_408,N_302,N_165);
nand U409 (N_409,In_230,N_326);
xnor U410 (N_410,N_337,N_364);
xor U411 (N_411,N_341,N_362);
nor U412 (N_412,N_173,N_236);
nand U413 (N_413,N_253,N_14);
and U414 (N_414,N_344,N_339);
nand U415 (N_415,N_300,In_410);
nand U416 (N_416,N_312,N_244);
nor U417 (N_417,N_327,N_372);
or U418 (N_418,N_371,N_269);
and U419 (N_419,N_56,N_374);
or U420 (N_420,N_354,N_238);
xnor U421 (N_421,N_290,N_355);
and U422 (N_422,N_313,N_282);
and U423 (N_423,N_303,N_258);
nor U424 (N_424,N_359,N_331);
xor U425 (N_425,N_346,N_311);
xor U426 (N_426,N_325,N_10);
nor U427 (N_427,N_351,N_310);
nand U428 (N_428,N_365,N_367);
and U429 (N_429,N_363,N_231);
nand U430 (N_430,In_252,N_356);
nand U431 (N_431,N_334,N_306);
nand U432 (N_432,N_271,N_323);
nor U433 (N_433,N_333,N_307);
and U434 (N_434,N_360,N_336);
nor U435 (N_435,N_340,In_339);
nand U436 (N_436,N_226,N_348);
xor U437 (N_437,N_305,N_366);
nand U438 (N_438,N_175,N_239);
nand U439 (N_439,N_48,N_303);
nand U440 (N_440,N_365,N_56);
nor U441 (N_441,N_365,N_303);
and U442 (N_442,N_282,N_356);
nand U443 (N_443,N_181,N_194);
nand U444 (N_444,N_194,N_332);
nand U445 (N_445,In_205,In_87);
nand U446 (N_446,N_247,N_338);
and U447 (N_447,N_277,N_319);
xor U448 (N_448,N_359,N_313);
and U449 (N_449,N_340,N_252);
nor U450 (N_450,N_377,N_444);
nor U451 (N_451,N_413,N_448);
nor U452 (N_452,N_418,N_386);
and U453 (N_453,N_405,N_383);
nand U454 (N_454,N_387,N_396);
nor U455 (N_455,N_378,N_408);
xnor U456 (N_456,N_390,N_423);
xnor U457 (N_457,N_394,N_401);
nand U458 (N_458,N_449,N_389);
and U459 (N_459,N_422,N_384);
xor U460 (N_460,N_425,N_417);
and U461 (N_461,N_379,N_400);
nand U462 (N_462,N_380,N_437);
and U463 (N_463,N_414,N_443);
nand U464 (N_464,N_430,N_436);
xnor U465 (N_465,N_398,N_428);
and U466 (N_466,N_438,N_375);
or U467 (N_467,N_431,N_433);
and U468 (N_468,N_420,N_381);
nor U469 (N_469,N_446,N_397);
and U470 (N_470,N_391,N_395);
nand U471 (N_471,N_424,N_382);
or U472 (N_472,N_415,N_392);
or U473 (N_473,N_412,N_439);
and U474 (N_474,N_407,N_404);
and U475 (N_475,N_435,N_406);
nand U476 (N_476,N_421,N_441);
nand U477 (N_477,N_416,N_427);
nand U478 (N_478,N_388,N_429);
xor U479 (N_479,N_376,N_411);
or U480 (N_480,N_399,N_409);
and U481 (N_481,N_410,N_426);
nand U482 (N_482,N_442,N_445);
nand U483 (N_483,N_432,N_419);
and U484 (N_484,N_440,N_447);
and U485 (N_485,N_393,N_385);
xnor U486 (N_486,N_402,N_403);
or U487 (N_487,N_434,N_403);
and U488 (N_488,N_446,N_398);
nor U489 (N_489,N_419,N_378);
or U490 (N_490,N_445,N_446);
xnor U491 (N_491,N_448,N_382);
xor U492 (N_492,N_390,N_424);
nor U493 (N_493,N_378,N_406);
xnor U494 (N_494,N_443,N_437);
or U495 (N_495,N_430,N_419);
nand U496 (N_496,N_433,N_399);
or U497 (N_497,N_408,N_445);
nand U498 (N_498,N_411,N_416);
xnor U499 (N_499,N_436,N_442);
or U500 (N_500,N_430,N_409);
nand U501 (N_501,N_426,N_389);
and U502 (N_502,N_417,N_398);
nand U503 (N_503,N_427,N_426);
xnor U504 (N_504,N_381,N_407);
nor U505 (N_505,N_423,N_421);
nand U506 (N_506,N_443,N_448);
or U507 (N_507,N_434,N_415);
nand U508 (N_508,N_443,N_384);
and U509 (N_509,N_401,N_410);
and U510 (N_510,N_387,N_382);
nor U511 (N_511,N_439,N_418);
and U512 (N_512,N_443,N_420);
nand U513 (N_513,N_440,N_381);
or U514 (N_514,N_380,N_424);
xor U515 (N_515,N_425,N_422);
nor U516 (N_516,N_403,N_395);
or U517 (N_517,N_440,N_408);
xor U518 (N_518,N_399,N_445);
nand U519 (N_519,N_386,N_445);
nand U520 (N_520,N_422,N_391);
xor U521 (N_521,N_443,N_408);
xnor U522 (N_522,N_428,N_425);
and U523 (N_523,N_415,N_420);
nand U524 (N_524,N_446,N_378);
nor U525 (N_525,N_504,N_512);
and U526 (N_526,N_523,N_501);
and U527 (N_527,N_496,N_491);
nor U528 (N_528,N_484,N_509);
nor U529 (N_529,N_461,N_522);
nand U530 (N_530,N_495,N_455);
nor U531 (N_531,N_459,N_465);
nor U532 (N_532,N_451,N_481);
nand U533 (N_533,N_499,N_500);
nand U534 (N_534,N_468,N_524);
xnor U535 (N_535,N_490,N_489);
nor U536 (N_536,N_485,N_514);
nor U537 (N_537,N_497,N_466);
nand U538 (N_538,N_510,N_478);
nand U539 (N_539,N_507,N_520);
xor U540 (N_540,N_483,N_521);
nor U541 (N_541,N_480,N_513);
nor U542 (N_542,N_457,N_511);
and U543 (N_543,N_498,N_488);
nor U544 (N_544,N_476,N_469);
and U545 (N_545,N_515,N_492);
or U546 (N_546,N_453,N_486);
and U547 (N_547,N_450,N_487);
nand U548 (N_548,N_518,N_505);
nand U549 (N_549,N_460,N_517);
and U550 (N_550,N_473,N_456);
and U551 (N_551,N_479,N_472);
and U552 (N_552,N_519,N_470);
or U553 (N_553,N_493,N_516);
xor U554 (N_554,N_502,N_506);
nor U555 (N_555,N_462,N_508);
or U556 (N_556,N_454,N_474);
nor U557 (N_557,N_503,N_458);
nor U558 (N_558,N_467,N_463);
nand U559 (N_559,N_482,N_471);
nand U560 (N_560,N_475,N_464);
and U561 (N_561,N_494,N_477);
xor U562 (N_562,N_452,N_465);
nor U563 (N_563,N_523,N_471);
nand U564 (N_564,N_462,N_505);
nor U565 (N_565,N_481,N_470);
nor U566 (N_566,N_512,N_451);
xor U567 (N_567,N_496,N_468);
or U568 (N_568,N_490,N_504);
nor U569 (N_569,N_477,N_456);
nand U570 (N_570,N_451,N_488);
and U571 (N_571,N_467,N_506);
xor U572 (N_572,N_469,N_492);
nor U573 (N_573,N_478,N_518);
nor U574 (N_574,N_515,N_524);
nor U575 (N_575,N_519,N_473);
nor U576 (N_576,N_465,N_480);
xor U577 (N_577,N_522,N_484);
nand U578 (N_578,N_524,N_517);
and U579 (N_579,N_483,N_475);
nand U580 (N_580,N_466,N_502);
and U581 (N_581,N_512,N_489);
nor U582 (N_582,N_498,N_452);
xor U583 (N_583,N_459,N_506);
nand U584 (N_584,N_497,N_501);
xor U585 (N_585,N_514,N_451);
or U586 (N_586,N_500,N_466);
xor U587 (N_587,N_486,N_454);
xor U588 (N_588,N_452,N_483);
and U589 (N_589,N_457,N_505);
or U590 (N_590,N_490,N_520);
xor U591 (N_591,N_522,N_485);
or U592 (N_592,N_500,N_507);
xnor U593 (N_593,N_507,N_471);
and U594 (N_594,N_456,N_493);
and U595 (N_595,N_494,N_478);
nand U596 (N_596,N_450,N_482);
or U597 (N_597,N_493,N_517);
nor U598 (N_598,N_472,N_450);
nand U599 (N_599,N_513,N_507);
or U600 (N_600,N_577,N_588);
nor U601 (N_601,N_589,N_543);
and U602 (N_602,N_591,N_548);
and U603 (N_603,N_535,N_586);
xor U604 (N_604,N_595,N_538);
or U605 (N_605,N_561,N_539);
and U606 (N_606,N_550,N_558);
xnor U607 (N_607,N_582,N_542);
and U608 (N_608,N_578,N_576);
or U609 (N_609,N_583,N_555);
and U610 (N_610,N_547,N_566);
nor U611 (N_611,N_537,N_534);
nand U612 (N_612,N_545,N_584);
or U613 (N_613,N_528,N_557);
nand U614 (N_614,N_570,N_574);
or U615 (N_615,N_530,N_556);
nand U616 (N_616,N_569,N_594);
or U617 (N_617,N_533,N_568);
nor U618 (N_618,N_532,N_549);
or U619 (N_619,N_585,N_529);
xor U620 (N_620,N_575,N_579);
and U621 (N_621,N_599,N_564);
nand U622 (N_622,N_559,N_525);
nor U623 (N_623,N_536,N_590);
nand U624 (N_624,N_563,N_531);
xor U625 (N_625,N_544,N_541);
xnor U626 (N_626,N_598,N_554);
xnor U627 (N_627,N_540,N_573);
nand U628 (N_628,N_565,N_571);
xnor U629 (N_629,N_527,N_562);
and U630 (N_630,N_597,N_592);
or U631 (N_631,N_572,N_581);
and U632 (N_632,N_551,N_553);
xor U633 (N_633,N_593,N_546);
and U634 (N_634,N_587,N_526);
nand U635 (N_635,N_560,N_552);
nand U636 (N_636,N_580,N_596);
xor U637 (N_637,N_567,N_582);
or U638 (N_638,N_581,N_561);
nor U639 (N_639,N_595,N_583);
and U640 (N_640,N_554,N_592);
or U641 (N_641,N_579,N_588);
nor U642 (N_642,N_575,N_545);
nand U643 (N_643,N_564,N_561);
and U644 (N_644,N_584,N_525);
nand U645 (N_645,N_526,N_564);
and U646 (N_646,N_575,N_558);
nor U647 (N_647,N_555,N_532);
or U648 (N_648,N_547,N_564);
or U649 (N_649,N_577,N_546);
and U650 (N_650,N_589,N_591);
nor U651 (N_651,N_593,N_548);
xnor U652 (N_652,N_554,N_588);
xor U653 (N_653,N_555,N_574);
xnor U654 (N_654,N_555,N_557);
xor U655 (N_655,N_574,N_571);
nand U656 (N_656,N_556,N_570);
nand U657 (N_657,N_594,N_540);
nand U658 (N_658,N_573,N_584);
xnor U659 (N_659,N_535,N_553);
or U660 (N_660,N_536,N_531);
xnor U661 (N_661,N_565,N_568);
nor U662 (N_662,N_571,N_529);
xnor U663 (N_663,N_543,N_557);
nand U664 (N_664,N_599,N_578);
or U665 (N_665,N_597,N_582);
nand U666 (N_666,N_534,N_558);
nand U667 (N_667,N_586,N_594);
and U668 (N_668,N_543,N_563);
nand U669 (N_669,N_599,N_533);
nand U670 (N_670,N_553,N_579);
or U671 (N_671,N_554,N_595);
or U672 (N_672,N_579,N_537);
nand U673 (N_673,N_568,N_548);
xnor U674 (N_674,N_589,N_564);
xor U675 (N_675,N_670,N_651);
xnor U676 (N_676,N_601,N_669);
nor U677 (N_677,N_613,N_635);
nand U678 (N_678,N_649,N_625);
xor U679 (N_679,N_622,N_671);
and U680 (N_680,N_602,N_659);
xor U681 (N_681,N_606,N_662);
or U682 (N_682,N_638,N_639);
and U683 (N_683,N_643,N_605);
and U684 (N_684,N_656,N_661);
xnor U685 (N_685,N_623,N_645);
nand U686 (N_686,N_652,N_648);
xnor U687 (N_687,N_673,N_636);
xor U688 (N_688,N_658,N_627);
or U689 (N_689,N_620,N_668);
and U690 (N_690,N_609,N_674);
and U691 (N_691,N_672,N_621);
or U692 (N_692,N_603,N_604);
xor U693 (N_693,N_647,N_626);
xor U694 (N_694,N_650,N_615);
nand U695 (N_695,N_663,N_667);
nand U696 (N_696,N_644,N_631);
or U697 (N_697,N_628,N_629);
nand U698 (N_698,N_634,N_611);
xor U699 (N_699,N_632,N_633);
or U700 (N_700,N_654,N_630);
nor U701 (N_701,N_610,N_655);
xnor U702 (N_702,N_657,N_624);
xnor U703 (N_703,N_607,N_640);
xor U704 (N_704,N_664,N_646);
and U705 (N_705,N_653,N_642);
nor U706 (N_706,N_660,N_612);
nand U707 (N_707,N_618,N_666);
or U708 (N_708,N_619,N_641);
and U709 (N_709,N_637,N_617);
nor U710 (N_710,N_600,N_665);
or U711 (N_711,N_608,N_616);
and U712 (N_712,N_614,N_610);
nand U713 (N_713,N_661,N_611);
or U714 (N_714,N_634,N_654);
or U715 (N_715,N_624,N_651);
nand U716 (N_716,N_618,N_625);
or U717 (N_717,N_646,N_665);
xor U718 (N_718,N_617,N_616);
nor U719 (N_719,N_635,N_661);
or U720 (N_720,N_605,N_651);
and U721 (N_721,N_664,N_667);
and U722 (N_722,N_619,N_636);
or U723 (N_723,N_629,N_606);
and U724 (N_724,N_607,N_616);
or U725 (N_725,N_616,N_614);
xor U726 (N_726,N_652,N_631);
or U727 (N_727,N_636,N_662);
and U728 (N_728,N_628,N_640);
xor U729 (N_729,N_609,N_658);
or U730 (N_730,N_654,N_629);
or U731 (N_731,N_668,N_669);
nor U732 (N_732,N_611,N_619);
nand U733 (N_733,N_612,N_644);
xnor U734 (N_734,N_658,N_662);
nand U735 (N_735,N_668,N_621);
xnor U736 (N_736,N_609,N_635);
and U737 (N_737,N_638,N_622);
xor U738 (N_738,N_650,N_622);
nor U739 (N_739,N_627,N_648);
or U740 (N_740,N_603,N_643);
xnor U741 (N_741,N_615,N_629);
and U742 (N_742,N_620,N_625);
xor U743 (N_743,N_614,N_635);
and U744 (N_744,N_633,N_612);
and U745 (N_745,N_655,N_669);
and U746 (N_746,N_666,N_624);
nor U747 (N_747,N_649,N_628);
xnor U748 (N_748,N_627,N_616);
nor U749 (N_749,N_661,N_673);
nand U750 (N_750,N_726,N_708);
nand U751 (N_751,N_709,N_696);
nor U752 (N_752,N_688,N_680);
and U753 (N_753,N_701,N_697);
nor U754 (N_754,N_719,N_715);
nor U755 (N_755,N_690,N_732);
or U756 (N_756,N_702,N_728);
nor U757 (N_757,N_699,N_687);
or U758 (N_758,N_675,N_738);
nor U759 (N_759,N_717,N_743);
xor U760 (N_760,N_716,N_722);
and U761 (N_761,N_689,N_734);
and U762 (N_762,N_693,N_706);
nand U763 (N_763,N_721,N_749);
nor U764 (N_764,N_703,N_686);
or U765 (N_765,N_746,N_705);
xnor U766 (N_766,N_678,N_730);
and U767 (N_767,N_679,N_745);
xnor U768 (N_768,N_739,N_698);
nor U769 (N_769,N_714,N_741);
nor U770 (N_770,N_684,N_718);
or U771 (N_771,N_692,N_731);
nand U772 (N_772,N_724,N_744);
nor U773 (N_773,N_713,N_707);
and U774 (N_774,N_683,N_723);
or U775 (N_775,N_681,N_682);
nor U776 (N_776,N_695,N_694);
nand U777 (N_777,N_742,N_735);
or U778 (N_778,N_748,N_736);
or U779 (N_779,N_710,N_685);
xnor U780 (N_780,N_740,N_737);
nand U781 (N_781,N_727,N_725);
and U782 (N_782,N_677,N_712);
xor U783 (N_783,N_720,N_691);
xnor U784 (N_784,N_747,N_733);
nand U785 (N_785,N_676,N_711);
nand U786 (N_786,N_700,N_704);
xnor U787 (N_787,N_729,N_717);
or U788 (N_788,N_747,N_694);
or U789 (N_789,N_700,N_699);
xor U790 (N_790,N_686,N_700);
nor U791 (N_791,N_679,N_738);
nand U792 (N_792,N_740,N_713);
nor U793 (N_793,N_675,N_710);
nor U794 (N_794,N_742,N_745);
or U795 (N_795,N_725,N_693);
nand U796 (N_796,N_686,N_708);
or U797 (N_797,N_711,N_742);
nand U798 (N_798,N_740,N_733);
nand U799 (N_799,N_714,N_716);
nand U800 (N_800,N_709,N_690);
xor U801 (N_801,N_702,N_746);
or U802 (N_802,N_744,N_694);
nor U803 (N_803,N_733,N_743);
or U804 (N_804,N_721,N_709);
nand U805 (N_805,N_745,N_733);
or U806 (N_806,N_692,N_719);
or U807 (N_807,N_700,N_721);
xnor U808 (N_808,N_714,N_743);
or U809 (N_809,N_720,N_690);
and U810 (N_810,N_710,N_712);
xor U811 (N_811,N_694,N_729);
and U812 (N_812,N_707,N_697);
and U813 (N_813,N_717,N_675);
nand U814 (N_814,N_724,N_746);
or U815 (N_815,N_703,N_725);
nor U816 (N_816,N_727,N_724);
nand U817 (N_817,N_697,N_696);
or U818 (N_818,N_693,N_729);
xor U819 (N_819,N_742,N_724);
xnor U820 (N_820,N_718,N_685);
nor U821 (N_821,N_720,N_717);
nand U822 (N_822,N_728,N_741);
xor U823 (N_823,N_693,N_728);
nor U824 (N_824,N_717,N_725);
and U825 (N_825,N_791,N_783);
and U826 (N_826,N_811,N_792);
xnor U827 (N_827,N_807,N_780);
or U828 (N_828,N_804,N_757);
nor U829 (N_829,N_789,N_771);
xor U830 (N_830,N_751,N_755);
and U831 (N_831,N_761,N_822);
xor U832 (N_832,N_754,N_794);
or U833 (N_833,N_803,N_798);
nor U834 (N_834,N_784,N_782);
xnor U835 (N_835,N_753,N_816);
nor U836 (N_836,N_764,N_775);
and U837 (N_837,N_820,N_772);
nor U838 (N_838,N_815,N_809);
or U839 (N_839,N_770,N_800);
nand U840 (N_840,N_752,N_769);
nand U841 (N_841,N_812,N_808);
and U842 (N_842,N_786,N_773);
nand U843 (N_843,N_790,N_787);
xnor U844 (N_844,N_806,N_767);
nor U845 (N_845,N_817,N_759);
and U846 (N_846,N_750,N_796);
or U847 (N_847,N_768,N_760);
xor U848 (N_848,N_801,N_793);
nor U849 (N_849,N_823,N_785);
and U850 (N_850,N_821,N_776);
or U851 (N_851,N_818,N_779);
or U852 (N_852,N_795,N_765);
xor U853 (N_853,N_788,N_756);
xnor U854 (N_854,N_762,N_758);
nand U855 (N_855,N_763,N_777);
or U856 (N_856,N_813,N_778);
or U857 (N_857,N_805,N_781);
xor U858 (N_858,N_819,N_766);
and U859 (N_859,N_774,N_810);
nand U860 (N_860,N_814,N_824);
or U861 (N_861,N_799,N_802);
nand U862 (N_862,N_797,N_776);
nand U863 (N_863,N_810,N_757);
and U864 (N_864,N_768,N_800);
and U865 (N_865,N_798,N_780);
nor U866 (N_866,N_794,N_812);
nor U867 (N_867,N_824,N_800);
nor U868 (N_868,N_765,N_823);
xnor U869 (N_869,N_768,N_817);
nor U870 (N_870,N_807,N_812);
xnor U871 (N_871,N_818,N_796);
nor U872 (N_872,N_757,N_800);
or U873 (N_873,N_755,N_811);
or U874 (N_874,N_750,N_794);
nand U875 (N_875,N_781,N_763);
or U876 (N_876,N_750,N_783);
xnor U877 (N_877,N_761,N_805);
nor U878 (N_878,N_774,N_752);
nor U879 (N_879,N_756,N_755);
or U880 (N_880,N_765,N_790);
xnor U881 (N_881,N_789,N_768);
xnor U882 (N_882,N_762,N_796);
nor U883 (N_883,N_754,N_803);
nand U884 (N_884,N_815,N_756);
or U885 (N_885,N_782,N_754);
xnor U886 (N_886,N_756,N_753);
or U887 (N_887,N_784,N_761);
nand U888 (N_888,N_812,N_781);
nand U889 (N_889,N_798,N_755);
or U890 (N_890,N_764,N_789);
xnor U891 (N_891,N_769,N_798);
and U892 (N_892,N_805,N_786);
or U893 (N_893,N_772,N_777);
nand U894 (N_894,N_792,N_783);
and U895 (N_895,N_821,N_808);
nand U896 (N_896,N_775,N_782);
xor U897 (N_897,N_823,N_781);
or U898 (N_898,N_804,N_814);
and U899 (N_899,N_801,N_812);
nor U900 (N_900,N_888,N_878);
xor U901 (N_901,N_861,N_869);
or U902 (N_902,N_879,N_865);
nand U903 (N_903,N_877,N_844);
and U904 (N_904,N_871,N_847);
and U905 (N_905,N_863,N_860);
nand U906 (N_906,N_825,N_842);
or U907 (N_907,N_854,N_899);
xor U908 (N_908,N_889,N_866);
or U909 (N_909,N_830,N_887);
xor U910 (N_910,N_839,N_835);
and U911 (N_911,N_848,N_841);
xor U912 (N_912,N_853,N_850);
and U913 (N_913,N_864,N_827);
nor U914 (N_914,N_834,N_891);
or U915 (N_915,N_894,N_831);
nor U916 (N_916,N_884,N_870);
and U917 (N_917,N_858,N_897);
nand U918 (N_918,N_880,N_836);
xnor U919 (N_919,N_837,N_845);
xnor U920 (N_920,N_859,N_849);
nand U921 (N_921,N_895,N_893);
or U922 (N_922,N_867,N_851);
nand U923 (N_923,N_882,N_868);
xor U924 (N_924,N_846,N_881);
nor U925 (N_925,N_856,N_857);
or U926 (N_926,N_873,N_892);
and U927 (N_927,N_829,N_828);
nand U928 (N_928,N_843,N_886);
xnor U929 (N_929,N_876,N_852);
nor U930 (N_930,N_872,N_875);
or U931 (N_931,N_898,N_838);
nor U932 (N_932,N_826,N_885);
or U933 (N_933,N_874,N_855);
or U934 (N_934,N_832,N_840);
or U935 (N_935,N_833,N_883);
or U936 (N_936,N_896,N_890);
nor U937 (N_937,N_862,N_890);
xnor U938 (N_938,N_849,N_845);
and U939 (N_939,N_826,N_889);
or U940 (N_940,N_839,N_888);
nand U941 (N_941,N_895,N_838);
and U942 (N_942,N_868,N_846);
and U943 (N_943,N_875,N_869);
nand U944 (N_944,N_829,N_838);
xor U945 (N_945,N_879,N_843);
or U946 (N_946,N_861,N_891);
and U947 (N_947,N_897,N_841);
xnor U948 (N_948,N_835,N_874);
nor U949 (N_949,N_864,N_870);
or U950 (N_950,N_836,N_844);
and U951 (N_951,N_867,N_874);
or U952 (N_952,N_877,N_880);
or U953 (N_953,N_855,N_889);
xnor U954 (N_954,N_867,N_831);
nor U955 (N_955,N_861,N_883);
or U956 (N_956,N_874,N_881);
and U957 (N_957,N_836,N_835);
and U958 (N_958,N_893,N_878);
nand U959 (N_959,N_855,N_890);
nand U960 (N_960,N_863,N_898);
or U961 (N_961,N_880,N_864);
nand U962 (N_962,N_868,N_858);
nor U963 (N_963,N_826,N_875);
nor U964 (N_964,N_860,N_830);
or U965 (N_965,N_884,N_846);
or U966 (N_966,N_891,N_897);
nor U967 (N_967,N_861,N_857);
and U968 (N_968,N_898,N_895);
or U969 (N_969,N_892,N_889);
nor U970 (N_970,N_868,N_879);
or U971 (N_971,N_894,N_830);
or U972 (N_972,N_889,N_878);
or U973 (N_973,N_872,N_835);
and U974 (N_974,N_857,N_855);
and U975 (N_975,N_918,N_957);
and U976 (N_976,N_917,N_949);
nand U977 (N_977,N_970,N_972);
or U978 (N_978,N_915,N_919);
and U979 (N_979,N_901,N_902);
or U980 (N_980,N_967,N_951);
or U981 (N_981,N_956,N_927);
and U982 (N_982,N_920,N_905);
xnor U983 (N_983,N_925,N_963);
nor U984 (N_984,N_935,N_955);
xor U985 (N_985,N_947,N_952);
and U986 (N_986,N_929,N_926);
and U987 (N_987,N_959,N_912);
and U988 (N_988,N_913,N_936);
xor U989 (N_989,N_974,N_940);
or U990 (N_990,N_934,N_916);
nand U991 (N_991,N_944,N_907);
nand U992 (N_992,N_923,N_938);
and U993 (N_993,N_969,N_962);
nor U994 (N_994,N_906,N_954);
nand U995 (N_995,N_900,N_928);
or U996 (N_996,N_904,N_922);
nand U997 (N_997,N_958,N_941);
and U998 (N_998,N_937,N_914);
nand U999 (N_999,N_964,N_961);
nor U1000 (N_1000,N_911,N_943);
nor U1001 (N_1001,N_939,N_971);
nand U1002 (N_1002,N_908,N_924);
xnor U1003 (N_1003,N_960,N_950);
xnor U1004 (N_1004,N_965,N_903);
or U1005 (N_1005,N_910,N_933);
or U1006 (N_1006,N_945,N_973);
xnor U1007 (N_1007,N_931,N_966);
xor U1008 (N_1008,N_909,N_968);
or U1009 (N_1009,N_921,N_942);
xnor U1010 (N_1010,N_932,N_930);
or U1011 (N_1011,N_953,N_948);
nand U1012 (N_1012,N_946,N_929);
and U1013 (N_1013,N_912,N_960);
or U1014 (N_1014,N_968,N_965);
nor U1015 (N_1015,N_949,N_954);
xnor U1016 (N_1016,N_963,N_930);
xnor U1017 (N_1017,N_939,N_904);
nor U1018 (N_1018,N_957,N_937);
xnor U1019 (N_1019,N_928,N_961);
or U1020 (N_1020,N_974,N_914);
nor U1021 (N_1021,N_959,N_952);
nand U1022 (N_1022,N_901,N_940);
nor U1023 (N_1023,N_965,N_936);
nand U1024 (N_1024,N_944,N_935);
nor U1025 (N_1025,N_911,N_915);
nor U1026 (N_1026,N_934,N_929);
nand U1027 (N_1027,N_956,N_904);
xor U1028 (N_1028,N_965,N_912);
or U1029 (N_1029,N_948,N_926);
and U1030 (N_1030,N_954,N_920);
or U1031 (N_1031,N_926,N_946);
nand U1032 (N_1032,N_961,N_914);
xnor U1033 (N_1033,N_955,N_934);
or U1034 (N_1034,N_961,N_927);
or U1035 (N_1035,N_956,N_967);
or U1036 (N_1036,N_901,N_922);
or U1037 (N_1037,N_959,N_935);
or U1038 (N_1038,N_917,N_902);
and U1039 (N_1039,N_949,N_907);
or U1040 (N_1040,N_924,N_968);
nor U1041 (N_1041,N_942,N_923);
nor U1042 (N_1042,N_974,N_960);
and U1043 (N_1043,N_908,N_917);
nand U1044 (N_1044,N_967,N_966);
and U1045 (N_1045,N_920,N_913);
xnor U1046 (N_1046,N_957,N_946);
or U1047 (N_1047,N_951,N_914);
and U1048 (N_1048,N_901,N_931);
or U1049 (N_1049,N_920,N_943);
or U1050 (N_1050,N_1016,N_1046);
xnor U1051 (N_1051,N_1031,N_1040);
and U1052 (N_1052,N_997,N_1035);
xor U1053 (N_1053,N_1001,N_1020);
and U1054 (N_1054,N_1023,N_975);
nand U1055 (N_1055,N_991,N_1036);
nand U1056 (N_1056,N_1038,N_1044);
or U1057 (N_1057,N_980,N_1022);
nor U1058 (N_1058,N_1037,N_1039);
xnor U1059 (N_1059,N_990,N_1005);
nand U1060 (N_1060,N_1004,N_1048);
nand U1061 (N_1061,N_977,N_978);
and U1062 (N_1062,N_986,N_1045);
xor U1063 (N_1063,N_1002,N_1029);
or U1064 (N_1064,N_1024,N_1034);
and U1065 (N_1065,N_988,N_1013);
nand U1066 (N_1066,N_1043,N_1028);
nand U1067 (N_1067,N_976,N_1003);
or U1068 (N_1068,N_1021,N_1033);
nor U1069 (N_1069,N_1042,N_989);
nor U1070 (N_1070,N_1019,N_993);
and U1071 (N_1071,N_1049,N_1015);
nor U1072 (N_1072,N_1010,N_1047);
or U1073 (N_1073,N_983,N_999);
or U1074 (N_1074,N_979,N_1041);
nand U1075 (N_1075,N_1006,N_981);
nand U1076 (N_1076,N_1007,N_996);
nand U1077 (N_1077,N_1014,N_1018);
and U1078 (N_1078,N_1011,N_1008);
nand U1079 (N_1079,N_984,N_1025);
or U1080 (N_1080,N_1009,N_995);
nand U1081 (N_1081,N_987,N_998);
and U1082 (N_1082,N_1026,N_985);
xnor U1083 (N_1083,N_1032,N_1000);
and U1084 (N_1084,N_1027,N_982);
and U1085 (N_1085,N_1017,N_992);
nor U1086 (N_1086,N_1030,N_994);
nor U1087 (N_1087,N_1012,N_1026);
nor U1088 (N_1088,N_983,N_988);
xnor U1089 (N_1089,N_1003,N_993);
nor U1090 (N_1090,N_1018,N_1019);
and U1091 (N_1091,N_1043,N_1038);
xor U1092 (N_1092,N_1036,N_1038);
or U1093 (N_1093,N_995,N_1033);
nor U1094 (N_1094,N_1016,N_1012);
or U1095 (N_1095,N_1012,N_1019);
xor U1096 (N_1096,N_992,N_1033);
xnor U1097 (N_1097,N_1007,N_1020);
nor U1098 (N_1098,N_1037,N_992);
xor U1099 (N_1099,N_1023,N_993);
nand U1100 (N_1100,N_1033,N_988);
or U1101 (N_1101,N_1043,N_997);
nand U1102 (N_1102,N_1025,N_998);
nand U1103 (N_1103,N_1027,N_987);
xnor U1104 (N_1104,N_983,N_1025);
nor U1105 (N_1105,N_1047,N_1036);
and U1106 (N_1106,N_980,N_1021);
nand U1107 (N_1107,N_1018,N_1010);
nand U1108 (N_1108,N_1004,N_1021);
xnor U1109 (N_1109,N_1042,N_992);
or U1110 (N_1110,N_1022,N_1006);
or U1111 (N_1111,N_1044,N_983);
nand U1112 (N_1112,N_1033,N_996);
or U1113 (N_1113,N_1026,N_982);
nand U1114 (N_1114,N_997,N_1010);
nand U1115 (N_1115,N_1039,N_1040);
nor U1116 (N_1116,N_1030,N_1049);
or U1117 (N_1117,N_983,N_1024);
or U1118 (N_1118,N_994,N_1020);
nor U1119 (N_1119,N_1045,N_1031);
or U1120 (N_1120,N_983,N_986);
or U1121 (N_1121,N_987,N_997);
nand U1122 (N_1122,N_1011,N_1000);
and U1123 (N_1123,N_1003,N_987);
nor U1124 (N_1124,N_1025,N_1021);
nand U1125 (N_1125,N_1093,N_1075);
xor U1126 (N_1126,N_1120,N_1115);
nand U1127 (N_1127,N_1058,N_1064);
nand U1128 (N_1128,N_1080,N_1091);
xor U1129 (N_1129,N_1116,N_1105);
nand U1130 (N_1130,N_1090,N_1078);
nor U1131 (N_1131,N_1063,N_1103);
and U1132 (N_1132,N_1099,N_1057);
and U1133 (N_1133,N_1104,N_1083);
nor U1134 (N_1134,N_1097,N_1052);
nand U1135 (N_1135,N_1106,N_1107);
and U1136 (N_1136,N_1109,N_1100);
nand U1137 (N_1137,N_1098,N_1101);
or U1138 (N_1138,N_1061,N_1094);
xnor U1139 (N_1139,N_1066,N_1053);
xnor U1140 (N_1140,N_1062,N_1055);
and U1141 (N_1141,N_1081,N_1050);
nor U1142 (N_1142,N_1095,N_1074);
nor U1143 (N_1143,N_1068,N_1110);
xnor U1144 (N_1144,N_1114,N_1102);
nand U1145 (N_1145,N_1112,N_1069);
nand U1146 (N_1146,N_1089,N_1117);
nor U1147 (N_1147,N_1067,N_1056);
nand U1148 (N_1148,N_1060,N_1119);
nor U1149 (N_1149,N_1118,N_1065);
and U1150 (N_1150,N_1084,N_1071);
or U1151 (N_1151,N_1092,N_1079);
nand U1152 (N_1152,N_1124,N_1108);
and U1153 (N_1153,N_1070,N_1077);
and U1154 (N_1154,N_1073,N_1123);
or U1155 (N_1155,N_1086,N_1096);
xor U1156 (N_1156,N_1085,N_1113);
xnor U1157 (N_1157,N_1054,N_1122);
or U1158 (N_1158,N_1076,N_1121);
xnor U1159 (N_1159,N_1111,N_1088);
and U1160 (N_1160,N_1051,N_1082);
xnor U1161 (N_1161,N_1087,N_1072);
or U1162 (N_1162,N_1059,N_1064);
xnor U1163 (N_1163,N_1090,N_1053);
or U1164 (N_1164,N_1106,N_1102);
xnor U1165 (N_1165,N_1059,N_1122);
and U1166 (N_1166,N_1054,N_1094);
nand U1167 (N_1167,N_1086,N_1089);
nand U1168 (N_1168,N_1114,N_1073);
or U1169 (N_1169,N_1075,N_1124);
and U1170 (N_1170,N_1110,N_1082);
nor U1171 (N_1171,N_1078,N_1074);
xnor U1172 (N_1172,N_1066,N_1120);
and U1173 (N_1173,N_1056,N_1099);
nand U1174 (N_1174,N_1100,N_1086);
and U1175 (N_1175,N_1121,N_1072);
xor U1176 (N_1176,N_1073,N_1100);
xnor U1177 (N_1177,N_1121,N_1078);
nand U1178 (N_1178,N_1055,N_1109);
or U1179 (N_1179,N_1104,N_1106);
nor U1180 (N_1180,N_1087,N_1076);
xnor U1181 (N_1181,N_1053,N_1095);
and U1182 (N_1182,N_1116,N_1091);
nand U1183 (N_1183,N_1060,N_1090);
nand U1184 (N_1184,N_1118,N_1119);
or U1185 (N_1185,N_1088,N_1119);
xor U1186 (N_1186,N_1069,N_1078);
xnor U1187 (N_1187,N_1102,N_1122);
nand U1188 (N_1188,N_1088,N_1115);
or U1189 (N_1189,N_1104,N_1080);
and U1190 (N_1190,N_1077,N_1091);
nor U1191 (N_1191,N_1082,N_1103);
xnor U1192 (N_1192,N_1108,N_1051);
xor U1193 (N_1193,N_1120,N_1051);
and U1194 (N_1194,N_1114,N_1058);
xnor U1195 (N_1195,N_1101,N_1067);
nand U1196 (N_1196,N_1101,N_1100);
and U1197 (N_1197,N_1057,N_1097);
and U1198 (N_1198,N_1082,N_1099);
or U1199 (N_1199,N_1095,N_1058);
or U1200 (N_1200,N_1192,N_1199);
or U1201 (N_1201,N_1138,N_1160);
or U1202 (N_1202,N_1176,N_1158);
or U1203 (N_1203,N_1151,N_1186);
nor U1204 (N_1204,N_1141,N_1197);
nand U1205 (N_1205,N_1131,N_1198);
or U1206 (N_1206,N_1195,N_1178);
nor U1207 (N_1207,N_1172,N_1165);
xnor U1208 (N_1208,N_1125,N_1169);
and U1209 (N_1209,N_1135,N_1194);
and U1210 (N_1210,N_1133,N_1184);
nand U1211 (N_1211,N_1136,N_1157);
or U1212 (N_1212,N_1166,N_1145);
or U1213 (N_1213,N_1147,N_1180);
or U1214 (N_1214,N_1167,N_1126);
and U1215 (N_1215,N_1161,N_1177);
nand U1216 (N_1216,N_1171,N_1159);
or U1217 (N_1217,N_1128,N_1146);
nand U1218 (N_1218,N_1173,N_1190);
xnor U1219 (N_1219,N_1164,N_1149);
nand U1220 (N_1220,N_1155,N_1189);
nand U1221 (N_1221,N_1170,N_1188);
or U1222 (N_1222,N_1144,N_1140);
and U1223 (N_1223,N_1181,N_1152);
or U1224 (N_1224,N_1153,N_1127);
nor U1225 (N_1225,N_1187,N_1134);
and U1226 (N_1226,N_1154,N_1183);
or U1227 (N_1227,N_1179,N_1130);
or U1228 (N_1228,N_1156,N_1168);
xor U1229 (N_1229,N_1196,N_1191);
nor U1230 (N_1230,N_1182,N_1137);
nand U1231 (N_1231,N_1148,N_1175);
xor U1232 (N_1232,N_1129,N_1143);
xor U1233 (N_1233,N_1174,N_1162);
or U1234 (N_1234,N_1142,N_1139);
xnor U1235 (N_1235,N_1150,N_1132);
and U1236 (N_1236,N_1163,N_1185);
nand U1237 (N_1237,N_1193,N_1187);
nor U1238 (N_1238,N_1147,N_1135);
nor U1239 (N_1239,N_1172,N_1157);
and U1240 (N_1240,N_1190,N_1164);
or U1241 (N_1241,N_1156,N_1199);
and U1242 (N_1242,N_1164,N_1182);
nand U1243 (N_1243,N_1133,N_1172);
xor U1244 (N_1244,N_1197,N_1137);
or U1245 (N_1245,N_1191,N_1141);
or U1246 (N_1246,N_1157,N_1158);
or U1247 (N_1247,N_1183,N_1187);
nand U1248 (N_1248,N_1172,N_1175);
or U1249 (N_1249,N_1175,N_1174);
or U1250 (N_1250,N_1181,N_1165);
xnor U1251 (N_1251,N_1143,N_1134);
or U1252 (N_1252,N_1139,N_1143);
nand U1253 (N_1253,N_1142,N_1167);
nand U1254 (N_1254,N_1125,N_1184);
nand U1255 (N_1255,N_1168,N_1192);
nor U1256 (N_1256,N_1184,N_1172);
xor U1257 (N_1257,N_1191,N_1190);
xnor U1258 (N_1258,N_1172,N_1162);
or U1259 (N_1259,N_1142,N_1170);
nor U1260 (N_1260,N_1196,N_1162);
and U1261 (N_1261,N_1136,N_1196);
or U1262 (N_1262,N_1135,N_1187);
or U1263 (N_1263,N_1193,N_1198);
nand U1264 (N_1264,N_1193,N_1185);
nand U1265 (N_1265,N_1143,N_1138);
and U1266 (N_1266,N_1155,N_1159);
or U1267 (N_1267,N_1171,N_1172);
and U1268 (N_1268,N_1191,N_1161);
nor U1269 (N_1269,N_1150,N_1156);
nand U1270 (N_1270,N_1176,N_1163);
or U1271 (N_1271,N_1169,N_1152);
xnor U1272 (N_1272,N_1186,N_1195);
and U1273 (N_1273,N_1130,N_1156);
nand U1274 (N_1274,N_1193,N_1192);
and U1275 (N_1275,N_1255,N_1243);
or U1276 (N_1276,N_1263,N_1261);
or U1277 (N_1277,N_1204,N_1257);
and U1278 (N_1278,N_1268,N_1230);
xor U1279 (N_1279,N_1241,N_1224);
nand U1280 (N_1280,N_1233,N_1253);
and U1281 (N_1281,N_1209,N_1217);
nand U1282 (N_1282,N_1245,N_1220);
or U1283 (N_1283,N_1254,N_1223);
or U1284 (N_1284,N_1212,N_1225);
nor U1285 (N_1285,N_1269,N_1266);
and U1286 (N_1286,N_1216,N_1265);
nand U1287 (N_1287,N_1264,N_1258);
nor U1288 (N_1288,N_1202,N_1203);
or U1289 (N_1289,N_1231,N_1222);
nor U1290 (N_1290,N_1246,N_1252);
nand U1291 (N_1291,N_1218,N_1206);
xor U1292 (N_1292,N_1229,N_1200);
or U1293 (N_1293,N_1244,N_1221);
or U1294 (N_1294,N_1274,N_1272);
nand U1295 (N_1295,N_1238,N_1256);
nor U1296 (N_1296,N_1267,N_1271);
or U1297 (N_1297,N_1227,N_1240);
and U1298 (N_1298,N_1237,N_1228);
or U1299 (N_1299,N_1235,N_1214);
nor U1300 (N_1300,N_1270,N_1207);
xnor U1301 (N_1301,N_1234,N_1249);
and U1302 (N_1302,N_1210,N_1201);
xnor U1303 (N_1303,N_1273,N_1205);
nor U1304 (N_1304,N_1232,N_1226);
xor U1305 (N_1305,N_1260,N_1219);
nor U1306 (N_1306,N_1208,N_1215);
nand U1307 (N_1307,N_1259,N_1262);
nor U1308 (N_1308,N_1239,N_1213);
or U1309 (N_1309,N_1251,N_1247);
nand U1310 (N_1310,N_1242,N_1211);
nand U1311 (N_1311,N_1250,N_1248);
and U1312 (N_1312,N_1236,N_1261);
xor U1313 (N_1313,N_1213,N_1206);
and U1314 (N_1314,N_1270,N_1253);
xor U1315 (N_1315,N_1208,N_1211);
and U1316 (N_1316,N_1255,N_1204);
or U1317 (N_1317,N_1236,N_1230);
nor U1318 (N_1318,N_1204,N_1220);
nand U1319 (N_1319,N_1206,N_1205);
and U1320 (N_1320,N_1214,N_1268);
or U1321 (N_1321,N_1237,N_1265);
nor U1322 (N_1322,N_1271,N_1213);
xor U1323 (N_1323,N_1242,N_1261);
and U1324 (N_1324,N_1243,N_1248);
xnor U1325 (N_1325,N_1212,N_1252);
xnor U1326 (N_1326,N_1259,N_1256);
xnor U1327 (N_1327,N_1237,N_1231);
xnor U1328 (N_1328,N_1207,N_1259);
and U1329 (N_1329,N_1266,N_1237);
and U1330 (N_1330,N_1207,N_1240);
and U1331 (N_1331,N_1265,N_1214);
xor U1332 (N_1332,N_1264,N_1223);
nand U1333 (N_1333,N_1218,N_1221);
nand U1334 (N_1334,N_1225,N_1208);
and U1335 (N_1335,N_1222,N_1250);
nand U1336 (N_1336,N_1214,N_1242);
xnor U1337 (N_1337,N_1204,N_1245);
xnor U1338 (N_1338,N_1228,N_1274);
nor U1339 (N_1339,N_1243,N_1212);
or U1340 (N_1340,N_1212,N_1247);
nand U1341 (N_1341,N_1269,N_1212);
xor U1342 (N_1342,N_1225,N_1213);
xnor U1343 (N_1343,N_1224,N_1253);
and U1344 (N_1344,N_1229,N_1245);
xor U1345 (N_1345,N_1259,N_1272);
or U1346 (N_1346,N_1217,N_1210);
xor U1347 (N_1347,N_1237,N_1220);
nand U1348 (N_1348,N_1220,N_1258);
nand U1349 (N_1349,N_1218,N_1254);
and U1350 (N_1350,N_1291,N_1334);
xnor U1351 (N_1351,N_1293,N_1303);
nand U1352 (N_1352,N_1287,N_1333);
nand U1353 (N_1353,N_1316,N_1288);
xnor U1354 (N_1354,N_1311,N_1315);
nor U1355 (N_1355,N_1297,N_1275);
nor U1356 (N_1356,N_1289,N_1349);
nor U1357 (N_1357,N_1302,N_1292);
and U1358 (N_1358,N_1306,N_1309);
or U1359 (N_1359,N_1321,N_1331);
nand U1360 (N_1360,N_1296,N_1323);
or U1361 (N_1361,N_1322,N_1282);
xor U1362 (N_1362,N_1336,N_1312);
nand U1363 (N_1363,N_1286,N_1328);
and U1364 (N_1364,N_1338,N_1324);
or U1365 (N_1365,N_1290,N_1325);
nor U1366 (N_1366,N_1305,N_1318);
or U1367 (N_1367,N_1283,N_1277);
or U1368 (N_1368,N_1280,N_1294);
or U1369 (N_1369,N_1342,N_1341);
nand U1370 (N_1370,N_1285,N_1276);
nand U1371 (N_1371,N_1348,N_1313);
nor U1372 (N_1372,N_1279,N_1347);
nor U1373 (N_1373,N_1340,N_1314);
xnor U1374 (N_1374,N_1330,N_1332);
nor U1375 (N_1375,N_1343,N_1326);
nor U1376 (N_1376,N_1301,N_1310);
nand U1377 (N_1377,N_1284,N_1298);
or U1378 (N_1378,N_1299,N_1327);
nand U1379 (N_1379,N_1281,N_1295);
and U1380 (N_1380,N_1300,N_1344);
nand U1381 (N_1381,N_1319,N_1339);
or U1382 (N_1382,N_1307,N_1329);
nand U1383 (N_1383,N_1337,N_1320);
and U1384 (N_1384,N_1345,N_1317);
and U1385 (N_1385,N_1346,N_1335);
nand U1386 (N_1386,N_1308,N_1278);
nor U1387 (N_1387,N_1304,N_1275);
and U1388 (N_1388,N_1275,N_1340);
nand U1389 (N_1389,N_1333,N_1311);
xor U1390 (N_1390,N_1319,N_1300);
nand U1391 (N_1391,N_1281,N_1298);
nor U1392 (N_1392,N_1335,N_1303);
nor U1393 (N_1393,N_1289,N_1342);
nor U1394 (N_1394,N_1316,N_1283);
nor U1395 (N_1395,N_1285,N_1314);
nor U1396 (N_1396,N_1322,N_1280);
xnor U1397 (N_1397,N_1317,N_1335);
and U1398 (N_1398,N_1275,N_1306);
nand U1399 (N_1399,N_1337,N_1306);
and U1400 (N_1400,N_1301,N_1315);
xnor U1401 (N_1401,N_1331,N_1282);
nand U1402 (N_1402,N_1313,N_1294);
and U1403 (N_1403,N_1277,N_1278);
nand U1404 (N_1404,N_1345,N_1342);
nor U1405 (N_1405,N_1279,N_1297);
and U1406 (N_1406,N_1323,N_1334);
xor U1407 (N_1407,N_1312,N_1292);
xor U1408 (N_1408,N_1290,N_1286);
and U1409 (N_1409,N_1337,N_1346);
or U1410 (N_1410,N_1319,N_1326);
nand U1411 (N_1411,N_1317,N_1303);
xor U1412 (N_1412,N_1287,N_1344);
nor U1413 (N_1413,N_1348,N_1323);
or U1414 (N_1414,N_1282,N_1309);
nor U1415 (N_1415,N_1298,N_1304);
and U1416 (N_1416,N_1305,N_1331);
xor U1417 (N_1417,N_1348,N_1286);
and U1418 (N_1418,N_1317,N_1347);
and U1419 (N_1419,N_1346,N_1312);
nand U1420 (N_1420,N_1283,N_1310);
and U1421 (N_1421,N_1338,N_1318);
or U1422 (N_1422,N_1344,N_1321);
xnor U1423 (N_1423,N_1299,N_1347);
or U1424 (N_1424,N_1294,N_1302);
or U1425 (N_1425,N_1423,N_1380);
nor U1426 (N_1426,N_1364,N_1361);
xnor U1427 (N_1427,N_1393,N_1383);
nor U1428 (N_1428,N_1353,N_1415);
or U1429 (N_1429,N_1386,N_1366);
nand U1430 (N_1430,N_1390,N_1387);
xor U1431 (N_1431,N_1352,N_1391);
nand U1432 (N_1432,N_1408,N_1395);
nor U1433 (N_1433,N_1369,N_1399);
nand U1434 (N_1434,N_1424,N_1370);
nor U1435 (N_1435,N_1379,N_1416);
or U1436 (N_1436,N_1407,N_1358);
or U1437 (N_1437,N_1394,N_1357);
nand U1438 (N_1438,N_1367,N_1373);
or U1439 (N_1439,N_1414,N_1365);
nand U1440 (N_1440,N_1363,N_1382);
nor U1441 (N_1441,N_1406,N_1374);
xnor U1442 (N_1442,N_1388,N_1418);
nor U1443 (N_1443,N_1400,N_1362);
nand U1444 (N_1444,N_1385,N_1372);
xnor U1445 (N_1445,N_1381,N_1409);
and U1446 (N_1446,N_1411,N_1376);
and U1447 (N_1447,N_1410,N_1368);
nand U1448 (N_1448,N_1378,N_1360);
and U1449 (N_1449,N_1354,N_1356);
xor U1450 (N_1450,N_1359,N_1404);
or U1451 (N_1451,N_1396,N_1413);
nor U1452 (N_1452,N_1350,N_1420);
and U1453 (N_1453,N_1419,N_1355);
xnor U1454 (N_1454,N_1405,N_1417);
nand U1455 (N_1455,N_1402,N_1398);
or U1456 (N_1456,N_1351,N_1397);
xnor U1457 (N_1457,N_1392,N_1375);
or U1458 (N_1458,N_1403,N_1371);
nor U1459 (N_1459,N_1384,N_1401);
nor U1460 (N_1460,N_1422,N_1412);
nor U1461 (N_1461,N_1421,N_1389);
or U1462 (N_1462,N_1377,N_1360);
nor U1463 (N_1463,N_1403,N_1406);
xor U1464 (N_1464,N_1375,N_1390);
or U1465 (N_1465,N_1372,N_1365);
or U1466 (N_1466,N_1415,N_1424);
nand U1467 (N_1467,N_1358,N_1359);
xor U1468 (N_1468,N_1419,N_1360);
nor U1469 (N_1469,N_1412,N_1386);
and U1470 (N_1470,N_1400,N_1415);
xnor U1471 (N_1471,N_1369,N_1411);
nand U1472 (N_1472,N_1406,N_1422);
nand U1473 (N_1473,N_1391,N_1395);
xor U1474 (N_1474,N_1358,N_1366);
nand U1475 (N_1475,N_1374,N_1368);
nor U1476 (N_1476,N_1405,N_1411);
and U1477 (N_1477,N_1410,N_1354);
nor U1478 (N_1478,N_1364,N_1352);
nor U1479 (N_1479,N_1408,N_1381);
nor U1480 (N_1480,N_1399,N_1382);
xnor U1481 (N_1481,N_1418,N_1407);
nand U1482 (N_1482,N_1351,N_1381);
and U1483 (N_1483,N_1409,N_1373);
nor U1484 (N_1484,N_1354,N_1383);
xor U1485 (N_1485,N_1375,N_1388);
and U1486 (N_1486,N_1415,N_1402);
or U1487 (N_1487,N_1372,N_1406);
xnor U1488 (N_1488,N_1358,N_1404);
or U1489 (N_1489,N_1387,N_1380);
nand U1490 (N_1490,N_1373,N_1356);
and U1491 (N_1491,N_1409,N_1411);
nor U1492 (N_1492,N_1413,N_1424);
nand U1493 (N_1493,N_1362,N_1391);
nand U1494 (N_1494,N_1369,N_1382);
or U1495 (N_1495,N_1413,N_1389);
or U1496 (N_1496,N_1360,N_1391);
nor U1497 (N_1497,N_1372,N_1423);
nand U1498 (N_1498,N_1370,N_1351);
and U1499 (N_1499,N_1418,N_1403);
and U1500 (N_1500,N_1485,N_1447);
nand U1501 (N_1501,N_1433,N_1488);
or U1502 (N_1502,N_1455,N_1432);
nand U1503 (N_1503,N_1476,N_1486);
nor U1504 (N_1504,N_1457,N_1434);
nand U1505 (N_1505,N_1425,N_1487);
xor U1506 (N_1506,N_1436,N_1495);
nor U1507 (N_1507,N_1440,N_1484);
nor U1508 (N_1508,N_1438,N_1470);
xor U1509 (N_1509,N_1472,N_1452);
nand U1510 (N_1510,N_1475,N_1449);
or U1511 (N_1511,N_1426,N_1458);
nor U1512 (N_1512,N_1490,N_1481);
nor U1513 (N_1513,N_1463,N_1429);
xor U1514 (N_1514,N_1446,N_1437);
or U1515 (N_1515,N_1451,N_1441);
xor U1516 (N_1516,N_1428,N_1461);
or U1517 (N_1517,N_1498,N_1480);
nand U1518 (N_1518,N_1499,N_1462);
nand U1519 (N_1519,N_1497,N_1482);
xnor U1520 (N_1520,N_1448,N_1427);
nand U1521 (N_1521,N_1435,N_1468);
nand U1522 (N_1522,N_1460,N_1466);
nor U1523 (N_1523,N_1492,N_1478);
xnor U1524 (N_1524,N_1430,N_1444);
or U1525 (N_1525,N_1442,N_1459);
xnor U1526 (N_1526,N_1469,N_1474);
xnor U1527 (N_1527,N_1473,N_1453);
and U1528 (N_1528,N_1454,N_1494);
and U1529 (N_1529,N_1464,N_1479);
or U1530 (N_1530,N_1477,N_1496);
nor U1531 (N_1531,N_1491,N_1439);
xor U1532 (N_1532,N_1483,N_1443);
or U1533 (N_1533,N_1431,N_1493);
and U1534 (N_1534,N_1465,N_1471);
nand U1535 (N_1535,N_1456,N_1450);
nand U1536 (N_1536,N_1489,N_1467);
nor U1537 (N_1537,N_1445,N_1473);
or U1538 (N_1538,N_1443,N_1425);
or U1539 (N_1539,N_1472,N_1441);
nor U1540 (N_1540,N_1478,N_1453);
xnor U1541 (N_1541,N_1497,N_1493);
nand U1542 (N_1542,N_1450,N_1477);
xnor U1543 (N_1543,N_1466,N_1434);
nand U1544 (N_1544,N_1429,N_1479);
nand U1545 (N_1545,N_1497,N_1468);
xnor U1546 (N_1546,N_1460,N_1491);
nor U1547 (N_1547,N_1466,N_1494);
xnor U1548 (N_1548,N_1491,N_1499);
nor U1549 (N_1549,N_1470,N_1443);
and U1550 (N_1550,N_1468,N_1457);
nand U1551 (N_1551,N_1433,N_1481);
nor U1552 (N_1552,N_1432,N_1444);
or U1553 (N_1553,N_1426,N_1439);
nand U1554 (N_1554,N_1499,N_1465);
and U1555 (N_1555,N_1450,N_1493);
nand U1556 (N_1556,N_1436,N_1430);
and U1557 (N_1557,N_1477,N_1441);
or U1558 (N_1558,N_1487,N_1432);
or U1559 (N_1559,N_1446,N_1453);
and U1560 (N_1560,N_1468,N_1425);
and U1561 (N_1561,N_1472,N_1425);
or U1562 (N_1562,N_1465,N_1444);
nor U1563 (N_1563,N_1459,N_1493);
nand U1564 (N_1564,N_1464,N_1448);
nand U1565 (N_1565,N_1428,N_1462);
nor U1566 (N_1566,N_1483,N_1425);
xor U1567 (N_1567,N_1441,N_1496);
nor U1568 (N_1568,N_1458,N_1427);
nand U1569 (N_1569,N_1434,N_1468);
and U1570 (N_1570,N_1475,N_1471);
or U1571 (N_1571,N_1433,N_1453);
or U1572 (N_1572,N_1455,N_1464);
nor U1573 (N_1573,N_1448,N_1428);
nor U1574 (N_1574,N_1476,N_1459);
nand U1575 (N_1575,N_1535,N_1557);
nor U1576 (N_1576,N_1545,N_1537);
nand U1577 (N_1577,N_1502,N_1572);
nor U1578 (N_1578,N_1536,N_1560);
xnor U1579 (N_1579,N_1539,N_1558);
nor U1580 (N_1580,N_1573,N_1541);
and U1581 (N_1581,N_1530,N_1534);
nor U1582 (N_1582,N_1548,N_1552);
nor U1583 (N_1583,N_1533,N_1544);
and U1584 (N_1584,N_1546,N_1523);
or U1585 (N_1585,N_1527,N_1569);
and U1586 (N_1586,N_1574,N_1570);
nand U1587 (N_1587,N_1531,N_1507);
nand U1588 (N_1588,N_1513,N_1562);
nor U1589 (N_1589,N_1571,N_1540);
xnor U1590 (N_1590,N_1559,N_1508);
nor U1591 (N_1591,N_1521,N_1503);
xnor U1592 (N_1592,N_1549,N_1506);
and U1593 (N_1593,N_1538,N_1517);
nand U1594 (N_1594,N_1514,N_1500);
xor U1595 (N_1595,N_1509,N_1554);
xor U1596 (N_1596,N_1511,N_1512);
or U1597 (N_1597,N_1567,N_1510);
xnor U1598 (N_1598,N_1543,N_1519);
or U1599 (N_1599,N_1551,N_1550);
and U1600 (N_1600,N_1505,N_1515);
nand U1601 (N_1601,N_1518,N_1524);
xnor U1602 (N_1602,N_1564,N_1532);
or U1603 (N_1603,N_1520,N_1501);
xnor U1604 (N_1604,N_1525,N_1568);
nand U1605 (N_1605,N_1563,N_1566);
xnor U1606 (N_1606,N_1516,N_1542);
nand U1607 (N_1607,N_1561,N_1504);
nor U1608 (N_1608,N_1555,N_1522);
nor U1609 (N_1609,N_1556,N_1526);
nand U1610 (N_1610,N_1553,N_1529);
nand U1611 (N_1611,N_1547,N_1528);
or U1612 (N_1612,N_1565,N_1570);
nand U1613 (N_1613,N_1534,N_1573);
or U1614 (N_1614,N_1519,N_1546);
and U1615 (N_1615,N_1541,N_1531);
or U1616 (N_1616,N_1572,N_1508);
nand U1617 (N_1617,N_1569,N_1564);
nor U1618 (N_1618,N_1548,N_1547);
nand U1619 (N_1619,N_1500,N_1570);
nand U1620 (N_1620,N_1522,N_1537);
or U1621 (N_1621,N_1528,N_1516);
nor U1622 (N_1622,N_1551,N_1500);
xor U1623 (N_1623,N_1544,N_1563);
or U1624 (N_1624,N_1516,N_1510);
nor U1625 (N_1625,N_1508,N_1528);
nand U1626 (N_1626,N_1548,N_1531);
xor U1627 (N_1627,N_1544,N_1501);
nand U1628 (N_1628,N_1507,N_1568);
or U1629 (N_1629,N_1554,N_1545);
xor U1630 (N_1630,N_1533,N_1540);
xnor U1631 (N_1631,N_1564,N_1519);
and U1632 (N_1632,N_1573,N_1550);
xor U1633 (N_1633,N_1518,N_1547);
xor U1634 (N_1634,N_1567,N_1553);
nor U1635 (N_1635,N_1515,N_1571);
nand U1636 (N_1636,N_1520,N_1523);
nor U1637 (N_1637,N_1550,N_1531);
nor U1638 (N_1638,N_1548,N_1559);
xnor U1639 (N_1639,N_1563,N_1568);
and U1640 (N_1640,N_1522,N_1514);
nor U1641 (N_1641,N_1544,N_1514);
nor U1642 (N_1642,N_1528,N_1560);
or U1643 (N_1643,N_1510,N_1562);
and U1644 (N_1644,N_1561,N_1549);
xnor U1645 (N_1645,N_1531,N_1559);
nand U1646 (N_1646,N_1505,N_1500);
nand U1647 (N_1647,N_1552,N_1567);
nor U1648 (N_1648,N_1533,N_1572);
nor U1649 (N_1649,N_1515,N_1544);
or U1650 (N_1650,N_1634,N_1619);
and U1651 (N_1651,N_1608,N_1640);
and U1652 (N_1652,N_1592,N_1649);
nand U1653 (N_1653,N_1599,N_1601);
or U1654 (N_1654,N_1631,N_1616);
and U1655 (N_1655,N_1637,N_1636);
xor U1656 (N_1656,N_1578,N_1623);
and U1657 (N_1657,N_1630,N_1588);
or U1658 (N_1658,N_1621,N_1643);
nand U1659 (N_1659,N_1629,N_1605);
or U1660 (N_1660,N_1596,N_1613);
and U1661 (N_1661,N_1593,N_1591);
nor U1662 (N_1662,N_1582,N_1618);
nand U1663 (N_1663,N_1627,N_1644);
or U1664 (N_1664,N_1603,N_1577);
nor U1665 (N_1665,N_1638,N_1625);
nand U1666 (N_1666,N_1598,N_1595);
and U1667 (N_1667,N_1609,N_1615);
nor U1668 (N_1668,N_1633,N_1624);
xnor U1669 (N_1669,N_1585,N_1635);
and U1670 (N_1670,N_1645,N_1579);
nand U1671 (N_1671,N_1586,N_1612);
xnor U1672 (N_1672,N_1587,N_1583);
nor U1673 (N_1673,N_1639,N_1620);
and U1674 (N_1674,N_1642,N_1641);
nand U1675 (N_1675,N_1576,N_1628);
and U1676 (N_1676,N_1575,N_1646);
nand U1677 (N_1677,N_1632,N_1580);
and U1678 (N_1678,N_1597,N_1590);
and U1679 (N_1679,N_1647,N_1614);
nand U1680 (N_1680,N_1602,N_1606);
or U1681 (N_1681,N_1589,N_1584);
and U1682 (N_1682,N_1611,N_1607);
nor U1683 (N_1683,N_1626,N_1600);
or U1684 (N_1684,N_1610,N_1617);
and U1685 (N_1685,N_1581,N_1604);
nor U1686 (N_1686,N_1594,N_1648);
or U1687 (N_1687,N_1622,N_1591);
and U1688 (N_1688,N_1581,N_1586);
nand U1689 (N_1689,N_1608,N_1610);
nand U1690 (N_1690,N_1601,N_1637);
nor U1691 (N_1691,N_1645,N_1632);
nand U1692 (N_1692,N_1579,N_1644);
nand U1693 (N_1693,N_1617,N_1626);
nand U1694 (N_1694,N_1625,N_1617);
nor U1695 (N_1695,N_1612,N_1580);
nand U1696 (N_1696,N_1598,N_1580);
nor U1697 (N_1697,N_1625,N_1645);
xor U1698 (N_1698,N_1596,N_1599);
and U1699 (N_1699,N_1640,N_1623);
nor U1700 (N_1700,N_1645,N_1623);
nand U1701 (N_1701,N_1610,N_1607);
nor U1702 (N_1702,N_1635,N_1599);
or U1703 (N_1703,N_1643,N_1624);
nor U1704 (N_1704,N_1636,N_1606);
nand U1705 (N_1705,N_1640,N_1603);
nor U1706 (N_1706,N_1608,N_1631);
and U1707 (N_1707,N_1600,N_1638);
xor U1708 (N_1708,N_1601,N_1584);
or U1709 (N_1709,N_1587,N_1584);
xor U1710 (N_1710,N_1628,N_1601);
or U1711 (N_1711,N_1643,N_1577);
xor U1712 (N_1712,N_1605,N_1581);
xnor U1713 (N_1713,N_1636,N_1628);
xnor U1714 (N_1714,N_1613,N_1648);
xnor U1715 (N_1715,N_1608,N_1632);
xnor U1716 (N_1716,N_1610,N_1628);
and U1717 (N_1717,N_1637,N_1641);
nand U1718 (N_1718,N_1643,N_1598);
xnor U1719 (N_1719,N_1606,N_1580);
and U1720 (N_1720,N_1605,N_1617);
or U1721 (N_1721,N_1617,N_1611);
nor U1722 (N_1722,N_1588,N_1576);
nor U1723 (N_1723,N_1646,N_1607);
xor U1724 (N_1724,N_1589,N_1646);
or U1725 (N_1725,N_1687,N_1661);
nand U1726 (N_1726,N_1698,N_1650);
xnor U1727 (N_1727,N_1679,N_1673);
and U1728 (N_1728,N_1707,N_1674);
xor U1729 (N_1729,N_1702,N_1655);
nor U1730 (N_1730,N_1690,N_1665);
nor U1731 (N_1731,N_1723,N_1718);
or U1732 (N_1732,N_1667,N_1706);
xor U1733 (N_1733,N_1704,N_1694);
nor U1734 (N_1734,N_1716,N_1703);
nor U1735 (N_1735,N_1684,N_1705);
or U1736 (N_1736,N_1685,N_1714);
and U1737 (N_1737,N_1708,N_1720);
nor U1738 (N_1738,N_1711,N_1683);
and U1739 (N_1739,N_1682,N_1656);
or U1740 (N_1740,N_1681,N_1651);
or U1741 (N_1741,N_1660,N_1680);
and U1742 (N_1742,N_1717,N_1715);
nor U1743 (N_1743,N_1713,N_1653);
and U1744 (N_1744,N_1664,N_1672);
xnor U1745 (N_1745,N_1701,N_1670);
nand U1746 (N_1746,N_1678,N_1677);
nor U1747 (N_1747,N_1658,N_1712);
xor U1748 (N_1748,N_1696,N_1659);
or U1749 (N_1749,N_1724,N_1675);
nor U1750 (N_1750,N_1699,N_1676);
or U1751 (N_1751,N_1662,N_1721);
xor U1752 (N_1752,N_1710,N_1693);
or U1753 (N_1753,N_1689,N_1669);
and U1754 (N_1754,N_1700,N_1657);
nor U1755 (N_1755,N_1671,N_1719);
nand U1756 (N_1756,N_1652,N_1688);
xnor U1757 (N_1757,N_1692,N_1686);
or U1758 (N_1758,N_1663,N_1722);
and U1759 (N_1759,N_1697,N_1666);
xor U1760 (N_1760,N_1691,N_1668);
and U1761 (N_1761,N_1654,N_1709);
nor U1762 (N_1762,N_1695,N_1713);
xnor U1763 (N_1763,N_1674,N_1657);
nand U1764 (N_1764,N_1715,N_1693);
and U1765 (N_1765,N_1705,N_1689);
nor U1766 (N_1766,N_1697,N_1660);
and U1767 (N_1767,N_1651,N_1707);
and U1768 (N_1768,N_1658,N_1690);
xnor U1769 (N_1769,N_1693,N_1670);
xnor U1770 (N_1770,N_1688,N_1721);
and U1771 (N_1771,N_1704,N_1705);
nand U1772 (N_1772,N_1696,N_1704);
and U1773 (N_1773,N_1652,N_1668);
nand U1774 (N_1774,N_1717,N_1663);
nor U1775 (N_1775,N_1698,N_1700);
or U1776 (N_1776,N_1656,N_1717);
nor U1777 (N_1777,N_1663,N_1724);
nand U1778 (N_1778,N_1694,N_1677);
nor U1779 (N_1779,N_1706,N_1716);
or U1780 (N_1780,N_1663,N_1686);
xor U1781 (N_1781,N_1704,N_1720);
and U1782 (N_1782,N_1721,N_1691);
nand U1783 (N_1783,N_1661,N_1706);
nor U1784 (N_1784,N_1714,N_1659);
xnor U1785 (N_1785,N_1669,N_1663);
nand U1786 (N_1786,N_1658,N_1715);
or U1787 (N_1787,N_1706,N_1697);
and U1788 (N_1788,N_1724,N_1716);
nor U1789 (N_1789,N_1654,N_1691);
or U1790 (N_1790,N_1710,N_1699);
nand U1791 (N_1791,N_1670,N_1672);
xnor U1792 (N_1792,N_1663,N_1676);
xor U1793 (N_1793,N_1681,N_1666);
nand U1794 (N_1794,N_1699,N_1682);
and U1795 (N_1795,N_1710,N_1683);
and U1796 (N_1796,N_1696,N_1669);
or U1797 (N_1797,N_1700,N_1715);
nand U1798 (N_1798,N_1717,N_1653);
nor U1799 (N_1799,N_1659,N_1655);
and U1800 (N_1800,N_1756,N_1743);
nor U1801 (N_1801,N_1774,N_1761);
nor U1802 (N_1802,N_1745,N_1752);
nor U1803 (N_1803,N_1737,N_1733);
nand U1804 (N_1804,N_1758,N_1740);
or U1805 (N_1805,N_1769,N_1798);
xor U1806 (N_1806,N_1783,N_1742);
xor U1807 (N_1807,N_1782,N_1792);
xor U1808 (N_1808,N_1754,N_1760);
nor U1809 (N_1809,N_1728,N_1730);
nand U1810 (N_1810,N_1781,N_1777);
xor U1811 (N_1811,N_1771,N_1789);
nor U1812 (N_1812,N_1747,N_1775);
xor U1813 (N_1813,N_1799,N_1770);
nand U1814 (N_1814,N_1746,N_1785);
and U1815 (N_1815,N_1751,N_1776);
nand U1816 (N_1816,N_1734,N_1757);
and U1817 (N_1817,N_1725,N_1741);
xor U1818 (N_1818,N_1795,N_1786);
or U1819 (N_1819,N_1759,N_1731);
nand U1820 (N_1820,N_1727,N_1764);
nor U1821 (N_1821,N_1778,N_1784);
nor U1822 (N_1822,N_1739,N_1762);
and U1823 (N_1823,N_1793,N_1790);
nor U1824 (N_1824,N_1726,N_1765);
and U1825 (N_1825,N_1772,N_1780);
nor U1826 (N_1826,N_1736,N_1787);
nand U1827 (N_1827,N_1768,N_1750);
nand U1828 (N_1828,N_1729,N_1796);
nand U1829 (N_1829,N_1763,N_1735);
xnor U1830 (N_1830,N_1797,N_1791);
nand U1831 (N_1831,N_1788,N_1766);
xnor U1832 (N_1832,N_1794,N_1732);
nand U1833 (N_1833,N_1744,N_1773);
and U1834 (N_1834,N_1749,N_1753);
xnor U1835 (N_1835,N_1779,N_1748);
nand U1836 (N_1836,N_1755,N_1738);
and U1837 (N_1837,N_1767,N_1766);
or U1838 (N_1838,N_1765,N_1747);
and U1839 (N_1839,N_1740,N_1760);
nor U1840 (N_1840,N_1794,N_1752);
nor U1841 (N_1841,N_1731,N_1749);
xnor U1842 (N_1842,N_1751,N_1779);
or U1843 (N_1843,N_1796,N_1770);
and U1844 (N_1844,N_1758,N_1733);
nor U1845 (N_1845,N_1747,N_1753);
and U1846 (N_1846,N_1794,N_1748);
nor U1847 (N_1847,N_1745,N_1778);
nor U1848 (N_1848,N_1772,N_1771);
or U1849 (N_1849,N_1752,N_1791);
nor U1850 (N_1850,N_1760,N_1735);
and U1851 (N_1851,N_1779,N_1732);
xor U1852 (N_1852,N_1799,N_1767);
nand U1853 (N_1853,N_1738,N_1743);
xnor U1854 (N_1854,N_1785,N_1728);
xor U1855 (N_1855,N_1775,N_1798);
nor U1856 (N_1856,N_1736,N_1784);
nor U1857 (N_1857,N_1793,N_1744);
xor U1858 (N_1858,N_1741,N_1791);
nand U1859 (N_1859,N_1725,N_1797);
nand U1860 (N_1860,N_1776,N_1799);
xor U1861 (N_1861,N_1798,N_1728);
nand U1862 (N_1862,N_1744,N_1740);
nand U1863 (N_1863,N_1778,N_1787);
and U1864 (N_1864,N_1794,N_1789);
xnor U1865 (N_1865,N_1745,N_1753);
nor U1866 (N_1866,N_1757,N_1777);
and U1867 (N_1867,N_1785,N_1784);
nand U1868 (N_1868,N_1747,N_1760);
and U1869 (N_1869,N_1755,N_1737);
xor U1870 (N_1870,N_1743,N_1744);
nor U1871 (N_1871,N_1798,N_1739);
xnor U1872 (N_1872,N_1785,N_1754);
or U1873 (N_1873,N_1782,N_1726);
nor U1874 (N_1874,N_1765,N_1755);
xnor U1875 (N_1875,N_1828,N_1874);
xor U1876 (N_1876,N_1804,N_1858);
xnor U1877 (N_1877,N_1853,N_1820);
nor U1878 (N_1878,N_1841,N_1844);
and U1879 (N_1879,N_1833,N_1851);
and U1880 (N_1880,N_1813,N_1812);
xor U1881 (N_1881,N_1817,N_1819);
or U1882 (N_1882,N_1800,N_1854);
nor U1883 (N_1883,N_1802,N_1827);
xnor U1884 (N_1884,N_1837,N_1815);
and U1885 (N_1885,N_1816,N_1801);
nand U1886 (N_1886,N_1863,N_1829);
xnor U1887 (N_1887,N_1869,N_1832);
nor U1888 (N_1888,N_1873,N_1834);
or U1889 (N_1889,N_1866,N_1814);
xnor U1890 (N_1890,N_1864,N_1803);
or U1891 (N_1891,N_1805,N_1865);
and U1892 (N_1892,N_1839,N_1808);
xnor U1893 (N_1893,N_1811,N_1846);
nor U1894 (N_1894,N_1870,N_1843);
or U1895 (N_1895,N_1809,N_1847);
xor U1896 (N_1896,N_1856,N_1842);
or U1897 (N_1897,N_1826,N_1859);
nor U1898 (N_1898,N_1818,N_1862);
or U1899 (N_1899,N_1848,N_1835);
xor U1900 (N_1900,N_1867,N_1861);
or U1901 (N_1901,N_1850,N_1831);
and U1902 (N_1902,N_1868,N_1845);
and U1903 (N_1903,N_1857,N_1810);
xnor U1904 (N_1904,N_1872,N_1806);
or U1905 (N_1905,N_1838,N_1871);
nor U1906 (N_1906,N_1840,N_1860);
nor U1907 (N_1907,N_1836,N_1821);
or U1908 (N_1908,N_1855,N_1807);
nand U1909 (N_1909,N_1825,N_1824);
or U1910 (N_1910,N_1823,N_1849);
nor U1911 (N_1911,N_1852,N_1822);
nor U1912 (N_1912,N_1830,N_1865);
nand U1913 (N_1913,N_1810,N_1855);
xor U1914 (N_1914,N_1826,N_1873);
xnor U1915 (N_1915,N_1865,N_1844);
and U1916 (N_1916,N_1870,N_1828);
nor U1917 (N_1917,N_1833,N_1848);
xnor U1918 (N_1918,N_1822,N_1816);
or U1919 (N_1919,N_1863,N_1835);
or U1920 (N_1920,N_1831,N_1834);
or U1921 (N_1921,N_1829,N_1831);
and U1922 (N_1922,N_1834,N_1806);
or U1923 (N_1923,N_1818,N_1836);
xnor U1924 (N_1924,N_1852,N_1815);
or U1925 (N_1925,N_1832,N_1822);
xor U1926 (N_1926,N_1821,N_1846);
or U1927 (N_1927,N_1830,N_1838);
and U1928 (N_1928,N_1801,N_1872);
nor U1929 (N_1929,N_1837,N_1822);
or U1930 (N_1930,N_1829,N_1848);
and U1931 (N_1931,N_1841,N_1837);
xor U1932 (N_1932,N_1848,N_1849);
or U1933 (N_1933,N_1820,N_1859);
or U1934 (N_1934,N_1871,N_1840);
xnor U1935 (N_1935,N_1848,N_1816);
and U1936 (N_1936,N_1818,N_1852);
xnor U1937 (N_1937,N_1873,N_1856);
nor U1938 (N_1938,N_1809,N_1866);
nor U1939 (N_1939,N_1835,N_1850);
and U1940 (N_1940,N_1811,N_1867);
nor U1941 (N_1941,N_1809,N_1873);
and U1942 (N_1942,N_1871,N_1818);
nor U1943 (N_1943,N_1861,N_1808);
or U1944 (N_1944,N_1811,N_1808);
or U1945 (N_1945,N_1826,N_1835);
xnor U1946 (N_1946,N_1845,N_1818);
nand U1947 (N_1947,N_1805,N_1826);
nor U1948 (N_1948,N_1810,N_1801);
or U1949 (N_1949,N_1838,N_1852);
xor U1950 (N_1950,N_1891,N_1926);
nor U1951 (N_1951,N_1903,N_1917);
or U1952 (N_1952,N_1880,N_1916);
xor U1953 (N_1953,N_1932,N_1904);
and U1954 (N_1954,N_1875,N_1897);
or U1955 (N_1955,N_1918,N_1899);
nor U1956 (N_1956,N_1889,N_1949);
nor U1957 (N_1957,N_1900,N_1901);
nand U1958 (N_1958,N_1943,N_1878);
nand U1959 (N_1959,N_1902,N_1948);
or U1960 (N_1960,N_1911,N_1944);
nor U1961 (N_1961,N_1939,N_1931);
or U1962 (N_1962,N_1887,N_1946);
and U1963 (N_1963,N_1922,N_1938);
nand U1964 (N_1964,N_1913,N_1907);
nand U1965 (N_1965,N_1914,N_1888);
and U1966 (N_1966,N_1929,N_1906);
or U1967 (N_1967,N_1947,N_1879);
or U1968 (N_1968,N_1928,N_1892);
nor U1969 (N_1969,N_1921,N_1908);
or U1970 (N_1970,N_1898,N_1890);
or U1971 (N_1971,N_1893,N_1881);
or U1972 (N_1972,N_1915,N_1883);
and U1973 (N_1973,N_1896,N_1940);
nor U1974 (N_1974,N_1941,N_1927);
nor U1975 (N_1975,N_1920,N_1925);
nor U1976 (N_1976,N_1909,N_1877);
and U1977 (N_1977,N_1930,N_1945);
xnor U1978 (N_1978,N_1894,N_1910);
nor U1979 (N_1979,N_1884,N_1886);
nor U1980 (N_1980,N_1924,N_1936);
nand U1981 (N_1981,N_1912,N_1942);
xnor U1982 (N_1982,N_1885,N_1933);
and U1983 (N_1983,N_1935,N_1937);
and U1984 (N_1984,N_1895,N_1919);
and U1985 (N_1985,N_1876,N_1934);
nor U1986 (N_1986,N_1923,N_1905);
nand U1987 (N_1987,N_1882,N_1889);
nand U1988 (N_1988,N_1919,N_1945);
nand U1989 (N_1989,N_1937,N_1898);
and U1990 (N_1990,N_1895,N_1892);
or U1991 (N_1991,N_1896,N_1930);
nor U1992 (N_1992,N_1886,N_1896);
nor U1993 (N_1993,N_1919,N_1892);
and U1994 (N_1994,N_1892,N_1896);
nand U1995 (N_1995,N_1929,N_1945);
xor U1996 (N_1996,N_1879,N_1938);
and U1997 (N_1997,N_1943,N_1937);
nand U1998 (N_1998,N_1916,N_1949);
or U1999 (N_1999,N_1946,N_1931);
and U2000 (N_2000,N_1912,N_1924);
and U2001 (N_2001,N_1883,N_1893);
nand U2002 (N_2002,N_1930,N_1919);
xor U2003 (N_2003,N_1927,N_1882);
and U2004 (N_2004,N_1932,N_1894);
and U2005 (N_2005,N_1923,N_1941);
or U2006 (N_2006,N_1894,N_1920);
nand U2007 (N_2007,N_1919,N_1910);
or U2008 (N_2008,N_1876,N_1937);
xor U2009 (N_2009,N_1882,N_1920);
and U2010 (N_2010,N_1888,N_1909);
xnor U2011 (N_2011,N_1925,N_1918);
and U2012 (N_2012,N_1894,N_1915);
nand U2013 (N_2013,N_1882,N_1885);
and U2014 (N_2014,N_1885,N_1912);
or U2015 (N_2015,N_1912,N_1879);
xor U2016 (N_2016,N_1938,N_1896);
nor U2017 (N_2017,N_1914,N_1886);
nand U2018 (N_2018,N_1878,N_1881);
nor U2019 (N_2019,N_1926,N_1928);
nor U2020 (N_2020,N_1933,N_1942);
or U2021 (N_2021,N_1940,N_1920);
nor U2022 (N_2022,N_1940,N_1923);
xor U2023 (N_2023,N_1937,N_1931);
nor U2024 (N_2024,N_1907,N_1927);
or U2025 (N_2025,N_2017,N_1976);
nor U2026 (N_2026,N_2023,N_1961);
xnor U2027 (N_2027,N_1966,N_1987);
nor U2028 (N_2028,N_1999,N_1972);
or U2029 (N_2029,N_2005,N_2020);
and U2030 (N_2030,N_1971,N_1969);
nor U2031 (N_2031,N_2003,N_2015);
and U2032 (N_2032,N_1980,N_1973);
xnor U2033 (N_2033,N_1952,N_2018);
nand U2034 (N_2034,N_1957,N_1992);
nor U2035 (N_2035,N_2019,N_1964);
nand U2036 (N_2036,N_1986,N_1981);
nor U2037 (N_2037,N_1955,N_1967);
nor U2038 (N_2038,N_2014,N_1959);
and U2039 (N_2039,N_2024,N_1956);
xnor U2040 (N_2040,N_1997,N_1991);
nand U2041 (N_2041,N_1974,N_1996);
or U2042 (N_2042,N_1960,N_2006);
nand U2043 (N_2043,N_2010,N_2007);
nand U2044 (N_2044,N_1989,N_2021);
nand U2045 (N_2045,N_2000,N_1950);
nand U2046 (N_2046,N_1951,N_1968);
nand U2047 (N_2047,N_2001,N_1963);
xnor U2048 (N_2048,N_2012,N_1995);
xnor U2049 (N_2049,N_1993,N_1962);
nor U2050 (N_2050,N_1979,N_1953);
or U2051 (N_2051,N_1977,N_2016);
xnor U2052 (N_2052,N_1998,N_2009);
nand U2053 (N_2053,N_1988,N_2002);
or U2054 (N_2054,N_2004,N_1994);
and U2055 (N_2055,N_2013,N_1982);
nor U2056 (N_2056,N_2011,N_1975);
or U2057 (N_2057,N_1985,N_1965);
nand U2058 (N_2058,N_1978,N_1970);
xnor U2059 (N_2059,N_1990,N_2008);
and U2060 (N_2060,N_1958,N_1984);
and U2061 (N_2061,N_2022,N_1983);
or U2062 (N_2062,N_1954,N_1991);
nand U2063 (N_2063,N_2017,N_1997);
xnor U2064 (N_2064,N_1968,N_2006);
nor U2065 (N_2065,N_2018,N_1962);
xnor U2066 (N_2066,N_1980,N_2015);
xnor U2067 (N_2067,N_1960,N_2020);
and U2068 (N_2068,N_1977,N_1990);
and U2069 (N_2069,N_1990,N_1965);
xnor U2070 (N_2070,N_1951,N_1958);
and U2071 (N_2071,N_1987,N_1974);
xnor U2072 (N_2072,N_1980,N_1968);
nand U2073 (N_2073,N_2017,N_1964);
nor U2074 (N_2074,N_1965,N_1970);
nor U2075 (N_2075,N_1967,N_2014);
and U2076 (N_2076,N_1997,N_1998);
and U2077 (N_2077,N_1981,N_1961);
and U2078 (N_2078,N_1950,N_1964);
xor U2079 (N_2079,N_2022,N_1959);
or U2080 (N_2080,N_2003,N_2012);
and U2081 (N_2081,N_1992,N_1986);
xnor U2082 (N_2082,N_2020,N_2001);
nand U2083 (N_2083,N_1985,N_1999);
xnor U2084 (N_2084,N_2000,N_1964);
nand U2085 (N_2085,N_1983,N_1967);
nand U2086 (N_2086,N_1974,N_1976);
xor U2087 (N_2087,N_1958,N_1971);
and U2088 (N_2088,N_1954,N_1970);
nor U2089 (N_2089,N_1972,N_2012);
nand U2090 (N_2090,N_2008,N_1963);
xnor U2091 (N_2091,N_1952,N_1995);
and U2092 (N_2092,N_1976,N_2023);
nand U2093 (N_2093,N_1967,N_1970);
xor U2094 (N_2094,N_1958,N_2003);
or U2095 (N_2095,N_1967,N_1964);
xor U2096 (N_2096,N_1988,N_1992);
nand U2097 (N_2097,N_2003,N_2010);
xnor U2098 (N_2098,N_1973,N_1978);
xor U2099 (N_2099,N_2000,N_1973);
or U2100 (N_2100,N_2055,N_2041);
and U2101 (N_2101,N_2082,N_2079);
nand U2102 (N_2102,N_2094,N_2070);
and U2103 (N_2103,N_2047,N_2044);
and U2104 (N_2104,N_2077,N_2075);
nor U2105 (N_2105,N_2091,N_2027);
xor U2106 (N_2106,N_2026,N_2053);
nand U2107 (N_2107,N_2029,N_2043);
nand U2108 (N_2108,N_2031,N_2067);
nor U2109 (N_2109,N_2085,N_2093);
or U2110 (N_2110,N_2042,N_2061);
nand U2111 (N_2111,N_2064,N_2095);
and U2112 (N_2112,N_2090,N_2046);
xor U2113 (N_2113,N_2034,N_2089);
xnor U2114 (N_2114,N_2065,N_2032);
or U2115 (N_2115,N_2050,N_2096);
xor U2116 (N_2116,N_2051,N_2038);
nor U2117 (N_2117,N_2037,N_2066);
nor U2118 (N_2118,N_2039,N_2098);
xor U2119 (N_2119,N_2059,N_2099);
nor U2120 (N_2120,N_2048,N_2057);
or U2121 (N_2121,N_2060,N_2056);
and U2122 (N_2122,N_2054,N_2097);
nand U2123 (N_2123,N_2058,N_2028);
nor U2124 (N_2124,N_2087,N_2081);
nor U2125 (N_2125,N_2083,N_2074);
xor U2126 (N_2126,N_2078,N_2076);
nor U2127 (N_2127,N_2080,N_2033);
nand U2128 (N_2128,N_2040,N_2068);
and U2129 (N_2129,N_2071,N_2084);
or U2130 (N_2130,N_2072,N_2049);
xor U2131 (N_2131,N_2030,N_2063);
or U2132 (N_2132,N_2045,N_2035);
or U2133 (N_2133,N_2052,N_2062);
and U2134 (N_2134,N_2073,N_2036);
xnor U2135 (N_2135,N_2088,N_2092);
or U2136 (N_2136,N_2086,N_2025);
or U2137 (N_2137,N_2069,N_2060);
xnor U2138 (N_2138,N_2072,N_2052);
nand U2139 (N_2139,N_2085,N_2063);
xor U2140 (N_2140,N_2043,N_2086);
and U2141 (N_2141,N_2054,N_2048);
nand U2142 (N_2142,N_2099,N_2056);
and U2143 (N_2143,N_2054,N_2051);
and U2144 (N_2144,N_2050,N_2034);
xor U2145 (N_2145,N_2060,N_2094);
or U2146 (N_2146,N_2050,N_2069);
nand U2147 (N_2147,N_2060,N_2066);
nor U2148 (N_2148,N_2028,N_2086);
nand U2149 (N_2149,N_2076,N_2090);
nor U2150 (N_2150,N_2054,N_2042);
nand U2151 (N_2151,N_2096,N_2028);
and U2152 (N_2152,N_2099,N_2064);
and U2153 (N_2153,N_2092,N_2027);
or U2154 (N_2154,N_2065,N_2095);
nor U2155 (N_2155,N_2039,N_2058);
nand U2156 (N_2156,N_2054,N_2036);
and U2157 (N_2157,N_2079,N_2032);
xnor U2158 (N_2158,N_2027,N_2028);
nor U2159 (N_2159,N_2092,N_2033);
or U2160 (N_2160,N_2074,N_2035);
xor U2161 (N_2161,N_2092,N_2089);
xor U2162 (N_2162,N_2082,N_2084);
nor U2163 (N_2163,N_2068,N_2045);
and U2164 (N_2164,N_2079,N_2048);
nand U2165 (N_2165,N_2053,N_2049);
and U2166 (N_2166,N_2049,N_2075);
and U2167 (N_2167,N_2094,N_2026);
and U2168 (N_2168,N_2050,N_2099);
nand U2169 (N_2169,N_2069,N_2081);
and U2170 (N_2170,N_2099,N_2044);
or U2171 (N_2171,N_2063,N_2082);
nand U2172 (N_2172,N_2076,N_2057);
nand U2173 (N_2173,N_2042,N_2096);
or U2174 (N_2174,N_2085,N_2054);
nand U2175 (N_2175,N_2124,N_2111);
and U2176 (N_2176,N_2121,N_2122);
and U2177 (N_2177,N_2148,N_2139);
xor U2178 (N_2178,N_2131,N_2166);
nor U2179 (N_2179,N_2144,N_2160);
or U2180 (N_2180,N_2154,N_2153);
xnor U2181 (N_2181,N_2109,N_2105);
xnor U2182 (N_2182,N_2103,N_2155);
nand U2183 (N_2183,N_2140,N_2150);
nor U2184 (N_2184,N_2116,N_2169);
xnor U2185 (N_2185,N_2151,N_2145);
or U2186 (N_2186,N_2164,N_2125);
or U2187 (N_2187,N_2152,N_2114);
nand U2188 (N_2188,N_2146,N_2119);
xnor U2189 (N_2189,N_2134,N_2168);
xnor U2190 (N_2190,N_2171,N_2115);
or U2191 (N_2191,N_2138,N_2107);
xnor U2192 (N_2192,N_2133,N_2128);
nor U2193 (N_2193,N_2126,N_2147);
or U2194 (N_2194,N_2101,N_2100);
nand U2195 (N_2195,N_2135,N_2143);
xor U2196 (N_2196,N_2127,N_2161);
and U2197 (N_2197,N_2137,N_2158);
nand U2198 (N_2198,N_2123,N_2163);
or U2199 (N_2199,N_2129,N_2104);
or U2200 (N_2200,N_2162,N_2156);
nor U2201 (N_2201,N_2165,N_2118);
xnor U2202 (N_2202,N_2170,N_2117);
nand U2203 (N_2203,N_2110,N_2142);
and U2204 (N_2204,N_2167,N_2173);
nand U2205 (N_2205,N_2113,N_2120);
nand U2206 (N_2206,N_2174,N_2141);
and U2207 (N_2207,N_2112,N_2130);
and U2208 (N_2208,N_2106,N_2136);
nor U2209 (N_2209,N_2102,N_2108);
xnor U2210 (N_2210,N_2159,N_2172);
nor U2211 (N_2211,N_2157,N_2132);
xnor U2212 (N_2212,N_2149,N_2101);
and U2213 (N_2213,N_2167,N_2109);
or U2214 (N_2214,N_2113,N_2134);
and U2215 (N_2215,N_2108,N_2101);
or U2216 (N_2216,N_2140,N_2129);
or U2217 (N_2217,N_2108,N_2166);
and U2218 (N_2218,N_2106,N_2137);
or U2219 (N_2219,N_2138,N_2119);
and U2220 (N_2220,N_2149,N_2152);
or U2221 (N_2221,N_2114,N_2132);
nor U2222 (N_2222,N_2113,N_2125);
or U2223 (N_2223,N_2114,N_2150);
xnor U2224 (N_2224,N_2104,N_2110);
nand U2225 (N_2225,N_2144,N_2112);
nor U2226 (N_2226,N_2151,N_2101);
nor U2227 (N_2227,N_2103,N_2102);
nor U2228 (N_2228,N_2103,N_2144);
and U2229 (N_2229,N_2161,N_2107);
or U2230 (N_2230,N_2152,N_2169);
nor U2231 (N_2231,N_2126,N_2100);
xnor U2232 (N_2232,N_2132,N_2144);
nand U2233 (N_2233,N_2168,N_2133);
and U2234 (N_2234,N_2144,N_2161);
xnor U2235 (N_2235,N_2144,N_2163);
or U2236 (N_2236,N_2141,N_2167);
nor U2237 (N_2237,N_2145,N_2122);
nand U2238 (N_2238,N_2113,N_2168);
nand U2239 (N_2239,N_2164,N_2173);
or U2240 (N_2240,N_2173,N_2131);
and U2241 (N_2241,N_2143,N_2111);
nand U2242 (N_2242,N_2166,N_2167);
xnor U2243 (N_2243,N_2113,N_2156);
and U2244 (N_2244,N_2103,N_2125);
or U2245 (N_2245,N_2163,N_2104);
nor U2246 (N_2246,N_2152,N_2139);
xor U2247 (N_2247,N_2171,N_2119);
or U2248 (N_2248,N_2120,N_2106);
nor U2249 (N_2249,N_2153,N_2119);
xor U2250 (N_2250,N_2197,N_2196);
or U2251 (N_2251,N_2190,N_2248);
or U2252 (N_2252,N_2208,N_2205);
xnor U2253 (N_2253,N_2204,N_2221);
xnor U2254 (N_2254,N_2189,N_2231);
xor U2255 (N_2255,N_2182,N_2233);
and U2256 (N_2256,N_2238,N_2193);
xor U2257 (N_2257,N_2178,N_2224);
or U2258 (N_2258,N_2249,N_2181);
nor U2259 (N_2259,N_2239,N_2247);
nand U2260 (N_2260,N_2226,N_2215);
nor U2261 (N_2261,N_2246,N_2232);
nand U2262 (N_2262,N_2211,N_2244);
nand U2263 (N_2263,N_2242,N_2187);
and U2264 (N_2264,N_2230,N_2235);
xnor U2265 (N_2265,N_2206,N_2228);
nand U2266 (N_2266,N_2183,N_2237);
or U2267 (N_2267,N_2202,N_2175);
nor U2268 (N_2268,N_2212,N_2214);
nor U2269 (N_2269,N_2188,N_2207);
nor U2270 (N_2270,N_2184,N_2201);
nor U2271 (N_2271,N_2245,N_2195);
nand U2272 (N_2272,N_2186,N_2222);
xor U2273 (N_2273,N_2203,N_2236);
nand U2274 (N_2274,N_2217,N_2225);
nand U2275 (N_2275,N_2191,N_2243);
nor U2276 (N_2276,N_2185,N_2240);
nor U2277 (N_2277,N_2199,N_2213);
or U2278 (N_2278,N_2218,N_2198);
or U2279 (N_2279,N_2216,N_2223);
xnor U2280 (N_2280,N_2176,N_2241);
nor U2281 (N_2281,N_2209,N_2192);
nor U2282 (N_2282,N_2227,N_2200);
and U2283 (N_2283,N_2210,N_2194);
and U2284 (N_2284,N_2219,N_2180);
nor U2285 (N_2285,N_2179,N_2177);
and U2286 (N_2286,N_2229,N_2234);
and U2287 (N_2287,N_2220,N_2185);
nor U2288 (N_2288,N_2208,N_2249);
xnor U2289 (N_2289,N_2229,N_2197);
nor U2290 (N_2290,N_2178,N_2238);
nand U2291 (N_2291,N_2220,N_2190);
nand U2292 (N_2292,N_2206,N_2190);
nor U2293 (N_2293,N_2202,N_2212);
and U2294 (N_2294,N_2198,N_2193);
nor U2295 (N_2295,N_2221,N_2195);
nand U2296 (N_2296,N_2179,N_2211);
nor U2297 (N_2297,N_2229,N_2210);
xor U2298 (N_2298,N_2217,N_2214);
nand U2299 (N_2299,N_2188,N_2184);
and U2300 (N_2300,N_2231,N_2203);
and U2301 (N_2301,N_2235,N_2184);
nand U2302 (N_2302,N_2187,N_2248);
or U2303 (N_2303,N_2242,N_2191);
and U2304 (N_2304,N_2202,N_2186);
nand U2305 (N_2305,N_2233,N_2200);
nand U2306 (N_2306,N_2239,N_2206);
or U2307 (N_2307,N_2196,N_2231);
or U2308 (N_2308,N_2183,N_2227);
nand U2309 (N_2309,N_2235,N_2218);
nand U2310 (N_2310,N_2211,N_2237);
and U2311 (N_2311,N_2224,N_2177);
and U2312 (N_2312,N_2229,N_2199);
nand U2313 (N_2313,N_2197,N_2231);
nand U2314 (N_2314,N_2211,N_2194);
xnor U2315 (N_2315,N_2193,N_2232);
or U2316 (N_2316,N_2198,N_2195);
nand U2317 (N_2317,N_2248,N_2195);
and U2318 (N_2318,N_2209,N_2182);
nor U2319 (N_2319,N_2245,N_2189);
or U2320 (N_2320,N_2229,N_2218);
nand U2321 (N_2321,N_2231,N_2239);
nand U2322 (N_2322,N_2247,N_2197);
xnor U2323 (N_2323,N_2219,N_2186);
xor U2324 (N_2324,N_2197,N_2184);
xnor U2325 (N_2325,N_2261,N_2254);
nor U2326 (N_2326,N_2324,N_2253);
or U2327 (N_2327,N_2263,N_2297);
nor U2328 (N_2328,N_2256,N_2271);
and U2329 (N_2329,N_2316,N_2270);
or U2330 (N_2330,N_2296,N_2302);
xor U2331 (N_2331,N_2260,N_2269);
nor U2332 (N_2332,N_2288,N_2265);
nand U2333 (N_2333,N_2251,N_2282);
nor U2334 (N_2334,N_2262,N_2268);
and U2335 (N_2335,N_2313,N_2323);
or U2336 (N_2336,N_2275,N_2295);
nor U2337 (N_2337,N_2298,N_2317);
nor U2338 (N_2338,N_2287,N_2320);
nand U2339 (N_2339,N_2278,N_2321);
nor U2340 (N_2340,N_2294,N_2283);
and U2341 (N_2341,N_2318,N_2274);
or U2342 (N_2342,N_2255,N_2307);
nand U2343 (N_2343,N_2314,N_2290);
and U2344 (N_2344,N_2315,N_2277);
and U2345 (N_2345,N_2259,N_2272);
xnor U2346 (N_2346,N_2305,N_2309);
and U2347 (N_2347,N_2299,N_2285);
xnor U2348 (N_2348,N_2284,N_2289);
and U2349 (N_2349,N_2304,N_2292);
and U2350 (N_2350,N_2280,N_2311);
and U2351 (N_2351,N_2291,N_2286);
xor U2352 (N_2352,N_2300,N_2301);
xor U2353 (N_2353,N_2312,N_2258);
xnor U2354 (N_2354,N_2266,N_2306);
or U2355 (N_2355,N_2257,N_2276);
nand U2356 (N_2356,N_2279,N_2281);
xnor U2357 (N_2357,N_2319,N_2250);
xnor U2358 (N_2358,N_2293,N_2267);
nand U2359 (N_2359,N_2273,N_2308);
nor U2360 (N_2360,N_2310,N_2322);
nand U2361 (N_2361,N_2264,N_2303);
or U2362 (N_2362,N_2252,N_2255);
or U2363 (N_2363,N_2252,N_2262);
xor U2364 (N_2364,N_2319,N_2261);
nor U2365 (N_2365,N_2313,N_2291);
or U2366 (N_2366,N_2278,N_2263);
nor U2367 (N_2367,N_2257,N_2300);
or U2368 (N_2368,N_2286,N_2297);
or U2369 (N_2369,N_2313,N_2251);
nand U2370 (N_2370,N_2275,N_2304);
xnor U2371 (N_2371,N_2283,N_2276);
nand U2372 (N_2372,N_2298,N_2295);
nor U2373 (N_2373,N_2309,N_2274);
or U2374 (N_2374,N_2277,N_2320);
xor U2375 (N_2375,N_2284,N_2273);
nor U2376 (N_2376,N_2321,N_2285);
nor U2377 (N_2377,N_2253,N_2278);
nand U2378 (N_2378,N_2308,N_2269);
or U2379 (N_2379,N_2295,N_2262);
nand U2380 (N_2380,N_2273,N_2299);
and U2381 (N_2381,N_2298,N_2293);
xnor U2382 (N_2382,N_2286,N_2306);
and U2383 (N_2383,N_2257,N_2258);
nor U2384 (N_2384,N_2279,N_2309);
xnor U2385 (N_2385,N_2307,N_2304);
xor U2386 (N_2386,N_2320,N_2307);
xnor U2387 (N_2387,N_2311,N_2283);
nor U2388 (N_2388,N_2287,N_2268);
nand U2389 (N_2389,N_2257,N_2296);
nand U2390 (N_2390,N_2257,N_2269);
nand U2391 (N_2391,N_2269,N_2275);
and U2392 (N_2392,N_2286,N_2319);
xnor U2393 (N_2393,N_2260,N_2273);
and U2394 (N_2394,N_2263,N_2311);
nor U2395 (N_2395,N_2257,N_2297);
nor U2396 (N_2396,N_2318,N_2272);
or U2397 (N_2397,N_2324,N_2289);
xnor U2398 (N_2398,N_2293,N_2257);
and U2399 (N_2399,N_2260,N_2267);
nor U2400 (N_2400,N_2367,N_2378);
xor U2401 (N_2401,N_2338,N_2325);
and U2402 (N_2402,N_2356,N_2348);
and U2403 (N_2403,N_2355,N_2357);
or U2404 (N_2404,N_2346,N_2333);
or U2405 (N_2405,N_2397,N_2366);
nand U2406 (N_2406,N_2369,N_2335);
nor U2407 (N_2407,N_2392,N_2387);
xor U2408 (N_2408,N_2375,N_2391);
and U2409 (N_2409,N_2388,N_2354);
nor U2410 (N_2410,N_2327,N_2352);
xnor U2411 (N_2411,N_2351,N_2339);
or U2412 (N_2412,N_2374,N_2363);
nor U2413 (N_2413,N_2362,N_2399);
or U2414 (N_2414,N_2398,N_2336);
nand U2415 (N_2415,N_2381,N_2389);
nand U2416 (N_2416,N_2353,N_2332);
and U2417 (N_2417,N_2393,N_2383);
nor U2418 (N_2418,N_2326,N_2347);
nand U2419 (N_2419,N_2394,N_2361);
or U2420 (N_2420,N_2384,N_2371);
or U2421 (N_2421,N_2379,N_2395);
or U2422 (N_2422,N_2341,N_2328);
and U2423 (N_2423,N_2386,N_2343);
or U2424 (N_2424,N_2364,N_2358);
and U2425 (N_2425,N_2370,N_2329);
or U2426 (N_2426,N_2350,N_2331);
and U2427 (N_2427,N_2349,N_2359);
or U2428 (N_2428,N_2385,N_2376);
and U2429 (N_2429,N_2344,N_2337);
nor U2430 (N_2430,N_2345,N_2377);
nor U2431 (N_2431,N_2340,N_2390);
nand U2432 (N_2432,N_2373,N_2382);
and U2433 (N_2433,N_2396,N_2342);
and U2434 (N_2434,N_2372,N_2380);
or U2435 (N_2435,N_2368,N_2365);
or U2436 (N_2436,N_2360,N_2330);
and U2437 (N_2437,N_2334,N_2344);
nand U2438 (N_2438,N_2325,N_2342);
nand U2439 (N_2439,N_2344,N_2332);
nand U2440 (N_2440,N_2341,N_2363);
or U2441 (N_2441,N_2354,N_2328);
and U2442 (N_2442,N_2362,N_2371);
or U2443 (N_2443,N_2373,N_2371);
nand U2444 (N_2444,N_2366,N_2389);
xnor U2445 (N_2445,N_2392,N_2373);
nand U2446 (N_2446,N_2370,N_2361);
xnor U2447 (N_2447,N_2353,N_2398);
nor U2448 (N_2448,N_2345,N_2389);
xor U2449 (N_2449,N_2382,N_2389);
and U2450 (N_2450,N_2350,N_2362);
nor U2451 (N_2451,N_2360,N_2340);
nand U2452 (N_2452,N_2380,N_2383);
or U2453 (N_2453,N_2390,N_2374);
nor U2454 (N_2454,N_2362,N_2377);
or U2455 (N_2455,N_2382,N_2380);
and U2456 (N_2456,N_2391,N_2384);
nor U2457 (N_2457,N_2379,N_2377);
nand U2458 (N_2458,N_2388,N_2390);
or U2459 (N_2459,N_2375,N_2386);
and U2460 (N_2460,N_2361,N_2385);
or U2461 (N_2461,N_2382,N_2325);
xor U2462 (N_2462,N_2399,N_2350);
nor U2463 (N_2463,N_2353,N_2373);
nor U2464 (N_2464,N_2352,N_2378);
nor U2465 (N_2465,N_2335,N_2358);
nand U2466 (N_2466,N_2338,N_2328);
nand U2467 (N_2467,N_2389,N_2327);
or U2468 (N_2468,N_2388,N_2335);
nand U2469 (N_2469,N_2328,N_2398);
or U2470 (N_2470,N_2327,N_2336);
and U2471 (N_2471,N_2397,N_2394);
or U2472 (N_2472,N_2339,N_2366);
and U2473 (N_2473,N_2343,N_2393);
xnor U2474 (N_2474,N_2383,N_2336);
nor U2475 (N_2475,N_2403,N_2469);
or U2476 (N_2476,N_2444,N_2414);
or U2477 (N_2477,N_2472,N_2439);
xor U2478 (N_2478,N_2409,N_2420);
xor U2479 (N_2479,N_2466,N_2452);
nor U2480 (N_2480,N_2461,N_2429);
nor U2481 (N_2481,N_2412,N_2437);
or U2482 (N_2482,N_2425,N_2405);
and U2483 (N_2483,N_2434,N_2458);
xnor U2484 (N_2484,N_2438,N_2448);
nand U2485 (N_2485,N_2449,N_2465);
and U2486 (N_2486,N_2443,N_2424);
nor U2487 (N_2487,N_2456,N_2459);
xor U2488 (N_2488,N_2428,N_2470);
nor U2489 (N_2489,N_2455,N_2407);
nand U2490 (N_2490,N_2401,N_2415);
xnor U2491 (N_2491,N_2411,N_2446);
and U2492 (N_2492,N_2436,N_2430);
and U2493 (N_2493,N_2408,N_2473);
and U2494 (N_2494,N_2447,N_2462);
nand U2495 (N_2495,N_2418,N_2410);
or U2496 (N_2496,N_2432,N_2433);
or U2497 (N_2497,N_2467,N_2426);
xnor U2498 (N_2498,N_2417,N_2402);
nor U2499 (N_2499,N_2460,N_2471);
nor U2500 (N_2500,N_2441,N_2400);
xnor U2501 (N_2501,N_2463,N_2404);
or U2502 (N_2502,N_2468,N_2450);
nand U2503 (N_2503,N_2431,N_2413);
xor U2504 (N_2504,N_2440,N_2442);
nor U2505 (N_2505,N_2474,N_2435);
or U2506 (N_2506,N_2451,N_2419);
or U2507 (N_2507,N_2427,N_2454);
nor U2508 (N_2508,N_2422,N_2421);
nor U2509 (N_2509,N_2457,N_2406);
nor U2510 (N_2510,N_2453,N_2423);
xnor U2511 (N_2511,N_2464,N_2445);
xnor U2512 (N_2512,N_2416,N_2467);
xor U2513 (N_2513,N_2446,N_2440);
nand U2514 (N_2514,N_2416,N_2431);
or U2515 (N_2515,N_2435,N_2468);
or U2516 (N_2516,N_2400,N_2416);
nor U2517 (N_2517,N_2465,N_2405);
nand U2518 (N_2518,N_2441,N_2464);
or U2519 (N_2519,N_2415,N_2416);
or U2520 (N_2520,N_2413,N_2429);
or U2521 (N_2521,N_2401,N_2417);
and U2522 (N_2522,N_2471,N_2451);
and U2523 (N_2523,N_2428,N_2422);
nand U2524 (N_2524,N_2442,N_2425);
and U2525 (N_2525,N_2443,N_2447);
nand U2526 (N_2526,N_2452,N_2429);
nand U2527 (N_2527,N_2413,N_2472);
nand U2528 (N_2528,N_2431,N_2452);
nor U2529 (N_2529,N_2440,N_2450);
xnor U2530 (N_2530,N_2405,N_2408);
nor U2531 (N_2531,N_2431,N_2445);
or U2532 (N_2532,N_2458,N_2471);
xor U2533 (N_2533,N_2461,N_2427);
xor U2534 (N_2534,N_2424,N_2432);
nand U2535 (N_2535,N_2457,N_2416);
or U2536 (N_2536,N_2438,N_2459);
xnor U2537 (N_2537,N_2411,N_2438);
and U2538 (N_2538,N_2461,N_2443);
and U2539 (N_2539,N_2410,N_2414);
or U2540 (N_2540,N_2412,N_2426);
nand U2541 (N_2541,N_2425,N_2435);
or U2542 (N_2542,N_2453,N_2400);
xnor U2543 (N_2543,N_2437,N_2462);
xnor U2544 (N_2544,N_2431,N_2414);
or U2545 (N_2545,N_2458,N_2431);
and U2546 (N_2546,N_2470,N_2471);
or U2547 (N_2547,N_2444,N_2472);
or U2548 (N_2548,N_2414,N_2437);
and U2549 (N_2549,N_2408,N_2416);
and U2550 (N_2550,N_2529,N_2523);
and U2551 (N_2551,N_2520,N_2521);
and U2552 (N_2552,N_2508,N_2493);
xnor U2553 (N_2553,N_2506,N_2512);
nand U2554 (N_2554,N_2505,N_2538);
nand U2555 (N_2555,N_2500,N_2504);
nand U2556 (N_2556,N_2507,N_2478);
nand U2557 (N_2557,N_2539,N_2537);
xnor U2558 (N_2558,N_2491,N_2499);
or U2559 (N_2559,N_2483,N_2525);
nor U2560 (N_2560,N_2502,N_2485);
nor U2561 (N_2561,N_2503,N_2541);
and U2562 (N_2562,N_2527,N_2482);
nand U2563 (N_2563,N_2479,N_2518);
and U2564 (N_2564,N_2494,N_2495);
nand U2565 (N_2565,N_2490,N_2498);
nor U2566 (N_2566,N_2497,N_2545);
nand U2567 (N_2567,N_2544,N_2510);
nor U2568 (N_2568,N_2522,N_2533);
xor U2569 (N_2569,N_2517,N_2531);
or U2570 (N_2570,N_2475,N_2519);
and U2571 (N_2571,N_2487,N_2496);
nor U2572 (N_2572,N_2536,N_2480);
nor U2573 (N_2573,N_2477,N_2484);
or U2574 (N_2574,N_2511,N_2492);
nor U2575 (N_2575,N_2509,N_2548);
nor U2576 (N_2576,N_2501,N_2549);
or U2577 (N_2577,N_2514,N_2513);
and U2578 (N_2578,N_2546,N_2540);
xor U2579 (N_2579,N_2515,N_2486);
and U2580 (N_2580,N_2535,N_2530);
xnor U2581 (N_2581,N_2488,N_2476);
or U2582 (N_2582,N_2532,N_2524);
and U2583 (N_2583,N_2516,N_2526);
xor U2584 (N_2584,N_2542,N_2481);
nor U2585 (N_2585,N_2547,N_2528);
nor U2586 (N_2586,N_2543,N_2489);
and U2587 (N_2587,N_2534,N_2528);
nand U2588 (N_2588,N_2486,N_2477);
and U2589 (N_2589,N_2526,N_2522);
xnor U2590 (N_2590,N_2482,N_2496);
nand U2591 (N_2591,N_2544,N_2485);
nand U2592 (N_2592,N_2487,N_2525);
and U2593 (N_2593,N_2486,N_2539);
xnor U2594 (N_2594,N_2480,N_2538);
nand U2595 (N_2595,N_2541,N_2498);
xnor U2596 (N_2596,N_2487,N_2547);
xnor U2597 (N_2597,N_2491,N_2476);
xnor U2598 (N_2598,N_2487,N_2541);
or U2599 (N_2599,N_2490,N_2478);
nand U2600 (N_2600,N_2495,N_2531);
and U2601 (N_2601,N_2486,N_2503);
nor U2602 (N_2602,N_2537,N_2547);
xor U2603 (N_2603,N_2493,N_2479);
xnor U2604 (N_2604,N_2506,N_2515);
xor U2605 (N_2605,N_2488,N_2493);
nor U2606 (N_2606,N_2514,N_2505);
or U2607 (N_2607,N_2538,N_2545);
or U2608 (N_2608,N_2476,N_2510);
and U2609 (N_2609,N_2547,N_2481);
xnor U2610 (N_2610,N_2548,N_2523);
nor U2611 (N_2611,N_2514,N_2482);
nand U2612 (N_2612,N_2528,N_2499);
and U2613 (N_2613,N_2548,N_2492);
and U2614 (N_2614,N_2530,N_2517);
and U2615 (N_2615,N_2492,N_2500);
or U2616 (N_2616,N_2514,N_2547);
nand U2617 (N_2617,N_2529,N_2541);
xnor U2618 (N_2618,N_2522,N_2483);
xor U2619 (N_2619,N_2536,N_2500);
and U2620 (N_2620,N_2517,N_2503);
nor U2621 (N_2621,N_2536,N_2537);
xnor U2622 (N_2622,N_2531,N_2526);
xor U2623 (N_2623,N_2544,N_2487);
or U2624 (N_2624,N_2508,N_2500);
or U2625 (N_2625,N_2569,N_2609);
and U2626 (N_2626,N_2617,N_2588);
xnor U2627 (N_2627,N_2599,N_2565);
nand U2628 (N_2628,N_2606,N_2557);
or U2629 (N_2629,N_2594,N_2611);
or U2630 (N_2630,N_2615,N_2579);
xnor U2631 (N_2631,N_2598,N_2624);
nand U2632 (N_2632,N_2576,N_2595);
nor U2633 (N_2633,N_2580,N_2553);
nand U2634 (N_2634,N_2570,N_2613);
nand U2635 (N_2635,N_2550,N_2555);
nor U2636 (N_2636,N_2614,N_2603);
nor U2637 (N_2637,N_2578,N_2558);
nor U2638 (N_2638,N_2593,N_2592);
nand U2639 (N_2639,N_2608,N_2623);
and U2640 (N_2640,N_2559,N_2620);
nor U2641 (N_2641,N_2618,N_2583);
nor U2642 (N_2642,N_2564,N_2590);
xor U2643 (N_2643,N_2556,N_2586);
and U2644 (N_2644,N_2602,N_2622);
nor U2645 (N_2645,N_2577,N_2610);
nand U2646 (N_2646,N_2563,N_2568);
nand U2647 (N_2647,N_2607,N_2596);
xnor U2648 (N_2648,N_2561,N_2619);
and U2649 (N_2649,N_2584,N_2562);
xnor U2650 (N_2650,N_2574,N_2552);
nor U2651 (N_2651,N_2612,N_2591);
nor U2652 (N_2652,N_2621,N_2605);
nor U2653 (N_2653,N_2566,N_2597);
and U2654 (N_2654,N_2573,N_2567);
or U2655 (N_2655,N_2551,N_2581);
or U2656 (N_2656,N_2601,N_2575);
xor U2657 (N_2657,N_2582,N_2554);
and U2658 (N_2658,N_2589,N_2600);
nand U2659 (N_2659,N_2585,N_2604);
nand U2660 (N_2660,N_2560,N_2587);
nand U2661 (N_2661,N_2571,N_2572);
and U2662 (N_2662,N_2616,N_2559);
nand U2663 (N_2663,N_2587,N_2592);
and U2664 (N_2664,N_2587,N_2609);
nor U2665 (N_2665,N_2581,N_2563);
nor U2666 (N_2666,N_2623,N_2605);
xor U2667 (N_2667,N_2605,N_2587);
xor U2668 (N_2668,N_2576,N_2581);
and U2669 (N_2669,N_2613,N_2568);
nand U2670 (N_2670,N_2622,N_2573);
and U2671 (N_2671,N_2560,N_2613);
nor U2672 (N_2672,N_2619,N_2557);
nand U2673 (N_2673,N_2581,N_2607);
nor U2674 (N_2674,N_2598,N_2593);
and U2675 (N_2675,N_2576,N_2555);
nor U2676 (N_2676,N_2584,N_2571);
xor U2677 (N_2677,N_2619,N_2554);
xor U2678 (N_2678,N_2604,N_2564);
nand U2679 (N_2679,N_2574,N_2589);
or U2680 (N_2680,N_2617,N_2620);
xnor U2681 (N_2681,N_2615,N_2554);
xor U2682 (N_2682,N_2557,N_2550);
nor U2683 (N_2683,N_2563,N_2561);
nand U2684 (N_2684,N_2621,N_2609);
xor U2685 (N_2685,N_2550,N_2620);
and U2686 (N_2686,N_2591,N_2578);
and U2687 (N_2687,N_2550,N_2613);
or U2688 (N_2688,N_2582,N_2590);
nand U2689 (N_2689,N_2623,N_2617);
nor U2690 (N_2690,N_2605,N_2603);
nand U2691 (N_2691,N_2586,N_2616);
or U2692 (N_2692,N_2559,N_2560);
or U2693 (N_2693,N_2555,N_2615);
xor U2694 (N_2694,N_2590,N_2611);
xnor U2695 (N_2695,N_2609,N_2565);
nor U2696 (N_2696,N_2595,N_2573);
and U2697 (N_2697,N_2584,N_2577);
or U2698 (N_2698,N_2585,N_2607);
xor U2699 (N_2699,N_2624,N_2582);
nor U2700 (N_2700,N_2692,N_2650);
xnor U2701 (N_2701,N_2670,N_2628);
and U2702 (N_2702,N_2661,N_2643);
nand U2703 (N_2703,N_2696,N_2674);
or U2704 (N_2704,N_2646,N_2651);
or U2705 (N_2705,N_2693,N_2630);
xor U2706 (N_2706,N_2648,N_2633);
or U2707 (N_2707,N_2662,N_2641);
nor U2708 (N_2708,N_2689,N_2697);
nor U2709 (N_2709,N_2672,N_2665);
nand U2710 (N_2710,N_2652,N_2666);
xnor U2711 (N_2711,N_2671,N_2626);
nand U2712 (N_2712,N_2685,N_2656);
and U2713 (N_2713,N_2642,N_2660);
or U2714 (N_2714,N_2635,N_2683);
nor U2715 (N_2715,N_2639,N_2676);
nand U2716 (N_2716,N_2686,N_2659);
nor U2717 (N_2717,N_2644,N_2673);
or U2718 (N_2718,N_2699,N_2679);
nand U2719 (N_2719,N_2636,N_2634);
xor U2720 (N_2720,N_2632,N_2647);
nand U2721 (N_2721,N_2658,N_2677);
and U2722 (N_2722,N_2653,N_2657);
or U2723 (N_2723,N_2654,N_2691);
nor U2724 (N_2724,N_2668,N_2631);
nor U2725 (N_2725,N_2645,N_2682);
xor U2726 (N_2726,N_2684,N_2698);
xor U2727 (N_2727,N_2664,N_2655);
nor U2728 (N_2728,N_2663,N_2629);
nor U2729 (N_2729,N_2625,N_2687);
nor U2730 (N_2730,N_2681,N_2694);
nand U2731 (N_2731,N_2640,N_2667);
nor U2732 (N_2732,N_2680,N_2688);
xnor U2733 (N_2733,N_2678,N_2638);
or U2734 (N_2734,N_2675,N_2627);
xor U2735 (N_2735,N_2649,N_2637);
or U2736 (N_2736,N_2690,N_2695);
nor U2737 (N_2737,N_2669,N_2639);
and U2738 (N_2738,N_2662,N_2682);
and U2739 (N_2739,N_2689,N_2699);
nand U2740 (N_2740,N_2685,N_2652);
and U2741 (N_2741,N_2657,N_2662);
nand U2742 (N_2742,N_2649,N_2628);
nor U2743 (N_2743,N_2685,N_2688);
and U2744 (N_2744,N_2684,N_2632);
xnor U2745 (N_2745,N_2685,N_2628);
and U2746 (N_2746,N_2675,N_2644);
and U2747 (N_2747,N_2685,N_2694);
and U2748 (N_2748,N_2650,N_2664);
nor U2749 (N_2749,N_2625,N_2679);
nor U2750 (N_2750,N_2680,N_2636);
nor U2751 (N_2751,N_2663,N_2635);
nand U2752 (N_2752,N_2687,N_2695);
and U2753 (N_2753,N_2679,N_2688);
nand U2754 (N_2754,N_2699,N_2632);
nor U2755 (N_2755,N_2639,N_2680);
xnor U2756 (N_2756,N_2697,N_2656);
xor U2757 (N_2757,N_2657,N_2692);
xnor U2758 (N_2758,N_2663,N_2653);
and U2759 (N_2759,N_2676,N_2683);
or U2760 (N_2760,N_2632,N_2678);
nor U2761 (N_2761,N_2649,N_2686);
nor U2762 (N_2762,N_2634,N_2669);
nor U2763 (N_2763,N_2639,N_2634);
or U2764 (N_2764,N_2684,N_2664);
and U2765 (N_2765,N_2658,N_2693);
xor U2766 (N_2766,N_2681,N_2687);
xor U2767 (N_2767,N_2681,N_2636);
nor U2768 (N_2768,N_2651,N_2641);
xnor U2769 (N_2769,N_2663,N_2688);
or U2770 (N_2770,N_2660,N_2648);
xor U2771 (N_2771,N_2633,N_2676);
xnor U2772 (N_2772,N_2657,N_2658);
and U2773 (N_2773,N_2646,N_2652);
nand U2774 (N_2774,N_2647,N_2638);
and U2775 (N_2775,N_2751,N_2741);
or U2776 (N_2776,N_2762,N_2709);
nor U2777 (N_2777,N_2712,N_2750);
or U2778 (N_2778,N_2715,N_2745);
and U2779 (N_2779,N_2757,N_2727);
nor U2780 (N_2780,N_2760,N_2702);
nand U2781 (N_2781,N_2763,N_2744);
and U2782 (N_2782,N_2724,N_2737);
nand U2783 (N_2783,N_2768,N_2723);
nor U2784 (N_2784,N_2746,N_2714);
or U2785 (N_2785,N_2710,N_2771);
nand U2786 (N_2786,N_2743,N_2703);
xnor U2787 (N_2787,N_2713,N_2726);
xnor U2788 (N_2788,N_2767,N_2718);
nand U2789 (N_2789,N_2752,N_2704);
nor U2790 (N_2790,N_2774,N_2705);
and U2791 (N_2791,N_2729,N_2761);
nor U2792 (N_2792,N_2730,N_2722);
xnor U2793 (N_2793,N_2749,N_2740);
or U2794 (N_2794,N_2773,N_2748);
xnor U2795 (N_2795,N_2735,N_2765);
xor U2796 (N_2796,N_2711,N_2739);
xor U2797 (N_2797,N_2756,N_2766);
or U2798 (N_2798,N_2755,N_2764);
and U2799 (N_2799,N_2721,N_2725);
nand U2800 (N_2800,N_2728,N_2747);
and U2801 (N_2801,N_2754,N_2758);
nand U2802 (N_2802,N_2708,N_2734);
xnor U2803 (N_2803,N_2753,N_2770);
or U2804 (N_2804,N_2700,N_2759);
and U2805 (N_2805,N_2769,N_2742);
xor U2806 (N_2806,N_2717,N_2772);
xor U2807 (N_2807,N_2701,N_2719);
or U2808 (N_2808,N_2720,N_2733);
xor U2809 (N_2809,N_2706,N_2731);
nor U2810 (N_2810,N_2738,N_2707);
nor U2811 (N_2811,N_2716,N_2736);
nand U2812 (N_2812,N_2732,N_2745);
or U2813 (N_2813,N_2772,N_2767);
and U2814 (N_2814,N_2765,N_2725);
xor U2815 (N_2815,N_2726,N_2723);
nand U2816 (N_2816,N_2734,N_2757);
or U2817 (N_2817,N_2750,N_2724);
nor U2818 (N_2818,N_2722,N_2770);
xor U2819 (N_2819,N_2705,N_2755);
xnor U2820 (N_2820,N_2753,N_2718);
xnor U2821 (N_2821,N_2766,N_2751);
and U2822 (N_2822,N_2723,N_2755);
or U2823 (N_2823,N_2733,N_2726);
nand U2824 (N_2824,N_2719,N_2770);
xnor U2825 (N_2825,N_2766,N_2762);
nor U2826 (N_2826,N_2719,N_2723);
and U2827 (N_2827,N_2758,N_2736);
xnor U2828 (N_2828,N_2709,N_2767);
xor U2829 (N_2829,N_2723,N_2733);
nor U2830 (N_2830,N_2739,N_2760);
and U2831 (N_2831,N_2770,N_2768);
nand U2832 (N_2832,N_2772,N_2749);
xnor U2833 (N_2833,N_2754,N_2763);
and U2834 (N_2834,N_2705,N_2721);
and U2835 (N_2835,N_2743,N_2773);
and U2836 (N_2836,N_2756,N_2736);
nand U2837 (N_2837,N_2766,N_2755);
nand U2838 (N_2838,N_2702,N_2748);
and U2839 (N_2839,N_2764,N_2706);
and U2840 (N_2840,N_2713,N_2717);
and U2841 (N_2841,N_2764,N_2747);
or U2842 (N_2842,N_2742,N_2712);
xnor U2843 (N_2843,N_2761,N_2756);
nor U2844 (N_2844,N_2708,N_2742);
nand U2845 (N_2845,N_2710,N_2705);
or U2846 (N_2846,N_2740,N_2751);
xor U2847 (N_2847,N_2724,N_2744);
and U2848 (N_2848,N_2726,N_2747);
nand U2849 (N_2849,N_2727,N_2718);
or U2850 (N_2850,N_2842,N_2783);
nand U2851 (N_2851,N_2793,N_2816);
nand U2852 (N_2852,N_2841,N_2798);
nand U2853 (N_2853,N_2784,N_2789);
xnor U2854 (N_2854,N_2838,N_2803);
nand U2855 (N_2855,N_2829,N_2827);
or U2856 (N_2856,N_2792,N_2788);
nor U2857 (N_2857,N_2823,N_2817);
nor U2858 (N_2858,N_2795,N_2837);
xnor U2859 (N_2859,N_2797,N_2787);
nor U2860 (N_2860,N_2780,N_2832);
and U2861 (N_2861,N_2848,N_2796);
xor U2862 (N_2862,N_2777,N_2779);
or U2863 (N_2863,N_2794,N_2843);
or U2864 (N_2864,N_2813,N_2775);
and U2865 (N_2865,N_2782,N_2800);
and U2866 (N_2866,N_2812,N_2786);
nand U2867 (N_2867,N_2820,N_2807);
xor U2868 (N_2868,N_2834,N_2825);
nand U2869 (N_2869,N_2845,N_2840);
or U2870 (N_2870,N_2831,N_2804);
or U2871 (N_2871,N_2806,N_2811);
nand U2872 (N_2872,N_2799,N_2822);
nand U2873 (N_2873,N_2828,N_2849);
and U2874 (N_2874,N_2844,N_2821);
or U2875 (N_2875,N_2778,N_2808);
nor U2876 (N_2876,N_2846,N_2785);
xor U2877 (N_2877,N_2802,N_2839);
xnor U2878 (N_2878,N_2781,N_2847);
nor U2879 (N_2879,N_2836,N_2810);
and U2880 (N_2880,N_2835,N_2824);
or U2881 (N_2881,N_2818,N_2801);
and U2882 (N_2882,N_2809,N_2790);
nand U2883 (N_2883,N_2819,N_2805);
or U2884 (N_2884,N_2830,N_2791);
nor U2885 (N_2885,N_2815,N_2826);
nand U2886 (N_2886,N_2776,N_2833);
xnor U2887 (N_2887,N_2814,N_2838);
xor U2888 (N_2888,N_2786,N_2845);
nand U2889 (N_2889,N_2800,N_2831);
and U2890 (N_2890,N_2778,N_2806);
or U2891 (N_2891,N_2786,N_2808);
xor U2892 (N_2892,N_2819,N_2809);
nand U2893 (N_2893,N_2777,N_2798);
nor U2894 (N_2894,N_2839,N_2798);
nor U2895 (N_2895,N_2780,N_2778);
nor U2896 (N_2896,N_2805,N_2848);
and U2897 (N_2897,N_2816,N_2797);
xor U2898 (N_2898,N_2791,N_2808);
nor U2899 (N_2899,N_2839,N_2843);
nor U2900 (N_2900,N_2778,N_2781);
nor U2901 (N_2901,N_2800,N_2848);
nand U2902 (N_2902,N_2842,N_2825);
xnor U2903 (N_2903,N_2787,N_2786);
nor U2904 (N_2904,N_2783,N_2837);
xnor U2905 (N_2905,N_2782,N_2806);
or U2906 (N_2906,N_2831,N_2807);
nor U2907 (N_2907,N_2783,N_2778);
nor U2908 (N_2908,N_2784,N_2788);
xnor U2909 (N_2909,N_2778,N_2795);
nand U2910 (N_2910,N_2780,N_2817);
nand U2911 (N_2911,N_2809,N_2805);
and U2912 (N_2912,N_2835,N_2781);
nand U2913 (N_2913,N_2823,N_2790);
or U2914 (N_2914,N_2837,N_2809);
or U2915 (N_2915,N_2815,N_2817);
nand U2916 (N_2916,N_2797,N_2844);
nand U2917 (N_2917,N_2802,N_2823);
nor U2918 (N_2918,N_2802,N_2836);
or U2919 (N_2919,N_2783,N_2843);
and U2920 (N_2920,N_2839,N_2775);
or U2921 (N_2921,N_2842,N_2793);
nor U2922 (N_2922,N_2817,N_2794);
xnor U2923 (N_2923,N_2821,N_2819);
nand U2924 (N_2924,N_2778,N_2846);
nand U2925 (N_2925,N_2906,N_2888);
and U2926 (N_2926,N_2891,N_2851);
or U2927 (N_2927,N_2870,N_2924);
nand U2928 (N_2928,N_2895,N_2857);
nand U2929 (N_2929,N_2872,N_2879);
xor U2930 (N_2930,N_2860,N_2919);
and U2931 (N_2931,N_2864,N_2877);
and U2932 (N_2932,N_2861,N_2905);
and U2933 (N_2933,N_2865,N_2907);
nand U2934 (N_2934,N_2913,N_2850);
and U2935 (N_2935,N_2887,N_2908);
nand U2936 (N_2936,N_2918,N_2854);
and U2937 (N_2937,N_2896,N_2917);
or U2938 (N_2938,N_2915,N_2890);
and U2939 (N_2939,N_2858,N_2880);
and U2940 (N_2940,N_2892,N_2873);
nor U2941 (N_2941,N_2889,N_2921);
xnor U2942 (N_2942,N_2902,N_2916);
and U2943 (N_2943,N_2867,N_2875);
nor U2944 (N_2944,N_2910,N_2912);
xor U2945 (N_2945,N_2894,N_2904);
xor U2946 (N_2946,N_2874,N_2871);
or U2947 (N_2947,N_2898,N_2881);
xor U2948 (N_2948,N_2901,N_2886);
and U2949 (N_2949,N_2909,N_2862);
or U2950 (N_2950,N_2922,N_2869);
nand U2951 (N_2951,N_2863,N_2893);
nor U2952 (N_2952,N_2920,N_2885);
or U2953 (N_2953,N_2878,N_2853);
or U2954 (N_2954,N_2884,N_2882);
nand U2955 (N_2955,N_2855,N_2923);
nor U2956 (N_2956,N_2866,N_2899);
nor U2957 (N_2957,N_2868,N_2859);
or U2958 (N_2958,N_2883,N_2897);
nand U2959 (N_2959,N_2911,N_2900);
or U2960 (N_2960,N_2914,N_2903);
or U2961 (N_2961,N_2856,N_2852);
xor U2962 (N_2962,N_2876,N_2879);
or U2963 (N_2963,N_2865,N_2885);
and U2964 (N_2964,N_2867,N_2923);
or U2965 (N_2965,N_2917,N_2864);
and U2966 (N_2966,N_2923,N_2921);
and U2967 (N_2967,N_2914,N_2852);
or U2968 (N_2968,N_2883,N_2862);
or U2969 (N_2969,N_2879,N_2917);
nor U2970 (N_2970,N_2873,N_2886);
or U2971 (N_2971,N_2916,N_2880);
and U2972 (N_2972,N_2859,N_2894);
nor U2973 (N_2973,N_2908,N_2862);
nand U2974 (N_2974,N_2869,N_2881);
and U2975 (N_2975,N_2872,N_2878);
or U2976 (N_2976,N_2883,N_2853);
and U2977 (N_2977,N_2892,N_2870);
xnor U2978 (N_2978,N_2870,N_2884);
or U2979 (N_2979,N_2893,N_2867);
or U2980 (N_2980,N_2897,N_2901);
nor U2981 (N_2981,N_2857,N_2912);
xor U2982 (N_2982,N_2892,N_2919);
nor U2983 (N_2983,N_2920,N_2905);
xnor U2984 (N_2984,N_2871,N_2868);
and U2985 (N_2985,N_2892,N_2908);
or U2986 (N_2986,N_2875,N_2886);
nand U2987 (N_2987,N_2893,N_2892);
nor U2988 (N_2988,N_2922,N_2919);
xnor U2989 (N_2989,N_2851,N_2869);
or U2990 (N_2990,N_2905,N_2915);
or U2991 (N_2991,N_2889,N_2884);
nor U2992 (N_2992,N_2924,N_2911);
nand U2993 (N_2993,N_2906,N_2889);
nor U2994 (N_2994,N_2882,N_2864);
xnor U2995 (N_2995,N_2851,N_2878);
or U2996 (N_2996,N_2918,N_2902);
nand U2997 (N_2997,N_2913,N_2864);
nand U2998 (N_2998,N_2862,N_2885);
and U2999 (N_2999,N_2905,N_2907);
nand UO_0 (O_0,N_2963,N_2994);
xnor UO_1 (O_1,N_2979,N_2951);
or UO_2 (O_2,N_2983,N_2950);
and UO_3 (O_3,N_2971,N_2928);
or UO_4 (O_4,N_2936,N_2961);
xnor UO_5 (O_5,N_2930,N_2996);
nor UO_6 (O_6,N_2962,N_2984);
and UO_7 (O_7,N_2932,N_2927);
and UO_8 (O_8,N_2958,N_2954);
nor UO_9 (O_9,N_2943,N_2947);
nand UO_10 (O_10,N_2948,N_2989);
nand UO_11 (O_11,N_2975,N_2973);
nand UO_12 (O_12,N_2997,N_2938);
nor UO_13 (O_13,N_2946,N_2985);
and UO_14 (O_14,N_2926,N_2974);
or UO_15 (O_15,N_2944,N_2978);
and UO_16 (O_16,N_2934,N_2945);
nand UO_17 (O_17,N_2937,N_2941);
and UO_18 (O_18,N_2988,N_2949);
and UO_19 (O_19,N_2929,N_2986);
xnor UO_20 (O_20,N_2955,N_2970);
nor UO_21 (O_21,N_2969,N_2999);
and UO_22 (O_22,N_2931,N_2939);
or UO_23 (O_23,N_2980,N_2991);
xnor UO_24 (O_24,N_2993,N_2953);
and UO_25 (O_25,N_2982,N_2965);
or UO_26 (O_26,N_2981,N_2952);
and UO_27 (O_27,N_2940,N_2964);
nor UO_28 (O_28,N_2968,N_2960);
nor UO_29 (O_29,N_2959,N_2935);
xor UO_30 (O_30,N_2933,N_2987);
xnor UO_31 (O_31,N_2956,N_2977);
nor UO_32 (O_32,N_2995,N_2972);
nor UO_33 (O_33,N_2957,N_2966);
nor UO_34 (O_34,N_2925,N_2992);
xor UO_35 (O_35,N_2998,N_2942);
or UO_36 (O_36,N_2976,N_2990);
or UO_37 (O_37,N_2967,N_2983);
or UO_38 (O_38,N_2936,N_2998);
nand UO_39 (O_39,N_2965,N_2985);
and UO_40 (O_40,N_2994,N_2978);
nor UO_41 (O_41,N_2928,N_2981);
or UO_42 (O_42,N_2988,N_2957);
nand UO_43 (O_43,N_2930,N_2925);
and UO_44 (O_44,N_2981,N_2956);
xor UO_45 (O_45,N_2975,N_2928);
or UO_46 (O_46,N_2946,N_2941);
or UO_47 (O_47,N_2940,N_2933);
nand UO_48 (O_48,N_2972,N_2979);
xor UO_49 (O_49,N_2995,N_2998);
nor UO_50 (O_50,N_2993,N_2951);
xor UO_51 (O_51,N_2994,N_2940);
xor UO_52 (O_52,N_2985,N_2984);
or UO_53 (O_53,N_2941,N_2986);
nand UO_54 (O_54,N_2959,N_2934);
or UO_55 (O_55,N_2939,N_2928);
nor UO_56 (O_56,N_2971,N_2970);
nand UO_57 (O_57,N_2988,N_2987);
xnor UO_58 (O_58,N_2992,N_2984);
and UO_59 (O_59,N_2974,N_2972);
nand UO_60 (O_60,N_2994,N_2936);
xnor UO_61 (O_61,N_2944,N_2969);
nand UO_62 (O_62,N_2985,N_2971);
nor UO_63 (O_63,N_2936,N_2973);
xor UO_64 (O_64,N_2967,N_2995);
and UO_65 (O_65,N_2927,N_2959);
nand UO_66 (O_66,N_2960,N_2952);
xor UO_67 (O_67,N_2945,N_2981);
xnor UO_68 (O_68,N_2987,N_2955);
nor UO_69 (O_69,N_2972,N_2993);
xor UO_70 (O_70,N_2962,N_2925);
and UO_71 (O_71,N_2966,N_2952);
or UO_72 (O_72,N_2947,N_2925);
or UO_73 (O_73,N_2953,N_2967);
and UO_74 (O_74,N_2944,N_2950);
nand UO_75 (O_75,N_2977,N_2984);
nand UO_76 (O_76,N_2981,N_2987);
and UO_77 (O_77,N_2929,N_2944);
nor UO_78 (O_78,N_2988,N_2950);
nand UO_79 (O_79,N_2997,N_2981);
or UO_80 (O_80,N_2927,N_2936);
nor UO_81 (O_81,N_2980,N_2972);
nand UO_82 (O_82,N_2929,N_2930);
and UO_83 (O_83,N_2949,N_2965);
or UO_84 (O_84,N_2968,N_2987);
or UO_85 (O_85,N_2966,N_2938);
nor UO_86 (O_86,N_2931,N_2991);
nand UO_87 (O_87,N_2978,N_2955);
and UO_88 (O_88,N_2994,N_2980);
xor UO_89 (O_89,N_2939,N_2943);
xnor UO_90 (O_90,N_2983,N_2943);
or UO_91 (O_91,N_2925,N_2984);
xor UO_92 (O_92,N_2975,N_2990);
xor UO_93 (O_93,N_2964,N_2928);
or UO_94 (O_94,N_2961,N_2950);
xor UO_95 (O_95,N_2972,N_2936);
and UO_96 (O_96,N_2977,N_2926);
nor UO_97 (O_97,N_2935,N_2976);
xor UO_98 (O_98,N_2954,N_2945);
and UO_99 (O_99,N_2961,N_2981);
nor UO_100 (O_100,N_2966,N_2943);
nand UO_101 (O_101,N_2993,N_2946);
and UO_102 (O_102,N_2949,N_2980);
nand UO_103 (O_103,N_2950,N_2984);
nand UO_104 (O_104,N_2970,N_2947);
nand UO_105 (O_105,N_2947,N_2968);
or UO_106 (O_106,N_2956,N_2965);
and UO_107 (O_107,N_2957,N_2981);
nand UO_108 (O_108,N_2972,N_2941);
nand UO_109 (O_109,N_2958,N_2959);
or UO_110 (O_110,N_2969,N_2983);
and UO_111 (O_111,N_2997,N_2968);
xnor UO_112 (O_112,N_2937,N_2942);
or UO_113 (O_113,N_2981,N_2991);
nand UO_114 (O_114,N_2960,N_2936);
or UO_115 (O_115,N_2927,N_2989);
xnor UO_116 (O_116,N_2945,N_2939);
nand UO_117 (O_117,N_2993,N_2938);
nand UO_118 (O_118,N_2976,N_2998);
or UO_119 (O_119,N_2940,N_2989);
xnor UO_120 (O_120,N_2969,N_2984);
nand UO_121 (O_121,N_2968,N_2939);
and UO_122 (O_122,N_2975,N_2947);
nand UO_123 (O_123,N_2979,N_2944);
or UO_124 (O_124,N_2966,N_2940);
nand UO_125 (O_125,N_2943,N_2960);
xor UO_126 (O_126,N_2946,N_2950);
nor UO_127 (O_127,N_2992,N_2956);
and UO_128 (O_128,N_2944,N_2972);
or UO_129 (O_129,N_2968,N_2932);
and UO_130 (O_130,N_2985,N_2996);
xor UO_131 (O_131,N_2958,N_2951);
or UO_132 (O_132,N_2990,N_2937);
xor UO_133 (O_133,N_2939,N_2996);
and UO_134 (O_134,N_2958,N_2978);
nand UO_135 (O_135,N_2962,N_2993);
or UO_136 (O_136,N_2952,N_2956);
or UO_137 (O_137,N_2946,N_2954);
and UO_138 (O_138,N_2970,N_2941);
and UO_139 (O_139,N_2953,N_2988);
xnor UO_140 (O_140,N_2980,N_2987);
xnor UO_141 (O_141,N_2979,N_2984);
nor UO_142 (O_142,N_2929,N_2997);
nand UO_143 (O_143,N_2986,N_2959);
and UO_144 (O_144,N_2987,N_2943);
xnor UO_145 (O_145,N_2940,N_2988);
nand UO_146 (O_146,N_2935,N_2930);
nor UO_147 (O_147,N_2945,N_2978);
nor UO_148 (O_148,N_2975,N_2959);
xnor UO_149 (O_149,N_2953,N_2930);
xnor UO_150 (O_150,N_2982,N_2974);
nor UO_151 (O_151,N_2925,N_2932);
xnor UO_152 (O_152,N_2973,N_2998);
nor UO_153 (O_153,N_2943,N_2967);
xnor UO_154 (O_154,N_2936,N_2977);
nor UO_155 (O_155,N_2934,N_2975);
nor UO_156 (O_156,N_2961,N_2984);
nand UO_157 (O_157,N_2944,N_2999);
xor UO_158 (O_158,N_2969,N_2998);
and UO_159 (O_159,N_2982,N_2934);
xor UO_160 (O_160,N_2960,N_2955);
nand UO_161 (O_161,N_2928,N_2993);
xnor UO_162 (O_162,N_2971,N_2930);
or UO_163 (O_163,N_2998,N_2949);
xnor UO_164 (O_164,N_2992,N_2930);
xor UO_165 (O_165,N_2933,N_2926);
nand UO_166 (O_166,N_2956,N_2987);
and UO_167 (O_167,N_2985,N_2969);
and UO_168 (O_168,N_2944,N_2928);
xor UO_169 (O_169,N_2956,N_2997);
nand UO_170 (O_170,N_2932,N_2939);
and UO_171 (O_171,N_2975,N_2972);
nand UO_172 (O_172,N_2947,N_2999);
xor UO_173 (O_173,N_2966,N_2937);
nor UO_174 (O_174,N_2994,N_2989);
and UO_175 (O_175,N_2954,N_2974);
xor UO_176 (O_176,N_2980,N_2940);
xor UO_177 (O_177,N_2929,N_2970);
and UO_178 (O_178,N_2938,N_2950);
or UO_179 (O_179,N_2964,N_2929);
and UO_180 (O_180,N_2926,N_2959);
nor UO_181 (O_181,N_2995,N_2945);
xor UO_182 (O_182,N_2925,N_2935);
nand UO_183 (O_183,N_2941,N_2985);
xor UO_184 (O_184,N_2969,N_2982);
nor UO_185 (O_185,N_2947,N_2989);
xnor UO_186 (O_186,N_2981,N_2962);
nand UO_187 (O_187,N_2966,N_2971);
and UO_188 (O_188,N_2968,N_2944);
nand UO_189 (O_189,N_2990,N_2928);
and UO_190 (O_190,N_2965,N_2932);
xor UO_191 (O_191,N_2928,N_2995);
or UO_192 (O_192,N_2988,N_2934);
and UO_193 (O_193,N_2939,N_2941);
or UO_194 (O_194,N_2931,N_2983);
xor UO_195 (O_195,N_2973,N_2976);
nor UO_196 (O_196,N_2954,N_2989);
nor UO_197 (O_197,N_2941,N_2929);
nor UO_198 (O_198,N_2987,N_2945);
and UO_199 (O_199,N_2948,N_2942);
and UO_200 (O_200,N_2973,N_2955);
xnor UO_201 (O_201,N_2989,N_2961);
and UO_202 (O_202,N_2973,N_2970);
nor UO_203 (O_203,N_2972,N_2968);
and UO_204 (O_204,N_2984,N_2933);
xnor UO_205 (O_205,N_2996,N_2969);
or UO_206 (O_206,N_2972,N_2933);
xnor UO_207 (O_207,N_2965,N_2960);
nor UO_208 (O_208,N_2937,N_2961);
nand UO_209 (O_209,N_2991,N_2938);
xor UO_210 (O_210,N_2980,N_2965);
xor UO_211 (O_211,N_2960,N_2962);
nand UO_212 (O_212,N_2956,N_2951);
or UO_213 (O_213,N_2927,N_2957);
nand UO_214 (O_214,N_2992,N_2933);
and UO_215 (O_215,N_2992,N_2971);
nand UO_216 (O_216,N_2972,N_2965);
nor UO_217 (O_217,N_2965,N_2941);
nand UO_218 (O_218,N_2986,N_2975);
or UO_219 (O_219,N_2970,N_2997);
xnor UO_220 (O_220,N_2988,N_2941);
xor UO_221 (O_221,N_2994,N_2969);
xor UO_222 (O_222,N_2978,N_2967);
and UO_223 (O_223,N_2999,N_2967);
nor UO_224 (O_224,N_2955,N_2956);
nand UO_225 (O_225,N_2996,N_2951);
or UO_226 (O_226,N_2998,N_2992);
nand UO_227 (O_227,N_2933,N_2981);
and UO_228 (O_228,N_2926,N_2953);
nor UO_229 (O_229,N_2975,N_2948);
nor UO_230 (O_230,N_2976,N_2969);
or UO_231 (O_231,N_2937,N_2958);
nor UO_232 (O_232,N_2936,N_2979);
nor UO_233 (O_233,N_2994,N_2960);
nor UO_234 (O_234,N_2956,N_2963);
xnor UO_235 (O_235,N_2972,N_2999);
nand UO_236 (O_236,N_2965,N_2988);
nand UO_237 (O_237,N_2965,N_2996);
nor UO_238 (O_238,N_2942,N_2939);
nand UO_239 (O_239,N_2929,N_2977);
nor UO_240 (O_240,N_2980,N_2956);
xnor UO_241 (O_241,N_2990,N_2942);
or UO_242 (O_242,N_2971,N_2993);
nand UO_243 (O_243,N_2966,N_2961);
nand UO_244 (O_244,N_2929,N_2994);
xnor UO_245 (O_245,N_2964,N_2930);
and UO_246 (O_246,N_2955,N_2986);
nor UO_247 (O_247,N_2945,N_2965);
nor UO_248 (O_248,N_2927,N_2977);
or UO_249 (O_249,N_2987,N_2992);
nor UO_250 (O_250,N_2996,N_2950);
nand UO_251 (O_251,N_2942,N_2952);
and UO_252 (O_252,N_2937,N_2928);
and UO_253 (O_253,N_2930,N_2956);
or UO_254 (O_254,N_2941,N_2975);
or UO_255 (O_255,N_2968,N_2953);
xor UO_256 (O_256,N_2927,N_2952);
and UO_257 (O_257,N_2978,N_2937);
or UO_258 (O_258,N_2936,N_2944);
and UO_259 (O_259,N_2961,N_2974);
or UO_260 (O_260,N_2974,N_2958);
and UO_261 (O_261,N_2990,N_2951);
nand UO_262 (O_262,N_2935,N_2977);
and UO_263 (O_263,N_2953,N_2944);
nor UO_264 (O_264,N_2975,N_2976);
nor UO_265 (O_265,N_2967,N_2938);
xor UO_266 (O_266,N_2970,N_2942);
nor UO_267 (O_267,N_2933,N_2982);
and UO_268 (O_268,N_2944,N_2956);
xnor UO_269 (O_269,N_2973,N_2974);
nand UO_270 (O_270,N_2957,N_2956);
or UO_271 (O_271,N_2990,N_2962);
nor UO_272 (O_272,N_2964,N_2981);
nor UO_273 (O_273,N_2983,N_2975);
nand UO_274 (O_274,N_2984,N_2954);
nor UO_275 (O_275,N_2926,N_2987);
nand UO_276 (O_276,N_2927,N_2962);
nand UO_277 (O_277,N_2929,N_2928);
xor UO_278 (O_278,N_2974,N_2955);
or UO_279 (O_279,N_2980,N_2976);
nand UO_280 (O_280,N_2926,N_2964);
and UO_281 (O_281,N_2985,N_2959);
nand UO_282 (O_282,N_2968,N_2952);
or UO_283 (O_283,N_2926,N_2948);
xnor UO_284 (O_284,N_2929,N_2960);
nand UO_285 (O_285,N_2930,N_2982);
nor UO_286 (O_286,N_2977,N_2940);
and UO_287 (O_287,N_2960,N_2975);
xnor UO_288 (O_288,N_2965,N_2975);
nor UO_289 (O_289,N_2930,N_2975);
and UO_290 (O_290,N_2933,N_2930);
nor UO_291 (O_291,N_2958,N_2942);
nand UO_292 (O_292,N_2931,N_2938);
and UO_293 (O_293,N_2932,N_2967);
or UO_294 (O_294,N_2940,N_2937);
nand UO_295 (O_295,N_2970,N_2934);
or UO_296 (O_296,N_2936,N_2988);
nand UO_297 (O_297,N_2968,N_2931);
or UO_298 (O_298,N_2999,N_2963);
nand UO_299 (O_299,N_2962,N_2974);
nand UO_300 (O_300,N_2953,N_2975);
nand UO_301 (O_301,N_2946,N_2944);
and UO_302 (O_302,N_2985,N_2953);
or UO_303 (O_303,N_2950,N_2964);
nand UO_304 (O_304,N_2979,N_2971);
and UO_305 (O_305,N_2958,N_2931);
nand UO_306 (O_306,N_2967,N_2958);
or UO_307 (O_307,N_2992,N_2957);
xor UO_308 (O_308,N_2993,N_2926);
xor UO_309 (O_309,N_2974,N_2949);
xor UO_310 (O_310,N_2974,N_2968);
nand UO_311 (O_311,N_2932,N_2969);
xnor UO_312 (O_312,N_2935,N_2993);
and UO_313 (O_313,N_2925,N_2960);
xor UO_314 (O_314,N_2945,N_2985);
and UO_315 (O_315,N_2975,N_2974);
nor UO_316 (O_316,N_2987,N_2939);
nand UO_317 (O_317,N_2997,N_2989);
or UO_318 (O_318,N_2963,N_2985);
and UO_319 (O_319,N_2961,N_2929);
xor UO_320 (O_320,N_2983,N_2925);
or UO_321 (O_321,N_2927,N_2940);
or UO_322 (O_322,N_2953,N_2948);
nor UO_323 (O_323,N_2964,N_2986);
or UO_324 (O_324,N_2947,N_2997);
or UO_325 (O_325,N_2989,N_2960);
nand UO_326 (O_326,N_2938,N_2981);
nand UO_327 (O_327,N_2953,N_2982);
nor UO_328 (O_328,N_2942,N_2975);
or UO_329 (O_329,N_2960,N_2982);
or UO_330 (O_330,N_2967,N_2929);
and UO_331 (O_331,N_2970,N_2999);
nand UO_332 (O_332,N_2937,N_2993);
nor UO_333 (O_333,N_2970,N_2993);
nor UO_334 (O_334,N_2925,N_2997);
xor UO_335 (O_335,N_2943,N_2993);
nor UO_336 (O_336,N_2925,N_2928);
or UO_337 (O_337,N_2976,N_2991);
nand UO_338 (O_338,N_2971,N_2987);
nor UO_339 (O_339,N_2931,N_2956);
xnor UO_340 (O_340,N_2964,N_2993);
or UO_341 (O_341,N_2985,N_2974);
nand UO_342 (O_342,N_2927,N_2976);
nor UO_343 (O_343,N_2930,N_2997);
nor UO_344 (O_344,N_2981,N_2963);
and UO_345 (O_345,N_2940,N_2942);
xor UO_346 (O_346,N_2964,N_2953);
nand UO_347 (O_347,N_2937,N_2981);
xnor UO_348 (O_348,N_2949,N_2963);
nand UO_349 (O_349,N_2996,N_2984);
nor UO_350 (O_350,N_2955,N_2942);
nor UO_351 (O_351,N_2988,N_2935);
nor UO_352 (O_352,N_2943,N_2975);
nor UO_353 (O_353,N_2983,N_2964);
or UO_354 (O_354,N_2992,N_2960);
nand UO_355 (O_355,N_2991,N_2959);
nand UO_356 (O_356,N_2986,N_2928);
and UO_357 (O_357,N_2963,N_2935);
or UO_358 (O_358,N_2941,N_2990);
and UO_359 (O_359,N_2929,N_2990);
xor UO_360 (O_360,N_2929,N_2958);
xnor UO_361 (O_361,N_2950,N_2940);
nand UO_362 (O_362,N_2960,N_2931);
nand UO_363 (O_363,N_2965,N_2957);
nand UO_364 (O_364,N_2944,N_2926);
and UO_365 (O_365,N_2997,N_2964);
or UO_366 (O_366,N_2959,N_2973);
or UO_367 (O_367,N_2984,N_2943);
nand UO_368 (O_368,N_2974,N_2941);
or UO_369 (O_369,N_2994,N_2965);
and UO_370 (O_370,N_2925,N_2950);
nand UO_371 (O_371,N_2977,N_2979);
nor UO_372 (O_372,N_2997,N_2967);
and UO_373 (O_373,N_2935,N_2933);
nand UO_374 (O_374,N_2945,N_2976);
or UO_375 (O_375,N_2952,N_2935);
or UO_376 (O_376,N_2967,N_2931);
xor UO_377 (O_377,N_2979,N_2976);
nand UO_378 (O_378,N_2965,N_2936);
xnor UO_379 (O_379,N_2993,N_2927);
nand UO_380 (O_380,N_2928,N_2946);
nand UO_381 (O_381,N_2977,N_2975);
and UO_382 (O_382,N_2947,N_2958);
nand UO_383 (O_383,N_2980,N_2990);
or UO_384 (O_384,N_2948,N_2941);
or UO_385 (O_385,N_2955,N_2976);
nand UO_386 (O_386,N_2960,N_2985);
and UO_387 (O_387,N_2928,N_2980);
nor UO_388 (O_388,N_2929,N_2946);
nand UO_389 (O_389,N_2961,N_2968);
nor UO_390 (O_390,N_2992,N_2979);
or UO_391 (O_391,N_2984,N_2929);
nor UO_392 (O_392,N_2926,N_2934);
and UO_393 (O_393,N_2995,N_2984);
or UO_394 (O_394,N_2959,N_2974);
nor UO_395 (O_395,N_2996,N_2963);
nor UO_396 (O_396,N_2968,N_2996);
or UO_397 (O_397,N_2942,N_2959);
xnor UO_398 (O_398,N_2934,N_2995);
or UO_399 (O_399,N_2931,N_2994);
nor UO_400 (O_400,N_2934,N_2987);
and UO_401 (O_401,N_2976,N_2964);
nor UO_402 (O_402,N_2968,N_2959);
and UO_403 (O_403,N_2986,N_2998);
and UO_404 (O_404,N_2977,N_2992);
and UO_405 (O_405,N_2994,N_2971);
xnor UO_406 (O_406,N_2988,N_2995);
nand UO_407 (O_407,N_2989,N_2943);
and UO_408 (O_408,N_2997,N_2962);
or UO_409 (O_409,N_2958,N_2938);
or UO_410 (O_410,N_2994,N_2972);
nor UO_411 (O_411,N_2940,N_2944);
or UO_412 (O_412,N_2937,N_2955);
and UO_413 (O_413,N_2989,N_2983);
and UO_414 (O_414,N_2942,N_2945);
nor UO_415 (O_415,N_2995,N_2973);
xor UO_416 (O_416,N_2995,N_2986);
nand UO_417 (O_417,N_2968,N_2930);
nand UO_418 (O_418,N_2945,N_2968);
xnor UO_419 (O_419,N_2932,N_2974);
nor UO_420 (O_420,N_2990,N_2977);
xor UO_421 (O_421,N_2947,N_2988);
xor UO_422 (O_422,N_2976,N_2960);
or UO_423 (O_423,N_2980,N_2958);
nor UO_424 (O_424,N_2951,N_2938);
nand UO_425 (O_425,N_2939,N_2986);
nand UO_426 (O_426,N_2963,N_2995);
xnor UO_427 (O_427,N_2939,N_2953);
or UO_428 (O_428,N_2943,N_2976);
nand UO_429 (O_429,N_2967,N_2994);
nor UO_430 (O_430,N_2983,N_2951);
nor UO_431 (O_431,N_2959,N_2957);
and UO_432 (O_432,N_2983,N_2945);
nor UO_433 (O_433,N_2928,N_2970);
or UO_434 (O_434,N_2948,N_2973);
and UO_435 (O_435,N_2930,N_2980);
and UO_436 (O_436,N_2970,N_2930);
xor UO_437 (O_437,N_2952,N_2995);
and UO_438 (O_438,N_2967,N_2952);
or UO_439 (O_439,N_2929,N_2996);
and UO_440 (O_440,N_2992,N_2934);
xor UO_441 (O_441,N_2968,N_2981);
nand UO_442 (O_442,N_2960,N_2979);
xnor UO_443 (O_443,N_2925,N_2977);
nor UO_444 (O_444,N_2974,N_2964);
xnor UO_445 (O_445,N_2952,N_2945);
nand UO_446 (O_446,N_2978,N_2927);
or UO_447 (O_447,N_2954,N_2944);
and UO_448 (O_448,N_2955,N_2975);
or UO_449 (O_449,N_2984,N_2994);
nor UO_450 (O_450,N_2967,N_2945);
and UO_451 (O_451,N_2993,N_2930);
nor UO_452 (O_452,N_2950,N_2987);
nand UO_453 (O_453,N_2951,N_2937);
nand UO_454 (O_454,N_2937,N_2985);
nand UO_455 (O_455,N_2939,N_2962);
or UO_456 (O_456,N_2934,N_2940);
and UO_457 (O_457,N_2966,N_2925);
nand UO_458 (O_458,N_2984,N_2991);
nor UO_459 (O_459,N_2985,N_2950);
and UO_460 (O_460,N_2954,N_2927);
nor UO_461 (O_461,N_2970,N_2945);
nand UO_462 (O_462,N_2929,N_2976);
nor UO_463 (O_463,N_2972,N_2986);
nor UO_464 (O_464,N_2957,N_2953);
xnor UO_465 (O_465,N_2925,N_2959);
nand UO_466 (O_466,N_2938,N_2956);
nand UO_467 (O_467,N_2957,N_2996);
and UO_468 (O_468,N_2994,N_2930);
nand UO_469 (O_469,N_2935,N_2926);
nor UO_470 (O_470,N_2943,N_2980);
and UO_471 (O_471,N_2970,N_2977);
xor UO_472 (O_472,N_2975,N_2958);
xnor UO_473 (O_473,N_2926,N_2976);
and UO_474 (O_474,N_2970,N_2932);
and UO_475 (O_475,N_2981,N_2965);
nand UO_476 (O_476,N_2999,N_2932);
and UO_477 (O_477,N_2948,N_2974);
or UO_478 (O_478,N_2939,N_2976);
xnor UO_479 (O_479,N_2998,N_2957);
or UO_480 (O_480,N_2969,N_2989);
and UO_481 (O_481,N_2981,N_2996);
or UO_482 (O_482,N_2970,N_2927);
nand UO_483 (O_483,N_2991,N_2972);
and UO_484 (O_484,N_2987,N_2935);
nor UO_485 (O_485,N_2947,N_2941);
nor UO_486 (O_486,N_2947,N_2948);
and UO_487 (O_487,N_2944,N_2958);
nand UO_488 (O_488,N_2971,N_2960);
nand UO_489 (O_489,N_2984,N_2946);
or UO_490 (O_490,N_2943,N_2988);
and UO_491 (O_491,N_2983,N_2996);
nor UO_492 (O_492,N_2982,N_2976);
xnor UO_493 (O_493,N_2985,N_2943);
or UO_494 (O_494,N_2985,N_2995);
nand UO_495 (O_495,N_2977,N_2946);
nand UO_496 (O_496,N_2962,N_2940);
or UO_497 (O_497,N_2975,N_2933);
xor UO_498 (O_498,N_2966,N_2959);
nor UO_499 (O_499,N_2941,N_2933);
endmodule