module basic_750_5000_1000_10_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_123,In_531);
or U1 (N_1,In_708,In_299);
nand U2 (N_2,In_29,In_518);
xnor U3 (N_3,In_167,In_651);
or U4 (N_4,In_185,In_241);
and U5 (N_5,In_196,In_364);
and U6 (N_6,In_13,In_749);
nand U7 (N_7,In_469,In_347);
xnor U8 (N_8,In_346,In_394);
nor U9 (N_9,In_319,In_546);
xnor U10 (N_10,In_431,In_204);
and U11 (N_11,In_164,In_127);
or U12 (N_12,In_214,In_344);
and U13 (N_13,In_149,In_609);
and U14 (N_14,In_624,In_338);
nand U15 (N_15,In_371,In_544);
nand U16 (N_16,In_705,In_276);
or U17 (N_17,In_361,In_331);
xnor U18 (N_18,In_390,In_577);
nor U19 (N_19,In_242,In_408);
and U20 (N_20,In_144,In_535);
xor U21 (N_21,In_122,In_261);
xor U22 (N_22,In_367,In_16);
nand U23 (N_23,In_666,In_642);
xnor U24 (N_24,In_124,In_567);
or U25 (N_25,In_262,In_215);
or U26 (N_26,In_86,In_505);
nand U27 (N_27,In_31,In_125);
or U28 (N_28,In_66,In_359);
and U29 (N_29,In_304,In_42);
nor U30 (N_30,In_392,In_134);
nor U31 (N_31,In_640,In_676);
xor U32 (N_32,In_418,In_322);
nor U33 (N_33,In_480,In_298);
nor U34 (N_34,In_73,In_499);
xor U35 (N_35,In_184,In_207);
nand U36 (N_36,In_658,In_107);
nand U37 (N_37,In_571,In_530);
and U38 (N_38,In_404,In_316);
and U39 (N_39,In_349,In_477);
xor U40 (N_40,In_116,In_324);
nand U41 (N_41,In_712,In_443);
xnor U42 (N_42,In_140,In_22);
or U43 (N_43,In_686,In_630);
nand U44 (N_44,In_46,In_635);
xor U45 (N_45,In_377,In_746);
nand U46 (N_46,In_447,In_315);
nand U47 (N_47,In_70,In_636);
or U48 (N_48,In_694,In_381);
or U49 (N_49,In_35,In_129);
and U50 (N_50,In_8,In_374);
nand U51 (N_51,In_646,In_0);
xor U52 (N_52,In_274,In_728);
or U53 (N_53,In_258,In_368);
or U54 (N_54,In_14,In_409);
xnor U55 (N_55,In_603,In_78);
and U56 (N_56,In_251,In_667);
nor U57 (N_57,In_302,In_143);
nand U58 (N_58,In_497,In_202);
or U59 (N_59,In_87,In_51);
nand U60 (N_60,In_575,In_190);
and U61 (N_61,In_662,In_482);
nand U62 (N_62,In_405,In_427);
or U63 (N_63,In_463,In_697);
xnor U64 (N_64,In_247,In_74);
and U65 (N_65,In_132,In_539);
and U66 (N_66,In_583,In_528);
or U67 (N_67,In_365,In_645);
nand U68 (N_68,In_668,In_740);
xor U69 (N_69,In_552,In_732);
or U70 (N_70,In_714,In_600);
or U71 (N_71,In_200,In_388);
or U72 (N_72,In_451,In_648);
nand U73 (N_73,In_62,In_201);
nand U74 (N_74,In_428,In_286);
nand U75 (N_75,In_7,In_594);
or U76 (N_76,In_671,In_300);
and U77 (N_77,In_317,In_227);
and U78 (N_78,In_67,In_513);
or U79 (N_79,In_681,In_734);
xnor U80 (N_80,In_456,In_631);
xnor U81 (N_81,In_670,In_586);
nor U82 (N_82,In_432,In_63);
xnor U83 (N_83,In_267,In_611);
nor U84 (N_84,In_5,In_625);
nor U85 (N_85,In_543,In_578);
nand U86 (N_86,In_706,In_395);
and U87 (N_87,In_101,In_506);
and U88 (N_88,In_689,In_3);
nand U89 (N_89,In_613,In_389);
and U90 (N_90,In_277,In_503);
or U91 (N_91,In_680,In_584);
and U92 (N_92,In_393,In_188);
and U93 (N_93,In_342,In_145);
or U94 (N_94,In_717,In_20);
nand U95 (N_95,In_629,In_307);
xor U96 (N_96,In_382,In_357);
or U97 (N_97,In_555,In_688);
and U98 (N_98,In_399,In_695);
and U99 (N_99,In_118,In_68);
nor U100 (N_100,In_417,In_446);
and U101 (N_101,In_572,In_454);
or U102 (N_102,In_654,In_219);
and U103 (N_103,In_719,In_605);
xor U104 (N_104,In_549,In_351);
xor U105 (N_105,In_11,In_142);
nand U106 (N_106,In_736,In_425);
xor U107 (N_107,In_103,In_72);
xnor U108 (N_108,In_228,In_633);
or U109 (N_109,In_474,In_453);
or U110 (N_110,In_353,In_157);
xor U111 (N_111,In_702,In_58);
nor U112 (N_112,In_147,In_71);
or U113 (N_113,In_591,In_641);
nand U114 (N_114,In_362,In_327);
and U115 (N_115,In_181,In_398);
nor U116 (N_116,In_683,In_461);
or U117 (N_117,In_108,In_486);
nand U118 (N_118,In_37,In_450);
nor U119 (N_119,In_597,In_715);
nor U120 (N_120,In_69,In_672);
or U121 (N_121,In_507,In_604);
and U122 (N_122,In_28,In_356);
nor U123 (N_123,In_363,In_592);
and U124 (N_124,In_350,In_311);
and U125 (N_125,In_239,In_560);
xor U126 (N_126,In_310,In_253);
and U127 (N_127,In_156,In_358);
xor U128 (N_128,In_150,In_723);
nor U129 (N_129,In_730,In_266);
nor U130 (N_130,In_523,In_620);
xnor U131 (N_131,In_64,In_509);
nand U132 (N_132,In_339,In_162);
xor U133 (N_133,In_55,In_334);
nand U134 (N_134,In_401,In_81);
nand U135 (N_135,In_738,In_716);
and U136 (N_136,In_91,In_416);
xor U137 (N_137,In_268,In_386);
nor U138 (N_138,In_669,In_95);
xor U139 (N_139,In_722,In_644);
or U140 (N_140,In_380,In_516);
xnor U141 (N_141,In_547,In_225);
and U142 (N_142,In_257,In_550);
nand U143 (N_143,In_429,In_387);
and U144 (N_144,In_490,In_366);
nand U145 (N_145,In_25,In_403);
nor U146 (N_146,In_665,In_186);
xor U147 (N_147,In_26,In_245);
nor U148 (N_148,In_218,In_385);
nor U149 (N_149,In_643,In_442);
and U150 (N_150,In_36,In_481);
nand U151 (N_151,In_301,In_373);
and U152 (N_152,In_685,In_663);
nand U153 (N_153,In_527,In_626);
nand U154 (N_154,In_551,In_472);
xnor U155 (N_155,In_97,In_287);
nor U156 (N_156,In_90,In_284);
nor U157 (N_157,In_83,In_158);
xor U158 (N_158,In_45,In_522);
xor U159 (N_159,In_121,In_698);
or U160 (N_160,In_397,In_565);
or U161 (N_161,In_606,In_440);
or U162 (N_162,In_217,In_47);
or U163 (N_163,In_462,In_283);
and U164 (N_164,In_569,In_588);
or U165 (N_165,In_660,In_153);
nor U166 (N_166,In_313,In_554);
xor U167 (N_167,In_294,In_263);
nand U168 (N_168,In_271,In_556);
nor U169 (N_169,In_93,In_748);
or U170 (N_170,In_514,In_508);
xnor U171 (N_171,In_109,In_79);
or U172 (N_172,In_724,In_98);
nor U173 (N_173,In_264,In_136);
nand U174 (N_174,In_259,In_59);
or U175 (N_175,In_618,In_690);
nand U176 (N_176,In_265,In_308);
nand U177 (N_177,In_92,In_691);
or U178 (N_178,In_221,In_407);
nand U179 (N_179,In_273,In_306);
or U180 (N_180,In_329,In_104);
nor U181 (N_181,In_573,In_384);
nor U182 (N_182,In_203,In_410);
xnor U183 (N_183,In_146,In_130);
and U184 (N_184,In_400,In_293);
and U185 (N_185,In_234,In_413);
and U186 (N_186,In_320,In_296);
nand U187 (N_187,In_679,In_585);
xnor U188 (N_188,In_187,In_449);
nor U189 (N_189,In_524,In_89);
and U190 (N_190,In_436,In_693);
and U191 (N_191,In_568,In_532);
or U192 (N_192,In_370,In_65);
nand U193 (N_193,In_533,In_161);
and U194 (N_194,In_488,In_209);
nor U195 (N_195,In_198,In_521);
nand U196 (N_196,In_598,In_699);
or U197 (N_197,In_468,In_191);
nand U198 (N_198,In_735,In_737);
xor U199 (N_199,In_484,In_321);
or U200 (N_200,In_17,In_421);
nor U201 (N_201,In_593,In_742);
xnor U202 (N_202,In_542,In_458);
and U203 (N_203,In_510,In_580);
or U204 (N_204,In_475,In_275);
nand U205 (N_205,In_733,In_595);
or U206 (N_206,In_673,In_596);
nor U207 (N_207,In_312,In_619);
and U208 (N_208,In_457,In_525);
and U209 (N_209,In_163,In_652);
and U210 (N_210,In_341,In_171);
or U211 (N_211,In_232,In_330);
nor U212 (N_212,In_113,In_402);
and U213 (N_213,In_529,In_56);
xnor U214 (N_214,In_224,In_272);
nor U215 (N_215,In_479,In_117);
nor U216 (N_216,In_169,In_376);
nor U217 (N_217,In_6,In_623);
xor U218 (N_218,In_700,In_483);
or U219 (N_219,In_415,In_659);
or U220 (N_220,In_574,In_195);
xor U221 (N_221,In_430,In_119);
and U222 (N_222,In_372,In_570);
and U223 (N_223,In_355,In_682);
nand U224 (N_224,In_411,In_696);
nand U225 (N_225,In_229,In_177);
nor U226 (N_226,In_725,In_538);
nand U227 (N_227,In_709,In_289);
or U228 (N_228,In_206,In_563);
nand U229 (N_229,In_57,In_579);
xor U230 (N_230,In_561,In_53);
nor U231 (N_231,In_664,In_435);
nand U232 (N_232,In_137,In_281);
or U233 (N_233,In_419,In_581);
and U234 (N_234,In_32,In_614);
nand U235 (N_235,In_343,In_291);
nand U236 (N_236,In_328,In_303);
or U237 (N_237,In_33,In_194);
and U238 (N_238,In_455,In_154);
nand U239 (N_239,In_470,In_621);
nand U240 (N_240,In_718,In_498);
or U241 (N_241,In_212,In_236);
nand U242 (N_242,In_354,In_332);
xor U243 (N_243,In_88,In_80);
nand U244 (N_244,In_174,In_617);
xor U245 (N_245,In_216,In_54);
and U246 (N_246,In_517,In_496);
or U247 (N_247,In_34,In_205);
or U248 (N_248,In_238,In_512);
xnor U249 (N_249,In_340,In_152);
and U250 (N_250,In_106,In_348);
or U251 (N_251,In_445,In_622);
nand U252 (N_252,In_252,In_237);
xnor U253 (N_253,In_255,In_278);
xnor U254 (N_254,In_471,In_48);
and U255 (N_255,In_165,In_27);
or U256 (N_256,In_60,In_260);
and U257 (N_257,In_433,In_638);
and U258 (N_258,In_396,In_444);
or U259 (N_259,In_39,In_40);
or U260 (N_260,In_323,In_138);
or U261 (N_261,In_222,In_473);
and U262 (N_262,In_540,In_412);
or U263 (N_263,In_230,In_30);
and U264 (N_264,In_710,In_459);
or U265 (N_265,In_305,In_352);
nor U266 (N_266,In_434,In_548);
nand U267 (N_267,In_96,In_170);
nand U268 (N_268,In_131,In_383);
nand U269 (N_269,In_254,In_420);
or U270 (N_270,In_628,In_369);
or U271 (N_271,In_173,In_82);
xnor U272 (N_272,In_279,In_166);
nand U273 (N_273,In_692,In_422);
and U274 (N_274,In_52,In_295);
nand U275 (N_275,In_4,In_661);
xnor U276 (N_276,In_677,In_208);
xor U277 (N_277,In_511,In_495);
or U278 (N_278,In_183,In_391);
or U279 (N_279,In_41,In_582);
or U280 (N_280,In_678,In_378);
and U281 (N_281,In_500,In_707);
nand U282 (N_282,In_112,In_494);
nand U283 (N_283,In_423,In_337);
or U284 (N_284,In_211,In_151);
nand U285 (N_285,In_438,In_375);
and U286 (N_286,In_178,In_210);
nand U287 (N_287,In_49,In_314);
nand U288 (N_288,In_126,In_610);
or U289 (N_289,In_226,In_44);
nand U290 (N_290,In_128,In_135);
xor U291 (N_291,In_587,In_657);
or U292 (N_292,In_612,In_487);
nor U293 (N_293,In_545,In_50);
nor U294 (N_294,In_566,In_231);
nor U295 (N_295,In_179,In_223);
and U296 (N_296,In_288,In_290);
and U297 (N_297,In_465,In_493);
nor U298 (N_298,In_192,In_720);
or U299 (N_299,In_627,In_655);
xnor U300 (N_300,In_674,In_590);
xor U301 (N_301,In_256,In_703);
or U302 (N_302,In_526,In_406);
nor U303 (N_303,In_653,In_537);
nand U304 (N_304,In_285,In_77);
and U305 (N_305,In_325,In_269);
and U306 (N_306,In_250,In_249);
nor U307 (N_307,In_489,In_309);
or U308 (N_308,In_426,In_75);
nand U309 (N_309,In_602,In_704);
nand U310 (N_310,In_564,In_12);
xor U311 (N_311,In_485,In_467);
xnor U312 (N_312,In_713,In_85);
nand U313 (N_313,In_19,In_159);
and U314 (N_314,In_632,In_9);
nor U315 (N_315,In_244,In_637);
or U316 (N_316,In_1,In_197);
or U317 (N_317,In_133,In_414);
and U318 (N_318,In_248,In_94);
nand U319 (N_319,In_105,In_519);
nor U320 (N_320,In_476,In_326);
nand U321 (N_321,In_448,In_739);
nand U322 (N_322,In_727,In_711);
and U323 (N_323,In_634,In_437);
and U324 (N_324,In_684,In_649);
and U325 (N_325,In_647,In_460);
nor U326 (N_326,In_576,In_452);
nand U327 (N_327,In_155,In_559);
nor U328 (N_328,In_160,In_18);
or U329 (N_329,In_84,In_336);
or U330 (N_330,In_541,In_189);
xor U331 (N_331,In_168,In_120);
and U332 (N_332,In_515,In_536);
xor U333 (N_333,In_360,In_608);
or U334 (N_334,In_491,In_193);
and U335 (N_335,In_199,In_607);
nor U336 (N_336,In_558,In_172);
xor U337 (N_337,In_599,In_318);
or U338 (N_338,In_182,In_701);
nor U339 (N_339,In_100,In_99);
xor U340 (N_340,In_333,In_520);
nor U341 (N_341,In_61,In_464);
and U342 (N_342,In_639,In_675);
or U343 (N_343,In_745,In_43);
and U344 (N_344,In_741,In_141);
and U345 (N_345,In_478,In_424);
nor U346 (N_346,In_656,In_601);
nand U347 (N_347,In_282,In_726);
and U348 (N_348,In_114,In_270);
nor U349 (N_349,In_115,In_102);
or U350 (N_350,In_687,In_492);
xor U351 (N_351,In_379,In_246);
nand U352 (N_352,In_233,In_501);
or U353 (N_353,In_76,In_297);
or U354 (N_354,In_345,In_615);
and U355 (N_355,In_213,In_466);
or U356 (N_356,In_553,In_721);
nand U357 (N_357,In_24,In_504);
nor U358 (N_358,In_441,In_439);
xor U359 (N_359,In_562,In_589);
nor U360 (N_360,In_729,In_38);
and U361 (N_361,In_15,In_111);
nand U362 (N_362,In_650,In_731);
xor U363 (N_363,In_10,In_175);
or U364 (N_364,In_21,In_176);
or U365 (N_365,In_148,In_280);
or U366 (N_366,In_23,In_139);
xnor U367 (N_367,In_335,In_616);
nor U368 (N_368,In_502,In_243);
and U369 (N_369,In_747,In_743);
xnor U370 (N_370,In_744,In_557);
nor U371 (N_371,In_110,In_2);
or U372 (N_372,In_235,In_240);
or U373 (N_373,In_180,In_292);
nand U374 (N_374,In_534,In_220);
and U375 (N_375,In_308,In_299);
nor U376 (N_376,In_293,In_227);
xnor U377 (N_377,In_438,In_105);
nand U378 (N_378,In_243,In_248);
xnor U379 (N_379,In_625,In_204);
nor U380 (N_380,In_600,In_498);
nand U381 (N_381,In_23,In_305);
nor U382 (N_382,In_507,In_399);
nor U383 (N_383,In_135,In_559);
and U384 (N_384,In_546,In_744);
or U385 (N_385,In_328,In_210);
xor U386 (N_386,In_440,In_667);
and U387 (N_387,In_438,In_705);
xnor U388 (N_388,In_5,In_310);
and U389 (N_389,In_17,In_274);
or U390 (N_390,In_178,In_346);
nand U391 (N_391,In_127,In_439);
xor U392 (N_392,In_104,In_97);
nand U393 (N_393,In_711,In_569);
nor U394 (N_394,In_659,In_30);
nand U395 (N_395,In_33,In_251);
nor U396 (N_396,In_616,In_512);
nor U397 (N_397,In_61,In_238);
or U398 (N_398,In_456,In_136);
and U399 (N_399,In_698,In_267);
xnor U400 (N_400,In_84,In_417);
xnor U401 (N_401,In_234,In_641);
xnor U402 (N_402,In_650,In_612);
xnor U403 (N_403,In_320,In_551);
nand U404 (N_404,In_455,In_384);
or U405 (N_405,In_223,In_38);
xor U406 (N_406,In_489,In_340);
nor U407 (N_407,In_515,In_382);
or U408 (N_408,In_28,In_572);
or U409 (N_409,In_35,In_726);
nand U410 (N_410,In_677,In_696);
or U411 (N_411,In_334,In_106);
xnor U412 (N_412,In_681,In_539);
nand U413 (N_413,In_320,In_610);
nand U414 (N_414,In_729,In_634);
nand U415 (N_415,In_177,In_300);
xnor U416 (N_416,In_271,In_717);
xor U417 (N_417,In_409,In_729);
or U418 (N_418,In_514,In_643);
or U419 (N_419,In_648,In_185);
or U420 (N_420,In_461,In_172);
nor U421 (N_421,In_542,In_200);
and U422 (N_422,In_72,In_694);
nor U423 (N_423,In_254,In_288);
or U424 (N_424,In_476,In_288);
nor U425 (N_425,In_684,In_162);
and U426 (N_426,In_520,In_36);
and U427 (N_427,In_78,In_469);
nand U428 (N_428,In_644,In_311);
or U429 (N_429,In_743,In_500);
xnor U430 (N_430,In_244,In_37);
nor U431 (N_431,In_245,In_403);
and U432 (N_432,In_604,In_366);
nor U433 (N_433,In_356,In_675);
xor U434 (N_434,In_92,In_312);
nor U435 (N_435,In_421,In_107);
and U436 (N_436,In_713,In_458);
xnor U437 (N_437,In_466,In_154);
or U438 (N_438,In_124,In_104);
or U439 (N_439,In_485,In_413);
nor U440 (N_440,In_563,In_651);
and U441 (N_441,In_581,In_456);
xnor U442 (N_442,In_447,In_209);
nand U443 (N_443,In_430,In_369);
nand U444 (N_444,In_77,In_162);
or U445 (N_445,In_77,In_120);
nand U446 (N_446,In_281,In_550);
and U447 (N_447,In_392,In_380);
xor U448 (N_448,In_94,In_289);
nor U449 (N_449,In_173,In_521);
nand U450 (N_450,In_511,In_567);
xnor U451 (N_451,In_277,In_596);
nor U452 (N_452,In_494,In_43);
xnor U453 (N_453,In_482,In_330);
xnor U454 (N_454,In_563,In_725);
or U455 (N_455,In_101,In_219);
nand U456 (N_456,In_473,In_314);
or U457 (N_457,In_442,In_518);
and U458 (N_458,In_27,In_411);
or U459 (N_459,In_480,In_125);
nor U460 (N_460,In_434,In_359);
and U461 (N_461,In_633,In_525);
nand U462 (N_462,In_316,In_592);
nor U463 (N_463,In_745,In_317);
and U464 (N_464,In_497,In_33);
nor U465 (N_465,In_434,In_612);
and U466 (N_466,In_435,In_136);
nand U467 (N_467,In_125,In_714);
or U468 (N_468,In_240,In_699);
nor U469 (N_469,In_604,In_128);
or U470 (N_470,In_153,In_648);
and U471 (N_471,In_464,In_352);
nand U472 (N_472,In_418,In_200);
nand U473 (N_473,In_526,In_163);
nor U474 (N_474,In_443,In_366);
and U475 (N_475,In_325,In_164);
xnor U476 (N_476,In_298,In_281);
nor U477 (N_477,In_231,In_629);
nor U478 (N_478,In_266,In_682);
nor U479 (N_479,In_96,In_77);
nor U480 (N_480,In_632,In_413);
and U481 (N_481,In_364,In_255);
and U482 (N_482,In_635,In_137);
xor U483 (N_483,In_368,In_624);
and U484 (N_484,In_312,In_630);
nor U485 (N_485,In_313,In_636);
nand U486 (N_486,In_372,In_289);
or U487 (N_487,In_38,In_181);
nand U488 (N_488,In_103,In_496);
xor U489 (N_489,In_376,In_483);
nand U490 (N_490,In_532,In_308);
and U491 (N_491,In_423,In_145);
xor U492 (N_492,In_457,In_559);
nor U493 (N_493,In_687,In_505);
nor U494 (N_494,In_398,In_449);
nand U495 (N_495,In_479,In_307);
and U496 (N_496,In_735,In_510);
nor U497 (N_497,In_137,In_523);
and U498 (N_498,In_184,In_227);
xnor U499 (N_499,In_483,In_556);
or U500 (N_500,N_249,N_135);
or U501 (N_501,N_468,N_293);
or U502 (N_502,N_403,N_40);
nor U503 (N_503,N_482,N_383);
nand U504 (N_504,N_147,N_319);
nand U505 (N_505,N_220,N_240);
and U506 (N_506,N_156,N_88);
nor U507 (N_507,N_51,N_260);
or U508 (N_508,N_358,N_284);
nor U509 (N_509,N_212,N_334);
and U510 (N_510,N_456,N_400);
nor U511 (N_511,N_179,N_31);
nand U512 (N_512,N_194,N_496);
nand U513 (N_513,N_123,N_155);
xor U514 (N_514,N_364,N_470);
nor U515 (N_515,N_116,N_306);
nor U516 (N_516,N_238,N_375);
or U517 (N_517,N_111,N_114);
and U518 (N_518,N_148,N_366);
nand U519 (N_519,N_22,N_187);
xnor U520 (N_520,N_303,N_413);
xnor U521 (N_521,N_416,N_139);
and U522 (N_522,N_232,N_140);
xnor U523 (N_523,N_189,N_442);
nand U524 (N_524,N_133,N_426);
nor U525 (N_525,N_9,N_34);
and U526 (N_526,N_425,N_331);
and U527 (N_527,N_85,N_8);
or U528 (N_528,N_107,N_268);
nor U529 (N_529,N_377,N_126);
and U530 (N_530,N_429,N_439);
nand U531 (N_531,N_1,N_11);
nand U532 (N_532,N_10,N_76);
nand U533 (N_533,N_282,N_315);
nand U534 (N_534,N_195,N_452);
nor U535 (N_535,N_352,N_33);
nor U536 (N_536,N_373,N_237);
and U537 (N_537,N_428,N_415);
xnor U538 (N_538,N_271,N_231);
and U539 (N_539,N_349,N_494);
or U540 (N_540,N_171,N_433);
nand U541 (N_541,N_69,N_41);
and U542 (N_542,N_434,N_299);
and U543 (N_543,N_185,N_124);
nand U544 (N_544,N_368,N_499);
xor U545 (N_545,N_45,N_217);
nor U546 (N_546,N_44,N_322);
xnor U547 (N_547,N_226,N_233);
xor U548 (N_548,N_254,N_42);
or U549 (N_549,N_277,N_180);
or U550 (N_550,N_317,N_491);
or U551 (N_551,N_227,N_363);
nand U552 (N_552,N_167,N_294);
or U553 (N_553,N_298,N_168);
or U554 (N_554,N_308,N_206);
and U555 (N_555,N_460,N_432);
or U556 (N_556,N_351,N_242);
or U557 (N_557,N_336,N_380);
nor U558 (N_558,N_483,N_143);
nand U559 (N_559,N_64,N_26);
and U560 (N_560,N_28,N_37);
or U561 (N_561,N_125,N_229);
or U562 (N_562,N_371,N_411);
and U563 (N_563,N_455,N_175);
nand U564 (N_564,N_397,N_49);
nand U565 (N_565,N_150,N_134);
or U566 (N_566,N_130,N_492);
or U567 (N_567,N_484,N_287);
nand U568 (N_568,N_63,N_154);
and U569 (N_569,N_197,N_296);
nand U570 (N_570,N_39,N_493);
nand U571 (N_571,N_477,N_219);
and U572 (N_572,N_313,N_353);
or U573 (N_573,N_53,N_476);
nor U574 (N_574,N_98,N_407);
or U575 (N_575,N_398,N_487);
nor U576 (N_576,N_208,N_58);
and U577 (N_577,N_152,N_142);
or U578 (N_578,N_326,N_486);
or U579 (N_579,N_356,N_186);
and U580 (N_580,N_448,N_77);
or U581 (N_581,N_246,N_419);
or U582 (N_582,N_279,N_228);
and U583 (N_583,N_52,N_191);
xor U584 (N_584,N_381,N_214);
nor U585 (N_585,N_245,N_19);
or U586 (N_586,N_234,N_113);
xor U587 (N_587,N_91,N_5);
nor U588 (N_588,N_17,N_347);
nor U589 (N_589,N_221,N_89);
nor U590 (N_590,N_387,N_138);
nor U591 (N_591,N_418,N_193);
or U592 (N_592,N_144,N_330);
nor U593 (N_593,N_263,N_151);
and U594 (N_594,N_164,N_471);
and U595 (N_595,N_201,N_361);
nor U596 (N_596,N_101,N_280);
and U597 (N_597,N_2,N_90);
xnor U598 (N_598,N_444,N_318);
or U599 (N_599,N_408,N_23);
nand U600 (N_600,N_495,N_273);
xor U601 (N_601,N_78,N_461);
xnor U602 (N_602,N_86,N_178);
or U603 (N_603,N_244,N_390);
or U604 (N_604,N_256,N_43);
nand U605 (N_605,N_73,N_176);
nor U606 (N_606,N_97,N_223);
nand U607 (N_607,N_453,N_0);
xor U608 (N_608,N_420,N_56);
and U609 (N_609,N_445,N_320);
xnor U610 (N_610,N_382,N_146);
nand U611 (N_611,N_261,N_203);
and U612 (N_612,N_450,N_474);
nand U613 (N_613,N_436,N_396);
nand U614 (N_614,N_462,N_100);
nand U615 (N_615,N_110,N_96);
nand U616 (N_616,N_449,N_61);
or U617 (N_617,N_278,N_106);
and U618 (N_618,N_286,N_57);
nand U619 (N_619,N_82,N_222);
nor U620 (N_620,N_129,N_490);
nand U621 (N_621,N_332,N_198);
nand U622 (N_622,N_20,N_120);
or U623 (N_623,N_71,N_392);
xor U624 (N_624,N_327,N_250);
or U625 (N_625,N_301,N_230);
xnor U626 (N_626,N_414,N_102);
and U627 (N_627,N_479,N_16);
or U628 (N_628,N_405,N_183);
xnor U629 (N_629,N_160,N_344);
nor U630 (N_630,N_269,N_87);
or U631 (N_631,N_399,N_35);
nand U632 (N_632,N_281,N_410);
xnor U633 (N_633,N_328,N_367);
xnor U634 (N_634,N_47,N_264);
nand U635 (N_635,N_55,N_431);
nand U636 (N_636,N_362,N_141);
or U637 (N_637,N_182,N_115);
xor U638 (N_638,N_170,N_412);
xnor U639 (N_639,N_14,N_12);
nand U640 (N_640,N_18,N_497);
xor U641 (N_641,N_437,N_251);
nand U642 (N_642,N_108,N_172);
xnor U643 (N_643,N_307,N_473);
nor U644 (N_644,N_389,N_395);
and U645 (N_645,N_488,N_13);
nand U646 (N_646,N_127,N_66);
xor U647 (N_647,N_209,N_59);
xnor U648 (N_648,N_354,N_292);
nand U649 (N_649,N_118,N_481);
xnor U650 (N_650,N_443,N_162);
nand U651 (N_651,N_104,N_302);
nand U652 (N_652,N_153,N_454);
and U653 (N_653,N_266,N_70);
xnor U654 (N_654,N_252,N_159);
nor U655 (N_655,N_305,N_321);
and U656 (N_656,N_391,N_360);
and U657 (N_657,N_489,N_385);
and U658 (N_658,N_333,N_190);
and U659 (N_659,N_80,N_25);
and U660 (N_660,N_215,N_99);
and U661 (N_661,N_235,N_128);
xor U662 (N_662,N_285,N_157);
nand U663 (N_663,N_169,N_247);
xnor U664 (N_664,N_204,N_446);
nor U665 (N_665,N_15,N_457);
xor U666 (N_666,N_469,N_374);
and U667 (N_667,N_253,N_174);
or U668 (N_668,N_424,N_402);
xor U669 (N_669,N_430,N_74);
nand U670 (N_670,N_6,N_467);
xor U671 (N_671,N_283,N_378);
xnor U672 (N_672,N_92,N_4);
or U673 (N_673,N_192,N_346);
and U674 (N_674,N_105,N_472);
or U675 (N_675,N_376,N_259);
nand U676 (N_676,N_357,N_29);
nand U677 (N_677,N_136,N_36);
or U678 (N_678,N_65,N_236);
nor U679 (N_679,N_161,N_304);
and U680 (N_680,N_276,N_475);
nor U681 (N_681,N_54,N_316);
nand U682 (N_682,N_274,N_365);
xnor U683 (N_683,N_337,N_24);
and U684 (N_684,N_132,N_7);
nand U685 (N_685,N_173,N_498);
and U686 (N_686,N_211,N_216);
nand U687 (N_687,N_325,N_202);
nand U688 (N_688,N_350,N_478);
and U689 (N_689,N_289,N_267);
or U690 (N_690,N_81,N_84);
or U691 (N_691,N_388,N_288);
nor U692 (N_692,N_213,N_137);
xnor U693 (N_693,N_393,N_441);
nor U694 (N_694,N_465,N_205);
and U695 (N_695,N_341,N_210);
and U696 (N_696,N_394,N_158);
xor U697 (N_697,N_94,N_75);
nor U698 (N_698,N_409,N_163);
nand U699 (N_699,N_272,N_48);
nand U700 (N_700,N_359,N_340);
nand U701 (N_701,N_262,N_112);
nor U702 (N_702,N_68,N_435);
xnor U703 (N_703,N_239,N_335);
nand U704 (N_704,N_311,N_270);
nor U705 (N_705,N_27,N_386);
xnor U706 (N_706,N_314,N_458);
and U707 (N_707,N_248,N_438);
xnor U708 (N_708,N_323,N_83);
and U709 (N_709,N_427,N_255);
or U710 (N_710,N_451,N_50);
xor U711 (N_711,N_224,N_309);
xnor U712 (N_712,N_370,N_67);
and U713 (N_713,N_463,N_384);
xnor U714 (N_714,N_131,N_200);
or U715 (N_715,N_422,N_46);
xnor U716 (N_716,N_149,N_21);
nand U717 (N_717,N_121,N_312);
or U718 (N_718,N_3,N_345);
xnor U719 (N_719,N_404,N_257);
and U720 (N_720,N_275,N_95);
nor U721 (N_721,N_79,N_348);
nor U722 (N_722,N_339,N_166);
xnor U723 (N_723,N_485,N_372);
or U724 (N_724,N_480,N_225);
xnor U725 (N_725,N_184,N_290);
nand U726 (N_726,N_300,N_177);
xor U727 (N_727,N_103,N_329);
or U728 (N_728,N_165,N_417);
and U729 (N_729,N_423,N_342);
or U730 (N_730,N_406,N_421);
nor U731 (N_731,N_199,N_379);
nor U732 (N_732,N_145,N_459);
nor U733 (N_733,N_369,N_243);
nand U734 (N_734,N_258,N_188);
nor U735 (N_735,N_32,N_310);
and U736 (N_736,N_265,N_109);
and U737 (N_737,N_122,N_241);
nor U738 (N_738,N_93,N_297);
nor U739 (N_739,N_295,N_218);
and U740 (N_740,N_38,N_62);
or U741 (N_741,N_291,N_440);
and U742 (N_742,N_466,N_447);
nor U743 (N_743,N_401,N_181);
nor U744 (N_744,N_338,N_196);
nor U745 (N_745,N_355,N_207);
and U746 (N_746,N_464,N_72);
and U747 (N_747,N_117,N_343);
xnor U748 (N_748,N_60,N_119);
nor U749 (N_749,N_324,N_30);
or U750 (N_750,N_328,N_6);
or U751 (N_751,N_179,N_468);
and U752 (N_752,N_466,N_15);
nor U753 (N_753,N_10,N_431);
and U754 (N_754,N_446,N_161);
nand U755 (N_755,N_37,N_355);
xor U756 (N_756,N_209,N_395);
xor U757 (N_757,N_335,N_303);
nand U758 (N_758,N_275,N_277);
and U759 (N_759,N_120,N_144);
nand U760 (N_760,N_35,N_397);
nor U761 (N_761,N_473,N_54);
and U762 (N_762,N_497,N_245);
nand U763 (N_763,N_209,N_230);
xor U764 (N_764,N_484,N_147);
or U765 (N_765,N_13,N_282);
nand U766 (N_766,N_135,N_229);
xor U767 (N_767,N_51,N_254);
nor U768 (N_768,N_464,N_19);
and U769 (N_769,N_322,N_249);
nor U770 (N_770,N_220,N_422);
and U771 (N_771,N_470,N_316);
and U772 (N_772,N_263,N_472);
nand U773 (N_773,N_222,N_385);
and U774 (N_774,N_36,N_75);
xnor U775 (N_775,N_404,N_65);
xnor U776 (N_776,N_481,N_52);
nor U777 (N_777,N_381,N_118);
or U778 (N_778,N_268,N_370);
and U779 (N_779,N_11,N_292);
xnor U780 (N_780,N_407,N_459);
and U781 (N_781,N_428,N_251);
or U782 (N_782,N_291,N_23);
nand U783 (N_783,N_157,N_135);
nor U784 (N_784,N_493,N_99);
nor U785 (N_785,N_431,N_14);
or U786 (N_786,N_422,N_167);
nand U787 (N_787,N_190,N_48);
or U788 (N_788,N_333,N_259);
and U789 (N_789,N_264,N_355);
xnor U790 (N_790,N_414,N_151);
and U791 (N_791,N_91,N_44);
xor U792 (N_792,N_233,N_179);
nand U793 (N_793,N_316,N_100);
or U794 (N_794,N_166,N_201);
nand U795 (N_795,N_102,N_160);
and U796 (N_796,N_329,N_451);
xnor U797 (N_797,N_339,N_27);
or U798 (N_798,N_225,N_5);
and U799 (N_799,N_481,N_448);
nor U800 (N_800,N_116,N_313);
and U801 (N_801,N_85,N_165);
or U802 (N_802,N_446,N_392);
nand U803 (N_803,N_427,N_244);
nor U804 (N_804,N_492,N_106);
nand U805 (N_805,N_240,N_469);
nand U806 (N_806,N_82,N_15);
nor U807 (N_807,N_248,N_157);
nor U808 (N_808,N_430,N_157);
nor U809 (N_809,N_96,N_24);
nand U810 (N_810,N_271,N_194);
and U811 (N_811,N_428,N_373);
and U812 (N_812,N_136,N_174);
and U813 (N_813,N_459,N_487);
or U814 (N_814,N_306,N_124);
nand U815 (N_815,N_455,N_52);
xor U816 (N_816,N_452,N_409);
nand U817 (N_817,N_233,N_192);
nand U818 (N_818,N_410,N_325);
and U819 (N_819,N_243,N_197);
nand U820 (N_820,N_154,N_134);
nor U821 (N_821,N_307,N_138);
or U822 (N_822,N_263,N_260);
nand U823 (N_823,N_76,N_471);
nand U824 (N_824,N_146,N_246);
or U825 (N_825,N_244,N_209);
nor U826 (N_826,N_423,N_337);
and U827 (N_827,N_226,N_242);
nand U828 (N_828,N_65,N_88);
xor U829 (N_829,N_183,N_417);
nor U830 (N_830,N_258,N_12);
or U831 (N_831,N_113,N_494);
xor U832 (N_832,N_4,N_357);
and U833 (N_833,N_35,N_39);
and U834 (N_834,N_292,N_269);
and U835 (N_835,N_167,N_438);
or U836 (N_836,N_377,N_84);
nand U837 (N_837,N_205,N_497);
and U838 (N_838,N_162,N_20);
nor U839 (N_839,N_388,N_497);
nor U840 (N_840,N_335,N_421);
xnor U841 (N_841,N_303,N_55);
nand U842 (N_842,N_312,N_278);
nand U843 (N_843,N_411,N_481);
nor U844 (N_844,N_53,N_396);
nand U845 (N_845,N_378,N_208);
or U846 (N_846,N_221,N_271);
and U847 (N_847,N_472,N_122);
nor U848 (N_848,N_59,N_160);
or U849 (N_849,N_387,N_173);
nor U850 (N_850,N_243,N_426);
or U851 (N_851,N_23,N_335);
xnor U852 (N_852,N_24,N_185);
nor U853 (N_853,N_341,N_216);
xor U854 (N_854,N_24,N_103);
and U855 (N_855,N_27,N_224);
nor U856 (N_856,N_144,N_446);
and U857 (N_857,N_113,N_419);
nor U858 (N_858,N_39,N_74);
xor U859 (N_859,N_300,N_145);
or U860 (N_860,N_24,N_397);
and U861 (N_861,N_257,N_354);
nand U862 (N_862,N_368,N_404);
xor U863 (N_863,N_233,N_411);
or U864 (N_864,N_78,N_211);
and U865 (N_865,N_329,N_148);
nand U866 (N_866,N_123,N_273);
and U867 (N_867,N_168,N_311);
xnor U868 (N_868,N_47,N_310);
nor U869 (N_869,N_326,N_125);
or U870 (N_870,N_366,N_242);
nand U871 (N_871,N_371,N_433);
or U872 (N_872,N_386,N_231);
and U873 (N_873,N_348,N_27);
or U874 (N_874,N_229,N_156);
nor U875 (N_875,N_193,N_233);
and U876 (N_876,N_175,N_104);
nor U877 (N_877,N_362,N_285);
nand U878 (N_878,N_403,N_451);
or U879 (N_879,N_305,N_20);
nor U880 (N_880,N_157,N_273);
nor U881 (N_881,N_81,N_200);
or U882 (N_882,N_116,N_182);
and U883 (N_883,N_410,N_330);
or U884 (N_884,N_403,N_325);
xnor U885 (N_885,N_249,N_126);
xor U886 (N_886,N_57,N_22);
or U887 (N_887,N_456,N_44);
xnor U888 (N_888,N_435,N_130);
nor U889 (N_889,N_381,N_430);
nand U890 (N_890,N_447,N_449);
and U891 (N_891,N_120,N_461);
xor U892 (N_892,N_392,N_240);
xor U893 (N_893,N_258,N_98);
xor U894 (N_894,N_419,N_479);
xor U895 (N_895,N_226,N_321);
or U896 (N_896,N_235,N_193);
or U897 (N_897,N_445,N_318);
nand U898 (N_898,N_339,N_334);
nand U899 (N_899,N_275,N_435);
nor U900 (N_900,N_19,N_446);
nor U901 (N_901,N_479,N_457);
xnor U902 (N_902,N_267,N_427);
or U903 (N_903,N_22,N_156);
or U904 (N_904,N_347,N_393);
and U905 (N_905,N_285,N_136);
or U906 (N_906,N_97,N_417);
or U907 (N_907,N_152,N_410);
and U908 (N_908,N_90,N_258);
or U909 (N_909,N_453,N_47);
nand U910 (N_910,N_487,N_195);
nand U911 (N_911,N_186,N_477);
xnor U912 (N_912,N_252,N_366);
nor U913 (N_913,N_447,N_9);
nand U914 (N_914,N_411,N_142);
nor U915 (N_915,N_173,N_75);
nor U916 (N_916,N_499,N_195);
xnor U917 (N_917,N_281,N_186);
or U918 (N_918,N_28,N_358);
and U919 (N_919,N_22,N_259);
nand U920 (N_920,N_231,N_113);
nor U921 (N_921,N_33,N_349);
xnor U922 (N_922,N_346,N_1);
xnor U923 (N_923,N_174,N_1);
nand U924 (N_924,N_284,N_46);
and U925 (N_925,N_54,N_398);
or U926 (N_926,N_329,N_55);
or U927 (N_927,N_26,N_220);
nor U928 (N_928,N_279,N_385);
or U929 (N_929,N_397,N_59);
nor U930 (N_930,N_403,N_51);
nand U931 (N_931,N_150,N_257);
or U932 (N_932,N_125,N_1);
nand U933 (N_933,N_118,N_394);
nand U934 (N_934,N_247,N_199);
xnor U935 (N_935,N_132,N_223);
and U936 (N_936,N_191,N_128);
and U937 (N_937,N_69,N_319);
nand U938 (N_938,N_322,N_342);
and U939 (N_939,N_266,N_75);
nand U940 (N_940,N_208,N_390);
and U941 (N_941,N_198,N_236);
or U942 (N_942,N_393,N_333);
nand U943 (N_943,N_389,N_407);
nand U944 (N_944,N_28,N_226);
and U945 (N_945,N_448,N_58);
nand U946 (N_946,N_7,N_22);
nor U947 (N_947,N_155,N_239);
or U948 (N_948,N_413,N_29);
nand U949 (N_949,N_63,N_189);
xnor U950 (N_950,N_26,N_271);
and U951 (N_951,N_144,N_25);
xor U952 (N_952,N_457,N_328);
nor U953 (N_953,N_196,N_49);
or U954 (N_954,N_263,N_63);
nor U955 (N_955,N_114,N_315);
xor U956 (N_956,N_219,N_9);
nor U957 (N_957,N_77,N_213);
nor U958 (N_958,N_250,N_251);
or U959 (N_959,N_232,N_496);
nand U960 (N_960,N_212,N_282);
nand U961 (N_961,N_42,N_437);
nand U962 (N_962,N_283,N_195);
nand U963 (N_963,N_333,N_26);
and U964 (N_964,N_248,N_406);
xor U965 (N_965,N_55,N_413);
nand U966 (N_966,N_364,N_201);
or U967 (N_967,N_154,N_281);
nand U968 (N_968,N_212,N_232);
nand U969 (N_969,N_174,N_243);
or U970 (N_970,N_486,N_50);
nand U971 (N_971,N_191,N_110);
or U972 (N_972,N_10,N_479);
xor U973 (N_973,N_328,N_107);
nor U974 (N_974,N_206,N_135);
nor U975 (N_975,N_93,N_401);
nor U976 (N_976,N_311,N_226);
nor U977 (N_977,N_74,N_181);
nand U978 (N_978,N_52,N_65);
and U979 (N_979,N_104,N_352);
nor U980 (N_980,N_134,N_315);
or U981 (N_981,N_152,N_30);
or U982 (N_982,N_175,N_7);
nand U983 (N_983,N_451,N_334);
xor U984 (N_984,N_464,N_50);
nor U985 (N_985,N_135,N_31);
xor U986 (N_986,N_63,N_58);
or U987 (N_987,N_152,N_27);
or U988 (N_988,N_177,N_454);
nand U989 (N_989,N_387,N_46);
nor U990 (N_990,N_203,N_88);
nor U991 (N_991,N_122,N_435);
or U992 (N_992,N_485,N_237);
and U993 (N_993,N_189,N_263);
or U994 (N_994,N_175,N_486);
nor U995 (N_995,N_57,N_474);
and U996 (N_996,N_292,N_22);
nand U997 (N_997,N_129,N_20);
and U998 (N_998,N_11,N_400);
nand U999 (N_999,N_203,N_366);
xnor U1000 (N_1000,N_944,N_608);
or U1001 (N_1001,N_807,N_664);
or U1002 (N_1002,N_739,N_534);
or U1003 (N_1003,N_956,N_886);
or U1004 (N_1004,N_697,N_943);
xor U1005 (N_1005,N_659,N_824);
or U1006 (N_1006,N_724,N_636);
and U1007 (N_1007,N_989,N_634);
nor U1008 (N_1008,N_810,N_707);
and U1009 (N_1009,N_730,N_996);
or U1010 (N_1010,N_966,N_702);
and U1011 (N_1011,N_889,N_825);
nor U1012 (N_1012,N_885,N_502);
xnor U1013 (N_1013,N_635,N_945);
or U1014 (N_1014,N_786,N_642);
and U1015 (N_1015,N_540,N_699);
nand U1016 (N_1016,N_719,N_839);
or U1017 (N_1017,N_845,N_892);
nor U1018 (N_1018,N_621,N_958);
or U1019 (N_1019,N_765,N_775);
nand U1020 (N_1020,N_850,N_604);
nor U1021 (N_1021,N_916,N_803);
or U1022 (N_1022,N_651,N_675);
nand U1023 (N_1023,N_835,N_998);
nand U1024 (N_1024,N_605,N_843);
nor U1025 (N_1025,N_617,N_537);
nand U1026 (N_1026,N_883,N_564);
nand U1027 (N_1027,N_973,N_764);
or U1028 (N_1028,N_787,N_682);
and U1029 (N_1029,N_976,N_923);
or U1030 (N_1030,N_523,N_901);
or U1031 (N_1031,N_586,N_629);
or U1032 (N_1032,N_934,N_967);
and U1033 (N_1033,N_565,N_587);
and U1034 (N_1034,N_832,N_551);
or U1035 (N_1035,N_672,N_789);
and U1036 (N_1036,N_962,N_828);
xnor U1037 (N_1037,N_653,N_715);
or U1038 (N_1038,N_741,N_555);
and U1039 (N_1039,N_802,N_578);
nand U1040 (N_1040,N_869,N_785);
nor U1041 (N_1041,N_530,N_856);
nand U1042 (N_1042,N_870,N_566);
nor U1043 (N_1043,N_932,N_581);
xnor U1044 (N_1044,N_713,N_718);
or U1045 (N_1045,N_854,N_696);
xnor U1046 (N_1046,N_960,N_689);
nand U1047 (N_1047,N_861,N_773);
nor U1048 (N_1048,N_542,N_595);
nor U1049 (N_1049,N_947,N_622);
nand U1050 (N_1050,N_738,N_579);
nand U1051 (N_1051,N_931,N_763);
and U1052 (N_1052,N_805,N_701);
and U1053 (N_1053,N_691,N_897);
and U1054 (N_1054,N_625,N_830);
and U1055 (N_1055,N_860,N_920);
xor U1056 (N_1056,N_567,N_937);
nand U1057 (N_1057,N_986,N_746);
nor U1058 (N_1058,N_528,N_949);
xnor U1059 (N_1059,N_547,N_592);
nor U1060 (N_1060,N_583,N_779);
xnor U1061 (N_1061,N_544,N_903);
and U1062 (N_1062,N_982,N_710);
or U1063 (N_1063,N_933,N_504);
nand U1064 (N_1064,N_963,N_831);
nand U1065 (N_1065,N_519,N_631);
and U1066 (N_1066,N_533,N_574);
xnor U1067 (N_1067,N_543,N_569);
nor U1068 (N_1068,N_965,N_927);
and U1069 (N_1069,N_538,N_734);
nor U1070 (N_1070,N_692,N_921);
nor U1071 (N_1071,N_627,N_859);
or U1072 (N_1072,N_576,N_979);
nand U1073 (N_1073,N_902,N_667);
nand U1074 (N_1074,N_541,N_950);
xor U1075 (N_1075,N_532,N_905);
and U1076 (N_1076,N_733,N_737);
or U1077 (N_1077,N_771,N_836);
and U1078 (N_1078,N_848,N_925);
nand U1079 (N_1079,N_678,N_681);
nor U1080 (N_1080,N_872,N_972);
or U1081 (N_1081,N_633,N_874);
nand U1082 (N_1082,N_751,N_781);
and U1083 (N_1083,N_614,N_968);
and U1084 (N_1084,N_849,N_558);
nor U1085 (N_1085,N_964,N_703);
xor U1086 (N_1086,N_743,N_646);
and U1087 (N_1087,N_783,N_990);
nand U1088 (N_1088,N_855,N_680);
nor U1089 (N_1089,N_811,N_531);
nand U1090 (N_1090,N_975,N_539);
xnor U1091 (N_1091,N_938,N_673);
and U1092 (N_1092,N_939,N_988);
nand U1093 (N_1093,N_603,N_914);
xor U1094 (N_1094,N_732,N_597);
and U1095 (N_1095,N_762,N_961);
nor U1096 (N_1096,N_879,N_900);
and U1097 (N_1097,N_750,N_867);
nor U1098 (N_1098,N_669,N_591);
nand U1099 (N_1099,N_782,N_767);
or U1100 (N_1100,N_521,N_674);
nor U1101 (N_1101,N_744,N_705);
xor U1102 (N_1102,N_690,N_501);
xnor U1103 (N_1103,N_894,N_709);
or U1104 (N_1104,N_814,N_818);
nor U1105 (N_1105,N_694,N_816);
xnor U1106 (N_1106,N_609,N_550);
or U1107 (N_1107,N_777,N_817);
nand U1108 (N_1108,N_891,N_645);
and U1109 (N_1109,N_992,N_655);
or U1110 (N_1110,N_529,N_695);
nor U1111 (N_1111,N_842,N_808);
xnor U1112 (N_1112,N_522,N_761);
and U1113 (N_1113,N_557,N_899);
and U1114 (N_1114,N_735,N_506);
nand U1115 (N_1115,N_729,N_706);
nand U1116 (N_1116,N_955,N_615);
and U1117 (N_1117,N_772,N_599);
nor U1118 (N_1118,N_797,N_851);
nor U1119 (N_1119,N_866,N_520);
and U1120 (N_1120,N_708,N_670);
xor U1121 (N_1121,N_942,N_554);
or U1122 (N_1122,N_910,N_712);
nand U1123 (N_1123,N_784,N_693);
nor U1124 (N_1124,N_753,N_776);
nor U1125 (N_1125,N_602,N_985);
nand U1126 (N_1126,N_868,N_911);
nor U1127 (N_1127,N_740,N_895);
nor U1128 (N_1128,N_683,N_801);
and U1129 (N_1129,N_560,N_823);
or U1130 (N_1130,N_676,N_846);
xor U1131 (N_1131,N_507,N_527);
or U1132 (N_1132,N_954,N_589);
or U1133 (N_1133,N_745,N_619);
nor U1134 (N_1134,N_834,N_953);
and U1135 (N_1135,N_686,N_922);
nand U1136 (N_1136,N_688,N_728);
xnor U1137 (N_1137,N_600,N_928);
or U1138 (N_1138,N_721,N_873);
or U1139 (N_1139,N_665,N_793);
xnor U1140 (N_1140,N_511,N_754);
nor U1141 (N_1141,N_720,N_607);
nand U1142 (N_1142,N_598,N_628);
and U1143 (N_1143,N_684,N_572);
or U1144 (N_1144,N_881,N_585);
nor U1145 (N_1145,N_792,N_906);
nor U1146 (N_1146,N_563,N_515);
nand U1147 (N_1147,N_637,N_747);
or U1148 (N_1148,N_644,N_526);
nand U1149 (N_1149,N_875,N_912);
nor U1150 (N_1150,N_641,N_913);
nand U1151 (N_1151,N_704,N_510);
nor U1152 (N_1152,N_829,N_601);
and U1153 (N_1153,N_853,N_714);
xnor U1154 (N_1154,N_974,N_623);
nand U1155 (N_1155,N_584,N_833);
and U1156 (N_1156,N_545,N_656);
and U1157 (N_1157,N_577,N_896);
nor U1158 (N_1158,N_722,N_748);
xnor U1159 (N_1159,N_984,N_610);
or U1160 (N_1160,N_878,N_582);
nand U1161 (N_1161,N_821,N_716);
and U1162 (N_1162,N_919,N_756);
nand U1163 (N_1163,N_970,N_685);
or U1164 (N_1164,N_915,N_800);
nand U1165 (N_1165,N_759,N_909);
or U1166 (N_1166,N_994,N_838);
xor U1167 (N_1167,N_570,N_826);
nand U1168 (N_1168,N_804,N_559);
and U1169 (N_1169,N_749,N_649);
nor U1170 (N_1170,N_500,N_661);
and U1171 (N_1171,N_790,N_995);
and U1172 (N_1172,N_548,N_606);
xor U1173 (N_1173,N_671,N_798);
xor U1174 (N_1174,N_711,N_679);
xnor U1175 (N_1175,N_552,N_788);
nand U1176 (N_1176,N_847,N_926);
and U1177 (N_1177,N_611,N_799);
nor U1178 (N_1178,N_517,N_524);
and U1179 (N_1179,N_717,N_546);
nand U1180 (N_1180,N_516,N_791);
nand U1181 (N_1181,N_930,N_725);
or U1182 (N_1182,N_991,N_503);
xnor U1183 (N_1183,N_654,N_536);
nor U1184 (N_1184,N_662,N_758);
nand U1185 (N_1185,N_650,N_620);
xnor U1186 (N_1186,N_727,N_580);
and U1187 (N_1187,N_638,N_640);
nor U1188 (N_1188,N_508,N_796);
nand U1189 (N_1189,N_888,N_575);
xor U1190 (N_1190,N_957,N_893);
xnor U1191 (N_1191,N_660,N_752);
and U1192 (N_1192,N_820,N_770);
xor U1193 (N_1193,N_884,N_700);
xor U1194 (N_1194,N_794,N_997);
nand U1195 (N_1195,N_766,N_723);
or U1196 (N_1196,N_827,N_971);
nand U1197 (N_1197,N_630,N_726);
nand U1198 (N_1198,N_588,N_907);
nand U1199 (N_1199,N_887,N_668);
xnor U1200 (N_1200,N_590,N_780);
and U1201 (N_1201,N_561,N_594);
or U1202 (N_1202,N_768,N_513);
nand U1203 (N_1203,N_935,N_882);
nor U1204 (N_1204,N_742,N_648);
and U1205 (N_1205,N_806,N_862);
nor U1206 (N_1206,N_917,N_898);
nand U1207 (N_1207,N_819,N_639);
xnor U1208 (N_1208,N_983,N_940);
or U1209 (N_1209,N_877,N_657);
nor U1210 (N_1210,N_731,N_999);
nand U1211 (N_1211,N_568,N_924);
or U1212 (N_1212,N_736,N_978);
or U1213 (N_1213,N_593,N_618);
nand U1214 (N_1214,N_774,N_813);
nor U1215 (N_1215,N_857,N_778);
nor U1216 (N_1216,N_929,N_556);
nand U1217 (N_1217,N_871,N_908);
xor U1218 (N_1218,N_769,N_553);
or U1219 (N_1219,N_815,N_535);
and U1220 (N_1220,N_571,N_936);
xnor U1221 (N_1221,N_946,N_858);
nor U1222 (N_1222,N_663,N_841);
nor U1223 (N_1223,N_624,N_795);
or U1224 (N_1224,N_948,N_865);
or U1225 (N_1225,N_941,N_647);
and U1226 (N_1226,N_509,N_549);
and U1227 (N_1227,N_677,N_525);
xnor U1228 (N_1228,N_837,N_863);
or U1229 (N_1229,N_981,N_658);
nand U1230 (N_1230,N_840,N_626);
and U1231 (N_1231,N_864,N_993);
or U1232 (N_1232,N_822,N_890);
xor U1233 (N_1233,N_632,N_844);
or U1234 (N_1234,N_977,N_505);
nand U1235 (N_1235,N_952,N_760);
xnor U1236 (N_1236,N_562,N_880);
nand U1237 (N_1237,N_809,N_613);
nor U1238 (N_1238,N_596,N_980);
nor U1239 (N_1239,N_573,N_757);
nand U1240 (N_1240,N_904,N_518);
nor U1241 (N_1241,N_612,N_987);
nor U1242 (N_1242,N_812,N_852);
nand U1243 (N_1243,N_951,N_512);
and U1244 (N_1244,N_969,N_666);
or U1245 (N_1245,N_959,N_698);
and U1246 (N_1246,N_755,N_918);
or U1247 (N_1247,N_616,N_643);
and U1248 (N_1248,N_514,N_652);
and U1249 (N_1249,N_687,N_876);
and U1250 (N_1250,N_859,N_530);
nand U1251 (N_1251,N_682,N_842);
xor U1252 (N_1252,N_934,N_835);
or U1253 (N_1253,N_908,N_938);
or U1254 (N_1254,N_729,N_856);
or U1255 (N_1255,N_756,N_898);
and U1256 (N_1256,N_819,N_774);
or U1257 (N_1257,N_533,N_870);
nand U1258 (N_1258,N_860,N_849);
nor U1259 (N_1259,N_834,N_747);
or U1260 (N_1260,N_858,N_805);
nor U1261 (N_1261,N_826,N_898);
xor U1262 (N_1262,N_531,N_881);
and U1263 (N_1263,N_953,N_788);
xnor U1264 (N_1264,N_703,N_543);
nor U1265 (N_1265,N_787,N_761);
xor U1266 (N_1266,N_976,N_787);
nor U1267 (N_1267,N_782,N_522);
nand U1268 (N_1268,N_739,N_730);
or U1269 (N_1269,N_526,N_561);
nor U1270 (N_1270,N_545,N_620);
nor U1271 (N_1271,N_757,N_739);
nor U1272 (N_1272,N_688,N_702);
nand U1273 (N_1273,N_953,N_543);
nor U1274 (N_1274,N_730,N_748);
or U1275 (N_1275,N_937,N_893);
nand U1276 (N_1276,N_651,N_996);
and U1277 (N_1277,N_773,N_708);
and U1278 (N_1278,N_645,N_545);
and U1279 (N_1279,N_888,N_698);
or U1280 (N_1280,N_800,N_566);
and U1281 (N_1281,N_507,N_998);
xor U1282 (N_1282,N_605,N_612);
or U1283 (N_1283,N_868,N_824);
nand U1284 (N_1284,N_552,N_695);
or U1285 (N_1285,N_967,N_606);
nor U1286 (N_1286,N_875,N_871);
or U1287 (N_1287,N_840,N_791);
nor U1288 (N_1288,N_878,N_713);
xnor U1289 (N_1289,N_553,N_826);
nor U1290 (N_1290,N_536,N_551);
xnor U1291 (N_1291,N_614,N_735);
nor U1292 (N_1292,N_564,N_899);
xor U1293 (N_1293,N_895,N_792);
or U1294 (N_1294,N_561,N_782);
nand U1295 (N_1295,N_685,N_825);
xor U1296 (N_1296,N_787,N_647);
xor U1297 (N_1297,N_898,N_721);
nand U1298 (N_1298,N_669,N_901);
xnor U1299 (N_1299,N_995,N_589);
nand U1300 (N_1300,N_527,N_920);
xnor U1301 (N_1301,N_994,N_915);
nand U1302 (N_1302,N_949,N_563);
nor U1303 (N_1303,N_863,N_919);
or U1304 (N_1304,N_911,N_994);
and U1305 (N_1305,N_675,N_536);
nor U1306 (N_1306,N_859,N_703);
nor U1307 (N_1307,N_760,N_706);
or U1308 (N_1308,N_932,N_628);
or U1309 (N_1309,N_974,N_646);
and U1310 (N_1310,N_721,N_953);
nand U1311 (N_1311,N_889,N_775);
nand U1312 (N_1312,N_792,N_666);
nand U1313 (N_1313,N_800,N_838);
xor U1314 (N_1314,N_932,N_907);
or U1315 (N_1315,N_755,N_630);
and U1316 (N_1316,N_791,N_584);
xnor U1317 (N_1317,N_663,N_657);
or U1318 (N_1318,N_665,N_786);
xnor U1319 (N_1319,N_751,N_881);
nand U1320 (N_1320,N_556,N_933);
nor U1321 (N_1321,N_625,N_633);
nor U1322 (N_1322,N_624,N_746);
xor U1323 (N_1323,N_532,N_951);
and U1324 (N_1324,N_885,N_985);
xor U1325 (N_1325,N_789,N_772);
nor U1326 (N_1326,N_964,N_811);
nor U1327 (N_1327,N_983,N_685);
and U1328 (N_1328,N_922,N_885);
and U1329 (N_1329,N_849,N_915);
xor U1330 (N_1330,N_832,N_645);
or U1331 (N_1331,N_870,N_654);
xor U1332 (N_1332,N_812,N_860);
xor U1333 (N_1333,N_557,N_784);
nand U1334 (N_1334,N_573,N_511);
nor U1335 (N_1335,N_652,N_855);
or U1336 (N_1336,N_849,N_953);
nor U1337 (N_1337,N_727,N_745);
nand U1338 (N_1338,N_758,N_706);
nor U1339 (N_1339,N_916,N_944);
and U1340 (N_1340,N_602,N_759);
and U1341 (N_1341,N_864,N_868);
nand U1342 (N_1342,N_647,N_927);
xor U1343 (N_1343,N_656,N_968);
or U1344 (N_1344,N_586,N_643);
or U1345 (N_1345,N_690,N_529);
and U1346 (N_1346,N_528,N_771);
and U1347 (N_1347,N_902,N_550);
xor U1348 (N_1348,N_721,N_658);
or U1349 (N_1349,N_898,N_889);
or U1350 (N_1350,N_847,N_916);
nor U1351 (N_1351,N_820,N_742);
nor U1352 (N_1352,N_541,N_626);
xor U1353 (N_1353,N_585,N_504);
or U1354 (N_1354,N_701,N_912);
nand U1355 (N_1355,N_759,N_886);
xor U1356 (N_1356,N_549,N_796);
nand U1357 (N_1357,N_681,N_593);
or U1358 (N_1358,N_706,N_583);
xor U1359 (N_1359,N_786,N_561);
and U1360 (N_1360,N_894,N_916);
nor U1361 (N_1361,N_646,N_900);
xnor U1362 (N_1362,N_585,N_796);
nand U1363 (N_1363,N_887,N_963);
and U1364 (N_1364,N_886,N_721);
or U1365 (N_1365,N_594,N_749);
nor U1366 (N_1366,N_815,N_605);
or U1367 (N_1367,N_645,N_772);
nor U1368 (N_1368,N_793,N_663);
and U1369 (N_1369,N_848,N_537);
or U1370 (N_1370,N_691,N_993);
or U1371 (N_1371,N_776,N_629);
xnor U1372 (N_1372,N_777,N_869);
nor U1373 (N_1373,N_870,N_914);
nand U1374 (N_1374,N_694,N_734);
xor U1375 (N_1375,N_525,N_714);
xnor U1376 (N_1376,N_794,N_871);
nor U1377 (N_1377,N_613,N_723);
or U1378 (N_1378,N_736,N_806);
xnor U1379 (N_1379,N_646,N_981);
nor U1380 (N_1380,N_714,N_827);
and U1381 (N_1381,N_795,N_519);
nand U1382 (N_1382,N_574,N_579);
xnor U1383 (N_1383,N_792,N_624);
xor U1384 (N_1384,N_554,N_848);
or U1385 (N_1385,N_764,N_921);
nand U1386 (N_1386,N_997,N_880);
xor U1387 (N_1387,N_934,N_546);
nand U1388 (N_1388,N_512,N_854);
and U1389 (N_1389,N_964,N_791);
nand U1390 (N_1390,N_600,N_722);
or U1391 (N_1391,N_925,N_637);
xor U1392 (N_1392,N_651,N_926);
and U1393 (N_1393,N_770,N_649);
nand U1394 (N_1394,N_663,N_678);
xor U1395 (N_1395,N_699,N_659);
nand U1396 (N_1396,N_540,N_850);
nand U1397 (N_1397,N_777,N_982);
nor U1398 (N_1398,N_587,N_519);
and U1399 (N_1399,N_840,N_624);
nor U1400 (N_1400,N_957,N_502);
xor U1401 (N_1401,N_769,N_790);
nor U1402 (N_1402,N_517,N_900);
xor U1403 (N_1403,N_912,N_841);
or U1404 (N_1404,N_766,N_596);
xor U1405 (N_1405,N_983,N_553);
and U1406 (N_1406,N_713,N_714);
or U1407 (N_1407,N_749,N_581);
nand U1408 (N_1408,N_635,N_889);
nor U1409 (N_1409,N_769,N_908);
nand U1410 (N_1410,N_646,N_616);
xor U1411 (N_1411,N_909,N_503);
xnor U1412 (N_1412,N_660,N_886);
or U1413 (N_1413,N_575,N_610);
and U1414 (N_1414,N_885,N_690);
nand U1415 (N_1415,N_530,N_786);
xor U1416 (N_1416,N_838,N_763);
nor U1417 (N_1417,N_881,N_737);
xnor U1418 (N_1418,N_556,N_920);
xnor U1419 (N_1419,N_856,N_906);
xnor U1420 (N_1420,N_577,N_649);
nand U1421 (N_1421,N_956,N_652);
and U1422 (N_1422,N_775,N_860);
xor U1423 (N_1423,N_887,N_713);
nand U1424 (N_1424,N_995,N_559);
xnor U1425 (N_1425,N_593,N_856);
and U1426 (N_1426,N_628,N_643);
nand U1427 (N_1427,N_533,N_539);
nor U1428 (N_1428,N_940,N_838);
xor U1429 (N_1429,N_674,N_667);
nand U1430 (N_1430,N_522,N_891);
or U1431 (N_1431,N_796,N_708);
nor U1432 (N_1432,N_738,N_665);
and U1433 (N_1433,N_523,N_647);
xor U1434 (N_1434,N_751,N_796);
or U1435 (N_1435,N_845,N_682);
and U1436 (N_1436,N_519,N_787);
or U1437 (N_1437,N_745,N_771);
or U1438 (N_1438,N_787,N_759);
nand U1439 (N_1439,N_590,N_824);
xor U1440 (N_1440,N_597,N_576);
and U1441 (N_1441,N_842,N_836);
and U1442 (N_1442,N_642,N_983);
nand U1443 (N_1443,N_500,N_823);
or U1444 (N_1444,N_699,N_869);
and U1445 (N_1445,N_941,N_908);
or U1446 (N_1446,N_506,N_571);
and U1447 (N_1447,N_800,N_589);
or U1448 (N_1448,N_565,N_659);
or U1449 (N_1449,N_904,N_656);
nand U1450 (N_1450,N_952,N_661);
nor U1451 (N_1451,N_567,N_582);
nand U1452 (N_1452,N_721,N_570);
nand U1453 (N_1453,N_927,N_834);
nand U1454 (N_1454,N_540,N_754);
nand U1455 (N_1455,N_850,N_666);
or U1456 (N_1456,N_872,N_523);
nand U1457 (N_1457,N_910,N_580);
nand U1458 (N_1458,N_865,N_708);
xnor U1459 (N_1459,N_949,N_531);
or U1460 (N_1460,N_522,N_556);
nor U1461 (N_1461,N_673,N_813);
nand U1462 (N_1462,N_971,N_952);
xnor U1463 (N_1463,N_512,N_513);
nor U1464 (N_1464,N_973,N_554);
nand U1465 (N_1465,N_599,N_752);
xnor U1466 (N_1466,N_638,N_632);
nor U1467 (N_1467,N_850,N_671);
xnor U1468 (N_1468,N_632,N_994);
or U1469 (N_1469,N_725,N_742);
and U1470 (N_1470,N_797,N_619);
nor U1471 (N_1471,N_924,N_809);
nand U1472 (N_1472,N_561,N_875);
nor U1473 (N_1473,N_895,N_530);
or U1474 (N_1474,N_873,N_577);
nor U1475 (N_1475,N_575,N_834);
xnor U1476 (N_1476,N_960,N_722);
or U1477 (N_1477,N_614,N_550);
xnor U1478 (N_1478,N_983,N_732);
nand U1479 (N_1479,N_790,N_825);
nand U1480 (N_1480,N_675,N_532);
nand U1481 (N_1481,N_684,N_581);
xnor U1482 (N_1482,N_990,N_533);
nor U1483 (N_1483,N_927,N_866);
xor U1484 (N_1484,N_849,N_975);
or U1485 (N_1485,N_756,N_862);
xor U1486 (N_1486,N_649,N_935);
nor U1487 (N_1487,N_663,N_910);
nand U1488 (N_1488,N_951,N_670);
or U1489 (N_1489,N_900,N_993);
or U1490 (N_1490,N_716,N_816);
nor U1491 (N_1491,N_534,N_519);
or U1492 (N_1492,N_875,N_643);
and U1493 (N_1493,N_704,N_942);
and U1494 (N_1494,N_597,N_999);
or U1495 (N_1495,N_513,N_805);
or U1496 (N_1496,N_755,N_905);
or U1497 (N_1497,N_663,N_609);
or U1498 (N_1498,N_833,N_988);
or U1499 (N_1499,N_966,N_779);
or U1500 (N_1500,N_1133,N_1478);
xnor U1501 (N_1501,N_1203,N_1319);
nand U1502 (N_1502,N_1099,N_1148);
nand U1503 (N_1503,N_1057,N_1171);
xnor U1504 (N_1504,N_1321,N_1042);
or U1505 (N_1505,N_1198,N_1205);
nor U1506 (N_1506,N_1410,N_1398);
and U1507 (N_1507,N_1139,N_1115);
nor U1508 (N_1508,N_1180,N_1156);
nor U1509 (N_1509,N_1263,N_1345);
xor U1510 (N_1510,N_1275,N_1300);
xnor U1511 (N_1511,N_1132,N_1040);
and U1512 (N_1512,N_1496,N_1187);
or U1513 (N_1513,N_1058,N_1073);
xnor U1514 (N_1514,N_1365,N_1480);
or U1515 (N_1515,N_1333,N_1189);
nor U1516 (N_1516,N_1165,N_1181);
nand U1517 (N_1517,N_1110,N_1092);
xor U1518 (N_1518,N_1352,N_1422);
or U1519 (N_1519,N_1491,N_1477);
and U1520 (N_1520,N_1046,N_1379);
xnor U1521 (N_1521,N_1395,N_1464);
and U1522 (N_1522,N_1453,N_1002);
and U1523 (N_1523,N_1388,N_1304);
xor U1524 (N_1524,N_1179,N_1278);
or U1525 (N_1525,N_1037,N_1079);
nor U1526 (N_1526,N_1201,N_1017);
xor U1527 (N_1527,N_1234,N_1141);
and U1528 (N_1528,N_1217,N_1430);
nor U1529 (N_1529,N_1396,N_1348);
xnor U1530 (N_1530,N_1355,N_1206);
or U1531 (N_1531,N_1039,N_1276);
xor U1532 (N_1532,N_1241,N_1380);
nor U1533 (N_1533,N_1183,N_1219);
or U1534 (N_1534,N_1003,N_1193);
nand U1535 (N_1535,N_1247,N_1339);
and U1536 (N_1536,N_1147,N_1415);
xnor U1537 (N_1537,N_1036,N_1296);
xor U1538 (N_1538,N_1486,N_1471);
nor U1539 (N_1539,N_1392,N_1439);
nand U1540 (N_1540,N_1474,N_1288);
and U1541 (N_1541,N_1063,N_1460);
nor U1542 (N_1542,N_1364,N_1083);
and U1543 (N_1543,N_1331,N_1213);
or U1544 (N_1544,N_1232,N_1377);
or U1545 (N_1545,N_1067,N_1235);
xnor U1546 (N_1546,N_1320,N_1294);
xor U1547 (N_1547,N_1318,N_1255);
nor U1548 (N_1548,N_1100,N_1218);
nor U1549 (N_1549,N_1479,N_1074);
or U1550 (N_1550,N_1428,N_1459);
xor U1551 (N_1551,N_1421,N_1382);
xor U1552 (N_1552,N_1363,N_1178);
nand U1553 (N_1553,N_1168,N_1055);
nand U1554 (N_1554,N_1495,N_1081);
nor U1555 (N_1555,N_1142,N_1243);
and U1556 (N_1556,N_1401,N_1314);
nor U1557 (N_1557,N_1476,N_1282);
nand U1558 (N_1558,N_1104,N_1118);
nand U1559 (N_1559,N_1208,N_1077);
nor U1560 (N_1560,N_1146,N_1116);
xnor U1561 (N_1561,N_1311,N_1256);
or U1562 (N_1562,N_1076,N_1498);
nand U1563 (N_1563,N_1440,N_1089);
or U1564 (N_1564,N_1335,N_1354);
and U1565 (N_1565,N_1358,N_1436);
nor U1566 (N_1566,N_1411,N_1091);
xnor U1567 (N_1567,N_1417,N_1405);
xnor U1568 (N_1568,N_1281,N_1093);
nand U1569 (N_1569,N_1001,N_1134);
xor U1570 (N_1570,N_1402,N_1023);
xnor U1571 (N_1571,N_1188,N_1145);
nor U1572 (N_1572,N_1420,N_1162);
or U1573 (N_1573,N_1293,N_1360);
xor U1574 (N_1574,N_1452,N_1324);
nand U1575 (N_1575,N_1197,N_1350);
nand U1576 (N_1576,N_1071,N_1466);
nand U1577 (N_1577,N_1385,N_1028);
xnor U1578 (N_1578,N_1468,N_1131);
nand U1579 (N_1579,N_1177,N_1284);
or U1580 (N_1580,N_1010,N_1397);
xor U1581 (N_1581,N_1418,N_1222);
nand U1582 (N_1582,N_1246,N_1386);
xnor U1583 (N_1583,N_1493,N_1435);
and U1584 (N_1584,N_1427,N_1049);
nor U1585 (N_1585,N_1112,N_1034);
nor U1586 (N_1586,N_1238,N_1357);
or U1587 (N_1587,N_1462,N_1429);
nor U1588 (N_1588,N_1444,N_1170);
nand U1589 (N_1589,N_1408,N_1259);
nor U1590 (N_1590,N_1064,N_1475);
xnor U1591 (N_1591,N_1458,N_1200);
and U1592 (N_1592,N_1406,N_1054);
or U1593 (N_1593,N_1223,N_1492);
nand U1594 (N_1594,N_1253,N_1119);
nand U1595 (N_1595,N_1024,N_1280);
or U1596 (N_1596,N_1102,N_1456);
or U1597 (N_1597,N_1048,N_1271);
nor U1598 (N_1598,N_1204,N_1370);
or U1599 (N_1599,N_1033,N_1220);
nand U1600 (N_1600,N_1457,N_1032);
nor U1601 (N_1601,N_1287,N_1065);
nand U1602 (N_1602,N_1260,N_1016);
or U1603 (N_1603,N_1265,N_1378);
xor U1604 (N_1604,N_1114,N_1268);
nor U1605 (N_1605,N_1409,N_1163);
and U1606 (N_1606,N_1394,N_1442);
and U1607 (N_1607,N_1096,N_1266);
nor U1608 (N_1608,N_1419,N_1214);
nand U1609 (N_1609,N_1356,N_1346);
nand U1610 (N_1610,N_1221,N_1233);
or U1611 (N_1611,N_1020,N_1309);
or U1612 (N_1612,N_1012,N_1006);
xnor U1613 (N_1613,N_1349,N_1375);
nand U1614 (N_1614,N_1251,N_1371);
nor U1615 (N_1615,N_1239,N_1191);
or U1616 (N_1616,N_1069,N_1080);
or U1617 (N_1617,N_1313,N_1196);
and U1618 (N_1618,N_1154,N_1323);
nand U1619 (N_1619,N_1490,N_1021);
nand U1620 (N_1620,N_1164,N_1261);
nor U1621 (N_1621,N_1025,N_1446);
xnor U1622 (N_1622,N_1128,N_1143);
xor U1623 (N_1623,N_1455,N_1270);
nand U1624 (N_1624,N_1240,N_1066);
xor U1625 (N_1625,N_1050,N_1085);
nand U1626 (N_1626,N_1144,N_1136);
nand U1627 (N_1627,N_1126,N_1431);
nand U1628 (N_1628,N_1315,N_1101);
nor U1629 (N_1629,N_1194,N_1307);
and U1630 (N_1630,N_1301,N_1332);
or U1631 (N_1631,N_1328,N_1072);
xnor U1632 (N_1632,N_1387,N_1122);
xor U1633 (N_1633,N_1159,N_1285);
and U1634 (N_1634,N_1123,N_1424);
nor U1635 (N_1635,N_1152,N_1433);
nor U1636 (N_1636,N_1111,N_1225);
nor U1637 (N_1637,N_1173,N_1400);
nor U1638 (N_1638,N_1264,N_1212);
xor U1639 (N_1639,N_1403,N_1082);
nand U1640 (N_1640,N_1224,N_1098);
or U1641 (N_1641,N_1423,N_1120);
xor U1642 (N_1642,N_1090,N_1105);
or U1643 (N_1643,N_1472,N_1237);
nor U1644 (N_1644,N_1150,N_1291);
xnor U1645 (N_1645,N_1202,N_1041);
and U1646 (N_1646,N_1393,N_1106);
xor U1647 (N_1647,N_1250,N_1044);
nand U1648 (N_1648,N_1267,N_1481);
or U1649 (N_1649,N_1153,N_1426);
xor U1650 (N_1650,N_1487,N_1340);
xnor U1651 (N_1651,N_1051,N_1008);
xor U1652 (N_1652,N_1438,N_1192);
and U1653 (N_1653,N_1390,N_1434);
or U1654 (N_1654,N_1155,N_1283);
nand U1655 (N_1655,N_1359,N_1022);
nor U1656 (N_1656,N_1445,N_1432);
or U1657 (N_1657,N_1094,N_1470);
xnor U1658 (N_1658,N_1229,N_1211);
and U1659 (N_1659,N_1329,N_1190);
nand U1660 (N_1660,N_1035,N_1108);
nor U1661 (N_1661,N_1000,N_1292);
nand U1662 (N_1662,N_1425,N_1277);
nand U1663 (N_1663,N_1075,N_1068);
xnor U1664 (N_1664,N_1011,N_1019);
or U1665 (N_1665,N_1448,N_1262);
nand U1666 (N_1666,N_1174,N_1404);
nand U1667 (N_1667,N_1447,N_1231);
and U1668 (N_1668,N_1373,N_1061);
nand U1669 (N_1669,N_1004,N_1416);
nand U1670 (N_1670,N_1306,N_1374);
and U1671 (N_1671,N_1412,N_1182);
or U1672 (N_1672,N_1485,N_1298);
and U1673 (N_1673,N_1351,N_1103);
xor U1674 (N_1674,N_1312,N_1451);
or U1675 (N_1675,N_1030,N_1184);
or U1676 (N_1676,N_1084,N_1245);
or U1677 (N_1677,N_1062,N_1299);
nand U1678 (N_1678,N_1242,N_1463);
or U1679 (N_1679,N_1052,N_1342);
nor U1680 (N_1680,N_1166,N_1443);
nor U1681 (N_1681,N_1169,N_1149);
or U1682 (N_1682,N_1322,N_1279);
nand U1683 (N_1683,N_1060,N_1316);
nand U1684 (N_1684,N_1140,N_1088);
nand U1685 (N_1685,N_1336,N_1244);
nand U1686 (N_1686,N_1249,N_1369);
nand U1687 (N_1687,N_1469,N_1199);
nand U1688 (N_1688,N_1384,N_1130);
nor U1689 (N_1689,N_1172,N_1461);
xnor U1690 (N_1690,N_1414,N_1043);
and U1691 (N_1691,N_1308,N_1347);
or U1692 (N_1692,N_1095,N_1195);
and U1693 (N_1693,N_1053,N_1047);
nor U1694 (N_1694,N_1027,N_1399);
nand U1695 (N_1695,N_1014,N_1361);
xor U1696 (N_1696,N_1018,N_1097);
xnor U1697 (N_1697,N_1209,N_1454);
and U1698 (N_1698,N_1302,N_1135);
nor U1699 (N_1699,N_1230,N_1167);
nand U1700 (N_1700,N_1059,N_1031);
or U1701 (N_1701,N_1029,N_1273);
xnor U1702 (N_1702,N_1482,N_1437);
and U1703 (N_1703,N_1107,N_1129);
or U1704 (N_1704,N_1009,N_1473);
or U1705 (N_1705,N_1407,N_1045);
or U1706 (N_1706,N_1254,N_1161);
nor U1707 (N_1707,N_1272,N_1158);
or U1708 (N_1708,N_1185,N_1327);
nor U1709 (N_1709,N_1227,N_1497);
nor U1710 (N_1710,N_1207,N_1344);
or U1711 (N_1711,N_1216,N_1137);
nor U1712 (N_1712,N_1372,N_1391);
or U1713 (N_1713,N_1269,N_1257);
nor U1714 (N_1714,N_1078,N_1038);
xor U1715 (N_1715,N_1087,N_1274);
or U1716 (N_1716,N_1305,N_1127);
or U1717 (N_1717,N_1286,N_1026);
nand U1718 (N_1718,N_1210,N_1337);
xor U1719 (N_1719,N_1343,N_1499);
xor U1720 (N_1720,N_1383,N_1289);
xor U1721 (N_1721,N_1215,N_1488);
nand U1722 (N_1722,N_1109,N_1236);
and U1723 (N_1723,N_1005,N_1389);
and U1724 (N_1724,N_1341,N_1013);
and U1725 (N_1725,N_1290,N_1228);
or U1726 (N_1726,N_1367,N_1441);
xnor U1727 (N_1727,N_1151,N_1157);
and U1728 (N_1728,N_1381,N_1317);
nor U1729 (N_1729,N_1226,N_1467);
and U1730 (N_1730,N_1124,N_1295);
or U1731 (N_1731,N_1334,N_1483);
or U1732 (N_1732,N_1449,N_1484);
and U1733 (N_1733,N_1489,N_1303);
nor U1734 (N_1734,N_1366,N_1330);
or U1735 (N_1735,N_1258,N_1368);
xor U1736 (N_1736,N_1176,N_1186);
or U1737 (N_1737,N_1450,N_1015);
nor U1738 (N_1738,N_1070,N_1325);
xnor U1739 (N_1739,N_1353,N_1125);
xor U1740 (N_1740,N_1117,N_1007);
and U1741 (N_1741,N_1248,N_1138);
and U1742 (N_1742,N_1465,N_1056);
xor U1743 (N_1743,N_1494,N_1086);
xnor U1744 (N_1744,N_1252,N_1160);
nor U1745 (N_1745,N_1121,N_1297);
or U1746 (N_1746,N_1310,N_1413);
and U1747 (N_1747,N_1326,N_1338);
or U1748 (N_1748,N_1175,N_1362);
xor U1749 (N_1749,N_1376,N_1113);
nand U1750 (N_1750,N_1254,N_1306);
or U1751 (N_1751,N_1089,N_1464);
nand U1752 (N_1752,N_1067,N_1256);
or U1753 (N_1753,N_1191,N_1435);
nand U1754 (N_1754,N_1370,N_1220);
or U1755 (N_1755,N_1157,N_1386);
or U1756 (N_1756,N_1288,N_1114);
nand U1757 (N_1757,N_1143,N_1287);
and U1758 (N_1758,N_1439,N_1199);
or U1759 (N_1759,N_1119,N_1438);
and U1760 (N_1760,N_1229,N_1366);
nand U1761 (N_1761,N_1121,N_1132);
and U1762 (N_1762,N_1224,N_1077);
or U1763 (N_1763,N_1403,N_1153);
xor U1764 (N_1764,N_1147,N_1229);
or U1765 (N_1765,N_1331,N_1361);
or U1766 (N_1766,N_1041,N_1465);
xor U1767 (N_1767,N_1198,N_1020);
nand U1768 (N_1768,N_1236,N_1157);
and U1769 (N_1769,N_1403,N_1286);
xor U1770 (N_1770,N_1379,N_1270);
and U1771 (N_1771,N_1119,N_1315);
xor U1772 (N_1772,N_1231,N_1115);
or U1773 (N_1773,N_1438,N_1388);
nor U1774 (N_1774,N_1166,N_1356);
nor U1775 (N_1775,N_1402,N_1217);
xor U1776 (N_1776,N_1034,N_1130);
xor U1777 (N_1777,N_1064,N_1430);
or U1778 (N_1778,N_1033,N_1139);
xor U1779 (N_1779,N_1331,N_1443);
nor U1780 (N_1780,N_1486,N_1109);
nand U1781 (N_1781,N_1104,N_1396);
or U1782 (N_1782,N_1411,N_1199);
and U1783 (N_1783,N_1452,N_1001);
or U1784 (N_1784,N_1195,N_1402);
and U1785 (N_1785,N_1083,N_1202);
nor U1786 (N_1786,N_1484,N_1293);
nor U1787 (N_1787,N_1294,N_1063);
nor U1788 (N_1788,N_1129,N_1288);
nor U1789 (N_1789,N_1446,N_1180);
nand U1790 (N_1790,N_1092,N_1254);
nand U1791 (N_1791,N_1131,N_1171);
and U1792 (N_1792,N_1242,N_1190);
nand U1793 (N_1793,N_1285,N_1495);
and U1794 (N_1794,N_1227,N_1339);
nor U1795 (N_1795,N_1408,N_1495);
nor U1796 (N_1796,N_1300,N_1179);
and U1797 (N_1797,N_1406,N_1229);
xnor U1798 (N_1798,N_1112,N_1170);
nor U1799 (N_1799,N_1166,N_1251);
or U1800 (N_1800,N_1165,N_1193);
and U1801 (N_1801,N_1357,N_1061);
and U1802 (N_1802,N_1493,N_1169);
nor U1803 (N_1803,N_1367,N_1115);
or U1804 (N_1804,N_1491,N_1445);
and U1805 (N_1805,N_1391,N_1307);
nand U1806 (N_1806,N_1460,N_1430);
xnor U1807 (N_1807,N_1010,N_1177);
nand U1808 (N_1808,N_1049,N_1290);
nand U1809 (N_1809,N_1203,N_1153);
xnor U1810 (N_1810,N_1082,N_1446);
xor U1811 (N_1811,N_1191,N_1123);
nand U1812 (N_1812,N_1013,N_1388);
nor U1813 (N_1813,N_1122,N_1172);
or U1814 (N_1814,N_1474,N_1042);
nand U1815 (N_1815,N_1149,N_1127);
or U1816 (N_1816,N_1033,N_1440);
nor U1817 (N_1817,N_1433,N_1079);
and U1818 (N_1818,N_1083,N_1395);
or U1819 (N_1819,N_1004,N_1153);
xnor U1820 (N_1820,N_1488,N_1485);
nand U1821 (N_1821,N_1228,N_1126);
nor U1822 (N_1822,N_1353,N_1455);
nor U1823 (N_1823,N_1374,N_1016);
xnor U1824 (N_1824,N_1435,N_1212);
nor U1825 (N_1825,N_1303,N_1253);
nand U1826 (N_1826,N_1408,N_1237);
or U1827 (N_1827,N_1300,N_1040);
nor U1828 (N_1828,N_1453,N_1455);
nor U1829 (N_1829,N_1259,N_1118);
xor U1830 (N_1830,N_1090,N_1295);
or U1831 (N_1831,N_1008,N_1072);
and U1832 (N_1832,N_1253,N_1008);
nand U1833 (N_1833,N_1198,N_1316);
nor U1834 (N_1834,N_1105,N_1247);
nor U1835 (N_1835,N_1179,N_1461);
xnor U1836 (N_1836,N_1037,N_1431);
nor U1837 (N_1837,N_1032,N_1030);
and U1838 (N_1838,N_1074,N_1483);
or U1839 (N_1839,N_1357,N_1391);
and U1840 (N_1840,N_1090,N_1129);
nor U1841 (N_1841,N_1247,N_1088);
and U1842 (N_1842,N_1490,N_1184);
nor U1843 (N_1843,N_1395,N_1038);
nand U1844 (N_1844,N_1473,N_1359);
or U1845 (N_1845,N_1361,N_1351);
or U1846 (N_1846,N_1281,N_1318);
nor U1847 (N_1847,N_1215,N_1019);
and U1848 (N_1848,N_1336,N_1203);
and U1849 (N_1849,N_1424,N_1195);
xor U1850 (N_1850,N_1422,N_1310);
and U1851 (N_1851,N_1144,N_1069);
xor U1852 (N_1852,N_1007,N_1274);
xnor U1853 (N_1853,N_1150,N_1492);
or U1854 (N_1854,N_1458,N_1253);
xor U1855 (N_1855,N_1225,N_1254);
and U1856 (N_1856,N_1314,N_1407);
or U1857 (N_1857,N_1333,N_1335);
nand U1858 (N_1858,N_1159,N_1444);
nor U1859 (N_1859,N_1006,N_1323);
or U1860 (N_1860,N_1373,N_1349);
nand U1861 (N_1861,N_1498,N_1301);
nand U1862 (N_1862,N_1315,N_1335);
or U1863 (N_1863,N_1377,N_1086);
or U1864 (N_1864,N_1024,N_1358);
xnor U1865 (N_1865,N_1056,N_1317);
xnor U1866 (N_1866,N_1489,N_1366);
nor U1867 (N_1867,N_1078,N_1020);
xnor U1868 (N_1868,N_1217,N_1453);
nand U1869 (N_1869,N_1403,N_1119);
or U1870 (N_1870,N_1304,N_1147);
or U1871 (N_1871,N_1385,N_1263);
or U1872 (N_1872,N_1132,N_1410);
nor U1873 (N_1873,N_1411,N_1444);
or U1874 (N_1874,N_1159,N_1152);
or U1875 (N_1875,N_1255,N_1249);
or U1876 (N_1876,N_1258,N_1447);
xor U1877 (N_1877,N_1067,N_1117);
nand U1878 (N_1878,N_1249,N_1195);
and U1879 (N_1879,N_1391,N_1395);
and U1880 (N_1880,N_1298,N_1308);
xnor U1881 (N_1881,N_1086,N_1364);
and U1882 (N_1882,N_1082,N_1346);
and U1883 (N_1883,N_1496,N_1034);
xnor U1884 (N_1884,N_1133,N_1148);
nand U1885 (N_1885,N_1384,N_1211);
and U1886 (N_1886,N_1003,N_1075);
nor U1887 (N_1887,N_1248,N_1457);
or U1888 (N_1888,N_1193,N_1305);
nand U1889 (N_1889,N_1191,N_1177);
xnor U1890 (N_1890,N_1091,N_1448);
and U1891 (N_1891,N_1424,N_1414);
nand U1892 (N_1892,N_1292,N_1094);
and U1893 (N_1893,N_1184,N_1453);
or U1894 (N_1894,N_1185,N_1173);
or U1895 (N_1895,N_1067,N_1419);
and U1896 (N_1896,N_1178,N_1387);
and U1897 (N_1897,N_1300,N_1072);
xnor U1898 (N_1898,N_1058,N_1191);
nor U1899 (N_1899,N_1198,N_1481);
xor U1900 (N_1900,N_1030,N_1425);
and U1901 (N_1901,N_1144,N_1046);
and U1902 (N_1902,N_1041,N_1261);
xor U1903 (N_1903,N_1169,N_1010);
nand U1904 (N_1904,N_1000,N_1474);
or U1905 (N_1905,N_1077,N_1493);
nor U1906 (N_1906,N_1171,N_1184);
and U1907 (N_1907,N_1046,N_1047);
and U1908 (N_1908,N_1021,N_1127);
and U1909 (N_1909,N_1403,N_1215);
nor U1910 (N_1910,N_1274,N_1422);
or U1911 (N_1911,N_1104,N_1464);
nand U1912 (N_1912,N_1338,N_1329);
nand U1913 (N_1913,N_1454,N_1252);
nor U1914 (N_1914,N_1126,N_1382);
nand U1915 (N_1915,N_1210,N_1218);
and U1916 (N_1916,N_1272,N_1481);
nand U1917 (N_1917,N_1295,N_1079);
and U1918 (N_1918,N_1026,N_1167);
or U1919 (N_1919,N_1004,N_1202);
or U1920 (N_1920,N_1144,N_1493);
or U1921 (N_1921,N_1379,N_1306);
or U1922 (N_1922,N_1334,N_1319);
and U1923 (N_1923,N_1040,N_1017);
nor U1924 (N_1924,N_1315,N_1419);
nand U1925 (N_1925,N_1208,N_1212);
xor U1926 (N_1926,N_1027,N_1439);
nor U1927 (N_1927,N_1212,N_1462);
xor U1928 (N_1928,N_1009,N_1008);
nor U1929 (N_1929,N_1019,N_1023);
xnor U1930 (N_1930,N_1137,N_1241);
nand U1931 (N_1931,N_1185,N_1362);
or U1932 (N_1932,N_1447,N_1165);
or U1933 (N_1933,N_1118,N_1115);
and U1934 (N_1934,N_1055,N_1155);
or U1935 (N_1935,N_1328,N_1327);
or U1936 (N_1936,N_1309,N_1204);
or U1937 (N_1937,N_1134,N_1254);
and U1938 (N_1938,N_1354,N_1421);
xor U1939 (N_1939,N_1376,N_1158);
or U1940 (N_1940,N_1117,N_1357);
xor U1941 (N_1941,N_1052,N_1343);
xor U1942 (N_1942,N_1208,N_1085);
nor U1943 (N_1943,N_1002,N_1108);
or U1944 (N_1944,N_1118,N_1033);
or U1945 (N_1945,N_1067,N_1481);
or U1946 (N_1946,N_1120,N_1480);
nand U1947 (N_1947,N_1166,N_1057);
and U1948 (N_1948,N_1452,N_1237);
nand U1949 (N_1949,N_1223,N_1471);
or U1950 (N_1950,N_1247,N_1447);
or U1951 (N_1951,N_1497,N_1237);
nand U1952 (N_1952,N_1423,N_1465);
or U1953 (N_1953,N_1490,N_1003);
or U1954 (N_1954,N_1451,N_1053);
nand U1955 (N_1955,N_1061,N_1309);
xor U1956 (N_1956,N_1051,N_1428);
nand U1957 (N_1957,N_1425,N_1268);
or U1958 (N_1958,N_1282,N_1097);
or U1959 (N_1959,N_1247,N_1388);
nand U1960 (N_1960,N_1090,N_1209);
or U1961 (N_1961,N_1327,N_1347);
and U1962 (N_1962,N_1202,N_1369);
xnor U1963 (N_1963,N_1008,N_1415);
and U1964 (N_1964,N_1237,N_1366);
nor U1965 (N_1965,N_1463,N_1062);
xnor U1966 (N_1966,N_1328,N_1397);
nand U1967 (N_1967,N_1028,N_1429);
and U1968 (N_1968,N_1225,N_1449);
and U1969 (N_1969,N_1380,N_1443);
or U1970 (N_1970,N_1112,N_1269);
or U1971 (N_1971,N_1346,N_1165);
or U1972 (N_1972,N_1281,N_1487);
nor U1973 (N_1973,N_1283,N_1234);
nor U1974 (N_1974,N_1268,N_1415);
nor U1975 (N_1975,N_1091,N_1353);
xnor U1976 (N_1976,N_1043,N_1302);
and U1977 (N_1977,N_1487,N_1384);
or U1978 (N_1978,N_1182,N_1270);
and U1979 (N_1979,N_1390,N_1246);
nor U1980 (N_1980,N_1187,N_1302);
and U1981 (N_1981,N_1040,N_1230);
nor U1982 (N_1982,N_1194,N_1222);
and U1983 (N_1983,N_1253,N_1012);
or U1984 (N_1984,N_1142,N_1368);
xor U1985 (N_1985,N_1328,N_1312);
nand U1986 (N_1986,N_1164,N_1338);
nor U1987 (N_1987,N_1443,N_1248);
xor U1988 (N_1988,N_1240,N_1229);
xnor U1989 (N_1989,N_1436,N_1308);
or U1990 (N_1990,N_1096,N_1021);
xnor U1991 (N_1991,N_1366,N_1087);
and U1992 (N_1992,N_1309,N_1180);
or U1993 (N_1993,N_1015,N_1148);
xor U1994 (N_1994,N_1370,N_1086);
and U1995 (N_1995,N_1213,N_1358);
nor U1996 (N_1996,N_1466,N_1288);
and U1997 (N_1997,N_1227,N_1289);
nand U1998 (N_1998,N_1033,N_1423);
xor U1999 (N_1999,N_1185,N_1457);
xnor U2000 (N_2000,N_1829,N_1552);
xnor U2001 (N_2001,N_1831,N_1738);
xnor U2002 (N_2002,N_1613,N_1793);
or U2003 (N_2003,N_1665,N_1630);
or U2004 (N_2004,N_1536,N_1694);
or U2005 (N_2005,N_1861,N_1688);
nand U2006 (N_2006,N_1847,N_1987);
and U2007 (N_2007,N_1983,N_1509);
xor U2008 (N_2008,N_1959,N_1689);
nand U2009 (N_2009,N_1669,N_1948);
or U2010 (N_2010,N_1743,N_1928);
and U2011 (N_2011,N_1652,N_1686);
and U2012 (N_2012,N_1964,N_1540);
xor U2013 (N_2013,N_1730,N_1742);
nand U2014 (N_2014,N_1558,N_1548);
or U2015 (N_2015,N_1655,N_1937);
xor U2016 (N_2016,N_1780,N_1549);
nand U2017 (N_2017,N_1758,N_1776);
and U2018 (N_2018,N_1573,N_1579);
or U2019 (N_2019,N_1707,N_1998);
nand U2020 (N_2020,N_1832,N_1988);
nor U2021 (N_2021,N_1551,N_1556);
and U2022 (N_2022,N_1524,N_1834);
xor U2023 (N_2023,N_1800,N_1868);
and U2024 (N_2024,N_1811,N_1699);
and U2025 (N_2025,N_1690,N_1892);
or U2026 (N_2026,N_1952,N_1646);
nor U2027 (N_2027,N_1866,N_1722);
and U2028 (N_2028,N_1601,N_1664);
nor U2029 (N_2029,N_1762,N_1781);
xnor U2030 (N_2030,N_1962,N_1640);
and U2031 (N_2031,N_1533,N_1715);
nand U2032 (N_2032,N_1666,N_1904);
nand U2033 (N_2033,N_1500,N_1812);
nand U2034 (N_2034,N_1783,N_1974);
and U2035 (N_2035,N_1663,N_1906);
xnor U2036 (N_2036,N_1969,N_1766);
or U2037 (N_2037,N_1817,N_1882);
nor U2038 (N_2038,N_1879,N_1873);
and U2039 (N_2039,N_1644,N_1550);
nand U2040 (N_2040,N_1735,N_1815);
nand U2041 (N_2041,N_1727,N_1858);
nand U2042 (N_2042,N_1836,N_1990);
and U2043 (N_2043,N_1567,N_1606);
xnor U2044 (N_2044,N_1583,N_1957);
nand U2045 (N_2045,N_1876,N_1810);
xnor U2046 (N_2046,N_1925,N_1502);
or U2047 (N_2047,N_1716,N_1534);
and U2048 (N_2048,N_1880,N_1750);
xor U2049 (N_2049,N_1641,N_1889);
and U2050 (N_2050,N_1599,N_1773);
nand U2051 (N_2051,N_1737,N_1823);
or U2052 (N_2052,N_1544,N_1872);
nand U2053 (N_2053,N_1513,N_1614);
or U2054 (N_2054,N_1845,N_1914);
and U2055 (N_2055,N_1569,N_1653);
nand U2056 (N_2056,N_1958,N_1616);
xor U2057 (N_2057,N_1572,N_1668);
and U2058 (N_2058,N_1701,N_1675);
or U2059 (N_2059,N_1989,N_1660);
nor U2060 (N_2060,N_1942,N_1886);
or U2061 (N_2061,N_1857,N_1752);
nand U2062 (N_2062,N_1725,N_1681);
xnor U2063 (N_2063,N_1710,N_1943);
or U2064 (N_2064,N_1504,N_1719);
and U2065 (N_2065,N_1803,N_1900);
or U2066 (N_2066,N_1765,N_1751);
and U2067 (N_2067,N_1764,N_1917);
xor U2068 (N_2068,N_1759,N_1687);
and U2069 (N_2069,N_1888,N_1867);
xnor U2070 (N_2070,N_1789,N_1907);
and U2071 (N_2071,N_1568,N_1902);
xnor U2072 (N_2072,N_1590,N_1594);
xor U2073 (N_2073,N_1932,N_1724);
or U2074 (N_2074,N_1931,N_1827);
and U2075 (N_2075,N_1506,N_1778);
nand U2076 (N_2076,N_1949,N_1680);
nand U2077 (N_2077,N_1887,N_1784);
nand U2078 (N_2078,N_1656,N_1945);
or U2079 (N_2079,N_1947,N_1704);
xor U2080 (N_2080,N_1825,N_1545);
nor U2081 (N_2081,N_1634,N_1624);
or U2082 (N_2082,N_1679,N_1537);
nor U2083 (N_2083,N_1794,N_1856);
or U2084 (N_2084,N_1961,N_1939);
or U2085 (N_2085,N_1553,N_1578);
nand U2086 (N_2086,N_1530,N_1515);
or U2087 (N_2087,N_1871,N_1982);
xor U2088 (N_2088,N_1560,N_1685);
nor U2089 (N_2089,N_1985,N_1520);
nand U2090 (N_2090,N_1518,N_1726);
nand U2091 (N_2091,N_1785,N_1527);
nor U2092 (N_2092,N_1673,N_1528);
xnor U2093 (N_2093,N_1977,N_1746);
nor U2094 (N_2094,N_1779,N_1582);
and U2095 (N_2095,N_1754,N_1870);
nand U2096 (N_2096,N_1993,N_1635);
nand U2097 (N_2097,N_1909,N_1531);
or U2098 (N_2098,N_1563,N_1960);
and U2099 (N_2099,N_1566,N_1884);
xor U2100 (N_2100,N_1562,N_1611);
xnor U2101 (N_2101,N_1649,N_1877);
and U2102 (N_2102,N_1539,N_1503);
nand U2103 (N_2103,N_1693,N_1542);
and U2104 (N_2104,N_1736,N_1878);
nor U2105 (N_2105,N_1901,N_1995);
nand U2106 (N_2106,N_1841,N_1721);
xor U2107 (N_2107,N_1881,N_1944);
or U2108 (N_2108,N_1950,N_1508);
and U2109 (N_2109,N_1755,N_1692);
nand U2110 (N_2110,N_1592,N_1547);
or U2111 (N_2111,N_1775,N_1529);
or U2112 (N_2112,N_1786,N_1820);
or U2113 (N_2113,N_1740,N_1729);
nand U2114 (N_2114,N_1731,N_1795);
xor U2115 (N_2115,N_1512,N_1670);
nand U2116 (N_2116,N_1637,N_1638);
and U2117 (N_2117,N_1580,N_1659);
nand U2118 (N_2118,N_1757,N_1849);
nand U2119 (N_2119,N_1797,N_1626);
and U2120 (N_2120,N_1564,N_1921);
or U2121 (N_2121,N_1851,N_1587);
or U2122 (N_2122,N_1593,N_1749);
and U2123 (N_2123,N_1602,N_1672);
and U2124 (N_2124,N_1862,N_1898);
nor U2125 (N_2125,N_1813,N_1926);
nand U2126 (N_2126,N_1767,N_1806);
nor U2127 (N_2127,N_1745,N_1523);
nor U2128 (N_2128,N_1922,N_1853);
xor U2129 (N_2129,N_1792,N_1585);
nor U2130 (N_2130,N_1541,N_1657);
and U2131 (N_2131,N_1891,N_1645);
nor U2132 (N_2132,N_1584,N_1991);
nor U2133 (N_2133,N_1621,N_1963);
xnor U2134 (N_2134,N_1604,N_1610);
nand U2135 (N_2135,N_1920,N_1627);
and U2136 (N_2136,N_1632,N_1554);
nand U2137 (N_2137,N_1896,N_1782);
and U2138 (N_2138,N_1835,N_1814);
xnor U2139 (N_2139,N_1935,N_1697);
and U2140 (N_2140,N_1575,N_1992);
xnor U2141 (N_2141,N_1658,N_1756);
nor U2142 (N_2142,N_1965,N_1865);
and U2143 (N_2143,N_1682,N_1966);
xnor U2144 (N_2144,N_1622,N_1801);
or U2145 (N_2145,N_1705,N_1608);
xor U2146 (N_2146,N_1739,N_1908);
or U2147 (N_2147,N_1702,N_1591);
or U2148 (N_2148,N_1543,N_1595);
nor U2149 (N_2149,N_1929,N_1696);
nand U2150 (N_2150,N_1863,N_1574);
nand U2151 (N_2151,N_1717,N_1984);
nand U2152 (N_2152,N_1761,N_1654);
nor U2153 (N_2153,N_1625,N_1631);
or U2154 (N_2154,N_1915,N_1748);
nand U2155 (N_2155,N_1796,N_1706);
or U2156 (N_2156,N_1581,N_1885);
nand U2157 (N_2157,N_1973,N_1890);
and U2158 (N_2158,N_1774,N_1517);
nor U2159 (N_2159,N_1830,N_1662);
nand U2160 (N_2160,N_1938,N_1596);
and U2161 (N_2161,N_1838,N_1674);
nand U2162 (N_2162,N_1953,N_1633);
nor U2163 (N_2163,N_1571,N_1712);
and U2164 (N_2164,N_1505,N_1916);
xor U2165 (N_2165,N_1521,N_1586);
xnor U2166 (N_2166,N_1994,N_1802);
nor U2167 (N_2167,N_1546,N_1507);
and U2168 (N_2168,N_1650,N_1522);
and U2169 (N_2169,N_1643,N_1623);
xor U2170 (N_2170,N_1532,N_1683);
and U2171 (N_2171,N_1526,N_1605);
nand U2172 (N_2172,N_1620,N_1833);
and U2173 (N_2173,N_1588,N_1874);
nor U2174 (N_2174,N_1570,N_1565);
xnor U2175 (N_2175,N_1760,N_1933);
or U2176 (N_2176,N_1981,N_1804);
and U2177 (N_2177,N_1733,N_1809);
nand U2178 (N_2178,N_1777,N_1855);
nand U2179 (N_2179,N_1609,N_1618);
nor U2180 (N_2180,N_1946,N_1589);
or U2181 (N_2181,N_1744,N_1818);
and U2182 (N_2182,N_1967,N_1846);
nor U2183 (N_2183,N_1918,N_1535);
nor U2184 (N_2184,N_1808,N_1919);
xor U2185 (N_2185,N_1600,N_1708);
and U2186 (N_2186,N_1923,N_1598);
and U2187 (N_2187,N_1839,N_1895);
or U2188 (N_2188,N_1559,N_1824);
nor U2189 (N_2189,N_1843,N_1629);
or U2190 (N_2190,N_1903,N_1805);
xnor U2191 (N_2191,N_1816,N_1768);
or U2192 (N_2192,N_1978,N_1511);
nand U2193 (N_2193,N_1648,N_1859);
xnor U2194 (N_2194,N_1875,N_1837);
nor U2195 (N_2195,N_1956,N_1951);
xor U2196 (N_2196,N_1869,N_1747);
nor U2197 (N_2197,N_1700,N_1741);
xnor U2198 (N_2198,N_1894,N_1864);
and U2199 (N_2199,N_1557,N_1713);
nor U2200 (N_2200,N_1698,N_1647);
xnor U2201 (N_2201,N_1799,N_1850);
nand U2202 (N_2202,N_1577,N_1999);
nor U2203 (N_2203,N_1597,N_1897);
and U2204 (N_2204,N_1753,N_1519);
and U2205 (N_2205,N_1684,N_1667);
or U2206 (N_2206,N_1671,N_1636);
or U2207 (N_2207,N_1927,N_1930);
nor U2208 (N_2208,N_1763,N_1561);
or U2209 (N_2209,N_1607,N_1997);
xor U2210 (N_2210,N_1910,N_1979);
xnor U2211 (N_2211,N_1819,N_1770);
nor U2212 (N_2212,N_1791,N_1612);
nand U2213 (N_2213,N_1842,N_1720);
and U2214 (N_2214,N_1828,N_1555);
and U2215 (N_2215,N_1912,N_1516);
and U2216 (N_2216,N_1976,N_1728);
nand U2217 (N_2217,N_1711,N_1514);
and U2218 (N_2218,N_1639,N_1787);
or U2219 (N_2219,N_1772,N_1714);
and U2220 (N_2220,N_1576,N_1854);
nand U2221 (N_2221,N_1691,N_1971);
and U2222 (N_2222,N_1678,N_1970);
nor U2223 (N_2223,N_1852,N_1771);
nand U2224 (N_2224,N_1538,N_1677);
xor U2225 (N_2225,N_1603,N_1883);
or U2226 (N_2226,N_1798,N_1996);
nor U2227 (N_2227,N_1899,N_1924);
and U2228 (N_2228,N_1893,N_1860);
xnor U2229 (N_2229,N_1619,N_1807);
xor U2230 (N_2230,N_1955,N_1934);
nor U2231 (N_2231,N_1734,N_1788);
nand U2232 (N_2232,N_1913,N_1525);
or U2233 (N_2233,N_1980,N_1936);
or U2234 (N_2234,N_1940,N_1954);
or U2235 (N_2235,N_1732,N_1972);
or U2236 (N_2236,N_1968,N_1510);
nor U2237 (N_2237,N_1840,N_1615);
or U2238 (N_2238,N_1790,N_1986);
nor U2239 (N_2239,N_1718,N_1661);
xnor U2240 (N_2240,N_1695,N_1975);
or U2241 (N_2241,N_1769,N_1703);
or U2242 (N_2242,N_1905,N_1651);
nand U2243 (N_2243,N_1822,N_1501);
xor U2244 (N_2244,N_1676,N_1642);
nor U2245 (N_2245,N_1826,N_1628);
nand U2246 (N_2246,N_1848,N_1709);
and U2247 (N_2247,N_1723,N_1821);
nand U2248 (N_2248,N_1941,N_1911);
or U2249 (N_2249,N_1844,N_1617);
and U2250 (N_2250,N_1506,N_1797);
and U2251 (N_2251,N_1834,N_1625);
nor U2252 (N_2252,N_1975,N_1946);
xor U2253 (N_2253,N_1758,N_1915);
xor U2254 (N_2254,N_1997,N_1549);
nand U2255 (N_2255,N_1783,N_1990);
or U2256 (N_2256,N_1641,N_1610);
or U2257 (N_2257,N_1584,N_1997);
and U2258 (N_2258,N_1976,N_1908);
and U2259 (N_2259,N_1928,N_1562);
nor U2260 (N_2260,N_1555,N_1962);
nor U2261 (N_2261,N_1615,N_1504);
nor U2262 (N_2262,N_1883,N_1558);
and U2263 (N_2263,N_1934,N_1727);
or U2264 (N_2264,N_1722,N_1959);
xor U2265 (N_2265,N_1508,N_1696);
or U2266 (N_2266,N_1670,N_1806);
xnor U2267 (N_2267,N_1915,N_1859);
nor U2268 (N_2268,N_1723,N_1625);
and U2269 (N_2269,N_1661,N_1700);
nor U2270 (N_2270,N_1676,N_1651);
or U2271 (N_2271,N_1539,N_1924);
and U2272 (N_2272,N_1700,N_1569);
xor U2273 (N_2273,N_1983,N_1550);
xor U2274 (N_2274,N_1822,N_1519);
nand U2275 (N_2275,N_1698,N_1507);
and U2276 (N_2276,N_1824,N_1882);
nand U2277 (N_2277,N_1725,N_1502);
xnor U2278 (N_2278,N_1866,N_1527);
and U2279 (N_2279,N_1829,N_1873);
and U2280 (N_2280,N_1506,N_1580);
nor U2281 (N_2281,N_1670,N_1797);
nand U2282 (N_2282,N_1551,N_1842);
and U2283 (N_2283,N_1657,N_1672);
and U2284 (N_2284,N_1548,N_1755);
nand U2285 (N_2285,N_1769,N_1545);
xnor U2286 (N_2286,N_1765,N_1738);
or U2287 (N_2287,N_1655,N_1548);
xnor U2288 (N_2288,N_1964,N_1920);
or U2289 (N_2289,N_1947,N_1715);
nand U2290 (N_2290,N_1550,N_1828);
nor U2291 (N_2291,N_1562,N_1595);
xor U2292 (N_2292,N_1825,N_1570);
xor U2293 (N_2293,N_1640,N_1738);
xnor U2294 (N_2294,N_1721,N_1663);
xor U2295 (N_2295,N_1933,N_1959);
nand U2296 (N_2296,N_1856,N_1820);
nor U2297 (N_2297,N_1554,N_1644);
nand U2298 (N_2298,N_1879,N_1943);
and U2299 (N_2299,N_1768,N_1676);
and U2300 (N_2300,N_1674,N_1809);
nor U2301 (N_2301,N_1508,N_1639);
and U2302 (N_2302,N_1641,N_1545);
and U2303 (N_2303,N_1657,N_1832);
xnor U2304 (N_2304,N_1822,N_1810);
and U2305 (N_2305,N_1761,N_1948);
xnor U2306 (N_2306,N_1628,N_1859);
nor U2307 (N_2307,N_1917,N_1527);
nor U2308 (N_2308,N_1968,N_1863);
or U2309 (N_2309,N_1665,N_1537);
nand U2310 (N_2310,N_1509,N_1814);
or U2311 (N_2311,N_1898,N_1732);
nor U2312 (N_2312,N_1927,N_1698);
and U2313 (N_2313,N_1761,N_1543);
nor U2314 (N_2314,N_1693,N_1886);
nand U2315 (N_2315,N_1915,N_1670);
nor U2316 (N_2316,N_1834,N_1634);
and U2317 (N_2317,N_1532,N_1579);
nand U2318 (N_2318,N_1813,N_1839);
nor U2319 (N_2319,N_1721,N_1803);
nor U2320 (N_2320,N_1670,N_1864);
nand U2321 (N_2321,N_1757,N_1905);
nor U2322 (N_2322,N_1675,N_1671);
and U2323 (N_2323,N_1938,N_1676);
xor U2324 (N_2324,N_1799,N_1952);
or U2325 (N_2325,N_1970,N_1831);
or U2326 (N_2326,N_1725,N_1691);
or U2327 (N_2327,N_1930,N_1811);
and U2328 (N_2328,N_1671,N_1644);
nor U2329 (N_2329,N_1674,N_1662);
nand U2330 (N_2330,N_1519,N_1817);
and U2331 (N_2331,N_1665,N_1616);
and U2332 (N_2332,N_1925,N_1616);
and U2333 (N_2333,N_1897,N_1732);
nor U2334 (N_2334,N_1992,N_1665);
nor U2335 (N_2335,N_1857,N_1799);
and U2336 (N_2336,N_1776,N_1571);
or U2337 (N_2337,N_1533,N_1878);
nand U2338 (N_2338,N_1778,N_1576);
nor U2339 (N_2339,N_1791,N_1543);
or U2340 (N_2340,N_1954,N_1644);
nand U2341 (N_2341,N_1998,N_1969);
xor U2342 (N_2342,N_1777,N_1553);
or U2343 (N_2343,N_1847,N_1525);
nand U2344 (N_2344,N_1807,N_1655);
xnor U2345 (N_2345,N_1650,N_1594);
xor U2346 (N_2346,N_1900,N_1870);
nand U2347 (N_2347,N_1970,N_1999);
nor U2348 (N_2348,N_1807,N_1586);
xnor U2349 (N_2349,N_1900,N_1907);
nand U2350 (N_2350,N_1951,N_1804);
nor U2351 (N_2351,N_1517,N_1745);
and U2352 (N_2352,N_1844,N_1759);
nor U2353 (N_2353,N_1922,N_1701);
and U2354 (N_2354,N_1719,N_1653);
xor U2355 (N_2355,N_1741,N_1767);
nand U2356 (N_2356,N_1741,N_1555);
nor U2357 (N_2357,N_1541,N_1804);
xor U2358 (N_2358,N_1532,N_1688);
and U2359 (N_2359,N_1951,N_1845);
xnor U2360 (N_2360,N_1997,N_1861);
or U2361 (N_2361,N_1665,N_1792);
and U2362 (N_2362,N_1521,N_1601);
xnor U2363 (N_2363,N_1653,N_1547);
and U2364 (N_2364,N_1872,N_1536);
nand U2365 (N_2365,N_1871,N_1764);
or U2366 (N_2366,N_1704,N_1899);
xor U2367 (N_2367,N_1788,N_1773);
xnor U2368 (N_2368,N_1953,N_1815);
and U2369 (N_2369,N_1742,N_1920);
or U2370 (N_2370,N_1893,N_1595);
nor U2371 (N_2371,N_1852,N_1717);
xor U2372 (N_2372,N_1503,N_1840);
or U2373 (N_2373,N_1597,N_1714);
nor U2374 (N_2374,N_1912,N_1908);
nor U2375 (N_2375,N_1686,N_1646);
xnor U2376 (N_2376,N_1541,N_1871);
nand U2377 (N_2377,N_1721,N_1633);
and U2378 (N_2378,N_1929,N_1978);
and U2379 (N_2379,N_1542,N_1870);
and U2380 (N_2380,N_1592,N_1767);
nand U2381 (N_2381,N_1616,N_1831);
or U2382 (N_2382,N_1710,N_1981);
nand U2383 (N_2383,N_1910,N_1958);
or U2384 (N_2384,N_1729,N_1628);
xnor U2385 (N_2385,N_1909,N_1658);
and U2386 (N_2386,N_1794,N_1792);
nand U2387 (N_2387,N_1604,N_1883);
nor U2388 (N_2388,N_1764,N_1695);
nor U2389 (N_2389,N_1752,N_1732);
nor U2390 (N_2390,N_1535,N_1919);
or U2391 (N_2391,N_1522,N_1513);
xor U2392 (N_2392,N_1945,N_1963);
xnor U2393 (N_2393,N_1648,N_1512);
nor U2394 (N_2394,N_1709,N_1772);
xnor U2395 (N_2395,N_1986,N_1749);
xnor U2396 (N_2396,N_1748,N_1867);
xnor U2397 (N_2397,N_1633,N_1854);
and U2398 (N_2398,N_1630,N_1703);
xnor U2399 (N_2399,N_1652,N_1838);
or U2400 (N_2400,N_1748,N_1589);
or U2401 (N_2401,N_1609,N_1674);
nand U2402 (N_2402,N_1869,N_1515);
nor U2403 (N_2403,N_1845,N_1915);
xor U2404 (N_2404,N_1558,N_1661);
xnor U2405 (N_2405,N_1823,N_1837);
or U2406 (N_2406,N_1601,N_1957);
nor U2407 (N_2407,N_1621,N_1657);
nor U2408 (N_2408,N_1787,N_1926);
and U2409 (N_2409,N_1559,N_1964);
xor U2410 (N_2410,N_1773,N_1886);
nand U2411 (N_2411,N_1867,N_1599);
and U2412 (N_2412,N_1628,N_1828);
nor U2413 (N_2413,N_1542,N_1546);
xnor U2414 (N_2414,N_1746,N_1649);
or U2415 (N_2415,N_1763,N_1940);
xnor U2416 (N_2416,N_1689,N_1609);
nand U2417 (N_2417,N_1759,N_1736);
nand U2418 (N_2418,N_1937,N_1600);
or U2419 (N_2419,N_1625,N_1646);
xor U2420 (N_2420,N_1614,N_1920);
nand U2421 (N_2421,N_1518,N_1934);
or U2422 (N_2422,N_1774,N_1983);
xor U2423 (N_2423,N_1801,N_1838);
nand U2424 (N_2424,N_1870,N_1764);
nor U2425 (N_2425,N_1916,N_1861);
nand U2426 (N_2426,N_1613,N_1827);
nor U2427 (N_2427,N_1518,N_1832);
or U2428 (N_2428,N_1569,N_1932);
or U2429 (N_2429,N_1697,N_1565);
nand U2430 (N_2430,N_1567,N_1871);
xor U2431 (N_2431,N_1574,N_1615);
and U2432 (N_2432,N_1792,N_1851);
and U2433 (N_2433,N_1670,N_1834);
xor U2434 (N_2434,N_1858,N_1503);
and U2435 (N_2435,N_1711,N_1740);
and U2436 (N_2436,N_1836,N_1694);
nor U2437 (N_2437,N_1865,N_1911);
nand U2438 (N_2438,N_1597,N_1789);
nand U2439 (N_2439,N_1503,N_1694);
nor U2440 (N_2440,N_1911,N_1818);
xor U2441 (N_2441,N_1664,N_1989);
nor U2442 (N_2442,N_1840,N_1732);
nor U2443 (N_2443,N_1515,N_1764);
or U2444 (N_2444,N_1799,N_1898);
xor U2445 (N_2445,N_1811,N_1531);
nor U2446 (N_2446,N_1892,N_1528);
nor U2447 (N_2447,N_1722,N_1770);
or U2448 (N_2448,N_1809,N_1938);
xnor U2449 (N_2449,N_1773,N_1614);
xnor U2450 (N_2450,N_1999,N_1934);
nor U2451 (N_2451,N_1882,N_1503);
and U2452 (N_2452,N_1663,N_1583);
nor U2453 (N_2453,N_1918,N_1908);
and U2454 (N_2454,N_1520,N_1652);
or U2455 (N_2455,N_1586,N_1753);
nor U2456 (N_2456,N_1682,N_1843);
nor U2457 (N_2457,N_1507,N_1705);
or U2458 (N_2458,N_1524,N_1514);
nor U2459 (N_2459,N_1634,N_1902);
nor U2460 (N_2460,N_1938,N_1683);
or U2461 (N_2461,N_1780,N_1666);
or U2462 (N_2462,N_1891,N_1705);
xnor U2463 (N_2463,N_1799,N_1938);
or U2464 (N_2464,N_1606,N_1602);
xnor U2465 (N_2465,N_1533,N_1528);
xor U2466 (N_2466,N_1630,N_1780);
or U2467 (N_2467,N_1710,N_1791);
nor U2468 (N_2468,N_1738,N_1959);
nor U2469 (N_2469,N_1541,N_1554);
or U2470 (N_2470,N_1916,N_1580);
xor U2471 (N_2471,N_1790,N_1646);
or U2472 (N_2472,N_1891,N_1803);
nand U2473 (N_2473,N_1631,N_1630);
nand U2474 (N_2474,N_1793,N_1598);
and U2475 (N_2475,N_1953,N_1859);
or U2476 (N_2476,N_1560,N_1858);
xnor U2477 (N_2477,N_1888,N_1980);
and U2478 (N_2478,N_1929,N_1703);
nand U2479 (N_2479,N_1761,N_1912);
or U2480 (N_2480,N_1580,N_1555);
nor U2481 (N_2481,N_1919,N_1769);
nand U2482 (N_2482,N_1585,N_1672);
and U2483 (N_2483,N_1826,N_1676);
and U2484 (N_2484,N_1625,N_1610);
or U2485 (N_2485,N_1987,N_1836);
nand U2486 (N_2486,N_1637,N_1873);
xnor U2487 (N_2487,N_1996,N_1516);
xor U2488 (N_2488,N_1791,N_1704);
and U2489 (N_2489,N_1990,N_1676);
and U2490 (N_2490,N_1752,N_1628);
nand U2491 (N_2491,N_1984,N_1989);
nand U2492 (N_2492,N_1695,N_1794);
nor U2493 (N_2493,N_1986,N_1750);
nor U2494 (N_2494,N_1855,N_1709);
nand U2495 (N_2495,N_1722,N_1973);
or U2496 (N_2496,N_1686,N_1871);
nand U2497 (N_2497,N_1557,N_1613);
nor U2498 (N_2498,N_1867,N_1568);
xor U2499 (N_2499,N_1964,N_1781);
or U2500 (N_2500,N_2300,N_2098);
and U2501 (N_2501,N_2186,N_2088);
and U2502 (N_2502,N_2283,N_2101);
xnor U2503 (N_2503,N_2016,N_2335);
xnor U2504 (N_2504,N_2245,N_2498);
nand U2505 (N_2505,N_2272,N_2151);
and U2506 (N_2506,N_2261,N_2127);
nand U2507 (N_2507,N_2441,N_2213);
xnor U2508 (N_2508,N_2246,N_2103);
xnor U2509 (N_2509,N_2327,N_2291);
xor U2510 (N_2510,N_2138,N_2466);
nand U2511 (N_2511,N_2275,N_2135);
nor U2512 (N_2512,N_2199,N_2323);
xnor U2513 (N_2513,N_2144,N_2414);
nand U2514 (N_2514,N_2375,N_2284);
or U2515 (N_2515,N_2399,N_2411);
nand U2516 (N_2516,N_2480,N_2294);
or U2517 (N_2517,N_2482,N_2126);
or U2518 (N_2518,N_2195,N_2171);
nor U2519 (N_2519,N_2212,N_2044);
xnor U2520 (N_2520,N_2439,N_2232);
xor U2521 (N_2521,N_2258,N_2386);
nand U2522 (N_2522,N_2393,N_2129);
nor U2523 (N_2523,N_2106,N_2351);
nand U2524 (N_2524,N_2379,N_2024);
and U2525 (N_2525,N_2249,N_2389);
and U2526 (N_2526,N_2167,N_2119);
or U2527 (N_2527,N_2049,N_2009);
and U2528 (N_2528,N_2188,N_2087);
and U2529 (N_2529,N_2125,N_2419);
nor U2530 (N_2530,N_2429,N_2421);
or U2531 (N_2531,N_2256,N_2054);
and U2532 (N_2532,N_2316,N_2394);
xnor U2533 (N_2533,N_2006,N_2209);
nor U2534 (N_2534,N_2180,N_2083);
and U2535 (N_2535,N_2364,N_2196);
xnor U2536 (N_2536,N_2168,N_2069);
nor U2537 (N_2537,N_2346,N_2056);
xor U2538 (N_2538,N_2432,N_2293);
nor U2539 (N_2539,N_2184,N_2035);
or U2540 (N_2540,N_2499,N_2365);
nor U2541 (N_2541,N_2207,N_2469);
and U2542 (N_2542,N_2002,N_2095);
and U2543 (N_2543,N_2325,N_2476);
nor U2544 (N_2544,N_2118,N_2107);
nand U2545 (N_2545,N_2005,N_2483);
nand U2546 (N_2546,N_2315,N_2128);
nor U2547 (N_2547,N_2440,N_2100);
and U2548 (N_2548,N_2001,N_2113);
nor U2549 (N_2549,N_2401,N_2084);
or U2550 (N_2550,N_2121,N_2430);
nand U2551 (N_2551,N_2241,N_2431);
or U2552 (N_2552,N_2099,N_2442);
nand U2553 (N_2553,N_2392,N_2165);
and U2554 (N_2554,N_2051,N_2285);
or U2555 (N_2555,N_2079,N_2175);
or U2556 (N_2556,N_2455,N_2475);
or U2557 (N_2557,N_2277,N_2021);
nor U2558 (N_2558,N_2355,N_2398);
or U2559 (N_2559,N_2090,N_2273);
and U2560 (N_2560,N_2173,N_2182);
xnor U2561 (N_2561,N_2307,N_2260);
nor U2562 (N_2562,N_2230,N_2486);
nand U2563 (N_2563,N_2117,N_2202);
nor U2564 (N_2564,N_2141,N_2048);
nand U2565 (N_2565,N_2003,N_2072);
xor U2566 (N_2566,N_2437,N_2022);
or U2567 (N_2567,N_2359,N_2336);
and U2568 (N_2568,N_2136,N_2251);
nor U2569 (N_2569,N_2221,N_2370);
or U2570 (N_2570,N_2176,N_2050);
nand U2571 (N_2571,N_2259,N_2211);
or U2572 (N_2572,N_2218,N_2491);
nor U2573 (N_2573,N_2114,N_2318);
and U2574 (N_2574,N_2362,N_2492);
xnor U2575 (N_2575,N_2229,N_2228);
nor U2576 (N_2576,N_2185,N_2381);
and U2577 (N_2577,N_2073,N_2013);
nor U2578 (N_2578,N_2155,N_2289);
nor U2579 (N_2579,N_2243,N_2080);
or U2580 (N_2580,N_2322,N_2027);
nand U2581 (N_2581,N_2280,N_2250);
nand U2582 (N_2582,N_2326,N_2481);
or U2583 (N_2583,N_2309,N_2342);
and U2584 (N_2584,N_2004,N_2148);
or U2585 (N_2585,N_2158,N_2248);
xnor U2586 (N_2586,N_2308,N_2093);
and U2587 (N_2587,N_2063,N_2296);
nor U2588 (N_2588,N_2410,N_2385);
and U2589 (N_2589,N_2029,N_2210);
nor U2590 (N_2590,N_2357,N_2298);
nand U2591 (N_2591,N_2270,N_2131);
and U2592 (N_2592,N_2060,N_2075);
nand U2593 (N_2593,N_2216,N_2488);
and U2594 (N_2594,N_2038,N_2062);
xnor U2595 (N_2595,N_2409,N_2124);
nor U2596 (N_2596,N_2434,N_2407);
nor U2597 (N_2597,N_2007,N_2337);
or U2598 (N_2598,N_2091,N_2425);
nor U2599 (N_2599,N_2467,N_2137);
nor U2600 (N_2600,N_2263,N_2052);
nor U2601 (N_2601,N_2462,N_2017);
or U2602 (N_2602,N_2164,N_2339);
and U2603 (N_2603,N_2019,N_2163);
and U2604 (N_2604,N_2169,N_2082);
xnor U2605 (N_2605,N_2329,N_2122);
or U2606 (N_2606,N_2478,N_2067);
nor U2607 (N_2607,N_2376,N_2380);
xnor U2608 (N_2608,N_2227,N_2404);
and U2609 (N_2609,N_2406,N_2239);
nor U2610 (N_2610,N_2479,N_2085);
and U2611 (N_2611,N_2402,N_2189);
and U2612 (N_2612,N_2115,N_2110);
nand U2613 (N_2613,N_2340,N_2426);
nand U2614 (N_2614,N_2485,N_2287);
nand U2615 (N_2615,N_2240,N_2142);
xnor U2616 (N_2616,N_2278,N_2383);
or U2617 (N_2617,N_2266,N_2147);
or U2618 (N_2618,N_2116,N_2094);
xnor U2619 (N_2619,N_2449,N_2276);
and U2620 (N_2620,N_2301,N_2178);
or U2621 (N_2621,N_2360,N_2153);
and U2622 (N_2622,N_2310,N_2053);
and U2623 (N_2623,N_2020,N_2377);
xnor U2624 (N_2624,N_2205,N_2015);
xor U2625 (N_2625,N_2368,N_2388);
nor U2626 (N_2626,N_2371,N_2254);
or U2627 (N_2627,N_2162,N_2448);
xor U2628 (N_2628,N_2288,N_2030);
and U2629 (N_2629,N_2460,N_2384);
nor U2630 (N_2630,N_2338,N_2233);
nor U2631 (N_2631,N_2474,N_2219);
nor U2632 (N_2632,N_2279,N_2252);
or U2633 (N_2633,N_2369,N_2343);
xor U2634 (N_2634,N_2495,N_2302);
nor U2635 (N_2635,N_2197,N_2281);
nand U2636 (N_2636,N_2292,N_2286);
nor U2637 (N_2637,N_2235,N_2299);
or U2638 (N_2638,N_2070,N_2000);
xor U2639 (N_2639,N_2076,N_2452);
and U2640 (N_2640,N_2472,N_2012);
xnor U2641 (N_2641,N_2156,N_2496);
nand U2642 (N_2642,N_2026,N_2011);
or U2643 (N_2643,N_2031,N_2344);
nand U2644 (N_2644,N_2317,N_2454);
or U2645 (N_2645,N_2313,N_2405);
and U2646 (N_2646,N_2459,N_2255);
xor U2647 (N_2647,N_2217,N_2191);
or U2648 (N_2648,N_2390,N_2133);
xnor U2649 (N_2649,N_2105,N_2428);
and U2650 (N_2650,N_2367,N_2304);
or U2651 (N_2651,N_2159,N_2174);
and U2652 (N_2652,N_2046,N_2071);
and U2653 (N_2653,N_2427,N_2413);
nand U2654 (N_2654,N_2477,N_2445);
nand U2655 (N_2655,N_2059,N_2161);
nand U2656 (N_2656,N_2305,N_2201);
nand U2657 (N_2657,N_2458,N_2081);
and U2658 (N_2658,N_2444,N_2424);
xor U2659 (N_2659,N_2181,N_2443);
nand U2660 (N_2660,N_2193,N_2214);
or U2661 (N_2661,N_2352,N_2416);
nand U2662 (N_2662,N_2366,N_2264);
and U2663 (N_2663,N_2215,N_2463);
nand U2664 (N_2664,N_2014,N_2403);
xor U2665 (N_2665,N_2297,N_2010);
xnor U2666 (N_2666,N_2055,N_2267);
nand U2667 (N_2667,N_2350,N_2047);
or U2668 (N_2668,N_2238,N_2490);
and U2669 (N_2669,N_2036,N_2420);
or U2670 (N_2670,N_2282,N_2374);
and U2671 (N_2671,N_2065,N_2331);
and U2672 (N_2672,N_2236,N_2453);
nand U2673 (N_2673,N_2349,N_2077);
nand U2674 (N_2674,N_2450,N_2032);
nor U2675 (N_2675,N_2456,N_2412);
nor U2676 (N_2676,N_2130,N_2311);
nand U2677 (N_2677,N_2111,N_2037);
and U2678 (N_2678,N_2231,N_2324);
nand U2679 (N_2679,N_2451,N_2008);
and U2680 (N_2680,N_2068,N_2089);
nor U2681 (N_2681,N_2348,N_2319);
or U2682 (N_2682,N_2493,N_2391);
nor U2683 (N_2683,N_2150,N_2358);
nor U2684 (N_2684,N_2226,N_2222);
nor U2685 (N_2685,N_2372,N_2320);
xor U2686 (N_2686,N_2224,N_2345);
or U2687 (N_2687,N_2435,N_2108);
and U2688 (N_2688,N_2166,N_2061);
and U2689 (N_2689,N_2058,N_2306);
nor U2690 (N_2690,N_2265,N_2200);
nand U2691 (N_2691,N_2045,N_2109);
nand U2692 (N_2692,N_2400,N_2314);
nand U2693 (N_2693,N_2271,N_2198);
nor U2694 (N_2694,N_2208,N_2187);
xor U2695 (N_2695,N_2387,N_2225);
and U2696 (N_2696,N_2157,N_2112);
nor U2697 (N_2697,N_2494,N_2041);
or U2698 (N_2698,N_2123,N_2033);
nand U2699 (N_2699,N_2097,N_2042);
and U2700 (N_2700,N_2134,N_2183);
nor U2701 (N_2701,N_2057,N_2465);
nor U2702 (N_2702,N_2417,N_2464);
nand U2703 (N_2703,N_2330,N_2312);
xnor U2704 (N_2704,N_2332,N_2034);
or U2705 (N_2705,N_2253,N_2146);
nand U2706 (N_2706,N_2023,N_2096);
or U2707 (N_2707,N_2237,N_2489);
nor U2708 (N_2708,N_2497,N_2074);
xor U2709 (N_2709,N_2356,N_2086);
or U2710 (N_2710,N_2039,N_2192);
and U2711 (N_2711,N_2220,N_2139);
or U2712 (N_2712,N_2064,N_2447);
nand U2713 (N_2713,N_2132,N_2018);
xor U2714 (N_2714,N_2484,N_2396);
and U2715 (N_2715,N_2242,N_2177);
xor U2716 (N_2716,N_2363,N_2204);
xnor U2717 (N_2717,N_2149,N_2234);
xor U2718 (N_2718,N_2382,N_2361);
nor U2719 (N_2719,N_2334,N_2223);
and U2720 (N_2720,N_2341,N_2154);
and U2721 (N_2721,N_2418,N_2333);
nand U2722 (N_2722,N_2152,N_2397);
nand U2723 (N_2723,N_2354,N_2028);
or U2724 (N_2724,N_2078,N_2347);
xnor U2725 (N_2725,N_2470,N_2143);
nand U2726 (N_2726,N_2247,N_2395);
and U2727 (N_2727,N_2257,N_2303);
or U2728 (N_2728,N_2269,N_2025);
xnor U2729 (N_2729,N_2433,N_2160);
and U2730 (N_2730,N_2203,N_2408);
xor U2731 (N_2731,N_2244,N_2066);
nor U2732 (N_2732,N_2274,N_2092);
nor U2733 (N_2733,N_2206,N_2487);
nor U2734 (N_2734,N_2194,N_2295);
and U2735 (N_2735,N_2104,N_2102);
xor U2736 (N_2736,N_2378,N_2415);
and U2737 (N_2737,N_2373,N_2268);
nand U2738 (N_2738,N_2473,N_2461);
nand U2739 (N_2739,N_2040,N_2043);
nand U2740 (N_2740,N_2170,N_2120);
and U2741 (N_2741,N_2436,N_2353);
or U2742 (N_2742,N_2321,N_2471);
and U2743 (N_2743,N_2422,N_2423);
nor U2744 (N_2744,N_2140,N_2290);
nand U2745 (N_2745,N_2190,N_2468);
nor U2746 (N_2746,N_2328,N_2446);
and U2747 (N_2747,N_2262,N_2457);
nor U2748 (N_2748,N_2172,N_2438);
xnor U2749 (N_2749,N_2145,N_2179);
or U2750 (N_2750,N_2205,N_2068);
xor U2751 (N_2751,N_2276,N_2338);
nor U2752 (N_2752,N_2217,N_2458);
and U2753 (N_2753,N_2330,N_2268);
xnor U2754 (N_2754,N_2222,N_2178);
or U2755 (N_2755,N_2198,N_2275);
xor U2756 (N_2756,N_2255,N_2238);
xnor U2757 (N_2757,N_2053,N_2126);
or U2758 (N_2758,N_2082,N_2407);
nor U2759 (N_2759,N_2001,N_2179);
nand U2760 (N_2760,N_2162,N_2289);
or U2761 (N_2761,N_2315,N_2019);
and U2762 (N_2762,N_2419,N_2355);
nor U2763 (N_2763,N_2432,N_2273);
or U2764 (N_2764,N_2107,N_2295);
xor U2765 (N_2765,N_2207,N_2333);
or U2766 (N_2766,N_2252,N_2483);
or U2767 (N_2767,N_2481,N_2216);
nand U2768 (N_2768,N_2205,N_2141);
and U2769 (N_2769,N_2103,N_2414);
xor U2770 (N_2770,N_2007,N_2228);
nand U2771 (N_2771,N_2245,N_2499);
xor U2772 (N_2772,N_2172,N_2243);
and U2773 (N_2773,N_2439,N_2211);
or U2774 (N_2774,N_2046,N_2237);
and U2775 (N_2775,N_2370,N_2397);
nor U2776 (N_2776,N_2124,N_2498);
and U2777 (N_2777,N_2324,N_2004);
and U2778 (N_2778,N_2451,N_2011);
nand U2779 (N_2779,N_2205,N_2206);
xor U2780 (N_2780,N_2147,N_2035);
xor U2781 (N_2781,N_2109,N_2139);
and U2782 (N_2782,N_2309,N_2156);
nand U2783 (N_2783,N_2495,N_2161);
and U2784 (N_2784,N_2245,N_2351);
nor U2785 (N_2785,N_2163,N_2161);
and U2786 (N_2786,N_2080,N_2137);
nand U2787 (N_2787,N_2187,N_2076);
and U2788 (N_2788,N_2247,N_2167);
or U2789 (N_2789,N_2000,N_2382);
xnor U2790 (N_2790,N_2239,N_2232);
nor U2791 (N_2791,N_2119,N_2310);
nor U2792 (N_2792,N_2165,N_2388);
nor U2793 (N_2793,N_2096,N_2339);
and U2794 (N_2794,N_2497,N_2458);
nor U2795 (N_2795,N_2493,N_2207);
and U2796 (N_2796,N_2337,N_2403);
and U2797 (N_2797,N_2310,N_2332);
or U2798 (N_2798,N_2171,N_2109);
nand U2799 (N_2799,N_2440,N_2321);
xnor U2800 (N_2800,N_2396,N_2439);
or U2801 (N_2801,N_2353,N_2477);
nand U2802 (N_2802,N_2369,N_2169);
nor U2803 (N_2803,N_2254,N_2462);
xnor U2804 (N_2804,N_2140,N_2399);
and U2805 (N_2805,N_2206,N_2071);
nand U2806 (N_2806,N_2429,N_2206);
nor U2807 (N_2807,N_2062,N_2129);
and U2808 (N_2808,N_2330,N_2429);
and U2809 (N_2809,N_2009,N_2495);
nor U2810 (N_2810,N_2194,N_2354);
xnor U2811 (N_2811,N_2164,N_2052);
nor U2812 (N_2812,N_2163,N_2403);
or U2813 (N_2813,N_2497,N_2073);
and U2814 (N_2814,N_2069,N_2072);
or U2815 (N_2815,N_2208,N_2473);
and U2816 (N_2816,N_2259,N_2001);
xor U2817 (N_2817,N_2485,N_2411);
nor U2818 (N_2818,N_2432,N_2177);
xnor U2819 (N_2819,N_2371,N_2242);
and U2820 (N_2820,N_2241,N_2286);
nand U2821 (N_2821,N_2036,N_2003);
or U2822 (N_2822,N_2278,N_2146);
xnor U2823 (N_2823,N_2311,N_2389);
nor U2824 (N_2824,N_2415,N_2397);
or U2825 (N_2825,N_2326,N_2220);
xnor U2826 (N_2826,N_2396,N_2385);
and U2827 (N_2827,N_2348,N_2124);
xnor U2828 (N_2828,N_2459,N_2472);
nand U2829 (N_2829,N_2305,N_2414);
and U2830 (N_2830,N_2302,N_2304);
nor U2831 (N_2831,N_2014,N_2233);
xor U2832 (N_2832,N_2397,N_2057);
nor U2833 (N_2833,N_2403,N_2011);
xnor U2834 (N_2834,N_2269,N_2477);
nand U2835 (N_2835,N_2063,N_2161);
and U2836 (N_2836,N_2268,N_2133);
or U2837 (N_2837,N_2007,N_2385);
nor U2838 (N_2838,N_2123,N_2433);
nor U2839 (N_2839,N_2117,N_2036);
xnor U2840 (N_2840,N_2349,N_2348);
or U2841 (N_2841,N_2041,N_2352);
nor U2842 (N_2842,N_2316,N_2218);
and U2843 (N_2843,N_2362,N_2140);
and U2844 (N_2844,N_2461,N_2328);
xor U2845 (N_2845,N_2023,N_2439);
xnor U2846 (N_2846,N_2233,N_2402);
or U2847 (N_2847,N_2343,N_2274);
nor U2848 (N_2848,N_2219,N_2161);
xnor U2849 (N_2849,N_2102,N_2323);
and U2850 (N_2850,N_2117,N_2328);
or U2851 (N_2851,N_2412,N_2337);
nor U2852 (N_2852,N_2028,N_2301);
and U2853 (N_2853,N_2143,N_2370);
nand U2854 (N_2854,N_2054,N_2418);
or U2855 (N_2855,N_2424,N_2390);
and U2856 (N_2856,N_2322,N_2451);
or U2857 (N_2857,N_2150,N_2161);
and U2858 (N_2858,N_2417,N_2076);
nor U2859 (N_2859,N_2401,N_2085);
xnor U2860 (N_2860,N_2456,N_2032);
or U2861 (N_2861,N_2055,N_2487);
or U2862 (N_2862,N_2194,N_2410);
xnor U2863 (N_2863,N_2194,N_2069);
or U2864 (N_2864,N_2235,N_2344);
xnor U2865 (N_2865,N_2296,N_2175);
nand U2866 (N_2866,N_2495,N_2097);
xnor U2867 (N_2867,N_2484,N_2439);
xnor U2868 (N_2868,N_2303,N_2237);
or U2869 (N_2869,N_2167,N_2166);
xnor U2870 (N_2870,N_2339,N_2466);
or U2871 (N_2871,N_2390,N_2048);
nor U2872 (N_2872,N_2285,N_2418);
or U2873 (N_2873,N_2330,N_2347);
xor U2874 (N_2874,N_2274,N_2025);
nand U2875 (N_2875,N_2189,N_2339);
xnor U2876 (N_2876,N_2308,N_2419);
and U2877 (N_2877,N_2327,N_2439);
or U2878 (N_2878,N_2344,N_2433);
xnor U2879 (N_2879,N_2450,N_2285);
and U2880 (N_2880,N_2458,N_2328);
nor U2881 (N_2881,N_2318,N_2423);
or U2882 (N_2882,N_2421,N_2098);
or U2883 (N_2883,N_2474,N_2194);
or U2884 (N_2884,N_2407,N_2053);
xor U2885 (N_2885,N_2020,N_2437);
and U2886 (N_2886,N_2024,N_2434);
xnor U2887 (N_2887,N_2450,N_2064);
nor U2888 (N_2888,N_2474,N_2132);
or U2889 (N_2889,N_2304,N_2419);
and U2890 (N_2890,N_2412,N_2010);
nor U2891 (N_2891,N_2304,N_2213);
or U2892 (N_2892,N_2053,N_2497);
nand U2893 (N_2893,N_2035,N_2103);
or U2894 (N_2894,N_2214,N_2114);
xor U2895 (N_2895,N_2125,N_2003);
and U2896 (N_2896,N_2400,N_2249);
nand U2897 (N_2897,N_2195,N_2028);
and U2898 (N_2898,N_2270,N_2165);
and U2899 (N_2899,N_2467,N_2122);
nor U2900 (N_2900,N_2349,N_2062);
or U2901 (N_2901,N_2194,N_2209);
and U2902 (N_2902,N_2285,N_2281);
nor U2903 (N_2903,N_2040,N_2190);
xnor U2904 (N_2904,N_2206,N_2066);
and U2905 (N_2905,N_2467,N_2304);
xnor U2906 (N_2906,N_2216,N_2467);
xnor U2907 (N_2907,N_2161,N_2108);
nand U2908 (N_2908,N_2484,N_2251);
xor U2909 (N_2909,N_2257,N_2264);
xor U2910 (N_2910,N_2076,N_2237);
and U2911 (N_2911,N_2494,N_2384);
nor U2912 (N_2912,N_2192,N_2431);
or U2913 (N_2913,N_2418,N_2360);
and U2914 (N_2914,N_2305,N_2179);
nand U2915 (N_2915,N_2051,N_2275);
nand U2916 (N_2916,N_2235,N_2343);
nor U2917 (N_2917,N_2007,N_2326);
nand U2918 (N_2918,N_2363,N_2173);
nor U2919 (N_2919,N_2213,N_2218);
xnor U2920 (N_2920,N_2150,N_2455);
and U2921 (N_2921,N_2244,N_2254);
xor U2922 (N_2922,N_2083,N_2460);
and U2923 (N_2923,N_2120,N_2271);
or U2924 (N_2924,N_2323,N_2173);
and U2925 (N_2925,N_2310,N_2252);
xnor U2926 (N_2926,N_2271,N_2159);
nor U2927 (N_2927,N_2317,N_2237);
nor U2928 (N_2928,N_2251,N_2114);
or U2929 (N_2929,N_2000,N_2244);
and U2930 (N_2930,N_2011,N_2090);
or U2931 (N_2931,N_2047,N_2053);
nand U2932 (N_2932,N_2156,N_2019);
or U2933 (N_2933,N_2119,N_2206);
or U2934 (N_2934,N_2366,N_2208);
or U2935 (N_2935,N_2260,N_2098);
nand U2936 (N_2936,N_2473,N_2412);
or U2937 (N_2937,N_2490,N_2041);
xnor U2938 (N_2938,N_2103,N_2012);
nand U2939 (N_2939,N_2239,N_2428);
nor U2940 (N_2940,N_2336,N_2176);
nor U2941 (N_2941,N_2020,N_2252);
nand U2942 (N_2942,N_2221,N_2257);
or U2943 (N_2943,N_2215,N_2089);
nor U2944 (N_2944,N_2368,N_2164);
and U2945 (N_2945,N_2478,N_2499);
xnor U2946 (N_2946,N_2115,N_2048);
and U2947 (N_2947,N_2452,N_2144);
nor U2948 (N_2948,N_2073,N_2010);
nor U2949 (N_2949,N_2487,N_2194);
nand U2950 (N_2950,N_2085,N_2097);
nor U2951 (N_2951,N_2095,N_2302);
xnor U2952 (N_2952,N_2483,N_2050);
nand U2953 (N_2953,N_2135,N_2380);
nand U2954 (N_2954,N_2497,N_2080);
or U2955 (N_2955,N_2043,N_2026);
nor U2956 (N_2956,N_2444,N_2033);
nor U2957 (N_2957,N_2129,N_2238);
nor U2958 (N_2958,N_2388,N_2010);
and U2959 (N_2959,N_2497,N_2420);
nor U2960 (N_2960,N_2450,N_2163);
xnor U2961 (N_2961,N_2129,N_2073);
nand U2962 (N_2962,N_2025,N_2075);
xnor U2963 (N_2963,N_2461,N_2056);
nand U2964 (N_2964,N_2405,N_2027);
nand U2965 (N_2965,N_2153,N_2459);
or U2966 (N_2966,N_2031,N_2133);
xor U2967 (N_2967,N_2171,N_2476);
or U2968 (N_2968,N_2302,N_2111);
nor U2969 (N_2969,N_2450,N_2392);
xnor U2970 (N_2970,N_2062,N_2401);
and U2971 (N_2971,N_2217,N_2471);
or U2972 (N_2972,N_2428,N_2258);
nand U2973 (N_2973,N_2374,N_2480);
xnor U2974 (N_2974,N_2104,N_2324);
and U2975 (N_2975,N_2377,N_2345);
nand U2976 (N_2976,N_2153,N_2492);
nor U2977 (N_2977,N_2106,N_2349);
and U2978 (N_2978,N_2438,N_2426);
nor U2979 (N_2979,N_2089,N_2485);
or U2980 (N_2980,N_2220,N_2211);
and U2981 (N_2981,N_2191,N_2309);
xor U2982 (N_2982,N_2006,N_2424);
xor U2983 (N_2983,N_2016,N_2352);
and U2984 (N_2984,N_2124,N_2363);
xnor U2985 (N_2985,N_2423,N_2092);
nand U2986 (N_2986,N_2080,N_2402);
xnor U2987 (N_2987,N_2209,N_2376);
and U2988 (N_2988,N_2402,N_2336);
nor U2989 (N_2989,N_2389,N_2025);
or U2990 (N_2990,N_2383,N_2020);
or U2991 (N_2991,N_2458,N_2279);
nand U2992 (N_2992,N_2279,N_2193);
and U2993 (N_2993,N_2276,N_2000);
nand U2994 (N_2994,N_2425,N_2415);
xnor U2995 (N_2995,N_2447,N_2430);
and U2996 (N_2996,N_2490,N_2044);
or U2997 (N_2997,N_2122,N_2344);
and U2998 (N_2998,N_2247,N_2053);
nor U2999 (N_2999,N_2318,N_2413);
nand U3000 (N_3000,N_2757,N_2525);
or U3001 (N_3001,N_2676,N_2886);
nor U3002 (N_3002,N_2873,N_2510);
nand U3003 (N_3003,N_2897,N_2541);
xnor U3004 (N_3004,N_2611,N_2581);
or U3005 (N_3005,N_2723,N_2702);
nor U3006 (N_3006,N_2855,N_2693);
and U3007 (N_3007,N_2952,N_2907);
nand U3008 (N_3008,N_2904,N_2953);
and U3009 (N_3009,N_2574,N_2863);
xnor U3010 (N_3010,N_2815,N_2782);
or U3011 (N_3011,N_2878,N_2721);
nor U3012 (N_3012,N_2982,N_2725);
or U3013 (N_3013,N_2658,N_2846);
and U3014 (N_3014,N_2979,N_2613);
nand U3015 (N_3015,N_2887,N_2675);
and U3016 (N_3016,N_2832,N_2728);
or U3017 (N_3017,N_2546,N_2970);
nor U3018 (N_3018,N_2866,N_2512);
nand U3019 (N_3019,N_2517,N_2939);
nand U3020 (N_3020,N_2857,N_2647);
nand U3021 (N_3021,N_2714,N_2841);
xor U3022 (N_3022,N_2854,N_2708);
xor U3023 (N_3023,N_2890,N_2666);
and U3024 (N_3024,N_2930,N_2687);
nand U3025 (N_3025,N_2899,N_2936);
and U3026 (N_3026,N_2769,N_2942);
or U3027 (N_3027,N_2995,N_2627);
nand U3028 (N_3028,N_2969,N_2635);
or U3029 (N_3029,N_2505,N_2926);
xor U3030 (N_3030,N_2888,N_2813);
or U3031 (N_3031,N_2508,N_2909);
xor U3032 (N_3032,N_2922,N_2754);
and U3033 (N_3033,N_2961,N_2649);
xor U3034 (N_3034,N_2641,N_2677);
and U3035 (N_3035,N_2957,N_2506);
and U3036 (N_3036,N_2535,N_2994);
nor U3037 (N_3037,N_2664,N_2685);
and U3038 (N_3038,N_2597,N_2968);
and U3039 (N_3039,N_2673,N_2612);
or U3040 (N_3040,N_2801,N_2738);
nand U3041 (N_3041,N_2730,N_2698);
nor U3042 (N_3042,N_2674,N_2780);
xnor U3043 (N_3043,N_2739,N_2646);
or U3044 (N_3044,N_2615,N_2981);
xor U3045 (N_3045,N_2853,N_2575);
xnor U3046 (N_3046,N_2683,N_2774);
and U3047 (N_3047,N_2937,N_2915);
and U3048 (N_3048,N_2614,N_2903);
or U3049 (N_3049,N_2644,N_2671);
xnor U3050 (N_3050,N_2959,N_2560);
nand U3051 (N_3051,N_2773,N_2638);
nor U3052 (N_3052,N_2564,N_2565);
xnor U3053 (N_3053,N_2912,N_2734);
nor U3054 (N_3054,N_2862,N_2806);
nor U3055 (N_3055,N_2713,N_2880);
and U3056 (N_3056,N_2819,N_2562);
or U3057 (N_3057,N_2944,N_2534);
and U3058 (N_3058,N_2705,N_2760);
nor U3059 (N_3059,N_2843,N_2761);
or U3060 (N_3060,N_2971,N_2567);
xor U3061 (N_3061,N_2703,N_2632);
and U3062 (N_3062,N_2607,N_2593);
nand U3063 (N_3063,N_2511,N_2945);
xnor U3064 (N_3064,N_2619,N_2672);
xnor U3065 (N_3065,N_2771,N_2849);
or U3066 (N_3066,N_2605,N_2755);
or U3067 (N_3067,N_2602,N_2777);
nor U3068 (N_3068,N_2758,N_2503);
nand U3069 (N_3069,N_2720,N_2695);
or U3070 (N_3070,N_2539,N_2621);
or U3071 (N_3071,N_2587,N_2962);
nand U3072 (N_3072,N_2872,N_2733);
xor U3073 (N_3073,N_2793,N_2642);
and U3074 (N_3074,N_2543,N_2988);
nand U3075 (N_3075,N_2515,N_2583);
or U3076 (N_3076,N_2894,N_2618);
xor U3077 (N_3077,N_2827,N_2833);
xnor U3078 (N_3078,N_2844,N_2622);
or U3079 (N_3079,N_2706,N_2501);
nor U3080 (N_3080,N_2779,N_2584);
and U3081 (N_3081,N_2648,N_2839);
and U3082 (N_3082,N_2579,N_2967);
nand U3083 (N_3083,N_2920,N_2617);
and U3084 (N_3084,N_2528,N_2608);
and U3085 (N_3085,N_2811,N_2568);
nor U3086 (N_3086,N_2657,N_2544);
nand U3087 (N_3087,N_2984,N_2913);
nand U3088 (N_3088,N_2788,N_2704);
and U3089 (N_3089,N_2557,N_2818);
nor U3090 (N_3090,N_2616,N_2652);
nand U3091 (N_3091,N_2835,N_2921);
or U3092 (N_3092,N_2591,N_2719);
nor U3093 (N_3093,N_2781,N_2716);
or U3094 (N_3094,N_2751,N_2566);
nand U3095 (N_3095,N_2885,N_2941);
and U3096 (N_3096,N_2975,N_2711);
or U3097 (N_3097,N_2786,N_2765);
and U3098 (N_3098,N_2661,N_2830);
and U3099 (N_3099,N_2669,N_2917);
nand U3100 (N_3100,N_2545,N_2604);
and U3101 (N_3101,N_2650,N_2729);
nand U3102 (N_3102,N_2883,N_2928);
or U3103 (N_3103,N_2825,N_2812);
and U3104 (N_3104,N_2516,N_2927);
and U3105 (N_3105,N_2736,N_2665);
or U3106 (N_3106,N_2750,N_2529);
xor U3107 (N_3107,N_2869,N_2845);
nor U3108 (N_3108,N_2993,N_2791);
or U3109 (N_3109,N_2831,N_2859);
nand U3110 (N_3110,N_2836,N_2923);
xor U3111 (N_3111,N_2856,N_2877);
nand U3112 (N_3112,N_2550,N_2804);
nand U3113 (N_3113,N_2884,N_2670);
xnor U3114 (N_3114,N_2542,N_2767);
and U3115 (N_3115,N_2752,N_2824);
or U3116 (N_3116,N_2983,N_2724);
nand U3117 (N_3117,N_2933,N_2893);
nor U3118 (N_3118,N_2655,N_2585);
xor U3119 (N_3119,N_2906,N_2807);
nand U3120 (N_3120,N_2861,N_2924);
and U3121 (N_3121,N_2947,N_2745);
and U3122 (N_3122,N_2643,N_2896);
xor U3123 (N_3123,N_2532,N_2998);
nand U3124 (N_3124,N_2783,N_2530);
and U3125 (N_3125,N_2690,N_2840);
and U3126 (N_3126,N_2697,N_2524);
xnor U3127 (N_3127,N_2951,N_2996);
nand U3128 (N_3128,N_2964,N_2868);
and U3129 (N_3129,N_2680,N_2556);
xor U3130 (N_3130,N_2829,N_2834);
or U3131 (N_3131,N_2805,N_2606);
and U3132 (N_3132,N_2974,N_2620);
nor U3133 (N_3133,N_2925,N_2688);
nor U3134 (N_3134,N_2571,N_2908);
nand U3135 (N_3135,N_2744,N_2691);
and U3136 (N_3136,N_2547,N_2814);
nand U3137 (N_3137,N_2989,N_2940);
and U3138 (N_3138,N_2727,N_2537);
or U3139 (N_3139,N_2701,N_2992);
and U3140 (N_3140,N_2502,N_2795);
xor U3141 (N_3141,N_2717,N_2514);
or U3142 (N_3142,N_2710,N_2743);
and U3143 (N_3143,N_2624,N_2722);
xor U3144 (N_3144,N_2916,N_2526);
nand U3145 (N_3145,N_2558,N_2826);
nor U3146 (N_3146,N_2582,N_2796);
xnor U3147 (N_3147,N_2946,N_2759);
xnor U3148 (N_3148,N_2965,N_2763);
or U3149 (N_3149,N_2871,N_2985);
nand U3150 (N_3150,N_2838,N_2726);
and U3151 (N_3151,N_2694,N_2918);
and U3152 (N_3152,N_2640,N_2934);
xnor U3153 (N_3153,N_2577,N_2569);
xor U3154 (N_3154,N_2681,N_2609);
nand U3155 (N_3155,N_2707,N_2910);
nor U3156 (N_3156,N_2990,N_2768);
nor U3157 (N_3157,N_2552,N_2789);
and U3158 (N_3158,N_2513,N_2696);
and U3159 (N_3159,N_2519,N_2784);
and U3160 (N_3160,N_2938,N_2889);
or U3161 (N_3161,N_2610,N_2803);
and U3162 (N_3162,N_2628,N_2631);
or U3163 (N_3163,N_2551,N_2527);
or U3164 (N_3164,N_2850,N_2949);
nand U3165 (N_3165,N_2559,N_2799);
xnor U3166 (N_3166,N_2678,N_2553);
and U3167 (N_3167,N_2592,N_2660);
or U3168 (N_3168,N_2712,N_2598);
or U3169 (N_3169,N_2601,N_2794);
nor U3170 (N_3170,N_2504,N_2764);
and U3171 (N_3171,N_2740,N_2822);
or U3172 (N_3172,N_2997,N_2828);
or U3173 (N_3173,N_2816,N_2538);
or U3174 (N_3174,N_2842,N_2977);
nor U3175 (N_3175,N_2639,N_2742);
or U3176 (N_3176,N_2563,N_2810);
or U3177 (N_3177,N_2797,N_2684);
and U3178 (N_3178,N_2561,N_2715);
or U3179 (N_3179,N_2895,N_2860);
and U3180 (N_3180,N_2548,N_2963);
nand U3181 (N_3181,N_2523,N_2596);
xor U3182 (N_3182,N_2570,N_2870);
xnor U3183 (N_3183,N_2507,N_2902);
and U3184 (N_3184,N_2914,N_2645);
nor U3185 (N_3185,N_2932,N_2879);
or U3186 (N_3186,N_2580,N_2966);
nor U3187 (N_3187,N_2654,N_2931);
xor U3188 (N_3188,N_2600,N_2858);
or U3189 (N_3189,N_2973,N_2662);
nor U3190 (N_3190,N_2817,N_2785);
nand U3191 (N_3191,N_2876,N_2522);
and U3192 (N_3192,N_2533,N_2972);
and U3193 (N_3193,N_2802,N_2589);
and U3194 (N_3194,N_2625,N_2875);
or U3195 (N_3195,N_2978,N_2536);
and U3196 (N_3196,N_2540,N_2656);
nor U3197 (N_3197,N_2573,N_2958);
and U3198 (N_3198,N_2776,N_2986);
nor U3199 (N_3199,N_2748,N_2766);
xnor U3200 (N_3200,N_2595,N_2731);
or U3201 (N_3201,N_2770,N_2699);
nor U3202 (N_3202,N_2689,N_2554);
and U3203 (N_3203,N_2864,N_2955);
or U3204 (N_3204,N_2787,N_2900);
or U3205 (N_3205,N_2882,N_2800);
xor U3206 (N_3206,N_2999,N_2901);
nor U3207 (N_3207,N_2629,N_2746);
nor U3208 (N_3208,N_2603,N_2848);
nand U3209 (N_3209,N_2549,N_2772);
xor U3210 (N_3210,N_2741,N_2623);
nor U3211 (N_3211,N_2987,N_2663);
or U3212 (N_3212,N_2633,N_2637);
and U3213 (N_3213,N_2960,N_2756);
nand U3214 (N_3214,N_2892,N_2948);
and U3215 (N_3215,N_2737,N_2572);
or U3216 (N_3216,N_2775,N_2837);
nand U3217 (N_3217,N_2881,N_2500);
nor U3218 (N_3218,N_2653,N_2935);
or U3219 (N_3219,N_2679,N_2991);
nor U3220 (N_3220,N_2700,N_2747);
and U3221 (N_3221,N_2667,N_2576);
nand U3222 (N_3222,N_2905,N_2753);
nand U3223 (N_3223,N_2867,N_2792);
nor U3224 (N_3224,N_2865,N_2943);
and U3225 (N_3225,N_2821,N_2976);
and U3226 (N_3226,N_2852,N_2518);
nor U3227 (N_3227,N_2709,N_2509);
and U3228 (N_3228,N_2590,N_2578);
xor U3229 (N_3229,N_2682,N_2762);
nand U3230 (N_3230,N_2586,N_2718);
xor U3231 (N_3231,N_2521,N_2891);
and U3232 (N_3232,N_2630,N_2809);
or U3233 (N_3233,N_2520,N_2735);
and U3234 (N_3234,N_2599,N_2594);
xnor U3235 (N_3235,N_2626,N_2588);
or U3236 (N_3236,N_2531,N_2808);
nand U3237 (N_3237,N_2929,N_2634);
nor U3238 (N_3238,N_2898,N_2851);
and U3239 (N_3239,N_2798,N_2954);
and U3240 (N_3240,N_2980,N_2956);
or U3241 (N_3241,N_2749,N_2820);
and U3242 (N_3242,N_2692,N_2555);
nor U3243 (N_3243,N_2659,N_2911);
nor U3244 (N_3244,N_2668,N_2636);
or U3245 (N_3245,N_2732,N_2651);
nand U3246 (N_3246,N_2874,N_2778);
nand U3247 (N_3247,N_2790,N_2919);
xor U3248 (N_3248,N_2686,N_2950);
or U3249 (N_3249,N_2847,N_2823);
xnor U3250 (N_3250,N_2999,N_2907);
or U3251 (N_3251,N_2598,N_2638);
nor U3252 (N_3252,N_2617,N_2712);
nand U3253 (N_3253,N_2902,N_2506);
or U3254 (N_3254,N_2872,N_2836);
or U3255 (N_3255,N_2585,N_2740);
nor U3256 (N_3256,N_2556,N_2944);
xnor U3257 (N_3257,N_2778,N_2653);
xor U3258 (N_3258,N_2704,N_2562);
and U3259 (N_3259,N_2950,N_2562);
xor U3260 (N_3260,N_2638,N_2872);
nor U3261 (N_3261,N_2936,N_2998);
nand U3262 (N_3262,N_2730,N_2834);
nor U3263 (N_3263,N_2883,N_2952);
nand U3264 (N_3264,N_2696,N_2937);
or U3265 (N_3265,N_2814,N_2900);
nor U3266 (N_3266,N_2847,N_2957);
xnor U3267 (N_3267,N_2900,N_2558);
nand U3268 (N_3268,N_2522,N_2631);
xnor U3269 (N_3269,N_2565,N_2537);
and U3270 (N_3270,N_2558,N_2637);
nor U3271 (N_3271,N_2733,N_2945);
or U3272 (N_3272,N_2961,N_2855);
nor U3273 (N_3273,N_2926,N_2698);
nor U3274 (N_3274,N_2539,N_2739);
nor U3275 (N_3275,N_2838,N_2702);
xnor U3276 (N_3276,N_2973,N_2712);
nor U3277 (N_3277,N_2952,N_2713);
and U3278 (N_3278,N_2729,N_2596);
or U3279 (N_3279,N_2723,N_2961);
and U3280 (N_3280,N_2922,N_2942);
nor U3281 (N_3281,N_2946,N_2823);
or U3282 (N_3282,N_2661,N_2561);
xor U3283 (N_3283,N_2650,N_2728);
nor U3284 (N_3284,N_2980,N_2602);
or U3285 (N_3285,N_2953,N_2910);
xnor U3286 (N_3286,N_2854,N_2582);
or U3287 (N_3287,N_2948,N_2936);
nor U3288 (N_3288,N_2947,N_2558);
and U3289 (N_3289,N_2584,N_2849);
nor U3290 (N_3290,N_2713,N_2793);
or U3291 (N_3291,N_2791,N_2795);
xor U3292 (N_3292,N_2767,N_2624);
nor U3293 (N_3293,N_2882,N_2962);
or U3294 (N_3294,N_2864,N_2605);
or U3295 (N_3295,N_2691,N_2526);
and U3296 (N_3296,N_2909,N_2791);
nand U3297 (N_3297,N_2536,N_2784);
nand U3298 (N_3298,N_2688,N_2961);
and U3299 (N_3299,N_2879,N_2547);
nor U3300 (N_3300,N_2639,N_2907);
and U3301 (N_3301,N_2994,N_2898);
nor U3302 (N_3302,N_2600,N_2996);
xnor U3303 (N_3303,N_2982,N_2726);
and U3304 (N_3304,N_2694,N_2637);
xnor U3305 (N_3305,N_2970,N_2552);
nand U3306 (N_3306,N_2639,N_2892);
nand U3307 (N_3307,N_2876,N_2513);
and U3308 (N_3308,N_2841,N_2842);
nor U3309 (N_3309,N_2990,N_2975);
nand U3310 (N_3310,N_2870,N_2999);
and U3311 (N_3311,N_2808,N_2718);
and U3312 (N_3312,N_2844,N_2824);
or U3313 (N_3313,N_2978,N_2604);
and U3314 (N_3314,N_2780,N_2611);
nand U3315 (N_3315,N_2599,N_2917);
and U3316 (N_3316,N_2914,N_2746);
nand U3317 (N_3317,N_2752,N_2575);
xor U3318 (N_3318,N_2630,N_2943);
or U3319 (N_3319,N_2671,N_2802);
or U3320 (N_3320,N_2814,N_2887);
nand U3321 (N_3321,N_2647,N_2951);
nor U3322 (N_3322,N_2528,N_2572);
and U3323 (N_3323,N_2874,N_2987);
xor U3324 (N_3324,N_2982,N_2501);
nor U3325 (N_3325,N_2673,N_2911);
xor U3326 (N_3326,N_2528,N_2764);
nor U3327 (N_3327,N_2929,N_2759);
and U3328 (N_3328,N_2840,N_2984);
nand U3329 (N_3329,N_2507,N_2839);
xor U3330 (N_3330,N_2671,N_2876);
nand U3331 (N_3331,N_2500,N_2816);
nor U3332 (N_3332,N_2515,N_2838);
or U3333 (N_3333,N_2506,N_2898);
nor U3334 (N_3334,N_2903,N_2738);
and U3335 (N_3335,N_2882,N_2749);
or U3336 (N_3336,N_2884,N_2530);
xnor U3337 (N_3337,N_2733,N_2692);
nor U3338 (N_3338,N_2631,N_2919);
nand U3339 (N_3339,N_2823,N_2978);
xor U3340 (N_3340,N_2849,N_2563);
xnor U3341 (N_3341,N_2557,N_2651);
and U3342 (N_3342,N_2622,N_2826);
nor U3343 (N_3343,N_2896,N_2654);
or U3344 (N_3344,N_2903,N_2833);
xor U3345 (N_3345,N_2864,N_2896);
nor U3346 (N_3346,N_2946,N_2518);
or U3347 (N_3347,N_2963,N_2873);
nor U3348 (N_3348,N_2659,N_2816);
nand U3349 (N_3349,N_2818,N_2512);
xnor U3350 (N_3350,N_2560,N_2666);
nand U3351 (N_3351,N_2832,N_2504);
or U3352 (N_3352,N_2706,N_2618);
and U3353 (N_3353,N_2777,N_2771);
or U3354 (N_3354,N_2848,N_2704);
xnor U3355 (N_3355,N_2591,N_2869);
and U3356 (N_3356,N_2748,N_2896);
nand U3357 (N_3357,N_2549,N_2559);
xor U3358 (N_3358,N_2692,N_2790);
nand U3359 (N_3359,N_2890,N_2795);
xor U3360 (N_3360,N_2572,N_2859);
and U3361 (N_3361,N_2559,N_2548);
nor U3362 (N_3362,N_2714,N_2621);
or U3363 (N_3363,N_2726,N_2677);
or U3364 (N_3364,N_2885,N_2520);
nand U3365 (N_3365,N_2593,N_2689);
or U3366 (N_3366,N_2615,N_2590);
or U3367 (N_3367,N_2630,N_2835);
nand U3368 (N_3368,N_2724,N_2933);
xor U3369 (N_3369,N_2712,N_2895);
or U3370 (N_3370,N_2885,N_2759);
and U3371 (N_3371,N_2530,N_2613);
and U3372 (N_3372,N_2602,N_2620);
nand U3373 (N_3373,N_2630,N_2612);
or U3374 (N_3374,N_2690,N_2882);
nand U3375 (N_3375,N_2722,N_2651);
nand U3376 (N_3376,N_2501,N_2692);
xor U3377 (N_3377,N_2572,N_2700);
nand U3378 (N_3378,N_2988,N_2907);
and U3379 (N_3379,N_2852,N_2976);
nand U3380 (N_3380,N_2777,N_2915);
or U3381 (N_3381,N_2543,N_2758);
or U3382 (N_3382,N_2651,N_2947);
or U3383 (N_3383,N_2865,N_2560);
nand U3384 (N_3384,N_2769,N_2653);
or U3385 (N_3385,N_2952,N_2640);
and U3386 (N_3386,N_2532,N_2639);
xnor U3387 (N_3387,N_2900,N_2908);
xnor U3388 (N_3388,N_2848,N_2998);
nor U3389 (N_3389,N_2552,N_2522);
or U3390 (N_3390,N_2970,N_2934);
or U3391 (N_3391,N_2534,N_2670);
or U3392 (N_3392,N_2628,N_2970);
xnor U3393 (N_3393,N_2929,N_2630);
or U3394 (N_3394,N_2547,N_2538);
nand U3395 (N_3395,N_2645,N_2809);
nand U3396 (N_3396,N_2583,N_2905);
xor U3397 (N_3397,N_2541,N_2973);
nor U3398 (N_3398,N_2981,N_2969);
or U3399 (N_3399,N_2814,N_2751);
and U3400 (N_3400,N_2517,N_2886);
and U3401 (N_3401,N_2871,N_2968);
or U3402 (N_3402,N_2976,N_2638);
xnor U3403 (N_3403,N_2883,N_2644);
nand U3404 (N_3404,N_2611,N_2615);
nor U3405 (N_3405,N_2844,N_2889);
nor U3406 (N_3406,N_2514,N_2726);
nor U3407 (N_3407,N_2634,N_2611);
nand U3408 (N_3408,N_2515,N_2976);
nand U3409 (N_3409,N_2510,N_2614);
xnor U3410 (N_3410,N_2549,N_2824);
and U3411 (N_3411,N_2845,N_2951);
nor U3412 (N_3412,N_2854,N_2888);
xnor U3413 (N_3413,N_2688,N_2623);
nand U3414 (N_3414,N_2530,N_2573);
or U3415 (N_3415,N_2838,N_2594);
and U3416 (N_3416,N_2762,N_2969);
or U3417 (N_3417,N_2766,N_2831);
or U3418 (N_3418,N_2838,N_2853);
or U3419 (N_3419,N_2820,N_2661);
or U3420 (N_3420,N_2508,N_2956);
nand U3421 (N_3421,N_2755,N_2819);
or U3422 (N_3422,N_2563,N_2959);
xor U3423 (N_3423,N_2661,N_2889);
and U3424 (N_3424,N_2808,N_2702);
nor U3425 (N_3425,N_2952,N_2597);
or U3426 (N_3426,N_2618,N_2846);
xor U3427 (N_3427,N_2884,N_2725);
and U3428 (N_3428,N_2758,N_2547);
nor U3429 (N_3429,N_2724,N_2526);
or U3430 (N_3430,N_2582,N_2552);
and U3431 (N_3431,N_2604,N_2655);
nand U3432 (N_3432,N_2827,N_2957);
and U3433 (N_3433,N_2654,N_2787);
and U3434 (N_3434,N_2823,N_2884);
nor U3435 (N_3435,N_2809,N_2848);
nand U3436 (N_3436,N_2670,N_2698);
nor U3437 (N_3437,N_2658,N_2563);
nor U3438 (N_3438,N_2979,N_2621);
or U3439 (N_3439,N_2707,N_2606);
and U3440 (N_3440,N_2529,N_2617);
xnor U3441 (N_3441,N_2628,N_2808);
nand U3442 (N_3442,N_2729,N_2613);
nand U3443 (N_3443,N_2575,N_2874);
xor U3444 (N_3444,N_2884,N_2761);
or U3445 (N_3445,N_2616,N_2950);
nand U3446 (N_3446,N_2946,N_2561);
nand U3447 (N_3447,N_2977,N_2778);
xnor U3448 (N_3448,N_2926,N_2557);
or U3449 (N_3449,N_2958,N_2792);
nand U3450 (N_3450,N_2801,N_2516);
nand U3451 (N_3451,N_2892,N_2786);
or U3452 (N_3452,N_2670,N_2806);
or U3453 (N_3453,N_2618,N_2780);
xor U3454 (N_3454,N_2631,N_2863);
nor U3455 (N_3455,N_2947,N_2916);
or U3456 (N_3456,N_2739,N_2574);
nand U3457 (N_3457,N_2720,N_2986);
xnor U3458 (N_3458,N_2978,N_2511);
or U3459 (N_3459,N_2976,N_2740);
or U3460 (N_3460,N_2704,N_2720);
or U3461 (N_3461,N_2522,N_2513);
nor U3462 (N_3462,N_2653,N_2945);
and U3463 (N_3463,N_2984,N_2936);
or U3464 (N_3464,N_2675,N_2796);
xor U3465 (N_3465,N_2743,N_2611);
or U3466 (N_3466,N_2660,N_2957);
and U3467 (N_3467,N_2749,N_2878);
or U3468 (N_3468,N_2848,N_2503);
xor U3469 (N_3469,N_2628,N_2725);
xor U3470 (N_3470,N_2818,N_2555);
nand U3471 (N_3471,N_2863,N_2722);
xnor U3472 (N_3472,N_2651,N_2582);
xnor U3473 (N_3473,N_2592,N_2852);
nand U3474 (N_3474,N_2575,N_2633);
xor U3475 (N_3475,N_2870,N_2691);
nor U3476 (N_3476,N_2873,N_2810);
nor U3477 (N_3477,N_2956,N_2948);
or U3478 (N_3478,N_2895,N_2988);
or U3479 (N_3479,N_2713,N_2972);
and U3480 (N_3480,N_2640,N_2759);
nand U3481 (N_3481,N_2584,N_2681);
nor U3482 (N_3482,N_2797,N_2695);
xor U3483 (N_3483,N_2716,N_2738);
nand U3484 (N_3484,N_2925,N_2666);
nand U3485 (N_3485,N_2559,N_2668);
or U3486 (N_3486,N_2889,N_2568);
and U3487 (N_3487,N_2628,N_2925);
or U3488 (N_3488,N_2974,N_2852);
nor U3489 (N_3489,N_2718,N_2769);
nor U3490 (N_3490,N_2883,N_2873);
nand U3491 (N_3491,N_2915,N_2813);
xor U3492 (N_3492,N_2884,N_2520);
nor U3493 (N_3493,N_2814,N_2697);
nor U3494 (N_3494,N_2563,N_2727);
xnor U3495 (N_3495,N_2814,N_2594);
nor U3496 (N_3496,N_2809,N_2871);
xor U3497 (N_3497,N_2941,N_2834);
or U3498 (N_3498,N_2524,N_2705);
xor U3499 (N_3499,N_2656,N_2560);
nand U3500 (N_3500,N_3251,N_3268);
and U3501 (N_3501,N_3063,N_3495);
and U3502 (N_3502,N_3307,N_3175);
or U3503 (N_3503,N_3472,N_3096);
xnor U3504 (N_3504,N_3166,N_3302);
nor U3505 (N_3505,N_3320,N_3270);
and U3506 (N_3506,N_3039,N_3443);
nor U3507 (N_3507,N_3120,N_3119);
and U3508 (N_3508,N_3460,N_3256);
nand U3509 (N_3509,N_3373,N_3296);
nand U3510 (N_3510,N_3125,N_3317);
xor U3511 (N_3511,N_3454,N_3093);
nand U3512 (N_3512,N_3441,N_3115);
nor U3513 (N_3513,N_3364,N_3319);
nand U3514 (N_3514,N_3086,N_3479);
nor U3515 (N_3515,N_3076,N_3034);
and U3516 (N_3516,N_3337,N_3062);
or U3517 (N_3517,N_3217,N_3171);
and U3518 (N_3518,N_3067,N_3097);
or U3519 (N_3519,N_3385,N_3211);
nand U3520 (N_3520,N_3196,N_3069);
or U3521 (N_3521,N_3066,N_3312);
nor U3522 (N_3522,N_3057,N_3498);
nand U3523 (N_3523,N_3085,N_3417);
and U3524 (N_3524,N_3293,N_3485);
nand U3525 (N_3525,N_3017,N_3071);
xnor U3526 (N_3526,N_3471,N_3224);
nor U3527 (N_3527,N_3225,N_3470);
or U3528 (N_3528,N_3316,N_3028);
nand U3529 (N_3529,N_3304,N_3160);
nand U3530 (N_3530,N_3235,N_3450);
nor U3531 (N_3531,N_3026,N_3099);
nand U3532 (N_3532,N_3018,N_3311);
nor U3533 (N_3533,N_3082,N_3052);
or U3534 (N_3534,N_3003,N_3007);
or U3535 (N_3535,N_3214,N_3167);
nor U3536 (N_3536,N_3269,N_3006);
and U3537 (N_3537,N_3328,N_3223);
nor U3538 (N_3538,N_3178,N_3087);
nor U3539 (N_3539,N_3045,N_3486);
xor U3540 (N_3540,N_3453,N_3103);
xnor U3541 (N_3541,N_3210,N_3291);
nor U3542 (N_3542,N_3469,N_3324);
nand U3543 (N_3543,N_3098,N_3239);
nor U3544 (N_3544,N_3174,N_3027);
or U3545 (N_3545,N_3231,N_3040);
nand U3546 (N_3546,N_3413,N_3083);
nand U3547 (N_3547,N_3163,N_3226);
or U3548 (N_3548,N_3355,N_3480);
nor U3549 (N_3549,N_3091,N_3016);
xor U3550 (N_3550,N_3019,N_3109);
or U3551 (N_3551,N_3271,N_3393);
nor U3552 (N_3552,N_3464,N_3213);
nor U3553 (N_3553,N_3327,N_3154);
nand U3554 (N_3554,N_3147,N_3287);
or U3555 (N_3555,N_3146,N_3064);
or U3556 (N_3556,N_3369,N_3134);
nor U3557 (N_3557,N_3037,N_3241);
or U3558 (N_3558,N_3477,N_3061);
or U3559 (N_3559,N_3199,N_3387);
nand U3560 (N_3560,N_3331,N_3212);
and U3561 (N_3561,N_3117,N_3168);
and U3562 (N_3562,N_3436,N_3132);
and U3563 (N_3563,N_3234,N_3151);
nand U3564 (N_3564,N_3145,N_3247);
nand U3565 (N_3565,N_3029,N_3333);
nor U3566 (N_3566,N_3164,N_3329);
nor U3567 (N_3567,N_3463,N_3411);
or U3568 (N_3568,N_3424,N_3130);
and U3569 (N_3569,N_3438,N_3338);
or U3570 (N_3570,N_3159,N_3065);
or U3571 (N_3571,N_3068,N_3105);
nand U3572 (N_3572,N_3140,N_3280);
and U3573 (N_3573,N_3216,N_3418);
and U3574 (N_3574,N_3092,N_3023);
xor U3575 (N_3575,N_3056,N_3272);
xnor U3576 (N_3576,N_3165,N_3158);
nand U3577 (N_3577,N_3194,N_3466);
xnor U3578 (N_3578,N_3395,N_3289);
and U3579 (N_3579,N_3310,N_3288);
xor U3580 (N_3580,N_3403,N_3357);
or U3581 (N_3581,N_3202,N_3384);
nor U3582 (N_3582,N_3397,N_3415);
nand U3583 (N_3583,N_3108,N_3070);
and U3584 (N_3584,N_3243,N_3010);
and U3585 (N_3585,N_3113,N_3255);
xor U3586 (N_3586,N_3394,N_3104);
nand U3587 (N_3587,N_3363,N_3282);
nand U3588 (N_3588,N_3425,N_3264);
nand U3589 (N_3589,N_3490,N_3123);
xnor U3590 (N_3590,N_3434,N_3177);
and U3591 (N_3591,N_3204,N_3346);
nand U3592 (N_3592,N_3230,N_3187);
and U3593 (N_3593,N_3491,N_3195);
or U3594 (N_3594,N_3143,N_3433);
xnor U3595 (N_3595,N_3439,N_3349);
xor U3596 (N_3596,N_3467,N_3347);
or U3597 (N_3597,N_3025,N_3376);
nor U3598 (N_3598,N_3414,N_3379);
nand U3599 (N_3599,N_3430,N_3481);
or U3600 (N_3600,N_3131,N_3127);
or U3601 (N_3601,N_3218,N_3049);
nand U3602 (N_3602,N_3351,N_3248);
nor U3603 (N_3603,N_3401,N_3493);
nor U3604 (N_3604,N_3257,N_3074);
xor U3605 (N_3605,N_3284,N_3445);
or U3606 (N_3606,N_3261,N_3184);
nand U3607 (N_3607,N_3406,N_3020);
nand U3608 (N_3608,N_3487,N_3170);
nor U3609 (N_3609,N_3221,N_3118);
nor U3610 (N_3610,N_3378,N_3303);
nor U3611 (N_3611,N_3153,N_3227);
or U3612 (N_3612,N_3262,N_3400);
or U3613 (N_3613,N_3141,N_3353);
or U3614 (N_3614,N_3295,N_3030);
nand U3615 (N_3615,N_3201,N_3238);
nor U3616 (N_3616,N_3339,N_3032);
xnor U3617 (N_3617,N_3455,N_3399);
and U3618 (N_3618,N_3022,N_3013);
or U3619 (N_3619,N_3048,N_3465);
and U3620 (N_3620,N_3047,N_3371);
or U3621 (N_3621,N_3322,N_3172);
nand U3622 (N_3622,N_3191,N_3391);
xnor U3623 (N_3623,N_3468,N_3309);
nand U3624 (N_3624,N_3451,N_3294);
and U3625 (N_3625,N_3366,N_3308);
and U3626 (N_3626,N_3041,N_3267);
xor U3627 (N_3627,N_3046,N_3169);
and U3628 (N_3628,N_3354,N_3220);
nor U3629 (N_3629,N_3273,N_3207);
or U3630 (N_3630,N_3419,N_3051);
nor U3631 (N_3631,N_3276,N_3180);
and U3632 (N_3632,N_3244,N_3054);
or U3633 (N_3633,N_3240,N_3462);
or U3634 (N_3634,N_3279,N_3435);
nor U3635 (N_3635,N_3050,N_3429);
nor U3636 (N_3636,N_3407,N_3292);
or U3637 (N_3637,N_3375,N_3044);
xor U3638 (N_3638,N_3405,N_3242);
xnor U3639 (N_3639,N_3356,N_3094);
nor U3640 (N_3640,N_3233,N_3330);
or U3641 (N_3641,N_3281,N_3428);
or U3642 (N_3642,N_3176,N_3388);
or U3643 (N_3643,N_3232,N_3249);
nand U3644 (N_3644,N_3344,N_3422);
xor U3645 (N_3645,N_3015,N_3404);
xnor U3646 (N_3646,N_3313,N_3408);
and U3647 (N_3647,N_3409,N_3260);
nand U3648 (N_3648,N_3421,N_3381);
and U3649 (N_3649,N_3183,N_3494);
xor U3650 (N_3650,N_3053,N_3205);
nand U3651 (N_3651,N_3423,N_3090);
or U3652 (N_3652,N_3265,N_3458);
xor U3653 (N_3653,N_3142,N_3150);
nand U3654 (N_3654,N_3081,N_3285);
nand U3655 (N_3655,N_3410,N_3473);
and U3656 (N_3656,N_3138,N_3186);
or U3657 (N_3657,N_3139,N_3386);
xor U3658 (N_3658,N_3058,N_3155);
or U3659 (N_3659,N_3124,N_3340);
or U3660 (N_3660,N_3301,N_3197);
xor U3661 (N_3661,N_3254,N_3345);
and U3662 (N_3662,N_3014,N_3444);
xnor U3663 (N_3663,N_3343,N_3283);
or U3664 (N_3664,N_3483,N_3002);
or U3665 (N_3665,N_3496,N_3215);
xnor U3666 (N_3666,N_3420,N_3365);
nand U3667 (N_3667,N_3121,N_3318);
and U3668 (N_3668,N_3306,N_3219);
and U3669 (N_3669,N_3358,N_3325);
xnor U3670 (N_3670,N_3489,N_3442);
nor U3671 (N_3671,N_3478,N_3208);
and U3672 (N_3672,N_3203,N_3278);
and U3673 (N_3673,N_3149,N_3334);
and U3674 (N_3674,N_3072,N_3352);
nand U3675 (N_3675,N_3416,N_3372);
nor U3676 (N_3676,N_3080,N_3370);
xor U3677 (N_3677,N_3259,N_3290);
nand U3678 (N_3678,N_3274,N_3059);
or U3679 (N_3679,N_3484,N_3396);
nand U3680 (N_3680,N_3088,N_3389);
nor U3681 (N_3681,N_3024,N_3055);
xor U3682 (N_3682,N_3456,N_3374);
nand U3683 (N_3683,N_3009,N_3162);
nor U3684 (N_3684,N_3367,N_3275);
xor U3685 (N_3685,N_3107,N_3122);
nor U3686 (N_3686,N_3152,N_3432);
nand U3687 (N_3687,N_3110,N_3181);
nand U3688 (N_3688,N_3136,N_3437);
nand U3689 (N_3689,N_3206,N_3342);
or U3690 (N_3690,N_3001,N_3263);
or U3691 (N_3691,N_3449,N_3488);
or U3692 (N_3692,N_3380,N_3360);
nand U3693 (N_3693,N_3193,N_3156);
nand U3694 (N_3694,N_3392,N_3229);
xor U3695 (N_3695,N_3298,N_3390);
xor U3696 (N_3696,N_3012,N_3335);
nor U3697 (N_3697,N_3446,N_3135);
or U3698 (N_3698,N_3297,N_3236);
nor U3699 (N_3699,N_3315,N_3431);
xnor U3700 (N_3700,N_3075,N_3101);
xnor U3701 (N_3701,N_3475,N_3161);
or U3702 (N_3702,N_3448,N_3209);
and U3703 (N_3703,N_3157,N_3021);
and U3704 (N_3704,N_3084,N_3137);
or U3705 (N_3705,N_3192,N_3182);
or U3706 (N_3706,N_3336,N_3499);
nand U3707 (N_3707,N_3476,N_3106);
xnor U3708 (N_3708,N_3368,N_3077);
and U3709 (N_3709,N_3185,N_3043);
xor U3710 (N_3710,N_3073,N_3008);
and U3711 (N_3711,N_3078,N_3111);
or U3712 (N_3712,N_3129,N_3079);
and U3713 (N_3713,N_3250,N_3482);
xor U3714 (N_3714,N_3200,N_3038);
nor U3715 (N_3715,N_3126,N_3412);
nand U3716 (N_3716,N_3042,N_3398);
and U3717 (N_3717,N_3252,N_3228);
or U3718 (N_3718,N_3457,N_3299);
or U3719 (N_3719,N_3492,N_3100);
nand U3720 (N_3720,N_3361,N_3440);
and U3721 (N_3721,N_3332,N_3095);
and U3722 (N_3722,N_3321,N_3362);
nor U3723 (N_3723,N_3102,N_3173);
nand U3724 (N_3724,N_3326,N_3033);
nand U3725 (N_3725,N_3253,N_3112);
or U3726 (N_3726,N_3350,N_3246);
xor U3727 (N_3727,N_3427,N_3277);
xnor U3728 (N_3728,N_3305,N_3198);
and U3729 (N_3729,N_3133,N_3089);
nor U3730 (N_3730,N_3148,N_3245);
and U3731 (N_3731,N_3036,N_3114);
nor U3732 (N_3732,N_3461,N_3383);
and U3733 (N_3733,N_3179,N_3258);
xor U3734 (N_3734,N_3035,N_3323);
or U3735 (N_3735,N_3426,N_3348);
xnor U3736 (N_3736,N_3314,N_3286);
nor U3737 (N_3737,N_3459,N_3266);
or U3738 (N_3738,N_3000,N_3447);
nor U3739 (N_3739,N_3031,N_3190);
and U3740 (N_3740,N_3004,N_3452);
nand U3741 (N_3741,N_3382,N_3116);
nor U3742 (N_3742,N_3237,N_3359);
nand U3743 (N_3743,N_3189,N_3144);
xor U3744 (N_3744,N_3011,N_3222);
nand U3745 (N_3745,N_3060,N_3128);
nand U3746 (N_3746,N_3474,N_3402);
and U3747 (N_3747,N_3377,N_3188);
nor U3748 (N_3748,N_3300,N_3005);
xnor U3749 (N_3749,N_3341,N_3497);
nor U3750 (N_3750,N_3426,N_3393);
xor U3751 (N_3751,N_3092,N_3411);
xnor U3752 (N_3752,N_3448,N_3056);
xor U3753 (N_3753,N_3213,N_3043);
nand U3754 (N_3754,N_3174,N_3146);
and U3755 (N_3755,N_3448,N_3112);
nand U3756 (N_3756,N_3074,N_3146);
or U3757 (N_3757,N_3438,N_3172);
or U3758 (N_3758,N_3393,N_3242);
and U3759 (N_3759,N_3054,N_3439);
and U3760 (N_3760,N_3386,N_3247);
or U3761 (N_3761,N_3295,N_3288);
nor U3762 (N_3762,N_3394,N_3107);
xnor U3763 (N_3763,N_3103,N_3403);
xnor U3764 (N_3764,N_3400,N_3228);
or U3765 (N_3765,N_3063,N_3067);
nand U3766 (N_3766,N_3406,N_3271);
nor U3767 (N_3767,N_3484,N_3277);
and U3768 (N_3768,N_3472,N_3109);
or U3769 (N_3769,N_3027,N_3162);
nand U3770 (N_3770,N_3196,N_3089);
or U3771 (N_3771,N_3457,N_3012);
nor U3772 (N_3772,N_3399,N_3099);
or U3773 (N_3773,N_3425,N_3024);
and U3774 (N_3774,N_3456,N_3251);
xor U3775 (N_3775,N_3490,N_3027);
and U3776 (N_3776,N_3311,N_3057);
nand U3777 (N_3777,N_3184,N_3166);
nor U3778 (N_3778,N_3115,N_3036);
nand U3779 (N_3779,N_3229,N_3283);
or U3780 (N_3780,N_3498,N_3407);
nor U3781 (N_3781,N_3182,N_3201);
nand U3782 (N_3782,N_3374,N_3489);
and U3783 (N_3783,N_3411,N_3397);
and U3784 (N_3784,N_3242,N_3046);
nand U3785 (N_3785,N_3372,N_3022);
nand U3786 (N_3786,N_3041,N_3045);
nand U3787 (N_3787,N_3290,N_3269);
xor U3788 (N_3788,N_3127,N_3279);
nand U3789 (N_3789,N_3193,N_3294);
and U3790 (N_3790,N_3359,N_3268);
or U3791 (N_3791,N_3358,N_3266);
or U3792 (N_3792,N_3216,N_3255);
nor U3793 (N_3793,N_3213,N_3354);
nor U3794 (N_3794,N_3251,N_3212);
nor U3795 (N_3795,N_3017,N_3101);
and U3796 (N_3796,N_3488,N_3427);
xnor U3797 (N_3797,N_3370,N_3236);
and U3798 (N_3798,N_3034,N_3094);
and U3799 (N_3799,N_3481,N_3282);
or U3800 (N_3800,N_3029,N_3265);
or U3801 (N_3801,N_3083,N_3386);
xnor U3802 (N_3802,N_3402,N_3089);
nand U3803 (N_3803,N_3173,N_3279);
or U3804 (N_3804,N_3199,N_3016);
or U3805 (N_3805,N_3329,N_3076);
xnor U3806 (N_3806,N_3197,N_3465);
nand U3807 (N_3807,N_3376,N_3265);
and U3808 (N_3808,N_3125,N_3450);
nand U3809 (N_3809,N_3221,N_3352);
and U3810 (N_3810,N_3015,N_3073);
xor U3811 (N_3811,N_3422,N_3119);
nor U3812 (N_3812,N_3423,N_3022);
nand U3813 (N_3813,N_3263,N_3055);
nor U3814 (N_3814,N_3151,N_3474);
and U3815 (N_3815,N_3219,N_3439);
and U3816 (N_3816,N_3254,N_3264);
xnor U3817 (N_3817,N_3011,N_3112);
or U3818 (N_3818,N_3223,N_3372);
nor U3819 (N_3819,N_3211,N_3274);
nor U3820 (N_3820,N_3446,N_3094);
xor U3821 (N_3821,N_3135,N_3322);
xnor U3822 (N_3822,N_3359,N_3090);
and U3823 (N_3823,N_3366,N_3382);
or U3824 (N_3824,N_3452,N_3027);
xnor U3825 (N_3825,N_3338,N_3394);
xor U3826 (N_3826,N_3058,N_3447);
and U3827 (N_3827,N_3078,N_3310);
nand U3828 (N_3828,N_3023,N_3051);
nor U3829 (N_3829,N_3435,N_3142);
nand U3830 (N_3830,N_3299,N_3041);
nor U3831 (N_3831,N_3499,N_3400);
nand U3832 (N_3832,N_3188,N_3053);
xor U3833 (N_3833,N_3002,N_3123);
and U3834 (N_3834,N_3247,N_3073);
and U3835 (N_3835,N_3054,N_3117);
and U3836 (N_3836,N_3004,N_3072);
xor U3837 (N_3837,N_3017,N_3326);
nor U3838 (N_3838,N_3276,N_3067);
nor U3839 (N_3839,N_3320,N_3395);
xnor U3840 (N_3840,N_3080,N_3248);
nor U3841 (N_3841,N_3272,N_3498);
or U3842 (N_3842,N_3495,N_3129);
and U3843 (N_3843,N_3007,N_3078);
nand U3844 (N_3844,N_3013,N_3036);
nand U3845 (N_3845,N_3365,N_3338);
nor U3846 (N_3846,N_3460,N_3109);
or U3847 (N_3847,N_3362,N_3238);
nand U3848 (N_3848,N_3135,N_3130);
or U3849 (N_3849,N_3292,N_3061);
nor U3850 (N_3850,N_3112,N_3348);
xor U3851 (N_3851,N_3188,N_3477);
and U3852 (N_3852,N_3218,N_3093);
nand U3853 (N_3853,N_3009,N_3170);
nand U3854 (N_3854,N_3394,N_3123);
nor U3855 (N_3855,N_3106,N_3421);
nor U3856 (N_3856,N_3123,N_3214);
or U3857 (N_3857,N_3291,N_3494);
xor U3858 (N_3858,N_3340,N_3293);
xor U3859 (N_3859,N_3024,N_3040);
or U3860 (N_3860,N_3265,N_3417);
xor U3861 (N_3861,N_3034,N_3153);
nor U3862 (N_3862,N_3277,N_3211);
and U3863 (N_3863,N_3305,N_3210);
xor U3864 (N_3864,N_3091,N_3078);
nor U3865 (N_3865,N_3203,N_3491);
and U3866 (N_3866,N_3199,N_3428);
nor U3867 (N_3867,N_3365,N_3005);
nor U3868 (N_3868,N_3413,N_3075);
nor U3869 (N_3869,N_3053,N_3206);
nand U3870 (N_3870,N_3116,N_3430);
and U3871 (N_3871,N_3477,N_3304);
or U3872 (N_3872,N_3311,N_3383);
and U3873 (N_3873,N_3258,N_3137);
nand U3874 (N_3874,N_3102,N_3270);
and U3875 (N_3875,N_3338,N_3481);
nand U3876 (N_3876,N_3376,N_3241);
nor U3877 (N_3877,N_3128,N_3206);
nor U3878 (N_3878,N_3396,N_3063);
nor U3879 (N_3879,N_3139,N_3010);
nor U3880 (N_3880,N_3248,N_3340);
nand U3881 (N_3881,N_3192,N_3259);
and U3882 (N_3882,N_3386,N_3192);
nor U3883 (N_3883,N_3278,N_3363);
xnor U3884 (N_3884,N_3263,N_3317);
nand U3885 (N_3885,N_3084,N_3493);
nor U3886 (N_3886,N_3059,N_3257);
and U3887 (N_3887,N_3207,N_3233);
or U3888 (N_3888,N_3066,N_3299);
or U3889 (N_3889,N_3483,N_3170);
xnor U3890 (N_3890,N_3141,N_3036);
nand U3891 (N_3891,N_3490,N_3452);
and U3892 (N_3892,N_3002,N_3277);
and U3893 (N_3893,N_3067,N_3440);
nor U3894 (N_3894,N_3114,N_3366);
nor U3895 (N_3895,N_3436,N_3345);
nor U3896 (N_3896,N_3054,N_3289);
nand U3897 (N_3897,N_3208,N_3376);
nor U3898 (N_3898,N_3082,N_3274);
xor U3899 (N_3899,N_3106,N_3403);
and U3900 (N_3900,N_3293,N_3093);
and U3901 (N_3901,N_3222,N_3089);
xor U3902 (N_3902,N_3008,N_3158);
or U3903 (N_3903,N_3419,N_3018);
nand U3904 (N_3904,N_3445,N_3157);
and U3905 (N_3905,N_3084,N_3291);
and U3906 (N_3906,N_3158,N_3412);
nor U3907 (N_3907,N_3467,N_3468);
nor U3908 (N_3908,N_3285,N_3382);
xor U3909 (N_3909,N_3393,N_3376);
and U3910 (N_3910,N_3132,N_3383);
nand U3911 (N_3911,N_3253,N_3179);
or U3912 (N_3912,N_3146,N_3057);
or U3913 (N_3913,N_3190,N_3345);
xor U3914 (N_3914,N_3042,N_3284);
nor U3915 (N_3915,N_3071,N_3447);
nand U3916 (N_3916,N_3309,N_3332);
or U3917 (N_3917,N_3365,N_3437);
nand U3918 (N_3918,N_3403,N_3359);
xnor U3919 (N_3919,N_3103,N_3199);
and U3920 (N_3920,N_3020,N_3157);
nor U3921 (N_3921,N_3324,N_3418);
xor U3922 (N_3922,N_3337,N_3316);
or U3923 (N_3923,N_3294,N_3322);
xor U3924 (N_3924,N_3408,N_3075);
and U3925 (N_3925,N_3276,N_3374);
xor U3926 (N_3926,N_3495,N_3090);
nor U3927 (N_3927,N_3317,N_3337);
nand U3928 (N_3928,N_3202,N_3167);
or U3929 (N_3929,N_3385,N_3439);
nand U3930 (N_3930,N_3469,N_3398);
nor U3931 (N_3931,N_3276,N_3167);
and U3932 (N_3932,N_3277,N_3477);
nand U3933 (N_3933,N_3331,N_3451);
nor U3934 (N_3934,N_3373,N_3490);
or U3935 (N_3935,N_3014,N_3169);
xor U3936 (N_3936,N_3427,N_3208);
nand U3937 (N_3937,N_3310,N_3447);
or U3938 (N_3938,N_3304,N_3343);
nand U3939 (N_3939,N_3370,N_3144);
xor U3940 (N_3940,N_3060,N_3075);
nor U3941 (N_3941,N_3272,N_3182);
xor U3942 (N_3942,N_3062,N_3077);
xnor U3943 (N_3943,N_3072,N_3367);
nor U3944 (N_3944,N_3335,N_3149);
or U3945 (N_3945,N_3101,N_3311);
or U3946 (N_3946,N_3269,N_3056);
or U3947 (N_3947,N_3196,N_3353);
xor U3948 (N_3948,N_3399,N_3296);
nor U3949 (N_3949,N_3343,N_3102);
nand U3950 (N_3950,N_3350,N_3101);
and U3951 (N_3951,N_3156,N_3102);
nor U3952 (N_3952,N_3197,N_3075);
nor U3953 (N_3953,N_3141,N_3326);
xor U3954 (N_3954,N_3087,N_3236);
nand U3955 (N_3955,N_3244,N_3249);
xnor U3956 (N_3956,N_3370,N_3004);
nand U3957 (N_3957,N_3330,N_3213);
xnor U3958 (N_3958,N_3402,N_3336);
or U3959 (N_3959,N_3197,N_3278);
nor U3960 (N_3960,N_3135,N_3481);
and U3961 (N_3961,N_3136,N_3287);
and U3962 (N_3962,N_3232,N_3472);
and U3963 (N_3963,N_3438,N_3201);
nand U3964 (N_3964,N_3229,N_3288);
nor U3965 (N_3965,N_3027,N_3185);
nand U3966 (N_3966,N_3434,N_3346);
and U3967 (N_3967,N_3269,N_3368);
xnor U3968 (N_3968,N_3084,N_3342);
and U3969 (N_3969,N_3240,N_3237);
or U3970 (N_3970,N_3098,N_3397);
xnor U3971 (N_3971,N_3343,N_3117);
or U3972 (N_3972,N_3339,N_3243);
xnor U3973 (N_3973,N_3419,N_3433);
nor U3974 (N_3974,N_3481,N_3494);
and U3975 (N_3975,N_3022,N_3391);
nor U3976 (N_3976,N_3277,N_3051);
nor U3977 (N_3977,N_3352,N_3117);
and U3978 (N_3978,N_3175,N_3436);
nor U3979 (N_3979,N_3029,N_3439);
and U3980 (N_3980,N_3285,N_3413);
or U3981 (N_3981,N_3268,N_3236);
and U3982 (N_3982,N_3448,N_3173);
xnor U3983 (N_3983,N_3087,N_3332);
nand U3984 (N_3984,N_3262,N_3011);
xor U3985 (N_3985,N_3060,N_3011);
nor U3986 (N_3986,N_3208,N_3196);
and U3987 (N_3987,N_3307,N_3044);
nor U3988 (N_3988,N_3258,N_3036);
xor U3989 (N_3989,N_3462,N_3312);
nor U3990 (N_3990,N_3460,N_3123);
nand U3991 (N_3991,N_3108,N_3188);
xor U3992 (N_3992,N_3293,N_3156);
nor U3993 (N_3993,N_3444,N_3028);
nor U3994 (N_3994,N_3005,N_3416);
or U3995 (N_3995,N_3095,N_3358);
and U3996 (N_3996,N_3198,N_3060);
nor U3997 (N_3997,N_3498,N_3287);
nand U3998 (N_3998,N_3242,N_3458);
or U3999 (N_3999,N_3283,N_3177);
or U4000 (N_4000,N_3658,N_3755);
and U4001 (N_4001,N_3620,N_3889);
nand U4002 (N_4002,N_3602,N_3756);
xor U4003 (N_4003,N_3703,N_3858);
xor U4004 (N_4004,N_3971,N_3509);
nand U4005 (N_4005,N_3920,N_3916);
xor U4006 (N_4006,N_3938,N_3593);
nor U4007 (N_4007,N_3805,N_3885);
xor U4008 (N_4008,N_3734,N_3564);
or U4009 (N_4009,N_3953,N_3757);
nor U4010 (N_4010,N_3753,N_3935);
nor U4011 (N_4011,N_3918,N_3599);
nand U4012 (N_4012,N_3614,N_3568);
or U4013 (N_4013,N_3868,N_3813);
nor U4014 (N_4014,N_3978,N_3771);
or U4015 (N_4015,N_3500,N_3989);
xnor U4016 (N_4016,N_3949,N_3644);
and U4017 (N_4017,N_3700,N_3711);
nand U4018 (N_4018,N_3555,N_3779);
xor U4019 (N_4019,N_3527,N_3514);
and U4020 (N_4020,N_3840,N_3901);
and U4021 (N_4021,N_3905,N_3824);
nand U4022 (N_4022,N_3639,N_3580);
nor U4023 (N_4023,N_3649,N_3997);
and U4024 (N_4024,N_3607,N_3957);
and U4025 (N_4025,N_3547,N_3590);
nor U4026 (N_4026,N_3859,N_3714);
and U4027 (N_4027,N_3936,N_3542);
xnor U4028 (N_4028,N_3860,N_3770);
and U4029 (N_4029,N_3972,N_3549);
nor U4030 (N_4030,N_3544,N_3876);
and U4031 (N_4031,N_3629,N_3750);
nand U4032 (N_4032,N_3809,N_3898);
nand U4033 (N_4033,N_3698,N_3654);
nand U4034 (N_4034,N_3672,N_3783);
and U4035 (N_4035,N_3583,N_3545);
nand U4036 (N_4036,N_3811,N_3834);
or U4037 (N_4037,N_3954,N_3837);
nand U4038 (N_4038,N_3626,N_3836);
nand U4039 (N_4039,N_3539,N_3791);
xnor U4040 (N_4040,N_3579,N_3922);
xnor U4041 (N_4041,N_3724,N_3694);
xnor U4042 (N_4042,N_3592,N_3899);
or U4043 (N_4043,N_3710,N_3759);
nand U4044 (N_4044,N_3526,N_3845);
nand U4045 (N_4045,N_3719,N_3796);
nor U4046 (N_4046,N_3529,N_3630);
xor U4047 (N_4047,N_3652,N_3910);
nor U4048 (N_4048,N_3820,N_3812);
xnor U4049 (N_4049,N_3578,N_3573);
and U4050 (N_4050,N_3660,N_3844);
nor U4051 (N_4051,N_3569,N_3541);
nand U4052 (N_4052,N_3926,N_3775);
nor U4053 (N_4053,N_3874,N_3650);
and U4054 (N_4054,N_3913,N_3793);
xor U4055 (N_4055,N_3553,N_3772);
and U4056 (N_4056,N_3729,N_3653);
or U4057 (N_4057,N_3778,N_3921);
and U4058 (N_4058,N_3713,N_3810);
xor U4059 (N_4059,N_3803,N_3659);
nor U4060 (N_4060,N_3673,N_3808);
and U4061 (N_4061,N_3690,N_3524);
nand U4062 (N_4062,N_3671,N_3645);
nand U4063 (N_4063,N_3675,N_3574);
and U4064 (N_4064,N_3937,N_3768);
nor U4065 (N_4065,N_3893,N_3882);
xnor U4066 (N_4066,N_3685,N_3795);
and U4067 (N_4067,N_3642,N_3571);
xor U4068 (N_4068,N_3847,N_3519);
or U4069 (N_4069,N_3502,N_3942);
xnor U4070 (N_4070,N_3745,N_3829);
or U4071 (N_4071,N_3956,N_3966);
nand U4072 (N_4072,N_3854,N_3537);
nand U4073 (N_4073,N_3631,N_3709);
and U4074 (N_4074,N_3737,N_3567);
xnor U4075 (N_4075,N_3951,N_3973);
xnor U4076 (N_4076,N_3941,N_3680);
nor U4077 (N_4077,N_3914,N_3843);
and U4078 (N_4078,N_3887,N_3990);
nor U4079 (N_4079,N_3561,N_3543);
xor U4080 (N_4080,N_3870,N_3604);
xnor U4081 (N_4081,N_3624,N_3738);
xnor U4082 (N_4082,N_3670,N_3739);
or U4083 (N_4083,N_3531,N_3979);
and U4084 (N_4084,N_3575,N_3548);
and U4085 (N_4085,N_3508,N_3666);
and U4086 (N_4086,N_3948,N_3589);
nand U4087 (N_4087,N_3704,N_3877);
nor U4088 (N_4088,N_3798,N_3640);
and U4089 (N_4089,N_3967,N_3934);
or U4090 (N_4090,N_3594,N_3760);
nor U4091 (N_4091,N_3864,N_3897);
nor U4092 (N_4092,N_3688,N_3754);
and U4093 (N_4093,N_3985,N_3781);
or U4094 (N_4094,N_3664,N_3695);
xor U4095 (N_4095,N_3689,N_3662);
nor U4096 (N_4096,N_3947,N_3528);
or U4097 (N_4097,N_3610,N_3977);
and U4098 (N_4098,N_3535,N_3881);
or U4099 (N_4099,N_3983,N_3655);
or U4100 (N_4100,N_3944,N_3988);
and U4101 (N_4101,N_3681,N_3702);
and U4102 (N_4102,N_3828,N_3651);
and U4103 (N_4103,N_3995,N_3731);
nand U4104 (N_4104,N_3582,N_3677);
nor U4105 (N_4105,N_3939,N_3904);
nor U4106 (N_4106,N_3776,N_3628);
xor U4107 (N_4107,N_3801,N_3924);
or U4108 (N_4108,N_3740,N_3974);
or U4109 (N_4109,N_3699,N_3999);
or U4110 (N_4110,N_3641,N_3758);
nand U4111 (N_4111,N_3678,N_3669);
and U4112 (N_4112,N_3512,N_3917);
nor U4113 (N_4113,N_3786,N_3965);
nor U4114 (N_4114,N_3552,N_3929);
and U4115 (N_4115,N_3510,N_3706);
nand U4116 (N_4116,N_3540,N_3987);
or U4117 (N_4117,N_3618,N_3521);
and U4118 (N_4118,N_3636,N_3902);
nor U4119 (N_4119,N_3741,N_3777);
nand U4120 (N_4120,N_3912,N_3853);
nor U4121 (N_4121,N_3832,N_3523);
xnor U4122 (N_4122,N_3743,N_3606);
or U4123 (N_4123,N_3839,N_3950);
xor U4124 (N_4124,N_3855,N_3908);
nand U4125 (N_4125,N_3998,N_3774);
nand U4126 (N_4126,N_3800,N_3852);
xor U4127 (N_4127,N_3621,N_3980);
nor U4128 (N_4128,N_3861,N_3577);
nand U4129 (N_4129,N_3835,N_3946);
and U4130 (N_4130,N_3895,N_3749);
nor U4131 (N_4131,N_3718,N_3605);
nand U4132 (N_4132,N_3925,N_3984);
nor U4133 (N_4133,N_3586,N_3520);
nor U4134 (N_4134,N_3866,N_3725);
or U4135 (N_4135,N_3851,N_3576);
and U4136 (N_4136,N_3674,N_3790);
and U4137 (N_4137,N_3727,N_3634);
and U4138 (N_4138,N_3560,N_3748);
nand U4139 (N_4139,N_3900,N_3525);
nand U4140 (N_4140,N_3906,N_3716);
and U4141 (N_4141,N_3533,N_3960);
and U4142 (N_4142,N_3815,N_3682);
nand U4143 (N_4143,N_3883,N_3684);
nor U4144 (N_4144,N_3572,N_3773);
nand U4145 (N_4145,N_3890,N_3814);
and U4146 (N_4146,N_3986,N_3735);
nor U4147 (N_4147,N_3615,N_3744);
xnor U4148 (N_4148,N_3687,N_3507);
nand U4149 (N_4149,N_3516,N_3693);
and U4150 (N_4150,N_3884,N_3964);
nor U4151 (N_4151,N_3538,N_3993);
or U4152 (N_4152,N_3976,N_3581);
xnor U4153 (N_4153,N_3804,N_3784);
or U4154 (N_4154,N_3970,N_3785);
xor U4155 (N_4155,N_3907,N_3848);
and U4156 (N_4156,N_3943,N_3728);
and U4157 (N_4157,N_3886,N_3879);
xor U4158 (N_4158,N_3816,N_3894);
nor U4159 (N_4159,N_3697,N_3932);
nand U4160 (N_4160,N_3888,N_3746);
and U4161 (N_4161,N_3780,N_3633);
or U4162 (N_4162,N_3518,N_3646);
and U4163 (N_4163,N_3969,N_3736);
xor U4164 (N_4164,N_3534,N_3647);
nand U4165 (N_4165,N_3873,N_3701);
and U4166 (N_4166,N_3720,N_3940);
or U4167 (N_4167,N_3517,N_3821);
nor U4168 (N_4168,N_3503,N_3915);
and U4169 (N_4169,N_3627,N_3846);
nor U4170 (N_4170,N_3763,N_3764);
nand U4171 (N_4171,N_3557,N_3849);
nor U4172 (N_4172,N_3788,N_3623);
or U4173 (N_4173,N_3807,N_3601);
xnor U4174 (N_4174,N_3504,N_3822);
xor U4175 (N_4175,N_3730,N_3665);
nor U4176 (N_4176,N_3871,N_3992);
nor U4177 (N_4177,N_3622,N_3705);
and U4178 (N_4178,N_3691,N_3612);
and U4179 (N_4179,N_3663,N_3600);
xor U4180 (N_4180,N_3625,N_3880);
nor U4181 (N_4181,N_3945,N_3769);
nor U4182 (N_4182,N_3676,N_3955);
nor U4183 (N_4183,N_3536,N_3732);
nand U4184 (N_4184,N_3862,N_3532);
xnor U4185 (N_4185,N_3668,N_3850);
nand U4186 (N_4186,N_3715,N_3818);
xnor U4187 (N_4187,N_3707,N_3721);
or U4188 (N_4188,N_3617,N_3733);
xor U4189 (N_4189,N_3863,N_3991);
nand U4190 (N_4190,N_3661,N_3891);
and U4191 (N_4191,N_3643,N_3648);
or U4192 (N_4192,N_3831,N_3981);
and U4193 (N_4193,N_3767,N_3588);
and U4194 (N_4194,N_3782,N_3930);
nor U4195 (N_4195,N_3513,N_3751);
or U4196 (N_4196,N_3546,N_3789);
or U4197 (N_4197,N_3869,N_3802);
nor U4198 (N_4198,N_3609,N_3562);
xor U4199 (N_4199,N_3952,N_3928);
xor U4200 (N_4200,N_3596,N_3657);
or U4201 (N_4201,N_3591,N_3530);
nor U4202 (N_4202,N_3505,N_3878);
and U4203 (N_4203,N_3996,N_3766);
nand U4204 (N_4204,N_3806,N_3686);
xnor U4205 (N_4205,N_3501,N_3867);
or U4206 (N_4206,N_3742,N_3556);
or U4207 (N_4207,N_3919,N_3827);
nor U4208 (N_4208,N_3968,N_3747);
xnor U4209 (N_4209,N_3717,N_3830);
or U4210 (N_4210,N_3522,N_3559);
or U4211 (N_4211,N_3723,N_3696);
nor U4212 (N_4212,N_3585,N_3558);
nand U4213 (N_4213,N_3823,N_3959);
nand U4214 (N_4214,N_3927,N_3616);
or U4215 (N_4215,N_3667,N_3911);
or U4216 (N_4216,N_3762,N_3598);
or U4217 (N_4217,N_3958,N_3683);
nor U4218 (N_4218,N_3975,N_3841);
xnor U4219 (N_4219,N_3825,N_3638);
and U4220 (N_4220,N_3563,N_3637);
xnor U4221 (N_4221,N_3817,N_3587);
nand U4222 (N_4222,N_3797,N_3799);
xnor U4223 (N_4223,N_3909,N_3708);
nand U4224 (N_4224,N_3565,N_3712);
nand U4225 (N_4225,N_3752,N_3597);
nand U4226 (N_4226,N_3875,N_3857);
and U4227 (N_4227,N_3515,N_3962);
and U4228 (N_4228,N_3963,N_3933);
or U4229 (N_4229,N_3872,N_3826);
xnor U4230 (N_4230,N_3679,N_3833);
nand U4231 (N_4231,N_3982,N_3961);
nand U4232 (N_4232,N_3765,N_3656);
nand U4233 (N_4233,N_3842,N_3692);
or U4234 (N_4234,N_3792,N_3819);
and U4235 (N_4235,N_3722,N_3584);
nor U4236 (N_4236,N_3896,N_3603);
nor U4237 (N_4237,N_3613,N_3856);
nand U4238 (N_4238,N_3923,N_3635);
or U4239 (N_4239,N_3619,N_3595);
and U4240 (N_4240,N_3892,N_3611);
nor U4241 (N_4241,N_3554,N_3794);
xnor U4242 (N_4242,N_3838,N_3787);
nor U4243 (N_4243,N_3570,N_3761);
or U4244 (N_4244,N_3551,N_3994);
or U4245 (N_4245,N_3865,N_3903);
xnor U4246 (N_4246,N_3566,N_3726);
nor U4247 (N_4247,N_3931,N_3511);
nand U4248 (N_4248,N_3632,N_3550);
nand U4249 (N_4249,N_3608,N_3506);
nor U4250 (N_4250,N_3821,N_3882);
nand U4251 (N_4251,N_3682,N_3873);
or U4252 (N_4252,N_3677,N_3644);
nor U4253 (N_4253,N_3572,N_3805);
nor U4254 (N_4254,N_3982,N_3956);
nor U4255 (N_4255,N_3632,N_3687);
or U4256 (N_4256,N_3955,N_3610);
nor U4257 (N_4257,N_3537,N_3558);
or U4258 (N_4258,N_3592,N_3710);
nand U4259 (N_4259,N_3609,N_3665);
or U4260 (N_4260,N_3866,N_3909);
nor U4261 (N_4261,N_3569,N_3955);
nor U4262 (N_4262,N_3524,N_3629);
xnor U4263 (N_4263,N_3734,N_3748);
nand U4264 (N_4264,N_3970,N_3645);
xor U4265 (N_4265,N_3855,N_3816);
nor U4266 (N_4266,N_3621,N_3778);
or U4267 (N_4267,N_3725,N_3541);
xnor U4268 (N_4268,N_3927,N_3791);
nor U4269 (N_4269,N_3685,N_3913);
or U4270 (N_4270,N_3715,N_3841);
and U4271 (N_4271,N_3514,N_3849);
and U4272 (N_4272,N_3662,N_3731);
nand U4273 (N_4273,N_3877,N_3812);
or U4274 (N_4274,N_3572,N_3802);
and U4275 (N_4275,N_3931,N_3854);
nor U4276 (N_4276,N_3856,N_3748);
nand U4277 (N_4277,N_3717,N_3537);
and U4278 (N_4278,N_3687,N_3868);
xnor U4279 (N_4279,N_3850,N_3989);
or U4280 (N_4280,N_3684,N_3613);
xnor U4281 (N_4281,N_3729,N_3954);
or U4282 (N_4282,N_3578,N_3971);
or U4283 (N_4283,N_3907,N_3674);
xnor U4284 (N_4284,N_3602,N_3728);
or U4285 (N_4285,N_3691,N_3816);
nand U4286 (N_4286,N_3959,N_3859);
and U4287 (N_4287,N_3650,N_3632);
and U4288 (N_4288,N_3670,N_3564);
or U4289 (N_4289,N_3942,N_3510);
nor U4290 (N_4290,N_3705,N_3822);
nor U4291 (N_4291,N_3620,N_3786);
xnor U4292 (N_4292,N_3699,N_3963);
xor U4293 (N_4293,N_3690,N_3782);
nor U4294 (N_4294,N_3556,N_3968);
nor U4295 (N_4295,N_3876,N_3504);
and U4296 (N_4296,N_3837,N_3852);
nand U4297 (N_4297,N_3816,N_3811);
nand U4298 (N_4298,N_3700,N_3914);
xor U4299 (N_4299,N_3913,N_3843);
or U4300 (N_4300,N_3668,N_3778);
xnor U4301 (N_4301,N_3976,N_3957);
nand U4302 (N_4302,N_3536,N_3574);
xnor U4303 (N_4303,N_3898,N_3566);
nor U4304 (N_4304,N_3549,N_3826);
nand U4305 (N_4305,N_3522,N_3517);
or U4306 (N_4306,N_3693,N_3737);
or U4307 (N_4307,N_3702,N_3563);
nor U4308 (N_4308,N_3915,N_3903);
and U4309 (N_4309,N_3922,N_3730);
and U4310 (N_4310,N_3920,N_3903);
and U4311 (N_4311,N_3691,N_3770);
xnor U4312 (N_4312,N_3711,N_3526);
or U4313 (N_4313,N_3799,N_3504);
or U4314 (N_4314,N_3670,N_3528);
and U4315 (N_4315,N_3653,N_3855);
nand U4316 (N_4316,N_3684,N_3681);
nor U4317 (N_4317,N_3861,N_3544);
and U4318 (N_4318,N_3951,N_3882);
or U4319 (N_4319,N_3933,N_3967);
or U4320 (N_4320,N_3517,N_3682);
xor U4321 (N_4321,N_3843,N_3560);
nand U4322 (N_4322,N_3831,N_3682);
and U4323 (N_4323,N_3537,N_3670);
and U4324 (N_4324,N_3813,N_3774);
or U4325 (N_4325,N_3779,N_3959);
or U4326 (N_4326,N_3545,N_3776);
xnor U4327 (N_4327,N_3753,N_3502);
nand U4328 (N_4328,N_3660,N_3829);
nand U4329 (N_4329,N_3757,N_3817);
nand U4330 (N_4330,N_3885,N_3559);
nor U4331 (N_4331,N_3713,N_3772);
or U4332 (N_4332,N_3945,N_3730);
nand U4333 (N_4333,N_3537,N_3933);
nor U4334 (N_4334,N_3897,N_3733);
nand U4335 (N_4335,N_3876,N_3545);
and U4336 (N_4336,N_3775,N_3783);
nor U4337 (N_4337,N_3967,N_3725);
xor U4338 (N_4338,N_3824,N_3517);
xor U4339 (N_4339,N_3731,N_3628);
xnor U4340 (N_4340,N_3741,N_3771);
and U4341 (N_4341,N_3527,N_3791);
xnor U4342 (N_4342,N_3749,N_3807);
nand U4343 (N_4343,N_3848,N_3965);
and U4344 (N_4344,N_3787,N_3685);
nand U4345 (N_4345,N_3692,N_3717);
or U4346 (N_4346,N_3762,N_3742);
nor U4347 (N_4347,N_3518,N_3923);
and U4348 (N_4348,N_3673,N_3970);
xor U4349 (N_4349,N_3670,N_3792);
nand U4350 (N_4350,N_3562,N_3810);
nand U4351 (N_4351,N_3792,N_3510);
or U4352 (N_4352,N_3763,N_3775);
xor U4353 (N_4353,N_3807,N_3536);
nor U4354 (N_4354,N_3761,N_3675);
xor U4355 (N_4355,N_3557,N_3535);
nand U4356 (N_4356,N_3545,N_3956);
nor U4357 (N_4357,N_3704,N_3775);
nor U4358 (N_4358,N_3652,N_3677);
or U4359 (N_4359,N_3679,N_3940);
nor U4360 (N_4360,N_3764,N_3613);
xnor U4361 (N_4361,N_3863,N_3809);
xnor U4362 (N_4362,N_3565,N_3575);
and U4363 (N_4363,N_3853,N_3516);
or U4364 (N_4364,N_3670,N_3607);
or U4365 (N_4365,N_3848,N_3704);
or U4366 (N_4366,N_3842,N_3901);
nand U4367 (N_4367,N_3736,N_3728);
or U4368 (N_4368,N_3813,N_3758);
xor U4369 (N_4369,N_3583,N_3586);
nor U4370 (N_4370,N_3755,N_3808);
xnor U4371 (N_4371,N_3932,N_3634);
xor U4372 (N_4372,N_3618,N_3614);
and U4373 (N_4373,N_3684,N_3519);
nor U4374 (N_4374,N_3988,N_3864);
xor U4375 (N_4375,N_3940,N_3871);
nand U4376 (N_4376,N_3720,N_3668);
and U4377 (N_4377,N_3735,N_3981);
nor U4378 (N_4378,N_3565,N_3704);
or U4379 (N_4379,N_3865,N_3501);
and U4380 (N_4380,N_3778,N_3982);
or U4381 (N_4381,N_3613,N_3769);
nor U4382 (N_4382,N_3713,N_3840);
nand U4383 (N_4383,N_3838,N_3525);
or U4384 (N_4384,N_3715,N_3772);
nand U4385 (N_4385,N_3843,N_3628);
nor U4386 (N_4386,N_3667,N_3881);
nor U4387 (N_4387,N_3594,N_3876);
and U4388 (N_4388,N_3746,N_3805);
nor U4389 (N_4389,N_3761,N_3647);
xor U4390 (N_4390,N_3567,N_3669);
or U4391 (N_4391,N_3845,N_3553);
nand U4392 (N_4392,N_3660,N_3896);
and U4393 (N_4393,N_3619,N_3739);
xnor U4394 (N_4394,N_3716,N_3736);
and U4395 (N_4395,N_3600,N_3893);
or U4396 (N_4396,N_3537,N_3591);
or U4397 (N_4397,N_3764,N_3862);
and U4398 (N_4398,N_3530,N_3886);
nor U4399 (N_4399,N_3532,N_3504);
and U4400 (N_4400,N_3608,N_3552);
nand U4401 (N_4401,N_3929,N_3606);
nand U4402 (N_4402,N_3815,N_3952);
xnor U4403 (N_4403,N_3635,N_3826);
xnor U4404 (N_4404,N_3606,N_3780);
nand U4405 (N_4405,N_3580,N_3761);
nand U4406 (N_4406,N_3778,N_3888);
nor U4407 (N_4407,N_3672,N_3596);
and U4408 (N_4408,N_3965,N_3881);
or U4409 (N_4409,N_3972,N_3507);
nand U4410 (N_4410,N_3583,N_3975);
or U4411 (N_4411,N_3634,N_3931);
nor U4412 (N_4412,N_3788,N_3524);
and U4413 (N_4413,N_3699,N_3525);
nand U4414 (N_4414,N_3673,N_3556);
and U4415 (N_4415,N_3931,N_3618);
and U4416 (N_4416,N_3658,N_3547);
xor U4417 (N_4417,N_3506,N_3818);
nand U4418 (N_4418,N_3775,N_3524);
nor U4419 (N_4419,N_3655,N_3610);
xnor U4420 (N_4420,N_3668,N_3763);
nor U4421 (N_4421,N_3670,N_3582);
nor U4422 (N_4422,N_3618,N_3717);
nand U4423 (N_4423,N_3581,N_3638);
nand U4424 (N_4424,N_3906,N_3980);
xor U4425 (N_4425,N_3854,N_3642);
or U4426 (N_4426,N_3886,N_3966);
xnor U4427 (N_4427,N_3900,N_3812);
nor U4428 (N_4428,N_3610,N_3904);
xnor U4429 (N_4429,N_3502,N_3877);
xor U4430 (N_4430,N_3523,N_3648);
nor U4431 (N_4431,N_3704,N_3884);
and U4432 (N_4432,N_3551,N_3770);
and U4433 (N_4433,N_3638,N_3726);
xnor U4434 (N_4434,N_3590,N_3822);
and U4435 (N_4435,N_3845,N_3906);
xnor U4436 (N_4436,N_3568,N_3530);
xnor U4437 (N_4437,N_3595,N_3523);
and U4438 (N_4438,N_3918,N_3862);
xnor U4439 (N_4439,N_3684,N_3915);
or U4440 (N_4440,N_3695,N_3705);
and U4441 (N_4441,N_3912,N_3724);
nor U4442 (N_4442,N_3709,N_3611);
or U4443 (N_4443,N_3921,N_3792);
and U4444 (N_4444,N_3661,N_3912);
or U4445 (N_4445,N_3814,N_3726);
xor U4446 (N_4446,N_3582,N_3675);
or U4447 (N_4447,N_3835,N_3850);
nor U4448 (N_4448,N_3596,N_3500);
xor U4449 (N_4449,N_3518,N_3898);
nand U4450 (N_4450,N_3704,N_3508);
xnor U4451 (N_4451,N_3699,N_3866);
xnor U4452 (N_4452,N_3711,N_3551);
or U4453 (N_4453,N_3659,N_3902);
or U4454 (N_4454,N_3822,N_3572);
nor U4455 (N_4455,N_3889,N_3962);
xor U4456 (N_4456,N_3987,N_3682);
and U4457 (N_4457,N_3701,N_3693);
xnor U4458 (N_4458,N_3674,N_3754);
nor U4459 (N_4459,N_3873,N_3833);
nand U4460 (N_4460,N_3594,N_3698);
and U4461 (N_4461,N_3850,N_3538);
nand U4462 (N_4462,N_3969,N_3821);
and U4463 (N_4463,N_3574,N_3818);
nand U4464 (N_4464,N_3686,N_3638);
nor U4465 (N_4465,N_3944,N_3582);
xnor U4466 (N_4466,N_3521,N_3510);
nand U4467 (N_4467,N_3913,N_3670);
nor U4468 (N_4468,N_3860,N_3513);
nand U4469 (N_4469,N_3542,N_3551);
nor U4470 (N_4470,N_3732,N_3914);
xor U4471 (N_4471,N_3959,N_3887);
nand U4472 (N_4472,N_3782,N_3662);
or U4473 (N_4473,N_3719,N_3905);
or U4474 (N_4474,N_3660,N_3920);
nand U4475 (N_4475,N_3713,N_3925);
and U4476 (N_4476,N_3993,N_3524);
nor U4477 (N_4477,N_3855,N_3937);
nand U4478 (N_4478,N_3615,N_3860);
nand U4479 (N_4479,N_3607,N_3707);
nor U4480 (N_4480,N_3893,N_3653);
xnor U4481 (N_4481,N_3648,N_3633);
and U4482 (N_4482,N_3586,N_3684);
nand U4483 (N_4483,N_3831,N_3867);
nand U4484 (N_4484,N_3723,N_3955);
and U4485 (N_4485,N_3733,N_3507);
or U4486 (N_4486,N_3558,N_3817);
xnor U4487 (N_4487,N_3732,N_3816);
and U4488 (N_4488,N_3518,N_3791);
or U4489 (N_4489,N_3705,N_3710);
nand U4490 (N_4490,N_3826,N_3797);
nor U4491 (N_4491,N_3902,N_3585);
and U4492 (N_4492,N_3833,N_3799);
xor U4493 (N_4493,N_3925,N_3959);
nor U4494 (N_4494,N_3584,N_3605);
xnor U4495 (N_4495,N_3721,N_3829);
or U4496 (N_4496,N_3785,N_3604);
xnor U4497 (N_4497,N_3627,N_3619);
and U4498 (N_4498,N_3927,N_3901);
nand U4499 (N_4499,N_3802,N_3822);
nand U4500 (N_4500,N_4477,N_4041);
nand U4501 (N_4501,N_4424,N_4339);
xnor U4502 (N_4502,N_4014,N_4389);
nor U4503 (N_4503,N_4430,N_4116);
and U4504 (N_4504,N_4354,N_4481);
nor U4505 (N_4505,N_4049,N_4406);
or U4506 (N_4506,N_4181,N_4179);
nand U4507 (N_4507,N_4268,N_4472);
nor U4508 (N_4508,N_4066,N_4242);
xor U4509 (N_4509,N_4064,N_4186);
and U4510 (N_4510,N_4250,N_4208);
xnor U4511 (N_4511,N_4375,N_4018);
nor U4512 (N_4512,N_4383,N_4396);
xnor U4513 (N_4513,N_4056,N_4391);
xor U4514 (N_4514,N_4478,N_4305);
nor U4515 (N_4515,N_4153,N_4190);
nor U4516 (N_4516,N_4008,N_4087);
and U4517 (N_4517,N_4351,N_4295);
and U4518 (N_4518,N_4281,N_4445);
and U4519 (N_4519,N_4042,N_4177);
and U4520 (N_4520,N_4244,N_4372);
and U4521 (N_4521,N_4310,N_4429);
xnor U4522 (N_4522,N_4058,N_4350);
or U4523 (N_4523,N_4228,N_4083);
nor U4524 (N_4524,N_4134,N_4456);
nand U4525 (N_4525,N_4303,N_4401);
and U4526 (N_4526,N_4100,N_4390);
nor U4527 (N_4527,N_4031,N_4026);
nor U4528 (N_4528,N_4203,N_4273);
xnor U4529 (N_4529,N_4357,N_4495);
and U4530 (N_4530,N_4236,N_4223);
nand U4531 (N_4531,N_4471,N_4076);
nor U4532 (N_4532,N_4157,N_4355);
nor U4533 (N_4533,N_4328,N_4422);
nor U4534 (N_4534,N_4297,N_4260);
nor U4535 (N_4535,N_4000,N_4394);
xor U4536 (N_4536,N_4262,N_4189);
xnor U4537 (N_4537,N_4413,N_4140);
nand U4538 (N_4538,N_4086,N_4493);
nor U4539 (N_4539,N_4377,N_4002);
and U4540 (N_4540,N_4022,N_4312);
xor U4541 (N_4541,N_4367,N_4443);
and U4542 (N_4542,N_4415,N_4340);
and U4543 (N_4543,N_4440,N_4419);
nand U4544 (N_4544,N_4338,N_4470);
or U4545 (N_4545,N_4194,N_4270);
nand U4546 (N_4546,N_4129,N_4165);
xor U4547 (N_4547,N_4015,N_4252);
nand U4548 (N_4548,N_4462,N_4089);
nand U4549 (N_4549,N_4239,N_4001);
nor U4550 (N_4550,N_4484,N_4095);
nand U4551 (N_4551,N_4258,N_4299);
nand U4552 (N_4552,N_4418,N_4011);
xnor U4553 (N_4553,N_4167,N_4040);
or U4554 (N_4554,N_4376,N_4085);
nand U4555 (N_4555,N_4274,N_4150);
or U4556 (N_4556,N_4004,N_4216);
and U4557 (N_4557,N_4352,N_4335);
or U4558 (N_4558,N_4021,N_4451);
xor U4559 (N_4559,N_4407,N_4233);
or U4560 (N_4560,N_4098,N_4173);
and U4561 (N_4561,N_4392,N_4143);
nand U4562 (N_4562,N_4183,N_4382);
or U4563 (N_4563,N_4046,N_4304);
or U4564 (N_4564,N_4154,N_4020);
or U4565 (N_4565,N_4205,N_4411);
xor U4566 (N_4566,N_4023,N_4084);
nand U4567 (N_4567,N_4296,N_4090);
xor U4568 (N_4568,N_4452,N_4290);
nor U4569 (N_4569,N_4346,N_4119);
xnor U4570 (N_4570,N_4038,N_4343);
or U4571 (N_4571,N_4264,N_4185);
nand U4572 (N_4572,N_4199,N_4210);
nand U4573 (N_4573,N_4436,N_4489);
or U4574 (N_4574,N_4044,N_4403);
nand U4575 (N_4575,N_4373,N_4218);
nand U4576 (N_4576,N_4212,N_4370);
nor U4577 (N_4577,N_4163,N_4192);
xnor U4578 (N_4578,N_4059,N_4364);
or U4579 (N_4579,N_4259,N_4423);
nor U4580 (N_4580,N_4490,N_4425);
nand U4581 (N_4581,N_4213,N_4149);
and U4582 (N_4582,N_4427,N_4234);
nand U4583 (N_4583,N_4444,N_4318);
nor U4584 (N_4584,N_4263,N_4385);
nor U4585 (N_4585,N_4457,N_4209);
nand U4586 (N_4586,N_4348,N_4169);
nand U4587 (N_4587,N_4308,N_4182);
nand U4588 (N_4588,N_4369,N_4298);
or U4589 (N_4589,N_4459,N_4077);
nand U4590 (N_4590,N_4317,N_4465);
and U4591 (N_4591,N_4243,N_4301);
and U4592 (N_4592,N_4287,N_4278);
nor U4593 (N_4593,N_4139,N_4068);
nand U4594 (N_4594,N_4421,N_4475);
and U4595 (N_4595,N_4334,N_4437);
nor U4596 (N_4596,N_4065,N_4039);
nor U4597 (N_4597,N_4285,N_4131);
xor U4598 (N_4598,N_4078,N_4349);
xnor U4599 (N_4599,N_4051,N_4446);
xnor U4600 (N_4600,N_4410,N_4055);
and U4601 (N_4601,N_4221,N_4237);
and U4602 (N_4602,N_4327,N_4034);
nand U4603 (N_4603,N_4017,N_4473);
nand U4604 (N_4604,N_4091,N_4126);
xor U4605 (N_4605,N_4045,N_4172);
xnor U4606 (N_4606,N_4107,N_4111);
and U4607 (N_4607,N_4109,N_4271);
nand U4608 (N_4608,N_4267,N_4054);
xnor U4609 (N_4609,N_4093,N_4013);
nand U4610 (N_4610,N_4487,N_4476);
and U4611 (N_4611,N_4247,N_4345);
or U4612 (N_4612,N_4479,N_4279);
xor U4613 (N_4613,N_4101,N_4442);
and U4614 (N_4614,N_4499,N_4144);
nor U4615 (N_4615,N_4099,N_4047);
or U4616 (N_4616,N_4486,N_4282);
or U4617 (N_4617,N_4070,N_4253);
xor U4618 (N_4618,N_4255,N_4012);
xor U4619 (N_4619,N_4032,N_4368);
xor U4620 (N_4620,N_4288,N_4151);
xor U4621 (N_4621,N_4311,N_4344);
nand U4622 (N_4622,N_4381,N_4329);
nor U4623 (N_4623,N_4409,N_4198);
nand U4624 (N_4624,N_4461,N_4016);
nor U4625 (N_4625,N_4324,N_4088);
nand U4626 (N_4626,N_4230,N_4130);
nand U4627 (N_4627,N_4359,N_4276);
nand U4628 (N_4628,N_4280,N_4166);
xnor U4629 (N_4629,N_4332,N_4314);
xnor U4630 (N_4630,N_4162,N_4191);
or U4631 (N_4631,N_4480,N_4283);
and U4632 (N_4632,N_4460,N_4148);
and U4633 (N_4633,N_4463,N_4482);
nor U4634 (N_4634,N_4112,N_4467);
or U4635 (N_4635,N_4306,N_4438);
or U4636 (N_4636,N_4062,N_4071);
or U4637 (N_4637,N_4206,N_4275);
nor U4638 (N_4638,N_4320,N_4196);
xnor U4639 (N_4639,N_4135,N_4245);
xnor U4640 (N_4640,N_4417,N_4171);
or U4641 (N_4641,N_4037,N_4384);
nor U4642 (N_4642,N_4175,N_4316);
xor U4643 (N_4643,N_4300,N_4399);
and U4644 (N_4644,N_4096,N_4204);
xor U4645 (N_4645,N_4257,N_4488);
or U4646 (N_4646,N_4050,N_4336);
or U4647 (N_4647,N_4426,N_4127);
xnor U4648 (N_4648,N_4072,N_4265);
nand U4649 (N_4649,N_4362,N_4374);
nand U4650 (N_4650,N_4118,N_4035);
nand U4651 (N_4651,N_4025,N_4269);
nor U4652 (N_4652,N_4075,N_4365);
nor U4653 (N_4653,N_4217,N_4128);
nor U4654 (N_4654,N_4067,N_4235);
or U4655 (N_4655,N_4284,N_4238);
or U4656 (N_4656,N_4103,N_4092);
xor U4657 (N_4657,N_4496,N_4497);
nand U4658 (N_4658,N_4207,N_4361);
xor U4659 (N_4659,N_4356,N_4358);
nand U4660 (N_4660,N_4286,N_4105);
or U4661 (N_4661,N_4492,N_4033);
and U4662 (N_4662,N_4138,N_4132);
xor U4663 (N_4663,N_4309,N_4319);
nor U4664 (N_4664,N_4498,N_4211);
or U4665 (N_4665,N_4420,N_4330);
or U4666 (N_4666,N_4435,N_4469);
xnor U4667 (N_4667,N_4387,N_4176);
nor U4668 (N_4668,N_4222,N_4102);
nand U4669 (N_4669,N_4048,N_4455);
and U4670 (N_4670,N_4184,N_4246);
or U4671 (N_4671,N_4395,N_4029);
xor U4672 (N_4672,N_4293,N_4024);
xnor U4673 (N_4673,N_4491,N_4404);
nand U4674 (N_4674,N_4082,N_4378);
or U4675 (N_4675,N_4069,N_4322);
and U4676 (N_4676,N_4178,N_4402);
xnor U4677 (N_4677,N_4219,N_4225);
or U4678 (N_4678,N_4454,N_4115);
or U4679 (N_4679,N_4168,N_4241);
nor U4680 (N_4680,N_4120,N_4214);
or U4681 (N_4681,N_4261,N_4123);
xnor U4682 (N_4682,N_4447,N_4122);
and U4683 (N_4683,N_4007,N_4379);
xor U4684 (N_4684,N_4360,N_4019);
xor U4685 (N_4685,N_4380,N_4152);
nand U4686 (N_4686,N_4197,N_4195);
and U4687 (N_4687,N_4081,N_4146);
nand U4688 (N_4688,N_4458,N_4405);
nand U4689 (N_4689,N_4159,N_4272);
or U4690 (N_4690,N_4448,N_4254);
or U4691 (N_4691,N_4202,N_4313);
xnor U4692 (N_4692,N_4124,N_4494);
nand U4693 (N_4693,N_4400,N_4028);
nand U4694 (N_4694,N_4333,N_4291);
and U4695 (N_4695,N_4043,N_4009);
or U4696 (N_4696,N_4468,N_4412);
or U4697 (N_4697,N_4227,N_4485);
and U4698 (N_4698,N_4439,N_4200);
and U4699 (N_4699,N_4441,N_4188);
nor U4700 (N_4700,N_4342,N_4450);
xnor U4701 (N_4701,N_4136,N_4057);
xnor U4702 (N_4702,N_4256,N_4158);
nor U4703 (N_4703,N_4156,N_4231);
xnor U4704 (N_4704,N_4408,N_4137);
and U4705 (N_4705,N_4155,N_4326);
nor U4706 (N_4706,N_4141,N_4170);
or U4707 (N_4707,N_4353,N_4226);
nor U4708 (N_4708,N_4347,N_4125);
and U4709 (N_4709,N_4398,N_4414);
xor U4710 (N_4710,N_4145,N_4073);
or U4711 (N_4711,N_4117,N_4164);
nand U4712 (N_4712,N_4315,N_4337);
nand U4713 (N_4713,N_4114,N_4121);
or U4714 (N_4714,N_4294,N_4113);
nand U4715 (N_4715,N_4321,N_4449);
and U4716 (N_4716,N_4393,N_4386);
or U4717 (N_4717,N_4010,N_4302);
and U4718 (N_4718,N_4464,N_4036);
or U4719 (N_4719,N_4060,N_4174);
xor U4720 (N_4720,N_4248,N_4266);
or U4721 (N_4721,N_4142,N_4193);
or U4722 (N_4722,N_4388,N_4079);
or U4723 (N_4723,N_4106,N_4292);
xor U4724 (N_4724,N_4277,N_4187);
nor U4725 (N_4725,N_4249,N_4363);
and U4726 (N_4726,N_4431,N_4307);
xor U4727 (N_4727,N_4289,N_4453);
and U4728 (N_4728,N_4104,N_4433);
nor U4729 (N_4729,N_4220,N_4331);
nand U4730 (N_4730,N_4063,N_4232);
nor U4731 (N_4731,N_4052,N_4416);
xnor U4732 (N_4732,N_4229,N_4428);
and U4733 (N_4733,N_4074,N_4432);
or U4734 (N_4734,N_4147,N_4240);
nor U4735 (N_4735,N_4466,N_4094);
nand U4736 (N_4736,N_4341,N_4474);
xor U4737 (N_4737,N_4201,N_4161);
or U4738 (N_4738,N_4030,N_4110);
nand U4739 (N_4739,N_4434,N_4097);
nor U4740 (N_4740,N_4133,N_4061);
or U4741 (N_4741,N_4027,N_4323);
nand U4742 (N_4742,N_4003,N_4108);
and U4743 (N_4743,N_4483,N_4160);
nand U4744 (N_4744,N_4006,N_4397);
nor U4745 (N_4745,N_4325,N_4371);
or U4746 (N_4746,N_4366,N_4180);
nor U4747 (N_4747,N_4215,N_4005);
nor U4748 (N_4748,N_4053,N_4251);
and U4749 (N_4749,N_4080,N_4224);
and U4750 (N_4750,N_4078,N_4123);
xnor U4751 (N_4751,N_4398,N_4423);
xnor U4752 (N_4752,N_4457,N_4255);
and U4753 (N_4753,N_4256,N_4306);
or U4754 (N_4754,N_4161,N_4271);
and U4755 (N_4755,N_4196,N_4052);
nor U4756 (N_4756,N_4291,N_4156);
xor U4757 (N_4757,N_4477,N_4171);
or U4758 (N_4758,N_4343,N_4193);
xnor U4759 (N_4759,N_4086,N_4242);
nor U4760 (N_4760,N_4312,N_4480);
or U4761 (N_4761,N_4076,N_4085);
xor U4762 (N_4762,N_4378,N_4323);
xor U4763 (N_4763,N_4067,N_4068);
and U4764 (N_4764,N_4043,N_4235);
xnor U4765 (N_4765,N_4445,N_4164);
nand U4766 (N_4766,N_4202,N_4015);
xnor U4767 (N_4767,N_4376,N_4081);
xnor U4768 (N_4768,N_4384,N_4330);
or U4769 (N_4769,N_4180,N_4057);
xor U4770 (N_4770,N_4023,N_4134);
and U4771 (N_4771,N_4163,N_4328);
or U4772 (N_4772,N_4474,N_4196);
or U4773 (N_4773,N_4172,N_4106);
or U4774 (N_4774,N_4319,N_4335);
nor U4775 (N_4775,N_4460,N_4471);
xnor U4776 (N_4776,N_4106,N_4140);
nor U4777 (N_4777,N_4326,N_4234);
nor U4778 (N_4778,N_4307,N_4439);
or U4779 (N_4779,N_4420,N_4069);
nor U4780 (N_4780,N_4452,N_4314);
nor U4781 (N_4781,N_4340,N_4380);
nand U4782 (N_4782,N_4473,N_4034);
nor U4783 (N_4783,N_4266,N_4285);
nor U4784 (N_4784,N_4269,N_4425);
or U4785 (N_4785,N_4204,N_4172);
and U4786 (N_4786,N_4192,N_4006);
xnor U4787 (N_4787,N_4347,N_4211);
and U4788 (N_4788,N_4462,N_4265);
nor U4789 (N_4789,N_4400,N_4158);
nand U4790 (N_4790,N_4352,N_4277);
and U4791 (N_4791,N_4039,N_4007);
nor U4792 (N_4792,N_4191,N_4293);
nand U4793 (N_4793,N_4149,N_4372);
nor U4794 (N_4794,N_4208,N_4113);
or U4795 (N_4795,N_4410,N_4402);
xor U4796 (N_4796,N_4205,N_4356);
nand U4797 (N_4797,N_4268,N_4029);
xor U4798 (N_4798,N_4249,N_4250);
nor U4799 (N_4799,N_4285,N_4272);
or U4800 (N_4800,N_4048,N_4318);
nand U4801 (N_4801,N_4196,N_4413);
xnor U4802 (N_4802,N_4336,N_4042);
xor U4803 (N_4803,N_4409,N_4152);
and U4804 (N_4804,N_4277,N_4336);
nand U4805 (N_4805,N_4234,N_4330);
nand U4806 (N_4806,N_4010,N_4149);
and U4807 (N_4807,N_4264,N_4084);
and U4808 (N_4808,N_4216,N_4193);
or U4809 (N_4809,N_4029,N_4461);
and U4810 (N_4810,N_4396,N_4015);
or U4811 (N_4811,N_4026,N_4122);
nor U4812 (N_4812,N_4379,N_4306);
nand U4813 (N_4813,N_4306,N_4406);
nand U4814 (N_4814,N_4459,N_4183);
and U4815 (N_4815,N_4195,N_4348);
or U4816 (N_4816,N_4027,N_4419);
nand U4817 (N_4817,N_4112,N_4083);
xor U4818 (N_4818,N_4194,N_4311);
nand U4819 (N_4819,N_4317,N_4199);
nor U4820 (N_4820,N_4217,N_4200);
and U4821 (N_4821,N_4053,N_4264);
and U4822 (N_4822,N_4121,N_4211);
or U4823 (N_4823,N_4227,N_4076);
xor U4824 (N_4824,N_4055,N_4001);
xnor U4825 (N_4825,N_4113,N_4424);
and U4826 (N_4826,N_4324,N_4475);
and U4827 (N_4827,N_4196,N_4078);
nor U4828 (N_4828,N_4045,N_4063);
nor U4829 (N_4829,N_4492,N_4133);
xor U4830 (N_4830,N_4257,N_4101);
and U4831 (N_4831,N_4104,N_4368);
or U4832 (N_4832,N_4126,N_4471);
nor U4833 (N_4833,N_4174,N_4480);
xnor U4834 (N_4834,N_4097,N_4043);
xor U4835 (N_4835,N_4232,N_4200);
and U4836 (N_4836,N_4042,N_4198);
or U4837 (N_4837,N_4038,N_4375);
nor U4838 (N_4838,N_4369,N_4457);
xor U4839 (N_4839,N_4214,N_4418);
nand U4840 (N_4840,N_4123,N_4380);
nand U4841 (N_4841,N_4166,N_4390);
nand U4842 (N_4842,N_4158,N_4006);
and U4843 (N_4843,N_4308,N_4277);
xnor U4844 (N_4844,N_4315,N_4498);
and U4845 (N_4845,N_4238,N_4278);
xnor U4846 (N_4846,N_4325,N_4227);
or U4847 (N_4847,N_4195,N_4455);
xnor U4848 (N_4848,N_4481,N_4051);
and U4849 (N_4849,N_4068,N_4224);
xnor U4850 (N_4850,N_4102,N_4150);
xor U4851 (N_4851,N_4065,N_4485);
nand U4852 (N_4852,N_4193,N_4450);
or U4853 (N_4853,N_4178,N_4143);
or U4854 (N_4854,N_4296,N_4355);
or U4855 (N_4855,N_4093,N_4372);
and U4856 (N_4856,N_4145,N_4244);
xnor U4857 (N_4857,N_4120,N_4096);
xor U4858 (N_4858,N_4290,N_4287);
nor U4859 (N_4859,N_4391,N_4368);
and U4860 (N_4860,N_4044,N_4303);
nor U4861 (N_4861,N_4004,N_4334);
nor U4862 (N_4862,N_4451,N_4102);
nand U4863 (N_4863,N_4205,N_4071);
nand U4864 (N_4864,N_4153,N_4257);
or U4865 (N_4865,N_4081,N_4069);
or U4866 (N_4866,N_4184,N_4066);
nand U4867 (N_4867,N_4313,N_4097);
xor U4868 (N_4868,N_4008,N_4130);
xnor U4869 (N_4869,N_4394,N_4380);
or U4870 (N_4870,N_4131,N_4325);
and U4871 (N_4871,N_4247,N_4115);
nor U4872 (N_4872,N_4029,N_4100);
and U4873 (N_4873,N_4377,N_4471);
nand U4874 (N_4874,N_4148,N_4084);
and U4875 (N_4875,N_4276,N_4040);
nor U4876 (N_4876,N_4054,N_4349);
xor U4877 (N_4877,N_4398,N_4303);
xnor U4878 (N_4878,N_4076,N_4173);
nor U4879 (N_4879,N_4289,N_4487);
nor U4880 (N_4880,N_4304,N_4061);
nor U4881 (N_4881,N_4131,N_4480);
nor U4882 (N_4882,N_4457,N_4193);
nand U4883 (N_4883,N_4487,N_4181);
or U4884 (N_4884,N_4267,N_4385);
nor U4885 (N_4885,N_4125,N_4311);
xor U4886 (N_4886,N_4161,N_4447);
nand U4887 (N_4887,N_4287,N_4041);
xor U4888 (N_4888,N_4314,N_4386);
and U4889 (N_4889,N_4495,N_4059);
or U4890 (N_4890,N_4189,N_4029);
nand U4891 (N_4891,N_4086,N_4413);
nand U4892 (N_4892,N_4265,N_4195);
xnor U4893 (N_4893,N_4054,N_4216);
nor U4894 (N_4894,N_4399,N_4289);
xor U4895 (N_4895,N_4169,N_4117);
xor U4896 (N_4896,N_4193,N_4029);
or U4897 (N_4897,N_4259,N_4106);
and U4898 (N_4898,N_4396,N_4081);
nand U4899 (N_4899,N_4102,N_4175);
or U4900 (N_4900,N_4026,N_4204);
xor U4901 (N_4901,N_4381,N_4224);
and U4902 (N_4902,N_4087,N_4499);
nor U4903 (N_4903,N_4446,N_4059);
or U4904 (N_4904,N_4493,N_4371);
nand U4905 (N_4905,N_4422,N_4360);
or U4906 (N_4906,N_4072,N_4490);
and U4907 (N_4907,N_4229,N_4390);
nand U4908 (N_4908,N_4334,N_4018);
xor U4909 (N_4909,N_4048,N_4235);
or U4910 (N_4910,N_4497,N_4266);
nor U4911 (N_4911,N_4009,N_4010);
nor U4912 (N_4912,N_4205,N_4198);
or U4913 (N_4913,N_4333,N_4163);
nand U4914 (N_4914,N_4465,N_4129);
xor U4915 (N_4915,N_4076,N_4380);
nand U4916 (N_4916,N_4128,N_4315);
or U4917 (N_4917,N_4343,N_4252);
nor U4918 (N_4918,N_4371,N_4175);
or U4919 (N_4919,N_4300,N_4171);
xnor U4920 (N_4920,N_4375,N_4117);
nand U4921 (N_4921,N_4279,N_4148);
nand U4922 (N_4922,N_4253,N_4334);
xnor U4923 (N_4923,N_4226,N_4030);
and U4924 (N_4924,N_4328,N_4310);
and U4925 (N_4925,N_4025,N_4259);
or U4926 (N_4926,N_4264,N_4044);
nand U4927 (N_4927,N_4491,N_4230);
nor U4928 (N_4928,N_4103,N_4441);
or U4929 (N_4929,N_4098,N_4448);
or U4930 (N_4930,N_4472,N_4245);
nand U4931 (N_4931,N_4105,N_4425);
nor U4932 (N_4932,N_4164,N_4249);
or U4933 (N_4933,N_4051,N_4279);
or U4934 (N_4934,N_4410,N_4474);
or U4935 (N_4935,N_4244,N_4499);
xor U4936 (N_4936,N_4298,N_4378);
nor U4937 (N_4937,N_4232,N_4086);
and U4938 (N_4938,N_4187,N_4178);
or U4939 (N_4939,N_4290,N_4084);
nand U4940 (N_4940,N_4268,N_4053);
and U4941 (N_4941,N_4372,N_4134);
nand U4942 (N_4942,N_4426,N_4117);
or U4943 (N_4943,N_4320,N_4267);
nand U4944 (N_4944,N_4383,N_4430);
or U4945 (N_4945,N_4373,N_4130);
or U4946 (N_4946,N_4487,N_4238);
xor U4947 (N_4947,N_4128,N_4317);
nand U4948 (N_4948,N_4254,N_4084);
nand U4949 (N_4949,N_4290,N_4270);
xor U4950 (N_4950,N_4337,N_4292);
or U4951 (N_4951,N_4044,N_4309);
or U4952 (N_4952,N_4416,N_4009);
xor U4953 (N_4953,N_4321,N_4337);
nand U4954 (N_4954,N_4353,N_4059);
and U4955 (N_4955,N_4037,N_4112);
nor U4956 (N_4956,N_4074,N_4354);
nor U4957 (N_4957,N_4407,N_4117);
xor U4958 (N_4958,N_4126,N_4101);
xor U4959 (N_4959,N_4043,N_4315);
xnor U4960 (N_4960,N_4325,N_4315);
or U4961 (N_4961,N_4094,N_4128);
nor U4962 (N_4962,N_4116,N_4097);
nor U4963 (N_4963,N_4057,N_4421);
nand U4964 (N_4964,N_4195,N_4138);
and U4965 (N_4965,N_4248,N_4077);
and U4966 (N_4966,N_4050,N_4422);
nor U4967 (N_4967,N_4314,N_4402);
xnor U4968 (N_4968,N_4015,N_4283);
nand U4969 (N_4969,N_4398,N_4168);
or U4970 (N_4970,N_4353,N_4227);
and U4971 (N_4971,N_4211,N_4450);
nor U4972 (N_4972,N_4248,N_4445);
or U4973 (N_4973,N_4280,N_4245);
nor U4974 (N_4974,N_4061,N_4044);
nor U4975 (N_4975,N_4206,N_4390);
or U4976 (N_4976,N_4384,N_4295);
xnor U4977 (N_4977,N_4116,N_4346);
nand U4978 (N_4978,N_4335,N_4271);
and U4979 (N_4979,N_4477,N_4001);
or U4980 (N_4980,N_4110,N_4253);
and U4981 (N_4981,N_4096,N_4248);
xnor U4982 (N_4982,N_4413,N_4430);
xor U4983 (N_4983,N_4431,N_4016);
nor U4984 (N_4984,N_4353,N_4086);
or U4985 (N_4985,N_4132,N_4314);
and U4986 (N_4986,N_4253,N_4022);
and U4987 (N_4987,N_4086,N_4355);
xor U4988 (N_4988,N_4363,N_4445);
or U4989 (N_4989,N_4093,N_4291);
and U4990 (N_4990,N_4358,N_4030);
and U4991 (N_4991,N_4482,N_4362);
nor U4992 (N_4992,N_4047,N_4350);
nand U4993 (N_4993,N_4034,N_4429);
nand U4994 (N_4994,N_4447,N_4160);
nand U4995 (N_4995,N_4057,N_4024);
xor U4996 (N_4996,N_4289,N_4140);
and U4997 (N_4997,N_4497,N_4227);
nand U4998 (N_4998,N_4152,N_4240);
nor U4999 (N_4999,N_4315,N_4234);
or UO_0 (O_0,N_4853,N_4887);
xnor UO_1 (O_1,N_4602,N_4601);
nor UO_2 (O_2,N_4535,N_4678);
nor UO_3 (O_3,N_4850,N_4574);
nand UO_4 (O_4,N_4950,N_4583);
nand UO_5 (O_5,N_4855,N_4573);
nand UO_6 (O_6,N_4849,N_4835);
xnor UO_7 (O_7,N_4620,N_4954);
or UO_8 (O_8,N_4694,N_4629);
xor UO_9 (O_9,N_4671,N_4902);
nand UO_10 (O_10,N_4893,N_4507);
xnor UO_11 (O_11,N_4895,N_4816);
nor UO_12 (O_12,N_4987,N_4843);
and UO_13 (O_13,N_4964,N_4988);
nor UO_14 (O_14,N_4758,N_4656);
xor UO_15 (O_15,N_4767,N_4534);
nand UO_16 (O_16,N_4996,N_4551);
nand UO_17 (O_17,N_4817,N_4719);
xnor UO_18 (O_18,N_4599,N_4703);
and UO_19 (O_19,N_4742,N_4577);
nor UO_20 (O_20,N_4709,N_4775);
or UO_21 (O_21,N_4857,N_4516);
nand UO_22 (O_22,N_4727,N_4809);
xnor UO_23 (O_23,N_4808,N_4744);
nand UO_24 (O_24,N_4822,N_4874);
or UO_25 (O_25,N_4943,N_4862);
nand UO_26 (O_26,N_4899,N_4877);
or UO_27 (O_27,N_4777,N_4802);
or UO_28 (O_28,N_4746,N_4548);
and UO_29 (O_29,N_4803,N_4870);
and UO_30 (O_30,N_4965,N_4948);
nor UO_31 (O_31,N_4969,N_4793);
nand UO_32 (O_32,N_4991,N_4582);
nor UO_33 (O_33,N_4995,N_4910);
and UO_34 (O_34,N_4641,N_4831);
xnor UO_35 (O_35,N_4651,N_4913);
xnor UO_36 (O_36,N_4596,N_4543);
or UO_37 (O_37,N_4962,N_4649);
and UO_38 (O_38,N_4662,N_4556);
xor UO_39 (O_39,N_4718,N_4733);
nand UO_40 (O_40,N_4559,N_4976);
and UO_41 (O_41,N_4890,N_4994);
nand UO_42 (O_42,N_4522,N_4806);
xnor UO_43 (O_43,N_4810,N_4589);
or UO_44 (O_44,N_4904,N_4798);
and UO_45 (O_45,N_4712,N_4915);
nand UO_46 (O_46,N_4732,N_4882);
nand UO_47 (O_47,N_4673,N_4754);
nand UO_48 (O_48,N_4832,N_4771);
nand UO_49 (O_49,N_4552,N_4829);
nand UO_50 (O_50,N_4918,N_4685);
or UO_51 (O_51,N_4700,N_4539);
and UO_52 (O_52,N_4749,N_4664);
xnor UO_53 (O_53,N_4823,N_4927);
or UO_54 (O_54,N_4977,N_4581);
xor UO_55 (O_55,N_4753,N_4680);
nand UO_56 (O_56,N_4542,N_4963);
xor UO_57 (O_57,N_4997,N_4676);
xor UO_58 (O_58,N_4936,N_4917);
or UO_59 (O_59,N_4686,N_4847);
xnor UO_60 (O_60,N_4666,N_4909);
nand UO_61 (O_61,N_4748,N_4511);
xnor UO_62 (O_62,N_4869,N_4638);
and UO_63 (O_63,N_4520,N_4725);
nor UO_64 (O_64,N_4799,N_4716);
nor UO_65 (O_65,N_4762,N_4989);
nor UO_66 (O_66,N_4568,N_4929);
nand UO_67 (O_67,N_4947,N_4624);
xor UO_68 (O_68,N_4878,N_4875);
nor UO_69 (O_69,N_4760,N_4827);
xor UO_70 (O_70,N_4611,N_4856);
xor UO_71 (O_71,N_4805,N_4634);
or UO_72 (O_72,N_4858,N_4532);
nor UO_73 (O_73,N_4691,N_4618);
nor UO_74 (O_74,N_4888,N_4654);
and UO_75 (O_75,N_4971,N_4630);
nand UO_76 (O_76,N_4687,N_4896);
nand UO_77 (O_77,N_4665,N_4587);
and UO_78 (O_78,N_4941,N_4627);
or UO_79 (O_79,N_4935,N_4966);
or UO_80 (O_80,N_4828,N_4815);
and UO_81 (O_81,N_4790,N_4538);
and UO_82 (O_82,N_4603,N_4713);
nand UO_83 (O_83,N_4766,N_4578);
nor UO_84 (O_84,N_4923,N_4655);
xnor UO_85 (O_85,N_4648,N_4722);
xnor UO_86 (O_86,N_4545,N_4571);
xnor UO_87 (O_87,N_4698,N_4759);
nand UO_88 (O_88,N_4839,N_4872);
nand UO_89 (O_89,N_4864,N_4961);
nand UO_90 (O_90,N_4531,N_4841);
or UO_91 (O_91,N_4852,N_4619);
xor UO_92 (O_92,N_4821,N_4824);
nand UO_93 (O_93,N_4788,N_4905);
nand UO_94 (O_94,N_4863,N_4818);
and UO_95 (O_95,N_4998,N_4702);
nand UO_96 (O_96,N_4787,N_4885);
xnor UO_97 (O_97,N_4770,N_4633);
nor UO_98 (O_98,N_4682,N_4595);
nor UO_99 (O_99,N_4974,N_4932);
xnor UO_100 (O_100,N_4859,N_4924);
and UO_101 (O_101,N_4679,N_4768);
nor UO_102 (O_102,N_4621,N_4773);
and UO_103 (O_103,N_4940,N_4562);
or UO_104 (O_104,N_4729,N_4956);
nor UO_105 (O_105,N_4616,N_4873);
nor UO_106 (O_106,N_4957,N_4693);
nor UO_107 (O_107,N_4764,N_4763);
nand UO_108 (O_108,N_4782,N_4741);
nand UO_109 (O_109,N_4623,N_4681);
and UO_110 (O_110,N_4570,N_4944);
and UO_111 (O_111,N_4569,N_4731);
and UO_112 (O_112,N_4642,N_4993);
or UO_113 (O_113,N_4541,N_4837);
and UO_114 (O_114,N_4509,N_4846);
or UO_115 (O_115,N_4825,N_4550);
nand UO_116 (O_116,N_4786,N_4696);
nand UO_117 (O_117,N_4636,N_4505);
xor UO_118 (O_118,N_4921,N_4527);
nor UO_119 (O_119,N_4783,N_4978);
and UO_120 (O_120,N_4892,N_4500);
xor UO_121 (O_121,N_4625,N_4980);
nor UO_122 (O_122,N_4736,N_4591);
xnor UO_123 (O_123,N_4675,N_4617);
nand UO_124 (O_124,N_4914,N_4695);
xor UO_125 (O_125,N_4519,N_4529);
xor UO_126 (O_126,N_4811,N_4756);
nand UO_127 (O_127,N_4774,N_4813);
nor UO_128 (O_128,N_4706,N_4939);
nand UO_129 (O_129,N_4743,N_4726);
nand UO_130 (O_130,N_4765,N_4622);
xnor UO_131 (O_131,N_4842,N_4593);
xor UO_132 (O_132,N_4946,N_4639);
nor UO_133 (O_133,N_4883,N_4643);
or UO_134 (O_134,N_4670,N_4886);
or UO_135 (O_135,N_4610,N_4645);
and UO_136 (O_136,N_4903,N_4724);
and UO_137 (O_137,N_4606,N_4515);
or UO_138 (O_138,N_4544,N_4644);
or UO_139 (O_139,N_4735,N_4547);
xor UO_140 (O_140,N_4584,N_4588);
xor UO_141 (O_141,N_4985,N_4684);
and UO_142 (O_142,N_4692,N_4851);
or UO_143 (O_143,N_4826,N_4973);
nand UO_144 (O_144,N_4563,N_4667);
xor UO_145 (O_145,N_4953,N_4751);
and UO_146 (O_146,N_4710,N_4845);
and UO_147 (O_147,N_4608,N_4501);
or UO_148 (O_148,N_4558,N_4897);
nor UO_149 (O_149,N_4580,N_4830);
or UO_150 (O_150,N_4757,N_4517);
or UO_151 (O_151,N_4592,N_4931);
and UO_152 (O_152,N_4502,N_4794);
or UO_153 (O_153,N_4715,N_4609);
or UO_154 (O_154,N_4785,N_4518);
nand UO_155 (O_155,N_4540,N_4983);
and UO_156 (O_156,N_4972,N_4945);
xnor UO_157 (O_157,N_4714,N_4881);
and UO_158 (O_158,N_4848,N_4791);
and UO_159 (O_159,N_4708,N_4912);
and UO_160 (O_160,N_4711,N_4510);
nor UO_161 (O_161,N_4553,N_4769);
nor UO_162 (O_162,N_4796,N_4546);
xor UO_163 (O_163,N_4807,N_4614);
xnor UO_164 (O_164,N_4720,N_4697);
nor UO_165 (O_165,N_4674,N_4958);
nor UO_166 (O_166,N_4524,N_4612);
nand UO_167 (O_167,N_4707,N_4779);
nor UO_168 (O_168,N_4761,N_4840);
xnor UO_169 (O_169,N_4801,N_4797);
or UO_170 (O_170,N_4868,N_4730);
xor UO_171 (O_171,N_4926,N_4672);
and UO_172 (O_172,N_4661,N_4683);
and UO_173 (O_173,N_4567,N_4523);
nand UO_174 (O_174,N_4631,N_4740);
and UO_175 (O_175,N_4804,N_4860);
xnor UO_176 (O_176,N_4723,N_4626);
nand UO_177 (O_177,N_4585,N_4663);
nor UO_178 (O_178,N_4704,N_4838);
and UO_179 (O_179,N_4861,N_4737);
nand UO_180 (O_180,N_4986,N_4615);
and UO_181 (O_181,N_4504,N_4554);
xor UO_182 (O_182,N_4508,N_4814);
or UO_183 (O_183,N_4772,N_4920);
nand UO_184 (O_184,N_4635,N_4594);
nand UO_185 (O_185,N_4982,N_4613);
nor UO_186 (O_186,N_4984,N_4652);
or UO_187 (O_187,N_4820,N_4833);
and UO_188 (O_188,N_4901,N_4650);
nand UO_189 (O_189,N_4975,N_4889);
nor UO_190 (O_190,N_4549,N_4640);
and UO_191 (O_191,N_4521,N_4659);
xnor UO_192 (O_192,N_4911,N_4530);
and UO_193 (O_193,N_4906,N_4955);
nand UO_194 (O_194,N_4526,N_4705);
or UO_195 (O_195,N_4503,N_4728);
nand UO_196 (O_196,N_4647,N_4560);
and UO_197 (O_197,N_4590,N_4628);
and UO_198 (O_198,N_4968,N_4572);
or UO_199 (O_199,N_4514,N_4689);
nand UO_200 (O_200,N_4999,N_4992);
nand UO_201 (O_201,N_4668,N_4699);
or UO_202 (O_202,N_4959,N_4506);
or UO_203 (O_203,N_4891,N_4739);
xor UO_204 (O_204,N_4836,N_4653);
and UO_205 (O_205,N_4928,N_4938);
nor UO_206 (O_206,N_4967,N_4717);
or UO_207 (O_207,N_4669,N_4907);
or UO_208 (O_208,N_4930,N_4605);
nor UO_209 (O_209,N_4747,N_4776);
xor UO_210 (O_210,N_4800,N_4933);
and UO_211 (O_211,N_4646,N_4604);
nand UO_212 (O_212,N_4781,N_4513);
xor UO_213 (O_213,N_4866,N_4898);
nor UO_214 (O_214,N_4784,N_4934);
and UO_215 (O_215,N_4894,N_4925);
or UO_216 (O_216,N_4949,N_4750);
nor UO_217 (O_217,N_4701,N_4755);
xnor UO_218 (O_218,N_4575,N_4792);
or UO_219 (O_219,N_4937,N_4512);
nor UO_220 (O_220,N_4780,N_4981);
and UO_221 (O_221,N_4844,N_4867);
xor UO_222 (O_222,N_4865,N_4597);
nand UO_223 (O_223,N_4880,N_4525);
nor UO_224 (O_224,N_4564,N_4970);
xor UO_225 (O_225,N_4637,N_4555);
nor UO_226 (O_226,N_4778,N_4677);
nor UO_227 (O_227,N_4900,N_4952);
xnor UO_228 (O_228,N_4879,N_4795);
xor UO_229 (O_229,N_4557,N_4688);
xnor UO_230 (O_230,N_4960,N_4942);
nor UO_231 (O_231,N_4979,N_4658);
xnor UO_232 (O_232,N_4632,N_4690);
or UO_233 (O_233,N_4876,N_4536);
and UO_234 (O_234,N_4752,N_4565);
nand UO_235 (O_235,N_4908,N_4579);
xor UO_236 (O_236,N_4834,N_4598);
and UO_237 (O_237,N_4789,N_4586);
xor UO_238 (O_238,N_4819,N_4561);
or UO_239 (O_239,N_4951,N_4738);
nor UO_240 (O_240,N_4576,N_4854);
and UO_241 (O_241,N_4537,N_4660);
and UO_242 (O_242,N_4528,N_4600);
xnor UO_243 (O_243,N_4657,N_4919);
or UO_244 (O_244,N_4533,N_4871);
and UO_245 (O_245,N_4566,N_4922);
or UO_246 (O_246,N_4990,N_4734);
nand UO_247 (O_247,N_4607,N_4721);
or UO_248 (O_248,N_4884,N_4812);
nor UO_249 (O_249,N_4745,N_4916);
and UO_250 (O_250,N_4540,N_4647);
nor UO_251 (O_251,N_4569,N_4788);
xnor UO_252 (O_252,N_4875,N_4691);
nand UO_253 (O_253,N_4744,N_4582);
or UO_254 (O_254,N_4809,N_4792);
nand UO_255 (O_255,N_4680,N_4593);
nand UO_256 (O_256,N_4587,N_4605);
and UO_257 (O_257,N_4877,N_4799);
or UO_258 (O_258,N_4775,N_4516);
nor UO_259 (O_259,N_4891,N_4736);
and UO_260 (O_260,N_4840,N_4996);
and UO_261 (O_261,N_4604,N_4631);
xor UO_262 (O_262,N_4757,N_4940);
nor UO_263 (O_263,N_4858,N_4999);
xor UO_264 (O_264,N_4987,N_4616);
and UO_265 (O_265,N_4778,N_4947);
and UO_266 (O_266,N_4999,N_4731);
nor UO_267 (O_267,N_4514,N_4747);
and UO_268 (O_268,N_4978,N_4540);
or UO_269 (O_269,N_4776,N_4933);
xor UO_270 (O_270,N_4542,N_4589);
or UO_271 (O_271,N_4711,N_4643);
nand UO_272 (O_272,N_4909,N_4615);
nand UO_273 (O_273,N_4709,N_4505);
nor UO_274 (O_274,N_4627,N_4695);
nand UO_275 (O_275,N_4898,N_4869);
or UO_276 (O_276,N_4979,N_4967);
xor UO_277 (O_277,N_4720,N_4700);
nand UO_278 (O_278,N_4569,N_4781);
nand UO_279 (O_279,N_4773,N_4695);
or UO_280 (O_280,N_4502,N_4958);
and UO_281 (O_281,N_4783,N_4523);
and UO_282 (O_282,N_4595,N_4753);
nor UO_283 (O_283,N_4620,N_4614);
or UO_284 (O_284,N_4672,N_4836);
xor UO_285 (O_285,N_4504,N_4737);
xnor UO_286 (O_286,N_4920,N_4805);
nand UO_287 (O_287,N_4651,N_4764);
and UO_288 (O_288,N_4949,N_4735);
and UO_289 (O_289,N_4648,N_4525);
and UO_290 (O_290,N_4936,N_4683);
xor UO_291 (O_291,N_4633,N_4530);
or UO_292 (O_292,N_4861,N_4702);
or UO_293 (O_293,N_4528,N_4814);
or UO_294 (O_294,N_4900,N_4529);
and UO_295 (O_295,N_4991,N_4897);
nand UO_296 (O_296,N_4528,N_4793);
xor UO_297 (O_297,N_4766,N_4591);
nand UO_298 (O_298,N_4502,N_4597);
nor UO_299 (O_299,N_4951,N_4757);
nand UO_300 (O_300,N_4854,N_4585);
and UO_301 (O_301,N_4725,N_4880);
and UO_302 (O_302,N_4623,N_4852);
nand UO_303 (O_303,N_4878,N_4978);
nor UO_304 (O_304,N_4690,N_4749);
and UO_305 (O_305,N_4857,N_4882);
xnor UO_306 (O_306,N_4734,N_4611);
nor UO_307 (O_307,N_4519,N_4986);
nand UO_308 (O_308,N_4573,N_4851);
nand UO_309 (O_309,N_4838,N_4527);
nor UO_310 (O_310,N_4977,N_4667);
or UO_311 (O_311,N_4931,N_4729);
or UO_312 (O_312,N_4940,N_4702);
and UO_313 (O_313,N_4625,N_4515);
and UO_314 (O_314,N_4528,N_4757);
or UO_315 (O_315,N_4871,N_4765);
or UO_316 (O_316,N_4863,N_4974);
nand UO_317 (O_317,N_4951,N_4901);
xnor UO_318 (O_318,N_4880,N_4979);
nor UO_319 (O_319,N_4528,N_4724);
or UO_320 (O_320,N_4676,N_4736);
and UO_321 (O_321,N_4838,N_4593);
xnor UO_322 (O_322,N_4576,N_4572);
and UO_323 (O_323,N_4880,N_4935);
xnor UO_324 (O_324,N_4516,N_4818);
and UO_325 (O_325,N_4597,N_4520);
or UO_326 (O_326,N_4951,N_4810);
and UO_327 (O_327,N_4519,N_4656);
xnor UO_328 (O_328,N_4633,N_4660);
nand UO_329 (O_329,N_4910,N_4571);
xnor UO_330 (O_330,N_4678,N_4684);
and UO_331 (O_331,N_4595,N_4738);
nor UO_332 (O_332,N_4905,N_4902);
and UO_333 (O_333,N_4807,N_4860);
xor UO_334 (O_334,N_4656,N_4713);
or UO_335 (O_335,N_4925,N_4582);
nand UO_336 (O_336,N_4629,N_4946);
nor UO_337 (O_337,N_4646,N_4866);
nand UO_338 (O_338,N_4817,N_4839);
nor UO_339 (O_339,N_4513,N_4692);
nand UO_340 (O_340,N_4765,N_4743);
xor UO_341 (O_341,N_4858,N_4957);
xnor UO_342 (O_342,N_4604,N_4560);
nand UO_343 (O_343,N_4707,N_4869);
nor UO_344 (O_344,N_4905,N_4618);
and UO_345 (O_345,N_4947,N_4997);
nand UO_346 (O_346,N_4913,N_4614);
xnor UO_347 (O_347,N_4910,N_4993);
or UO_348 (O_348,N_4580,N_4677);
nand UO_349 (O_349,N_4520,N_4872);
xor UO_350 (O_350,N_4781,N_4599);
nand UO_351 (O_351,N_4580,N_4813);
and UO_352 (O_352,N_4715,N_4970);
nor UO_353 (O_353,N_4640,N_4892);
nand UO_354 (O_354,N_4709,N_4958);
or UO_355 (O_355,N_4741,N_4970);
xor UO_356 (O_356,N_4595,N_4711);
or UO_357 (O_357,N_4866,N_4869);
xor UO_358 (O_358,N_4600,N_4672);
or UO_359 (O_359,N_4850,N_4949);
or UO_360 (O_360,N_4840,N_4740);
nor UO_361 (O_361,N_4778,N_4946);
xnor UO_362 (O_362,N_4951,N_4794);
xnor UO_363 (O_363,N_4887,N_4744);
nor UO_364 (O_364,N_4671,N_4667);
xnor UO_365 (O_365,N_4940,N_4597);
xnor UO_366 (O_366,N_4509,N_4616);
nand UO_367 (O_367,N_4932,N_4756);
and UO_368 (O_368,N_4938,N_4891);
or UO_369 (O_369,N_4787,N_4657);
xor UO_370 (O_370,N_4616,N_4833);
xor UO_371 (O_371,N_4906,N_4898);
nor UO_372 (O_372,N_4526,N_4897);
nand UO_373 (O_373,N_4527,N_4544);
xnor UO_374 (O_374,N_4859,N_4709);
xor UO_375 (O_375,N_4786,N_4668);
nand UO_376 (O_376,N_4967,N_4877);
and UO_377 (O_377,N_4720,N_4681);
nand UO_378 (O_378,N_4881,N_4585);
or UO_379 (O_379,N_4645,N_4865);
nand UO_380 (O_380,N_4676,N_4884);
nor UO_381 (O_381,N_4917,N_4850);
and UO_382 (O_382,N_4573,N_4516);
nand UO_383 (O_383,N_4519,N_4546);
or UO_384 (O_384,N_4607,N_4895);
nor UO_385 (O_385,N_4838,N_4904);
or UO_386 (O_386,N_4772,N_4784);
nor UO_387 (O_387,N_4503,N_4953);
nor UO_388 (O_388,N_4600,N_4756);
nand UO_389 (O_389,N_4779,N_4678);
xnor UO_390 (O_390,N_4929,N_4883);
xnor UO_391 (O_391,N_4606,N_4503);
xnor UO_392 (O_392,N_4735,N_4505);
and UO_393 (O_393,N_4506,N_4918);
nor UO_394 (O_394,N_4997,N_4875);
nor UO_395 (O_395,N_4654,N_4616);
and UO_396 (O_396,N_4888,N_4892);
nor UO_397 (O_397,N_4942,N_4581);
nand UO_398 (O_398,N_4752,N_4874);
and UO_399 (O_399,N_4840,N_4598);
xnor UO_400 (O_400,N_4704,N_4707);
nor UO_401 (O_401,N_4622,N_4727);
and UO_402 (O_402,N_4975,N_4539);
or UO_403 (O_403,N_4748,N_4796);
nand UO_404 (O_404,N_4973,N_4687);
nand UO_405 (O_405,N_4711,N_4566);
xnor UO_406 (O_406,N_4590,N_4769);
xor UO_407 (O_407,N_4505,N_4655);
nand UO_408 (O_408,N_4682,N_4711);
or UO_409 (O_409,N_4736,N_4713);
and UO_410 (O_410,N_4766,N_4864);
nand UO_411 (O_411,N_4773,N_4853);
xor UO_412 (O_412,N_4864,N_4510);
or UO_413 (O_413,N_4547,N_4604);
nand UO_414 (O_414,N_4665,N_4764);
nor UO_415 (O_415,N_4834,N_4654);
and UO_416 (O_416,N_4543,N_4662);
or UO_417 (O_417,N_4740,N_4802);
nor UO_418 (O_418,N_4901,N_4700);
or UO_419 (O_419,N_4543,N_4732);
and UO_420 (O_420,N_4567,N_4606);
or UO_421 (O_421,N_4765,N_4712);
xnor UO_422 (O_422,N_4727,N_4623);
xnor UO_423 (O_423,N_4887,N_4627);
xor UO_424 (O_424,N_4897,N_4890);
or UO_425 (O_425,N_4733,N_4854);
nand UO_426 (O_426,N_4575,N_4713);
or UO_427 (O_427,N_4739,N_4984);
xnor UO_428 (O_428,N_4889,N_4708);
or UO_429 (O_429,N_4715,N_4506);
nand UO_430 (O_430,N_4545,N_4634);
or UO_431 (O_431,N_4889,N_4569);
xor UO_432 (O_432,N_4693,N_4840);
and UO_433 (O_433,N_4545,N_4626);
and UO_434 (O_434,N_4823,N_4861);
or UO_435 (O_435,N_4681,N_4974);
or UO_436 (O_436,N_4816,N_4953);
nand UO_437 (O_437,N_4820,N_4616);
nor UO_438 (O_438,N_4814,N_4647);
xor UO_439 (O_439,N_4956,N_4548);
nor UO_440 (O_440,N_4884,N_4723);
or UO_441 (O_441,N_4879,N_4532);
and UO_442 (O_442,N_4745,N_4669);
and UO_443 (O_443,N_4780,N_4699);
xnor UO_444 (O_444,N_4864,N_4954);
or UO_445 (O_445,N_4760,N_4928);
nand UO_446 (O_446,N_4985,N_4613);
and UO_447 (O_447,N_4970,N_4559);
and UO_448 (O_448,N_4589,N_4837);
nand UO_449 (O_449,N_4608,N_4550);
xor UO_450 (O_450,N_4630,N_4524);
or UO_451 (O_451,N_4714,N_4522);
nor UO_452 (O_452,N_4603,N_4824);
and UO_453 (O_453,N_4804,N_4686);
xnor UO_454 (O_454,N_4670,N_4956);
or UO_455 (O_455,N_4897,N_4671);
nand UO_456 (O_456,N_4755,N_4910);
xor UO_457 (O_457,N_4861,N_4589);
or UO_458 (O_458,N_4623,N_4788);
nand UO_459 (O_459,N_4685,N_4689);
xnor UO_460 (O_460,N_4534,N_4728);
and UO_461 (O_461,N_4682,N_4920);
xor UO_462 (O_462,N_4965,N_4545);
nor UO_463 (O_463,N_4699,N_4620);
and UO_464 (O_464,N_4626,N_4738);
and UO_465 (O_465,N_4678,N_4984);
xor UO_466 (O_466,N_4767,N_4623);
nor UO_467 (O_467,N_4773,N_4569);
xor UO_468 (O_468,N_4638,N_4946);
or UO_469 (O_469,N_4763,N_4868);
or UO_470 (O_470,N_4852,N_4703);
or UO_471 (O_471,N_4994,N_4677);
and UO_472 (O_472,N_4530,N_4916);
xnor UO_473 (O_473,N_4771,N_4553);
and UO_474 (O_474,N_4980,N_4714);
xnor UO_475 (O_475,N_4832,N_4550);
xnor UO_476 (O_476,N_4741,N_4566);
nand UO_477 (O_477,N_4514,N_4809);
xnor UO_478 (O_478,N_4591,N_4581);
nor UO_479 (O_479,N_4693,N_4536);
or UO_480 (O_480,N_4782,N_4784);
and UO_481 (O_481,N_4944,N_4500);
nor UO_482 (O_482,N_4597,N_4602);
and UO_483 (O_483,N_4916,N_4520);
or UO_484 (O_484,N_4993,N_4983);
and UO_485 (O_485,N_4652,N_4923);
nor UO_486 (O_486,N_4752,N_4962);
or UO_487 (O_487,N_4956,N_4810);
or UO_488 (O_488,N_4922,N_4963);
xnor UO_489 (O_489,N_4847,N_4818);
nand UO_490 (O_490,N_4970,N_4762);
nand UO_491 (O_491,N_4506,N_4602);
nor UO_492 (O_492,N_4935,N_4916);
nor UO_493 (O_493,N_4901,N_4921);
xnor UO_494 (O_494,N_4985,N_4801);
nand UO_495 (O_495,N_4695,N_4815);
or UO_496 (O_496,N_4711,N_4692);
or UO_497 (O_497,N_4818,N_4751);
or UO_498 (O_498,N_4812,N_4720);
and UO_499 (O_499,N_4802,N_4961);
nor UO_500 (O_500,N_4662,N_4613);
nor UO_501 (O_501,N_4857,N_4887);
or UO_502 (O_502,N_4828,N_4662);
nor UO_503 (O_503,N_4980,N_4569);
xnor UO_504 (O_504,N_4574,N_4826);
xor UO_505 (O_505,N_4979,N_4857);
nand UO_506 (O_506,N_4583,N_4725);
nor UO_507 (O_507,N_4801,N_4947);
nor UO_508 (O_508,N_4839,N_4544);
or UO_509 (O_509,N_4593,N_4630);
xnor UO_510 (O_510,N_4888,N_4881);
nand UO_511 (O_511,N_4645,N_4758);
and UO_512 (O_512,N_4686,N_4931);
nor UO_513 (O_513,N_4742,N_4811);
and UO_514 (O_514,N_4619,N_4716);
or UO_515 (O_515,N_4819,N_4796);
nor UO_516 (O_516,N_4771,N_4829);
xnor UO_517 (O_517,N_4784,N_4949);
and UO_518 (O_518,N_4910,N_4989);
nand UO_519 (O_519,N_4935,N_4767);
nor UO_520 (O_520,N_4776,N_4553);
and UO_521 (O_521,N_4982,N_4781);
and UO_522 (O_522,N_4575,N_4927);
and UO_523 (O_523,N_4944,N_4614);
nor UO_524 (O_524,N_4519,N_4750);
nand UO_525 (O_525,N_4999,N_4662);
and UO_526 (O_526,N_4935,N_4641);
or UO_527 (O_527,N_4607,N_4692);
nand UO_528 (O_528,N_4863,N_4887);
nor UO_529 (O_529,N_4716,N_4782);
nor UO_530 (O_530,N_4821,N_4888);
or UO_531 (O_531,N_4844,N_4719);
xnor UO_532 (O_532,N_4873,N_4904);
xnor UO_533 (O_533,N_4654,N_4718);
nand UO_534 (O_534,N_4847,N_4727);
or UO_535 (O_535,N_4667,N_4878);
xor UO_536 (O_536,N_4674,N_4669);
or UO_537 (O_537,N_4997,N_4894);
and UO_538 (O_538,N_4904,N_4846);
xnor UO_539 (O_539,N_4618,N_4548);
nor UO_540 (O_540,N_4790,N_4540);
or UO_541 (O_541,N_4686,N_4873);
nand UO_542 (O_542,N_4993,N_4913);
xnor UO_543 (O_543,N_4746,N_4831);
xor UO_544 (O_544,N_4558,N_4809);
nand UO_545 (O_545,N_4542,N_4796);
xnor UO_546 (O_546,N_4548,N_4555);
xnor UO_547 (O_547,N_4514,N_4864);
nand UO_548 (O_548,N_4994,N_4723);
or UO_549 (O_549,N_4545,N_4800);
or UO_550 (O_550,N_4905,N_4625);
or UO_551 (O_551,N_4808,N_4954);
nor UO_552 (O_552,N_4664,N_4561);
and UO_553 (O_553,N_4969,N_4702);
nand UO_554 (O_554,N_4628,N_4612);
nor UO_555 (O_555,N_4531,N_4517);
nand UO_556 (O_556,N_4543,N_4518);
or UO_557 (O_557,N_4620,N_4992);
and UO_558 (O_558,N_4880,N_4515);
nand UO_559 (O_559,N_4546,N_4753);
and UO_560 (O_560,N_4935,N_4938);
nand UO_561 (O_561,N_4613,N_4505);
or UO_562 (O_562,N_4932,N_4577);
xor UO_563 (O_563,N_4729,N_4786);
nand UO_564 (O_564,N_4578,N_4707);
nor UO_565 (O_565,N_4575,N_4635);
nor UO_566 (O_566,N_4987,N_4762);
xor UO_567 (O_567,N_4628,N_4665);
xnor UO_568 (O_568,N_4693,N_4588);
or UO_569 (O_569,N_4873,N_4832);
nor UO_570 (O_570,N_4868,N_4528);
and UO_571 (O_571,N_4911,N_4658);
nand UO_572 (O_572,N_4715,N_4713);
nor UO_573 (O_573,N_4949,N_4939);
nand UO_574 (O_574,N_4527,N_4926);
or UO_575 (O_575,N_4600,N_4984);
nor UO_576 (O_576,N_4726,N_4821);
nor UO_577 (O_577,N_4520,N_4841);
nand UO_578 (O_578,N_4973,N_4907);
nor UO_579 (O_579,N_4901,N_4933);
or UO_580 (O_580,N_4899,N_4950);
nor UO_581 (O_581,N_4788,N_4690);
or UO_582 (O_582,N_4712,N_4598);
and UO_583 (O_583,N_4895,N_4578);
and UO_584 (O_584,N_4837,N_4908);
and UO_585 (O_585,N_4529,N_4516);
nand UO_586 (O_586,N_4715,N_4957);
xor UO_587 (O_587,N_4900,N_4741);
nor UO_588 (O_588,N_4962,N_4689);
nor UO_589 (O_589,N_4587,N_4785);
nor UO_590 (O_590,N_4723,N_4649);
nand UO_591 (O_591,N_4973,N_4981);
nand UO_592 (O_592,N_4556,N_4641);
or UO_593 (O_593,N_4993,N_4848);
nand UO_594 (O_594,N_4960,N_4850);
xor UO_595 (O_595,N_4853,N_4698);
xor UO_596 (O_596,N_4811,N_4840);
and UO_597 (O_597,N_4615,N_4625);
or UO_598 (O_598,N_4818,N_4990);
or UO_599 (O_599,N_4796,N_4526);
nor UO_600 (O_600,N_4589,N_4852);
nor UO_601 (O_601,N_4545,N_4769);
or UO_602 (O_602,N_4512,N_4545);
and UO_603 (O_603,N_4982,N_4558);
nor UO_604 (O_604,N_4727,N_4522);
nand UO_605 (O_605,N_4689,N_4619);
or UO_606 (O_606,N_4872,N_4681);
xor UO_607 (O_607,N_4958,N_4518);
nand UO_608 (O_608,N_4834,N_4570);
nand UO_609 (O_609,N_4547,N_4558);
nand UO_610 (O_610,N_4545,N_4854);
or UO_611 (O_611,N_4885,N_4589);
and UO_612 (O_612,N_4895,N_4604);
nand UO_613 (O_613,N_4763,N_4713);
and UO_614 (O_614,N_4518,N_4981);
nand UO_615 (O_615,N_4503,N_4897);
and UO_616 (O_616,N_4539,N_4834);
nand UO_617 (O_617,N_4620,N_4672);
or UO_618 (O_618,N_4678,N_4914);
nand UO_619 (O_619,N_4588,N_4847);
nand UO_620 (O_620,N_4511,N_4974);
xnor UO_621 (O_621,N_4868,N_4971);
xnor UO_622 (O_622,N_4873,N_4975);
nor UO_623 (O_623,N_4577,N_4653);
or UO_624 (O_624,N_4810,N_4808);
nor UO_625 (O_625,N_4887,N_4534);
nand UO_626 (O_626,N_4519,N_4874);
xnor UO_627 (O_627,N_4642,N_4740);
or UO_628 (O_628,N_4704,N_4938);
xnor UO_629 (O_629,N_4846,N_4789);
xnor UO_630 (O_630,N_4872,N_4852);
or UO_631 (O_631,N_4927,N_4748);
nor UO_632 (O_632,N_4685,N_4659);
nand UO_633 (O_633,N_4942,N_4506);
or UO_634 (O_634,N_4819,N_4916);
or UO_635 (O_635,N_4990,N_4882);
nand UO_636 (O_636,N_4608,N_4643);
nor UO_637 (O_637,N_4559,N_4878);
nor UO_638 (O_638,N_4767,N_4692);
nor UO_639 (O_639,N_4707,N_4618);
xor UO_640 (O_640,N_4894,N_4927);
and UO_641 (O_641,N_4625,N_4651);
nor UO_642 (O_642,N_4610,N_4964);
nor UO_643 (O_643,N_4679,N_4996);
or UO_644 (O_644,N_4656,N_4934);
and UO_645 (O_645,N_4909,N_4699);
nand UO_646 (O_646,N_4995,N_4641);
xnor UO_647 (O_647,N_4684,N_4844);
nand UO_648 (O_648,N_4670,N_4687);
nand UO_649 (O_649,N_4612,N_4615);
or UO_650 (O_650,N_4911,N_4734);
nor UO_651 (O_651,N_4869,N_4527);
xor UO_652 (O_652,N_4671,N_4925);
and UO_653 (O_653,N_4861,N_4758);
xor UO_654 (O_654,N_4895,N_4884);
nand UO_655 (O_655,N_4787,N_4977);
nand UO_656 (O_656,N_4751,N_4557);
xnor UO_657 (O_657,N_4555,N_4807);
and UO_658 (O_658,N_4567,N_4592);
xnor UO_659 (O_659,N_4771,N_4654);
nand UO_660 (O_660,N_4890,N_4996);
and UO_661 (O_661,N_4797,N_4536);
and UO_662 (O_662,N_4576,N_4955);
nor UO_663 (O_663,N_4540,N_4997);
xor UO_664 (O_664,N_4989,N_4674);
and UO_665 (O_665,N_4848,N_4938);
and UO_666 (O_666,N_4509,N_4864);
or UO_667 (O_667,N_4959,N_4872);
and UO_668 (O_668,N_4851,N_4705);
and UO_669 (O_669,N_4998,N_4860);
xor UO_670 (O_670,N_4509,N_4932);
or UO_671 (O_671,N_4992,N_4687);
nand UO_672 (O_672,N_4919,N_4766);
nor UO_673 (O_673,N_4769,N_4827);
xor UO_674 (O_674,N_4550,N_4701);
and UO_675 (O_675,N_4739,N_4953);
or UO_676 (O_676,N_4796,N_4588);
and UO_677 (O_677,N_4890,N_4900);
nor UO_678 (O_678,N_4795,N_4705);
xor UO_679 (O_679,N_4669,N_4719);
nor UO_680 (O_680,N_4635,N_4988);
xnor UO_681 (O_681,N_4903,N_4934);
xor UO_682 (O_682,N_4669,N_4805);
xnor UO_683 (O_683,N_4563,N_4539);
or UO_684 (O_684,N_4885,N_4611);
xnor UO_685 (O_685,N_4701,N_4521);
xor UO_686 (O_686,N_4777,N_4502);
nand UO_687 (O_687,N_4997,N_4718);
and UO_688 (O_688,N_4877,N_4624);
and UO_689 (O_689,N_4809,N_4922);
or UO_690 (O_690,N_4703,N_4953);
and UO_691 (O_691,N_4860,N_4828);
nand UO_692 (O_692,N_4940,N_4541);
nor UO_693 (O_693,N_4808,N_4631);
and UO_694 (O_694,N_4841,N_4655);
xnor UO_695 (O_695,N_4918,N_4938);
xnor UO_696 (O_696,N_4613,N_4739);
xnor UO_697 (O_697,N_4524,N_4842);
and UO_698 (O_698,N_4608,N_4797);
or UO_699 (O_699,N_4620,N_4671);
or UO_700 (O_700,N_4738,N_4814);
or UO_701 (O_701,N_4739,N_4732);
or UO_702 (O_702,N_4666,N_4824);
or UO_703 (O_703,N_4873,N_4798);
nor UO_704 (O_704,N_4968,N_4971);
nand UO_705 (O_705,N_4511,N_4623);
or UO_706 (O_706,N_4876,N_4769);
nor UO_707 (O_707,N_4642,N_4641);
and UO_708 (O_708,N_4828,N_4791);
nand UO_709 (O_709,N_4576,N_4825);
nor UO_710 (O_710,N_4804,N_4857);
and UO_711 (O_711,N_4776,N_4843);
xor UO_712 (O_712,N_4743,N_4860);
nand UO_713 (O_713,N_4942,N_4918);
and UO_714 (O_714,N_4919,N_4525);
nor UO_715 (O_715,N_4774,N_4653);
xor UO_716 (O_716,N_4994,N_4797);
or UO_717 (O_717,N_4931,N_4785);
and UO_718 (O_718,N_4614,N_4794);
nor UO_719 (O_719,N_4995,N_4895);
xnor UO_720 (O_720,N_4567,N_4950);
xor UO_721 (O_721,N_4516,N_4537);
or UO_722 (O_722,N_4932,N_4596);
and UO_723 (O_723,N_4864,N_4702);
xor UO_724 (O_724,N_4575,N_4836);
or UO_725 (O_725,N_4669,N_4532);
or UO_726 (O_726,N_4774,N_4621);
nand UO_727 (O_727,N_4703,N_4908);
nand UO_728 (O_728,N_4999,N_4723);
nand UO_729 (O_729,N_4607,N_4540);
nor UO_730 (O_730,N_4752,N_4620);
nand UO_731 (O_731,N_4669,N_4883);
or UO_732 (O_732,N_4815,N_4953);
xnor UO_733 (O_733,N_4572,N_4861);
nor UO_734 (O_734,N_4533,N_4998);
or UO_735 (O_735,N_4989,N_4912);
nand UO_736 (O_736,N_4863,N_4864);
xor UO_737 (O_737,N_4898,N_4723);
xnor UO_738 (O_738,N_4544,N_4871);
and UO_739 (O_739,N_4865,N_4570);
or UO_740 (O_740,N_4818,N_4528);
and UO_741 (O_741,N_4564,N_4777);
xor UO_742 (O_742,N_4767,N_4875);
or UO_743 (O_743,N_4671,N_4960);
nor UO_744 (O_744,N_4946,N_4650);
nand UO_745 (O_745,N_4607,N_4739);
and UO_746 (O_746,N_4845,N_4778);
nand UO_747 (O_747,N_4977,N_4674);
xnor UO_748 (O_748,N_4921,N_4964);
and UO_749 (O_749,N_4708,N_4879);
nand UO_750 (O_750,N_4735,N_4675);
and UO_751 (O_751,N_4719,N_4604);
nor UO_752 (O_752,N_4636,N_4514);
or UO_753 (O_753,N_4863,N_4938);
and UO_754 (O_754,N_4554,N_4680);
and UO_755 (O_755,N_4912,N_4669);
or UO_756 (O_756,N_4570,N_4915);
nor UO_757 (O_757,N_4685,N_4823);
nand UO_758 (O_758,N_4767,N_4913);
xor UO_759 (O_759,N_4885,N_4571);
nand UO_760 (O_760,N_4889,N_4944);
nor UO_761 (O_761,N_4661,N_4783);
xor UO_762 (O_762,N_4596,N_4980);
nand UO_763 (O_763,N_4620,N_4691);
and UO_764 (O_764,N_4712,N_4725);
nand UO_765 (O_765,N_4754,N_4991);
nor UO_766 (O_766,N_4669,N_4551);
nand UO_767 (O_767,N_4610,N_4640);
nand UO_768 (O_768,N_4950,N_4761);
xor UO_769 (O_769,N_4536,N_4520);
nand UO_770 (O_770,N_4682,N_4961);
nand UO_771 (O_771,N_4501,N_4563);
nand UO_772 (O_772,N_4615,N_4719);
nor UO_773 (O_773,N_4962,N_4958);
nand UO_774 (O_774,N_4656,N_4779);
xnor UO_775 (O_775,N_4735,N_4794);
or UO_776 (O_776,N_4636,N_4658);
or UO_777 (O_777,N_4565,N_4726);
nand UO_778 (O_778,N_4667,N_4568);
and UO_779 (O_779,N_4678,N_4810);
or UO_780 (O_780,N_4644,N_4874);
or UO_781 (O_781,N_4700,N_4535);
or UO_782 (O_782,N_4890,N_4723);
nand UO_783 (O_783,N_4957,N_4649);
and UO_784 (O_784,N_4960,N_4808);
nand UO_785 (O_785,N_4615,N_4839);
nand UO_786 (O_786,N_4735,N_4975);
and UO_787 (O_787,N_4658,N_4634);
nor UO_788 (O_788,N_4706,N_4880);
and UO_789 (O_789,N_4517,N_4656);
xor UO_790 (O_790,N_4821,N_4738);
and UO_791 (O_791,N_4935,N_4918);
xnor UO_792 (O_792,N_4567,N_4538);
and UO_793 (O_793,N_4623,N_4576);
or UO_794 (O_794,N_4935,N_4867);
and UO_795 (O_795,N_4542,N_4593);
and UO_796 (O_796,N_4537,N_4947);
xnor UO_797 (O_797,N_4579,N_4734);
nand UO_798 (O_798,N_4604,N_4591);
nor UO_799 (O_799,N_4546,N_4620);
nand UO_800 (O_800,N_4831,N_4525);
xor UO_801 (O_801,N_4826,N_4851);
nor UO_802 (O_802,N_4688,N_4859);
or UO_803 (O_803,N_4907,N_4836);
nor UO_804 (O_804,N_4723,N_4674);
and UO_805 (O_805,N_4591,N_4995);
nor UO_806 (O_806,N_4561,N_4734);
xor UO_807 (O_807,N_4613,N_4758);
and UO_808 (O_808,N_4736,N_4909);
nand UO_809 (O_809,N_4586,N_4850);
nor UO_810 (O_810,N_4678,N_4971);
or UO_811 (O_811,N_4674,N_4964);
nand UO_812 (O_812,N_4608,N_4939);
xnor UO_813 (O_813,N_4813,N_4845);
and UO_814 (O_814,N_4999,N_4925);
nand UO_815 (O_815,N_4688,N_4862);
xor UO_816 (O_816,N_4734,N_4774);
or UO_817 (O_817,N_4945,N_4728);
xnor UO_818 (O_818,N_4745,N_4667);
and UO_819 (O_819,N_4923,N_4718);
nor UO_820 (O_820,N_4680,N_4771);
and UO_821 (O_821,N_4959,N_4546);
xor UO_822 (O_822,N_4796,N_4541);
and UO_823 (O_823,N_4675,N_4672);
or UO_824 (O_824,N_4980,N_4990);
xor UO_825 (O_825,N_4898,N_4612);
nand UO_826 (O_826,N_4806,N_4734);
and UO_827 (O_827,N_4605,N_4955);
xnor UO_828 (O_828,N_4580,N_4641);
nand UO_829 (O_829,N_4512,N_4825);
or UO_830 (O_830,N_4845,N_4693);
nor UO_831 (O_831,N_4665,N_4957);
nand UO_832 (O_832,N_4775,N_4766);
nor UO_833 (O_833,N_4608,N_4554);
nand UO_834 (O_834,N_4919,N_4970);
and UO_835 (O_835,N_4520,N_4616);
xnor UO_836 (O_836,N_4895,N_4828);
or UO_837 (O_837,N_4538,N_4634);
xnor UO_838 (O_838,N_4963,N_4880);
xnor UO_839 (O_839,N_4950,N_4843);
nand UO_840 (O_840,N_4902,N_4862);
or UO_841 (O_841,N_4621,N_4909);
xor UO_842 (O_842,N_4985,N_4779);
and UO_843 (O_843,N_4593,N_4898);
or UO_844 (O_844,N_4553,N_4652);
and UO_845 (O_845,N_4535,N_4830);
xor UO_846 (O_846,N_4670,N_4917);
or UO_847 (O_847,N_4627,N_4677);
nor UO_848 (O_848,N_4784,N_4503);
nand UO_849 (O_849,N_4739,N_4752);
xor UO_850 (O_850,N_4974,N_4742);
or UO_851 (O_851,N_4921,N_4552);
and UO_852 (O_852,N_4884,N_4724);
and UO_853 (O_853,N_4583,N_4860);
nand UO_854 (O_854,N_4897,N_4841);
and UO_855 (O_855,N_4681,N_4936);
or UO_856 (O_856,N_4823,N_4671);
nand UO_857 (O_857,N_4831,N_4652);
or UO_858 (O_858,N_4751,N_4877);
and UO_859 (O_859,N_4644,N_4797);
and UO_860 (O_860,N_4825,N_4789);
and UO_861 (O_861,N_4744,N_4766);
xor UO_862 (O_862,N_4580,N_4593);
nand UO_863 (O_863,N_4559,N_4617);
nand UO_864 (O_864,N_4989,N_4637);
nor UO_865 (O_865,N_4746,N_4687);
nand UO_866 (O_866,N_4574,N_4891);
or UO_867 (O_867,N_4886,N_4782);
xor UO_868 (O_868,N_4869,N_4678);
xor UO_869 (O_869,N_4754,N_4762);
and UO_870 (O_870,N_4520,N_4810);
nand UO_871 (O_871,N_4944,N_4738);
nor UO_872 (O_872,N_4687,N_4590);
nor UO_873 (O_873,N_4927,N_4510);
nor UO_874 (O_874,N_4679,N_4888);
and UO_875 (O_875,N_4940,N_4634);
and UO_876 (O_876,N_4799,N_4625);
nand UO_877 (O_877,N_4939,N_4607);
xor UO_878 (O_878,N_4880,N_4774);
nand UO_879 (O_879,N_4635,N_4636);
xnor UO_880 (O_880,N_4546,N_4843);
or UO_881 (O_881,N_4526,N_4782);
nor UO_882 (O_882,N_4847,N_4747);
xor UO_883 (O_883,N_4976,N_4693);
and UO_884 (O_884,N_4501,N_4828);
nor UO_885 (O_885,N_4531,N_4952);
nor UO_886 (O_886,N_4611,N_4779);
nand UO_887 (O_887,N_4540,N_4701);
xnor UO_888 (O_888,N_4872,N_4518);
or UO_889 (O_889,N_4896,N_4545);
nand UO_890 (O_890,N_4728,N_4699);
nor UO_891 (O_891,N_4696,N_4758);
xnor UO_892 (O_892,N_4801,N_4613);
nand UO_893 (O_893,N_4890,N_4962);
nor UO_894 (O_894,N_4689,N_4874);
nor UO_895 (O_895,N_4522,N_4945);
nand UO_896 (O_896,N_4642,N_4761);
nor UO_897 (O_897,N_4507,N_4535);
nor UO_898 (O_898,N_4580,N_4968);
nor UO_899 (O_899,N_4949,N_4550);
nor UO_900 (O_900,N_4581,N_4963);
nor UO_901 (O_901,N_4717,N_4843);
and UO_902 (O_902,N_4870,N_4531);
or UO_903 (O_903,N_4989,N_4723);
or UO_904 (O_904,N_4991,N_4619);
nor UO_905 (O_905,N_4904,N_4733);
or UO_906 (O_906,N_4865,N_4501);
xnor UO_907 (O_907,N_4560,N_4813);
and UO_908 (O_908,N_4927,N_4766);
and UO_909 (O_909,N_4951,N_4716);
xnor UO_910 (O_910,N_4716,N_4976);
xnor UO_911 (O_911,N_4595,N_4876);
and UO_912 (O_912,N_4970,N_4651);
nand UO_913 (O_913,N_4727,N_4807);
and UO_914 (O_914,N_4604,N_4790);
and UO_915 (O_915,N_4549,N_4515);
nor UO_916 (O_916,N_4603,N_4591);
and UO_917 (O_917,N_4845,N_4584);
and UO_918 (O_918,N_4770,N_4740);
xnor UO_919 (O_919,N_4501,N_4909);
xnor UO_920 (O_920,N_4884,N_4563);
xnor UO_921 (O_921,N_4529,N_4946);
nand UO_922 (O_922,N_4705,N_4778);
xnor UO_923 (O_923,N_4552,N_4948);
nor UO_924 (O_924,N_4663,N_4922);
nand UO_925 (O_925,N_4588,N_4695);
or UO_926 (O_926,N_4989,N_4521);
or UO_927 (O_927,N_4675,N_4519);
nand UO_928 (O_928,N_4925,N_4604);
xor UO_929 (O_929,N_4967,N_4922);
or UO_930 (O_930,N_4502,N_4801);
nand UO_931 (O_931,N_4671,N_4855);
and UO_932 (O_932,N_4959,N_4744);
xnor UO_933 (O_933,N_4534,N_4805);
or UO_934 (O_934,N_4695,N_4887);
nor UO_935 (O_935,N_4823,N_4840);
nor UO_936 (O_936,N_4819,N_4823);
xor UO_937 (O_937,N_4807,N_4625);
or UO_938 (O_938,N_4714,N_4618);
nand UO_939 (O_939,N_4621,N_4519);
and UO_940 (O_940,N_4756,N_4504);
or UO_941 (O_941,N_4904,N_4754);
xor UO_942 (O_942,N_4807,N_4578);
nor UO_943 (O_943,N_4678,N_4768);
or UO_944 (O_944,N_4752,N_4648);
nand UO_945 (O_945,N_4730,N_4699);
xor UO_946 (O_946,N_4773,N_4884);
or UO_947 (O_947,N_4943,N_4591);
nand UO_948 (O_948,N_4900,N_4715);
nand UO_949 (O_949,N_4618,N_4530);
nor UO_950 (O_950,N_4945,N_4674);
and UO_951 (O_951,N_4746,N_4841);
or UO_952 (O_952,N_4630,N_4985);
xnor UO_953 (O_953,N_4511,N_4885);
or UO_954 (O_954,N_4558,N_4599);
nand UO_955 (O_955,N_4713,N_4535);
and UO_956 (O_956,N_4608,N_4515);
xor UO_957 (O_957,N_4708,N_4785);
xor UO_958 (O_958,N_4570,N_4780);
and UO_959 (O_959,N_4603,N_4864);
xnor UO_960 (O_960,N_4958,N_4683);
or UO_961 (O_961,N_4697,N_4506);
or UO_962 (O_962,N_4820,N_4831);
nand UO_963 (O_963,N_4985,N_4512);
xnor UO_964 (O_964,N_4692,N_4611);
and UO_965 (O_965,N_4839,N_4954);
nor UO_966 (O_966,N_4563,N_4670);
nor UO_967 (O_967,N_4900,N_4612);
and UO_968 (O_968,N_4849,N_4697);
and UO_969 (O_969,N_4735,N_4920);
nor UO_970 (O_970,N_4799,N_4862);
xnor UO_971 (O_971,N_4631,N_4907);
or UO_972 (O_972,N_4857,N_4525);
xor UO_973 (O_973,N_4833,N_4995);
or UO_974 (O_974,N_4722,N_4848);
nor UO_975 (O_975,N_4634,N_4514);
or UO_976 (O_976,N_4833,N_4904);
nor UO_977 (O_977,N_4568,N_4938);
xor UO_978 (O_978,N_4670,N_4577);
nor UO_979 (O_979,N_4709,N_4518);
nand UO_980 (O_980,N_4708,N_4678);
xnor UO_981 (O_981,N_4948,N_4915);
nand UO_982 (O_982,N_4953,N_4725);
nand UO_983 (O_983,N_4500,N_4889);
nor UO_984 (O_984,N_4642,N_4817);
or UO_985 (O_985,N_4876,N_4501);
and UO_986 (O_986,N_4705,N_4942);
nor UO_987 (O_987,N_4850,N_4555);
nor UO_988 (O_988,N_4523,N_4728);
xnor UO_989 (O_989,N_4613,N_4626);
xor UO_990 (O_990,N_4998,N_4899);
or UO_991 (O_991,N_4915,N_4809);
nand UO_992 (O_992,N_4995,N_4523);
and UO_993 (O_993,N_4716,N_4802);
xnor UO_994 (O_994,N_4794,N_4724);
nand UO_995 (O_995,N_4985,N_4578);
or UO_996 (O_996,N_4942,N_4598);
nand UO_997 (O_997,N_4852,N_4944);
nor UO_998 (O_998,N_4823,N_4965);
nor UO_999 (O_999,N_4526,N_4864);
endmodule