module basic_2000_20000_2500_40_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_1029,In_1190);
nand U1 (N_1,In_858,In_24);
and U2 (N_2,In_1183,In_1570);
and U3 (N_3,In_1701,In_767);
xnor U4 (N_4,In_998,In_351);
or U5 (N_5,In_1810,In_1678);
nor U6 (N_6,In_1192,In_985);
and U7 (N_7,In_1344,In_1267);
nor U8 (N_8,In_301,In_1543);
nor U9 (N_9,In_1459,In_1776);
nor U10 (N_10,In_1057,In_457);
or U11 (N_11,In_745,In_996);
and U12 (N_12,In_1974,In_1979);
xnor U13 (N_13,In_342,In_678);
xnor U14 (N_14,In_1823,In_1608);
nor U15 (N_15,In_336,In_674);
or U16 (N_16,In_1067,In_1493);
or U17 (N_17,In_1902,In_448);
nor U18 (N_18,In_785,In_790);
or U19 (N_19,In_406,In_1405);
or U20 (N_20,In_1603,In_1573);
nand U21 (N_21,In_832,In_1085);
nor U22 (N_22,In_1504,In_1754);
and U23 (N_23,In_496,In_868);
or U24 (N_24,In_1772,In_1592);
and U25 (N_25,In_140,In_234);
xnor U26 (N_26,In_999,In_219);
nand U27 (N_27,In_601,In_1092);
and U28 (N_28,In_1956,In_704);
xor U29 (N_29,In_1855,In_1071);
or U30 (N_30,In_1125,In_1893);
or U31 (N_31,In_501,In_10);
or U32 (N_32,In_886,In_1926);
and U33 (N_33,In_165,In_565);
xnor U34 (N_34,In_300,In_1294);
nor U35 (N_35,In_1006,In_1891);
xor U36 (N_36,In_407,In_1640);
nor U37 (N_37,In_839,In_1312);
nor U38 (N_38,In_420,In_1295);
and U39 (N_39,In_1909,In_1148);
and U40 (N_40,In_1717,In_1545);
and U41 (N_41,In_310,In_396);
xor U42 (N_42,In_1491,In_1691);
nand U43 (N_43,In_375,In_1673);
nand U44 (N_44,In_600,In_1601);
and U45 (N_45,In_294,In_1900);
nor U46 (N_46,In_632,In_841);
xnor U47 (N_47,In_8,In_1554);
nand U48 (N_48,In_722,In_1813);
and U49 (N_49,In_676,In_166);
and U50 (N_50,In_810,In_987);
and U51 (N_51,In_1099,In_932);
nand U52 (N_52,In_459,In_1866);
or U53 (N_53,In_1858,In_1273);
nand U54 (N_54,In_1164,In_520);
nand U55 (N_55,In_1381,In_504);
and U56 (N_56,In_1895,In_603);
xnor U57 (N_57,In_700,In_312);
nor U58 (N_58,In_107,In_837);
and U59 (N_59,In_1515,In_1809);
nand U60 (N_60,In_1285,In_126);
xor U61 (N_61,In_1774,In_432);
or U62 (N_62,In_919,In_874);
nand U63 (N_63,In_626,In_355);
and U64 (N_64,In_694,In_1685);
or U65 (N_65,In_951,In_1014);
nor U66 (N_66,In_1366,In_307);
xor U67 (N_67,In_1734,In_1654);
or U68 (N_68,In_763,In_833);
nor U69 (N_69,In_1886,In_945);
or U70 (N_70,In_713,In_1216);
and U71 (N_71,In_428,In_1093);
nor U72 (N_72,In_1751,In_1514);
and U73 (N_73,In_1311,In_575);
nor U74 (N_74,In_1676,In_1781);
and U75 (N_75,In_1972,In_792);
nand U76 (N_76,In_612,In_887);
xnor U77 (N_77,In_404,In_1477);
nor U78 (N_78,In_1013,In_321);
and U79 (N_79,In_71,In_619);
and U80 (N_80,In_1547,In_31);
nor U81 (N_81,In_1506,In_395);
nor U82 (N_82,In_750,In_820);
nor U83 (N_83,In_954,In_1338);
or U84 (N_84,In_818,In_1779);
and U85 (N_85,In_559,In_156);
xnor U86 (N_86,In_655,In_1869);
or U87 (N_87,In_1200,In_22);
nand U88 (N_88,In_1523,In_550);
xor U89 (N_89,In_167,In_807);
and U90 (N_90,In_1474,In_1602);
nor U91 (N_91,In_1137,In_563);
and U92 (N_92,In_374,In_37);
nor U93 (N_93,In_1769,In_1121);
or U94 (N_94,In_215,In_1532);
and U95 (N_95,In_123,In_667);
nor U96 (N_96,In_445,In_1144);
and U97 (N_97,In_353,In_150);
nor U98 (N_98,In_341,In_1320);
nor U99 (N_99,In_693,In_1931);
or U100 (N_100,In_794,In_109);
and U101 (N_101,In_1213,In_1198);
xnor U102 (N_102,In_1430,In_1173);
xor U103 (N_103,In_1923,In_1243);
nand U104 (N_104,In_884,In_689);
nor U105 (N_105,In_1229,In_196);
xor U106 (N_106,In_203,In_613);
nor U107 (N_107,In_1332,In_392);
xnor U108 (N_108,In_1594,In_831);
xnor U109 (N_109,In_471,In_617);
nor U110 (N_110,In_828,In_1143);
nor U111 (N_111,In_178,In_553);
nor U112 (N_112,In_524,In_1871);
nand U113 (N_113,In_1537,In_939);
nor U114 (N_114,In_1916,In_387);
xor U115 (N_115,In_1657,In_528);
or U116 (N_116,In_182,In_222);
nand U117 (N_117,In_1560,In_174);
nor U118 (N_118,In_510,In_1083);
and U119 (N_119,In_1921,In_105);
xnor U120 (N_120,In_1520,In_724);
nor U121 (N_121,In_606,In_946);
xor U122 (N_122,In_1385,In_1262);
or U123 (N_123,In_51,In_1157);
and U124 (N_124,In_1833,In_1806);
nor U125 (N_125,In_1363,In_1845);
nand U126 (N_126,In_598,In_350);
or U127 (N_127,In_1933,In_1219);
xnor U128 (N_128,In_229,In_1282);
and U129 (N_129,In_475,In_296);
xnor U130 (N_130,In_1720,In_1829);
xor U131 (N_131,In_1114,In_1432);
xnor U132 (N_132,In_369,In_1470);
and U133 (N_133,In_86,In_656);
nor U134 (N_134,In_1724,In_1945);
or U135 (N_135,In_1204,In_611);
nand U136 (N_136,In_1247,In_1087);
or U137 (N_137,In_1647,In_1703);
xor U138 (N_138,In_1302,In_904);
or U139 (N_139,In_335,In_200);
nand U140 (N_140,In_882,In_231);
nor U141 (N_141,In_79,In_492);
and U142 (N_142,In_1863,In_1374);
nand U143 (N_143,In_1175,In_1544);
and U144 (N_144,In_1924,In_444);
nand U145 (N_145,In_1737,In_1787);
and U146 (N_146,In_899,In_652);
or U147 (N_147,In_1696,In_771);
nor U148 (N_148,In_1670,In_1815);
and U149 (N_149,In_1788,In_394);
xor U150 (N_150,In_777,In_188);
nand U151 (N_151,In_212,In_1770);
xor U152 (N_152,In_153,In_703);
nor U153 (N_153,In_1558,In_1429);
nor U154 (N_154,In_639,In_835);
nand U155 (N_155,In_1347,In_218);
or U156 (N_156,In_1874,In_1202);
nor U157 (N_157,In_786,In_1596);
and U158 (N_158,In_1934,In_25);
nor U159 (N_159,In_1847,In_1453);
and U160 (N_160,In_737,In_1726);
and U161 (N_161,In_881,In_190);
and U162 (N_162,In_1290,In_357);
nand U163 (N_163,In_930,In_823);
and U164 (N_164,In_1919,In_1220);
and U165 (N_165,In_1153,In_1605);
xor U166 (N_166,In_1010,In_356);
nor U167 (N_167,In_1998,In_303);
or U168 (N_168,In_93,In_329);
nor U169 (N_169,In_263,In_938);
xnor U170 (N_170,In_1653,In_1988);
and U171 (N_171,In_850,In_1380);
and U172 (N_172,In_1476,In_1797);
xnor U173 (N_173,In_813,In_1613);
nor U174 (N_174,In_430,In_244);
and U175 (N_175,In_684,In_615);
xnor U176 (N_176,In_217,In_1040);
nand U177 (N_177,In_1597,In_633);
or U178 (N_178,In_423,In_1086);
nor U179 (N_179,In_408,In_585);
nor U180 (N_180,In_112,In_1034);
nand U181 (N_181,In_458,In_1619);
nor U182 (N_182,In_1709,In_122);
or U183 (N_183,In_378,In_1637);
xnor U184 (N_184,In_1076,In_900);
or U185 (N_185,In_1616,In_1671);
or U186 (N_186,In_427,In_685);
xor U187 (N_187,In_1897,In_266);
or U188 (N_188,In_172,In_1394);
or U189 (N_189,In_1827,In_108);
xnor U190 (N_190,In_1343,In_1281);
and U191 (N_191,In_1349,In_1237);
and U192 (N_192,In_1700,In_1912);
xnor U193 (N_193,In_1584,In_509);
or U194 (N_194,In_1880,In_1463);
nand U195 (N_195,In_1288,In_869);
xnor U196 (N_196,In_1860,In_663);
xor U197 (N_197,In_1599,In_1208);
and U198 (N_198,In_368,In_1796);
or U199 (N_199,In_711,In_1830);
or U200 (N_200,In_1231,In_1283);
and U201 (N_201,In_867,In_1120);
and U202 (N_202,In_1705,In_1245);
or U203 (N_203,In_959,In_1254);
xnor U204 (N_204,In_758,In_1929);
and U205 (N_205,In_1064,In_242);
xor U206 (N_206,In_669,In_1728);
xor U207 (N_207,In_670,In_592);
and U208 (N_208,In_1206,In_1449);
nor U209 (N_209,In_1882,In_449);
xor U210 (N_210,In_1509,In_1910);
nor U211 (N_211,In_579,In_1334);
nand U212 (N_212,In_1081,In_915);
or U213 (N_213,In_1595,In_1066);
xnor U214 (N_214,In_1309,In_16);
or U215 (N_215,In_1350,In_717);
and U216 (N_216,In_1741,In_805);
and U217 (N_217,In_686,In_1170);
xor U218 (N_218,In_1364,In_1588);
nor U219 (N_219,In_1759,In_534);
or U220 (N_220,In_829,In_1488);
or U221 (N_221,In_173,In_610);
nor U222 (N_222,In_1318,In_1140);
nand U223 (N_223,In_339,In_735);
or U224 (N_224,In_1090,In_776);
xnor U225 (N_225,In_1244,In_246);
nand U226 (N_226,In_232,In_587);
nor U227 (N_227,In_290,In_1328);
nor U228 (N_228,In_326,In_485);
nor U229 (N_229,In_84,In_1358);
or U230 (N_230,In_1511,In_1854);
and U231 (N_231,In_488,In_812);
xor U232 (N_232,In_808,In_1186);
nor U233 (N_233,In_224,In_936);
nor U234 (N_234,In_1296,In_46);
and U235 (N_235,In_1324,In_861);
xnor U236 (N_236,In_718,In_625);
or U237 (N_237,In_1339,In_1398);
xor U238 (N_238,In_1005,In_1433);
nor U239 (N_239,In_1417,In_1443);
or U240 (N_240,In_903,In_556);
or U241 (N_241,In_1379,In_1128);
or U242 (N_242,In_913,In_1714);
nor U243 (N_243,In_283,In_741);
nor U244 (N_244,In_822,In_1913);
and U245 (N_245,In_1444,In_1939);
and U246 (N_246,In_104,In_1775);
and U247 (N_247,In_584,In_997);
and U248 (N_248,In_943,In_1961);
and U249 (N_249,In_431,In_1825);
nand U250 (N_250,In_1335,In_209);
nand U251 (N_251,In_1628,In_14);
and U252 (N_252,In_309,In_0);
or U253 (N_253,In_1305,In_1533);
xor U254 (N_254,In_132,In_1549);
and U255 (N_255,In_605,In_1473);
nor U256 (N_256,In_546,In_415);
or U257 (N_257,In_1329,In_1760);
and U258 (N_258,In_791,In_262);
xor U259 (N_259,In_1160,In_1408);
nand U260 (N_260,In_1008,In_1950);
or U261 (N_261,In_1261,In_1053);
and U262 (N_262,In_1614,In_1710);
nor U263 (N_263,In_1315,In_1373);
xor U264 (N_264,In_762,In_705);
and U265 (N_265,In_1074,In_1842);
nor U266 (N_266,In_1421,In_1069);
nand U267 (N_267,In_865,In_549);
nor U268 (N_268,In_1356,In_1036);
and U269 (N_269,In_41,In_1957);
and U270 (N_270,In_422,In_1032);
nor U271 (N_271,In_966,In_564);
nor U272 (N_272,In_1994,In_917);
nor U273 (N_273,In_1227,In_1745);
or U274 (N_274,In_964,In_637);
nor U275 (N_275,In_732,In_49);
nor U276 (N_276,In_80,In_484);
nand U277 (N_277,In_57,In_1181);
and U278 (N_278,In_1807,In_382);
nor U279 (N_279,In_1765,In_1098);
or U280 (N_280,In_1841,In_235);
or U281 (N_281,In_749,In_384);
xnor U282 (N_282,In_541,In_738);
nor U283 (N_283,In_346,In_184);
xor U284 (N_284,In_1031,In_1660);
xor U285 (N_285,In_163,In_463);
nand U286 (N_286,In_586,In_747);
and U287 (N_287,In_281,In_538);
nor U288 (N_288,In_1451,In_1415);
nor U289 (N_289,In_1481,In_1423);
nand U290 (N_290,In_1413,In_1650);
and U291 (N_291,In_1968,In_1611);
nor U292 (N_292,In_1983,In_1702);
and U293 (N_293,In_1757,In_844);
nor U294 (N_294,In_1753,In_77);
nor U295 (N_295,In_434,In_1027);
and U296 (N_296,In_1041,In_1351);
and U297 (N_297,In_802,In_784);
nand U298 (N_298,In_358,In_1412);
nor U299 (N_299,In_1655,In_277);
or U300 (N_300,In_1591,In_1659);
and U301 (N_301,In_755,In_1145);
nand U302 (N_302,In_1191,In_620);
or U303 (N_303,In_1308,In_171);
nand U304 (N_304,In_1297,In_500);
and U305 (N_305,In_1359,In_1428);
nand U306 (N_306,In_1284,In_1836);
nand U307 (N_307,In_662,In_852);
nor U308 (N_308,In_1538,In_54);
nand U309 (N_309,In_1264,In_1452);
nand U310 (N_310,In_1630,In_1130);
and U311 (N_311,In_855,In_214);
nor U312 (N_312,In_521,In_142);
nor U313 (N_313,In_1049,In_1127);
nor U314 (N_314,In_474,In_1168);
xor U315 (N_315,In_349,In_29);
and U316 (N_316,In_816,In_780);
or U317 (N_317,In_795,In_533);
or U318 (N_318,In_118,In_1859);
xnor U319 (N_319,In_161,In_1684);
nand U320 (N_320,In_1265,In_890);
or U321 (N_321,In_1068,In_443);
nand U322 (N_322,In_1814,In_1579);
and U323 (N_323,In_896,In_1583);
xor U324 (N_324,In_1156,In_421);
and U325 (N_325,In_590,In_1821);
and U326 (N_326,In_1489,In_716);
or U327 (N_327,In_1188,In_419);
or U328 (N_328,In_1773,In_1028);
xnor U329 (N_329,In_977,In_177);
nand U330 (N_330,In_806,In_895);
xnor U331 (N_331,In_1299,In_1868);
nand U332 (N_332,In_1211,In_1341);
and U333 (N_333,In_687,In_748);
and U334 (N_334,In_59,In_920);
and U335 (N_335,In_1623,In_284);
and U336 (N_336,In_1197,In_410);
and U337 (N_337,In_1632,In_1426);
or U338 (N_338,In_1557,In_1508);
or U339 (N_339,In_75,In_1954);
xnor U340 (N_340,In_1325,In_250);
or U341 (N_341,In_1536,In_1436);
or U342 (N_342,In_906,In_1958);
xor U343 (N_343,In_1326,In_1292);
nor U344 (N_344,In_1711,In_390);
xor U345 (N_345,In_1952,In_1870);
and U346 (N_346,In_712,In_877);
nor U347 (N_347,In_1060,In_1203);
and U348 (N_348,In_388,In_983);
and U349 (N_349,In_1030,In_562);
or U350 (N_350,In_1486,In_1944);
xnor U351 (N_351,In_253,In_1688);
nor U352 (N_352,In_468,In_532);
or U353 (N_353,In_48,In_441);
nand U354 (N_354,In_1903,In_1963);
or U355 (N_355,In_146,In_20);
or U356 (N_356,In_513,In_682);
and U357 (N_357,In_1925,In_27);
nand U358 (N_358,In_101,In_769);
and U359 (N_359,In_1510,In_931);
xnor U360 (N_360,In_1990,In_1758);
nor U361 (N_361,In_1025,In_1499);
or U362 (N_362,In_1503,In_1966);
or U363 (N_363,In_846,In_45);
and U364 (N_364,In_1877,In_824);
and U365 (N_365,In_811,In_537);
or U366 (N_366,In_379,In_1377);
nor U367 (N_367,In_69,In_1755);
or U368 (N_368,In_657,In_1675);
nor U369 (N_369,In_186,In_1620);
nor U370 (N_370,In_1340,In_258);
nand U371 (N_371,In_1468,In_642);
or U372 (N_372,In_187,In_1906);
and U373 (N_373,In_757,In_481);
xnor U374 (N_374,In_1686,In_1166);
nand U375 (N_375,In_1484,In_653);
xor U376 (N_376,In_1995,In_120);
xnor U377 (N_377,In_1763,In_143);
nand U378 (N_378,In_1849,In_1624);
nor U379 (N_379,In_58,In_486);
nor U380 (N_380,In_1795,In_154);
and U381 (N_381,In_1445,In_23);
or U382 (N_382,In_1985,In_331);
xor U383 (N_383,In_95,In_1141);
and U384 (N_384,In_1269,In_1310);
or U385 (N_385,In_1004,In_1690);
or U386 (N_386,In_1593,In_1246);
nand U387 (N_387,In_1680,In_1942);
nor U388 (N_388,In_561,In_1865);
or U389 (N_389,In_1885,In_498);
and U390 (N_390,In_1565,In_1852);
and U391 (N_391,In_539,In_1330);
xnor U392 (N_392,In_1798,In_1129);
nor U393 (N_393,In_627,In_1276);
or U394 (N_394,In_380,In_117);
or U395 (N_395,In_1996,In_413);
nor U396 (N_396,In_1274,In_1023);
nand U397 (N_397,In_1879,In_1035);
or U398 (N_398,In_1839,In_55);
nand U399 (N_399,In_1406,In_1563);
or U400 (N_400,In_1255,In_479);
xor U401 (N_401,In_87,In_551);
nor U402 (N_402,In_1179,In_1643);
or U403 (N_403,In_1577,In_761);
nand U404 (N_404,In_1662,In_742);
nor U405 (N_405,In_1975,In_894);
nor U406 (N_406,In_1138,In_6);
xnor U407 (N_407,In_238,In_345);
xor U408 (N_408,In_1492,In_1762);
nor U409 (N_409,In_1250,In_1997);
nand U410 (N_410,In_401,In_292);
and U411 (N_411,In_1124,In_455);
nand U412 (N_412,In_1768,In_1258);
nand U413 (N_413,In_452,In_450);
and U414 (N_414,In_53,In_1420);
xor U415 (N_415,In_333,In_683);
or U416 (N_416,In_1749,In_111);
or U417 (N_417,In_106,In_950);
and U418 (N_418,In_892,In_1861);
nand U419 (N_419,In_1930,In_1884);
nor U420 (N_420,In_1892,In_1189);
nor U421 (N_421,In_466,In_1740);
nand U422 (N_422,In_1331,In_1824);
nor U423 (N_423,In_1947,In_860);
and U424 (N_424,In_1345,In_1552);
nand U425 (N_425,In_323,In_298);
nand U426 (N_426,In_287,In_759);
nand U427 (N_427,In_1722,In_52);
xnor U428 (N_428,In_988,In_1050);
xnor U429 (N_429,In_594,In_1981);
nand U430 (N_430,In_522,In_297);
or U431 (N_431,In_1362,In_1001);
or U432 (N_432,In_1915,In_982);
nand U433 (N_433,In_26,In_672);
or U434 (N_434,In_1615,In_337);
nand U435 (N_435,In_990,In_183);
xor U436 (N_436,In_385,In_168);
or U437 (N_437,In_1840,In_1002);
nand U438 (N_438,In_1372,In_1626);
or U439 (N_439,In_609,In_871);
and U440 (N_440,In_644,In_1392);
nor U441 (N_441,In_1382,In_347);
and U442 (N_442,In_905,In_596);
xnor U443 (N_443,In_873,In_1908);
nand U444 (N_444,In_815,In_961);
nor U445 (N_445,In_1395,In_181);
nor U446 (N_446,In_1802,In_1646);
nand U447 (N_447,In_1907,In_1631);
or U448 (N_448,In_70,In_328);
xor U449 (N_449,In_502,In_1525);
nor U450 (N_450,In_544,In_1209);
nand U451 (N_451,In_195,In_1464);
nor U452 (N_452,In_416,In_487);
nor U453 (N_453,In_447,In_372);
and U454 (N_454,In_1419,In_1386);
and U455 (N_455,In_1977,In_876);
and U456 (N_456,In_1529,In_872);
and U457 (N_457,In_1117,In_1941);
xor U458 (N_458,In_426,In_1289);
and U459 (N_459,In_680,In_113);
xor U460 (N_460,In_194,In_373);
and U461 (N_461,In_1521,In_1911);
xor U462 (N_462,In_293,In_654);
xor U463 (N_463,In_754,In_1546);
xnor U464 (N_464,In_313,In_1007);
and U465 (N_465,In_1946,In_1832);
or U466 (N_466,In_456,In_343);
or U467 (N_467,In_1404,In_1948);
nand U468 (N_468,In_885,In_1959);
and U469 (N_469,In_1550,In_1820);
xnor U470 (N_470,In_993,In_1649);
and U471 (N_471,In_972,In_189);
nand U472 (N_472,In_1073,In_1712);
or U473 (N_473,In_1495,In_640);
nand U474 (N_474,In_1039,In_1991);
and U475 (N_475,In_169,In_1771);
nand U476 (N_476,In_723,In_523);
and U477 (N_477,In_207,In_542);
or U478 (N_478,In_679,In_949);
or U479 (N_479,In_237,In_578);
or U480 (N_480,In_1767,In_360);
nand U481 (N_481,In_702,In_147);
and U482 (N_482,In_125,In_1618);
nand U483 (N_483,In_840,In_1864);
xor U484 (N_484,In_1287,In_1883);
and U485 (N_485,In_1812,In_446);
and U486 (N_486,In_412,In_304);
nor U487 (N_487,In_1816,In_1058);
nor U488 (N_488,In_1078,In_650);
or U489 (N_489,In_740,In_100);
nand U490 (N_490,In_89,In_478);
xor U491 (N_491,In_692,In_267);
and U492 (N_492,In_260,In_1964);
or U493 (N_493,In_288,In_1727);
nor U494 (N_494,In_1427,In_1410);
nor U495 (N_495,In_1185,In_1169);
nand U496 (N_496,In_916,In_854);
xor U497 (N_497,In_1642,In_1526);
and U498 (N_498,In_1844,In_221);
xnor U499 (N_499,In_7,In_1600);
and U500 (N_500,In_1391,In_1713);
xnor U501 (N_501,N_48,In_213);
xnor U502 (N_502,In_773,N_343);
xnor U503 (N_503,In_1890,N_11);
nand U504 (N_504,In_1411,In_1578);
and U505 (N_505,N_465,N_82);
nand U506 (N_506,In_941,N_391);
nor U507 (N_507,N_14,In_760);
nand U508 (N_508,N_194,N_90);
or U509 (N_509,In_1682,In_256);
nor U510 (N_510,N_395,In_614);
nor U511 (N_511,In_1454,In_1277);
nor U512 (N_512,In_1656,N_65);
nand U513 (N_513,N_172,N_466);
nand U514 (N_514,In_1176,N_443);
and U515 (N_515,N_58,In_540);
nand U516 (N_516,N_220,N_486);
nor U517 (N_517,In_1791,In_1633);
and U518 (N_518,In_103,In_536);
and U519 (N_519,In_464,In_13);
and U520 (N_520,In_1735,N_269);
nor U521 (N_521,In_783,In_73);
and U522 (N_522,N_420,N_254);
or U523 (N_523,In_923,In_1752);
or U524 (N_524,In_1725,In_12);
and U525 (N_525,N_95,In_1011);
or U526 (N_526,In_1252,In_1218);
nand U527 (N_527,In_362,In_204);
nor U528 (N_528,In_505,N_185);
xnor U529 (N_529,In_1803,N_318);
nor U530 (N_530,N_436,N_334);
or U531 (N_531,In_1161,In_102);
xor U532 (N_532,In_47,In_1665);
nor U533 (N_533,N_402,In_1012);
and U534 (N_534,In_766,In_361);
nand U535 (N_535,N_227,N_474);
xor U536 (N_536,In_1784,N_68);
xor U537 (N_537,In_1111,In_82);
xor U538 (N_538,In_175,In_1167);
xnor U539 (N_539,In_1571,N_175);
or U540 (N_540,N_215,In_1441);
or U541 (N_541,N_419,In_889);
or U542 (N_542,In_247,In_418);
xnor U543 (N_543,N_31,In_99);
nand U544 (N_544,In_1920,In_1249);
and U545 (N_545,In_708,In_74);
nor U546 (N_546,In_241,In_1052);
and U547 (N_547,In_1112,In_220);
nand U548 (N_548,In_719,In_170);
nor U549 (N_549,In_17,N_271);
and U550 (N_550,N_96,In_734);
xnor U551 (N_551,In_1314,In_1695);
nand U552 (N_552,N_446,In_136);
nand U553 (N_553,N_8,In_696);
or U554 (N_554,In_548,N_26);
and U555 (N_555,N_481,In_582);
nor U556 (N_556,In_746,N_358);
xor U557 (N_557,N_107,N_5);
nor U558 (N_558,N_331,In_1524);
or U559 (N_559,In_1540,In_1790);
and U560 (N_560,In_825,In_273);
nand U561 (N_561,N_206,In_302);
nor U562 (N_562,In_128,N_428);
or U563 (N_563,N_405,In_1178);
xor U564 (N_564,In_133,In_583);
nand U565 (N_565,In_843,N_74);
nor U566 (N_566,N_484,In_963);
nand U567 (N_567,In_1739,In_1253);
and U568 (N_568,In_1743,N_429);
or U569 (N_569,In_589,In_1106);
nand U570 (N_570,In_727,N_21);
xor U571 (N_571,In_397,In_442);
xnor U572 (N_572,In_701,In_1786);
nand U573 (N_573,N_339,In_233);
nor U574 (N_574,In_1542,In_1539);
or U575 (N_575,In_1103,N_388);
and U576 (N_576,N_151,N_114);
nor U577 (N_577,N_246,In_1699);
and U578 (N_578,N_119,In_334);
xor U579 (N_579,N_273,In_1898);
xor U580 (N_580,N_417,In_1465);
xor U581 (N_581,In_1021,In_781);
xor U582 (N_582,In_127,In_516);
and U583 (N_583,In_1355,N_201);
and U584 (N_584,N_311,N_150);
and U585 (N_585,N_132,N_4);
and U586 (N_586,In_470,In_1187);
nand U587 (N_587,N_463,In_1361);
and U588 (N_588,In_1555,N_208);
nor U589 (N_589,In_1609,In_1482);
or U590 (N_590,In_607,In_1396);
nor U591 (N_591,In_85,In_42);
nor U592 (N_592,In_1694,In_285);
nand U593 (N_593,In_1096,In_252);
or U594 (N_594,In_666,N_156);
nand U595 (N_595,In_311,In_436);
nor U596 (N_596,In_1848,N_492);
nor U597 (N_597,N_469,N_319);
nor U598 (N_598,In_1580,In_50);
nor U599 (N_599,In_1306,In_148);
nand U600 (N_600,N_401,In_36);
xor U601 (N_601,N_448,N_332);
or U602 (N_602,N_360,N_221);
nor U603 (N_603,In_1872,N_476);
nand U604 (N_604,N_346,In_192);
nor U605 (N_605,N_37,In_1462);
xor U606 (N_606,In_1561,N_413);
nand U607 (N_607,N_441,In_879);
nor U608 (N_608,In_199,N_71);
nor U609 (N_609,N_310,N_345);
or U610 (N_610,In_270,In_489);
nand U611 (N_611,In_695,In_1467);
and U612 (N_612,In_744,In_665);
and U613 (N_613,In_710,N_421);
nand U614 (N_614,In_1376,In_324);
or U615 (N_615,In_503,In_411);
nor U616 (N_616,In_1777,In_78);
nor U617 (N_617,N_171,In_1617);
and U618 (N_618,N_27,N_479);
or U619 (N_619,In_554,In_671);
or U620 (N_620,N_181,In_1046);
and U621 (N_621,N_35,In_1371);
or U622 (N_622,In_1123,N_385);
xnor U623 (N_623,In_1697,In_1055);
xor U624 (N_624,In_743,In_878);
nand U625 (N_625,N_293,In_1024);
or U626 (N_626,In_417,In_1980);
nand U627 (N_627,In_1418,In_1606);
nand U628 (N_628,In_1992,N_88);
xnor U629 (N_629,In_67,N_426);
and U630 (N_630,In_135,N_362);
or U631 (N_631,In_1478,In_1512);
nand U632 (N_632,In_1077,In_739);
nand U633 (N_633,In_1748,In_90);
nor U634 (N_634,In_1687,N_392);
and U635 (N_635,In_1519,In_1182);
xor U636 (N_636,In_364,In_1360);
nor U637 (N_637,In_1955,In_391);
and U638 (N_638,In_155,In_254);
xnor U639 (N_639,In_1088,In_145);
nor U640 (N_640,In_1692,In_1065);
xnor U641 (N_641,N_316,In_636);
nand U642 (N_642,In_306,N_209);
and U643 (N_643,N_3,In_688);
xnor U644 (N_644,In_1736,N_79);
nor U645 (N_645,N_471,N_279);
nor U646 (N_646,In_979,In_56);
and U647 (N_647,In_1894,In_965);
xnor U648 (N_648,In_409,In_97);
and U649 (N_649,In_1707,N_349);
and U650 (N_650,N_296,N_39);
xor U651 (N_651,In_1575,In_1517);
or U652 (N_652,N_255,In_1610);
nor U653 (N_653,In_299,In_1147);
or U654 (N_654,N_178,N_376);
xnor U655 (N_655,In_1063,In_1733);
nand U656 (N_656,In_1993,In_1108);
or U657 (N_657,In_555,In_1199);
or U658 (N_658,N_307,In_1982);
nand U659 (N_659,In_291,In_1193);
and U660 (N_660,N_280,N_399);
nor U661 (N_661,In_1152,N_406);
and U662 (N_662,N_60,In_1469);
xor U663 (N_663,N_439,In_1223);
xnor U664 (N_664,In_1846,N_485);
or U665 (N_665,In_864,In_1317);
or U666 (N_666,In_847,In_201);
xnor U667 (N_667,In_1976,In_641);
nor U668 (N_668,In_1447,In_1446);
nor U669 (N_669,N_118,In_782);
nor U670 (N_670,N_112,In_1230);
and U671 (N_671,In_910,In_921);
or U672 (N_672,In_315,N_472);
or U673 (N_673,N_93,In_134);
nor U674 (N_674,N_387,In_1887);
nor U675 (N_675,In_658,In_517);
nor U676 (N_676,In_1159,N_184);
nand U677 (N_677,In_918,N_289);
xnor U678 (N_678,In_1574,In_1016);
xor U679 (N_679,In_901,N_435);
or U680 (N_680,In_1801,In_386);
xor U681 (N_681,N_249,In_1072);
nor U682 (N_682,In_1256,N_383);
and U683 (N_683,In_518,In_530);
nand U684 (N_684,In_573,N_84);
nor U685 (N_685,N_449,N_287);
or U686 (N_686,In_897,In_1501);
or U687 (N_687,In_1319,In_9);
nand U688 (N_688,In_1037,In_506);
and U689 (N_689,In_1800,In_756);
or U690 (N_690,In_1416,N_497);
or U691 (N_691,N_62,N_368);
nand U692 (N_692,In_571,In_72);
nor U693 (N_693,In_491,N_453);
nand U694 (N_694,N_251,N_142);
nor U695 (N_695,N_214,In_371);
or U696 (N_696,In_709,In_621);
nor U697 (N_697,In_924,In_19);
or U698 (N_698,In_1215,N_72);
or U699 (N_699,In_995,In_305);
xor U700 (N_700,N_414,In_1940);
or U701 (N_701,In_992,N_258);
and U702 (N_702,In_1978,N_63);
nand U703 (N_703,N_372,In_1100);
nor U704 (N_704,In_129,N_92);
or U705 (N_705,In_937,In_570);
or U706 (N_706,In_994,In_1224);
xnor U707 (N_707,N_105,In_1407);
xnor U708 (N_708,In_857,N_285);
and U709 (N_709,In_893,N_136);
or U710 (N_710,In_476,In_2);
nor U711 (N_711,N_330,In_922);
or U712 (N_712,In_497,In_124);
and U713 (N_713,In_1422,In_591);
nor U714 (N_714,In_1251,N_243);
xnor U715 (N_715,In_1587,In_856);
or U716 (N_716,In_1598,In_1280);
nand U717 (N_717,N_19,In_631);
nand U718 (N_718,In_1518,In_927);
nor U719 (N_719,N_245,In_902);
nand U720 (N_720,In_96,N_212);
nor U721 (N_721,N_315,N_430);
xor U722 (N_722,In_1582,N_393);
or U723 (N_723,N_217,In_1142);
xnor U724 (N_724,In_249,In_1764);
xnor U725 (N_725,In_942,In_593);
xnor U726 (N_726,In_275,In_64);
nor U727 (N_727,In_1180,In_1047);
or U728 (N_728,N_238,In_366);
or U729 (N_729,In_1922,In_567);
xor U730 (N_730,N_149,N_305);
nand U731 (N_731,In_208,In_1918);
or U732 (N_732,In_527,In_308);
or U733 (N_733,In_1516,In_1971);
xnor U734 (N_734,In_974,In_1937);
and U735 (N_735,In_797,N_355);
nor U736 (N_736,In_715,N_361);
and U737 (N_737,In_453,In_259);
or U738 (N_738,N_10,N_94);
nand U739 (N_739,N_216,N_329);
nor U740 (N_740,In_677,In_1572);
or U741 (N_741,In_158,N_478);
nand U742 (N_742,In_535,N_291);
and U743 (N_743,In_753,In_1116);
nor U744 (N_744,In_1853,In_66);
or U745 (N_745,In_1048,In_834);
or U746 (N_746,N_232,In_1652);
xnor U747 (N_747,In_1805,N_226);
nand U748 (N_748,In_849,In_1778);
and U749 (N_749,N_468,In_1018);
and U750 (N_750,In_1834,In_1399);
nor U751 (N_751,N_0,In_1303);
or U752 (N_752,In_1466,N_23);
xor U753 (N_753,N_442,In_332);
nor U754 (N_754,In_482,N_344);
or U755 (N_755,N_22,In_279);
nor U756 (N_756,In_967,In_1850);
xnor U757 (N_757,In_1732,In_1901);
nor U758 (N_758,N_317,N_261);
nand U759 (N_759,N_241,In_461);
nand U760 (N_760,N_371,In_1062);
or U761 (N_761,N_108,N_290);
nand U762 (N_762,N_374,N_43);
nor U763 (N_763,In_1369,In_958);
xor U764 (N_764,In_399,N_67);
or U765 (N_765,In_1424,In_568);
nor U766 (N_766,N_301,In_1286);
and U767 (N_767,N_166,N_129);
nand U768 (N_768,In_1586,In_286);
nor U769 (N_769,In_228,In_1528);
or U770 (N_770,In_1149,In_1742);
xnor U771 (N_771,In_451,N_459);
or U772 (N_772,N_496,N_83);
nand U773 (N_773,In_318,N_244);
or U774 (N_774,In_1271,In_1534);
and U775 (N_775,In_1119,N_297);
and U776 (N_776,In_236,In_180);
nor U777 (N_777,In_1683,In_661);
or U778 (N_778,In_185,In_1502);
or U779 (N_779,In_1818,N_121);
nand U780 (N_780,In_162,In_1738);
and U781 (N_781,N_135,In_1401);
nand U782 (N_782,In_425,In_1101);
and U783 (N_783,In_1936,In_1681);
nand U784 (N_784,In_547,N_440);
and U785 (N_785,In_149,N_2);
and U786 (N_786,In_572,In_898);
nand U787 (N_787,In_1851,In_1126);
xor U788 (N_788,In_630,N_54);
nor U789 (N_789,In_1163,In_525);
or U790 (N_790,N_18,In_1837);
nand U791 (N_791,In_1935,In_1475);
and U792 (N_792,N_1,In_1293);
nand U793 (N_793,N_382,In_1095);
xnor U794 (N_794,N_404,In_768);
or U795 (N_795,In_827,In_1228);
xnor U796 (N_796,In_44,In_370);
and U797 (N_797,In_986,In_1857);
and U798 (N_798,In_515,In_1020);
or U799 (N_799,In_1548,N_120);
nand U800 (N_800,In_529,N_61);
or U801 (N_801,N_288,In_519);
and U802 (N_802,N_342,In_330);
nand U803 (N_803,In_248,In_137);
or U804 (N_804,In_772,In_731);
nor U805 (N_805,N_354,N_462);
nand U806 (N_806,In_92,In_1989);
and U807 (N_807,N_64,N_51);
xor U808 (N_808,N_42,In_1240);
and U809 (N_809,N_81,N_190);
or U810 (N_810,N_263,N_375);
nor U811 (N_811,In_348,In_1634);
nor U812 (N_812,In_405,N_126);
nor U813 (N_813,N_9,N_30);
xnor U814 (N_814,In_1661,In_1625);
xnor U815 (N_815,In_1397,In_1490);
xnor U816 (N_816,In_1999,In_1146);
and U817 (N_817,In_1987,N_262);
nand U818 (N_818,N_408,In_1154);
nand U819 (N_819,N_321,In_314);
or U820 (N_820,In_809,In_467);
or U821 (N_821,In_354,In_956);
nor U822 (N_822,In_1434,In_1402);
nor U823 (N_823,In_1856,In_63);
and U824 (N_824,N_259,N_12);
nor U825 (N_825,In_121,In_1232);
nor U826 (N_826,N_434,N_66);
xnor U827 (N_827,N_490,In_775);
xor U828 (N_828,In_325,In_638);
and U829 (N_829,In_851,In_1105);
and U830 (N_830,In_1435,In_1794);
and U831 (N_831,N_341,In_1);
nand U832 (N_832,N_487,In_216);
or U833 (N_833,In_1607,N_53);
or U834 (N_834,In_729,N_56);
nor U835 (N_835,In_978,In_651);
nor U836 (N_836,N_286,N_353);
nand U837 (N_837,In_1115,In_1564);
or U838 (N_838,In_1496,In_1107);
nand U839 (N_839,In_1097,N_138);
or U840 (N_840,In_629,In_230);
and U841 (N_841,In_1638,In_659);
nand U842 (N_842,In_1667,N_451);
or U843 (N_843,In_493,N_44);
and U844 (N_844,In_953,N_223);
nand U845 (N_845,In_276,N_454);
or U846 (N_846,In_1905,N_266);
xor U847 (N_847,In_159,In_1715);
and U848 (N_848,In_91,In_690);
or U849 (N_849,N_70,In_675);
nor U850 (N_850,In_268,In_465);
nor U851 (N_851,In_933,In_1522);
nand U852 (N_852,N_230,N_489);
and U853 (N_853,N_427,In_1967);
nor U854 (N_854,N_205,In_726);
and U855 (N_855,In_1225,In_1505);
nand U856 (N_856,In_1747,N_445);
and U857 (N_857,N_187,N_41);
or U858 (N_858,N_295,N_398);
nand U859 (N_859,In_1875,In_647);
nand U860 (N_860,N_106,In_499);
xor U861 (N_861,N_122,In_821);
nor U862 (N_862,In_265,N_160);
xnor U863 (N_863,In_1056,In_1497);
xor U864 (N_864,In_912,In_352);
xnor U865 (N_865,N_304,In_1914);
nand U866 (N_866,In_1943,In_531);
xor U867 (N_867,In_367,N_335);
xnor U868 (N_868,In_210,N_7);
nand U869 (N_869,N_473,In_1513);
or U870 (N_870,N_247,In_1442);
and U871 (N_871,In_1214,In_1793);
and U872 (N_872,N_379,In_698);
xnor U873 (N_873,In_1368,N_165);
nand U874 (N_874,N_173,N_275);
and U875 (N_875,N_91,In_1448);
or U876 (N_876,In_622,In_1089);
or U877 (N_877,In_634,In_940);
nand U878 (N_878,N_158,In_198);
nand U879 (N_879,In_960,In_1651);
and U880 (N_880,In_891,In_398);
nor U881 (N_881,In_1400,N_225);
xnor U882 (N_882,In_648,N_277);
or U883 (N_883,In_1375,N_153);
nand U884 (N_884,In_1756,In_282);
xnor U885 (N_885,N_491,In_1403);
nand U886 (N_886,In_1627,N_274);
nand U887 (N_887,In_557,N_45);
nor U888 (N_888,N_394,N_483);
xnor U889 (N_889,In_728,N_250);
or U890 (N_890,N_400,In_577);
nor U891 (N_891,In_35,In_1226);
xor U892 (N_892,N_298,In_566);
nor U893 (N_893,In_1541,In_68);
xnor U894 (N_894,In_511,In_494);
xnor U895 (N_895,In_730,In_801);
nand U896 (N_896,In_389,N_320);
nor U897 (N_897,In_1235,In_1082);
and U898 (N_898,In_34,N_357);
and U899 (N_899,In_490,In_1414);
nand U900 (N_900,N_425,N_437);
and U901 (N_901,N_86,In_483);
nand U902 (N_902,N_219,In_798);
or U903 (N_903,N_218,In_914);
nand U904 (N_904,N_364,In_1015);
nor U905 (N_905,In_1110,In_1313);
and U906 (N_906,In_778,N_369);
or U907 (N_907,N_28,N_299);
or U908 (N_908,In_870,In_1471);
and U909 (N_909,In_576,In_193);
xor U910 (N_910,In_803,N_239);
nand U911 (N_911,In_1450,In_1689);
xor U912 (N_912,In_1817,N_6);
and U913 (N_913,N_306,In_202);
nand U914 (N_914,N_424,N_157);
and U915 (N_915,In_1456,In_1109);
xor U916 (N_916,N_377,In_1298);
xor U917 (N_917,In_197,N_412);
nand U918 (N_918,In_580,N_240);
nor U919 (N_919,N_124,N_235);
or U920 (N_920,In_1367,In_1136);
and U921 (N_921,In_1862,In_1664);
nand U922 (N_922,In_1437,In_1241);
nor U923 (N_923,N_416,In_1026);
xor U924 (N_924,In_1819,In_968);
nand U925 (N_925,In_628,N_231);
nand U926 (N_926,In_883,In_673);
or U927 (N_927,In_1531,N_183);
and U928 (N_928,In_4,In_1612);
nor U929 (N_929,In_402,In_28);
xor U930 (N_930,N_333,In_645);
nor U931 (N_931,In_1438,In_1899);
xor U932 (N_932,N_104,In_289);
and U933 (N_933,In_793,In_1641);
and U934 (N_934,In_736,In_796);
nand U935 (N_935,In_344,In_1174);
nor U936 (N_936,In_435,In_261);
xor U937 (N_937,In_764,In_1393);
nand U938 (N_938,In_1500,In_1196);
or U939 (N_939,N_99,N_75);
xnor U940 (N_940,N_55,In_1693);
nor U941 (N_941,In_1207,In_1822);
and U942 (N_942,In_1337,In_116);
nand U943 (N_943,In_1387,In_1257);
nand U944 (N_944,In_1304,N_170);
xor U945 (N_945,N_85,N_347);
nand U946 (N_946,In_1569,In_1431);
or U947 (N_947,In_1730,N_267);
nand U948 (N_948,In_1045,N_109);
xor U949 (N_949,In_838,In_907);
nor U950 (N_950,In_271,In_1059);
xnor U951 (N_951,In_119,In_1960);
nand U952 (N_952,N_363,In_765);
xnor U953 (N_953,In_1719,In_473);
xor U954 (N_954,N_242,In_733);
or U955 (N_955,N_270,N_116);
nor U956 (N_956,N_284,In_616);
and U957 (N_957,N_326,In_1731);
xnor U958 (N_958,In_971,N_340);
or U959 (N_959,In_789,In_206);
or U960 (N_960,In_1205,N_103);
or U961 (N_961,N_176,In_264);
or U962 (N_962,In_1965,N_155);
and U963 (N_963,N_352,In_130);
nor U964 (N_964,N_47,In_316);
nand U965 (N_965,In_526,N_20);
nor U966 (N_966,N_438,In_1485);
nor U967 (N_967,In_1384,In_1780);
nand U968 (N_968,In_94,In_814);
nor U969 (N_969,In_552,In_1838);
xnor U970 (N_970,In_439,In_1783);
and U971 (N_971,In_1480,In_1195);
or U972 (N_972,N_101,N_407);
or U973 (N_973,In_1483,N_204);
and U974 (N_974,N_164,In_1984);
and U975 (N_975,In_240,In_1698);
nor U976 (N_976,In_599,In_1969);
xnor U977 (N_977,In_934,In_65);
nand U978 (N_978,In_1268,In_969);
nor U979 (N_979,N_137,In_98);
nand U980 (N_980,In_1718,N_80);
nand U981 (N_981,In_131,In_1336);
xor U982 (N_982,In_1342,In_1217);
xor U983 (N_983,N_193,In_595);
nand U984 (N_984,In_836,N_131);
and U985 (N_985,N_97,In_991);
xnor U986 (N_986,In_33,In_1263);
nor U987 (N_987,In_649,In_691);
xnor U988 (N_988,In_1316,N_161);
nand U989 (N_989,N_495,In_1291);
nor U990 (N_990,In_681,In_623);
or U991 (N_991,In_1162,In_1888);
nand U992 (N_992,In_512,N_234);
nor U993 (N_993,In_507,In_1789);
nand U994 (N_994,N_309,In_160);
xnor U995 (N_995,In_5,In_376);
or U996 (N_996,In_88,N_467);
or U997 (N_997,In_1150,In_1951);
or U998 (N_998,N_198,In_888);
nand U999 (N_999,N_313,In_788);
nor U1000 (N_1000,N_982,In_545);
xnor U1001 (N_1001,N_908,N_791);
and U1002 (N_1002,In_152,N_800);
xor U1003 (N_1003,In_980,In_1896);
xor U1004 (N_1004,N_710,N_24);
xnor U1005 (N_1005,N_779,N_732);
xor U1006 (N_1006,N_759,In_984);
nand U1007 (N_1007,In_227,N_946);
nand U1008 (N_1008,N_646,N_228);
xor U1009 (N_1009,N_337,N_849);
or U1010 (N_1010,N_415,N_885);
and U1011 (N_1011,N_620,N_550);
and U1012 (N_1012,In_1135,N_786);
xor U1013 (N_1013,In_1357,In_1389);
nand U1014 (N_1014,N_773,N_544);
nand U1015 (N_1015,In_110,In_1113);
and U1016 (N_1016,In_1084,N_698);
xor U1017 (N_1017,N_650,N_76);
and U1018 (N_1018,N_962,N_582);
xor U1019 (N_1019,N_639,N_411);
and U1020 (N_1020,N_785,N_995);
xnor U1021 (N_1021,N_568,N_50);
nor U1022 (N_1022,N_203,In_543);
and U1023 (N_1023,In_191,N_324);
nand U1024 (N_1024,In_1383,N_963);
xor U1025 (N_1025,In_205,N_644);
nor U1026 (N_1026,N_551,In_1461);
or U1027 (N_1027,In_15,N_713);
xnor U1028 (N_1028,N_747,N_906);
xor U1029 (N_1029,In_955,In_141);
nor U1030 (N_1030,N_706,N_629);
nor U1031 (N_1031,N_742,In_1171);
nor U1032 (N_1032,N_148,N_115);
xor U1033 (N_1033,N_889,N_770);
nand U1034 (N_1034,In_1669,N_303);
nor U1035 (N_1035,N_986,In_1766);
or U1036 (N_1036,N_678,N_621);
or U1037 (N_1037,N_192,N_769);
or U1038 (N_1038,N_359,N_702);
nand U1039 (N_1039,N_622,N_824);
nor U1040 (N_1040,In_1409,N_565);
and U1041 (N_1041,N_676,N_826);
xnor U1042 (N_1042,N_850,In_643);
nand U1043 (N_1043,In_460,In_1706);
and U1044 (N_1044,N_971,N_979);
xor U1045 (N_1045,N_127,N_147);
xnor U1046 (N_1046,In_383,In_1139);
xor U1047 (N_1047,N_739,In_1581);
and U1048 (N_1048,N_527,N_662);
xor U1049 (N_1049,In_225,N_977);
xnor U1050 (N_1050,N_588,N_859);
or U1051 (N_1051,In_799,In_1043);
xor U1052 (N_1052,In_32,In_251);
nor U1053 (N_1053,N_877,N_546);
and U1054 (N_1054,N_510,N_422);
nand U1055 (N_1055,In_779,N_926);
and U1056 (N_1056,In_597,In_508);
nand U1057 (N_1057,N_776,N_664);
and U1058 (N_1058,N_883,In_1388);
and U1059 (N_1059,N_822,N_512);
nand U1060 (N_1060,N_924,N_34);
nand U1061 (N_1061,N_938,In_1804);
or U1062 (N_1062,N_370,In_1644);
xnor U1063 (N_1063,N_925,N_852);
nor U1064 (N_1064,N_923,N_870);
xor U1065 (N_1065,In_243,N_488);
or U1066 (N_1066,N_874,N_456);
nor U1067 (N_1067,In_76,N_878);
nor U1068 (N_1068,In_1177,In_929);
and U1069 (N_1069,In_866,In_1075);
nor U1070 (N_1070,N_450,In_558);
nor U1071 (N_1071,N_180,N_757);
xor U1072 (N_1072,N_222,In_646);
nand U1073 (N_1073,In_819,In_440);
xor U1074 (N_1074,In_1042,N_33);
or U1075 (N_1075,N_111,N_145);
and U1076 (N_1076,N_672,N_990);
or U1077 (N_1077,N_827,N_500);
and U1078 (N_1078,N_853,N_452);
nand U1079 (N_1079,In_1233,N_820);
and U1080 (N_1080,N_915,N_981);
or U1081 (N_1081,N_559,N_300);
nand U1082 (N_1082,N_720,N_681);
or U1083 (N_1083,In_381,N_579);
nand U1084 (N_1084,In_1553,N_433);
nor U1085 (N_1085,N_89,In_1639);
nor U1086 (N_1086,N_934,N_760);
or U1087 (N_1087,N_688,In_624);
nor U1088 (N_1088,N_252,N_677);
xnor U1089 (N_1089,In_338,In_1352);
or U1090 (N_1090,N_139,In_1390);
and U1091 (N_1091,In_1165,N_736);
nor U1092 (N_1092,In_1761,N_403);
xor U1093 (N_1093,N_756,N_17);
nand U1094 (N_1094,N_631,In_975);
xor U1095 (N_1095,N_470,N_789);
or U1096 (N_1096,N_236,N_632);
or U1097 (N_1097,In_1279,In_255);
or U1098 (N_1098,In_317,In_1354);
xor U1099 (N_1099,N_969,N_944);
nand U1100 (N_1100,N_207,N_817);
or U1101 (N_1101,N_593,N_77);
nor U1102 (N_1102,N_767,N_577);
xor U1103 (N_1103,N_538,N_911);
and U1104 (N_1104,N_685,In_817);
nand U1105 (N_1105,In_239,In_1457);
or U1106 (N_1106,N_684,In_1876);
and U1107 (N_1107,N_768,N_848);
xnor U1108 (N_1108,N_525,N_802);
nand U1109 (N_1109,In_1266,N_366);
nor U1110 (N_1110,N_692,N_932);
nand U1111 (N_1111,In_81,In_1567);
nand U1112 (N_1112,N_587,N_953);
nand U1113 (N_1113,In_1527,In_1808);
or U1114 (N_1114,In_1327,N_673);
nor U1115 (N_1115,N_507,N_741);
and U1116 (N_1116,In_257,In_115);
and U1117 (N_1117,N_952,N_46);
or U1118 (N_1118,In_1260,N_256);
nand U1119 (N_1119,In_1589,In_908);
nand U1120 (N_1120,In_1826,In_1022);
nand U1121 (N_1121,N_516,N_560);
nand U1122 (N_1122,In_400,In_668);
nor U1123 (N_1123,N_169,N_188);
and U1124 (N_1124,N_987,N_968);
or U1125 (N_1125,In_327,N_947);
or U1126 (N_1126,N_807,N_133);
nand U1127 (N_1127,N_573,N_994);
or U1128 (N_1128,N_502,N_536);
nand U1129 (N_1129,N_787,N_530);
xnor U1130 (N_1130,In_377,N_647);
xnor U1131 (N_1131,N_323,N_809);
xnor U1132 (N_1132,In_1986,N_888);
and U1133 (N_1133,N_567,N_49);
xor U1134 (N_1134,N_73,N_998);
xnor U1135 (N_1135,In_770,N_976);
xor U1136 (N_1136,N_945,N_322);
nor U1137 (N_1137,N_199,N_197);
nor U1138 (N_1138,N_195,In_1102);
nor U1139 (N_1139,N_144,N_113);
and U1140 (N_1140,In_1708,In_1307);
and U1141 (N_1141,In_495,N_522);
or U1142 (N_1142,In_1079,N_754);
nand U1143 (N_1143,N_746,N_726);
and U1144 (N_1144,N_993,N_397);
or U1145 (N_1145,In_1668,N_856);
or U1146 (N_1146,In_1238,N_542);
nor U1147 (N_1147,N_380,N_956);
nor U1148 (N_1148,In_1744,In_1132);
and U1149 (N_1149,N_740,In_1184);
nor U1150 (N_1150,In_1248,N_618);
or U1151 (N_1151,In_1151,In_602);
or U1152 (N_1152,N_584,N_771);
or U1153 (N_1153,In_1458,N_253);
xor U1154 (N_1154,In_1663,N_814);
or U1155 (N_1155,In_1242,N_890);
xnor U1156 (N_1156,N_294,N_117);
nor U1157 (N_1157,N_520,N_737);
or U1158 (N_1158,N_583,N_795);
nor U1159 (N_1159,N_832,In_1750);
nand U1160 (N_1160,N_655,N_130);
nand U1161 (N_1161,In_40,N_634);
or U1162 (N_1162,N_918,N_928);
xor U1163 (N_1163,In_1507,In_403);
nor U1164 (N_1164,N_803,N_237);
xor U1165 (N_1165,N_661,N_16);
xor U1166 (N_1166,N_606,N_59);
and U1167 (N_1167,In_1889,In_1716);
and U1168 (N_1168,N_186,In_1629);
nor U1169 (N_1169,In_18,N_863);
nand U1170 (N_1170,N_873,N_917);
and U1171 (N_1171,In_1938,N_989);
or U1172 (N_1172,N_914,N_654);
and U1173 (N_1173,In_1038,N_886);
nand U1174 (N_1174,In_280,In_138);
xnor U1175 (N_1175,N_87,N_959);
and U1176 (N_1176,In_948,N_703);
nor U1177 (N_1177,N_174,In_1017);
nand U1178 (N_1178,N_973,N_141);
xor U1179 (N_1179,N_966,N_841);
nor U1180 (N_1180,N_282,In_800);
nand U1181 (N_1181,N_901,N_838);
and U1182 (N_1182,N_781,In_1019);
and U1183 (N_1183,N_858,N_640);
xor U1184 (N_1184,In_1917,N_864);
nand U1185 (N_1185,N_338,N_52);
and U1186 (N_1186,In_574,N_682);
nand U1187 (N_1187,N_576,N_506);
or U1188 (N_1188,N_605,N_920);
or U1189 (N_1189,N_997,N_553);
nor U1190 (N_1190,In_804,N_964);
and U1191 (N_1191,N_784,In_144);
and U1192 (N_1192,In_1091,N_764);
or U1193 (N_1193,In_875,In_911);
nor U1194 (N_1194,N_978,N_880);
xor U1195 (N_1195,In_1321,In_1439);
or U1196 (N_1196,N_327,N_733);
or U1197 (N_1197,In_1158,N_669);
xnor U1198 (N_1198,N_816,In_787);
or U1199 (N_1199,N_229,In_720);
nor U1200 (N_1200,In_472,N_447);
or U1201 (N_1201,N_750,N_302);
nor U1202 (N_1202,N_515,N_819);
and U1203 (N_1203,N_929,N_700);
nor U1204 (N_1204,N_735,In_272);
nand U1205 (N_1205,N_941,In_269);
and U1206 (N_1206,N_721,In_714);
nor U1207 (N_1207,In_1604,In_1155);
xor U1208 (N_1208,N_558,In_1635);
nand U1209 (N_1209,In_62,In_320);
and U1210 (N_1210,N_666,In_604);
xnor U1211 (N_1211,N_724,N_260);
or U1212 (N_1212,N_690,N_608);
and U1213 (N_1213,N_694,N_460);
nand U1214 (N_1214,In_1658,N_948);
xor U1215 (N_1215,N_611,In_1323);
nor U1216 (N_1216,N_540,N_566);
nand U1217 (N_1217,In_1333,N_991);
xor U1218 (N_1218,In_1556,N_179);
and U1219 (N_1219,N_796,N_931);
nor U1220 (N_1220,N_815,N_102);
xor U1221 (N_1221,N_701,N_257);
nor U1222 (N_1222,N_813,In_1346);
xnor U1223 (N_1223,In_721,N_69);
nor U1224 (N_1224,In_725,N_143);
nand U1225 (N_1225,In_1054,In_699);
nand U1226 (N_1226,N_630,N_896);
or U1227 (N_1227,N_716,In_1094);
or U1228 (N_1228,N_389,N_868);
and U1229 (N_1229,N_867,N_182);
xor U1230 (N_1230,N_312,In_635);
xor U1231 (N_1231,N_482,N_835);
nor U1232 (N_1232,In_1194,N_825);
and U1233 (N_1233,N_752,In_1666);
nor U1234 (N_1234,N_604,In_1272);
or U1235 (N_1235,N_774,In_1878);
nand U1236 (N_1236,N_935,In_319);
xnor U1237 (N_1237,N_163,N_649);
or U1238 (N_1238,In_1831,In_480);
and U1239 (N_1239,N_351,N_665);
or U1240 (N_1240,N_903,N_823);
nand U1241 (N_1241,In_952,In_1953);
or U1242 (N_1242,In_1551,N_78);
or U1243 (N_1243,In_1723,N_248);
and U1244 (N_1244,N_900,N_999);
nand U1245 (N_1245,N_727,In_1792);
nor U1246 (N_1246,N_25,N_725);
nand U1247 (N_1247,N_589,In_176);
nand U1248 (N_1248,In_1455,N_758);
nand U1249 (N_1249,In_569,N_638);
nand U1250 (N_1250,N_348,N_580);
xor U1251 (N_1251,N_578,N_992);
or U1252 (N_1252,N_851,N_818);
nor U1253 (N_1253,N_658,N_32);
and U1254 (N_1254,N_40,N_569);
nor U1255 (N_1255,N_719,N_775);
and U1256 (N_1256,N_381,N_350);
nand U1257 (N_1257,N_475,In_1278);
or U1258 (N_1258,N_591,N_937);
nor U1259 (N_1259,N_575,N_722);
or U1260 (N_1260,In_1070,N_140);
or U1261 (N_1261,In_454,N_603);
nand U1262 (N_1262,In_1835,N_596);
and U1263 (N_1263,N_533,In_3);
and U1264 (N_1264,In_845,N_613);
or U1265 (N_1265,In_438,N_793);
xor U1266 (N_1266,In_1033,In_981);
nor U1267 (N_1267,N_975,N_547);
or U1268 (N_1268,N_610,N_879);
nor U1269 (N_1269,In_925,In_560);
and U1270 (N_1270,N_927,In_1498);
xor U1271 (N_1271,N_829,N_477);
or U1272 (N_1272,N_633,N_704);
xor U1273 (N_1273,N_891,N_892);
and U1274 (N_1274,N_955,N_783);
nor U1275 (N_1275,N_810,N_555);
and U1276 (N_1276,N_919,In_211);
or U1277 (N_1277,N_532,N_529);
and U1278 (N_1278,N_950,N_523);
and U1279 (N_1279,N_36,In_157);
or U1280 (N_1280,N_519,N_461);
and U1281 (N_1281,In_1172,In_1568);
xor U1282 (N_1282,N_612,N_499);
and U1283 (N_1283,In_1479,In_226);
and U1284 (N_1284,N_882,N_872);
or U1285 (N_1285,N_562,N_687);
nor U1286 (N_1286,N_278,In_880);
nor U1287 (N_1287,N_680,N_146);
or U1288 (N_1288,N_281,N_432);
nor U1289 (N_1289,N_862,N_730);
xor U1290 (N_1290,N_524,In_1679);
or U1291 (N_1291,In_1970,In_1621);
nand U1292 (N_1292,In_697,In_1973);
or U1293 (N_1293,In_1000,In_1270);
xor U1294 (N_1294,In_1259,N_696);
xnor U1295 (N_1295,In_278,N_561);
and U1296 (N_1296,N_902,N_623);
xor U1297 (N_1297,N_15,N_899);
nor U1298 (N_1298,In_664,N_939);
nand U1299 (N_1299,N_942,N_745);
nor U1300 (N_1300,N_834,N_233);
nor U1301 (N_1301,In_660,N_196);
xnor U1302 (N_1302,N_907,In_957);
nand U1303 (N_1303,N_125,In_1585);
xor U1304 (N_1304,N_695,In_909);
and U1305 (N_1305,N_548,N_686);
or U1306 (N_1306,N_659,In_1932);
or U1307 (N_1307,In_414,N_731);
nand U1308 (N_1308,N_390,N_714);
nand U1309 (N_1309,In_926,N_861);
xor U1310 (N_1310,N_980,In_1472);
and U1311 (N_1311,N_586,In_863);
xor U1312 (N_1312,N_884,In_1118);
and U1313 (N_1313,In_1003,N_554);
nand U1314 (N_1314,N_844,N_636);
and U1315 (N_1315,N_689,N_373);
nor U1316 (N_1316,In_223,In_433);
or U1317 (N_1317,N_840,N_961);
nand U1318 (N_1318,N_152,N_693);
and U1319 (N_1319,N_799,N_642);
nor U1320 (N_1320,N_794,In_707);
or U1321 (N_1321,In_1530,N_431);
nor U1322 (N_1322,N_656,N_396);
nor U1323 (N_1323,In_30,N_843);
and U1324 (N_1324,N_660,N_110);
and U1325 (N_1325,N_806,In_1636);
or U1326 (N_1326,N_585,N_857);
and U1327 (N_1327,N_675,N_189);
and U1328 (N_1328,N_276,N_895);
nand U1329 (N_1329,In_139,N_641);
nand U1330 (N_1330,N_913,In_1785);
xor U1331 (N_1331,In_1672,N_13);
and U1332 (N_1332,In_1425,N_602);
xnor U1333 (N_1333,N_831,N_833);
or U1334 (N_1334,In_1782,N_763);
or U1335 (N_1335,In_365,In_164);
xnor U1336 (N_1336,In_1236,In_1009);
and U1337 (N_1337,In_340,In_947);
nand U1338 (N_1338,N_805,In_618);
or U1339 (N_1339,N_691,N_905);
xnor U1340 (N_1340,In_39,In_774);
or U1341 (N_1341,N_571,In_1061);
nor U1342 (N_1342,N_921,In_862);
xor U1343 (N_1343,N_985,N_984);
nand U1344 (N_1344,N_869,N_974);
xor U1345 (N_1345,N_951,N_916);
and U1346 (N_1346,N_607,In_1904);
nor U1347 (N_1347,N_777,N_526);
and U1348 (N_1348,In_1460,N_539);
xor U1349 (N_1349,In_1928,N_683);
xnor U1350 (N_1350,N_811,In_1051);
and U1351 (N_1351,N_755,In_588);
and U1352 (N_1352,In_842,In_1949);
nand U1353 (N_1353,N_821,N_797);
nand U1354 (N_1354,N_581,N_528);
and U1355 (N_1355,N_808,N_513);
xor U1356 (N_1356,N_556,N_699);
nor U1357 (N_1357,In_826,In_1799);
or U1358 (N_1358,N_210,In_1365);
nor U1359 (N_1359,N_667,In_848);
xnor U1360 (N_1360,N_729,N_455);
and U1361 (N_1361,N_423,N_983);
nor U1362 (N_1362,N_534,In_1843);
nand U1363 (N_1363,In_274,N_712);
xnor U1364 (N_1364,N_904,N_887);
nand U1365 (N_1365,In_928,N_875);
and U1366 (N_1366,N_616,N_378);
and U1367 (N_1367,N_871,N_609);
nand U1368 (N_1368,N_893,In_1353);
nand U1369 (N_1369,In_970,N_625);
and U1370 (N_1370,N_778,N_940);
nand U1371 (N_1371,N_521,In_514);
nor U1372 (N_1372,In_608,N_480);
and U1373 (N_1373,In_1828,N_386);
or U1374 (N_1374,In_1645,N_57);
and U1375 (N_1375,In_830,N_508);
or U1376 (N_1376,N_846,In_60);
nand U1377 (N_1377,In_151,N_563);
and U1378 (N_1378,In_1867,In_1535);
nand U1379 (N_1379,In_1133,In_1566);
nand U1380 (N_1380,N_458,N_464);
xor U1381 (N_1381,N_325,In_245);
nand U1382 (N_1382,N_909,In_706);
or U1383 (N_1383,In_1300,N_707);
and U1384 (N_1384,N_854,N_628);
and U1385 (N_1385,N_504,In_322);
nor U1386 (N_1386,N_782,N_367);
nand U1387 (N_1387,N_762,N_648);
xnor U1388 (N_1388,N_549,N_498);
and U1389 (N_1389,In_1131,N_272);
nor U1390 (N_1390,N_705,N_828);
nand U1391 (N_1391,N_365,In_1301);
and U1392 (N_1392,N_624,N_635);
xor U1393 (N_1393,N_744,N_511);
or U1394 (N_1394,N_29,In_1873);
xor U1395 (N_1395,N_493,N_600);
and U1396 (N_1396,In_61,N_501);
xnor U1397 (N_1397,In_1487,N_211);
or U1398 (N_1398,N_409,In_1622);
nor U1399 (N_1399,N_418,N_328);
or U1400 (N_1400,N_598,N_788);
xnor U1401 (N_1401,N_936,N_972);
nor U1402 (N_1402,N_619,N_38);
nor U1403 (N_1403,N_615,N_202);
or U1404 (N_1404,N_651,N_564);
and U1405 (N_1405,N_283,N_200);
nand U1406 (N_1406,N_715,In_1562);
nand U1407 (N_1407,In_1677,N_595);
and U1408 (N_1408,In_1044,In_751);
nand U1409 (N_1409,N_457,In_38);
xor U1410 (N_1410,N_592,N_517);
and U1411 (N_1411,N_711,In_1322);
and U1412 (N_1412,N_761,N_224);
and U1413 (N_1413,N_765,N_123);
nor U1414 (N_1414,N_749,In_989);
xnor U1415 (N_1415,N_162,N_792);
nor U1416 (N_1416,N_743,N_356);
nor U1417 (N_1417,N_531,N_537);
and U1418 (N_1418,In_1962,In_853);
xnor U1419 (N_1419,In_859,In_1378);
or U1420 (N_1420,In_1811,N_100);
or U1421 (N_1421,In_295,N_922);
and U1422 (N_1422,N_967,N_264);
and U1423 (N_1423,In_1746,N_599);
and U1424 (N_1424,N_541,N_855);
and U1425 (N_1425,N_697,N_866);
and U1426 (N_1426,N_842,In_114);
nand U1427 (N_1427,N_865,N_134);
or U1428 (N_1428,In_437,In_1927);
nor U1429 (N_1429,N_943,N_790);
or U1430 (N_1430,N_753,N_860);
nand U1431 (N_1431,In_1729,N_717);
or U1432 (N_1432,N_751,N_626);
xnor U1433 (N_1433,N_679,N_912);
nand U1434 (N_1434,In_1674,N_545);
or U1435 (N_1435,N_574,N_960);
and U1436 (N_1436,In_1559,N_594);
nor U1437 (N_1437,N_268,In_752);
nor U1438 (N_1438,In_1212,N_876);
nand U1439 (N_1439,N_535,N_670);
xnor U1440 (N_1440,N_748,In_973);
nand U1441 (N_1441,N_191,N_552);
or U1442 (N_1442,N_177,N_898);
or U1443 (N_1443,N_723,N_954);
nor U1444 (N_1444,N_627,In_11);
and U1445 (N_1445,N_503,N_709);
nor U1446 (N_1446,In_1576,N_652);
and U1447 (N_1447,N_988,N_839);
nand U1448 (N_1448,N_772,In_424);
nor U1449 (N_1449,N_663,In_83);
nand U1450 (N_1450,N_590,N_336);
and U1451 (N_1451,N_597,In_1210);
xor U1452 (N_1452,N_801,N_668);
and U1453 (N_1453,N_804,N_965);
or U1454 (N_1454,N_766,In_1704);
and U1455 (N_1455,N_514,N_718);
xor U1456 (N_1456,N_798,In_43);
nand U1457 (N_1457,In_1494,N_410);
and U1458 (N_1458,In_1881,In_462);
or U1459 (N_1459,N_505,In_1234);
xnor U1460 (N_1460,N_637,N_812);
or U1461 (N_1461,N_444,N_957);
nand U1462 (N_1462,N_881,N_657);
and U1463 (N_1463,N_933,N_830);
nor U1464 (N_1464,N_836,N_728);
and U1465 (N_1465,N_128,N_572);
xnor U1466 (N_1466,In_1440,N_98);
nor U1467 (N_1467,N_958,N_557);
nor U1468 (N_1468,N_308,In_1370);
and U1469 (N_1469,In_935,N_653);
nor U1470 (N_1470,N_894,N_614);
nand U1471 (N_1471,N_292,In_477);
xnor U1472 (N_1472,N_996,N_601);
nor U1473 (N_1473,N_671,In_581);
nor U1474 (N_1474,In_1239,N_154);
nand U1475 (N_1475,In_469,N_543);
and U1476 (N_1476,N_167,In_976);
xor U1477 (N_1477,N_897,N_384);
nor U1478 (N_1478,In_962,In_363);
nor U1479 (N_1479,In_1222,N_738);
xor U1480 (N_1480,N_674,In_1348);
and U1481 (N_1481,In_1221,In_1080);
and U1482 (N_1482,N_837,N_518);
and U1483 (N_1483,In_1275,N_910);
or U1484 (N_1484,In_1122,N_314);
xor U1485 (N_1485,N_645,In_21);
nor U1486 (N_1486,N_847,In_944);
or U1487 (N_1487,N_509,N_780);
or U1488 (N_1488,N_265,N_970);
nand U1489 (N_1489,In_1134,In_1201);
and U1490 (N_1490,N_570,N_213);
nor U1491 (N_1491,N_168,N_617);
and U1492 (N_1492,N_159,N_845);
xor U1493 (N_1493,In_359,N_930);
nor U1494 (N_1494,N_494,In_393);
xnor U1495 (N_1495,In_179,In_1590);
nand U1496 (N_1496,In_429,N_643);
xnor U1497 (N_1497,N_949,In_1104);
or U1498 (N_1498,In_1721,In_1648);
xnor U1499 (N_1499,N_734,N_708);
nor U1500 (N_1500,N_1155,N_1383);
or U1501 (N_1501,N_1231,N_1330);
nor U1502 (N_1502,N_1176,N_1397);
nor U1503 (N_1503,N_1360,N_1237);
nor U1504 (N_1504,N_1484,N_1347);
and U1505 (N_1505,N_1234,N_1499);
and U1506 (N_1506,N_1122,N_1151);
xnor U1507 (N_1507,N_1346,N_1097);
xor U1508 (N_1508,N_1281,N_1453);
nand U1509 (N_1509,N_1295,N_1195);
nand U1510 (N_1510,N_1404,N_1197);
nor U1511 (N_1511,N_1171,N_1389);
nor U1512 (N_1512,N_1180,N_1410);
xnor U1513 (N_1513,N_1233,N_1049);
nor U1514 (N_1514,N_1487,N_1370);
and U1515 (N_1515,N_1223,N_1392);
nand U1516 (N_1516,N_1262,N_1343);
or U1517 (N_1517,N_1304,N_1002);
nand U1518 (N_1518,N_1057,N_1078);
xor U1519 (N_1519,N_1293,N_1428);
nor U1520 (N_1520,N_1104,N_1110);
nand U1521 (N_1521,N_1280,N_1378);
or U1522 (N_1522,N_1296,N_1429);
xor U1523 (N_1523,N_1124,N_1481);
nor U1524 (N_1524,N_1163,N_1433);
and U1525 (N_1525,N_1409,N_1339);
nor U1526 (N_1526,N_1337,N_1322);
or U1527 (N_1527,N_1201,N_1353);
nor U1528 (N_1528,N_1047,N_1158);
nand U1529 (N_1529,N_1417,N_1006);
nor U1530 (N_1530,N_1044,N_1040);
nor U1531 (N_1531,N_1270,N_1113);
or U1532 (N_1532,N_1148,N_1077);
nor U1533 (N_1533,N_1308,N_1174);
xor U1534 (N_1534,N_1468,N_1272);
and U1535 (N_1535,N_1001,N_1140);
nor U1536 (N_1536,N_1451,N_1016);
nor U1537 (N_1537,N_1119,N_1082);
xnor U1538 (N_1538,N_1394,N_1412);
xnor U1539 (N_1539,N_1246,N_1442);
or U1540 (N_1540,N_1048,N_1166);
nor U1541 (N_1541,N_1000,N_1460);
nor U1542 (N_1542,N_1291,N_1208);
nor U1543 (N_1543,N_1472,N_1385);
and U1544 (N_1544,N_1284,N_1015);
and U1545 (N_1545,N_1011,N_1477);
and U1546 (N_1546,N_1116,N_1440);
or U1547 (N_1547,N_1161,N_1127);
or U1548 (N_1548,N_1269,N_1445);
and U1549 (N_1549,N_1479,N_1178);
or U1550 (N_1550,N_1108,N_1213);
nand U1551 (N_1551,N_1135,N_1379);
nor U1552 (N_1552,N_1265,N_1075);
or U1553 (N_1553,N_1323,N_1074);
nand U1554 (N_1554,N_1035,N_1186);
or U1555 (N_1555,N_1061,N_1375);
xor U1556 (N_1556,N_1482,N_1091);
and U1557 (N_1557,N_1391,N_1098);
and U1558 (N_1558,N_1107,N_1138);
nand U1559 (N_1559,N_1117,N_1332);
nand U1560 (N_1560,N_1421,N_1111);
xor U1561 (N_1561,N_1088,N_1256);
or U1562 (N_1562,N_1368,N_1087);
xor U1563 (N_1563,N_1042,N_1465);
xnor U1564 (N_1564,N_1357,N_1260);
nor U1565 (N_1565,N_1317,N_1434);
xnor U1566 (N_1566,N_1448,N_1229);
nand U1567 (N_1567,N_1286,N_1399);
and U1568 (N_1568,N_1261,N_1149);
nor U1569 (N_1569,N_1452,N_1130);
and U1570 (N_1570,N_1418,N_1214);
or U1571 (N_1571,N_1287,N_1244);
nand U1572 (N_1572,N_1402,N_1446);
nor U1573 (N_1573,N_1069,N_1141);
nand U1574 (N_1574,N_1093,N_1463);
nor U1575 (N_1575,N_1250,N_1050);
or U1576 (N_1576,N_1466,N_1150);
nand U1577 (N_1577,N_1356,N_1145);
and U1578 (N_1578,N_1039,N_1019);
xnor U1579 (N_1579,N_1315,N_1311);
xor U1580 (N_1580,N_1471,N_1457);
or U1581 (N_1581,N_1289,N_1172);
nor U1582 (N_1582,N_1338,N_1187);
and U1583 (N_1583,N_1080,N_1247);
nor U1584 (N_1584,N_1121,N_1393);
nand U1585 (N_1585,N_1026,N_1090);
or U1586 (N_1586,N_1407,N_1012);
nand U1587 (N_1587,N_1480,N_1419);
nor U1588 (N_1588,N_1314,N_1345);
xor U1589 (N_1589,N_1106,N_1297);
xnor U1590 (N_1590,N_1328,N_1386);
xor U1591 (N_1591,N_1263,N_1240);
nor U1592 (N_1592,N_1342,N_1408);
or U1593 (N_1593,N_1305,N_1251);
nor U1594 (N_1594,N_1344,N_1177);
nor U1595 (N_1595,N_1126,N_1198);
xnor U1596 (N_1596,N_1156,N_1268);
nand U1597 (N_1597,N_1303,N_1365);
and U1598 (N_1598,N_1222,N_1013);
or U1599 (N_1599,N_1199,N_1051);
nand U1600 (N_1600,N_1420,N_1063);
xor U1601 (N_1601,N_1257,N_1207);
nor U1602 (N_1602,N_1219,N_1205);
and U1603 (N_1603,N_1059,N_1381);
xnor U1604 (N_1604,N_1239,N_1079);
nor U1605 (N_1605,N_1228,N_1153);
and U1606 (N_1606,N_1041,N_1449);
xnor U1607 (N_1607,N_1029,N_1254);
nor U1608 (N_1608,N_1046,N_1206);
nor U1609 (N_1609,N_1190,N_1462);
or U1610 (N_1610,N_1227,N_1105);
or U1611 (N_1611,N_1003,N_1025);
xor U1612 (N_1612,N_1133,N_1355);
and U1613 (N_1613,N_1363,N_1175);
or U1614 (N_1614,N_1225,N_1324);
or U1615 (N_1615,N_1298,N_1004);
or U1616 (N_1616,N_1089,N_1492);
nand U1617 (N_1617,N_1009,N_1266);
or U1618 (N_1618,N_1341,N_1109);
xor U1619 (N_1619,N_1081,N_1065);
xor U1620 (N_1620,N_1470,N_1132);
nand U1621 (N_1621,N_1264,N_1157);
or U1622 (N_1622,N_1327,N_1200);
and U1623 (N_1623,N_1497,N_1243);
xor U1624 (N_1624,N_1181,N_1070);
or U1625 (N_1625,N_1045,N_1160);
or U1626 (N_1626,N_1486,N_1095);
and U1627 (N_1627,N_1218,N_1183);
nor U1628 (N_1628,N_1437,N_1024);
or U1629 (N_1629,N_1401,N_1242);
nor U1630 (N_1630,N_1249,N_1066);
xnor U1631 (N_1631,N_1060,N_1068);
or U1632 (N_1632,N_1489,N_1278);
or U1633 (N_1633,N_1120,N_1372);
or U1634 (N_1634,N_1137,N_1101);
nand U1635 (N_1635,N_1350,N_1292);
and U1636 (N_1636,N_1493,N_1396);
nor U1637 (N_1637,N_1475,N_1474);
nand U1638 (N_1638,N_1351,N_1196);
nand U1639 (N_1639,N_1435,N_1364);
nand U1640 (N_1640,N_1403,N_1152);
xnor U1641 (N_1641,N_1425,N_1458);
or U1642 (N_1642,N_1123,N_1274);
xnor U1643 (N_1643,N_1114,N_1191);
nor U1644 (N_1644,N_1216,N_1329);
xor U1645 (N_1645,N_1320,N_1469);
nor U1646 (N_1646,N_1326,N_1043);
nor U1647 (N_1647,N_1055,N_1390);
xor U1648 (N_1648,N_1348,N_1100);
xor U1649 (N_1649,N_1333,N_1221);
and U1650 (N_1650,N_1165,N_1302);
nor U1651 (N_1651,N_1491,N_1125);
or U1652 (N_1652,N_1212,N_1014);
and U1653 (N_1653,N_1321,N_1131);
xor U1654 (N_1654,N_1112,N_1352);
xnor U1655 (N_1655,N_1032,N_1439);
nor U1656 (N_1656,N_1056,N_1283);
nand U1657 (N_1657,N_1224,N_1427);
xor U1658 (N_1658,N_1118,N_1170);
nor U1659 (N_1659,N_1300,N_1294);
and U1660 (N_1660,N_1159,N_1400);
nor U1661 (N_1661,N_1373,N_1473);
nand U1662 (N_1662,N_1167,N_1371);
nor U1663 (N_1663,N_1173,N_1414);
xor U1664 (N_1664,N_1426,N_1358);
and U1665 (N_1665,N_1217,N_1236);
nand U1666 (N_1666,N_1349,N_1232);
or U1667 (N_1667,N_1255,N_1277);
xor U1668 (N_1668,N_1279,N_1192);
nand U1669 (N_1669,N_1495,N_1144);
nand U1670 (N_1670,N_1496,N_1354);
xnor U1671 (N_1671,N_1276,N_1031);
and U1672 (N_1672,N_1142,N_1147);
nor U1673 (N_1673,N_1245,N_1275);
xnor U1674 (N_1674,N_1430,N_1388);
and U1675 (N_1675,N_1395,N_1028);
or U1676 (N_1676,N_1136,N_1424);
and U1677 (N_1677,N_1115,N_1454);
nor U1678 (N_1678,N_1189,N_1488);
xor U1679 (N_1679,N_1362,N_1444);
or U1680 (N_1680,N_1238,N_1464);
xor U1681 (N_1681,N_1335,N_1010);
nor U1682 (N_1682,N_1406,N_1182);
or U1683 (N_1683,N_1058,N_1083);
nor U1684 (N_1684,N_1164,N_1387);
nand U1685 (N_1685,N_1382,N_1282);
xor U1686 (N_1686,N_1476,N_1184);
nand U1687 (N_1687,N_1316,N_1129);
nor U1688 (N_1688,N_1377,N_1052);
or U1689 (N_1689,N_1072,N_1154);
nor U1690 (N_1690,N_1490,N_1361);
or U1691 (N_1691,N_1483,N_1215);
and U1692 (N_1692,N_1193,N_1094);
nor U1693 (N_1693,N_1441,N_1102);
nand U1694 (N_1694,N_1498,N_1485);
xor U1695 (N_1695,N_1005,N_1443);
and U1696 (N_1696,N_1271,N_1384);
and U1697 (N_1697,N_1204,N_1096);
or U1698 (N_1698,N_1134,N_1053);
nor U1699 (N_1699,N_1331,N_1461);
nand U1700 (N_1700,N_1139,N_1415);
or U1701 (N_1701,N_1030,N_1459);
xor U1702 (N_1702,N_1038,N_1027);
or U1703 (N_1703,N_1202,N_1252);
nor U1704 (N_1704,N_1423,N_1084);
and U1705 (N_1705,N_1007,N_1253);
or U1706 (N_1706,N_1413,N_1336);
xor U1707 (N_1707,N_1285,N_1467);
and U1708 (N_1708,N_1076,N_1241);
or U1709 (N_1709,N_1021,N_1325);
and U1710 (N_1710,N_1367,N_1008);
nand U1711 (N_1711,N_1220,N_1034);
and U1712 (N_1712,N_1235,N_1494);
nor U1713 (N_1713,N_1169,N_1376);
xor U1714 (N_1714,N_1313,N_1073);
and U1715 (N_1715,N_1017,N_1455);
or U1716 (N_1716,N_1299,N_1103);
nor U1717 (N_1717,N_1194,N_1023);
nand U1718 (N_1718,N_1301,N_1450);
and U1719 (N_1719,N_1185,N_1064);
xor U1720 (N_1720,N_1211,N_1310);
and U1721 (N_1721,N_1062,N_1022);
xnor U1722 (N_1722,N_1312,N_1306);
nor U1723 (N_1723,N_1456,N_1359);
xnor U1724 (N_1724,N_1307,N_1288);
nor U1725 (N_1725,N_1478,N_1340);
nor U1726 (N_1726,N_1248,N_1309);
and U1727 (N_1727,N_1411,N_1020);
or U1728 (N_1728,N_1162,N_1273);
nand U1729 (N_1729,N_1416,N_1374);
and U1730 (N_1730,N_1398,N_1209);
xnor U1731 (N_1731,N_1099,N_1188);
xnor U1732 (N_1732,N_1226,N_1432);
and U1733 (N_1733,N_1405,N_1036);
or U1734 (N_1734,N_1085,N_1168);
and U1735 (N_1735,N_1033,N_1071);
nor U1736 (N_1736,N_1179,N_1380);
and U1737 (N_1737,N_1267,N_1067);
xnor U1738 (N_1738,N_1203,N_1054);
and U1739 (N_1739,N_1334,N_1146);
or U1740 (N_1740,N_1431,N_1230);
or U1741 (N_1741,N_1447,N_1369);
or U1742 (N_1742,N_1086,N_1092);
or U1743 (N_1743,N_1259,N_1290);
nand U1744 (N_1744,N_1366,N_1128);
nor U1745 (N_1745,N_1143,N_1438);
or U1746 (N_1746,N_1258,N_1210);
nor U1747 (N_1747,N_1436,N_1319);
or U1748 (N_1748,N_1037,N_1018);
or U1749 (N_1749,N_1422,N_1318);
xnor U1750 (N_1750,N_1322,N_1241);
nor U1751 (N_1751,N_1044,N_1353);
nor U1752 (N_1752,N_1328,N_1424);
or U1753 (N_1753,N_1457,N_1199);
nor U1754 (N_1754,N_1087,N_1146);
nand U1755 (N_1755,N_1141,N_1212);
xor U1756 (N_1756,N_1392,N_1051);
and U1757 (N_1757,N_1140,N_1110);
xnor U1758 (N_1758,N_1249,N_1239);
or U1759 (N_1759,N_1108,N_1174);
or U1760 (N_1760,N_1348,N_1359);
nand U1761 (N_1761,N_1050,N_1120);
xor U1762 (N_1762,N_1268,N_1482);
nor U1763 (N_1763,N_1068,N_1393);
or U1764 (N_1764,N_1358,N_1109);
xor U1765 (N_1765,N_1133,N_1333);
xor U1766 (N_1766,N_1277,N_1200);
nand U1767 (N_1767,N_1323,N_1446);
or U1768 (N_1768,N_1201,N_1063);
nand U1769 (N_1769,N_1201,N_1277);
or U1770 (N_1770,N_1051,N_1030);
xnor U1771 (N_1771,N_1098,N_1362);
xor U1772 (N_1772,N_1394,N_1460);
and U1773 (N_1773,N_1037,N_1124);
nand U1774 (N_1774,N_1362,N_1062);
nand U1775 (N_1775,N_1218,N_1084);
and U1776 (N_1776,N_1495,N_1387);
nand U1777 (N_1777,N_1371,N_1296);
nand U1778 (N_1778,N_1160,N_1458);
or U1779 (N_1779,N_1311,N_1414);
or U1780 (N_1780,N_1087,N_1448);
nor U1781 (N_1781,N_1375,N_1276);
nor U1782 (N_1782,N_1013,N_1302);
or U1783 (N_1783,N_1304,N_1364);
xor U1784 (N_1784,N_1010,N_1092);
nor U1785 (N_1785,N_1324,N_1070);
nor U1786 (N_1786,N_1396,N_1002);
or U1787 (N_1787,N_1266,N_1244);
xnor U1788 (N_1788,N_1115,N_1190);
and U1789 (N_1789,N_1345,N_1304);
and U1790 (N_1790,N_1199,N_1368);
nand U1791 (N_1791,N_1367,N_1144);
and U1792 (N_1792,N_1066,N_1494);
nand U1793 (N_1793,N_1326,N_1327);
and U1794 (N_1794,N_1455,N_1340);
xnor U1795 (N_1795,N_1341,N_1352);
nand U1796 (N_1796,N_1288,N_1445);
xor U1797 (N_1797,N_1133,N_1347);
nor U1798 (N_1798,N_1153,N_1315);
xnor U1799 (N_1799,N_1432,N_1404);
nand U1800 (N_1800,N_1495,N_1460);
nand U1801 (N_1801,N_1126,N_1210);
nor U1802 (N_1802,N_1076,N_1126);
nand U1803 (N_1803,N_1138,N_1007);
xnor U1804 (N_1804,N_1321,N_1269);
or U1805 (N_1805,N_1292,N_1225);
and U1806 (N_1806,N_1308,N_1191);
or U1807 (N_1807,N_1303,N_1447);
and U1808 (N_1808,N_1364,N_1105);
or U1809 (N_1809,N_1208,N_1082);
or U1810 (N_1810,N_1308,N_1208);
nand U1811 (N_1811,N_1240,N_1381);
xor U1812 (N_1812,N_1152,N_1005);
or U1813 (N_1813,N_1322,N_1009);
and U1814 (N_1814,N_1184,N_1180);
xnor U1815 (N_1815,N_1289,N_1112);
nand U1816 (N_1816,N_1295,N_1486);
nor U1817 (N_1817,N_1474,N_1130);
nand U1818 (N_1818,N_1154,N_1118);
and U1819 (N_1819,N_1064,N_1180);
xor U1820 (N_1820,N_1238,N_1414);
or U1821 (N_1821,N_1392,N_1498);
nand U1822 (N_1822,N_1285,N_1203);
and U1823 (N_1823,N_1378,N_1038);
nand U1824 (N_1824,N_1157,N_1408);
xnor U1825 (N_1825,N_1398,N_1199);
and U1826 (N_1826,N_1075,N_1450);
nor U1827 (N_1827,N_1148,N_1305);
xnor U1828 (N_1828,N_1181,N_1462);
nor U1829 (N_1829,N_1194,N_1341);
nand U1830 (N_1830,N_1302,N_1485);
xor U1831 (N_1831,N_1022,N_1271);
xnor U1832 (N_1832,N_1069,N_1102);
nand U1833 (N_1833,N_1169,N_1471);
and U1834 (N_1834,N_1234,N_1399);
xor U1835 (N_1835,N_1137,N_1049);
and U1836 (N_1836,N_1407,N_1117);
xnor U1837 (N_1837,N_1051,N_1027);
xnor U1838 (N_1838,N_1368,N_1117);
xor U1839 (N_1839,N_1059,N_1246);
or U1840 (N_1840,N_1432,N_1272);
xnor U1841 (N_1841,N_1169,N_1396);
nand U1842 (N_1842,N_1436,N_1070);
xnor U1843 (N_1843,N_1201,N_1026);
nor U1844 (N_1844,N_1468,N_1360);
or U1845 (N_1845,N_1100,N_1409);
xor U1846 (N_1846,N_1169,N_1381);
nor U1847 (N_1847,N_1490,N_1212);
and U1848 (N_1848,N_1134,N_1448);
nand U1849 (N_1849,N_1309,N_1275);
or U1850 (N_1850,N_1054,N_1312);
and U1851 (N_1851,N_1483,N_1223);
nor U1852 (N_1852,N_1481,N_1266);
or U1853 (N_1853,N_1243,N_1152);
xnor U1854 (N_1854,N_1476,N_1292);
or U1855 (N_1855,N_1068,N_1380);
nor U1856 (N_1856,N_1476,N_1294);
nor U1857 (N_1857,N_1337,N_1094);
nor U1858 (N_1858,N_1330,N_1181);
nand U1859 (N_1859,N_1431,N_1030);
and U1860 (N_1860,N_1062,N_1106);
nor U1861 (N_1861,N_1425,N_1448);
or U1862 (N_1862,N_1088,N_1421);
nor U1863 (N_1863,N_1019,N_1444);
nor U1864 (N_1864,N_1014,N_1402);
xnor U1865 (N_1865,N_1208,N_1413);
xnor U1866 (N_1866,N_1067,N_1125);
nand U1867 (N_1867,N_1061,N_1224);
or U1868 (N_1868,N_1435,N_1437);
nand U1869 (N_1869,N_1143,N_1181);
or U1870 (N_1870,N_1089,N_1333);
nand U1871 (N_1871,N_1482,N_1340);
and U1872 (N_1872,N_1134,N_1172);
xor U1873 (N_1873,N_1208,N_1436);
nand U1874 (N_1874,N_1138,N_1290);
nor U1875 (N_1875,N_1251,N_1411);
nor U1876 (N_1876,N_1259,N_1236);
or U1877 (N_1877,N_1132,N_1137);
or U1878 (N_1878,N_1438,N_1157);
nand U1879 (N_1879,N_1136,N_1139);
and U1880 (N_1880,N_1014,N_1425);
xor U1881 (N_1881,N_1024,N_1000);
or U1882 (N_1882,N_1328,N_1036);
and U1883 (N_1883,N_1066,N_1214);
xor U1884 (N_1884,N_1444,N_1212);
and U1885 (N_1885,N_1092,N_1446);
nand U1886 (N_1886,N_1067,N_1362);
or U1887 (N_1887,N_1035,N_1455);
or U1888 (N_1888,N_1287,N_1185);
xnor U1889 (N_1889,N_1127,N_1461);
nor U1890 (N_1890,N_1399,N_1021);
and U1891 (N_1891,N_1297,N_1122);
and U1892 (N_1892,N_1080,N_1201);
nand U1893 (N_1893,N_1128,N_1328);
nand U1894 (N_1894,N_1031,N_1497);
nor U1895 (N_1895,N_1169,N_1421);
nand U1896 (N_1896,N_1450,N_1296);
and U1897 (N_1897,N_1067,N_1068);
nor U1898 (N_1898,N_1478,N_1319);
nand U1899 (N_1899,N_1441,N_1483);
and U1900 (N_1900,N_1073,N_1457);
and U1901 (N_1901,N_1287,N_1219);
and U1902 (N_1902,N_1065,N_1373);
and U1903 (N_1903,N_1012,N_1360);
xor U1904 (N_1904,N_1339,N_1493);
nor U1905 (N_1905,N_1061,N_1131);
xnor U1906 (N_1906,N_1149,N_1427);
or U1907 (N_1907,N_1013,N_1067);
nor U1908 (N_1908,N_1093,N_1355);
or U1909 (N_1909,N_1314,N_1482);
nor U1910 (N_1910,N_1360,N_1271);
and U1911 (N_1911,N_1149,N_1333);
nand U1912 (N_1912,N_1472,N_1157);
and U1913 (N_1913,N_1469,N_1460);
and U1914 (N_1914,N_1443,N_1180);
and U1915 (N_1915,N_1000,N_1187);
and U1916 (N_1916,N_1345,N_1211);
xor U1917 (N_1917,N_1218,N_1045);
or U1918 (N_1918,N_1392,N_1035);
nor U1919 (N_1919,N_1405,N_1136);
or U1920 (N_1920,N_1195,N_1425);
and U1921 (N_1921,N_1380,N_1424);
nor U1922 (N_1922,N_1129,N_1002);
nand U1923 (N_1923,N_1223,N_1447);
nand U1924 (N_1924,N_1419,N_1001);
or U1925 (N_1925,N_1301,N_1211);
nand U1926 (N_1926,N_1305,N_1441);
xor U1927 (N_1927,N_1353,N_1220);
xor U1928 (N_1928,N_1267,N_1406);
nor U1929 (N_1929,N_1214,N_1049);
nor U1930 (N_1930,N_1011,N_1224);
nor U1931 (N_1931,N_1297,N_1080);
nor U1932 (N_1932,N_1148,N_1245);
and U1933 (N_1933,N_1340,N_1499);
nand U1934 (N_1934,N_1485,N_1028);
xnor U1935 (N_1935,N_1391,N_1191);
and U1936 (N_1936,N_1141,N_1404);
nand U1937 (N_1937,N_1106,N_1095);
nor U1938 (N_1938,N_1039,N_1307);
and U1939 (N_1939,N_1321,N_1222);
nor U1940 (N_1940,N_1046,N_1280);
nor U1941 (N_1941,N_1396,N_1043);
nand U1942 (N_1942,N_1442,N_1274);
nand U1943 (N_1943,N_1271,N_1478);
nor U1944 (N_1944,N_1073,N_1176);
and U1945 (N_1945,N_1345,N_1199);
or U1946 (N_1946,N_1057,N_1035);
nor U1947 (N_1947,N_1103,N_1286);
nor U1948 (N_1948,N_1174,N_1054);
or U1949 (N_1949,N_1067,N_1390);
or U1950 (N_1950,N_1288,N_1048);
and U1951 (N_1951,N_1201,N_1420);
nand U1952 (N_1952,N_1489,N_1492);
or U1953 (N_1953,N_1084,N_1181);
and U1954 (N_1954,N_1474,N_1123);
nand U1955 (N_1955,N_1362,N_1395);
or U1956 (N_1956,N_1016,N_1240);
nor U1957 (N_1957,N_1328,N_1298);
and U1958 (N_1958,N_1041,N_1294);
nor U1959 (N_1959,N_1322,N_1190);
and U1960 (N_1960,N_1207,N_1093);
nor U1961 (N_1961,N_1092,N_1039);
nand U1962 (N_1962,N_1327,N_1015);
or U1963 (N_1963,N_1409,N_1451);
nand U1964 (N_1964,N_1412,N_1156);
nor U1965 (N_1965,N_1459,N_1344);
xor U1966 (N_1966,N_1076,N_1036);
nor U1967 (N_1967,N_1211,N_1462);
or U1968 (N_1968,N_1412,N_1210);
xor U1969 (N_1969,N_1206,N_1069);
xor U1970 (N_1970,N_1312,N_1010);
and U1971 (N_1971,N_1206,N_1470);
nand U1972 (N_1972,N_1332,N_1021);
or U1973 (N_1973,N_1420,N_1376);
nand U1974 (N_1974,N_1350,N_1157);
nor U1975 (N_1975,N_1412,N_1237);
and U1976 (N_1976,N_1048,N_1014);
xor U1977 (N_1977,N_1392,N_1279);
xnor U1978 (N_1978,N_1349,N_1322);
and U1979 (N_1979,N_1037,N_1202);
or U1980 (N_1980,N_1450,N_1326);
nor U1981 (N_1981,N_1232,N_1263);
nand U1982 (N_1982,N_1170,N_1377);
or U1983 (N_1983,N_1272,N_1381);
and U1984 (N_1984,N_1278,N_1355);
and U1985 (N_1985,N_1335,N_1421);
or U1986 (N_1986,N_1406,N_1487);
nand U1987 (N_1987,N_1004,N_1337);
or U1988 (N_1988,N_1458,N_1184);
nand U1989 (N_1989,N_1118,N_1414);
nor U1990 (N_1990,N_1338,N_1040);
nor U1991 (N_1991,N_1237,N_1372);
nand U1992 (N_1992,N_1217,N_1416);
and U1993 (N_1993,N_1217,N_1006);
xnor U1994 (N_1994,N_1179,N_1292);
and U1995 (N_1995,N_1248,N_1012);
xor U1996 (N_1996,N_1372,N_1309);
xnor U1997 (N_1997,N_1134,N_1226);
xor U1998 (N_1998,N_1118,N_1401);
nor U1999 (N_1999,N_1104,N_1355);
or U2000 (N_2000,N_1617,N_1738);
xor U2001 (N_2001,N_1635,N_1852);
or U2002 (N_2002,N_1554,N_1891);
or U2003 (N_2003,N_1991,N_1704);
nand U2004 (N_2004,N_1589,N_1681);
and U2005 (N_2005,N_1646,N_1702);
or U2006 (N_2006,N_1524,N_1552);
and U2007 (N_2007,N_1748,N_1625);
or U2008 (N_2008,N_1680,N_1880);
nor U2009 (N_2009,N_1531,N_1587);
xnor U2010 (N_2010,N_1515,N_1919);
or U2011 (N_2011,N_1930,N_1546);
or U2012 (N_2012,N_1613,N_1932);
nand U2013 (N_2013,N_1964,N_1507);
nor U2014 (N_2014,N_1923,N_1514);
xnor U2015 (N_2015,N_1595,N_1869);
xnor U2016 (N_2016,N_1715,N_1761);
or U2017 (N_2017,N_1872,N_1870);
or U2018 (N_2018,N_1945,N_1720);
xor U2019 (N_2019,N_1741,N_1770);
xnor U2020 (N_2020,N_1679,N_1569);
or U2021 (N_2021,N_1745,N_1944);
nand U2022 (N_2022,N_1574,N_1961);
nand U2023 (N_2023,N_1754,N_1746);
nor U2024 (N_2024,N_1585,N_1801);
or U2025 (N_2025,N_1901,N_1751);
nor U2026 (N_2026,N_1753,N_1717);
nand U2027 (N_2027,N_1830,N_1955);
nand U2028 (N_2028,N_1951,N_1672);
nor U2029 (N_2029,N_1573,N_1980);
or U2030 (N_2030,N_1785,N_1674);
or U2031 (N_2031,N_1547,N_1892);
and U2032 (N_2032,N_1757,N_1520);
nor U2033 (N_2033,N_1643,N_1926);
and U2034 (N_2034,N_1533,N_1927);
nand U2035 (N_2035,N_1975,N_1953);
or U2036 (N_2036,N_1744,N_1800);
nand U2037 (N_2037,N_1823,N_1827);
or U2038 (N_2038,N_1752,N_1576);
and U2039 (N_2039,N_1548,N_1645);
and U2040 (N_2040,N_1593,N_1619);
xor U2041 (N_2041,N_1950,N_1972);
and U2042 (N_2042,N_1984,N_1854);
and U2043 (N_2043,N_1504,N_1959);
xor U2044 (N_2044,N_1659,N_1556);
xnor U2045 (N_2045,N_1652,N_1934);
or U2046 (N_2046,N_1665,N_1618);
xnor U2047 (N_2047,N_1671,N_1612);
nand U2048 (N_2048,N_1764,N_1749);
xor U2049 (N_2049,N_1883,N_1815);
xnor U2050 (N_2050,N_1884,N_1712);
nor U2051 (N_2051,N_1867,N_1620);
or U2052 (N_2052,N_1530,N_1796);
xnor U2053 (N_2053,N_1897,N_1843);
xor U2054 (N_2054,N_1729,N_1793);
or U2055 (N_2055,N_1648,N_1722);
or U2056 (N_2056,N_1724,N_1970);
xnor U2057 (N_2057,N_1896,N_1816);
xor U2058 (N_2058,N_1505,N_1624);
nor U2059 (N_2059,N_1621,N_1839);
nor U2060 (N_2060,N_1765,N_1543);
and U2061 (N_2061,N_1693,N_1733);
nand U2062 (N_2062,N_1868,N_1769);
or U2063 (N_2063,N_1632,N_1539);
or U2064 (N_2064,N_1900,N_1644);
nor U2065 (N_2065,N_1798,N_1538);
nand U2066 (N_2066,N_1881,N_1965);
and U2067 (N_2067,N_1615,N_1791);
xnor U2068 (N_2068,N_1565,N_1985);
nand U2069 (N_2069,N_1701,N_1571);
nand U2070 (N_2070,N_1802,N_1545);
nor U2071 (N_2071,N_1768,N_1756);
xor U2072 (N_2072,N_1521,N_1570);
xor U2073 (N_2073,N_1998,N_1963);
or U2074 (N_2074,N_1694,N_1703);
and U2075 (N_2075,N_1656,N_1856);
nor U2076 (N_2076,N_1536,N_1588);
nor U2077 (N_2077,N_1742,N_1853);
or U2078 (N_2078,N_1949,N_1647);
xnor U2079 (N_2079,N_1805,N_1699);
xor U2080 (N_2080,N_1669,N_1684);
or U2081 (N_2081,N_1821,N_1808);
xor U2082 (N_2082,N_1562,N_1928);
xor U2083 (N_2083,N_1845,N_1825);
and U2084 (N_2084,N_1590,N_1713);
nand U2085 (N_2085,N_1627,N_1996);
and U2086 (N_2086,N_1743,N_1610);
nand U2087 (N_2087,N_1732,N_1654);
or U2088 (N_2088,N_1875,N_1534);
and U2089 (N_2089,N_1954,N_1682);
xor U2090 (N_2090,N_1766,N_1509);
nand U2091 (N_2091,N_1831,N_1807);
or U2092 (N_2092,N_1568,N_1982);
or U2093 (N_2093,N_1916,N_1990);
and U2094 (N_2094,N_1542,N_1526);
nor U2095 (N_2095,N_1885,N_1760);
and U2096 (N_2096,N_1506,N_1908);
nand U2097 (N_2097,N_1976,N_1832);
or U2098 (N_2098,N_1550,N_1792);
xnor U2099 (N_2099,N_1687,N_1818);
or U2100 (N_2100,N_1572,N_1979);
xnor U2101 (N_2101,N_1931,N_1859);
and U2102 (N_2102,N_1634,N_1826);
and U2103 (N_2103,N_1567,N_1555);
xnor U2104 (N_2104,N_1940,N_1840);
or U2105 (N_2105,N_1773,N_1824);
or U2106 (N_2106,N_1862,N_1532);
xnor U2107 (N_2107,N_1952,N_1636);
nor U2108 (N_2108,N_1683,N_1782);
nor U2109 (N_2109,N_1913,N_1622);
nand U2110 (N_2110,N_1605,N_1561);
nor U2111 (N_2111,N_1688,N_1566);
nand U2112 (N_2112,N_1778,N_1731);
and U2113 (N_2113,N_1811,N_1977);
nand U2114 (N_2114,N_1658,N_1623);
xor U2115 (N_2115,N_1762,N_1692);
or U2116 (N_2116,N_1657,N_1700);
nor U2117 (N_2117,N_1783,N_1600);
xor U2118 (N_2118,N_1829,N_1997);
nand U2119 (N_2119,N_1810,N_1956);
or U2120 (N_2120,N_1591,N_1988);
nand U2121 (N_2121,N_1660,N_1563);
and U2122 (N_2122,N_1895,N_1850);
or U2123 (N_2123,N_1864,N_1708);
nand U2124 (N_2124,N_1834,N_1544);
xor U2125 (N_2125,N_1887,N_1609);
or U2126 (N_2126,N_1912,N_1989);
or U2127 (N_2127,N_1848,N_1642);
and U2128 (N_2128,N_1718,N_1836);
or U2129 (N_2129,N_1966,N_1915);
nand U2130 (N_2130,N_1999,N_1835);
nand U2131 (N_2131,N_1637,N_1725);
xor U2132 (N_2132,N_1781,N_1763);
nor U2133 (N_2133,N_1938,N_1558);
or U2134 (N_2134,N_1626,N_1597);
and U2135 (N_2135,N_1819,N_1886);
and U2136 (N_2136,N_1677,N_1847);
nor U2137 (N_2137,N_1678,N_1594);
nand U2138 (N_2138,N_1935,N_1747);
or U2139 (N_2139,N_1633,N_1858);
nor U2140 (N_2140,N_1871,N_1986);
nand U2141 (N_2141,N_1511,N_1902);
nor U2142 (N_2142,N_1501,N_1795);
nand U2143 (N_2143,N_1513,N_1601);
xnor U2144 (N_2144,N_1776,N_1673);
and U2145 (N_2145,N_1994,N_1812);
and U2146 (N_2146,N_1780,N_1535);
and U2147 (N_2147,N_1933,N_1641);
or U2148 (N_2148,N_1734,N_1523);
and U2149 (N_2149,N_1592,N_1596);
xor U2150 (N_2150,N_1987,N_1579);
nand U2151 (N_2151,N_1920,N_1728);
and U2152 (N_2152,N_1664,N_1861);
nor U2153 (N_2153,N_1936,N_1755);
or U2154 (N_2154,N_1981,N_1960);
nand U2155 (N_2155,N_1500,N_1817);
nor U2156 (N_2156,N_1578,N_1974);
nand U2157 (N_2157,N_1968,N_1516);
and U2158 (N_2158,N_1517,N_1640);
nor U2159 (N_2159,N_1958,N_1921);
or U2160 (N_2160,N_1549,N_1586);
nor U2161 (N_2161,N_1750,N_1606);
or U2162 (N_2162,N_1925,N_1759);
and U2163 (N_2163,N_1696,N_1604);
nor U2164 (N_2164,N_1559,N_1739);
nor U2165 (N_2165,N_1978,N_1851);
or U2166 (N_2166,N_1584,N_1833);
and U2167 (N_2167,N_1685,N_1525);
nor U2168 (N_2168,N_1894,N_1789);
xnor U2169 (N_2169,N_1577,N_1842);
xor U2170 (N_2170,N_1638,N_1607);
or U2171 (N_2171,N_1502,N_1690);
xnor U2172 (N_2172,N_1518,N_1865);
and U2173 (N_2173,N_1799,N_1828);
nor U2174 (N_2174,N_1608,N_1860);
or U2175 (N_2175,N_1527,N_1969);
nor U2176 (N_2176,N_1857,N_1855);
nor U2177 (N_2177,N_1522,N_1602);
nand U2178 (N_2178,N_1794,N_1649);
xor U2179 (N_2179,N_1772,N_1719);
and U2180 (N_2180,N_1777,N_1670);
nor U2181 (N_2181,N_1797,N_1909);
nor U2182 (N_2182,N_1758,N_1663);
nand U2183 (N_2183,N_1710,N_1846);
or U2184 (N_2184,N_1992,N_1689);
or U2185 (N_2185,N_1714,N_1631);
nor U2186 (N_2186,N_1922,N_1804);
and U2187 (N_2187,N_1598,N_1771);
nand U2188 (N_2188,N_1866,N_1735);
xnor U2189 (N_2189,N_1786,N_1813);
nand U2190 (N_2190,N_1676,N_1614);
nor U2191 (N_2191,N_1879,N_1557);
nand U2192 (N_2192,N_1560,N_1906);
or U2193 (N_2193,N_1695,N_1726);
nor U2194 (N_2194,N_1943,N_1603);
nand U2195 (N_2195,N_1779,N_1639);
nor U2196 (N_2196,N_1904,N_1727);
nand U2197 (N_2197,N_1564,N_1971);
or U2198 (N_2198,N_1903,N_1873);
xor U2199 (N_2199,N_1551,N_1877);
or U2200 (N_2200,N_1820,N_1924);
nand U2201 (N_2201,N_1888,N_1941);
and U2202 (N_2202,N_1939,N_1993);
xnor U2203 (N_2203,N_1787,N_1705);
xnor U2204 (N_2204,N_1874,N_1918);
and U2205 (N_2205,N_1893,N_1540);
xor U2206 (N_2206,N_1882,N_1973);
xnor U2207 (N_2207,N_1774,N_1937);
nor U2208 (N_2208,N_1721,N_1711);
xor U2209 (N_2209,N_1698,N_1995);
or U2210 (N_2210,N_1723,N_1611);
nand U2211 (N_2211,N_1575,N_1898);
and U2212 (N_2212,N_1775,N_1946);
xnor U2213 (N_2213,N_1790,N_1806);
nand U2214 (N_2214,N_1662,N_1616);
nor U2215 (N_2215,N_1983,N_1653);
and U2216 (N_2216,N_1730,N_1709);
or U2217 (N_2217,N_1890,N_1863);
xnor U2218 (N_2218,N_1844,N_1841);
or U2219 (N_2219,N_1707,N_1706);
nor U2220 (N_2220,N_1675,N_1914);
xnor U2221 (N_2221,N_1528,N_1508);
or U2222 (N_2222,N_1822,N_1716);
xor U2223 (N_2223,N_1737,N_1767);
and U2224 (N_2224,N_1962,N_1668);
xnor U2225 (N_2225,N_1512,N_1876);
and U2226 (N_2226,N_1667,N_1630);
or U2227 (N_2227,N_1686,N_1553);
nand U2228 (N_2228,N_1581,N_1838);
nor U2229 (N_2229,N_1510,N_1948);
nand U2230 (N_2230,N_1583,N_1736);
and U2231 (N_2231,N_1967,N_1907);
and U2232 (N_2232,N_1929,N_1814);
nand U2233 (N_2233,N_1905,N_1837);
or U2234 (N_2234,N_1503,N_1917);
or U2235 (N_2235,N_1628,N_1942);
nor U2236 (N_2236,N_1537,N_1651);
nor U2237 (N_2237,N_1899,N_1655);
nand U2238 (N_2238,N_1529,N_1580);
and U2239 (N_2239,N_1519,N_1889);
or U2240 (N_2240,N_1666,N_1911);
nand U2241 (N_2241,N_1788,N_1878);
xnor U2242 (N_2242,N_1650,N_1803);
nand U2243 (N_2243,N_1947,N_1541);
and U2244 (N_2244,N_1691,N_1582);
xor U2245 (N_2245,N_1740,N_1599);
and U2246 (N_2246,N_1809,N_1910);
and U2247 (N_2247,N_1661,N_1784);
xor U2248 (N_2248,N_1697,N_1629);
xor U2249 (N_2249,N_1849,N_1957);
or U2250 (N_2250,N_1778,N_1881);
nand U2251 (N_2251,N_1845,N_1691);
nor U2252 (N_2252,N_1662,N_1890);
and U2253 (N_2253,N_1675,N_1894);
or U2254 (N_2254,N_1780,N_1884);
xnor U2255 (N_2255,N_1752,N_1958);
xnor U2256 (N_2256,N_1551,N_1765);
xnor U2257 (N_2257,N_1813,N_1847);
nor U2258 (N_2258,N_1569,N_1669);
nor U2259 (N_2259,N_1924,N_1607);
nand U2260 (N_2260,N_1619,N_1925);
and U2261 (N_2261,N_1859,N_1987);
nor U2262 (N_2262,N_1602,N_1660);
and U2263 (N_2263,N_1598,N_1605);
or U2264 (N_2264,N_1614,N_1536);
nor U2265 (N_2265,N_1534,N_1755);
nor U2266 (N_2266,N_1585,N_1905);
xnor U2267 (N_2267,N_1731,N_1900);
nand U2268 (N_2268,N_1902,N_1606);
nand U2269 (N_2269,N_1630,N_1970);
or U2270 (N_2270,N_1757,N_1611);
nand U2271 (N_2271,N_1709,N_1574);
and U2272 (N_2272,N_1570,N_1629);
nor U2273 (N_2273,N_1628,N_1756);
nor U2274 (N_2274,N_1602,N_1549);
nor U2275 (N_2275,N_1770,N_1644);
nor U2276 (N_2276,N_1760,N_1935);
xnor U2277 (N_2277,N_1831,N_1703);
xor U2278 (N_2278,N_1760,N_1981);
nand U2279 (N_2279,N_1508,N_1930);
xnor U2280 (N_2280,N_1712,N_1732);
or U2281 (N_2281,N_1975,N_1806);
xnor U2282 (N_2282,N_1662,N_1898);
xor U2283 (N_2283,N_1795,N_1772);
nand U2284 (N_2284,N_1690,N_1562);
and U2285 (N_2285,N_1821,N_1965);
nor U2286 (N_2286,N_1566,N_1657);
nand U2287 (N_2287,N_1811,N_1928);
nor U2288 (N_2288,N_1995,N_1632);
nor U2289 (N_2289,N_1767,N_1515);
xnor U2290 (N_2290,N_1570,N_1677);
or U2291 (N_2291,N_1791,N_1892);
nand U2292 (N_2292,N_1917,N_1910);
or U2293 (N_2293,N_1804,N_1703);
xor U2294 (N_2294,N_1980,N_1691);
xor U2295 (N_2295,N_1906,N_1876);
and U2296 (N_2296,N_1693,N_1704);
or U2297 (N_2297,N_1554,N_1566);
nor U2298 (N_2298,N_1603,N_1666);
nor U2299 (N_2299,N_1556,N_1611);
and U2300 (N_2300,N_1977,N_1758);
nand U2301 (N_2301,N_1518,N_1805);
nor U2302 (N_2302,N_1539,N_1903);
nor U2303 (N_2303,N_1691,N_1711);
and U2304 (N_2304,N_1940,N_1810);
nand U2305 (N_2305,N_1697,N_1855);
and U2306 (N_2306,N_1996,N_1925);
nand U2307 (N_2307,N_1770,N_1897);
or U2308 (N_2308,N_1879,N_1830);
nand U2309 (N_2309,N_1773,N_1650);
xnor U2310 (N_2310,N_1802,N_1816);
nand U2311 (N_2311,N_1502,N_1820);
or U2312 (N_2312,N_1956,N_1680);
nand U2313 (N_2313,N_1985,N_1754);
xnor U2314 (N_2314,N_1906,N_1923);
nand U2315 (N_2315,N_1601,N_1782);
xnor U2316 (N_2316,N_1970,N_1794);
nand U2317 (N_2317,N_1533,N_1629);
xnor U2318 (N_2318,N_1652,N_1540);
xnor U2319 (N_2319,N_1642,N_1908);
nand U2320 (N_2320,N_1667,N_1593);
nor U2321 (N_2321,N_1909,N_1734);
nand U2322 (N_2322,N_1747,N_1616);
xnor U2323 (N_2323,N_1908,N_1852);
or U2324 (N_2324,N_1698,N_1598);
xor U2325 (N_2325,N_1500,N_1820);
and U2326 (N_2326,N_1853,N_1682);
and U2327 (N_2327,N_1986,N_1876);
or U2328 (N_2328,N_1889,N_1650);
nor U2329 (N_2329,N_1762,N_1864);
nand U2330 (N_2330,N_1593,N_1645);
nor U2331 (N_2331,N_1968,N_1572);
nand U2332 (N_2332,N_1807,N_1522);
nor U2333 (N_2333,N_1667,N_1561);
or U2334 (N_2334,N_1876,N_1582);
nor U2335 (N_2335,N_1540,N_1920);
nand U2336 (N_2336,N_1947,N_1586);
and U2337 (N_2337,N_1989,N_1608);
xor U2338 (N_2338,N_1551,N_1853);
nor U2339 (N_2339,N_1576,N_1659);
or U2340 (N_2340,N_1791,N_1859);
xnor U2341 (N_2341,N_1828,N_1776);
nor U2342 (N_2342,N_1854,N_1703);
nor U2343 (N_2343,N_1778,N_1856);
nand U2344 (N_2344,N_1546,N_1818);
or U2345 (N_2345,N_1915,N_1684);
xnor U2346 (N_2346,N_1839,N_1712);
or U2347 (N_2347,N_1606,N_1726);
nand U2348 (N_2348,N_1720,N_1956);
nand U2349 (N_2349,N_1972,N_1543);
nor U2350 (N_2350,N_1984,N_1990);
nand U2351 (N_2351,N_1821,N_1857);
and U2352 (N_2352,N_1673,N_1574);
nor U2353 (N_2353,N_1611,N_1886);
or U2354 (N_2354,N_1841,N_1957);
and U2355 (N_2355,N_1529,N_1905);
or U2356 (N_2356,N_1729,N_1774);
nand U2357 (N_2357,N_1605,N_1821);
and U2358 (N_2358,N_1711,N_1651);
or U2359 (N_2359,N_1588,N_1606);
or U2360 (N_2360,N_1907,N_1550);
or U2361 (N_2361,N_1938,N_1886);
nand U2362 (N_2362,N_1534,N_1848);
nand U2363 (N_2363,N_1842,N_1916);
xor U2364 (N_2364,N_1780,N_1723);
and U2365 (N_2365,N_1852,N_1597);
nor U2366 (N_2366,N_1849,N_1752);
and U2367 (N_2367,N_1879,N_1776);
nor U2368 (N_2368,N_1620,N_1509);
nand U2369 (N_2369,N_1735,N_1628);
and U2370 (N_2370,N_1630,N_1803);
and U2371 (N_2371,N_1988,N_1847);
xnor U2372 (N_2372,N_1613,N_1570);
or U2373 (N_2373,N_1682,N_1985);
nor U2374 (N_2374,N_1752,N_1573);
and U2375 (N_2375,N_1726,N_1646);
xor U2376 (N_2376,N_1757,N_1713);
nand U2377 (N_2377,N_1503,N_1637);
nor U2378 (N_2378,N_1816,N_1948);
xor U2379 (N_2379,N_1909,N_1726);
xor U2380 (N_2380,N_1626,N_1782);
and U2381 (N_2381,N_1992,N_1952);
or U2382 (N_2382,N_1936,N_1695);
or U2383 (N_2383,N_1508,N_1824);
and U2384 (N_2384,N_1735,N_1851);
nor U2385 (N_2385,N_1845,N_1552);
or U2386 (N_2386,N_1847,N_1804);
and U2387 (N_2387,N_1744,N_1905);
or U2388 (N_2388,N_1705,N_1517);
and U2389 (N_2389,N_1641,N_1980);
xor U2390 (N_2390,N_1632,N_1838);
xor U2391 (N_2391,N_1895,N_1587);
nand U2392 (N_2392,N_1615,N_1966);
xor U2393 (N_2393,N_1852,N_1610);
nand U2394 (N_2394,N_1824,N_1502);
and U2395 (N_2395,N_1946,N_1796);
xor U2396 (N_2396,N_1881,N_1788);
xnor U2397 (N_2397,N_1662,N_1629);
or U2398 (N_2398,N_1899,N_1929);
and U2399 (N_2399,N_1539,N_1898);
and U2400 (N_2400,N_1772,N_1928);
and U2401 (N_2401,N_1942,N_1677);
xnor U2402 (N_2402,N_1568,N_1895);
xor U2403 (N_2403,N_1881,N_1971);
or U2404 (N_2404,N_1902,N_1517);
or U2405 (N_2405,N_1926,N_1517);
or U2406 (N_2406,N_1620,N_1834);
xor U2407 (N_2407,N_1969,N_1521);
nand U2408 (N_2408,N_1599,N_1869);
and U2409 (N_2409,N_1995,N_1908);
and U2410 (N_2410,N_1534,N_1760);
xnor U2411 (N_2411,N_1541,N_1827);
or U2412 (N_2412,N_1662,N_1604);
and U2413 (N_2413,N_1567,N_1694);
xor U2414 (N_2414,N_1963,N_1767);
or U2415 (N_2415,N_1784,N_1734);
nand U2416 (N_2416,N_1628,N_1955);
and U2417 (N_2417,N_1941,N_1929);
xnor U2418 (N_2418,N_1644,N_1713);
nor U2419 (N_2419,N_1962,N_1834);
nand U2420 (N_2420,N_1576,N_1833);
xor U2421 (N_2421,N_1943,N_1806);
or U2422 (N_2422,N_1743,N_1899);
nand U2423 (N_2423,N_1588,N_1884);
nand U2424 (N_2424,N_1567,N_1737);
or U2425 (N_2425,N_1637,N_1678);
xnor U2426 (N_2426,N_1794,N_1925);
nand U2427 (N_2427,N_1966,N_1601);
or U2428 (N_2428,N_1984,N_1590);
and U2429 (N_2429,N_1885,N_1706);
and U2430 (N_2430,N_1579,N_1614);
nor U2431 (N_2431,N_1845,N_1756);
or U2432 (N_2432,N_1862,N_1963);
nand U2433 (N_2433,N_1566,N_1905);
or U2434 (N_2434,N_1548,N_1792);
xnor U2435 (N_2435,N_1719,N_1649);
nor U2436 (N_2436,N_1807,N_1886);
nor U2437 (N_2437,N_1876,N_1620);
nor U2438 (N_2438,N_1661,N_1619);
or U2439 (N_2439,N_1574,N_1664);
xnor U2440 (N_2440,N_1943,N_1503);
and U2441 (N_2441,N_1534,N_1780);
or U2442 (N_2442,N_1514,N_1830);
nand U2443 (N_2443,N_1738,N_1970);
and U2444 (N_2444,N_1863,N_1884);
and U2445 (N_2445,N_1671,N_1819);
or U2446 (N_2446,N_1916,N_1806);
nand U2447 (N_2447,N_1711,N_1945);
and U2448 (N_2448,N_1735,N_1725);
or U2449 (N_2449,N_1604,N_1740);
nand U2450 (N_2450,N_1699,N_1755);
nand U2451 (N_2451,N_1628,N_1567);
and U2452 (N_2452,N_1610,N_1964);
xor U2453 (N_2453,N_1627,N_1603);
and U2454 (N_2454,N_1866,N_1573);
nand U2455 (N_2455,N_1862,N_1816);
xnor U2456 (N_2456,N_1525,N_1818);
nor U2457 (N_2457,N_1575,N_1733);
and U2458 (N_2458,N_1853,N_1816);
xor U2459 (N_2459,N_1567,N_1580);
or U2460 (N_2460,N_1508,N_1891);
or U2461 (N_2461,N_1791,N_1607);
nand U2462 (N_2462,N_1992,N_1573);
or U2463 (N_2463,N_1687,N_1637);
nor U2464 (N_2464,N_1876,N_1579);
and U2465 (N_2465,N_1865,N_1771);
and U2466 (N_2466,N_1848,N_1517);
xnor U2467 (N_2467,N_1796,N_1751);
and U2468 (N_2468,N_1874,N_1964);
or U2469 (N_2469,N_1672,N_1965);
or U2470 (N_2470,N_1754,N_1704);
nor U2471 (N_2471,N_1991,N_1598);
xnor U2472 (N_2472,N_1500,N_1779);
nor U2473 (N_2473,N_1528,N_1620);
and U2474 (N_2474,N_1753,N_1676);
and U2475 (N_2475,N_1690,N_1967);
xnor U2476 (N_2476,N_1728,N_1629);
or U2477 (N_2477,N_1956,N_1962);
or U2478 (N_2478,N_1620,N_1860);
nand U2479 (N_2479,N_1861,N_1629);
and U2480 (N_2480,N_1737,N_1743);
xor U2481 (N_2481,N_1644,N_1593);
xnor U2482 (N_2482,N_1745,N_1542);
nand U2483 (N_2483,N_1839,N_1634);
or U2484 (N_2484,N_1963,N_1996);
nand U2485 (N_2485,N_1512,N_1543);
nor U2486 (N_2486,N_1763,N_1874);
nand U2487 (N_2487,N_1843,N_1541);
nand U2488 (N_2488,N_1586,N_1640);
nand U2489 (N_2489,N_1854,N_1929);
nor U2490 (N_2490,N_1555,N_1702);
or U2491 (N_2491,N_1748,N_1734);
nor U2492 (N_2492,N_1502,N_1756);
xor U2493 (N_2493,N_1712,N_1619);
xor U2494 (N_2494,N_1552,N_1873);
xor U2495 (N_2495,N_1760,N_1622);
and U2496 (N_2496,N_1736,N_1988);
or U2497 (N_2497,N_1801,N_1760);
xor U2498 (N_2498,N_1579,N_1706);
xor U2499 (N_2499,N_1919,N_1725);
xor U2500 (N_2500,N_2230,N_2021);
and U2501 (N_2501,N_2302,N_2389);
nor U2502 (N_2502,N_2191,N_2170);
xor U2503 (N_2503,N_2109,N_2199);
nand U2504 (N_2504,N_2373,N_2332);
xor U2505 (N_2505,N_2227,N_2487);
and U2506 (N_2506,N_2308,N_2384);
nand U2507 (N_2507,N_2448,N_2045);
nand U2508 (N_2508,N_2040,N_2043);
nand U2509 (N_2509,N_2229,N_2125);
or U2510 (N_2510,N_2347,N_2435);
xor U2511 (N_2511,N_2479,N_2374);
xnor U2512 (N_2512,N_2190,N_2341);
and U2513 (N_2513,N_2258,N_2097);
xnor U2514 (N_2514,N_2102,N_2242);
xnor U2515 (N_2515,N_2322,N_2355);
xor U2516 (N_2516,N_2444,N_2124);
nor U2517 (N_2517,N_2052,N_2391);
nand U2518 (N_2518,N_2395,N_2012);
and U2519 (N_2519,N_2293,N_2168);
nor U2520 (N_2520,N_2113,N_2066);
nand U2521 (N_2521,N_2343,N_2305);
and U2522 (N_2522,N_2336,N_2408);
nand U2523 (N_2523,N_2120,N_2018);
xor U2524 (N_2524,N_2006,N_2110);
and U2525 (N_2525,N_2091,N_2087);
xnor U2526 (N_2526,N_2453,N_2264);
or U2527 (N_2527,N_2153,N_2425);
nand U2528 (N_2528,N_2237,N_2112);
nor U2529 (N_2529,N_2461,N_2300);
and U2530 (N_2530,N_2495,N_2096);
nor U2531 (N_2531,N_2318,N_2064);
and U2532 (N_2532,N_2286,N_2457);
or U2533 (N_2533,N_2416,N_2010);
or U2534 (N_2534,N_2131,N_2345);
and U2535 (N_2535,N_2001,N_2253);
xnor U2536 (N_2536,N_2086,N_2438);
nor U2537 (N_2537,N_2314,N_2164);
nor U2538 (N_2538,N_2002,N_2289);
nor U2539 (N_2539,N_2447,N_2205);
xor U2540 (N_2540,N_2081,N_2259);
xnor U2541 (N_2541,N_2411,N_2019);
and U2542 (N_2542,N_2261,N_2419);
or U2543 (N_2543,N_2246,N_2366);
xor U2544 (N_2544,N_2026,N_2069);
nand U2545 (N_2545,N_2030,N_2173);
xnor U2546 (N_2546,N_2197,N_2148);
nand U2547 (N_2547,N_2473,N_2492);
or U2548 (N_2548,N_2111,N_2491);
xnor U2549 (N_2549,N_2126,N_2134);
nand U2550 (N_2550,N_2020,N_2195);
nand U2551 (N_2551,N_2218,N_2100);
nor U2552 (N_2552,N_2428,N_2455);
nor U2553 (N_2553,N_2059,N_2372);
and U2554 (N_2554,N_2454,N_2079);
xor U2555 (N_2555,N_2145,N_2339);
or U2556 (N_2556,N_2203,N_2039);
and U2557 (N_2557,N_2114,N_2049);
nand U2558 (N_2558,N_2418,N_2443);
or U2559 (N_2559,N_2046,N_2015);
and U2560 (N_2560,N_2146,N_2144);
nor U2561 (N_2561,N_2274,N_2279);
and U2562 (N_2562,N_2141,N_2223);
xor U2563 (N_2563,N_2304,N_2121);
nand U2564 (N_2564,N_2239,N_2252);
and U2565 (N_2565,N_2474,N_2149);
xnor U2566 (N_2566,N_2159,N_2247);
nor U2567 (N_2567,N_2422,N_2234);
xnor U2568 (N_2568,N_2061,N_2367);
or U2569 (N_2569,N_2370,N_2358);
or U2570 (N_2570,N_2349,N_2353);
nand U2571 (N_2571,N_2053,N_2270);
nor U2572 (N_2572,N_2430,N_2310);
xor U2573 (N_2573,N_2468,N_2179);
nand U2574 (N_2574,N_2129,N_2160);
nand U2575 (N_2575,N_2417,N_2137);
and U2576 (N_2576,N_2445,N_2003);
nor U2577 (N_2577,N_2449,N_2285);
nor U2578 (N_2578,N_2094,N_2232);
nand U2579 (N_2579,N_2278,N_2499);
xor U2580 (N_2580,N_2276,N_2426);
xnor U2581 (N_2581,N_2017,N_2470);
and U2582 (N_2582,N_2210,N_2014);
xnor U2583 (N_2583,N_2241,N_2383);
nor U2584 (N_2584,N_2004,N_2140);
and U2585 (N_2585,N_2334,N_2090);
and U2586 (N_2586,N_2397,N_2496);
xnor U2587 (N_2587,N_2362,N_2065);
nor U2588 (N_2588,N_2167,N_2044);
xor U2589 (N_2589,N_2078,N_2007);
nand U2590 (N_2590,N_2188,N_2378);
or U2591 (N_2591,N_2238,N_2316);
nand U2592 (N_2592,N_2363,N_2421);
or U2593 (N_2593,N_2452,N_2333);
nand U2594 (N_2594,N_2055,N_2284);
or U2595 (N_2595,N_2122,N_2398);
nand U2596 (N_2596,N_2151,N_2072);
or U2597 (N_2597,N_2023,N_2268);
nor U2598 (N_2598,N_2233,N_2106);
or U2599 (N_2599,N_2209,N_2458);
nand U2600 (N_2600,N_2317,N_2387);
and U2601 (N_2601,N_2471,N_2104);
or U2602 (N_2602,N_2360,N_2000);
xnor U2603 (N_2603,N_2409,N_2335);
and U2604 (N_2604,N_2181,N_2208);
or U2605 (N_2605,N_2375,N_2291);
and U2606 (N_2606,N_2295,N_2415);
xnor U2607 (N_2607,N_2163,N_2287);
and U2608 (N_2608,N_2108,N_2074);
and U2609 (N_2609,N_2182,N_2076);
or U2610 (N_2610,N_2156,N_2013);
nor U2611 (N_2611,N_2342,N_2150);
nand U2612 (N_2612,N_2005,N_2154);
and U2613 (N_2613,N_2257,N_2290);
nand U2614 (N_2614,N_2269,N_2123);
nor U2615 (N_2615,N_2202,N_2338);
or U2616 (N_2616,N_2364,N_2119);
xnor U2617 (N_2617,N_2138,N_2369);
xor U2618 (N_2618,N_2174,N_2051);
xnor U2619 (N_2619,N_2215,N_2396);
or U2620 (N_2620,N_2117,N_2207);
xor U2621 (N_2621,N_2427,N_2147);
or U2622 (N_2622,N_2399,N_2486);
and U2623 (N_2623,N_2143,N_2288);
and U2624 (N_2624,N_2319,N_2033);
and U2625 (N_2625,N_2410,N_2429);
or U2626 (N_2626,N_2184,N_2282);
nor U2627 (N_2627,N_2099,N_2325);
or U2628 (N_2628,N_2206,N_2324);
xnor U2629 (N_2629,N_2371,N_2381);
and U2630 (N_2630,N_2472,N_2498);
or U2631 (N_2631,N_2357,N_2477);
or U2632 (N_2632,N_2404,N_2235);
or U2633 (N_2633,N_2344,N_2062);
nand U2634 (N_2634,N_2077,N_2193);
and U2635 (N_2635,N_2058,N_2073);
or U2636 (N_2636,N_2323,N_2437);
nor U2637 (N_2637,N_2130,N_2490);
nand U2638 (N_2638,N_2228,N_2216);
nand U2639 (N_2639,N_2480,N_2315);
nand U2640 (N_2640,N_2194,N_2393);
nand U2641 (N_2641,N_2189,N_2068);
and U2642 (N_2642,N_2440,N_2166);
and U2643 (N_2643,N_2254,N_2424);
nand U2644 (N_2644,N_2475,N_2298);
nand U2645 (N_2645,N_2158,N_2027);
nor U2646 (N_2646,N_2272,N_2379);
xnor U2647 (N_2647,N_2326,N_2225);
or U2648 (N_2648,N_2089,N_2420);
nand U2649 (N_2649,N_2183,N_2083);
xnor U2650 (N_2650,N_2459,N_2331);
nand U2651 (N_2651,N_2054,N_2266);
xor U2652 (N_2652,N_2361,N_2465);
nor U2653 (N_2653,N_2376,N_2400);
xnor U2654 (N_2654,N_2031,N_2301);
and U2655 (N_2655,N_2201,N_2297);
and U2656 (N_2656,N_2139,N_2497);
nand U2657 (N_2657,N_2439,N_2101);
xor U2658 (N_2658,N_2296,N_2115);
nor U2659 (N_2659,N_2463,N_2098);
xnor U2660 (N_2660,N_2243,N_2390);
and U2661 (N_2661,N_2456,N_2180);
or U2662 (N_2662,N_2277,N_2165);
nand U2663 (N_2663,N_2133,N_2385);
or U2664 (N_2664,N_2403,N_2142);
and U2665 (N_2665,N_2063,N_2405);
and U2666 (N_2666,N_2161,N_2103);
xnor U2667 (N_2667,N_2280,N_2292);
xor U2668 (N_2668,N_2032,N_2309);
or U2669 (N_2669,N_2155,N_2231);
or U2670 (N_2670,N_2485,N_2388);
and U2671 (N_2671,N_2359,N_2483);
xnor U2672 (N_2672,N_2434,N_2263);
or U2673 (N_2673,N_2025,N_2116);
nor U2674 (N_2674,N_2407,N_2135);
nor U2675 (N_2675,N_2350,N_2368);
and U2676 (N_2676,N_2313,N_2037);
nand U2677 (N_2677,N_2084,N_2041);
or U2678 (N_2678,N_2082,N_2431);
xnor U2679 (N_2679,N_2198,N_2303);
or U2680 (N_2680,N_2494,N_2450);
xor U2681 (N_2681,N_2071,N_2050);
nand U2682 (N_2682,N_2219,N_2035);
xor U2683 (N_2683,N_2320,N_2009);
or U2684 (N_2684,N_2478,N_2481);
or U2685 (N_2685,N_2392,N_2176);
nand U2686 (N_2686,N_2105,N_2451);
or U2687 (N_2687,N_2067,N_2414);
or U2688 (N_2688,N_2187,N_2070);
and U2689 (N_2689,N_2432,N_2047);
and U2690 (N_2690,N_2249,N_2482);
or U2691 (N_2691,N_2011,N_2008);
nand U2692 (N_2692,N_2406,N_2401);
xor U2693 (N_2693,N_2251,N_2356);
nand U2694 (N_2694,N_2446,N_2256);
and U2695 (N_2695,N_2213,N_2107);
xnor U2696 (N_2696,N_2024,N_2060);
nand U2697 (N_2697,N_2281,N_2330);
nor U2698 (N_2698,N_2036,N_2132);
nor U2699 (N_2699,N_2224,N_2307);
xor U2700 (N_2700,N_2245,N_2192);
nand U2701 (N_2701,N_2283,N_2136);
xor U2702 (N_2702,N_2214,N_2057);
nor U2703 (N_2703,N_2016,N_2321);
xor U2704 (N_2704,N_2244,N_2412);
or U2705 (N_2705,N_2413,N_2042);
xor U2706 (N_2706,N_2311,N_2460);
and U2707 (N_2707,N_2299,N_2466);
or U2708 (N_2708,N_2354,N_2394);
or U2709 (N_2709,N_2493,N_2436);
nor U2710 (N_2710,N_2088,N_2221);
or U2711 (N_2711,N_2157,N_2172);
and U2712 (N_2712,N_2380,N_2352);
or U2713 (N_2713,N_2464,N_2034);
nor U2714 (N_2714,N_2346,N_2095);
xor U2715 (N_2715,N_2211,N_2178);
and U2716 (N_2716,N_2348,N_2265);
or U2717 (N_2717,N_2423,N_2469);
nand U2718 (N_2718,N_2260,N_2382);
nand U2719 (N_2719,N_2248,N_2175);
and U2720 (N_2720,N_2441,N_2275);
nand U2721 (N_2721,N_2328,N_2177);
or U2722 (N_2722,N_2196,N_2271);
and U2723 (N_2723,N_2029,N_2075);
and U2724 (N_2724,N_2226,N_2294);
nor U2725 (N_2725,N_2340,N_2171);
and U2726 (N_2726,N_2489,N_2212);
nand U2727 (N_2727,N_2092,N_2222);
and U2728 (N_2728,N_2377,N_2169);
nand U2729 (N_2729,N_2250,N_2093);
or U2730 (N_2730,N_2267,N_2118);
or U2731 (N_2731,N_2152,N_2262);
nand U2732 (N_2732,N_2022,N_2337);
xor U2733 (N_2733,N_2128,N_2240);
or U2734 (N_2734,N_2402,N_2186);
nor U2735 (N_2735,N_2306,N_2204);
and U2736 (N_2736,N_2329,N_2028);
nor U2737 (N_2737,N_2162,N_2386);
and U2738 (N_2738,N_2236,N_2351);
or U2739 (N_2739,N_2365,N_2255);
nor U2740 (N_2740,N_2467,N_2048);
nor U2741 (N_2741,N_2327,N_2217);
xor U2742 (N_2742,N_2085,N_2273);
nand U2743 (N_2743,N_2127,N_2442);
nand U2744 (N_2744,N_2056,N_2200);
nand U2745 (N_2745,N_2488,N_2312);
nand U2746 (N_2746,N_2080,N_2038);
nor U2747 (N_2747,N_2220,N_2476);
or U2748 (N_2748,N_2185,N_2484);
nor U2749 (N_2749,N_2433,N_2462);
nor U2750 (N_2750,N_2443,N_2060);
or U2751 (N_2751,N_2361,N_2400);
xnor U2752 (N_2752,N_2204,N_2272);
and U2753 (N_2753,N_2355,N_2039);
xnor U2754 (N_2754,N_2106,N_2144);
xnor U2755 (N_2755,N_2194,N_2398);
nand U2756 (N_2756,N_2207,N_2267);
and U2757 (N_2757,N_2403,N_2112);
xnor U2758 (N_2758,N_2469,N_2127);
and U2759 (N_2759,N_2207,N_2086);
or U2760 (N_2760,N_2054,N_2081);
xor U2761 (N_2761,N_2122,N_2498);
and U2762 (N_2762,N_2135,N_2074);
and U2763 (N_2763,N_2305,N_2222);
nor U2764 (N_2764,N_2134,N_2028);
and U2765 (N_2765,N_2359,N_2158);
nand U2766 (N_2766,N_2478,N_2371);
nor U2767 (N_2767,N_2019,N_2001);
nand U2768 (N_2768,N_2354,N_2121);
and U2769 (N_2769,N_2191,N_2278);
nand U2770 (N_2770,N_2224,N_2302);
or U2771 (N_2771,N_2296,N_2352);
and U2772 (N_2772,N_2266,N_2229);
or U2773 (N_2773,N_2220,N_2482);
xor U2774 (N_2774,N_2456,N_2206);
and U2775 (N_2775,N_2274,N_2427);
and U2776 (N_2776,N_2386,N_2328);
or U2777 (N_2777,N_2274,N_2311);
nor U2778 (N_2778,N_2016,N_2088);
or U2779 (N_2779,N_2003,N_2379);
nor U2780 (N_2780,N_2221,N_2070);
or U2781 (N_2781,N_2345,N_2399);
or U2782 (N_2782,N_2271,N_2252);
and U2783 (N_2783,N_2438,N_2290);
nor U2784 (N_2784,N_2358,N_2463);
xnor U2785 (N_2785,N_2052,N_2024);
or U2786 (N_2786,N_2261,N_2282);
and U2787 (N_2787,N_2221,N_2214);
or U2788 (N_2788,N_2338,N_2074);
xnor U2789 (N_2789,N_2021,N_2342);
xnor U2790 (N_2790,N_2047,N_2159);
xnor U2791 (N_2791,N_2014,N_2415);
or U2792 (N_2792,N_2352,N_2035);
nor U2793 (N_2793,N_2316,N_2021);
nand U2794 (N_2794,N_2381,N_2486);
xor U2795 (N_2795,N_2154,N_2050);
nor U2796 (N_2796,N_2013,N_2140);
xnor U2797 (N_2797,N_2385,N_2458);
xnor U2798 (N_2798,N_2142,N_2326);
xor U2799 (N_2799,N_2174,N_2181);
xor U2800 (N_2800,N_2349,N_2285);
xnor U2801 (N_2801,N_2249,N_2102);
nor U2802 (N_2802,N_2448,N_2103);
nand U2803 (N_2803,N_2055,N_2408);
nand U2804 (N_2804,N_2232,N_2003);
and U2805 (N_2805,N_2011,N_2001);
nand U2806 (N_2806,N_2316,N_2205);
xor U2807 (N_2807,N_2266,N_2295);
xnor U2808 (N_2808,N_2446,N_2476);
xor U2809 (N_2809,N_2129,N_2228);
nand U2810 (N_2810,N_2129,N_2072);
or U2811 (N_2811,N_2442,N_2280);
and U2812 (N_2812,N_2027,N_2162);
or U2813 (N_2813,N_2104,N_2162);
xnor U2814 (N_2814,N_2146,N_2433);
nor U2815 (N_2815,N_2471,N_2089);
nor U2816 (N_2816,N_2465,N_2144);
or U2817 (N_2817,N_2162,N_2099);
and U2818 (N_2818,N_2071,N_2341);
nor U2819 (N_2819,N_2076,N_2301);
xor U2820 (N_2820,N_2386,N_2482);
nand U2821 (N_2821,N_2380,N_2023);
xor U2822 (N_2822,N_2217,N_2181);
or U2823 (N_2823,N_2179,N_2101);
nor U2824 (N_2824,N_2473,N_2278);
or U2825 (N_2825,N_2203,N_2210);
or U2826 (N_2826,N_2470,N_2070);
nor U2827 (N_2827,N_2127,N_2245);
xor U2828 (N_2828,N_2340,N_2407);
or U2829 (N_2829,N_2378,N_2386);
or U2830 (N_2830,N_2014,N_2125);
xor U2831 (N_2831,N_2017,N_2032);
or U2832 (N_2832,N_2329,N_2475);
nor U2833 (N_2833,N_2214,N_2093);
nor U2834 (N_2834,N_2227,N_2065);
or U2835 (N_2835,N_2006,N_2305);
or U2836 (N_2836,N_2138,N_2056);
nand U2837 (N_2837,N_2253,N_2015);
xnor U2838 (N_2838,N_2030,N_2064);
xnor U2839 (N_2839,N_2060,N_2201);
nor U2840 (N_2840,N_2096,N_2083);
nand U2841 (N_2841,N_2407,N_2466);
or U2842 (N_2842,N_2103,N_2166);
or U2843 (N_2843,N_2061,N_2352);
and U2844 (N_2844,N_2417,N_2313);
or U2845 (N_2845,N_2223,N_2383);
nand U2846 (N_2846,N_2444,N_2237);
or U2847 (N_2847,N_2231,N_2050);
and U2848 (N_2848,N_2232,N_2474);
nor U2849 (N_2849,N_2049,N_2020);
nand U2850 (N_2850,N_2224,N_2278);
and U2851 (N_2851,N_2249,N_2337);
nor U2852 (N_2852,N_2293,N_2167);
and U2853 (N_2853,N_2414,N_2192);
and U2854 (N_2854,N_2480,N_2182);
xor U2855 (N_2855,N_2003,N_2211);
nor U2856 (N_2856,N_2221,N_2395);
nor U2857 (N_2857,N_2445,N_2430);
nand U2858 (N_2858,N_2411,N_2383);
nand U2859 (N_2859,N_2244,N_2347);
or U2860 (N_2860,N_2003,N_2086);
nand U2861 (N_2861,N_2356,N_2249);
xnor U2862 (N_2862,N_2286,N_2315);
nand U2863 (N_2863,N_2170,N_2133);
and U2864 (N_2864,N_2079,N_2480);
or U2865 (N_2865,N_2068,N_2148);
nand U2866 (N_2866,N_2345,N_2227);
and U2867 (N_2867,N_2215,N_2426);
xnor U2868 (N_2868,N_2444,N_2328);
and U2869 (N_2869,N_2453,N_2390);
xor U2870 (N_2870,N_2231,N_2307);
and U2871 (N_2871,N_2249,N_2411);
and U2872 (N_2872,N_2336,N_2389);
and U2873 (N_2873,N_2030,N_2239);
nand U2874 (N_2874,N_2314,N_2027);
nand U2875 (N_2875,N_2478,N_2216);
nand U2876 (N_2876,N_2022,N_2417);
or U2877 (N_2877,N_2471,N_2466);
nand U2878 (N_2878,N_2235,N_2005);
xor U2879 (N_2879,N_2396,N_2059);
xnor U2880 (N_2880,N_2021,N_2129);
nor U2881 (N_2881,N_2036,N_2406);
nor U2882 (N_2882,N_2043,N_2346);
and U2883 (N_2883,N_2265,N_2241);
nand U2884 (N_2884,N_2012,N_2498);
and U2885 (N_2885,N_2410,N_2269);
xor U2886 (N_2886,N_2469,N_2042);
or U2887 (N_2887,N_2274,N_2314);
nand U2888 (N_2888,N_2081,N_2431);
nand U2889 (N_2889,N_2219,N_2048);
and U2890 (N_2890,N_2126,N_2453);
nand U2891 (N_2891,N_2093,N_2225);
and U2892 (N_2892,N_2044,N_2090);
nand U2893 (N_2893,N_2033,N_2451);
xor U2894 (N_2894,N_2377,N_2099);
xnor U2895 (N_2895,N_2061,N_2123);
nand U2896 (N_2896,N_2235,N_2492);
or U2897 (N_2897,N_2245,N_2043);
nor U2898 (N_2898,N_2272,N_2290);
nor U2899 (N_2899,N_2469,N_2068);
xnor U2900 (N_2900,N_2078,N_2214);
and U2901 (N_2901,N_2049,N_2229);
and U2902 (N_2902,N_2091,N_2327);
or U2903 (N_2903,N_2332,N_2468);
nor U2904 (N_2904,N_2435,N_2100);
xnor U2905 (N_2905,N_2092,N_2209);
or U2906 (N_2906,N_2493,N_2207);
or U2907 (N_2907,N_2346,N_2008);
and U2908 (N_2908,N_2018,N_2374);
or U2909 (N_2909,N_2331,N_2477);
and U2910 (N_2910,N_2145,N_2207);
xnor U2911 (N_2911,N_2157,N_2303);
nor U2912 (N_2912,N_2318,N_2488);
nor U2913 (N_2913,N_2022,N_2067);
or U2914 (N_2914,N_2208,N_2107);
nand U2915 (N_2915,N_2357,N_2429);
nand U2916 (N_2916,N_2448,N_2398);
nand U2917 (N_2917,N_2026,N_2335);
xnor U2918 (N_2918,N_2291,N_2002);
and U2919 (N_2919,N_2352,N_2408);
or U2920 (N_2920,N_2392,N_2184);
xnor U2921 (N_2921,N_2028,N_2491);
xor U2922 (N_2922,N_2211,N_2329);
or U2923 (N_2923,N_2017,N_2264);
xnor U2924 (N_2924,N_2419,N_2331);
nor U2925 (N_2925,N_2094,N_2496);
nor U2926 (N_2926,N_2324,N_2008);
and U2927 (N_2927,N_2016,N_2060);
xnor U2928 (N_2928,N_2042,N_2075);
nor U2929 (N_2929,N_2388,N_2288);
or U2930 (N_2930,N_2143,N_2097);
xnor U2931 (N_2931,N_2457,N_2052);
xnor U2932 (N_2932,N_2219,N_2405);
xnor U2933 (N_2933,N_2480,N_2170);
nor U2934 (N_2934,N_2332,N_2355);
or U2935 (N_2935,N_2427,N_2292);
or U2936 (N_2936,N_2310,N_2238);
and U2937 (N_2937,N_2091,N_2383);
xor U2938 (N_2938,N_2141,N_2142);
xnor U2939 (N_2939,N_2020,N_2487);
or U2940 (N_2940,N_2438,N_2403);
or U2941 (N_2941,N_2000,N_2458);
nor U2942 (N_2942,N_2062,N_2102);
xor U2943 (N_2943,N_2283,N_2166);
xnor U2944 (N_2944,N_2385,N_2041);
nor U2945 (N_2945,N_2468,N_2256);
and U2946 (N_2946,N_2181,N_2037);
nor U2947 (N_2947,N_2139,N_2006);
nand U2948 (N_2948,N_2020,N_2120);
xor U2949 (N_2949,N_2369,N_2208);
and U2950 (N_2950,N_2198,N_2318);
or U2951 (N_2951,N_2141,N_2320);
xnor U2952 (N_2952,N_2326,N_2375);
or U2953 (N_2953,N_2316,N_2498);
and U2954 (N_2954,N_2010,N_2400);
nor U2955 (N_2955,N_2118,N_2027);
and U2956 (N_2956,N_2192,N_2416);
and U2957 (N_2957,N_2168,N_2477);
or U2958 (N_2958,N_2298,N_2183);
and U2959 (N_2959,N_2266,N_2269);
nand U2960 (N_2960,N_2178,N_2470);
xnor U2961 (N_2961,N_2241,N_2314);
and U2962 (N_2962,N_2130,N_2212);
xor U2963 (N_2963,N_2178,N_2142);
xnor U2964 (N_2964,N_2199,N_2076);
xnor U2965 (N_2965,N_2457,N_2395);
xor U2966 (N_2966,N_2442,N_2205);
nor U2967 (N_2967,N_2208,N_2321);
nor U2968 (N_2968,N_2307,N_2148);
nor U2969 (N_2969,N_2180,N_2108);
nor U2970 (N_2970,N_2386,N_2408);
or U2971 (N_2971,N_2059,N_2226);
or U2972 (N_2972,N_2442,N_2023);
nand U2973 (N_2973,N_2034,N_2373);
and U2974 (N_2974,N_2391,N_2271);
or U2975 (N_2975,N_2204,N_2077);
xor U2976 (N_2976,N_2356,N_2054);
nand U2977 (N_2977,N_2324,N_2301);
nand U2978 (N_2978,N_2261,N_2414);
and U2979 (N_2979,N_2171,N_2317);
or U2980 (N_2980,N_2235,N_2135);
nor U2981 (N_2981,N_2058,N_2311);
and U2982 (N_2982,N_2327,N_2015);
xnor U2983 (N_2983,N_2472,N_2168);
nand U2984 (N_2984,N_2282,N_2004);
xnor U2985 (N_2985,N_2295,N_2015);
nand U2986 (N_2986,N_2452,N_2250);
nor U2987 (N_2987,N_2356,N_2196);
and U2988 (N_2988,N_2249,N_2495);
xor U2989 (N_2989,N_2415,N_2327);
nor U2990 (N_2990,N_2499,N_2406);
xnor U2991 (N_2991,N_2100,N_2114);
nor U2992 (N_2992,N_2339,N_2361);
and U2993 (N_2993,N_2096,N_2059);
xor U2994 (N_2994,N_2144,N_2209);
nor U2995 (N_2995,N_2226,N_2328);
nand U2996 (N_2996,N_2262,N_2076);
nor U2997 (N_2997,N_2386,N_2136);
or U2998 (N_2998,N_2062,N_2480);
or U2999 (N_2999,N_2214,N_2395);
nor U3000 (N_3000,N_2944,N_2586);
or U3001 (N_3001,N_2688,N_2817);
nor U3002 (N_3002,N_2909,N_2749);
or U3003 (N_3003,N_2813,N_2916);
xnor U3004 (N_3004,N_2747,N_2739);
and U3005 (N_3005,N_2553,N_2700);
xor U3006 (N_3006,N_2927,N_2743);
xnor U3007 (N_3007,N_2849,N_2830);
nand U3008 (N_3008,N_2685,N_2973);
nand U3009 (N_3009,N_2615,N_2926);
and U3010 (N_3010,N_2925,N_2882);
nand U3011 (N_3011,N_2782,N_2801);
or U3012 (N_3012,N_2578,N_2567);
nor U3013 (N_3013,N_2737,N_2772);
nand U3014 (N_3014,N_2562,N_2694);
nor U3015 (N_3015,N_2512,N_2731);
nand U3016 (N_3016,N_2533,N_2758);
nor U3017 (N_3017,N_2940,N_2796);
nor U3018 (N_3018,N_2552,N_2554);
xor U3019 (N_3019,N_2910,N_2707);
xor U3020 (N_3020,N_2955,N_2629);
nand U3021 (N_3021,N_2844,N_2899);
or U3022 (N_3022,N_2762,N_2996);
xor U3023 (N_3023,N_2814,N_2886);
nand U3024 (N_3024,N_2682,N_2756);
or U3025 (N_3025,N_2654,N_2861);
or U3026 (N_3026,N_2866,N_2744);
xnor U3027 (N_3027,N_2676,N_2712);
xor U3028 (N_3028,N_2865,N_2537);
or U3029 (N_3029,N_2600,N_2661);
and U3030 (N_3030,N_2528,N_2810);
nand U3031 (N_3031,N_2568,N_2767);
or U3032 (N_3032,N_2757,N_2729);
and U3033 (N_3033,N_2859,N_2559);
or U3034 (N_3034,N_2594,N_2690);
or U3035 (N_3035,N_2799,N_2970);
and U3036 (N_3036,N_2705,N_2632);
xnor U3037 (N_3037,N_2995,N_2623);
nand U3038 (N_3038,N_2991,N_2900);
or U3039 (N_3039,N_2691,N_2887);
nand U3040 (N_3040,N_2603,N_2986);
or U3041 (N_3041,N_2523,N_2922);
and U3042 (N_3042,N_2888,N_2826);
nor U3043 (N_3043,N_2583,N_2725);
nand U3044 (N_3044,N_2842,N_2863);
nor U3045 (N_3045,N_2630,N_2589);
nand U3046 (N_3046,N_2823,N_2565);
nor U3047 (N_3047,N_2873,N_2638);
and U3048 (N_3048,N_2961,N_2500);
and U3049 (N_3049,N_2716,N_2531);
xnor U3050 (N_3050,N_2677,N_2893);
and U3051 (N_3051,N_2896,N_2805);
or U3052 (N_3052,N_2972,N_2645);
and U3053 (N_3053,N_2894,N_2585);
xnor U3054 (N_3054,N_2543,N_2641);
xor U3055 (N_3055,N_2652,N_2546);
or U3056 (N_3056,N_2903,N_2878);
xnor U3057 (N_3057,N_2699,N_2526);
and U3058 (N_3058,N_2644,N_2975);
or U3059 (N_3059,N_2597,N_2722);
nand U3060 (N_3060,N_2858,N_2579);
or U3061 (N_3061,N_2720,N_2530);
or U3062 (N_3062,N_2981,N_2669);
nor U3063 (N_3063,N_2588,N_2934);
nand U3064 (N_3064,N_2704,N_2768);
nand U3065 (N_3065,N_2607,N_2511);
nand U3066 (N_3066,N_2697,N_2658);
nand U3067 (N_3067,N_2764,N_2908);
or U3068 (N_3068,N_2924,N_2785);
nand U3069 (N_3069,N_2804,N_2748);
nand U3070 (N_3070,N_2673,N_2634);
or U3071 (N_3071,N_2751,N_2990);
nor U3072 (N_3072,N_2501,N_2897);
and U3073 (N_3073,N_2733,N_2773);
or U3074 (N_3074,N_2879,N_2904);
nor U3075 (N_3075,N_2642,N_2602);
xnor U3076 (N_3076,N_2506,N_2633);
nand U3077 (N_3077,N_2891,N_2867);
or U3078 (N_3078,N_2920,N_2941);
nand U3079 (N_3079,N_2755,N_2754);
nand U3080 (N_3080,N_2587,N_2846);
nand U3081 (N_3081,N_2971,N_2693);
nor U3082 (N_3082,N_2529,N_2779);
nand U3083 (N_3083,N_2809,N_2932);
nor U3084 (N_3084,N_2957,N_2983);
xor U3085 (N_3085,N_2811,N_2540);
xor U3086 (N_3086,N_2752,N_2774);
nand U3087 (N_3087,N_2798,N_2794);
or U3088 (N_3088,N_2678,N_2636);
or U3089 (N_3089,N_2667,N_2734);
and U3090 (N_3090,N_2832,N_2592);
nor U3091 (N_3091,N_2787,N_2509);
xnor U3092 (N_3092,N_2890,N_2624);
nor U3093 (N_3093,N_2596,N_2692);
xnor U3094 (N_3094,N_2946,N_2706);
xnor U3095 (N_3095,N_2614,N_2640);
xor U3096 (N_3096,N_2982,N_2988);
xnor U3097 (N_3097,N_2542,N_2591);
xnor U3098 (N_3098,N_2848,N_2833);
nor U3099 (N_3099,N_2679,N_2545);
and U3100 (N_3100,N_2503,N_2837);
nor U3101 (N_3101,N_2876,N_2763);
or U3102 (N_3102,N_2558,N_2680);
nand U3103 (N_3103,N_2561,N_2571);
xor U3104 (N_3104,N_2675,N_2617);
or U3105 (N_3105,N_2637,N_2839);
nand U3106 (N_3106,N_2776,N_2732);
and U3107 (N_3107,N_2959,N_2821);
and U3108 (N_3108,N_2956,N_2939);
and U3109 (N_3109,N_2648,N_2777);
nand U3110 (N_3110,N_2980,N_2761);
nand U3111 (N_3111,N_2504,N_2831);
nor U3112 (N_3112,N_2539,N_2871);
and U3113 (N_3113,N_2812,N_2619);
nand U3114 (N_3114,N_2574,N_2760);
nor U3115 (N_3115,N_2918,N_2953);
nand U3116 (N_3116,N_2513,N_2827);
nor U3117 (N_3117,N_2917,N_2627);
and U3118 (N_3118,N_2551,N_2605);
nor U3119 (N_3119,N_2783,N_2874);
and U3120 (N_3120,N_2911,N_2958);
xor U3121 (N_3121,N_2989,N_2740);
and U3122 (N_3122,N_2789,N_2723);
and U3123 (N_3123,N_2780,N_2936);
xor U3124 (N_3124,N_2681,N_2853);
or U3125 (N_3125,N_2771,N_2881);
xnor U3126 (N_3126,N_2610,N_2807);
nand U3127 (N_3127,N_2517,N_2951);
or U3128 (N_3128,N_2854,N_2660);
or U3129 (N_3129,N_2584,N_2687);
xnor U3130 (N_3130,N_2670,N_2581);
nand U3131 (N_3131,N_2902,N_2913);
or U3132 (N_3132,N_2883,N_2836);
nor U3133 (N_3133,N_2599,N_2671);
and U3134 (N_3134,N_2626,N_2666);
xnor U3135 (N_3135,N_2895,N_2570);
nand U3136 (N_3136,N_2505,N_2514);
nor U3137 (N_3137,N_2672,N_2516);
nor U3138 (N_3138,N_2819,N_2905);
nand U3139 (N_3139,N_2822,N_2901);
or U3140 (N_3140,N_2689,N_2525);
or U3141 (N_3141,N_2736,N_2575);
and U3142 (N_3142,N_2820,N_2683);
nor U3143 (N_3143,N_2742,N_2993);
or U3144 (N_3144,N_2595,N_2829);
and U3145 (N_3145,N_2622,N_2938);
and U3146 (N_3146,N_2719,N_2727);
and U3147 (N_3147,N_2963,N_2611);
or U3148 (N_3148,N_2835,N_2869);
nor U3149 (N_3149,N_2745,N_2872);
nand U3150 (N_3150,N_2816,N_2862);
nor U3151 (N_3151,N_2977,N_2802);
and U3152 (N_3152,N_2766,N_2532);
xnor U3153 (N_3153,N_2519,N_2770);
nor U3154 (N_3154,N_2750,N_2639);
and U3155 (N_3155,N_2884,N_2850);
nor U3156 (N_3156,N_2527,N_2663);
xnor U3157 (N_3157,N_2928,N_2741);
or U3158 (N_3158,N_2618,N_2730);
nand U3159 (N_3159,N_2684,N_2717);
nor U3160 (N_3160,N_2714,N_2952);
and U3161 (N_3161,N_2549,N_2793);
xor U3162 (N_3162,N_2664,N_2643);
nor U3163 (N_3163,N_2696,N_2650);
nand U3164 (N_3164,N_2709,N_2984);
nand U3165 (N_3165,N_2948,N_2686);
and U3166 (N_3166,N_2702,N_2608);
nand U3167 (N_3167,N_2778,N_2753);
xnor U3168 (N_3168,N_2759,N_2838);
nor U3169 (N_3169,N_2724,N_2557);
nand U3170 (N_3170,N_2590,N_2978);
and U3171 (N_3171,N_2856,N_2803);
or U3172 (N_3172,N_2877,N_2535);
and U3173 (N_3173,N_2646,N_2815);
and U3174 (N_3174,N_2792,N_2933);
and U3175 (N_3175,N_2541,N_2668);
and U3176 (N_3176,N_2576,N_2653);
nor U3177 (N_3177,N_2828,N_2655);
nor U3178 (N_3178,N_2788,N_2651);
xor U3179 (N_3179,N_2797,N_2912);
nand U3180 (N_3180,N_2647,N_2864);
xnor U3181 (N_3181,N_2659,N_2715);
nand U3182 (N_3182,N_2572,N_2987);
or U3183 (N_3183,N_2889,N_2547);
and U3184 (N_3184,N_2808,N_2609);
and U3185 (N_3185,N_2840,N_2612);
or U3186 (N_3186,N_2577,N_2507);
nand U3187 (N_3187,N_2601,N_2847);
nor U3188 (N_3188,N_2875,N_2649);
xnor U3189 (N_3189,N_2931,N_2855);
and U3190 (N_3190,N_2781,N_2937);
xor U3191 (N_3191,N_2580,N_2915);
nor U3192 (N_3192,N_2845,N_2985);
xnor U3193 (N_3193,N_2502,N_2962);
nand U3194 (N_3194,N_2930,N_2965);
and U3195 (N_3195,N_2998,N_2906);
or U3196 (N_3196,N_2538,N_2746);
or U3197 (N_3197,N_2818,N_2999);
nand U3198 (N_3198,N_2631,N_2536);
nor U3199 (N_3199,N_2674,N_2573);
xnor U3200 (N_3200,N_2735,N_2942);
xnor U3201 (N_3201,N_2726,N_2784);
xor U3202 (N_3202,N_2738,N_2775);
nor U3203 (N_3203,N_2665,N_2698);
nand U3204 (N_3204,N_2966,N_2979);
xnor U3205 (N_3205,N_2919,N_2834);
and U3206 (N_3206,N_2510,N_2907);
xnor U3207 (N_3207,N_2976,N_2518);
and U3208 (N_3208,N_2695,N_2728);
nand U3209 (N_3209,N_2824,N_2870);
nand U3210 (N_3210,N_2949,N_2885);
and U3211 (N_3211,N_2974,N_2713);
and U3212 (N_3212,N_2593,N_2620);
or U3213 (N_3213,N_2524,N_2613);
or U3214 (N_3214,N_2769,N_2969);
and U3215 (N_3215,N_2521,N_2954);
xnor U3216 (N_3216,N_2656,N_2923);
xor U3217 (N_3217,N_2950,N_2947);
xor U3218 (N_3218,N_2968,N_2604);
and U3219 (N_3219,N_2943,N_2843);
and U3220 (N_3220,N_2564,N_2520);
xnor U3221 (N_3221,N_2566,N_2625);
nand U3222 (N_3222,N_2967,N_2786);
or U3223 (N_3223,N_2534,N_2563);
nand U3224 (N_3224,N_2701,N_2935);
xnor U3225 (N_3225,N_2851,N_2711);
nor U3226 (N_3226,N_2544,N_2662);
and U3227 (N_3227,N_2825,N_2550);
xnor U3228 (N_3228,N_2857,N_2628);
nand U3229 (N_3229,N_2721,N_2791);
nand U3230 (N_3230,N_2522,N_2582);
xnor U3231 (N_3231,N_2598,N_2635);
nand U3232 (N_3232,N_2841,N_2606);
nor U3233 (N_3233,N_2994,N_2795);
nand U3234 (N_3234,N_2703,N_2997);
or U3235 (N_3235,N_2892,N_2560);
nor U3236 (N_3236,N_2616,N_2555);
or U3237 (N_3237,N_2868,N_2852);
or U3238 (N_3238,N_2718,N_2914);
and U3239 (N_3239,N_2992,N_2765);
or U3240 (N_3240,N_2921,N_2548);
or U3241 (N_3241,N_2860,N_2964);
xor U3242 (N_3242,N_2945,N_2657);
nand U3243 (N_3243,N_2708,N_2556);
nand U3244 (N_3244,N_2710,N_2880);
xnor U3245 (N_3245,N_2800,N_2898);
nor U3246 (N_3246,N_2929,N_2508);
nand U3247 (N_3247,N_2621,N_2790);
nor U3248 (N_3248,N_2515,N_2569);
and U3249 (N_3249,N_2960,N_2806);
xor U3250 (N_3250,N_2995,N_2611);
nand U3251 (N_3251,N_2955,N_2831);
xnor U3252 (N_3252,N_2601,N_2524);
nand U3253 (N_3253,N_2763,N_2948);
nor U3254 (N_3254,N_2746,N_2680);
or U3255 (N_3255,N_2784,N_2823);
nand U3256 (N_3256,N_2534,N_2863);
nor U3257 (N_3257,N_2529,N_2911);
xor U3258 (N_3258,N_2994,N_2761);
xor U3259 (N_3259,N_2922,N_2888);
xor U3260 (N_3260,N_2617,N_2723);
nor U3261 (N_3261,N_2704,N_2701);
and U3262 (N_3262,N_2745,N_2631);
and U3263 (N_3263,N_2880,N_2989);
nor U3264 (N_3264,N_2954,N_2844);
nand U3265 (N_3265,N_2657,N_2881);
or U3266 (N_3266,N_2701,N_2897);
or U3267 (N_3267,N_2565,N_2560);
nor U3268 (N_3268,N_2501,N_2553);
or U3269 (N_3269,N_2819,N_2981);
nor U3270 (N_3270,N_2988,N_2896);
xnor U3271 (N_3271,N_2901,N_2549);
nor U3272 (N_3272,N_2941,N_2559);
nand U3273 (N_3273,N_2799,N_2671);
or U3274 (N_3274,N_2701,N_2623);
or U3275 (N_3275,N_2599,N_2561);
nand U3276 (N_3276,N_2864,N_2559);
and U3277 (N_3277,N_2782,N_2731);
nand U3278 (N_3278,N_2883,N_2954);
nand U3279 (N_3279,N_2552,N_2748);
nor U3280 (N_3280,N_2805,N_2960);
nand U3281 (N_3281,N_2617,N_2938);
nand U3282 (N_3282,N_2525,N_2723);
or U3283 (N_3283,N_2787,N_2919);
and U3284 (N_3284,N_2799,N_2786);
nor U3285 (N_3285,N_2871,N_2687);
nor U3286 (N_3286,N_2838,N_2861);
nor U3287 (N_3287,N_2773,N_2653);
or U3288 (N_3288,N_2774,N_2805);
or U3289 (N_3289,N_2538,N_2596);
and U3290 (N_3290,N_2915,N_2941);
and U3291 (N_3291,N_2599,N_2817);
and U3292 (N_3292,N_2551,N_2501);
nand U3293 (N_3293,N_2771,N_2781);
nand U3294 (N_3294,N_2507,N_2612);
nand U3295 (N_3295,N_2613,N_2958);
xor U3296 (N_3296,N_2992,N_2998);
xor U3297 (N_3297,N_2501,N_2560);
or U3298 (N_3298,N_2522,N_2717);
or U3299 (N_3299,N_2609,N_2773);
and U3300 (N_3300,N_2567,N_2886);
and U3301 (N_3301,N_2842,N_2644);
or U3302 (N_3302,N_2836,N_2732);
xor U3303 (N_3303,N_2595,N_2726);
xnor U3304 (N_3304,N_2580,N_2906);
nor U3305 (N_3305,N_2729,N_2921);
nand U3306 (N_3306,N_2598,N_2828);
and U3307 (N_3307,N_2853,N_2578);
and U3308 (N_3308,N_2551,N_2522);
nand U3309 (N_3309,N_2547,N_2903);
or U3310 (N_3310,N_2531,N_2597);
nand U3311 (N_3311,N_2924,N_2672);
xnor U3312 (N_3312,N_2791,N_2736);
and U3313 (N_3313,N_2752,N_2824);
nor U3314 (N_3314,N_2949,N_2592);
and U3315 (N_3315,N_2825,N_2969);
nor U3316 (N_3316,N_2623,N_2501);
nand U3317 (N_3317,N_2702,N_2630);
and U3318 (N_3318,N_2677,N_2542);
nand U3319 (N_3319,N_2728,N_2853);
nand U3320 (N_3320,N_2877,N_2580);
and U3321 (N_3321,N_2997,N_2528);
xor U3322 (N_3322,N_2712,N_2811);
xnor U3323 (N_3323,N_2806,N_2640);
nor U3324 (N_3324,N_2939,N_2934);
or U3325 (N_3325,N_2512,N_2932);
xor U3326 (N_3326,N_2775,N_2878);
nor U3327 (N_3327,N_2590,N_2689);
xnor U3328 (N_3328,N_2938,N_2681);
nand U3329 (N_3329,N_2522,N_2736);
nand U3330 (N_3330,N_2578,N_2850);
or U3331 (N_3331,N_2989,N_2656);
xnor U3332 (N_3332,N_2719,N_2866);
or U3333 (N_3333,N_2937,N_2555);
nand U3334 (N_3334,N_2925,N_2731);
nand U3335 (N_3335,N_2690,N_2816);
xor U3336 (N_3336,N_2511,N_2904);
or U3337 (N_3337,N_2663,N_2632);
nand U3338 (N_3338,N_2663,N_2820);
and U3339 (N_3339,N_2978,N_2531);
xnor U3340 (N_3340,N_2504,N_2735);
nand U3341 (N_3341,N_2737,N_2712);
xor U3342 (N_3342,N_2566,N_2951);
nand U3343 (N_3343,N_2672,N_2957);
or U3344 (N_3344,N_2562,N_2650);
or U3345 (N_3345,N_2850,N_2988);
and U3346 (N_3346,N_2746,N_2882);
nor U3347 (N_3347,N_2870,N_2644);
nor U3348 (N_3348,N_2517,N_2882);
or U3349 (N_3349,N_2648,N_2865);
xnor U3350 (N_3350,N_2852,N_2854);
nand U3351 (N_3351,N_2936,N_2652);
nor U3352 (N_3352,N_2704,N_2697);
nor U3353 (N_3353,N_2628,N_2920);
and U3354 (N_3354,N_2672,N_2804);
or U3355 (N_3355,N_2944,N_2890);
or U3356 (N_3356,N_2961,N_2696);
or U3357 (N_3357,N_2691,N_2722);
and U3358 (N_3358,N_2590,N_2775);
xnor U3359 (N_3359,N_2783,N_2646);
nand U3360 (N_3360,N_2956,N_2964);
or U3361 (N_3361,N_2650,N_2768);
nor U3362 (N_3362,N_2684,N_2785);
xnor U3363 (N_3363,N_2758,N_2585);
xor U3364 (N_3364,N_2727,N_2507);
nor U3365 (N_3365,N_2597,N_2997);
and U3366 (N_3366,N_2896,N_2571);
nand U3367 (N_3367,N_2611,N_2946);
xnor U3368 (N_3368,N_2507,N_2769);
and U3369 (N_3369,N_2508,N_2883);
and U3370 (N_3370,N_2992,N_2958);
nor U3371 (N_3371,N_2981,N_2820);
or U3372 (N_3372,N_2690,N_2744);
nor U3373 (N_3373,N_2965,N_2617);
and U3374 (N_3374,N_2886,N_2613);
nor U3375 (N_3375,N_2944,N_2870);
nor U3376 (N_3376,N_2890,N_2758);
or U3377 (N_3377,N_2869,N_2536);
xnor U3378 (N_3378,N_2682,N_2654);
xnor U3379 (N_3379,N_2627,N_2613);
xor U3380 (N_3380,N_2656,N_2685);
nor U3381 (N_3381,N_2503,N_2936);
nand U3382 (N_3382,N_2657,N_2544);
and U3383 (N_3383,N_2709,N_2701);
xor U3384 (N_3384,N_2610,N_2930);
nor U3385 (N_3385,N_2618,N_2765);
xnor U3386 (N_3386,N_2526,N_2917);
or U3387 (N_3387,N_2871,N_2872);
or U3388 (N_3388,N_2847,N_2650);
or U3389 (N_3389,N_2568,N_2532);
xor U3390 (N_3390,N_2884,N_2938);
nor U3391 (N_3391,N_2973,N_2510);
nor U3392 (N_3392,N_2808,N_2824);
nor U3393 (N_3393,N_2978,N_2977);
nand U3394 (N_3394,N_2500,N_2700);
xor U3395 (N_3395,N_2928,N_2667);
nor U3396 (N_3396,N_2607,N_2899);
or U3397 (N_3397,N_2772,N_2797);
and U3398 (N_3398,N_2990,N_2871);
nand U3399 (N_3399,N_2851,N_2765);
or U3400 (N_3400,N_2638,N_2859);
and U3401 (N_3401,N_2714,N_2963);
nand U3402 (N_3402,N_2639,N_2980);
nor U3403 (N_3403,N_2543,N_2683);
nand U3404 (N_3404,N_2825,N_2861);
or U3405 (N_3405,N_2725,N_2930);
xor U3406 (N_3406,N_2964,N_2574);
xnor U3407 (N_3407,N_2928,N_2633);
xnor U3408 (N_3408,N_2678,N_2599);
nor U3409 (N_3409,N_2677,N_2974);
xor U3410 (N_3410,N_2569,N_2889);
nand U3411 (N_3411,N_2794,N_2570);
and U3412 (N_3412,N_2984,N_2731);
and U3413 (N_3413,N_2614,N_2516);
or U3414 (N_3414,N_2933,N_2604);
and U3415 (N_3415,N_2907,N_2536);
nand U3416 (N_3416,N_2938,N_2654);
nand U3417 (N_3417,N_2756,N_2986);
nand U3418 (N_3418,N_2577,N_2900);
or U3419 (N_3419,N_2647,N_2683);
and U3420 (N_3420,N_2987,N_2772);
nor U3421 (N_3421,N_2533,N_2915);
nand U3422 (N_3422,N_2844,N_2672);
nor U3423 (N_3423,N_2973,N_2731);
nand U3424 (N_3424,N_2937,N_2925);
xnor U3425 (N_3425,N_2848,N_2949);
or U3426 (N_3426,N_2572,N_2586);
xnor U3427 (N_3427,N_2812,N_2748);
or U3428 (N_3428,N_2536,N_2696);
or U3429 (N_3429,N_2991,N_2804);
xor U3430 (N_3430,N_2753,N_2665);
xor U3431 (N_3431,N_2666,N_2916);
and U3432 (N_3432,N_2923,N_2916);
or U3433 (N_3433,N_2651,N_2886);
nand U3434 (N_3434,N_2795,N_2792);
and U3435 (N_3435,N_2719,N_2998);
and U3436 (N_3436,N_2757,N_2601);
and U3437 (N_3437,N_2915,N_2511);
nand U3438 (N_3438,N_2901,N_2921);
nand U3439 (N_3439,N_2550,N_2708);
nand U3440 (N_3440,N_2554,N_2954);
nand U3441 (N_3441,N_2625,N_2826);
and U3442 (N_3442,N_2770,N_2572);
nor U3443 (N_3443,N_2522,N_2503);
xnor U3444 (N_3444,N_2923,N_2822);
and U3445 (N_3445,N_2938,N_2661);
and U3446 (N_3446,N_2997,N_2902);
or U3447 (N_3447,N_2530,N_2760);
nand U3448 (N_3448,N_2954,N_2899);
xnor U3449 (N_3449,N_2866,N_2767);
nand U3450 (N_3450,N_2513,N_2887);
or U3451 (N_3451,N_2961,N_2748);
and U3452 (N_3452,N_2613,N_2876);
xnor U3453 (N_3453,N_2519,N_2508);
xnor U3454 (N_3454,N_2558,N_2709);
or U3455 (N_3455,N_2877,N_2953);
nand U3456 (N_3456,N_2545,N_2949);
and U3457 (N_3457,N_2966,N_2575);
xor U3458 (N_3458,N_2786,N_2663);
nor U3459 (N_3459,N_2664,N_2704);
xor U3460 (N_3460,N_2795,N_2562);
or U3461 (N_3461,N_2771,N_2953);
nand U3462 (N_3462,N_2991,N_2687);
and U3463 (N_3463,N_2636,N_2711);
nand U3464 (N_3464,N_2866,N_2606);
and U3465 (N_3465,N_2732,N_2888);
or U3466 (N_3466,N_2669,N_2631);
or U3467 (N_3467,N_2795,N_2572);
xor U3468 (N_3468,N_2519,N_2965);
nand U3469 (N_3469,N_2562,N_2739);
nand U3470 (N_3470,N_2938,N_2983);
nor U3471 (N_3471,N_2618,N_2586);
nand U3472 (N_3472,N_2866,N_2724);
nor U3473 (N_3473,N_2751,N_2674);
or U3474 (N_3474,N_2973,N_2942);
xor U3475 (N_3475,N_2936,N_2599);
or U3476 (N_3476,N_2862,N_2984);
and U3477 (N_3477,N_2906,N_2770);
or U3478 (N_3478,N_2506,N_2920);
and U3479 (N_3479,N_2805,N_2551);
or U3480 (N_3480,N_2588,N_2864);
nand U3481 (N_3481,N_2852,N_2984);
or U3482 (N_3482,N_2644,N_2527);
nand U3483 (N_3483,N_2838,N_2933);
nor U3484 (N_3484,N_2940,N_2538);
nand U3485 (N_3485,N_2734,N_2851);
and U3486 (N_3486,N_2886,N_2906);
nand U3487 (N_3487,N_2634,N_2910);
nand U3488 (N_3488,N_2800,N_2604);
xnor U3489 (N_3489,N_2893,N_2871);
or U3490 (N_3490,N_2547,N_2939);
xnor U3491 (N_3491,N_2537,N_2811);
and U3492 (N_3492,N_2680,N_2887);
xnor U3493 (N_3493,N_2755,N_2870);
nand U3494 (N_3494,N_2742,N_2597);
nor U3495 (N_3495,N_2688,N_2842);
and U3496 (N_3496,N_2928,N_2777);
nand U3497 (N_3497,N_2906,N_2705);
or U3498 (N_3498,N_2983,N_2729);
or U3499 (N_3499,N_2927,N_2506);
nor U3500 (N_3500,N_3248,N_3189);
and U3501 (N_3501,N_3169,N_3315);
and U3502 (N_3502,N_3026,N_3013);
and U3503 (N_3503,N_3359,N_3267);
nand U3504 (N_3504,N_3014,N_3203);
or U3505 (N_3505,N_3022,N_3141);
nor U3506 (N_3506,N_3133,N_3295);
nand U3507 (N_3507,N_3045,N_3184);
and U3508 (N_3508,N_3010,N_3447);
xnor U3509 (N_3509,N_3361,N_3050);
xnor U3510 (N_3510,N_3320,N_3216);
nand U3511 (N_3511,N_3490,N_3424);
or U3512 (N_3512,N_3180,N_3019);
or U3513 (N_3513,N_3164,N_3426);
and U3514 (N_3514,N_3163,N_3266);
or U3515 (N_3515,N_3365,N_3255);
nor U3516 (N_3516,N_3410,N_3431);
and U3517 (N_3517,N_3155,N_3479);
nor U3518 (N_3518,N_3339,N_3336);
or U3519 (N_3519,N_3448,N_3429);
nor U3520 (N_3520,N_3367,N_3331);
nand U3521 (N_3521,N_3226,N_3212);
xnor U3522 (N_3522,N_3389,N_3038);
xor U3523 (N_3523,N_3103,N_3222);
and U3524 (N_3524,N_3435,N_3159);
nor U3525 (N_3525,N_3296,N_3415);
and U3526 (N_3526,N_3351,N_3093);
xor U3527 (N_3527,N_3001,N_3033);
or U3528 (N_3528,N_3208,N_3258);
and U3529 (N_3529,N_3004,N_3337);
nand U3530 (N_3530,N_3385,N_3340);
nor U3531 (N_3531,N_3171,N_3003);
nand U3532 (N_3532,N_3275,N_3186);
nand U3533 (N_3533,N_3039,N_3236);
nand U3534 (N_3534,N_3006,N_3297);
nor U3535 (N_3535,N_3495,N_3356);
nor U3536 (N_3536,N_3127,N_3303);
xnor U3537 (N_3537,N_3412,N_3061);
xnor U3538 (N_3538,N_3404,N_3069);
nand U3539 (N_3539,N_3397,N_3288);
nor U3540 (N_3540,N_3423,N_3346);
xor U3541 (N_3541,N_3059,N_3342);
xnor U3542 (N_3542,N_3284,N_3441);
or U3543 (N_3543,N_3058,N_3480);
xor U3544 (N_3544,N_3371,N_3108);
or U3545 (N_3545,N_3172,N_3048);
nor U3546 (N_3546,N_3292,N_3129);
xnor U3547 (N_3547,N_3040,N_3273);
or U3548 (N_3548,N_3185,N_3017);
nor U3549 (N_3549,N_3140,N_3378);
or U3550 (N_3550,N_3433,N_3082);
nand U3551 (N_3551,N_3230,N_3009);
and U3552 (N_3552,N_3488,N_3400);
or U3553 (N_3553,N_3221,N_3406);
or U3554 (N_3554,N_3139,N_3213);
xnor U3555 (N_3555,N_3096,N_3386);
and U3556 (N_3556,N_3076,N_3244);
or U3557 (N_3557,N_3228,N_3262);
xnor U3558 (N_3558,N_3482,N_3047);
nand U3559 (N_3559,N_3131,N_3224);
and U3560 (N_3560,N_3478,N_3051);
nand U3561 (N_3561,N_3135,N_3408);
and U3562 (N_3562,N_3160,N_3193);
or U3563 (N_3563,N_3064,N_3483);
and U3564 (N_3564,N_3298,N_3115);
and U3565 (N_3565,N_3265,N_3138);
and U3566 (N_3566,N_3156,N_3421);
nor U3567 (N_3567,N_3062,N_3489);
nor U3568 (N_3568,N_3436,N_3143);
nor U3569 (N_3569,N_3344,N_3316);
or U3570 (N_3570,N_3176,N_3036);
nor U3571 (N_3571,N_3493,N_3387);
nand U3572 (N_3572,N_3375,N_3217);
xor U3573 (N_3573,N_3350,N_3179);
or U3574 (N_3574,N_3381,N_3335);
nor U3575 (N_3575,N_3465,N_3285);
and U3576 (N_3576,N_3041,N_3154);
xor U3577 (N_3577,N_3293,N_3084);
and U3578 (N_3578,N_3147,N_3321);
xnor U3579 (N_3579,N_3243,N_3027);
xnor U3580 (N_3580,N_3153,N_3025);
and U3581 (N_3581,N_3341,N_3268);
xnor U3582 (N_3582,N_3308,N_3332);
nor U3583 (N_3583,N_3121,N_3126);
nand U3584 (N_3584,N_3473,N_3496);
nor U3585 (N_3585,N_3376,N_3491);
or U3586 (N_3586,N_3130,N_3099);
nor U3587 (N_3587,N_3471,N_3328);
nor U3588 (N_3588,N_3205,N_3440);
and U3589 (N_3589,N_3043,N_3204);
nor U3590 (N_3590,N_3391,N_3007);
nor U3591 (N_3591,N_3401,N_3157);
nand U3592 (N_3592,N_3362,N_3072);
nor U3593 (N_3593,N_3149,N_3023);
or U3594 (N_3594,N_3369,N_3498);
or U3595 (N_3595,N_3366,N_3252);
nand U3596 (N_3596,N_3452,N_3283);
and U3597 (N_3597,N_3466,N_3111);
nand U3598 (N_3598,N_3263,N_3420);
or U3599 (N_3599,N_3458,N_3460);
nand U3600 (N_3600,N_3067,N_3449);
or U3601 (N_3601,N_3301,N_3112);
xor U3602 (N_3602,N_3167,N_3427);
or U3603 (N_3603,N_3097,N_3459);
nand U3604 (N_3604,N_3246,N_3322);
nand U3605 (N_3605,N_3233,N_3110);
nand U3606 (N_3606,N_3188,N_3355);
or U3607 (N_3607,N_3462,N_3291);
nor U3608 (N_3608,N_3150,N_3117);
nand U3609 (N_3609,N_3383,N_3286);
nand U3610 (N_3610,N_3242,N_3046);
or U3611 (N_3611,N_3005,N_3271);
and U3612 (N_3612,N_3409,N_3118);
nand U3613 (N_3613,N_3403,N_3486);
nand U3614 (N_3614,N_3054,N_3313);
nor U3615 (N_3615,N_3497,N_3094);
nand U3616 (N_3616,N_3183,N_3100);
nand U3617 (N_3617,N_3148,N_3077);
nand U3618 (N_3618,N_3021,N_3114);
and U3619 (N_3619,N_3227,N_3095);
or U3620 (N_3620,N_3090,N_3294);
nand U3621 (N_3621,N_3442,N_3463);
xnor U3622 (N_3622,N_3310,N_3151);
or U3623 (N_3623,N_3398,N_3124);
nor U3624 (N_3624,N_3457,N_3254);
or U3625 (N_3625,N_3201,N_3210);
and U3626 (N_3626,N_3231,N_3195);
xnor U3627 (N_3627,N_3395,N_3166);
nand U3628 (N_3628,N_3128,N_3334);
nor U3629 (N_3629,N_3261,N_3053);
xnor U3630 (N_3630,N_3287,N_3079);
xnor U3631 (N_3631,N_3187,N_3085);
or U3632 (N_3632,N_3223,N_3312);
and U3633 (N_3633,N_3469,N_3134);
nand U3634 (N_3634,N_3065,N_3309);
nor U3635 (N_3635,N_3029,N_3152);
xnor U3636 (N_3636,N_3345,N_3178);
or U3637 (N_3637,N_3274,N_3434);
or U3638 (N_3638,N_3439,N_3063);
or U3639 (N_3639,N_3073,N_3354);
xnor U3640 (N_3640,N_3087,N_3414);
xor U3641 (N_3641,N_3107,N_3030);
nor U3642 (N_3642,N_3468,N_3250);
or U3643 (N_3643,N_3174,N_3113);
or U3644 (N_3644,N_3158,N_3240);
nor U3645 (N_3645,N_3372,N_3136);
xor U3646 (N_3646,N_3052,N_3206);
or U3647 (N_3647,N_3422,N_3215);
or U3648 (N_3648,N_3338,N_3477);
xor U3649 (N_3649,N_3417,N_3430);
xnor U3650 (N_3650,N_3137,N_3333);
nor U3651 (N_3651,N_3349,N_3437);
and U3652 (N_3652,N_3330,N_3481);
and U3653 (N_3653,N_3390,N_3299);
xor U3654 (N_3654,N_3235,N_3253);
or U3655 (N_3655,N_3011,N_3081);
nand U3656 (N_3656,N_3306,N_3125);
and U3657 (N_3657,N_3144,N_3234);
nor U3658 (N_3658,N_3220,N_3015);
and U3659 (N_3659,N_3008,N_3419);
xnor U3660 (N_3660,N_3088,N_3120);
xnor U3661 (N_3661,N_3453,N_3277);
or U3662 (N_3662,N_3380,N_3194);
and U3663 (N_3663,N_3492,N_3162);
or U3664 (N_3664,N_3199,N_3476);
xor U3665 (N_3665,N_3302,N_3499);
nor U3666 (N_3666,N_3105,N_3374);
and U3667 (N_3667,N_3360,N_3260);
xor U3668 (N_3668,N_3211,N_3307);
xor U3669 (N_3669,N_3425,N_3405);
nor U3670 (N_3670,N_3413,N_3247);
and U3671 (N_3671,N_3239,N_3494);
nand U3672 (N_3672,N_3057,N_3200);
nor U3673 (N_3673,N_3122,N_3173);
xor U3674 (N_3674,N_3259,N_3074);
or U3675 (N_3675,N_3445,N_3384);
xor U3676 (N_3676,N_3289,N_3470);
nand U3677 (N_3677,N_3080,N_3024);
and U3678 (N_3678,N_3418,N_3256);
xnor U3679 (N_3679,N_3232,N_3218);
or U3680 (N_3680,N_3348,N_3245);
xor U3681 (N_3681,N_3379,N_3055);
nand U3682 (N_3682,N_3060,N_3300);
or U3683 (N_3683,N_3446,N_3323);
and U3684 (N_3684,N_3407,N_3119);
nand U3685 (N_3685,N_3329,N_3165);
nand U3686 (N_3686,N_3035,N_3443);
xor U3687 (N_3687,N_3388,N_3270);
xnor U3688 (N_3688,N_3311,N_3197);
nand U3689 (N_3689,N_3319,N_3363);
and U3690 (N_3690,N_3382,N_3209);
nor U3691 (N_3691,N_3091,N_3318);
nand U3692 (N_3692,N_3432,N_3000);
or U3693 (N_3693,N_3214,N_3392);
and U3694 (N_3694,N_3190,N_3416);
and U3695 (N_3695,N_3237,N_3281);
xnor U3696 (N_3696,N_3475,N_3402);
xor U3697 (N_3697,N_3279,N_3106);
xor U3698 (N_3698,N_3347,N_3399);
xnor U3699 (N_3699,N_3450,N_3451);
nor U3700 (N_3700,N_3317,N_3394);
nor U3701 (N_3701,N_3467,N_3264);
or U3702 (N_3702,N_3358,N_3002);
or U3703 (N_3703,N_3249,N_3191);
and U3704 (N_3704,N_3049,N_3198);
or U3705 (N_3705,N_3364,N_3377);
nand U3706 (N_3706,N_3086,N_3168);
or U3707 (N_3707,N_3474,N_3042);
nand U3708 (N_3708,N_3028,N_3177);
and U3709 (N_3709,N_3037,N_3304);
xnor U3710 (N_3710,N_3428,N_3464);
or U3711 (N_3711,N_3083,N_3327);
or U3712 (N_3712,N_3207,N_3098);
nor U3713 (N_3713,N_3225,N_3444);
nand U3714 (N_3714,N_3132,N_3101);
nand U3715 (N_3715,N_3078,N_3182);
nand U3716 (N_3716,N_3070,N_3251);
nand U3717 (N_3717,N_3229,N_3326);
and U3718 (N_3718,N_3370,N_3343);
nor U3719 (N_3719,N_3487,N_3305);
nand U3720 (N_3720,N_3280,N_3196);
nand U3721 (N_3721,N_3170,N_3241);
or U3722 (N_3722,N_3109,N_3357);
and U3723 (N_3723,N_3068,N_3352);
nand U3724 (N_3724,N_3373,N_3012);
and U3725 (N_3725,N_3145,N_3123);
nor U3726 (N_3726,N_3353,N_3438);
xnor U3727 (N_3727,N_3456,N_3142);
xor U3728 (N_3728,N_3238,N_3272);
xor U3729 (N_3729,N_3102,N_3146);
or U3730 (N_3730,N_3368,N_3325);
and U3731 (N_3731,N_3269,N_3089);
and U3732 (N_3732,N_3018,N_3219);
xnor U3733 (N_3733,N_3393,N_3104);
nor U3734 (N_3734,N_3181,N_3202);
xnor U3735 (N_3735,N_3016,N_3192);
and U3736 (N_3736,N_3276,N_3071);
nand U3737 (N_3737,N_3075,N_3454);
nand U3738 (N_3738,N_3290,N_3324);
xnor U3739 (N_3739,N_3455,N_3034);
nor U3740 (N_3740,N_3175,N_3032);
nor U3741 (N_3741,N_3257,N_3472);
xnor U3742 (N_3742,N_3116,N_3396);
nand U3743 (N_3743,N_3411,N_3092);
or U3744 (N_3744,N_3020,N_3161);
xnor U3745 (N_3745,N_3056,N_3066);
nor U3746 (N_3746,N_3484,N_3485);
xnor U3747 (N_3747,N_3044,N_3278);
nand U3748 (N_3748,N_3031,N_3282);
nand U3749 (N_3749,N_3461,N_3314);
xnor U3750 (N_3750,N_3142,N_3092);
nand U3751 (N_3751,N_3123,N_3459);
and U3752 (N_3752,N_3365,N_3484);
nor U3753 (N_3753,N_3107,N_3048);
xnor U3754 (N_3754,N_3152,N_3467);
nand U3755 (N_3755,N_3483,N_3083);
or U3756 (N_3756,N_3327,N_3255);
nand U3757 (N_3757,N_3150,N_3115);
or U3758 (N_3758,N_3316,N_3079);
or U3759 (N_3759,N_3107,N_3366);
nor U3760 (N_3760,N_3174,N_3202);
nor U3761 (N_3761,N_3073,N_3175);
and U3762 (N_3762,N_3380,N_3263);
or U3763 (N_3763,N_3437,N_3463);
nor U3764 (N_3764,N_3208,N_3322);
xnor U3765 (N_3765,N_3034,N_3078);
nor U3766 (N_3766,N_3264,N_3435);
and U3767 (N_3767,N_3308,N_3289);
nand U3768 (N_3768,N_3363,N_3141);
or U3769 (N_3769,N_3309,N_3031);
and U3770 (N_3770,N_3415,N_3023);
xor U3771 (N_3771,N_3099,N_3412);
nand U3772 (N_3772,N_3094,N_3380);
nand U3773 (N_3773,N_3265,N_3209);
xor U3774 (N_3774,N_3337,N_3042);
nand U3775 (N_3775,N_3265,N_3339);
nor U3776 (N_3776,N_3465,N_3019);
nor U3777 (N_3777,N_3197,N_3132);
or U3778 (N_3778,N_3050,N_3473);
or U3779 (N_3779,N_3365,N_3296);
xor U3780 (N_3780,N_3428,N_3397);
and U3781 (N_3781,N_3459,N_3052);
and U3782 (N_3782,N_3163,N_3046);
or U3783 (N_3783,N_3166,N_3432);
nor U3784 (N_3784,N_3006,N_3266);
nor U3785 (N_3785,N_3283,N_3060);
or U3786 (N_3786,N_3484,N_3205);
xnor U3787 (N_3787,N_3395,N_3234);
or U3788 (N_3788,N_3128,N_3062);
nor U3789 (N_3789,N_3255,N_3166);
or U3790 (N_3790,N_3415,N_3495);
xor U3791 (N_3791,N_3240,N_3404);
or U3792 (N_3792,N_3177,N_3475);
nor U3793 (N_3793,N_3288,N_3484);
nor U3794 (N_3794,N_3222,N_3164);
xnor U3795 (N_3795,N_3387,N_3118);
nor U3796 (N_3796,N_3213,N_3281);
and U3797 (N_3797,N_3190,N_3341);
and U3798 (N_3798,N_3339,N_3226);
nand U3799 (N_3799,N_3329,N_3110);
or U3800 (N_3800,N_3035,N_3428);
and U3801 (N_3801,N_3087,N_3240);
and U3802 (N_3802,N_3041,N_3436);
nand U3803 (N_3803,N_3320,N_3483);
or U3804 (N_3804,N_3016,N_3434);
or U3805 (N_3805,N_3189,N_3430);
or U3806 (N_3806,N_3026,N_3295);
nor U3807 (N_3807,N_3321,N_3265);
and U3808 (N_3808,N_3404,N_3419);
nand U3809 (N_3809,N_3148,N_3226);
nor U3810 (N_3810,N_3179,N_3072);
nor U3811 (N_3811,N_3159,N_3042);
nor U3812 (N_3812,N_3171,N_3286);
or U3813 (N_3813,N_3368,N_3314);
or U3814 (N_3814,N_3213,N_3136);
nand U3815 (N_3815,N_3103,N_3400);
nand U3816 (N_3816,N_3306,N_3052);
xor U3817 (N_3817,N_3195,N_3378);
and U3818 (N_3818,N_3268,N_3310);
nand U3819 (N_3819,N_3386,N_3291);
xor U3820 (N_3820,N_3332,N_3127);
nand U3821 (N_3821,N_3257,N_3173);
nand U3822 (N_3822,N_3049,N_3061);
and U3823 (N_3823,N_3485,N_3421);
xnor U3824 (N_3824,N_3008,N_3357);
nand U3825 (N_3825,N_3247,N_3497);
nor U3826 (N_3826,N_3003,N_3125);
or U3827 (N_3827,N_3120,N_3482);
and U3828 (N_3828,N_3232,N_3017);
nand U3829 (N_3829,N_3253,N_3000);
and U3830 (N_3830,N_3133,N_3289);
nand U3831 (N_3831,N_3202,N_3381);
or U3832 (N_3832,N_3067,N_3008);
or U3833 (N_3833,N_3158,N_3297);
xnor U3834 (N_3834,N_3449,N_3117);
or U3835 (N_3835,N_3420,N_3018);
or U3836 (N_3836,N_3053,N_3214);
and U3837 (N_3837,N_3017,N_3008);
nand U3838 (N_3838,N_3022,N_3265);
nand U3839 (N_3839,N_3403,N_3325);
or U3840 (N_3840,N_3116,N_3182);
nand U3841 (N_3841,N_3018,N_3269);
nor U3842 (N_3842,N_3359,N_3246);
nand U3843 (N_3843,N_3250,N_3014);
nand U3844 (N_3844,N_3293,N_3285);
xor U3845 (N_3845,N_3116,N_3402);
xor U3846 (N_3846,N_3461,N_3438);
xnor U3847 (N_3847,N_3493,N_3366);
xor U3848 (N_3848,N_3282,N_3008);
xor U3849 (N_3849,N_3336,N_3392);
xnor U3850 (N_3850,N_3018,N_3432);
and U3851 (N_3851,N_3265,N_3331);
and U3852 (N_3852,N_3114,N_3333);
nor U3853 (N_3853,N_3421,N_3455);
or U3854 (N_3854,N_3400,N_3089);
and U3855 (N_3855,N_3218,N_3032);
or U3856 (N_3856,N_3030,N_3047);
and U3857 (N_3857,N_3350,N_3365);
nand U3858 (N_3858,N_3245,N_3137);
and U3859 (N_3859,N_3197,N_3155);
xnor U3860 (N_3860,N_3446,N_3075);
nand U3861 (N_3861,N_3449,N_3289);
nand U3862 (N_3862,N_3350,N_3150);
nand U3863 (N_3863,N_3302,N_3267);
xnor U3864 (N_3864,N_3082,N_3360);
or U3865 (N_3865,N_3171,N_3179);
nand U3866 (N_3866,N_3058,N_3400);
or U3867 (N_3867,N_3380,N_3169);
xor U3868 (N_3868,N_3346,N_3167);
nor U3869 (N_3869,N_3258,N_3084);
nor U3870 (N_3870,N_3430,N_3492);
xor U3871 (N_3871,N_3081,N_3393);
nand U3872 (N_3872,N_3261,N_3498);
nand U3873 (N_3873,N_3205,N_3430);
xnor U3874 (N_3874,N_3489,N_3047);
nor U3875 (N_3875,N_3430,N_3401);
and U3876 (N_3876,N_3094,N_3488);
xnor U3877 (N_3877,N_3030,N_3086);
nor U3878 (N_3878,N_3115,N_3245);
xor U3879 (N_3879,N_3259,N_3362);
nand U3880 (N_3880,N_3277,N_3473);
nand U3881 (N_3881,N_3412,N_3359);
nand U3882 (N_3882,N_3320,N_3363);
xor U3883 (N_3883,N_3364,N_3264);
or U3884 (N_3884,N_3360,N_3136);
and U3885 (N_3885,N_3368,N_3077);
nor U3886 (N_3886,N_3001,N_3158);
or U3887 (N_3887,N_3044,N_3161);
and U3888 (N_3888,N_3280,N_3363);
or U3889 (N_3889,N_3089,N_3257);
or U3890 (N_3890,N_3284,N_3181);
or U3891 (N_3891,N_3297,N_3457);
xor U3892 (N_3892,N_3394,N_3028);
xnor U3893 (N_3893,N_3475,N_3179);
and U3894 (N_3894,N_3380,N_3178);
xnor U3895 (N_3895,N_3104,N_3285);
nand U3896 (N_3896,N_3408,N_3452);
nor U3897 (N_3897,N_3337,N_3494);
or U3898 (N_3898,N_3255,N_3273);
or U3899 (N_3899,N_3318,N_3322);
nand U3900 (N_3900,N_3072,N_3097);
nor U3901 (N_3901,N_3223,N_3436);
and U3902 (N_3902,N_3091,N_3307);
xor U3903 (N_3903,N_3156,N_3414);
and U3904 (N_3904,N_3252,N_3423);
nand U3905 (N_3905,N_3004,N_3194);
nand U3906 (N_3906,N_3143,N_3077);
xor U3907 (N_3907,N_3215,N_3154);
nor U3908 (N_3908,N_3021,N_3096);
nand U3909 (N_3909,N_3490,N_3393);
xor U3910 (N_3910,N_3219,N_3072);
or U3911 (N_3911,N_3178,N_3208);
nand U3912 (N_3912,N_3160,N_3166);
or U3913 (N_3913,N_3219,N_3226);
nor U3914 (N_3914,N_3292,N_3089);
xnor U3915 (N_3915,N_3209,N_3263);
nand U3916 (N_3916,N_3014,N_3348);
or U3917 (N_3917,N_3315,N_3018);
nor U3918 (N_3918,N_3267,N_3129);
nand U3919 (N_3919,N_3279,N_3227);
nand U3920 (N_3920,N_3281,N_3488);
nand U3921 (N_3921,N_3350,N_3073);
nor U3922 (N_3922,N_3243,N_3129);
nor U3923 (N_3923,N_3267,N_3336);
nand U3924 (N_3924,N_3150,N_3483);
nand U3925 (N_3925,N_3343,N_3143);
nand U3926 (N_3926,N_3088,N_3232);
and U3927 (N_3927,N_3247,N_3480);
and U3928 (N_3928,N_3147,N_3202);
nor U3929 (N_3929,N_3012,N_3124);
nand U3930 (N_3930,N_3420,N_3264);
or U3931 (N_3931,N_3064,N_3130);
and U3932 (N_3932,N_3229,N_3355);
nor U3933 (N_3933,N_3046,N_3257);
or U3934 (N_3934,N_3350,N_3356);
or U3935 (N_3935,N_3263,N_3085);
nand U3936 (N_3936,N_3339,N_3095);
and U3937 (N_3937,N_3166,N_3477);
nand U3938 (N_3938,N_3255,N_3015);
xor U3939 (N_3939,N_3045,N_3485);
or U3940 (N_3940,N_3280,N_3337);
xor U3941 (N_3941,N_3127,N_3115);
or U3942 (N_3942,N_3296,N_3290);
nand U3943 (N_3943,N_3364,N_3205);
nor U3944 (N_3944,N_3453,N_3146);
xnor U3945 (N_3945,N_3265,N_3137);
xnor U3946 (N_3946,N_3250,N_3072);
nand U3947 (N_3947,N_3402,N_3028);
and U3948 (N_3948,N_3224,N_3102);
and U3949 (N_3949,N_3068,N_3464);
nand U3950 (N_3950,N_3428,N_3354);
or U3951 (N_3951,N_3081,N_3083);
or U3952 (N_3952,N_3066,N_3021);
or U3953 (N_3953,N_3366,N_3125);
or U3954 (N_3954,N_3131,N_3236);
nand U3955 (N_3955,N_3411,N_3393);
xnor U3956 (N_3956,N_3260,N_3320);
or U3957 (N_3957,N_3335,N_3474);
nand U3958 (N_3958,N_3191,N_3235);
nor U3959 (N_3959,N_3434,N_3272);
and U3960 (N_3960,N_3318,N_3242);
and U3961 (N_3961,N_3216,N_3363);
and U3962 (N_3962,N_3147,N_3287);
nand U3963 (N_3963,N_3156,N_3309);
or U3964 (N_3964,N_3126,N_3201);
nand U3965 (N_3965,N_3332,N_3055);
or U3966 (N_3966,N_3309,N_3203);
and U3967 (N_3967,N_3005,N_3269);
or U3968 (N_3968,N_3182,N_3396);
and U3969 (N_3969,N_3043,N_3221);
nor U3970 (N_3970,N_3380,N_3122);
nor U3971 (N_3971,N_3276,N_3370);
nor U3972 (N_3972,N_3289,N_3218);
or U3973 (N_3973,N_3021,N_3260);
xor U3974 (N_3974,N_3491,N_3242);
nor U3975 (N_3975,N_3000,N_3269);
and U3976 (N_3976,N_3089,N_3336);
and U3977 (N_3977,N_3093,N_3053);
or U3978 (N_3978,N_3063,N_3130);
and U3979 (N_3979,N_3395,N_3042);
nor U3980 (N_3980,N_3159,N_3017);
nor U3981 (N_3981,N_3215,N_3205);
nand U3982 (N_3982,N_3389,N_3046);
or U3983 (N_3983,N_3161,N_3133);
or U3984 (N_3984,N_3171,N_3407);
nor U3985 (N_3985,N_3010,N_3467);
xor U3986 (N_3986,N_3139,N_3127);
and U3987 (N_3987,N_3125,N_3379);
nand U3988 (N_3988,N_3326,N_3242);
or U3989 (N_3989,N_3315,N_3256);
or U3990 (N_3990,N_3456,N_3315);
or U3991 (N_3991,N_3000,N_3053);
nor U3992 (N_3992,N_3070,N_3026);
nand U3993 (N_3993,N_3432,N_3170);
or U3994 (N_3994,N_3243,N_3060);
xor U3995 (N_3995,N_3444,N_3036);
nand U3996 (N_3996,N_3336,N_3278);
or U3997 (N_3997,N_3257,N_3421);
xnor U3998 (N_3998,N_3236,N_3416);
or U3999 (N_3999,N_3098,N_3019);
and U4000 (N_4000,N_3529,N_3612);
nor U4001 (N_4001,N_3822,N_3941);
or U4002 (N_4002,N_3886,N_3979);
or U4003 (N_4003,N_3732,N_3658);
nor U4004 (N_4004,N_3827,N_3974);
nor U4005 (N_4005,N_3729,N_3851);
nor U4006 (N_4006,N_3640,N_3889);
xnor U4007 (N_4007,N_3964,N_3701);
nor U4008 (N_4008,N_3998,N_3774);
xnor U4009 (N_4009,N_3662,N_3962);
or U4010 (N_4010,N_3965,N_3652);
and U4011 (N_4011,N_3504,N_3923);
nand U4012 (N_4012,N_3837,N_3800);
xor U4013 (N_4013,N_3747,N_3560);
nand U4014 (N_4014,N_3770,N_3871);
nand U4015 (N_4015,N_3509,N_3565);
or U4016 (N_4016,N_3860,N_3666);
or U4017 (N_4017,N_3826,N_3870);
nand U4018 (N_4018,N_3792,N_3862);
and U4019 (N_4019,N_3702,N_3823);
nor U4020 (N_4020,N_3634,N_3916);
or U4021 (N_4021,N_3879,N_3756);
nand U4022 (N_4022,N_3785,N_3734);
nor U4023 (N_4023,N_3989,N_3737);
nand U4024 (N_4024,N_3550,N_3901);
xor U4025 (N_4025,N_3523,N_3791);
nor U4026 (N_4026,N_3766,N_3745);
xnor U4027 (N_4027,N_3997,N_3781);
and U4028 (N_4028,N_3939,N_3794);
xor U4029 (N_4029,N_3543,N_3632);
nand U4030 (N_4030,N_3859,N_3542);
xor U4031 (N_4031,N_3709,N_3643);
nand U4032 (N_4032,N_3651,N_3602);
nor U4033 (N_4033,N_3842,N_3703);
or U4034 (N_4034,N_3668,N_3821);
nor U4035 (N_4035,N_3858,N_3783);
or U4036 (N_4036,N_3960,N_3637);
xor U4037 (N_4037,N_3516,N_3674);
xnor U4038 (N_4038,N_3510,N_3888);
or U4039 (N_4039,N_3636,N_3708);
nor U4040 (N_4040,N_3515,N_3679);
nand U4041 (N_4041,N_3804,N_3771);
nand U4042 (N_4042,N_3660,N_3948);
xnor U4043 (N_4043,N_3784,N_3790);
or U4044 (N_4044,N_3900,N_3743);
nor U4045 (N_4045,N_3567,N_3593);
nand U4046 (N_4046,N_3587,N_3868);
xnor U4047 (N_4047,N_3929,N_3852);
and U4048 (N_4048,N_3921,N_3564);
nor U4049 (N_4049,N_3548,N_3557);
xor U4050 (N_4050,N_3915,N_3810);
nand U4051 (N_4051,N_3677,N_3591);
nor U4052 (N_4052,N_3907,N_3749);
and U4053 (N_4053,N_3933,N_3838);
xnor U4054 (N_4054,N_3502,N_3511);
nor U4055 (N_4055,N_3973,N_3932);
nor U4056 (N_4056,N_3795,N_3902);
xnor U4057 (N_4057,N_3608,N_3891);
and U4058 (N_4058,N_3648,N_3811);
or U4059 (N_4059,N_3746,N_3569);
nand U4060 (N_4060,N_3622,N_3953);
and U4061 (N_4061,N_3796,N_3958);
and U4062 (N_4062,N_3914,N_3554);
xor U4063 (N_4063,N_3725,N_3806);
and U4064 (N_4064,N_3688,N_3667);
or U4065 (N_4065,N_3968,N_3903);
nor U4066 (N_4066,N_3620,N_3803);
nor U4067 (N_4067,N_3831,N_3911);
nand U4068 (N_4068,N_3546,N_3656);
xor U4069 (N_4069,N_3893,N_3683);
xor U4070 (N_4070,N_3573,N_3589);
nand U4071 (N_4071,N_3857,N_3697);
nand U4072 (N_4072,N_3592,N_3522);
nand U4073 (N_4073,N_3987,N_3559);
or U4074 (N_4074,N_3944,N_3954);
and U4075 (N_4075,N_3580,N_3536);
nand U4076 (N_4076,N_3887,N_3633);
nand U4077 (N_4077,N_3830,N_3981);
or U4078 (N_4078,N_3990,N_3758);
and U4079 (N_4079,N_3604,N_3969);
xnor U4080 (N_4080,N_3897,N_3614);
nand U4081 (N_4081,N_3575,N_3844);
or U4082 (N_4082,N_3527,N_3928);
nand U4083 (N_4083,N_3563,N_3676);
and U4084 (N_4084,N_3878,N_3556);
nand U4085 (N_4085,N_3584,N_3684);
or U4086 (N_4086,N_3751,N_3918);
nor U4087 (N_4087,N_3807,N_3805);
nor U4088 (N_4088,N_3707,N_3909);
or U4089 (N_4089,N_3999,N_3854);
nand U4090 (N_4090,N_3750,N_3936);
nand U4091 (N_4091,N_3711,N_3699);
and U4092 (N_4092,N_3541,N_3847);
nand U4093 (N_4093,N_3599,N_3943);
nand U4094 (N_4094,N_3736,N_3904);
or U4095 (N_4095,N_3812,N_3910);
and U4096 (N_4096,N_3621,N_3908);
and U4097 (N_4097,N_3874,N_3512);
or U4098 (N_4098,N_3663,N_3764);
and U4099 (N_4099,N_3585,N_3927);
nor U4100 (N_4100,N_3572,N_3789);
or U4101 (N_4101,N_3877,N_3996);
or U4102 (N_4102,N_3627,N_3582);
xor U4103 (N_4103,N_3884,N_3881);
nor U4104 (N_4104,N_3984,N_3947);
and U4105 (N_4105,N_3982,N_3514);
xor U4106 (N_4106,N_3742,N_3892);
or U4107 (N_4107,N_3978,N_3661);
xnor U4108 (N_4108,N_3664,N_3649);
nor U4109 (N_4109,N_3946,N_3988);
or U4110 (N_4110,N_3603,N_3722);
nand U4111 (N_4111,N_3906,N_3839);
nor U4112 (N_4112,N_3534,N_3972);
nand U4113 (N_4113,N_3595,N_3727);
or U4114 (N_4114,N_3720,N_3586);
nor U4115 (N_4115,N_3547,N_3519);
or U4116 (N_4116,N_3779,N_3617);
nand U4117 (N_4117,N_3925,N_3912);
nor U4118 (N_4118,N_3957,N_3562);
or U4119 (N_4119,N_3873,N_3829);
and U4120 (N_4120,N_3520,N_3672);
nor U4121 (N_4121,N_3930,N_3619);
nor U4122 (N_4122,N_3966,N_3850);
nand U4123 (N_4123,N_3815,N_3682);
nor U4124 (N_4124,N_3898,N_3931);
xor U4125 (N_4125,N_3865,N_3687);
nand U4126 (N_4126,N_3501,N_3977);
and U4127 (N_4127,N_3773,N_3517);
nor U4128 (N_4128,N_3721,N_3757);
nand U4129 (N_4129,N_3601,N_3882);
nand U4130 (N_4130,N_3814,N_3505);
xnor U4131 (N_4131,N_3880,N_3647);
nor U4132 (N_4132,N_3574,N_3583);
xnor U4133 (N_4133,N_3710,N_3872);
and U4134 (N_4134,N_3670,N_3924);
nand U4135 (N_4135,N_3626,N_3824);
nand U4136 (N_4136,N_3740,N_3638);
xnor U4137 (N_4137,N_3739,N_3995);
nand U4138 (N_4138,N_3855,N_3681);
nand U4139 (N_4139,N_3846,N_3856);
nor U4140 (N_4140,N_3919,N_3959);
and U4141 (N_4141,N_3600,N_3577);
nand U4142 (N_4142,N_3945,N_3700);
nand U4143 (N_4143,N_3561,N_3528);
nand U4144 (N_4144,N_3816,N_3728);
and U4145 (N_4145,N_3698,N_3993);
nand U4146 (N_4146,N_3864,N_3714);
xnor U4147 (N_4147,N_3926,N_3802);
and U4148 (N_4148,N_3705,N_3539);
and U4149 (N_4149,N_3994,N_3853);
and U4150 (N_4150,N_3980,N_3685);
and U4151 (N_4151,N_3738,N_3654);
nand U4152 (N_4152,N_3733,N_3956);
xnor U4153 (N_4153,N_3594,N_3691);
nor U4154 (N_4154,N_3678,N_3761);
nor U4155 (N_4155,N_3861,N_3799);
and U4156 (N_4156,N_3503,N_3537);
nand U4157 (N_4157,N_3639,N_3798);
nor U4158 (N_4158,N_3545,N_3975);
nand U4159 (N_4159,N_3793,N_3631);
xnor U4160 (N_4160,N_3843,N_3553);
xnor U4161 (N_4161,N_3935,N_3775);
xor U4162 (N_4162,N_3768,N_3992);
xor U4163 (N_4163,N_3835,N_3724);
nand U4164 (N_4164,N_3832,N_3748);
or U4165 (N_4165,N_3942,N_3950);
nand U4166 (N_4166,N_3610,N_3726);
and U4167 (N_4167,N_3730,N_3540);
nand U4168 (N_4168,N_3712,N_3611);
and U4169 (N_4169,N_3849,N_3646);
and U4170 (N_4170,N_3544,N_3778);
nand U4171 (N_4171,N_3955,N_3623);
xor U4172 (N_4172,N_3571,N_3665);
xor U4173 (N_4173,N_3976,N_3508);
nor U4174 (N_4174,N_3616,N_3890);
nor U4175 (N_4175,N_3716,N_3940);
nor U4176 (N_4176,N_3717,N_3922);
and U4177 (N_4177,N_3809,N_3876);
xor U4178 (N_4178,N_3963,N_3533);
and U4179 (N_4179,N_3971,N_3762);
or U4180 (N_4180,N_3776,N_3841);
nand U4181 (N_4181,N_3566,N_3613);
and U4182 (N_4182,N_3549,N_3767);
or U4183 (N_4183,N_3753,N_3820);
or U4184 (N_4184,N_3629,N_3744);
nor U4185 (N_4185,N_3624,N_3840);
and U4186 (N_4186,N_3513,N_3787);
or U4187 (N_4187,N_3695,N_3506);
nor U4188 (N_4188,N_3644,N_3895);
xnor U4189 (N_4189,N_3763,N_3741);
nor U4190 (N_4190,N_3780,N_3706);
nor U4191 (N_4191,N_3905,N_3769);
nand U4192 (N_4192,N_3524,N_3597);
or U4193 (N_4193,N_3680,N_3917);
nor U4194 (N_4194,N_3535,N_3570);
and U4195 (N_4195,N_3590,N_3719);
nand U4196 (N_4196,N_3568,N_3818);
or U4197 (N_4197,N_3689,N_3949);
and U4198 (N_4198,N_3713,N_3913);
nand U4199 (N_4199,N_3967,N_3635);
xor U4200 (N_4200,N_3754,N_3653);
nor U4201 (N_4201,N_3521,N_3836);
nor U4202 (N_4202,N_3828,N_3937);
nand U4203 (N_4203,N_3723,N_3645);
nor U4204 (N_4204,N_3531,N_3985);
and U4205 (N_4205,N_3525,N_3866);
or U4206 (N_4206,N_3755,N_3867);
xnor U4207 (N_4207,N_3983,N_3801);
xor U4208 (N_4208,N_3817,N_3938);
nand U4209 (N_4209,N_3615,N_3883);
nand U4210 (N_4210,N_3786,N_3777);
or U4211 (N_4211,N_3715,N_3552);
xor U4212 (N_4212,N_3692,N_3690);
nor U4213 (N_4213,N_3605,N_3551);
nor U4214 (N_4214,N_3788,N_3782);
or U4215 (N_4215,N_3628,N_3899);
and U4216 (N_4216,N_3759,N_3875);
nor U4217 (N_4217,N_3693,N_3704);
xnor U4218 (N_4218,N_3991,N_3869);
xor U4219 (N_4219,N_3833,N_3657);
xor U4220 (N_4220,N_3530,N_3641);
or U4221 (N_4221,N_3659,N_3538);
or U4222 (N_4222,N_3675,N_3834);
or U4223 (N_4223,N_3607,N_3673);
and U4224 (N_4224,N_3618,N_3718);
and U4225 (N_4225,N_3885,N_3696);
or U4226 (N_4226,N_3951,N_3500);
nand U4227 (N_4227,N_3848,N_3532);
or U4228 (N_4228,N_3797,N_3808);
nor U4229 (N_4229,N_3986,N_3819);
nand U4230 (N_4230,N_3894,N_3694);
nor U4231 (N_4231,N_3606,N_3558);
nand U4232 (N_4232,N_3518,N_3845);
or U4233 (N_4233,N_3669,N_3596);
nand U4234 (N_4234,N_3642,N_3579);
xor U4235 (N_4235,N_3507,N_3609);
and U4236 (N_4236,N_3735,N_3526);
xnor U4237 (N_4237,N_3952,N_3813);
xor U4238 (N_4238,N_3555,N_3731);
xnor U4239 (N_4239,N_3625,N_3760);
nand U4240 (N_4240,N_3863,N_3576);
or U4241 (N_4241,N_3650,N_3686);
nand U4242 (N_4242,N_3671,N_3934);
nand U4243 (N_4243,N_3655,N_3588);
nor U4244 (N_4244,N_3970,N_3920);
or U4245 (N_4245,N_3825,N_3581);
nand U4246 (N_4246,N_3896,N_3598);
and U4247 (N_4247,N_3752,N_3578);
nor U4248 (N_4248,N_3630,N_3765);
or U4249 (N_4249,N_3961,N_3772);
nor U4250 (N_4250,N_3701,N_3916);
xnor U4251 (N_4251,N_3977,N_3578);
and U4252 (N_4252,N_3862,N_3775);
and U4253 (N_4253,N_3633,N_3562);
and U4254 (N_4254,N_3783,N_3551);
nand U4255 (N_4255,N_3673,N_3816);
nor U4256 (N_4256,N_3589,N_3781);
xor U4257 (N_4257,N_3574,N_3521);
or U4258 (N_4258,N_3721,N_3891);
nand U4259 (N_4259,N_3707,N_3557);
nor U4260 (N_4260,N_3852,N_3804);
or U4261 (N_4261,N_3945,N_3704);
nand U4262 (N_4262,N_3939,N_3620);
xnor U4263 (N_4263,N_3523,N_3594);
nand U4264 (N_4264,N_3828,N_3507);
nand U4265 (N_4265,N_3920,N_3729);
xor U4266 (N_4266,N_3536,N_3659);
or U4267 (N_4267,N_3759,N_3855);
nor U4268 (N_4268,N_3702,N_3736);
xnor U4269 (N_4269,N_3840,N_3785);
nor U4270 (N_4270,N_3503,N_3867);
nand U4271 (N_4271,N_3517,N_3976);
and U4272 (N_4272,N_3898,N_3940);
xor U4273 (N_4273,N_3985,N_3779);
xor U4274 (N_4274,N_3819,N_3981);
or U4275 (N_4275,N_3796,N_3536);
xnor U4276 (N_4276,N_3937,N_3693);
xor U4277 (N_4277,N_3858,N_3710);
nand U4278 (N_4278,N_3759,N_3794);
nand U4279 (N_4279,N_3612,N_3599);
and U4280 (N_4280,N_3753,N_3945);
nor U4281 (N_4281,N_3960,N_3924);
xnor U4282 (N_4282,N_3538,N_3964);
nand U4283 (N_4283,N_3796,N_3747);
nand U4284 (N_4284,N_3910,N_3642);
nand U4285 (N_4285,N_3551,N_3615);
nand U4286 (N_4286,N_3601,N_3970);
or U4287 (N_4287,N_3876,N_3780);
nor U4288 (N_4288,N_3581,N_3611);
xor U4289 (N_4289,N_3916,N_3647);
or U4290 (N_4290,N_3957,N_3917);
or U4291 (N_4291,N_3668,N_3696);
nor U4292 (N_4292,N_3624,N_3860);
or U4293 (N_4293,N_3518,N_3868);
xor U4294 (N_4294,N_3778,N_3909);
nand U4295 (N_4295,N_3726,N_3601);
and U4296 (N_4296,N_3843,N_3747);
xnor U4297 (N_4297,N_3682,N_3785);
and U4298 (N_4298,N_3566,N_3802);
or U4299 (N_4299,N_3592,N_3561);
and U4300 (N_4300,N_3799,N_3896);
xor U4301 (N_4301,N_3597,N_3902);
nand U4302 (N_4302,N_3694,N_3501);
xor U4303 (N_4303,N_3776,N_3982);
and U4304 (N_4304,N_3963,N_3991);
xnor U4305 (N_4305,N_3680,N_3527);
nand U4306 (N_4306,N_3892,N_3712);
nand U4307 (N_4307,N_3724,N_3532);
and U4308 (N_4308,N_3610,N_3579);
nand U4309 (N_4309,N_3646,N_3508);
nor U4310 (N_4310,N_3800,N_3566);
nor U4311 (N_4311,N_3513,N_3554);
and U4312 (N_4312,N_3591,N_3759);
nor U4313 (N_4313,N_3519,N_3766);
or U4314 (N_4314,N_3724,N_3577);
and U4315 (N_4315,N_3728,N_3517);
nor U4316 (N_4316,N_3773,N_3644);
xnor U4317 (N_4317,N_3503,N_3746);
or U4318 (N_4318,N_3594,N_3618);
and U4319 (N_4319,N_3865,N_3816);
xor U4320 (N_4320,N_3629,N_3578);
and U4321 (N_4321,N_3658,N_3879);
and U4322 (N_4322,N_3881,N_3534);
nand U4323 (N_4323,N_3534,N_3917);
nand U4324 (N_4324,N_3797,N_3577);
nor U4325 (N_4325,N_3609,N_3893);
nor U4326 (N_4326,N_3635,N_3585);
nor U4327 (N_4327,N_3535,N_3854);
nand U4328 (N_4328,N_3676,N_3753);
and U4329 (N_4329,N_3577,N_3719);
nor U4330 (N_4330,N_3603,N_3519);
nand U4331 (N_4331,N_3847,N_3719);
nor U4332 (N_4332,N_3566,N_3845);
and U4333 (N_4333,N_3803,N_3685);
nor U4334 (N_4334,N_3538,N_3891);
and U4335 (N_4335,N_3622,N_3813);
or U4336 (N_4336,N_3765,N_3847);
nor U4337 (N_4337,N_3510,N_3753);
nor U4338 (N_4338,N_3999,N_3888);
nand U4339 (N_4339,N_3603,N_3629);
xor U4340 (N_4340,N_3869,N_3510);
or U4341 (N_4341,N_3689,N_3978);
nor U4342 (N_4342,N_3504,N_3866);
and U4343 (N_4343,N_3944,N_3712);
or U4344 (N_4344,N_3979,N_3659);
or U4345 (N_4345,N_3831,N_3703);
or U4346 (N_4346,N_3943,N_3869);
xnor U4347 (N_4347,N_3607,N_3728);
xor U4348 (N_4348,N_3582,N_3846);
nand U4349 (N_4349,N_3684,N_3567);
xnor U4350 (N_4350,N_3791,N_3744);
or U4351 (N_4351,N_3970,N_3688);
or U4352 (N_4352,N_3621,N_3832);
nand U4353 (N_4353,N_3913,N_3536);
nor U4354 (N_4354,N_3679,N_3523);
and U4355 (N_4355,N_3712,N_3839);
or U4356 (N_4356,N_3501,N_3792);
nand U4357 (N_4357,N_3517,N_3519);
or U4358 (N_4358,N_3892,N_3651);
nand U4359 (N_4359,N_3901,N_3629);
xor U4360 (N_4360,N_3930,N_3549);
xnor U4361 (N_4361,N_3586,N_3981);
nor U4362 (N_4362,N_3975,N_3942);
nor U4363 (N_4363,N_3705,N_3875);
and U4364 (N_4364,N_3956,N_3935);
nor U4365 (N_4365,N_3724,N_3662);
xnor U4366 (N_4366,N_3571,N_3910);
xnor U4367 (N_4367,N_3945,N_3999);
xor U4368 (N_4368,N_3760,N_3765);
nor U4369 (N_4369,N_3923,N_3647);
nor U4370 (N_4370,N_3568,N_3976);
nor U4371 (N_4371,N_3851,N_3599);
nand U4372 (N_4372,N_3777,N_3521);
xnor U4373 (N_4373,N_3705,N_3745);
nor U4374 (N_4374,N_3720,N_3591);
nor U4375 (N_4375,N_3698,N_3928);
nor U4376 (N_4376,N_3638,N_3898);
and U4377 (N_4377,N_3715,N_3623);
nor U4378 (N_4378,N_3701,N_3968);
or U4379 (N_4379,N_3976,N_3614);
nor U4380 (N_4380,N_3586,N_3640);
and U4381 (N_4381,N_3844,N_3615);
or U4382 (N_4382,N_3737,N_3947);
and U4383 (N_4383,N_3782,N_3818);
or U4384 (N_4384,N_3541,N_3586);
xnor U4385 (N_4385,N_3941,N_3672);
or U4386 (N_4386,N_3789,N_3750);
nor U4387 (N_4387,N_3742,N_3519);
nor U4388 (N_4388,N_3993,N_3749);
xor U4389 (N_4389,N_3515,N_3653);
xnor U4390 (N_4390,N_3896,N_3638);
nand U4391 (N_4391,N_3717,N_3888);
nand U4392 (N_4392,N_3726,N_3758);
and U4393 (N_4393,N_3718,N_3624);
nand U4394 (N_4394,N_3886,N_3672);
nor U4395 (N_4395,N_3555,N_3784);
nand U4396 (N_4396,N_3963,N_3941);
or U4397 (N_4397,N_3943,N_3951);
xor U4398 (N_4398,N_3548,N_3549);
nand U4399 (N_4399,N_3770,N_3863);
or U4400 (N_4400,N_3542,N_3996);
nor U4401 (N_4401,N_3743,N_3653);
nor U4402 (N_4402,N_3516,N_3705);
nand U4403 (N_4403,N_3565,N_3673);
or U4404 (N_4404,N_3512,N_3563);
nand U4405 (N_4405,N_3835,N_3935);
xnor U4406 (N_4406,N_3847,N_3877);
xor U4407 (N_4407,N_3919,N_3742);
nand U4408 (N_4408,N_3965,N_3926);
nor U4409 (N_4409,N_3638,N_3982);
or U4410 (N_4410,N_3636,N_3838);
nand U4411 (N_4411,N_3502,N_3581);
nand U4412 (N_4412,N_3615,N_3788);
xor U4413 (N_4413,N_3769,N_3941);
nor U4414 (N_4414,N_3714,N_3830);
nor U4415 (N_4415,N_3523,N_3945);
and U4416 (N_4416,N_3920,N_3755);
or U4417 (N_4417,N_3969,N_3516);
nand U4418 (N_4418,N_3676,N_3751);
and U4419 (N_4419,N_3538,N_3970);
or U4420 (N_4420,N_3976,N_3748);
xor U4421 (N_4421,N_3765,N_3638);
and U4422 (N_4422,N_3711,N_3695);
and U4423 (N_4423,N_3606,N_3727);
and U4424 (N_4424,N_3859,N_3882);
xor U4425 (N_4425,N_3823,N_3973);
xor U4426 (N_4426,N_3925,N_3847);
or U4427 (N_4427,N_3601,N_3959);
and U4428 (N_4428,N_3532,N_3755);
xor U4429 (N_4429,N_3624,N_3646);
xor U4430 (N_4430,N_3861,N_3679);
or U4431 (N_4431,N_3753,N_3562);
xor U4432 (N_4432,N_3996,N_3953);
and U4433 (N_4433,N_3807,N_3531);
nand U4434 (N_4434,N_3842,N_3667);
and U4435 (N_4435,N_3618,N_3950);
xor U4436 (N_4436,N_3751,N_3810);
and U4437 (N_4437,N_3615,N_3740);
nor U4438 (N_4438,N_3745,N_3618);
and U4439 (N_4439,N_3584,N_3919);
nor U4440 (N_4440,N_3829,N_3550);
nand U4441 (N_4441,N_3503,N_3562);
nand U4442 (N_4442,N_3921,N_3568);
and U4443 (N_4443,N_3759,N_3874);
nor U4444 (N_4444,N_3839,N_3543);
xor U4445 (N_4445,N_3763,N_3894);
or U4446 (N_4446,N_3900,N_3602);
nor U4447 (N_4447,N_3906,N_3880);
nand U4448 (N_4448,N_3924,N_3735);
and U4449 (N_4449,N_3906,N_3838);
nor U4450 (N_4450,N_3884,N_3746);
nor U4451 (N_4451,N_3629,N_3736);
and U4452 (N_4452,N_3729,N_3823);
and U4453 (N_4453,N_3966,N_3574);
or U4454 (N_4454,N_3554,N_3994);
xor U4455 (N_4455,N_3603,N_3667);
xor U4456 (N_4456,N_3562,N_3990);
xnor U4457 (N_4457,N_3748,N_3503);
or U4458 (N_4458,N_3806,N_3836);
xnor U4459 (N_4459,N_3606,N_3981);
nand U4460 (N_4460,N_3628,N_3831);
nand U4461 (N_4461,N_3941,N_3852);
and U4462 (N_4462,N_3618,N_3674);
nand U4463 (N_4463,N_3703,N_3933);
or U4464 (N_4464,N_3937,N_3891);
and U4465 (N_4465,N_3840,N_3735);
nor U4466 (N_4466,N_3654,N_3922);
nor U4467 (N_4467,N_3673,N_3711);
nor U4468 (N_4468,N_3705,N_3823);
nor U4469 (N_4469,N_3890,N_3571);
and U4470 (N_4470,N_3697,N_3874);
nor U4471 (N_4471,N_3504,N_3798);
nor U4472 (N_4472,N_3876,N_3629);
and U4473 (N_4473,N_3776,N_3975);
nor U4474 (N_4474,N_3830,N_3548);
or U4475 (N_4475,N_3735,N_3588);
nand U4476 (N_4476,N_3652,N_3892);
nor U4477 (N_4477,N_3665,N_3655);
nand U4478 (N_4478,N_3501,N_3918);
xor U4479 (N_4479,N_3822,N_3580);
and U4480 (N_4480,N_3886,N_3992);
nor U4481 (N_4481,N_3762,N_3852);
nor U4482 (N_4482,N_3984,N_3704);
or U4483 (N_4483,N_3924,N_3748);
xor U4484 (N_4484,N_3591,N_3776);
xor U4485 (N_4485,N_3733,N_3572);
and U4486 (N_4486,N_3742,N_3959);
and U4487 (N_4487,N_3729,N_3915);
nor U4488 (N_4488,N_3776,N_3567);
or U4489 (N_4489,N_3992,N_3713);
xor U4490 (N_4490,N_3816,N_3855);
nor U4491 (N_4491,N_3817,N_3582);
and U4492 (N_4492,N_3878,N_3733);
nand U4493 (N_4493,N_3604,N_3508);
nand U4494 (N_4494,N_3914,N_3961);
nand U4495 (N_4495,N_3929,N_3922);
xor U4496 (N_4496,N_3521,N_3906);
and U4497 (N_4497,N_3629,N_3880);
xor U4498 (N_4498,N_3983,N_3648);
xor U4499 (N_4499,N_3960,N_3554);
nor U4500 (N_4500,N_4154,N_4089);
and U4501 (N_4501,N_4477,N_4123);
and U4502 (N_4502,N_4458,N_4475);
xor U4503 (N_4503,N_4131,N_4230);
xnor U4504 (N_4504,N_4207,N_4020);
nand U4505 (N_4505,N_4085,N_4061);
or U4506 (N_4506,N_4428,N_4215);
or U4507 (N_4507,N_4030,N_4220);
nor U4508 (N_4508,N_4057,N_4361);
xor U4509 (N_4509,N_4111,N_4217);
xnor U4510 (N_4510,N_4375,N_4423);
xor U4511 (N_4511,N_4022,N_4434);
or U4512 (N_4512,N_4199,N_4024);
or U4513 (N_4513,N_4441,N_4415);
xnor U4514 (N_4514,N_4260,N_4334);
xnor U4515 (N_4515,N_4106,N_4476);
nor U4516 (N_4516,N_4234,N_4086);
and U4517 (N_4517,N_4093,N_4406);
nor U4518 (N_4518,N_4042,N_4281);
nor U4519 (N_4519,N_4147,N_4074);
xnor U4520 (N_4520,N_4311,N_4454);
or U4521 (N_4521,N_4425,N_4456);
nand U4522 (N_4522,N_4046,N_4376);
or U4523 (N_4523,N_4470,N_4305);
nor U4524 (N_4524,N_4318,N_4274);
nand U4525 (N_4525,N_4211,N_4254);
and U4526 (N_4526,N_4485,N_4065);
nor U4527 (N_4527,N_4180,N_4322);
and U4528 (N_4528,N_4262,N_4276);
xor U4529 (N_4529,N_4480,N_4269);
and U4530 (N_4530,N_4188,N_4248);
nor U4531 (N_4531,N_4080,N_4390);
or U4532 (N_4532,N_4295,N_4342);
nand U4533 (N_4533,N_4224,N_4320);
xnor U4534 (N_4534,N_4356,N_4031);
xnor U4535 (N_4535,N_4364,N_4142);
xor U4536 (N_4536,N_4279,N_4077);
xor U4537 (N_4537,N_4102,N_4383);
nor U4538 (N_4538,N_4385,N_4448);
xnor U4539 (N_4539,N_4256,N_4268);
xor U4540 (N_4540,N_4330,N_4007);
and U4541 (N_4541,N_4414,N_4003);
nand U4542 (N_4542,N_4328,N_4360);
nor U4543 (N_4543,N_4138,N_4422);
xor U4544 (N_4544,N_4097,N_4001);
nand U4545 (N_4545,N_4076,N_4208);
xnor U4546 (N_4546,N_4244,N_4405);
nor U4547 (N_4547,N_4150,N_4186);
nand U4548 (N_4548,N_4017,N_4229);
or U4549 (N_4549,N_4228,N_4047);
or U4550 (N_4550,N_4484,N_4430);
or U4551 (N_4551,N_4108,N_4298);
and U4552 (N_4552,N_4403,N_4416);
and U4553 (N_4553,N_4225,N_4253);
nand U4554 (N_4554,N_4049,N_4200);
nand U4555 (N_4555,N_4058,N_4408);
xnor U4556 (N_4556,N_4381,N_4034);
xor U4557 (N_4557,N_4117,N_4303);
xnor U4558 (N_4558,N_4148,N_4399);
or U4559 (N_4559,N_4005,N_4206);
nand U4560 (N_4560,N_4327,N_4349);
or U4561 (N_4561,N_4073,N_4446);
nor U4562 (N_4562,N_4026,N_4426);
nand U4563 (N_4563,N_4095,N_4407);
or U4564 (N_4564,N_4272,N_4099);
nor U4565 (N_4565,N_4395,N_4280);
or U4566 (N_4566,N_4339,N_4167);
xnor U4567 (N_4567,N_4120,N_4092);
and U4568 (N_4568,N_4310,N_4023);
xor U4569 (N_4569,N_4125,N_4323);
nor U4570 (N_4570,N_4198,N_4233);
and U4571 (N_4571,N_4402,N_4166);
nor U4572 (N_4572,N_4165,N_4341);
nor U4573 (N_4573,N_4453,N_4488);
nor U4574 (N_4574,N_4331,N_4210);
and U4575 (N_4575,N_4445,N_4014);
or U4576 (N_4576,N_4388,N_4384);
nand U4577 (N_4577,N_4245,N_4124);
and U4578 (N_4578,N_4185,N_4370);
and U4579 (N_4579,N_4401,N_4421);
xor U4580 (N_4580,N_4437,N_4343);
or U4581 (N_4581,N_4435,N_4292);
and U4582 (N_4582,N_4393,N_4240);
xnor U4583 (N_4583,N_4169,N_4377);
or U4584 (N_4584,N_4155,N_4235);
nor U4585 (N_4585,N_4372,N_4288);
nor U4586 (N_4586,N_4241,N_4359);
and U4587 (N_4587,N_4460,N_4491);
xor U4588 (N_4588,N_4348,N_4033);
and U4589 (N_4589,N_4252,N_4151);
nor U4590 (N_4590,N_4338,N_4496);
nor U4591 (N_4591,N_4152,N_4139);
nand U4592 (N_4592,N_4038,N_4010);
and U4593 (N_4593,N_4202,N_4451);
nor U4594 (N_4594,N_4177,N_4133);
and U4595 (N_4595,N_4469,N_4144);
nor U4596 (N_4596,N_4392,N_4329);
nand U4597 (N_4597,N_4203,N_4071);
nor U4598 (N_4598,N_4140,N_4326);
and U4599 (N_4599,N_4096,N_4110);
xor U4600 (N_4600,N_4366,N_4025);
xnor U4601 (N_4601,N_4231,N_4270);
and U4602 (N_4602,N_4069,N_4127);
or U4603 (N_4603,N_4221,N_4365);
nand U4604 (N_4604,N_4483,N_4345);
nor U4605 (N_4605,N_4119,N_4373);
nand U4606 (N_4606,N_4389,N_4450);
nand U4607 (N_4607,N_4255,N_4337);
nor U4608 (N_4608,N_4251,N_4145);
xor U4609 (N_4609,N_4287,N_4143);
nand U4610 (N_4610,N_4227,N_4013);
nor U4611 (N_4611,N_4209,N_4194);
xor U4612 (N_4612,N_4420,N_4018);
nor U4613 (N_4613,N_4053,N_4216);
xor U4614 (N_4614,N_4094,N_4316);
or U4615 (N_4615,N_4352,N_4498);
xor U4616 (N_4616,N_4293,N_4126);
or U4617 (N_4617,N_4019,N_4171);
nand U4618 (N_4618,N_4101,N_4465);
nand U4619 (N_4619,N_4482,N_4467);
or U4620 (N_4620,N_4478,N_4149);
xnor U4621 (N_4621,N_4232,N_4321);
or U4622 (N_4622,N_4083,N_4045);
and U4623 (N_4623,N_4387,N_4246);
nor U4624 (N_4624,N_4357,N_4090);
nand U4625 (N_4625,N_4201,N_4457);
xor U4626 (N_4626,N_4249,N_4055);
or U4627 (N_4627,N_4427,N_4137);
and U4628 (N_4628,N_4213,N_4452);
xnor U4629 (N_4629,N_4205,N_4346);
nand U4630 (N_4630,N_4223,N_4442);
nor U4631 (N_4631,N_4162,N_4409);
or U4632 (N_4632,N_4391,N_4317);
nand U4633 (N_4633,N_4439,N_4164);
and U4634 (N_4634,N_4075,N_4079);
nand U4635 (N_4635,N_4052,N_4494);
or U4636 (N_4636,N_4489,N_4344);
nor U4637 (N_4637,N_4369,N_4297);
and U4638 (N_4638,N_4474,N_4059);
nand U4639 (N_4639,N_4347,N_4159);
xor U4640 (N_4640,N_4394,N_4492);
xor U4641 (N_4641,N_4011,N_4168);
or U4642 (N_4642,N_4146,N_4006);
xnor U4643 (N_4643,N_4064,N_4072);
and U4644 (N_4644,N_4187,N_4134);
nor U4645 (N_4645,N_4463,N_4319);
nor U4646 (N_4646,N_4265,N_4218);
nand U4647 (N_4647,N_4130,N_4037);
or U4648 (N_4648,N_4307,N_4333);
nor U4649 (N_4649,N_4471,N_4275);
or U4650 (N_4650,N_4433,N_4060);
and U4651 (N_4651,N_4091,N_4473);
and U4652 (N_4652,N_4160,N_4178);
nand U4653 (N_4653,N_4012,N_4109);
or U4654 (N_4654,N_4367,N_4002);
nor U4655 (N_4655,N_4301,N_4189);
nor U4656 (N_4656,N_4340,N_4068);
nand U4657 (N_4657,N_4300,N_4000);
and U4658 (N_4658,N_4379,N_4290);
nor U4659 (N_4659,N_4196,N_4258);
xor U4660 (N_4660,N_4410,N_4063);
nor U4661 (N_4661,N_4294,N_4156);
or U4662 (N_4662,N_4497,N_4040);
or U4663 (N_4663,N_4259,N_4462);
nand U4664 (N_4664,N_4009,N_4157);
nor U4665 (N_4665,N_4335,N_4056);
and U4666 (N_4666,N_4257,N_4067);
and U4667 (N_4667,N_4495,N_4100);
nand U4668 (N_4668,N_4044,N_4172);
nand U4669 (N_4669,N_4029,N_4035);
and U4670 (N_4670,N_4039,N_4070);
or U4671 (N_4671,N_4132,N_4192);
nor U4672 (N_4672,N_4499,N_4237);
nor U4673 (N_4673,N_4115,N_4313);
nand U4674 (N_4674,N_4242,N_4112);
nand U4675 (N_4675,N_4479,N_4459);
and U4676 (N_4676,N_4179,N_4176);
xor U4677 (N_4677,N_4141,N_4250);
and U4678 (N_4678,N_4461,N_4308);
or U4679 (N_4679,N_4136,N_4214);
nor U4680 (N_4680,N_4368,N_4267);
nand U4681 (N_4681,N_4153,N_4028);
nor U4682 (N_4682,N_4411,N_4008);
nor U4683 (N_4683,N_4332,N_4336);
xor U4684 (N_4684,N_4066,N_4443);
nand U4685 (N_4685,N_4116,N_4247);
or U4686 (N_4686,N_4299,N_4417);
nor U4687 (N_4687,N_4400,N_4264);
xnor U4688 (N_4688,N_4487,N_4418);
xnor U4689 (N_4689,N_4184,N_4312);
nand U4690 (N_4690,N_4266,N_4078);
nand U4691 (N_4691,N_4173,N_4449);
nand U4692 (N_4692,N_4291,N_4174);
or U4693 (N_4693,N_4122,N_4350);
xnor U4694 (N_4694,N_4404,N_4436);
nand U4695 (N_4695,N_4314,N_4382);
nor U4696 (N_4696,N_4325,N_4296);
nand U4697 (N_4697,N_4380,N_4243);
nand U4698 (N_4698,N_4324,N_4397);
xor U4699 (N_4699,N_4353,N_4191);
xnor U4700 (N_4700,N_4396,N_4161);
nand U4701 (N_4701,N_4118,N_4486);
or U4702 (N_4702,N_4273,N_4204);
nor U4703 (N_4703,N_4289,N_4043);
xor U4704 (N_4704,N_4398,N_4238);
or U4705 (N_4705,N_4355,N_4105);
and U4706 (N_4706,N_4444,N_4413);
xor U4707 (N_4707,N_4371,N_4424);
or U4708 (N_4708,N_4468,N_4284);
or U4709 (N_4709,N_4197,N_4429);
xnor U4710 (N_4710,N_4278,N_4087);
nand U4711 (N_4711,N_4374,N_4032);
and U4712 (N_4712,N_4190,N_4440);
nor U4713 (N_4713,N_4195,N_4062);
nand U4714 (N_4714,N_4129,N_4081);
xnor U4715 (N_4715,N_4236,N_4107);
nand U4716 (N_4716,N_4103,N_4113);
and U4717 (N_4717,N_4193,N_4048);
nand U4718 (N_4718,N_4283,N_4464);
nor U4719 (N_4719,N_4114,N_4098);
nand U4720 (N_4720,N_4277,N_4175);
nor U4721 (N_4721,N_4158,N_4309);
xnor U4722 (N_4722,N_4104,N_4490);
nor U4723 (N_4723,N_4447,N_4304);
nand U4724 (N_4724,N_4466,N_4182);
or U4725 (N_4725,N_4431,N_4302);
or U4726 (N_4726,N_4082,N_4472);
xor U4727 (N_4727,N_4084,N_4282);
nor U4728 (N_4728,N_4219,N_4351);
nor U4729 (N_4729,N_4050,N_4412);
nor U4730 (N_4730,N_4362,N_4054);
nand U4731 (N_4731,N_4239,N_4163);
or U4732 (N_4732,N_4419,N_4432);
nand U4733 (N_4733,N_4121,N_4261);
nor U4734 (N_4734,N_4306,N_4271);
or U4735 (N_4735,N_4226,N_4021);
nand U4736 (N_4736,N_4015,N_4088);
nor U4737 (N_4737,N_4016,N_4027);
nor U4738 (N_4738,N_4285,N_4222);
nand U4739 (N_4739,N_4481,N_4354);
nor U4740 (N_4740,N_4315,N_4455);
xnor U4741 (N_4741,N_4263,N_4212);
and U4742 (N_4742,N_4358,N_4181);
xor U4743 (N_4743,N_4183,N_4386);
or U4744 (N_4744,N_4051,N_4363);
nor U4745 (N_4745,N_4135,N_4286);
xnor U4746 (N_4746,N_4438,N_4493);
nor U4747 (N_4747,N_4004,N_4170);
and U4748 (N_4748,N_4041,N_4036);
or U4749 (N_4749,N_4378,N_4128);
nand U4750 (N_4750,N_4049,N_4320);
and U4751 (N_4751,N_4088,N_4345);
and U4752 (N_4752,N_4385,N_4004);
nor U4753 (N_4753,N_4429,N_4098);
xor U4754 (N_4754,N_4021,N_4288);
or U4755 (N_4755,N_4387,N_4074);
nand U4756 (N_4756,N_4210,N_4316);
and U4757 (N_4757,N_4181,N_4495);
and U4758 (N_4758,N_4497,N_4403);
nor U4759 (N_4759,N_4261,N_4101);
and U4760 (N_4760,N_4273,N_4143);
or U4761 (N_4761,N_4486,N_4117);
nand U4762 (N_4762,N_4187,N_4254);
nand U4763 (N_4763,N_4491,N_4290);
xnor U4764 (N_4764,N_4146,N_4136);
nand U4765 (N_4765,N_4070,N_4103);
nor U4766 (N_4766,N_4419,N_4316);
nand U4767 (N_4767,N_4000,N_4293);
and U4768 (N_4768,N_4356,N_4407);
nor U4769 (N_4769,N_4435,N_4021);
or U4770 (N_4770,N_4276,N_4418);
nor U4771 (N_4771,N_4022,N_4432);
nand U4772 (N_4772,N_4066,N_4440);
xnor U4773 (N_4773,N_4096,N_4135);
nand U4774 (N_4774,N_4012,N_4085);
or U4775 (N_4775,N_4440,N_4254);
or U4776 (N_4776,N_4089,N_4011);
xor U4777 (N_4777,N_4081,N_4464);
and U4778 (N_4778,N_4147,N_4366);
and U4779 (N_4779,N_4003,N_4300);
nand U4780 (N_4780,N_4427,N_4416);
nor U4781 (N_4781,N_4169,N_4078);
or U4782 (N_4782,N_4380,N_4144);
nor U4783 (N_4783,N_4163,N_4160);
or U4784 (N_4784,N_4434,N_4158);
nor U4785 (N_4785,N_4316,N_4391);
nor U4786 (N_4786,N_4477,N_4107);
or U4787 (N_4787,N_4014,N_4097);
and U4788 (N_4788,N_4162,N_4015);
or U4789 (N_4789,N_4412,N_4280);
nand U4790 (N_4790,N_4297,N_4403);
nor U4791 (N_4791,N_4479,N_4357);
or U4792 (N_4792,N_4268,N_4208);
or U4793 (N_4793,N_4168,N_4093);
nor U4794 (N_4794,N_4126,N_4038);
nand U4795 (N_4795,N_4024,N_4293);
nor U4796 (N_4796,N_4465,N_4099);
xor U4797 (N_4797,N_4493,N_4463);
nor U4798 (N_4798,N_4285,N_4104);
xor U4799 (N_4799,N_4012,N_4411);
nand U4800 (N_4800,N_4104,N_4033);
or U4801 (N_4801,N_4156,N_4075);
nor U4802 (N_4802,N_4367,N_4220);
and U4803 (N_4803,N_4390,N_4246);
and U4804 (N_4804,N_4017,N_4202);
or U4805 (N_4805,N_4108,N_4474);
nand U4806 (N_4806,N_4344,N_4400);
and U4807 (N_4807,N_4228,N_4314);
nor U4808 (N_4808,N_4192,N_4129);
nand U4809 (N_4809,N_4483,N_4365);
and U4810 (N_4810,N_4158,N_4297);
or U4811 (N_4811,N_4003,N_4466);
nand U4812 (N_4812,N_4031,N_4455);
xnor U4813 (N_4813,N_4183,N_4421);
nor U4814 (N_4814,N_4254,N_4259);
nand U4815 (N_4815,N_4375,N_4027);
or U4816 (N_4816,N_4476,N_4354);
and U4817 (N_4817,N_4109,N_4341);
nand U4818 (N_4818,N_4197,N_4066);
nand U4819 (N_4819,N_4435,N_4464);
xor U4820 (N_4820,N_4277,N_4129);
or U4821 (N_4821,N_4231,N_4360);
xor U4822 (N_4822,N_4403,N_4292);
or U4823 (N_4823,N_4432,N_4010);
or U4824 (N_4824,N_4458,N_4038);
or U4825 (N_4825,N_4055,N_4026);
nand U4826 (N_4826,N_4143,N_4189);
xnor U4827 (N_4827,N_4446,N_4136);
and U4828 (N_4828,N_4320,N_4056);
nand U4829 (N_4829,N_4326,N_4170);
and U4830 (N_4830,N_4125,N_4056);
nor U4831 (N_4831,N_4177,N_4490);
nand U4832 (N_4832,N_4270,N_4073);
xor U4833 (N_4833,N_4337,N_4028);
nor U4834 (N_4834,N_4128,N_4448);
or U4835 (N_4835,N_4255,N_4447);
and U4836 (N_4836,N_4243,N_4441);
xor U4837 (N_4837,N_4145,N_4490);
or U4838 (N_4838,N_4212,N_4178);
and U4839 (N_4839,N_4375,N_4133);
or U4840 (N_4840,N_4155,N_4050);
nor U4841 (N_4841,N_4440,N_4358);
xnor U4842 (N_4842,N_4170,N_4123);
and U4843 (N_4843,N_4268,N_4141);
nor U4844 (N_4844,N_4237,N_4178);
nor U4845 (N_4845,N_4094,N_4351);
and U4846 (N_4846,N_4326,N_4304);
or U4847 (N_4847,N_4275,N_4297);
xor U4848 (N_4848,N_4394,N_4289);
nand U4849 (N_4849,N_4481,N_4170);
nor U4850 (N_4850,N_4119,N_4382);
or U4851 (N_4851,N_4035,N_4243);
nor U4852 (N_4852,N_4144,N_4065);
xor U4853 (N_4853,N_4024,N_4079);
and U4854 (N_4854,N_4288,N_4472);
nand U4855 (N_4855,N_4274,N_4172);
and U4856 (N_4856,N_4133,N_4157);
xor U4857 (N_4857,N_4190,N_4362);
nand U4858 (N_4858,N_4051,N_4095);
nand U4859 (N_4859,N_4022,N_4050);
and U4860 (N_4860,N_4040,N_4159);
nand U4861 (N_4861,N_4205,N_4176);
nor U4862 (N_4862,N_4313,N_4482);
nor U4863 (N_4863,N_4268,N_4043);
xnor U4864 (N_4864,N_4225,N_4369);
xnor U4865 (N_4865,N_4230,N_4455);
nor U4866 (N_4866,N_4406,N_4311);
nor U4867 (N_4867,N_4470,N_4257);
or U4868 (N_4868,N_4127,N_4493);
nor U4869 (N_4869,N_4237,N_4167);
xor U4870 (N_4870,N_4176,N_4168);
and U4871 (N_4871,N_4024,N_4321);
and U4872 (N_4872,N_4359,N_4264);
nand U4873 (N_4873,N_4181,N_4458);
or U4874 (N_4874,N_4024,N_4330);
nand U4875 (N_4875,N_4182,N_4400);
xnor U4876 (N_4876,N_4177,N_4314);
or U4877 (N_4877,N_4463,N_4498);
xnor U4878 (N_4878,N_4498,N_4401);
and U4879 (N_4879,N_4138,N_4395);
and U4880 (N_4880,N_4431,N_4009);
nor U4881 (N_4881,N_4008,N_4152);
nor U4882 (N_4882,N_4402,N_4371);
or U4883 (N_4883,N_4307,N_4121);
nand U4884 (N_4884,N_4272,N_4189);
and U4885 (N_4885,N_4322,N_4072);
xor U4886 (N_4886,N_4079,N_4342);
nor U4887 (N_4887,N_4421,N_4093);
nor U4888 (N_4888,N_4345,N_4105);
nand U4889 (N_4889,N_4101,N_4278);
and U4890 (N_4890,N_4064,N_4160);
and U4891 (N_4891,N_4014,N_4033);
xnor U4892 (N_4892,N_4308,N_4313);
xor U4893 (N_4893,N_4488,N_4024);
nand U4894 (N_4894,N_4366,N_4243);
xnor U4895 (N_4895,N_4248,N_4139);
and U4896 (N_4896,N_4309,N_4455);
nor U4897 (N_4897,N_4290,N_4303);
and U4898 (N_4898,N_4224,N_4047);
nor U4899 (N_4899,N_4344,N_4330);
nand U4900 (N_4900,N_4280,N_4359);
nand U4901 (N_4901,N_4297,N_4436);
xor U4902 (N_4902,N_4254,N_4231);
or U4903 (N_4903,N_4196,N_4127);
nand U4904 (N_4904,N_4325,N_4335);
or U4905 (N_4905,N_4425,N_4449);
xor U4906 (N_4906,N_4268,N_4228);
nand U4907 (N_4907,N_4266,N_4100);
or U4908 (N_4908,N_4368,N_4040);
xnor U4909 (N_4909,N_4384,N_4340);
nand U4910 (N_4910,N_4487,N_4244);
xor U4911 (N_4911,N_4287,N_4020);
or U4912 (N_4912,N_4212,N_4326);
xor U4913 (N_4913,N_4056,N_4483);
xnor U4914 (N_4914,N_4019,N_4160);
nand U4915 (N_4915,N_4189,N_4393);
nand U4916 (N_4916,N_4162,N_4101);
xor U4917 (N_4917,N_4325,N_4456);
nor U4918 (N_4918,N_4252,N_4035);
and U4919 (N_4919,N_4189,N_4116);
xnor U4920 (N_4920,N_4301,N_4383);
nand U4921 (N_4921,N_4468,N_4362);
nand U4922 (N_4922,N_4499,N_4043);
xnor U4923 (N_4923,N_4354,N_4406);
nand U4924 (N_4924,N_4444,N_4279);
nor U4925 (N_4925,N_4421,N_4439);
xnor U4926 (N_4926,N_4241,N_4180);
xor U4927 (N_4927,N_4165,N_4003);
or U4928 (N_4928,N_4113,N_4329);
nand U4929 (N_4929,N_4153,N_4295);
or U4930 (N_4930,N_4251,N_4204);
xor U4931 (N_4931,N_4183,N_4126);
and U4932 (N_4932,N_4404,N_4431);
nor U4933 (N_4933,N_4422,N_4478);
nor U4934 (N_4934,N_4287,N_4345);
nand U4935 (N_4935,N_4008,N_4108);
and U4936 (N_4936,N_4457,N_4405);
xnor U4937 (N_4937,N_4489,N_4114);
xnor U4938 (N_4938,N_4221,N_4177);
and U4939 (N_4939,N_4484,N_4280);
and U4940 (N_4940,N_4483,N_4112);
and U4941 (N_4941,N_4320,N_4417);
xor U4942 (N_4942,N_4385,N_4386);
nor U4943 (N_4943,N_4107,N_4394);
and U4944 (N_4944,N_4132,N_4295);
nand U4945 (N_4945,N_4398,N_4104);
nand U4946 (N_4946,N_4391,N_4164);
xnor U4947 (N_4947,N_4117,N_4289);
or U4948 (N_4948,N_4155,N_4044);
or U4949 (N_4949,N_4299,N_4221);
nor U4950 (N_4950,N_4367,N_4357);
xnor U4951 (N_4951,N_4005,N_4257);
and U4952 (N_4952,N_4097,N_4171);
nor U4953 (N_4953,N_4443,N_4401);
nand U4954 (N_4954,N_4056,N_4102);
nor U4955 (N_4955,N_4241,N_4324);
and U4956 (N_4956,N_4014,N_4385);
nor U4957 (N_4957,N_4495,N_4202);
or U4958 (N_4958,N_4193,N_4403);
or U4959 (N_4959,N_4283,N_4149);
and U4960 (N_4960,N_4071,N_4476);
nand U4961 (N_4961,N_4077,N_4242);
xnor U4962 (N_4962,N_4373,N_4440);
xor U4963 (N_4963,N_4303,N_4095);
nor U4964 (N_4964,N_4310,N_4273);
xnor U4965 (N_4965,N_4212,N_4334);
or U4966 (N_4966,N_4044,N_4140);
nor U4967 (N_4967,N_4099,N_4300);
nand U4968 (N_4968,N_4034,N_4054);
or U4969 (N_4969,N_4173,N_4055);
xnor U4970 (N_4970,N_4019,N_4331);
xor U4971 (N_4971,N_4179,N_4347);
nor U4972 (N_4972,N_4379,N_4496);
and U4973 (N_4973,N_4391,N_4023);
and U4974 (N_4974,N_4498,N_4106);
nor U4975 (N_4975,N_4310,N_4041);
nor U4976 (N_4976,N_4087,N_4162);
and U4977 (N_4977,N_4022,N_4141);
xor U4978 (N_4978,N_4408,N_4280);
and U4979 (N_4979,N_4472,N_4395);
nand U4980 (N_4980,N_4023,N_4361);
nor U4981 (N_4981,N_4168,N_4212);
or U4982 (N_4982,N_4370,N_4075);
or U4983 (N_4983,N_4298,N_4442);
or U4984 (N_4984,N_4071,N_4187);
nand U4985 (N_4985,N_4351,N_4053);
nor U4986 (N_4986,N_4369,N_4149);
and U4987 (N_4987,N_4131,N_4367);
nand U4988 (N_4988,N_4044,N_4100);
nor U4989 (N_4989,N_4064,N_4281);
xor U4990 (N_4990,N_4117,N_4357);
nand U4991 (N_4991,N_4409,N_4385);
or U4992 (N_4992,N_4366,N_4080);
nand U4993 (N_4993,N_4014,N_4222);
or U4994 (N_4994,N_4288,N_4010);
or U4995 (N_4995,N_4462,N_4129);
and U4996 (N_4996,N_4337,N_4473);
xor U4997 (N_4997,N_4256,N_4438);
or U4998 (N_4998,N_4290,N_4232);
nand U4999 (N_4999,N_4265,N_4081);
xor U5000 (N_5000,N_4587,N_4844);
and U5001 (N_5001,N_4725,N_4934);
nand U5002 (N_5002,N_4797,N_4639);
and U5003 (N_5003,N_4562,N_4822);
or U5004 (N_5004,N_4666,N_4632);
or U5005 (N_5005,N_4712,N_4554);
or U5006 (N_5006,N_4594,N_4978);
and U5007 (N_5007,N_4746,N_4915);
and U5008 (N_5008,N_4843,N_4876);
nand U5009 (N_5009,N_4741,N_4714);
or U5010 (N_5010,N_4709,N_4858);
nand U5011 (N_5011,N_4667,N_4793);
nand U5012 (N_5012,N_4513,N_4648);
and U5013 (N_5013,N_4547,N_4987);
or U5014 (N_5014,N_4592,N_4745);
nor U5015 (N_5015,N_4734,N_4806);
xor U5016 (N_5016,N_4574,N_4864);
nand U5017 (N_5017,N_4724,N_4925);
or U5018 (N_5018,N_4726,N_4600);
nor U5019 (N_5019,N_4583,N_4560);
nand U5020 (N_5020,N_4754,N_4750);
xnor U5021 (N_5021,N_4658,N_4768);
xnor U5022 (N_5022,N_4718,N_4581);
nand U5023 (N_5023,N_4846,N_4707);
or U5024 (N_5024,N_4875,N_4857);
xnor U5025 (N_5025,N_4696,N_4553);
nand U5026 (N_5026,N_4802,N_4789);
nand U5027 (N_5027,N_4898,N_4663);
nor U5028 (N_5028,N_4653,N_4737);
and U5029 (N_5029,N_4956,N_4928);
nor U5030 (N_5030,N_4706,N_4609);
nor U5031 (N_5031,N_4952,N_4633);
or U5032 (N_5032,N_4816,N_4539);
and U5033 (N_5033,N_4540,N_4739);
nor U5034 (N_5034,N_4983,N_4975);
and U5035 (N_5035,N_4618,N_4660);
or U5036 (N_5036,N_4919,N_4577);
xnor U5037 (N_5037,N_4603,N_4941);
nor U5038 (N_5038,N_4635,N_4736);
and U5039 (N_5039,N_4519,N_4527);
nor U5040 (N_5040,N_4572,N_4917);
or U5041 (N_5041,N_4582,N_4868);
nor U5042 (N_5042,N_4533,N_4828);
and U5043 (N_5043,N_4637,N_4644);
nand U5044 (N_5044,N_4955,N_4926);
nor U5045 (N_5045,N_4505,N_4848);
and U5046 (N_5046,N_4508,N_4701);
or U5047 (N_5047,N_4555,N_4931);
and U5048 (N_5048,N_4524,N_4728);
nor U5049 (N_5049,N_4812,N_4591);
or U5050 (N_5050,N_4971,N_4944);
xnor U5051 (N_5051,N_4954,N_4872);
nand U5052 (N_5052,N_4589,N_4881);
xor U5053 (N_5053,N_4845,N_4780);
or U5054 (N_5054,N_4831,N_4570);
nand U5055 (N_5055,N_4690,N_4897);
nor U5056 (N_5056,N_4715,N_4579);
and U5057 (N_5057,N_4762,N_4966);
xnor U5058 (N_5058,N_4650,N_4847);
nor U5059 (N_5059,N_4672,N_4853);
and U5060 (N_5060,N_4604,N_4902);
xnor U5061 (N_5061,N_4886,N_4622);
xnor U5062 (N_5062,N_4567,N_4814);
and U5063 (N_5063,N_4766,N_4520);
or U5064 (N_5064,N_4504,N_4751);
and U5065 (N_5065,N_4948,N_4962);
or U5066 (N_5066,N_4891,N_4534);
nor U5067 (N_5067,N_4601,N_4636);
nand U5068 (N_5068,N_4733,N_4871);
nor U5069 (N_5069,N_4748,N_4883);
and U5070 (N_5070,N_4985,N_4757);
xnor U5071 (N_5071,N_4970,N_4564);
and U5072 (N_5072,N_4783,N_4835);
and U5073 (N_5073,N_4628,N_4861);
nand U5074 (N_5074,N_4964,N_4984);
or U5075 (N_5075,N_4957,N_4959);
nand U5076 (N_5076,N_4924,N_4998);
xnor U5077 (N_5077,N_4829,N_4680);
nand U5078 (N_5078,N_4824,N_4683);
xor U5079 (N_5079,N_4758,N_4731);
xor U5080 (N_5080,N_4986,N_4598);
nor U5081 (N_5081,N_4640,N_4590);
xor U5082 (N_5082,N_4907,N_4646);
nand U5083 (N_5083,N_4870,N_4665);
and U5084 (N_5084,N_4961,N_4935);
xor U5085 (N_5085,N_4550,N_4638);
or U5086 (N_5086,N_4990,N_4662);
and U5087 (N_5087,N_4760,N_4947);
nand U5088 (N_5088,N_4951,N_4630);
xor U5089 (N_5089,N_4918,N_4624);
xor U5090 (N_5090,N_4677,N_4652);
nor U5091 (N_5091,N_4526,N_4634);
nand U5092 (N_5092,N_4867,N_4874);
xor U5093 (N_5093,N_4992,N_4509);
or U5094 (N_5094,N_4813,N_4626);
nand U5095 (N_5095,N_4788,N_4958);
nor U5096 (N_5096,N_4989,N_4997);
or U5097 (N_5097,N_4791,N_4865);
and U5098 (N_5098,N_4890,N_4573);
nor U5099 (N_5099,N_4825,N_4960);
and U5100 (N_5100,N_4596,N_4777);
nor U5101 (N_5101,N_4950,N_4586);
or U5102 (N_5102,N_4521,N_4700);
nor U5103 (N_5103,N_4972,N_4805);
nor U5104 (N_5104,N_4559,N_4678);
nor U5105 (N_5105,N_4675,N_4682);
nor U5106 (N_5106,N_4608,N_4568);
xnor U5107 (N_5107,N_4514,N_4536);
nor U5108 (N_5108,N_4765,N_4548);
nand U5109 (N_5109,N_4885,N_4647);
and U5110 (N_5110,N_4896,N_4982);
or U5111 (N_5111,N_4738,N_4676);
and U5112 (N_5112,N_4691,N_4545);
xor U5113 (N_5113,N_4641,N_4838);
and U5114 (N_5114,N_4617,N_4742);
or U5115 (N_5115,N_4999,N_4673);
nand U5116 (N_5116,N_4702,N_4878);
nor U5117 (N_5117,N_4921,N_4827);
nor U5118 (N_5118,N_4588,N_4723);
nor U5119 (N_5119,N_4749,N_4819);
nor U5120 (N_5120,N_4859,N_4879);
nor U5121 (N_5121,N_4784,N_4786);
nand U5122 (N_5122,N_4535,N_4727);
or U5123 (N_5123,N_4730,N_4551);
xor U5124 (N_5124,N_4599,N_4882);
xor U5125 (N_5125,N_4597,N_4889);
xor U5126 (N_5126,N_4770,N_4798);
xnor U5127 (N_5127,N_4967,N_4576);
xnor U5128 (N_5128,N_4595,N_4888);
nor U5129 (N_5129,N_4654,N_4538);
and U5130 (N_5130,N_4721,N_4785);
nor U5131 (N_5131,N_4979,N_4656);
nor U5132 (N_5132,N_4507,N_4942);
nand U5133 (N_5133,N_4720,N_4580);
and U5134 (N_5134,N_4991,N_4887);
or U5135 (N_5135,N_4914,N_4856);
nor U5136 (N_5136,N_4541,N_4556);
nor U5137 (N_5137,N_4929,N_4779);
nor U5138 (N_5138,N_4500,N_4674);
nand U5139 (N_5139,N_4523,N_4661);
nand U5140 (N_5140,N_4605,N_4968);
xor U5141 (N_5141,N_4900,N_4906);
nor U5142 (N_5142,N_4818,N_4965);
nor U5143 (N_5143,N_4512,N_4552);
xnor U5144 (N_5144,N_4933,N_4826);
nor U5145 (N_5145,N_4710,N_4804);
and U5146 (N_5146,N_4855,N_4893);
and U5147 (N_5147,N_4688,N_4940);
nor U5148 (N_5148,N_4877,N_4518);
nor U5149 (N_5149,N_4761,N_4558);
nand U5150 (N_5150,N_4894,N_4773);
nor U5151 (N_5151,N_4963,N_4629);
and U5152 (N_5152,N_4860,N_4543);
and U5153 (N_5153,N_4530,N_4616);
nor U5154 (N_5154,N_4930,N_4911);
xor U5155 (N_5155,N_4842,N_4722);
or U5156 (N_5156,N_4615,N_4685);
and U5157 (N_5157,N_4912,N_4664);
xor U5158 (N_5158,N_4800,N_4927);
nor U5159 (N_5159,N_4585,N_4790);
nor U5160 (N_5160,N_4695,N_4895);
and U5161 (N_5161,N_4620,N_4980);
xor U5162 (N_5162,N_4981,N_4953);
or U5163 (N_5163,N_4692,N_4566);
or U5164 (N_5164,N_4515,N_4631);
nand U5165 (N_5165,N_4913,N_4973);
nor U5166 (N_5166,N_4901,N_4516);
or U5167 (N_5167,N_4936,N_4621);
xor U5168 (N_5168,N_4905,N_4899);
and U5169 (N_5169,N_4625,N_4923);
nor U5170 (N_5170,N_4995,N_4694);
and U5171 (N_5171,N_4510,N_4686);
and U5172 (N_5172,N_4670,N_4781);
or U5173 (N_5173,N_4852,N_4502);
nor U5174 (N_5174,N_4866,N_4612);
nand U5175 (N_5175,N_4776,N_4840);
xor U5176 (N_5176,N_4854,N_4892);
or U5177 (N_5177,N_4943,N_4668);
or U5178 (N_5178,N_4528,N_4795);
xor U5179 (N_5179,N_4969,N_4809);
nor U5180 (N_5180,N_4529,N_4546);
and U5181 (N_5181,N_4732,N_4703);
or U5182 (N_5182,N_4873,N_4904);
nor U5183 (N_5183,N_4503,N_4849);
nand U5184 (N_5184,N_4837,N_4763);
nand U5185 (N_5185,N_4974,N_4922);
or U5186 (N_5186,N_4833,N_4920);
and U5187 (N_5187,N_4544,N_4775);
nand U5188 (N_5188,N_4810,N_4705);
nor U5189 (N_5189,N_4764,N_4735);
xor U5190 (N_5190,N_4561,N_4988);
or U5191 (N_5191,N_4778,N_4704);
and U5192 (N_5192,N_4657,N_4708);
or U5193 (N_5193,N_4651,N_4711);
nand U5194 (N_5194,N_4501,N_4697);
or U5195 (N_5195,N_4817,N_4549);
and U5196 (N_5196,N_4698,N_4994);
nand U5197 (N_5197,N_4611,N_4755);
nor U5198 (N_5198,N_4531,N_4681);
and U5199 (N_5199,N_4659,N_4832);
xnor U5200 (N_5200,N_4836,N_4569);
or U5201 (N_5201,N_4578,N_4839);
and U5202 (N_5202,N_4506,N_4627);
nor U5203 (N_5203,N_4740,N_4932);
and U5204 (N_5204,N_4643,N_4850);
and U5205 (N_5205,N_4851,N_4719);
nand U5206 (N_5206,N_4799,N_4769);
nand U5207 (N_5207,N_4649,N_4908);
or U5208 (N_5208,N_4747,N_4614);
and U5209 (N_5209,N_4880,N_4939);
and U5210 (N_5210,N_4687,N_4977);
nand U5211 (N_5211,N_4794,N_4787);
or U5212 (N_5212,N_4532,N_4863);
and U5213 (N_5213,N_4811,N_4606);
or U5214 (N_5214,N_4807,N_4689);
or U5215 (N_5215,N_4642,N_4772);
nor U5216 (N_5216,N_4949,N_4623);
nor U5217 (N_5217,N_4542,N_4909);
or U5218 (N_5218,N_4537,N_4684);
nand U5219 (N_5219,N_4938,N_4815);
nor U5220 (N_5220,N_4993,N_4593);
xnor U5221 (N_5221,N_4602,N_4699);
xor U5222 (N_5222,N_4525,N_4743);
or U5223 (N_5223,N_4752,N_4759);
or U5224 (N_5224,N_4910,N_4821);
and U5225 (N_5225,N_4571,N_4796);
xor U5226 (N_5226,N_4830,N_4803);
xor U5227 (N_5227,N_4729,N_4884);
nand U5228 (N_5228,N_4565,N_4903);
xnor U5229 (N_5229,N_4679,N_4841);
xnor U5230 (N_5230,N_4820,N_4575);
and U5231 (N_5231,N_4834,N_4713);
and U5232 (N_5232,N_4945,N_4693);
nor U5233 (N_5233,N_4607,N_4767);
and U5234 (N_5234,N_4613,N_4916);
nor U5235 (N_5235,N_4753,N_4996);
xnor U5236 (N_5236,N_4645,N_4584);
and U5237 (N_5237,N_4869,N_4717);
or U5238 (N_5238,N_4522,N_4610);
and U5239 (N_5239,N_4716,N_4774);
nand U5240 (N_5240,N_4976,N_4801);
nand U5241 (N_5241,N_4655,N_4671);
nand U5242 (N_5242,N_4937,N_4771);
or U5243 (N_5243,N_4619,N_4563);
nand U5244 (N_5244,N_4782,N_4511);
nand U5245 (N_5245,N_4557,N_4946);
or U5246 (N_5246,N_4744,N_4808);
or U5247 (N_5247,N_4862,N_4517);
nand U5248 (N_5248,N_4669,N_4823);
and U5249 (N_5249,N_4792,N_4756);
or U5250 (N_5250,N_4768,N_4843);
nor U5251 (N_5251,N_4608,N_4762);
or U5252 (N_5252,N_4988,N_4582);
nor U5253 (N_5253,N_4662,N_4707);
nand U5254 (N_5254,N_4937,N_4521);
or U5255 (N_5255,N_4815,N_4893);
xor U5256 (N_5256,N_4814,N_4556);
nor U5257 (N_5257,N_4811,N_4845);
nand U5258 (N_5258,N_4647,N_4822);
nand U5259 (N_5259,N_4510,N_4772);
or U5260 (N_5260,N_4907,N_4892);
and U5261 (N_5261,N_4615,N_4759);
and U5262 (N_5262,N_4852,N_4980);
or U5263 (N_5263,N_4854,N_4708);
nand U5264 (N_5264,N_4941,N_4541);
or U5265 (N_5265,N_4618,N_4826);
nand U5266 (N_5266,N_4898,N_4983);
and U5267 (N_5267,N_4661,N_4814);
and U5268 (N_5268,N_4543,N_4873);
nand U5269 (N_5269,N_4510,N_4623);
xor U5270 (N_5270,N_4915,N_4654);
or U5271 (N_5271,N_4885,N_4672);
or U5272 (N_5272,N_4977,N_4785);
or U5273 (N_5273,N_4678,N_4978);
and U5274 (N_5274,N_4587,N_4935);
or U5275 (N_5275,N_4592,N_4762);
nor U5276 (N_5276,N_4507,N_4933);
and U5277 (N_5277,N_4811,N_4841);
nand U5278 (N_5278,N_4736,N_4672);
xor U5279 (N_5279,N_4839,N_4670);
and U5280 (N_5280,N_4749,N_4908);
nor U5281 (N_5281,N_4515,N_4809);
nor U5282 (N_5282,N_4536,N_4703);
nand U5283 (N_5283,N_4879,N_4690);
xnor U5284 (N_5284,N_4584,N_4512);
nor U5285 (N_5285,N_4658,N_4851);
or U5286 (N_5286,N_4808,N_4802);
or U5287 (N_5287,N_4776,N_4580);
nand U5288 (N_5288,N_4925,N_4761);
nor U5289 (N_5289,N_4668,N_4639);
nor U5290 (N_5290,N_4842,N_4633);
and U5291 (N_5291,N_4810,N_4597);
nor U5292 (N_5292,N_4756,N_4589);
and U5293 (N_5293,N_4523,N_4706);
nor U5294 (N_5294,N_4979,N_4755);
or U5295 (N_5295,N_4606,N_4738);
nor U5296 (N_5296,N_4952,N_4558);
or U5297 (N_5297,N_4926,N_4671);
or U5298 (N_5298,N_4812,N_4519);
xor U5299 (N_5299,N_4724,N_4670);
nor U5300 (N_5300,N_4758,N_4950);
nand U5301 (N_5301,N_4727,N_4663);
or U5302 (N_5302,N_4928,N_4595);
or U5303 (N_5303,N_4785,N_4729);
and U5304 (N_5304,N_4562,N_4710);
and U5305 (N_5305,N_4519,N_4952);
or U5306 (N_5306,N_4534,N_4763);
or U5307 (N_5307,N_4648,N_4552);
and U5308 (N_5308,N_4673,N_4957);
nor U5309 (N_5309,N_4660,N_4815);
or U5310 (N_5310,N_4643,N_4546);
and U5311 (N_5311,N_4848,N_4644);
or U5312 (N_5312,N_4955,N_4709);
nand U5313 (N_5313,N_4789,N_4673);
nand U5314 (N_5314,N_4524,N_4840);
nor U5315 (N_5315,N_4598,N_4787);
or U5316 (N_5316,N_4990,N_4559);
or U5317 (N_5317,N_4938,N_4967);
nand U5318 (N_5318,N_4988,N_4563);
and U5319 (N_5319,N_4734,N_4886);
nor U5320 (N_5320,N_4651,N_4891);
and U5321 (N_5321,N_4517,N_4547);
nor U5322 (N_5322,N_4877,N_4935);
or U5323 (N_5323,N_4638,N_4791);
xnor U5324 (N_5324,N_4809,N_4954);
or U5325 (N_5325,N_4526,N_4789);
nor U5326 (N_5326,N_4906,N_4544);
nor U5327 (N_5327,N_4811,N_4626);
and U5328 (N_5328,N_4794,N_4546);
nor U5329 (N_5329,N_4573,N_4589);
nor U5330 (N_5330,N_4673,N_4943);
xor U5331 (N_5331,N_4591,N_4733);
and U5332 (N_5332,N_4638,N_4621);
nand U5333 (N_5333,N_4590,N_4964);
and U5334 (N_5334,N_4615,N_4870);
nand U5335 (N_5335,N_4596,N_4690);
or U5336 (N_5336,N_4992,N_4986);
or U5337 (N_5337,N_4586,N_4799);
xnor U5338 (N_5338,N_4956,N_4856);
nor U5339 (N_5339,N_4630,N_4793);
nor U5340 (N_5340,N_4799,N_4740);
or U5341 (N_5341,N_4501,N_4762);
xor U5342 (N_5342,N_4959,N_4999);
nor U5343 (N_5343,N_4765,N_4859);
nand U5344 (N_5344,N_4749,N_4688);
nand U5345 (N_5345,N_4665,N_4954);
and U5346 (N_5346,N_4613,N_4920);
or U5347 (N_5347,N_4611,N_4880);
xor U5348 (N_5348,N_4725,N_4714);
xnor U5349 (N_5349,N_4993,N_4634);
xor U5350 (N_5350,N_4865,N_4523);
nor U5351 (N_5351,N_4772,N_4764);
xor U5352 (N_5352,N_4807,N_4821);
nand U5353 (N_5353,N_4580,N_4746);
and U5354 (N_5354,N_4919,N_4548);
nor U5355 (N_5355,N_4968,N_4671);
xnor U5356 (N_5356,N_4661,N_4734);
or U5357 (N_5357,N_4521,N_4918);
and U5358 (N_5358,N_4787,N_4718);
or U5359 (N_5359,N_4787,N_4944);
and U5360 (N_5360,N_4529,N_4598);
or U5361 (N_5361,N_4813,N_4572);
nand U5362 (N_5362,N_4786,N_4796);
and U5363 (N_5363,N_4648,N_4651);
xor U5364 (N_5364,N_4556,N_4900);
xnor U5365 (N_5365,N_4928,N_4977);
and U5366 (N_5366,N_4580,N_4716);
or U5367 (N_5367,N_4763,N_4933);
or U5368 (N_5368,N_4804,N_4540);
or U5369 (N_5369,N_4815,N_4879);
or U5370 (N_5370,N_4832,N_4959);
or U5371 (N_5371,N_4699,N_4595);
or U5372 (N_5372,N_4509,N_4829);
nor U5373 (N_5373,N_4549,N_4667);
xnor U5374 (N_5374,N_4821,N_4757);
nand U5375 (N_5375,N_4514,N_4728);
and U5376 (N_5376,N_4936,N_4534);
nor U5377 (N_5377,N_4650,N_4569);
xor U5378 (N_5378,N_4993,N_4850);
nor U5379 (N_5379,N_4952,N_4879);
xnor U5380 (N_5380,N_4704,N_4910);
and U5381 (N_5381,N_4532,N_4633);
xor U5382 (N_5382,N_4663,N_4592);
or U5383 (N_5383,N_4609,N_4551);
xor U5384 (N_5384,N_4695,N_4857);
nand U5385 (N_5385,N_4712,N_4822);
or U5386 (N_5386,N_4714,N_4929);
xnor U5387 (N_5387,N_4598,N_4608);
xnor U5388 (N_5388,N_4837,N_4988);
nand U5389 (N_5389,N_4574,N_4677);
nor U5390 (N_5390,N_4588,N_4706);
and U5391 (N_5391,N_4714,N_4648);
or U5392 (N_5392,N_4692,N_4859);
or U5393 (N_5393,N_4585,N_4827);
and U5394 (N_5394,N_4831,N_4997);
or U5395 (N_5395,N_4572,N_4962);
nand U5396 (N_5396,N_4897,N_4765);
nand U5397 (N_5397,N_4885,N_4734);
nand U5398 (N_5398,N_4644,N_4757);
nor U5399 (N_5399,N_4959,N_4753);
nand U5400 (N_5400,N_4978,N_4896);
nand U5401 (N_5401,N_4563,N_4906);
nand U5402 (N_5402,N_4802,N_4525);
or U5403 (N_5403,N_4632,N_4647);
nand U5404 (N_5404,N_4863,N_4614);
or U5405 (N_5405,N_4684,N_4768);
or U5406 (N_5406,N_4737,N_4823);
or U5407 (N_5407,N_4716,N_4675);
nor U5408 (N_5408,N_4981,N_4906);
nand U5409 (N_5409,N_4747,N_4709);
xnor U5410 (N_5410,N_4821,N_4615);
xnor U5411 (N_5411,N_4737,N_4966);
and U5412 (N_5412,N_4797,N_4757);
xor U5413 (N_5413,N_4996,N_4615);
xnor U5414 (N_5414,N_4691,N_4987);
nand U5415 (N_5415,N_4536,N_4753);
nand U5416 (N_5416,N_4972,N_4721);
and U5417 (N_5417,N_4762,N_4796);
nand U5418 (N_5418,N_4917,N_4819);
and U5419 (N_5419,N_4552,N_4905);
xnor U5420 (N_5420,N_4863,N_4877);
nand U5421 (N_5421,N_4723,N_4843);
nand U5422 (N_5422,N_4863,N_4779);
xor U5423 (N_5423,N_4847,N_4524);
and U5424 (N_5424,N_4630,N_4925);
and U5425 (N_5425,N_4820,N_4577);
nor U5426 (N_5426,N_4819,N_4671);
or U5427 (N_5427,N_4581,N_4855);
nor U5428 (N_5428,N_4660,N_4859);
nand U5429 (N_5429,N_4989,N_4719);
nand U5430 (N_5430,N_4544,N_4630);
or U5431 (N_5431,N_4637,N_4711);
xor U5432 (N_5432,N_4705,N_4545);
xor U5433 (N_5433,N_4744,N_4663);
or U5434 (N_5434,N_4608,N_4784);
or U5435 (N_5435,N_4987,N_4522);
or U5436 (N_5436,N_4825,N_4681);
nor U5437 (N_5437,N_4753,N_4756);
xor U5438 (N_5438,N_4991,N_4796);
or U5439 (N_5439,N_4517,N_4717);
and U5440 (N_5440,N_4731,N_4923);
nand U5441 (N_5441,N_4912,N_4544);
nand U5442 (N_5442,N_4896,N_4812);
xnor U5443 (N_5443,N_4917,N_4803);
or U5444 (N_5444,N_4650,N_4923);
or U5445 (N_5445,N_4641,N_4949);
nor U5446 (N_5446,N_4655,N_4971);
or U5447 (N_5447,N_4832,N_4765);
and U5448 (N_5448,N_4850,N_4818);
nor U5449 (N_5449,N_4696,N_4626);
nand U5450 (N_5450,N_4773,N_4520);
nor U5451 (N_5451,N_4818,N_4830);
and U5452 (N_5452,N_4674,N_4539);
xnor U5453 (N_5453,N_4821,N_4643);
xnor U5454 (N_5454,N_4798,N_4720);
xor U5455 (N_5455,N_4617,N_4548);
xor U5456 (N_5456,N_4558,N_4567);
nand U5457 (N_5457,N_4665,N_4934);
and U5458 (N_5458,N_4552,N_4996);
and U5459 (N_5459,N_4956,N_4507);
nand U5460 (N_5460,N_4890,N_4756);
or U5461 (N_5461,N_4796,N_4831);
nor U5462 (N_5462,N_4798,N_4847);
xor U5463 (N_5463,N_4502,N_4806);
xnor U5464 (N_5464,N_4670,N_4751);
nor U5465 (N_5465,N_4875,N_4941);
nand U5466 (N_5466,N_4698,N_4704);
or U5467 (N_5467,N_4778,N_4877);
xor U5468 (N_5468,N_4927,N_4617);
nor U5469 (N_5469,N_4532,N_4543);
nor U5470 (N_5470,N_4669,N_4558);
or U5471 (N_5471,N_4505,N_4657);
or U5472 (N_5472,N_4584,N_4536);
nand U5473 (N_5473,N_4818,N_4664);
and U5474 (N_5474,N_4699,N_4574);
xnor U5475 (N_5475,N_4598,N_4964);
and U5476 (N_5476,N_4755,N_4511);
nand U5477 (N_5477,N_4626,N_4924);
nand U5478 (N_5478,N_4553,N_4708);
xor U5479 (N_5479,N_4675,N_4763);
nand U5480 (N_5480,N_4579,N_4758);
nand U5481 (N_5481,N_4651,N_4877);
nand U5482 (N_5482,N_4933,N_4905);
nor U5483 (N_5483,N_4773,N_4866);
xnor U5484 (N_5484,N_4887,N_4560);
xor U5485 (N_5485,N_4624,N_4587);
xnor U5486 (N_5486,N_4655,N_4955);
xnor U5487 (N_5487,N_4742,N_4869);
and U5488 (N_5488,N_4897,N_4693);
xnor U5489 (N_5489,N_4712,N_4770);
and U5490 (N_5490,N_4800,N_4679);
xor U5491 (N_5491,N_4616,N_4986);
and U5492 (N_5492,N_4822,N_4793);
nand U5493 (N_5493,N_4900,N_4707);
xor U5494 (N_5494,N_4946,N_4751);
or U5495 (N_5495,N_4738,N_4695);
nand U5496 (N_5496,N_4775,N_4971);
nand U5497 (N_5497,N_4960,N_4748);
nand U5498 (N_5498,N_4564,N_4821);
nor U5499 (N_5499,N_4726,N_4758);
or U5500 (N_5500,N_5108,N_5372);
and U5501 (N_5501,N_5375,N_5203);
nor U5502 (N_5502,N_5141,N_5050);
xnor U5503 (N_5503,N_5148,N_5397);
nor U5504 (N_5504,N_5335,N_5303);
or U5505 (N_5505,N_5059,N_5448);
or U5506 (N_5506,N_5469,N_5330);
nand U5507 (N_5507,N_5009,N_5462);
and U5508 (N_5508,N_5013,N_5274);
and U5509 (N_5509,N_5112,N_5069);
xnor U5510 (N_5510,N_5295,N_5022);
nand U5511 (N_5511,N_5074,N_5019);
nand U5512 (N_5512,N_5166,N_5422);
nor U5513 (N_5513,N_5136,N_5264);
xnor U5514 (N_5514,N_5197,N_5045);
nand U5515 (N_5515,N_5114,N_5273);
and U5516 (N_5516,N_5037,N_5284);
or U5517 (N_5517,N_5426,N_5380);
nand U5518 (N_5518,N_5470,N_5345);
nand U5519 (N_5519,N_5368,N_5007);
nor U5520 (N_5520,N_5178,N_5119);
or U5521 (N_5521,N_5127,N_5350);
nand U5522 (N_5522,N_5058,N_5106);
or U5523 (N_5523,N_5493,N_5400);
or U5524 (N_5524,N_5078,N_5023);
or U5525 (N_5525,N_5488,N_5055);
nor U5526 (N_5526,N_5256,N_5317);
or U5527 (N_5527,N_5246,N_5314);
and U5528 (N_5528,N_5235,N_5447);
or U5529 (N_5529,N_5441,N_5340);
nor U5530 (N_5530,N_5071,N_5233);
nand U5531 (N_5531,N_5213,N_5103);
and U5532 (N_5532,N_5301,N_5001);
nor U5533 (N_5533,N_5424,N_5461);
nor U5534 (N_5534,N_5239,N_5205);
nor U5535 (N_5535,N_5128,N_5428);
and U5536 (N_5536,N_5342,N_5229);
or U5537 (N_5537,N_5320,N_5234);
or U5538 (N_5538,N_5312,N_5124);
or U5539 (N_5539,N_5225,N_5449);
nand U5540 (N_5540,N_5398,N_5404);
and U5541 (N_5541,N_5355,N_5433);
nor U5542 (N_5542,N_5297,N_5248);
nand U5543 (N_5543,N_5220,N_5268);
xnor U5544 (N_5544,N_5016,N_5231);
nor U5545 (N_5545,N_5145,N_5053);
xnor U5546 (N_5546,N_5362,N_5221);
nand U5547 (N_5547,N_5215,N_5173);
nor U5548 (N_5548,N_5155,N_5249);
nand U5549 (N_5549,N_5206,N_5430);
xnor U5550 (N_5550,N_5219,N_5230);
and U5551 (N_5551,N_5082,N_5432);
or U5552 (N_5552,N_5434,N_5327);
nor U5553 (N_5553,N_5495,N_5125);
and U5554 (N_5554,N_5113,N_5321);
and U5555 (N_5555,N_5122,N_5222);
and U5556 (N_5556,N_5391,N_5170);
xor U5557 (N_5557,N_5167,N_5476);
nand U5558 (N_5558,N_5253,N_5478);
nand U5559 (N_5559,N_5172,N_5459);
xor U5560 (N_5560,N_5263,N_5420);
and U5561 (N_5561,N_5138,N_5472);
or U5562 (N_5562,N_5280,N_5269);
xor U5563 (N_5563,N_5392,N_5323);
and U5564 (N_5564,N_5457,N_5440);
xnor U5565 (N_5565,N_5384,N_5159);
xor U5566 (N_5566,N_5004,N_5279);
xor U5567 (N_5567,N_5387,N_5287);
nand U5568 (N_5568,N_5099,N_5410);
and U5569 (N_5569,N_5032,N_5150);
or U5570 (N_5570,N_5336,N_5346);
xor U5571 (N_5571,N_5183,N_5395);
xor U5572 (N_5572,N_5038,N_5160);
xor U5573 (N_5573,N_5110,N_5043);
nand U5574 (N_5574,N_5438,N_5024);
and U5575 (N_5575,N_5014,N_5405);
nand U5576 (N_5576,N_5157,N_5188);
xnor U5577 (N_5577,N_5083,N_5463);
nand U5578 (N_5578,N_5111,N_5423);
and U5579 (N_5579,N_5015,N_5146);
nand U5580 (N_5580,N_5065,N_5254);
nor U5581 (N_5581,N_5326,N_5349);
and U5582 (N_5582,N_5169,N_5139);
nand U5583 (N_5583,N_5091,N_5465);
xnor U5584 (N_5584,N_5409,N_5377);
nor U5585 (N_5585,N_5067,N_5338);
xnor U5586 (N_5586,N_5270,N_5008);
or U5587 (N_5587,N_5399,N_5494);
nor U5588 (N_5588,N_5369,N_5105);
nor U5589 (N_5589,N_5218,N_5238);
and U5590 (N_5590,N_5163,N_5406);
nand U5591 (N_5591,N_5289,N_5176);
nor U5592 (N_5592,N_5277,N_5095);
and U5593 (N_5593,N_5240,N_5285);
xor U5594 (N_5594,N_5307,N_5325);
nor U5595 (N_5595,N_5418,N_5131);
nand U5596 (N_5596,N_5018,N_5356);
nor U5597 (N_5597,N_5484,N_5204);
or U5598 (N_5598,N_5132,N_5278);
or U5599 (N_5599,N_5208,N_5480);
or U5600 (N_5600,N_5427,N_5028);
nand U5601 (N_5601,N_5390,N_5026);
or U5602 (N_5602,N_5475,N_5396);
or U5603 (N_5603,N_5115,N_5195);
and U5604 (N_5604,N_5223,N_5352);
xor U5605 (N_5605,N_5381,N_5093);
nor U5606 (N_5606,N_5033,N_5079);
and U5607 (N_5607,N_5002,N_5492);
xor U5608 (N_5608,N_5247,N_5177);
nand U5609 (N_5609,N_5121,N_5416);
nand U5610 (N_5610,N_5486,N_5070);
or U5611 (N_5611,N_5066,N_5304);
and U5612 (N_5612,N_5436,N_5389);
or U5613 (N_5613,N_5064,N_5408);
xor U5614 (N_5614,N_5452,N_5156);
xor U5615 (N_5615,N_5034,N_5360);
nand U5616 (N_5616,N_5378,N_5097);
nor U5617 (N_5617,N_5437,N_5481);
nor U5618 (N_5618,N_5193,N_5134);
nand U5619 (N_5619,N_5123,N_5084);
xnor U5620 (N_5620,N_5000,N_5102);
and U5621 (N_5621,N_5402,N_5187);
and U5622 (N_5622,N_5107,N_5394);
nand U5623 (N_5623,N_5021,N_5151);
and U5624 (N_5624,N_5011,N_5162);
nand U5625 (N_5625,N_5057,N_5149);
xor U5626 (N_5626,N_5421,N_5444);
and U5627 (N_5627,N_5451,N_5242);
xor U5628 (N_5628,N_5454,N_5228);
nand U5629 (N_5629,N_5044,N_5025);
nand U5630 (N_5630,N_5168,N_5499);
nand U5631 (N_5631,N_5199,N_5383);
xnor U5632 (N_5632,N_5226,N_5036);
nand U5633 (N_5633,N_5089,N_5094);
nor U5634 (N_5634,N_5029,N_5407);
nor U5635 (N_5635,N_5329,N_5047);
or U5636 (N_5636,N_5117,N_5224);
nor U5637 (N_5637,N_5450,N_5485);
xor U5638 (N_5638,N_5458,N_5257);
and U5639 (N_5639,N_5140,N_5196);
or U5640 (N_5640,N_5184,N_5347);
or U5641 (N_5641,N_5147,N_5243);
xnor U5642 (N_5642,N_5386,N_5049);
and U5643 (N_5643,N_5361,N_5051);
nor U5644 (N_5644,N_5241,N_5498);
xor U5645 (N_5645,N_5088,N_5217);
nor U5646 (N_5646,N_5190,N_5275);
xnor U5647 (N_5647,N_5339,N_5265);
xor U5648 (N_5648,N_5298,N_5186);
nor U5649 (N_5649,N_5258,N_5046);
and U5650 (N_5650,N_5137,N_5471);
nor U5651 (N_5651,N_5490,N_5343);
nor U5652 (N_5652,N_5439,N_5161);
xor U5653 (N_5653,N_5216,N_5191);
nor U5654 (N_5654,N_5294,N_5308);
nand U5655 (N_5655,N_5042,N_5101);
xnor U5656 (N_5656,N_5332,N_5429);
nor U5657 (N_5657,N_5453,N_5291);
or U5658 (N_5658,N_5376,N_5385);
and U5659 (N_5659,N_5425,N_5096);
nor U5660 (N_5660,N_5006,N_5266);
nand U5661 (N_5661,N_5282,N_5181);
or U5662 (N_5662,N_5061,N_5063);
nand U5663 (N_5663,N_5252,N_5133);
xor U5664 (N_5664,N_5153,N_5272);
nand U5665 (N_5665,N_5413,N_5482);
nand U5666 (N_5666,N_5367,N_5473);
or U5667 (N_5667,N_5309,N_5202);
or U5668 (N_5668,N_5299,N_5292);
or U5669 (N_5669,N_5306,N_5316);
or U5670 (N_5670,N_5035,N_5143);
nand U5671 (N_5671,N_5371,N_5142);
nor U5672 (N_5672,N_5179,N_5086);
xor U5673 (N_5673,N_5185,N_5322);
nand U5674 (N_5674,N_5087,N_5017);
xnor U5675 (N_5675,N_5466,N_5040);
or U5676 (N_5676,N_5041,N_5062);
and U5677 (N_5677,N_5474,N_5232);
xor U5678 (N_5678,N_5353,N_5468);
nand U5679 (N_5679,N_5445,N_5180);
xnor U5680 (N_5680,N_5075,N_5104);
and U5681 (N_5681,N_5417,N_5003);
nor U5682 (N_5682,N_5250,N_5048);
nor U5683 (N_5683,N_5302,N_5401);
nor U5684 (N_5684,N_5175,N_5194);
nor U5685 (N_5685,N_5085,N_5158);
xor U5686 (N_5686,N_5374,N_5118);
and U5687 (N_5687,N_5271,N_5039);
xor U5688 (N_5688,N_5311,N_5348);
nor U5689 (N_5689,N_5276,N_5318);
nand U5690 (N_5690,N_5259,N_5479);
nor U5691 (N_5691,N_5286,N_5331);
xor U5692 (N_5692,N_5251,N_5100);
nand U5693 (N_5693,N_5054,N_5333);
xnor U5694 (N_5694,N_5456,N_5477);
nor U5695 (N_5695,N_5363,N_5487);
and U5696 (N_5696,N_5431,N_5315);
xnor U5697 (N_5697,N_5443,N_5357);
nor U5698 (N_5698,N_5060,N_5092);
nor U5699 (N_5699,N_5341,N_5351);
or U5700 (N_5700,N_5344,N_5152);
and U5701 (N_5701,N_5373,N_5198);
nor U5702 (N_5702,N_5379,N_5164);
nand U5703 (N_5703,N_5260,N_5403);
nor U5704 (N_5704,N_5244,N_5077);
xnor U5705 (N_5705,N_5319,N_5261);
nand U5706 (N_5706,N_5283,N_5245);
nor U5707 (N_5707,N_5300,N_5328);
and U5708 (N_5708,N_5366,N_5154);
or U5709 (N_5709,N_5237,N_5435);
xnor U5710 (N_5710,N_5210,N_5255);
xor U5711 (N_5711,N_5189,N_5056);
xor U5712 (N_5712,N_5460,N_5337);
xnor U5713 (N_5713,N_5030,N_5411);
nor U5714 (N_5714,N_5171,N_5135);
nand U5715 (N_5715,N_5120,N_5382);
xor U5716 (N_5716,N_5020,N_5081);
nor U5717 (N_5717,N_5227,N_5489);
nand U5718 (N_5718,N_5415,N_5412);
or U5719 (N_5719,N_5209,N_5214);
xor U5720 (N_5720,N_5174,N_5281);
or U5721 (N_5721,N_5358,N_5491);
and U5722 (N_5722,N_5098,N_5052);
xor U5723 (N_5723,N_5012,N_5109);
nor U5724 (N_5724,N_5073,N_5305);
nor U5725 (N_5725,N_5116,N_5496);
or U5726 (N_5726,N_5354,N_5334);
xnor U5727 (N_5727,N_5010,N_5467);
nor U5728 (N_5728,N_5296,N_5211);
nor U5729 (N_5729,N_5293,N_5455);
nand U5730 (N_5730,N_5201,N_5005);
or U5731 (N_5731,N_5072,N_5324);
nand U5732 (N_5732,N_5370,N_5365);
or U5733 (N_5733,N_5364,N_5090);
xor U5734 (N_5734,N_5144,N_5027);
nor U5735 (N_5735,N_5483,N_5313);
and U5736 (N_5736,N_5236,N_5419);
nor U5737 (N_5737,N_5129,N_5290);
or U5738 (N_5738,N_5442,N_5165);
nor U5739 (N_5739,N_5192,N_5200);
xor U5740 (N_5740,N_5182,N_5464);
and U5741 (N_5741,N_5414,N_5388);
nand U5742 (N_5742,N_5068,N_5310);
and U5743 (N_5743,N_5130,N_5207);
and U5744 (N_5744,N_5076,N_5288);
xor U5745 (N_5745,N_5080,N_5267);
or U5746 (N_5746,N_5393,N_5446);
xnor U5747 (N_5747,N_5359,N_5497);
or U5748 (N_5748,N_5212,N_5126);
nor U5749 (N_5749,N_5031,N_5262);
or U5750 (N_5750,N_5268,N_5189);
or U5751 (N_5751,N_5083,N_5258);
nand U5752 (N_5752,N_5098,N_5347);
and U5753 (N_5753,N_5144,N_5347);
nand U5754 (N_5754,N_5151,N_5271);
or U5755 (N_5755,N_5074,N_5340);
or U5756 (N_5756,N_5122,N_5084);
nor U5757 (N_5757,N_5441,N_5277);
nor U5758 (N_5758,N_5391,N_5208);
xnor U5759 (N_5759,N_5309,N_5180);
nand U5760 (N_5760,N_5049,N_5462);
nand U5761 (N_5761,N_5414,N_5221);
or U5762 (N_5762,N_5295,N_5362);
nand U5763 (N_5763,N_5457,N_5048);
and U5764 (N_5764,N_5250,N_5199);
nor U5765 (N_5765,N_5154,N_5432);
xnor U5766 (N_5766,N_5192,N_5280);
nor U5767 (N_5767,N_5334,N_5454);
and U5768 (N_5768,N_5148,N_5054);
xnor U5769 (N_5769,N_5068,N_5081);
and U5770 (N_5770,N_5113,N_5364);
or U5771 (N_5771,N_5255,N_5432);
nor U5772 (N_5772,N_5297,N_5147);
nor U5773 (N_5773,N_5145,N_5086);
xor U5774 (N_5774,N_5431,N_5260);
and U5775 (N_5775,N_5459,N_5160);
nor U5776 (N_5776,N_5298,N_5432);
and U5777 (N_5777,N_5446,N_5051);
or U5778 (N_5778,N_5193,N_5127);
nand U5779 (N_5779,N_5399,N_5168);
xor U5780 (N_5780,N_5006,N_5390);
or U5781 (N_5781,N_5449,N_5140);
or U5782 (N_5782,N_5104,N_5155);
and U5783 (N_5783,N_5481,N_5220);
and U5784 (N_5784,N_5316,N_5157);
and U5785 (N_5785,N_5476,N_5359);
and U5786 (N_5786,N_5165,N_5459);
nor U5787 (N_5787,N_5445,N_5403);
nand U5788 (N_5788,N_5422,N_5191);
nand U5789 (N_5789,N_5342,N_5479);
and U5790 (N_5790,N_5279,N_5250);
and U5791 (N_5791,N_5326,N_5271);
nand U5792 (N_5792,N_5122,N_5219);
nor U5793 (N_5793,N_5092,N_5205);
nand U5794 (N_5794,N_5473,N_5270);
nand U5795 (N_5795,N_5430,N_5232);
or U5796 (N_5796,N_5080,N_5448);
xor U5797 (N_5797,N_5211,N_5337);
and U5798 (N_5798,N_5423,N_5352);
or U5799 (N_5799,N_5109,N_5082);
or U5800 (N_5800,N_5040,N_5313);
nand U5801 (N_5801,N_5472,N_5221);
or U5802 (N_5802,N_5192,N_5215);
nor U5803 (N_5803,N_5458,N_5122);
or U5804 (N_5804,N_5468,N_5403);
or U5805 (N_5805,N_5419,N_5280);
nand U5806 (N_5806,N_5261,N_5399);
nand U5807 (N_5807,N_5370,N_5343);
and U5808 (N_5808,N_5261,N_5051);
xnor U5809 (N_5809,N_5257,N_5471);
nand U5810 (N_5810,N_5243,N_5029);
nand U5811 (N_5811,N_5106,N_5008);
xor U5812 (N_5812,N_5281,N_5280);
nand U5813 (N_5813,N_5041,N_5400);
xnor U5814 (N_5814,N_5064,N_5076);
nand U5815 (N_5815,N_5068,N_5071);
or U5816 (N_5816,N_5374,N_5364);
xnor U5817 (N_5817,N_5469,N_5278);
and U5818 (N_5818,N_5074,N_5199);
or U5819 (N_5819,N_5448,N_5460);
nor U5820 (N_5820,N_5329,N_5461);
and U5821 (N_5821,N_5150,N_5492);
nor U5822 (N_5822,N_5039,N_5261);
nand U5823 (N_5823,N_5071,N_5228);
nor U5824 (N_5824,N_5375,N_5019);
nand U5825 (N_5825,N_5400,N_5183);
and U5826 (N_5826,N_5198,N_5090);
nand U5827 (N_5827,N_5153,N_5459);
nor U5828 (N_5828,N_5145,N_5290);
xor U5829 (N_5829,N_5393,N_5460);
and U5830 (N_5830,N_5462,N_5309);
nand U5831 (N_5831,N_5293,N_5191);
nor U5832 (N_5832,N_5019,N_5101);
xnor U5833 (N_5833,N_5408,N_5032);
or U5834 (N_5834,N_5171,N_5155);
or U5835 (N_5835,N_5037,N_5408);
nand U5836 (N_5836,N_5409,N_5292);
nand U5837 (N_5837,N_5017,N_5266);
and U5838 (N_5838,N_5115,N_5295);
or U5839 (N_5839,N_5013,N_5489);
or U5840 (N_5840,N_5395,N_5311);
and U5841 (N_5841,N_5103,N_5456);
nand U5842 (N_5842,N_5126,N_5133);
or U5843 (N_5843,N_5296,N_5344);
nand U5844 (N_5844,N_5153,N_5062);
xnor U5845 (N_5845,N_5151,N_5346);
nor U5846 (N_5846,N_5079,N_5493);
nor U5847 (N_5847,N_5007,N_5419);
xnor U5848 (N_5848,N_5236,N_5324);
xnor U5849 (N_5849,N_5051,N_5284);
nand U5850 (N_5850,N_5201,N_5088);
xnor U5851 (N_5851,N_5253,N_5013);
or U5852 (N_5852,N_5147,N_5304);
or U5853 (N_5853,N_5184,N_5265);
or U5854 (N_5854,N_5049,N_5116);
and U5855 (N_5855,N_5176,N_5413);
xnor U5856 (N_5856,N_5174,N_5085);
nor U5857 (N_5857,N_5169,N_5151);
nor U5858 (N_5858,N_5353,N_5065);
nand U5859 (N_5859,N_5125,N_5351);
nor U5860 (N_5860,N_5389,N_5419);
xnor U5861 (N_5861,N_5330,N_5416);
or U5862 (N_5862,N_5172,N_5160);
nand U5863 (N_5863,N_5448,N_5363);
and U5864 (N_5864,N_5170,N_5019);
xor U5865 (N_5865,N_5402,N_5056);
nor U5866 (N_5866,N_5099,N_5433);
nand U5867 (N_5867,N_5112,N_5443);
xor U5868 (N_5868,N_5123,N_5027);
or U5869 (N_5869,N_5236,N_5335);
or U5870 (N_5870,N_5124,N_5332);
xnor U5871 (N_5871,N_5157,N_5407);
or U5872 (N_5872,N_5278,N_5220);
or U5873 (N_5873,N_5058,N_5358);
or U5874 (N_5874,N_5058,N_5090);
or U5875 (N_5875,N_5187,N_5277);
xnor U5876 (N_5876,N_5202,N_5407);
and U5877 (N_5877,N_5042,N_5014);
nor U5878 (N_5878,N_5153,N_5189);
xor U5879 (N_5879,N_5040,N_5496);
and U5880 (N_5880,N_5304,N_5250);
nand U5881 (N_5881,N_5095,N_5060);
nor U5882 (N_5882,N_5222,N_5386);
or U5883 (N_5883,N_5197,N_5175);
nand U5884 (N_5884,N_5040,N_5353);
nand U5885 (N_5885,N_5303,N_5169);
and U5886 (N_5886,N_5010,N_5306);
or U5887 (N_5887,N_5484,N_5241);
or U5888 (N_5888,N_5218,N_5202);
xnor U5889 (N_5889,N_5322,N_5224);
nand U5890 (N_5890,N_5360,N_5292);
nand U5891 (N_5891,N_5280,N_5152);
nand U5892 (N_5892,N_5306,N_5006);
xnor U5893 (N_5893,N_5051,N_5472);
nor U5894 (N_5894,N_5068,N_5095);
nor U5895 (N_5895,N_5006,N_5302);
xnor U5896 (N_5896,N_5150,N_5221);
nor U5897 (N_5897,N_5327,N_5482);
nor U5898 (N_5898,N_5429,N_5054);
xnor U5899 (N_5899,N_5046,N_5134);
and U5900 (N_5900,N_5238,N_5378);
and U5901 (N_5901,N_5053,N_5478);
nor U5902 (N_5902,N_5455,N_5072);
xnor U5903 (N_5903,N_5451,N_5327);
or U5904 (N_5904,N_5466,N_5073);
nand U5905 (N_5905,N_5493,N_5144);
or U5906 (N_5906,N_5437,N_5069);
nor U5907 (N_5907,N_5227,N_5052);
and U5908 (N_5908,N_5013,N_5327);
nand U5909 (N_5909,N_5411,N_5276);
nor U5910 (N_5910,N_5015,N_5134);
and U5911 (N_5911,N_5436,N_5013);
or U5912 (N_5912,N_5192,N_5026);
or U5913 (N_5913,N_5263,N_5042);
or U5914 (N_5914,N_5151,N_5190);
or U5915 (N_5915,N_5462,N_5135);
and U5916 (N_5916,N_5235,N_5239);
nor U5917 (N_5917,N_5174,N_5188);
or U5918 (N_5918,N_5304,N_5102);
nor U5919 (N_5919,N_5449,N_5360);
xnor U5920 (N_5920,N_5144,N_5486);
nand U5921 (N_5921,N_5339,N_5122);
nor U5922 (N_5922,N_5260,N_5065);
xnor U5923 (N_5923,N_5052,N_5314);
xnor U5924 (N_5924,N_5474,N_5348);
xnor U5925 (N_5925,N_5008,N_5168);
or U5926 (N_5926,N_5058,N_5322);
nor U5927 (N_5927,N_5000,N_5413);
nand U5928 (N_5928,N_5255,N_5079);
or U5929 (N_5929,N_5404,N_5178);
nor U5930 (N_5930,N_5035,N_5318);
and U5931 (N_5931,N_5161,N_5174);
nand U5932 (N_5932,N_5293,N_5451);
nor U5933 (N_5933,N_5162,N_5026);
xnor U5934 (N_5934,N_5282,N_5246);
xnor U5935 (N_5935,N_5106,N_5485);
or U5936 (N_5936,N_5282,N_5070);
xnor U5937 (N_5937,N_5054,N_5393);
nand U5938 (N_5938,N_5278,N_5356);
nor U5939 (N_5939,N_5070,N_5259);
nand U5940 (N_5940,N_5160,N_5153);
nand U5941 (N_5941,N_5127,N_5207);
nor U5942 (N_5942,N_5173,N_5048);
nand U5943 (N_5943,N_5358,N_5128);
and U5944 (N_5944,N_5331,N_5255);
nand U5945 (N_5945,N_5182,N_5221);
and U5946 (N_5946,N_5109,N_5010);
xnor U5947 (N_5947,N_5414,N_5210);
xnor U5948 (N_5948,N_5484,N_5188);
or U5949 (N_5949,N_5022,N_5053);
nand U5950 (N_5950,N_5264,N_5499);
and U5951 (N_5951,N_5479,N_5232);
nand U5952 (N_5952,N_5350,N_5419);
nor U5953 (N_5953,N_5230,N_5239);
nand U5954 (N_5954,N_5018,N_5169);
nand U5955 (N_5955,N_5245,N_5325);
and U5956 (N_5956,N_5469,N_5248);
nor U5957 (N_5957,N_5367,N_5006);
xnor U5958 (N_5958,N_5291,N_5486);
nand U5959 (N_5959,N_5246,N_5243);
nor U5960 (N_5960,N_5369,N_5182);
xnor U5961 (N_5961,N_5060,N_5371);
or U5962 (N_5962,N_5068,N_5177);
nor U5963 (N_5963,N_5296,N_5430);
and U5964 (N_5964,N_5151,N_5088);
nand U5965 (N_5965,N_5237,N_5352);
xnor U5966 (N_5966,N_5327,N_5352);
xor U5967 (N_5967,N_5047,N_5392);
nor U5968 (N_5968,N_5192,N_5291);
and U5969 (N_5969,N_5191,N_5330);
and U5970 (N_5970,N_5328,N_5232);
or U5971 (N_5971,N_5315,N_5179);
nand U5972 (N_5972,N_5187,N_5204);
and U5973 (N_5973,N_5431,N_5048);
xor U5974 (N_5974,N_5346,N_5426);
and U5975 (N_5975,N_5346,N_5400);
or U5976 (N_5976,N_5187,N_5337);
and U5977 (N_5977,N_5111,N_5147);
nor U5978 (N_5978,N_5150,N_5071);
and U5979 (N_5979,N_5156,N_5444);
xor U5980 (N_5980,N_5412,N_5242);
nor U5981 (N_5981,N_5242,N_5392);
nor U5982 (N_5982,N_5389,N_5281);
nor U5983 (N_5983,N_5401,N_5061);
nor U5984 (N_5984,N_5218,N_5162);
nor U5985 (N_5985,N_5104,N_5487);
nand U5986 (N_5986,N_5001,N_5463);
or U5987 (N_5987,N_5112,N_5049);
nor U5988 (N_5988,N_5195,N_5094);
and U5989 (N_5989,N_5320,N_5475);
xnor U5990 (N_5990,N_5111,N_5210);
nor U5991 (N_5991,N_5015,N_5247);
and U5992 (N_5992,N_5417,N_5066);
xor U5993 (N_5993,N_5210,N_5059);
or U5994 (N_5994,N_5371,N_5292);
nor U5995 (N_5995,N_5010,N_5114);
nand U5996 (N_5996,N_5289,N_5378);
and U5997 (N_5997,N_5351,N_5183);
nand U5998 (N_5998,N_5026,N_5331);
and U5999 (N_5999,N_5037,N_5205);
xnor U6000 (N_6000,N_5971,N_5636);
nand U6001 (N_6001,N_5561,N_5877);
and U6002 (N_6002,N_5967,N_5667);
or U6003 (N_6003,N_5943,N_5835);
or U6004 (N_6004,N_5859,N_5534);
nand U6005 (N_6005,N_5870,N_5676);
or U6006 (N_6006,N_5840,N_5749);
or U6007 (N_6007,N_5845,N_5539);
and U6008 (N_6008,N_5926,N_5730);
and U6009 (N_6009,N_5989,N_5772);
nand U6010 (N_6010,N_5819,N_5898);
nand U6011 (N_6011,N_5707,N_5856);
or U6012 (N_6012,N_5950,N_5713);
and U6013 (N_6013,N_5661,N_5813);
xor U6014 (N_6014,N_5654,N_5701);
xnor U6015 (N_6015,N_5564,N_5987);
or U6016 (N_6016,N_5585,N_5786);
nand U6017 (N_6017,N_5921,N_5928);
or U6018 (N_6018,N_5526,N_5611);
nor U6019 (N_6019,N_5597,N_5900);
nand U6020 (N_6020,N_5640,N_5836);
nor U6021 (N_6021,N_5624,N_5897);
or U6022 (N_6022,N_5711,N_5522);
and U6023 (N_6023,N_5861,N_5664);
nand U6024 (N_6024,N_5691,N_5718);
or U6025 (N_6025,N_5988,N_5940);
and U6026 (N_6026,N_5991,N_5964);
or U6027 (N_6027,N_5675,N_5797);
and U6028 (N_6028,N_5885,N_5717);
xnor U6029 (N_6029,N_5848,N_5773);
or U6030 (N_6030,N_5603,N_5849);
and U6031 (N_6031,N_5830,N_5951);
nor U6032 (N_6032,N_5532,N_5947);
nand U6033 (N_6033,N_5702,N_5710);
nor U6034 (N_6034,N_5756,N_5604);
nand U6035 (N_6035,N_5720,N_5591);
nor U6036 (N_6036,N_5980,N_5925);
or U6037 (N_6037,N_5891,N_5868);
xnor U6038 (N_6038,N_5945,N_5789);
nand U6039 (N_6039,N_5699,N_5931);
nor U6040 (N_6040,N_5686,N_5714);
and U6041 (N_6041,N_5761,N_5540);
xnor U6042 (N_6042,N_5935,N_5723);
or U6043 (N_6043,N_5649,N_5847);
or U6044 (N_6044,N_5792,N_5906);
nand U6045 (N_6045,N_5937,N_5881);
xor U6046 (N_6046,N_5765,N_5796);
xnor U6047 (N_6047,N_5529,N_5893);
nor U6048 (N_6048,N_5791,N_5729);
or U6049 (N_6049,N_5975,N_5703);
xor U6050 (N_6050,N_5501,N_5787);
xnor U6051 (N_6051,N_5504,N_5509);
nor U6052 (N_6052,N_5584,N_5630);
xnor U6053 (N_6053,N_5565,N_5735);
nand U6054 (N_6054,N_5556,N_5875);
nor U6055 (N_6055,N_5957,N_5531);
xor U6056 (N_6056,N_5569,N_5721);
nand U6057 (N_6057,N_5738,N_5758);
nand U6058 (N_6058,N_5650,N_5916);
xnor U6059 (N_6059,N_5606,N_5521);
nand U6060 (N_6060,N_5719,N_5913);
or U6061 (N_6061,N_5983,N_5985);
xnor U6062 (N_6062,N_5764,N_5645);
or U6063 (N_6063,N_5642,N_5660);
and U6064 (N_6064,N_5579,N_5523);
and U6065 (N_6065,N_5613,N_5958);
or U6066 (N_6066,N_5737,N_5771);
or U6067 (N_6067,N_5984,N_5644);
and U6068 (N_6068,N_5551,N_5949);
nor U6069 (N_6069,N_5862,N_5618);
or U6070 (N_6070,N_5995,N_5709);
nor U6071 (N_6071,N_5511,N_5643);
nor U6072 (N_6072,N_5956,N_5646);
nor U6073 (N_6073,N_5527,N_5700);
nand U6074 (N_6074,N_5927,N_5508);
nand U6075 (N_6075,N_5982,N_5586);
and U6076 (N_6076,N_5879,N_5939);
or U6077 (N_6077,N_5750,N_5742);
and U6078 (N_6078,N_5555,N_5566);
and U6079 (N_6079,N_5576,N_5571);
and U6080 (N_6080,N_5657,N_5651);
or U6081 (N_6081,N_5697,N_5970);
or U6082 (N_6082,N_5652,N_5878);
or U6083 (N_6083,N_5770,N_5778);
or U6084 (N_6084,N_5823,N_5816);
nor U6085 (N_6085,N_5692,N_5938);
nand U6086 (N_6086,N_5903,N_5623);
nor U6087 (N_6087,N_5743,N_5588);
nand U6088 (N_6088,N_5698,N_5766);
nor U6089 (N_6089,N_5860,N_5788);
nand U6090 (N_6090,N_5963,N_5635);
or U6091 (N_6091,N_5867,N_5972);
nor U6092 (N_6092,N_5615,N_5799);
and U6093 (N_6093,N_5994,N_5929);
xnor U6094 (N_6094,N_5869,N_5594);
xnor U6095 (N_6095,N_5874,N_5533);
or U6096 (N_6096,N_5593,N_5706);
or U6097 (N_6097,N_5517,N_5768);
or U6098 (N_6098,N_5748,N_5932);
and U6099 (N_6099,N_5827,N_5844);
xor U6100 (N_6100,N_5923,N_5577);
and U6101 (N_6101,N_5818,N_5518);
nor U6102 (N_6102,N_5582,N_5689);
and U6103 (N_6103,N_5690,N_5670);
nand U6104 (N_6104,N_5996,N_5519);
xnor U6105 (N_6105,N_5658,N_5560);
and U6106 (N_6106,N_5696,N_5866);
nor U6107 (N_6107,N_5863,N_5887);
and U6108 (N_6108,N_5746,N_5888);
xnor U6109 (N_6109,N_5922,N_5662);
and U6110 (N_6110,N_5685,N_5572);
xor U6111 (N_6111,N_5815,N_5632);
nor U6112 (N_6112,N_5600,N_5965);
xnor U6113 (N_6113,N_5781,N_5920);
and U6114 (N_6114,N_5802,N_5824);
or U6115 (N_6115,N_5633,N_5677);
or U6116 (N_6116,N_5784,N_5812);
and U6117 (N_6117,N_5679,N_5776);
nand U6118 (N_6118,N_5548,N_5678);
nor U6119 (N_6119,N_5736,N_5727);
xor U6120 (N_6120,N_5790,N_5538);
xnor U6121 (N_6121,N_5656,N_5915);
and U6122 (N_6122,N_5934,N_5933);
xnor U6123 (N_6123,N_5575,N_5598);
nand U6124 (N_6124,N_5946,N_5782);
or U6125 (N_6125,N_5568,N_5545);
and U6126 (N_6126,N_5552,N_5687);
and U6127 (N_6127,N_5546,N_5665);
nand U6128 (N_6128,N_5841,N_5858);
or U6129 (N_6129,N_5514,N_5744);
xnor U6130 (N_6130,N_5745,N_5919);
nand U6131 (N_6131,N_5739,N_5864);
nand U6132 (N_6132,N_5638,N_5528);
or U6133 (N_6133,N_5506,N_5833);
nand U6134 (N_6134,N_5831,N_5828);
xor U6135 (N_6135,N_5592,N_5674);
nand U6136 (N_6136,N_5631,N_5754);
xnor U6137 (N_6137,N_5637,N_5639);
xor U6138 (N_6138,N_5974,N_5554);
nor U6139 (N_6139,N_5977,N_5890);
and U6140 (N_6140,N_5805,N_5608);
xnor U6141 (N_6141,N_5952,N_5502);
nor U6142 (N_6142,N_5751,N_5904);
or U6143 (N_6143,N_5948,N_5817);
xnor U6144 (N_6144,N_5850,N_5684);
or U6145 (N_6145,N_5857,N_5587);
xnor U6146 (N_6146,N_5562,N_5590);
and U6147 (N_6147,N_5680,N_5852);
or U6148 (N_6148,N_5820,N_5992);
nand U6149 (N_6149,N_5894,N_5581);
and U6150 (N_6150,N_5614,N_5801);
xor U6151 (N_6151,N_5693,N_5601);
nor U6152 (N_6152,N_5541,N_5573);
nand U6153 (N_6153,N_5990,N_5973);
or U6154 (N_6154,N_5871,N_5808);
nand U6155 (N_6155,N_5780,N_5580);
and U6156 (N_6156,N_5741,N_5912);
or U6157 (N_6157,N_5978,N_5825);
or U6158 (N_6158,N_5663,N_5682);
xnor U6159 (N_6159,N_5671,N_5503);
nor U6160 (N_6160,N_5648,N_5583);
nor U6161 (N_6161,N_5883,N_5832);
nor U6162 (N_6162,N_5872,N_5954);
nand U6163 (N_6163,N_5753,N_5767);
nor U6164 (N_6164,N_5821,N_5837);
nor U6165 (N_6165,N_5999,N_5769);
or U6166 (N_6166,N_5549,N_5513);
or U6167 (N_6167,N_5731,N_5524);
xor U6168 (N_6168,N_5733,N_5607);
nand U6169 (N_6169,N_5843,N_5793);
and U6170 (N_6170,N_5694,N_5734);
nand U6171 (N_6171,N_5617,N_5629);
nand U6172 (N_6172,N_5838,N_5627);
and U6173 (N_6173,N_5775,N_5763);
or U6174 (N_6174,N_5798,N_5616);
or U6175 (N_6175,N_5537,N_5563);
xor U6176 (N_6176,N_5530,N_5909);
nand U6177 (N_6177,N_5804,N_5732);
and U6178 (N_6178,N_5889,N_5882);
xnor U6179 (N_6179,N_5961,N_5621);
and U6180 (N_6180,N_5774,N_5515);
and U6181 (N_6181,N_5612,N_5544);
xor U6182 (N_6182,N_5578,N_5704);
and U6183 (N_6183,N_5558,N_5892);
nor U6184 (N_6184,N_5553,N_5854);
xnor U6185 (N_6185,N_5683,N_5899);
xnor U6186 (N_6186,N_5966,N_5647);
nor U6187 (N_6187,N_5902,N_5777);
xnor U6188 (N_6188,N_5557,N_5543);
nor U6189 (N_6189,N_5542,N_5550);
or U6190 (N_6190,N_5814,N_5986);
nor U6191 (N_6191,N_5596,N_5811);
xnor U6192 (N_6192,N_5525,N_5510);
nand U6193 (N_6193,N_5512,N_5655);
nand U6194 (N_6194,N_5785,N_5896);
xnor U6195 (N_6195,N_5567,N_5705);
nor U6196 (N_6196,N_5998,N_5634);
and U6197 (N_6197,N_5747,N_5884);
nand U6198 (N_6198,N_5779,N_5880);
or U6199 (N_6199,N_5976,N_5834);
nor U6200 (N_6200,N_5979,N_5800);
or U6201 (N_6201,N_5944,N_5851);
xor U6202 (N_6202,N_5806,N_5936);
or U6203 (N_6203,N_5842,N_5993);
nand U6204 (N_6204,N_5911,N_5803);
nand U6205 (N_6205,N_5942,N_5917);
nor U6206 (N_6206,N_5535,N_5599);
nand U6207 (N_6207,N_5873,N_5914);
xor U6208 (N_6208,N_5895,N_5570);
xor U6209 (N_6209,N_5725,N_5997);
nand U6210 (N_6210,N_5901,N_5740);
xnor U6211 (N_6211,N_5609,N_5688);
nand U6212 (N_6212,N_5829,N_5726);
nand U6213 (N_6213,N_5955,N_5622);
and U6214 (N_6214,N_5905,N_5516);
and U6215 (N_6215,N_5716,N_5853);
nand U6216 (N_6216,N_5547,N_5960);
and U6217 (N_6217,N_5620,N_5619);
and U6218 (N_6218,N_5759,N_5809);
and U6219 (N_6219,N_5795,N_5672);
or U6220 (N_6220,N_5595,N_5783);
nand U6221 (N_6221,N_5762,N_5755);
or U6222 (N_6222,N_5959,N_5695);
xnor U6223 (N_6223,N_5953,N_5826);
nor U6224 (N_6224,N_5628,N_5536);
or U6225 (N_6225,N_5941,N_5669);
nor U6226 (N_6226,N_5507,N_5810);
and U6227 (N_6227,N_5641,N_5668);
xor U6228 (N_6228,N_5886,N_5822);
or U6229 (N_6229,N_5605,N_5855);
and U6230 (N_6230,N_5715,N_5500);
nor U6231 (N_6231,N_5918,N_5981);
xnor U6232 (N_6232,N_5760,N_5625);
or U6233 (N_6233,N_5968,N_5907);
or U6234 (N_6234,N_5924,N_5910);
nand U6235 (N_6235,N_5589,N_5757);
xnor U6236 (N_6236,N_5722,N_5807);
nor U6237 (N_6237,N_5505,N_5659);
nor U6238 (N_6238,N_5673,N_5908);
nor U6239 (N_6239,N_5610,N_5962);
xor U6240 (N_6240,N_5752,N_5839);
nand U6241 (N_6241,N_5846,N_5724);
and U6242 (N_6242,N_5865,N_5559);
or U6243 (N_6243,N_5681,N_5602);
nand U6244 (N_6244,N_5969,N_5794);
nor U6245 (N_6245,N_5728,N_5653);
and U6246 (N_6246,N_5520,N_5708);
or U6247 (N_6247,N_5666,N_5876);
xnor U6248 (N_6248,N_5712,N_5574);
nor U6249 (N_6249,N_5930,N_5626);
nand U6250 (N_6250,N_5503,N_5720);
xor U6251 (N_6251,N_5965,N_5727);
and U6252 (N_6252,N_5976,N_5553);
xnor U6253 (N_6253,N_5638,N_5918);
xor U6254 (N_6254,N_5871,N_5575);
nand U6255 (N_6255,N_5825,N_5570);
nor U6256 (N_6256,N_5968,N_5991);
or U6257 (N_6257,N_5967,N_5801);
or U6258 (N_6258,N_5521,N_5687);
nand U6259 (N_6259,N_5592,N_5544);
or U6260 (N_6260,N_5590,N_5868);
or U6261 (N_6261,N_5934,N_5866);
xor U6262 (N_6262,N_5543,N_5783);
xnor U6263 (N_6263,N_5585,N_5560);
xnor U6264 (N_6264,N_5745,N_5910);
xor U6265 (N_6265,N_5716,N_5965);
nor U6266 (N_6266,N_5923,N_5727);
xnor U6267 (N_6267,N_5505,N_5694);
and U6268 (N_6268,N_5995,N_5784);
nor U6269 (N_6269,N_5777,N_5545);
or U6270 (N_6270,N_5720,N_5913);
or U6271 (N_6271,N_5929,N_5999);
nor U6272 (N_6272,N_5680,N_5876);
and U6273 (N_6273,N_5658,N_5599);
xor U6274 (N_6274,N_5914,N_5633);
and U6275 (N_6275,N_5626,N_5562);
nor U6276 (N_6276,N_5812,N_5972);
nand U6277 (N_6277,N_5540,N_5723);
nor U6278 (N_6278,N_5918,N_5812);
and U6279 (N_6279,N_5959,N_5551);
nand U6280 (N_6280,N_5682,N_5508);
and U6281 (N_6281,N_5551,N_5670);
xor U6282 (N_6282,N_5802,N_5646);
nand U6283 (N_6283,N_5556,N_5950);
nor U6284 (N_6284,N_5654,N_5640);
xnor U6285 (N_6285,N_5673,N_5792);
nand U6286 (N_6286,N_5705,N_5791);
xor U6287 (N_6287,N_5877,N_5646);
nand U6288 (N_6288,N_5889,N_5852);
or U6289 (N_6289,N_5869,N_5677);
or U6290 (N_6290,N_5716,N_5842);
and U6291 (N_6291,N_5678,N_5634);
and U6292 (N_6292,N_5632,N_5619);
and U6293 (N_6293,N_5580,N_5769);
nand U6294 (N_6294,N_5992,N_5583);
xor U6295 (N_6295,N_5837,N_5858);
and U6296 (N_6296,N_5603,N_5551);
or U6297 (N_6297,N_5638,N_5694);
or U6298 (N_6298,N_5869,N_5705);
xor U6299 (N_6299,N_5772,N_5705);
xnor U6300 (N_6300,N_5850,N_5977);
or U6301 (N_6301,N_5801,N_5961);
nor U6302 (N_6302,N_5540,N_5620);
and U6303 (N_6303,N_5527,N_5999);
nor U6304 (N_6304,N_5826,N_5500);
xnor U6305 (N_6305,N_5925,N_5994);
or U6306 (N_6306,N_5731,N_5844);
and U6307 (N_6307,N_5569,N_5555);
nand U6308 (N_6308,N_5861,N_5545);
nor U6309 (N_6309,N_5561,N_5862);
nor U6310 (N_6310,N_5826,N_5643);
xnor U6311 (N_6311,N_5566,N_5610);
nor U6312 (N_6312,N_5623,N_5844);
or U6313 (N_6313,N_5874,N_5543);
nor U6314 (N_6314,N_5692,N_5701);
xor U6315 (N_6315,N_5766,N_5703);
xor U6316 (N_6316,N_5805,N_5573);
and U6317 (N_6317,N_5899,N_5659);
nand U6318 (N_6318,N_5773,N_5737);
xnor U6319 (N_6319,N_5539,N_5542);
and U6320 (N_6320,N_5862,N_5530);
xor U6321 (N_6321,N_5579,N_5712);
xnor U6322 (N_6322,N_5684,N_5691);
nand U6323 (N_6323,N_5571,N_5895);
or U6324 (N_6324,N_5726,N_5537);
xor U6325 (N_6325,N_5727,N_5992);
nand U6326 (N_6326,N_5971,N_5701);
nand U6327 (N_6327,N_5963,N_5920);
xor U6328 (N_6328,N_5710,N_5569);
and U6329 (N_6329,N_5817,N_5995);
and U6330 (N_6330,N_5823,N_5634);
and U6331 (N_6331,N_5674,N_5974);
xor U6332 (N_6332,N_5542,N_5829);
or U6333 (N_6333,N_5770,N_5697);
xnor U6334 (N_6334,N_5871,N_5864);
xnor U6335 (N_6335,N_5811,N_5765);
or U6336 (N_6336,N_5831,N_5542);
nor U6337 (N_6337,N_5839,N_5543);
and U6338 (N_6338,N_5760,N_5970);
and U6339 (N_6339,N_5927,N_5727);
and U6340 (N_6340,N_5763,N_5737);
and U6341 (N_6341,N_5939,N_5551);
xnor U6342 (N_6342,N_5912,N_5807);
xnor U6343 (N_6343,N_5966,N_5658);
nor U6344 (N_6344,N_5982,N_5974);
nand U6345 (N_6345,N_5677,N_5854);
xor U6346 (N_6346,N_5752,N_5857);
xor U6347 (N_6347,N_5667,N_5981);
nor U6348 (N_6348,N_5795,N_5516);
nand U6349 (N_6349,N_5953,N_5664);
and U6350 (N_6350,N_5520,N_5610);
xnor U6351 (N_6351,N_5589,N_5730);
xnor U6352 (N_6352,N_5653,N_5505);
xor U6353 (N_6353,N_5520,N_5522);
or U6354 (N_6354,N_5697,N_5894);
nand U6355 (N_6355,N_5706,N_5568);
xnor U6356 (N_6356,N_5505,N_5667);
nor U6357 (N_6357,N_5780,N_5749);
nor U6358 (N_6358,N_5965,N_5659);
xor U6359 (N_6359,N_5772,N_5875);
xnor U6360 (N_6360,N_5954,N_5764);
or U6361 (N_6361,N_5945,N_5738);
xnor U6362 (N_6362,N_5893,N_5965);
xnor U6363 (N_6363,N_5554,N_5840);
nand U6364 (N_6364,N_5990,N_5650);
xnor U6365 (N_6365,N_5626,N_5660);
nor U6366 (N_6366,N_5900,N_5908);
nand U6367 (N_6367,N_5778,N_5967);
nand U6368 (N_6368,N_5733,N_5712);
nand U6369 (N_6369,N_5779,N_5633);
nor U6370 (N_6370,N_5558,N_5516);
nand U6371 (N_6371,N_5606,N_5613);
or U6372 (N_6372,N_5514,N_5893);
and U6373 (N_6373,N_5884,N_5854);
and U6374 (N_6374,N_5589,N_5542);
xor U6375 (N_6375,N_5877,N_5624);
nand U6376 (N_6376,N_5788,N_5871);
and U6377 (N_6377,N_5831,N_5953);
or U6378 (N_6378,N_5892,N_5775);
or U6379 (N_6379,N_5998,N_5854);
xor U6380 (N_6380,N_5780,N_5545);
nand U6381 (N_6381,N_5639,N_5647);
or U6382 (N_6382,N_5500,N_5765);
or U6383 (N_6383,N_5963,N_5928);
and U6384 (N_6384,N_5757,N_5819);
nand U6385 (N_6385,N_5722,N_5548);
nand U6386 (N_6386,N_5511,N_5942);
xor U6387 (N_6387,N_5927,N_5860);
xnor U6388 (N_6388,N_5805,N_5786);
xnor U6389 (N_6389,N_5955,N_5772);
nand U6390 (N_6390,N_5998,N_5609);
and U6391 (N_6391,N_5545,N_5823);
or U6392 (N_6392,N_5873,N_5650);
xor U6393 (N_6393,N_5726,N_5785);
xor U6394 (N_6394,N_5856,N_5532);
nand U6395 (N_6395,N_5650,N_5522);
nor U6396 (N_6396,N_5694,N_5871);
nand U6397 (N_6397,N_5617,N_5965);
nor U6398 (N_6398,N_5933,N_5800);
nor U6399 (N_6399,N_5725,N_5847);
nor U6400 (N_6400,N_5810,N_5753);
nor U6401 (N_6401,N_5683,N_5596);
nor U6402 (N_6402,N_5500,N_5589);
nand U6403 (N_6403,N_5775,N_5604);
nand U6404 (N_6404,N_5760,N_5972);
nor U6405 (N_6405,N_5900,N_5901);
and U6406 (N_6406,N_5532,N_5751);
and U6407 (N_6407,N_5910,N_5849);
or U6408 (N_6408,N_5797,N_5515);
nand U6409 (N_6409,N_5705,N_5718);
nor U6410 (N_6410,N_5824,N_5782);
and U6411 (N_6411,N_5954,N_5806);
nand U6412 (N_6412,N_5919,N_5690);
xor U6413 (N_6413,N_5852,N_5948);
xnor U6414 (N_6414,N_5883,N_5568);
or U6415 (N_6415,N_5756,N_5548);
xor U6416 (N_6416,N_5692,N_5782);
or U6417 (N_6417,N_5687,N_5597);
nor U6418 (N_6418,N_5794,N_5971);
nand U6419 (N_6419,N_5976,N_5663);
nand U6420 (N_6420,N_5715,N_5989);
or U6421 (N_6421,N_5559,N_5575);
or U6422 (N_6422,N_5663,N_5932);
xnor U6423 (N_6423,N_5756,N_5916);
and U6424 (N_6424,N_5737,N_5784);
xor U6425 (N_6425,N_5793,N_5913);
nand U6426 (N_6426,N_5958,N_5749);
nand U6427 (N_6427,N_5999,N_5945);
or U6428 (N_6428,N_5880,N_5881);
nor U6429 (N_6429,N_5620,N_5748);
nor U6430 (N_6430,N_5811,N_5534);
or U6431 (N_6431,N_5878,N_5703);
or U6432 (N_6432,N_5559,N_5693);
nand U6433 (N_6433,N_5719,N_5577);
or U6434 (N_6434,N_5642,N_5716);
nand U6435 (N_6435,N_5627,N_5839);
nor U6436 (N_6436,N_5642,N_5696);
and U6437 (N_6437,N_5819,N_5525);
nor U6438 (N_6438,N_5543,N_5951);
xor U6439 (N_6439,N_5848,N_5799);
nand U6440 (N_6440,N_5748,N_5686);
and U6441 (N_6441,N_5746,N_5824);
and U6442 (N_6442,N_5961,N_5738);
and U6443 (N_6443,N_5991,N_5628);
or U6444 (N_6444,N_5819,N_5761);
and U6445 (N_6445,N_5936,N_5909);
and U6446 (N_6446,N_5841,N_5906);
or U6447 (N_6447,N_5877,N_5575);
nand U6448 (N_6448,N_5712,N_5528);
xor U6449 (N_6449,N_5914,N_5614);
nand U6450 (N_6450,N_5617,N_5917);
nor U6451 (N_6451,N_5924,N_5836);
nor U6452 (N_6452,N_5702,N_5527);
or U6453 (N_6453,N_5743,N_5723);
or U6454 (N_6454,N_5869,N_5688);
nor U6455 (N_6455,N_5693,N_5909);
xnor U6456 (N_6456,N_5530,N_5563);
and U6457 (N_6457,N_5512,N_5695);
or U6458 (N_6458,N_5618,N_5764);
nor U6459 (N_6459,N_5522,N_5600);
nor U6460 (N_6460,N_5746,N_5835);
or U6461 (N_6461,N_5777,N_5760);
xnor U6462 (N_6462,N_5541,N_5917);
or U6463 (N_6463,N_5713,N_5599);
and U6464 (N_6464,N_5593,N_5723);
xnor U6465 (N_6465,N_5907,N_5749);
nand U6466 (N_6466,N_5991,N_5901);
nand U6467 (N_6467,N_5799,N_5890);
xor U6468 (N_6468,N_5854,N_5605);
nand U6469 (N_6469,N_5734,N_5526);
or U6470 (N_6470,N_5596,N_5711);
and U6471 (N_6471,N_5554,N_5659);
nand U6472 (N_6472,N_5615,N_5695);
xor U6473 (N_6473,N_5816,N_5927);
xor U6474 (N_6474,N_5817,N_5522);
and U6475 (N_6475,N_5895,N_5744);
or U6476 (N_6476,N_5503,N_5920);
and U6477 (N_6477,N_5515,N_5738);
nor U6478 (N_6478,N_5694,N_5818);
nand U6479 (N_6479,N_5672,N_5754);
or U6480 (N_6480,N_5965,N_5628);
nor U6481 (N_6481,N_5668,N_5531);
nor U6482 (N_6482,N_5559,N_5773);
or U6483 (N_6483,N_5662,N_5967);
xor U6484 (N_6484,N_5752,N_5780);
or U6485 (N_6485,N_5621,N_5856);
nand U6486 (N_6486,N_5539,N_5826);
and U6487 (N_6487,N_5523,N_5851);
and U6488 (N_6488,N_5500,N_5671);
nand U6489 (N_6489,N_5743,N_5860);
xor U6490 (N_6490,N_5587,N_5521);
and U6491 (N_6491,N_5650,N_5929);
xnor U6492 (N_6492,N_5649,N_5973);
xnor U6493 (N_6493,N_5816,N_5669);
and U6494 (N_6494,N_5694,N_5785);
nand U6495 (N_6495,N_5980,N_5704);
and U6496 (N_6496,N_5615,N_5840);
xor U6497 (N_6497,N_5759,N_5838);
xnor U6498 (N_6498,N_5672,N_5858);
xor U6499 (N_6499,N_5594,N_5646);
and U6500 (N_6500,N_6129,N_6297);
xor U6501 (N_6501,N_6212,N_6101);
nand U6502 (N_6502,N_6321,N_6193);
nand U6503 (N_6503,N_6493,N_6279);
nand U6504 (N_6504,N_6487,N_6417);
nor U6505 (N_6505,N_6220,N_6026);
xnor U6506 (N_6506,N_6239,N_6082);
or U6507 (N_6507,N_6485,N_6073);
nand U6508 (N_6508,N_6430,N_6243);
xnor U6509 (N_6509,N_6259,N_6453);
nand U6510 (N_6510,N_6048,N_6252);
and U6511 (N_6511,N_6363,N_6158);
xor U6512 (N_6512,N_6123,N_6071);
xor U6513 (N_6513,N_6164,N_6432);
xor U6514 (N_6514,N_6383,N_6402);
and U6515 (N_6515,N_6157,N_6401);
or U6516 (N_6516,N_6240,N_6277);
or U6517 (N_6517,N_6392,N_6037);
nand U6518 (N_6518,N_6056,N_6325);
and U6519 (N_6519,N_6312,N_6358);
or U6520 (N_6520,N_6246,N_6078);
nand U6521 (N_6521,N_6200,N_6340);
or U6522 (N_6522,N_6378,N_6084);
nor U6523 (N_6523,N_6475,N_6036);
or U6524 (N_6524,N_6008,N_6142);
or U6525 (N_6525,N_6218,N_6127);
nand U6526 (N_6526,N_6155,N_6159);
xor U6527 (N_6527,N_6199,N_6107);
xnor U6528 (N_6528,N_6484,N_6054);
nand U6529 (N_6529,N_6172,N_6278);
nand U6530 (N_6530,N_6264,N_6244);
and U6531 (N_6531,N_6188,N_6347);
xnor U6532 (N_6532,N_6028,N_6290);
nor U6533 (N_6533,N_6115,N_6119);
and U6534 (N_6534,N_6330,N_6310);
xor U6535 (N_6535,N_6085,N_6125);
nor U6536 (N_6536,N_6474,N_6272);
or U6537 (N_6537,N_6300,N_6380);
and U6538 (N_6538,N_6138,N_6012);
nor U6539 (N_6539,N_6455,N_6447);
nand U6540 (N_6540,N_6260,N_6134);
xor U6541 (N_6541,N_6361,N_6480);
nand U6542 (N_6542,N_6019,N_6496);
nor U6543 (N_6543,N_6209,N_6150);
or U6544 (N_6544,N_6110,N_6191);
and U6545 (N_6545,N_6175,N_6092);
nor U6546 (N_6546,N_6359,N_6268);
nor U6547 (N_6547,N_6385,N_6441);
nor U6548 (N_6548,N_6370,N_6444);
xnor U6549 (N_6549,N_6381,N_6439);
and U6550 (N_6550,N_6041,N_6492);
nand U6551 (N_6551,N_6423,N_6215);
or U6552 (N_6552,N_6117,N_6059);
nor U6553 (N_6553,N_6067,N_6341);
xor U6554 (N_6554,N_6372,N_6466);
xor U6555 (N_6555,N_6324,N_6214);
nand U6556 (N_6556,N_6418,N_6154);
nor U6557 (N_6557,N_6309,N_6088);
nand U6558 (N_6558,N_6346,N_6050);
nand U6559 (N_6559,N_6433,N_6343);
or U6560 (N_6560,N_6288,N_6305);
and U6561 (N_6561,N_6186,N_6201);
or U6562 (N_6562,N_6436,N_6491);
nor U6563 (N_6563,N_6398,N_6327);
nand U6564 (N_6564,N_6425,N_6420);
nand U6565 (N_6565,N_6061,N_6038);
nand U6566 (N_6566,N_6494,N_6421);
xnor U6567 (N_6567,N_6454,N_6431);
nor U6568 (N_6568,N_6018,N_6499);
xor U6569 (N_6569,N_6224,N_6292);
nand U6570 (N_6570,N_6234,N_6409);
or U6571 (N_6571,N_6146,N_6250);
nand U6572 (N_6572,N_6002,N_6195);
and U6573 (N_6573,N_6253,N_6202);
nor U6574 (N_6574,N_6350,N_6000);
and U6575 (N_6575,N_6360,N_6263);
nand U6576 (N_6576,N_6072,N_6400);
xor U6577 (N_6577,N_6130,N_6091);
nor U6578 (N_6578,N_6017,N_6062);
xor U6579 (N_6579,N_6303,N_6351);
nor U6580 (N_6580,N_6304,N_6096);
nor U6581 (N_6581,N_6083,N_6483);
xnor U6582 (N_6582,N_6355,N_6404);
or U6583 (N_6583,N_6233,N_6414);
nand U6584 (N_6584,N_6294,N_6098);
xor U6585 (N_6585,N_6276,N_6226);
nand U6586 (N_6586,N_6367,N_6094);
and U6587 (N_6587,N_6395,N_6034);
or U6588 (N_6588,N_6261,N_6319);
and U6589 (N_6589,N_6365,N_6227);
and U6590 (N_6590,N_6255,N_6296);
nor U6591 (N_6591,N_6316,N_6030);
nor U6592 (N_6592,N_6489,N_6176);
nor U6593 (N_6593,N_6289,N_6055);
and U6594 (N_6594,N_6419,N_6333);
and U6595 (N_6595,N_6205,N_6219);
or U6596 (N_6596,N_6497,N_6063);
or U6597 (N_6597,N_6032,N_6011);
xnor U6598 (N_6598,N_6147,N_6258);
or U6599 (N_6599,N_6122,N_6245);
xor U6600 (N_6600,N_6165,N_6238);
nand U6601 (N_6601,N_6376,N_6043);
nand U6602 (N_6602,N_6407,N_6352);
nand U6603 (N_6603,N_6462,N_6449);
and U6604 (N_6604,N_6095,N_6016);
or U6605 (N_6605,N_6076,N_6477);
or U6606 (N_6606,N_6197,N_6135);
or U6607 (N_6607,N_6457,N_6223);
or U6608 (N_6608,N_6314,N_6044);
and U6609 (N_6609,N_6208,N_6295);
xor U6610 (N_6610,N_6459,N_6058);
and U6611 (N_6611,N_6266,N_6174);
xnor U6612 (N_6612,N_6178,N_6473);
xnor U6613 (N_6613,N_6315,N_6232);
and U6614 (N_6614,N_6006,N_6302);
or U6615 (N_6615,N_6495,N_6410);
or U6616 (N_6616,N_6120,N_6105);
xnor U6617 (N_6617,N_6111,N_6068);
and U6618 (N_6618,N_6481,N_6039);
nand U6619 (N_6619,N_6133,N_6229);
xnor U6620 (N_6620,N_6162,N_6015);
nor U6621 (N_6621,N_6356,N_6131);
nor U6622 (N_6622,N_6198,N_6031);
xor U6623 (N_6623,N_6136,N_6060);
and U6624 (N_6624,N_6116,N_6438);
xnor U6625 (N_6625,N_6113,N_6287);
xor U6626 (N_6626,N_6013,N_6090);
nand U6627 (N_6627,N_6241,N_6160);
and U6628 (N_6628,N_6328,N_6149);
nand U6629 (N_6629,N_6190,N_6332);
nand U6630 (N_6630,N_6153,N_6403);
nand U6631 (N_6631,N_6336,N_6445);
nor U6632 (N_6632,N_6440,N_6464);
xnor U6633 (N_6633,N_6128,N_6326);
xnor U6634 (N_6634,N_6033,N_6099);
and U6635 (N_6635,N_6482,N_6397);
xnor U6636 (N_6636,N_6235,N_6374);
and U6637 (N_6637,N_6311,N_6124);
and U6638 (N_6638,N_6331,N_6424);
and U6639 (N_6639,N_6348,N_6411);
and U6640 (N_6640,N_6075,N_6163);
xnor U6641 (N_6641,N_6298,N_6161);
and U6642 (N_6642,N_6422,N_6339);
nand U6643 (N_6643,N_6269,N_6051);
xnor U6644 (N_6644,N_6443,N_6437);
nand U6645 (N_6645,N_6353,N_6387);
xnor U6646 (N_6646,N_6184,N_6283);
nor U6647 (N_6647,N_6318,N_6181);
nand U6648 (N_6648,N_6470,N_6183);
nor U6649 (N_6649,N_6435,N_6046);
nand U6650 (N_6650,N_6427,N_6415);
nand U6651 (N_6651,N_6396,N_6104);
or U6652 (N_6652,N_6114,N_6079);
and U6653 (N_6653,N_6069,N_6247);
nor U6654 (N_6654,N_6179,N_6313);
or U6655 (N_6655,N_6393,N_6384);
nor U6656 (N_6656,N_6293,N_6177);
nand U6657 (N_6657,N_6299,N_6486);
xor U6658 (N_6658,N_6320,N_6121);
nand U6659 (N_6659,N_6335,N_6093);
or U6660 (N_6660,N_6004,N_6057);
nand U6661 (N_6661,N_6389,N_6369);
nor U6662 (N_6662,N_6074,N_6362);
nand U6663 (N_6663,N_6007,N_6140);
and U6664 (N_6664,N_6003,N_6132);
or U6665 (N_6665,N_6498,N_6463);
xor U6666 (N_6666,N_6391,N_6109);
xnor U6667 (N_6667,N_6284,N_6364);
xnor U6668 (N_6668,N_6009,N_6025);
and U6669 (N_6669,N_6210,N_6373);
nand U6670 (N_6670,N_6194,N_6211);
nand U6671 (N_6671,N_6461,N_6458);
nor U6672 (N_6672,N_6413,N_6189);
nand U6673 (N_6673,N_6040,N_6257);
xnor U6674 (N_6674,N_6468,N_6027);
or U6675 (N_6675,N_6467,N_6322);
nand U6676 (N_6676,N_6291,N_6274);
xor U6677 (N_6677,N_6399,N_6452);
nor U6678 (N_6678,N_6187,N_6213);
or U6679 (N_6679,N_6426,N_6080);
xor U6680 (N_6680,N_6196,N_6102);
xnor U6681 (N_6681,N_6371,N_6171);
and U6682 (N_6682,N_6014,N_6029);
and U6683 (N_6683,N_6236,N_6379);
and U6684 (N_6684,N_6286,N_6377);
and U6685 (N_6685,N_6045,N_6180);
and U6686 (N_6686,N_6023,N_6207);
xnor U6687 (N_6687,N_6273,N_6206);
xnor U6688 (N_6688,N_6216,N_6262);
or U6689 (N_6689,N_6329,N_6428);
nor U6690 (N_6690,N_6412,N_6170);
xnor U6691 (N_6691,N_6275,N_6388);
xor U6692 (N_6692,N_6448,N_6471);
or U6693 (N_6693,N_6167,N_6256);
or U6694 (N_6694,N_6143,N_6429);
or U6695 (N_6695,N_6137,N_6228);
nor U6696 (N_6696,N_6070,N_6490);
xor U6697 (N_6697,N_6087,N_6386);
nor U6698 (N_6698,N_6456,N_6222);
nand U6699 (N_6699,N_6203,N_6173);
xnor U6700 (N_6700,N_6152,N_6145);
or U6701 (N_6701,N_6156,N_6368);
or U6702 (N_6702,N_6406,N_6345);
nand U6703 (N_6703,N_6024,N_6271);
nand U6704 (N_6704,N_6408,N_6465);
nor U6705 (N_6705,N_6103,N_6344);
and U6706 (N_6706,N_6066,N_6390);
or U6707 (N_6707,N_6020,N_6141);
nand U6708 (N_6708,N_6488,N_6281);
xnor U6709 (N_6709,N_6469,N_6342);
xnor U6710 (N_6710,N_6139,N_6478);
nor U6711 (N_6711,N_6118,N_6151);
nor U6712 (N_6712,N_6001,N_6450);
nand U6713 (N_6713,N_6416,N_6472);
or U6714 (N_6714,N_6230,N_6254);
xnor U6715 (N_6715,N_6451,N_6285);
nand U6716 (N_6716,N_6077,N_6357);
and U6717 (N_6717,N_6221,N_6112);
and U6718 (N_6718,N_6394,N_6168);
and U6719 (N_6719,N_6185,N_6021);
or U6720 (N_6720,N_6405,N_6144);
or U6721 (N_6721,N_6064,N_6005);
nand U6722 (N_6722,N_6204,N_6089);
or U6723 (N_6723,N_6334,N_6349);
nand U6724 (N_6724,N_6042,N_6446);
or U6725 (N_6725,N_6047,N_6337);
xnor U6726 (N_6726,N_6280,N_6265);
xor U6727 (N_6727,N_6479,N_6086);
and U6728 (N_6728,N_6049,N_6251);
nand U6729 (N_6729,N_6081,N_6053);
or U6730 (N_6730,N_6267,N_6192);
nor U6731 (N_6731,N_6307,N_6231);
or U6732 (N_6732,N_6148,N_6052);
nand U6733 (N_6733,N_6382,N_6354);
or U6734 (N_6734,N_6182,N_6225);
and U6735 (N_6735,N_6442,N_6169);
nand U6736 (N_6736,N_6323,N_6126);
and U6737 (N_6737,N_6476,N_6306);
nand U6738 (N_6738,N_6106,N_6248);
or U6739 (N_6739,N_6282,N_6237);
or U6740 (N_6740,N_6010,N_6317);
xnor U6741 (N_6741,N_6366,N_6217);
xor U6742 (N_6742,N_6022,N_6166);
nor U6743 (N_6743,N_6460,N_6270);
and U6744 (N_6744,N_6249,N_6035);
nor U6745 (N_6745,N_6375,N_6338);
nor U6746 (N_6746,N_6308,N_6108);
nor U6747 (N_6747,N_6065,N_6100);
and U6748 (N_6748,N_6301,N_6434);
or U6749 (N_6749,N_6097,N_6242);
nand U6750 (N_6750,N_6256,N_6459);
nor U6751 (N_6751,N_6325,N_6049);
nand U6752 (N_6752,N_6261,N_6100);
nor U6753 (N_6753,N_6195,N_6324);
xor U6754 (N_6754,N_6207,N_6162);
nand U6755 (N_6755,N_6008,N_6477);
and U6756 (N_6756,N_6283,N_6451);
and U6757 (N_6757,N_6310,N_6392);
nand U6758 (N_6758,N_6434,N_6273);
xnor U6759 (N_6759,N_6282,N_6214);
and U6760 (N_6760,N_6195,N_6223);
nand U6761 (N_6761,N_6341,N_6362);
nand U6762 (N_6762,N_6077,N_6150);
xor U6763 (N_6763,N_6004,N_6197);
xor U6764 (N_6764,N_6413,N_6053);
or U6765 (N_6765,N_6014,N_6203);
nor U6766 (N_6766,N_6001,N_6174);
nand U6767 (N_6767,N_6106,N_6168);
and U6768 (N_6768,N_6195,N_6268);
and U6769 (N_6769,N_6462,N_6362);
or U6770 (N_6770,N_6495,N_6254);
or U6771 (N_6771,N_6037,N_6046);
and U6772 (N_6772,N_6481,N_6131);
nor U6773 (N_6773,N_6495,N_6117);
and U6774 (N_6774,N_6318,N_6140);
and U6775 (N_6775,N_6249,N_6258);
or U6776 (N_6776,N_6319,N_6291);
nor U6777 (N_6777,N_6086,N_6199);
or U6778 (N_6778,N_6093,N_6279);
or U6779 (N_6779,N_6124,N_6165);
or U6780 (N_6780,N_6496,N_6474);
or U6781 (N_6781,N_6478,N_6026);
nand U6782 (N_6782,N_6033,N_6475);
and U6783 (N_6783,N_6179,N_6299);
and U6784 (N_6784,N_6269,N_6271);
nor U6785 (N_6785,N_6438,N_6071);
and U6786 (N_6786,N_6223,N_6336);
xor U6787 (N_6787,N_6238,N_6042);
nor U6788 (N_6788,N_6402,N_6149);
or U6789 (N_6789,N_6488,N_6124);
nor U6790 (N_6790,N_6362,N_6436);
xnor U6791 (N_6791,N_6038,N_6170);
nand U6792 (N_6792,N_6444,N_6214);
nand U6793 (N_6793,N_6045,N_6138);
nand U6794 (N_6794,N_6104,N_6230);
and U6795 (N_6795,N_6204,N_6262);
xnor U6796 (N_6796,N_6335,N_6127);
and U6797 (N_6797,N_6286,N_6445);
xnor U6798 (N_6798,N_6018,N_6445);
xnor U6799 (N_6799,N_6010,N_6345);
and U6800 (N_6800,N_6009,N_6234);
and U6801 (N_6801,N_6344,N_6260);
nor U6802 (N_6802,N_6427,N_6364);
nand U6803 (N_6803,N_6420,N_6166);
and U6804 (N_6804,N_6417,N_6372);
xnor U6805 (N_6805,N_6411,N_6187);
nand U6806 (N_6806,N_6275,N_6474);
or U6807 (N_6807,N_6355,N_6186);
and U6808 (N_6808,N_6475,N_6258);
or U6809 (N_6809,N_6342,N_6165);
or U6810 (N_6810,N_6010,N_6198);
nor U6811 (N_6811,N_6050,N_6465);
and U6812 (N_6812,N_6119,N_6145);
nor U6813 (N_6813,N_6253,N_6340);
xnor U6814 (N_6814,N_6211,N_6475);
and U6815 (N_6815,N_6153,N_6013);
nand U6816 (N_6816,N_6224,N_6432);
xnor U6817 (N_6817,N_6276,N_6092);
xor U6818 (N_6818,N_6417,N_6412);
xor U6819 (N_6819,N_6036,N_6470);
xor U6820 (N_6820,N_6324,N_6102);
or U6821 (N_6821,N_6495,N_6022);
xnor U6822 (N_6822,N_6096,N_6171);
nand U6823 (N_6823,N_6298,N_6281);
and U6824 (N_6824,N_6218,N_6371);
and U6825 (N_6825,N_6483,N_6427);
nand U6826 (N_6826,N_6170,N_6091);
xnor U6827 (N_6827,N_6424,N_6394);
or U6828 (N_6828,N_6282,N_6488);
nand U6829 (N_6829,N_6055,N_6314);
or U6830 (N_6830,N_6124,N_6475);
and U6831 (N_6831,N_6060,N_6020);
xnor U6832 (N_6832,N_6286,N_6289);
nor U6833 (N_6833,N_6222,N_6338);
and U6834 (N_6834,N_6180,N_6275);
or U6835 (N_6835,N_6014,N_6230);
and U6836 (N_6836,N_6383,N_6421);
xnor U6837 (N_6837,N_6381,N_6174);
and U6838 (N_6838,N_6163,N_6171);
xnor U6839 (N_6839,N_6317,N_6006);
nand U6840 (N_6840,N_6082,N_6262);
or U6841 (N_6841,N_6270,N_6085);
and U6842 (N_6842,N_6204,N_6172);
nand U6843 (N_6843,N_6278,N_6318);
and U6844 (N_6844,N_6329,N_6019);
and U6845 (N_6845,N_6438,N_6461);
or U6846 (N_6846,N_6464,N_6163);
or U6847 (N_6847,N_6248,N_6490);
nor U6848 (N_6848,N_6297,N_6092);
nand U6849 (N_6849,N_6124,N_6006);
and U6850 (N_6850,N_6299,N_6249);
or U6851 (N_6851,N_6407,N_6270);
nor U6852 (N_6852,N_6333,N_6096);
nand U6853 (N_6853,N_6310,N_6064);
xor U6854 (N_6854,N_6429,N_6129);
xor U6855 (N_6855,N_6406,N_6440);
or U6856 (N_6856,N_6129,N_6092);
xor U6857 (N_6857,N_6287,N_6144);
or U6858 (N_6858,N_6196,N_6439);
nor U6859 (N_6859,N_6062,N_6484);
and U6860 (N_6860,N_6328,N_6004);
nand U6861 (N_6861,N_6324,N_6403);
nand U6862 (N_6862,N_6485,N_6151);
xnor U6863 (N_6863,N_6259,N_6125);
xnor U6864 (N_6864,N_6005,N_6205);
xnor U6865 (N_6865,N_6332,N_6411);
and U6866 (N_6866,N_6199,N_6451);
and U6867 (N_6867,N_6238,N_6163);
nor U6868 (N_6868,N_6112,N_6416);
and U6869 (N_6869,N_6193,N_6448);
nor U6870 (N_6870,N_6076,N_6128);
xor U6871 (N_6871,N_6039,N_6279);
xor U6872 (N_6872,N_6274,N_6024);
nor U6873 (N_6873,N_6387,N_6368);
and U6874 (N_6874,N_6412,N_6199);
xnor U6875 (N_6875,N_6174,N_6483);
nor U6876 (N_6876,N_6077,N_6456);
nand U6877 (N_6877,N_6065,N_6172);
and U6878 (N_6878,N_6108,N_6336);
or U6879 (N_6879,N_6005,N_6187);
and U6880 (N_6880,N_6034,N_6067);
nand U6881 (N_6881,N_6075,N_6148);
nand U6882 (N_6882,N_6356,N_6251);
xnor U6883 (N_6883,N_6292,N_6002);
xnor U6884 (N_6884,N_6030,N_6167);
and U6885 (N_6885,N_6149,N_6354);
nand U6886 (N_6886,N_6110,N_6195);
nand U6887 (N_6887,N_6311,N_6308);
nand U6888 (N_6888,N_6062,N_6312);
xnor U6889 (N_6889,N_6144,N_6314);
nor U6890 (N_6890,N_6489,N_6359);
xnor U6891 (N_6891,N_6344,N_6206);
xor U6892 (N_6892,N_6379,N_6084);
xnor U6893 (N_6893,N_6354,N_6405);
and U6894 (N_6894,N_6358,N_6258);
xor U6895 (N_6895,N_6306,N_6340);
nor U6896 (N_6896,N_6201,N_6077);
nand U6897 (N_6897,N_6204,N_6373);
or U6898 (N_6898,N_6442,N_6004);
nand U6899 (N_6899,N_6120,N_6204);
xor U6900 (N_6900,N_6315,N_6342);
nor U6901 (N_6901,N_6288,N_6027);
or U6902 (N_6902,N_6258,N_6107);
nand U6903 (N_6903,N_6098,N_6420);
xor U6904 (N_6904,N_6137,N_6020);
nand U6905 (N_6905,N_6145,N_6416);
or U6906 (N_6906,N_6015,N_6290);
nor U6907 (N_6907,N_6197,N_6289);
and U6908 (N_6908,N_6359,N_6216);
or U6909 (N_6909,N_6450,N_6068);
nor U6910 (N_6910,N_6046,N_6388);
xor U6911 (N_6911,N_6178,N_6138);
nand U6912 (N_6912,N_6411,N_6134);
nand U6913 (N_6913,N_6415,N_6333);
nand U6914 (N_6914,N_6062,N_6133);
and U6915 (N_6915,N_6296,N_6305);
nand U6916 (N_6916,N_6254,N_6000);
nand U6917 (N_6917,N_6252,N_6457);
or U6918 (N_6918,N_6280,N_6194);
and U6919 (N_6919,N_6094,N_6373);
nand U6920 (N_6920,N_6000,N_6337);
or U6921 (N_6921,N_6225,N_6479);
nand U6922 (N_6922,N_6012,N_6023);
xnor U6923 (N_6923,N_6402,N_6411);
or U6924 (N_6924,N_6398,N_6184);
and U6925 (N_6925,N_6442,N_6159);
nand U6926 (N_6926,N_6122,N_6102);
nand U6927 (N_6927,N_6490,N_6117);
nand U6928 (N_6928,N_6314,N_6240);
and U6929 (N_6929,N_6454,N_6089);
nand U6930 (N_6930,N_6452,N_6412);
nand U6931 (N_6931,N_6291,N_6246);
or U6932 (N_6932,N_6328,N_6107);
xnor U6933 (N_6933,N_6433,N_6363);
or U6934 (N_6934,N_6227,N_6393);
and U6935 (N_6935,N_6353,N_6195);
nor U6936 (N_6936,N_6037,N_6397);
xnor U6937 (N_6937,N_6402,N_6365);
and U6938 (N_6938,N_6128,N_6107);
xnor U6939 (N_6939,N_6361,N_6371);
and U6940 (N_6940,N_6211,N_6390);
and U6941 (N_6941,N_6185,N_6305);
or U6942 (N_6942,N_6310,N_6168);
nor U6943 (N_6943,N_6113,N_6098);
nor U6944 (N_6944,N_6489,N_6258);
or U6945 (N_6945,N_6213,N_6343);
nand U6946 (N_6946,N_6000,N_6351);
nor U6947 (N_6947,N_6071,N_6128);
xnor U6948 (N_6948,N_6425,N_6423);
or U6949 (N_6949,N_6123,N_6095);
xnor U6950 (N_6950,N_6386,N_6411);
nor U6951 (N_6951,N_6457,N_6461);
xnor U6952 (N_6952,N_6224,N_6477);
nand U6953 (N_6953,N_6191,N_6427);
nand U6954 (N_6954,N_6012,N_6318);
nor U6955 (N_6955,N_6491,N_6256);
nand U6956 (N_6956,N_6417,N_6303);
nand U6957 (N_6957,N_6275,N_6368);
nor U6958 (N_6958,N_6406,N_6439);
and U6959 (N_6959,N_6133,N_6466);
xnor U6960 (N_6960,N_6243,N_6144);
and U6961 (N_6961,N_6236,N_6461);
xnor U6962 (N_6962,N_6005,N_6173);
nand U6963 (N_6963,N_6291,N_6021);
and U6964 (N_6964,N_6238,N_6098);
nand U6965 (N_6965,N_6463,N_6209);
or U6966 (N_6966,N_6049,N_6168);
nor U6967 (N_6967,N_6236,N_6149);
xnor U6968 (N_6968,N_6210,N_6484);
nand U6969 (N_6969,N_6439,N_6024);
xor U6970 (N_6970,N_6100,N_6271);
nand U6971 (N_6971,N_6133,N_6249);
nand U6972 (N_6972,N_6394,N_6277);
and U6973 (N_6973,N_6103,N_6273);
and U6974 (N_6974,N_6031,N_6106);
xnor U6975 (N_6975,N_6119,N_6335);
xnor U6976 (N_6976,N_6325,N_6001);
and U6977 (N_6977,N_6455,N_6254);
or U6978 (N_6978,N_6334,N_6301);
nand U6979 (N_6979,N_6407,N_6320);
and U6980 (N_6980,N_6321,N_6235);
xnor U6981 (N_6981,N_6232,N_6199);
and U6982 (N_6982,N_6158,N_6438);
nand U6983 (N_6983,N_6347,N_6254);
nand U6984 (N_6984,N_6067,N_6227);
nand U6985 (N_6985,N_6053,N_6409);
nand U6986 (N_6986,N_6041,N_6355);
and U6987 (N_6987,N_6105,N_6412);
and U6988 (N_6988,N_6220,N_6322);
or U6989 (N_6989,N_6048,N_6184);
or U6990 (N_6990,N_6416,N_6277);
xor U6991 (N_6991,N_6244,N_6250);
xnor U6992 (N_6992,N_6453,N_6160);
xor U6993 (N_6993,N_6051,N_6169);
and U6994 (N_6994,N_6113,N_6425);
nand U6995 (N_6995,N_6415,N_6017);
nor U6996 (N_6996,N_6032,N_6325);
nand U6997 (N_6997,N_6187,N_6359);
or U6998 (N_6998,N_6223,N_6094);
or U6999 (N_6999,N_6089,N_6179);
nand U7000 (N_7000,N_6579,N_6650);
and U7001 (N_7001,N_6715,N_6874);
nor U7002 (N_7002,N_6887,N_6990);
nor U7003 (N_7003,N_6672,N_6625);
and U7004 (N_7004,N_6534,N_6519);
nand U7005 (N_7005,N_6555,N_6881);
or U7006 (N_7006,N_6586,N_6687);
nor U7007 (N_7007,N_6578,N_6627);
nand U7008 (N_7008,N_6820,N_6802);
and U7009 (N_7009,N_6969,N_6637);
and U7010 (N_7010,N_6686,N_6634);
nand U7011 (N_7011,N_6930,N_6681);
and U7012 (N_7012,N_6948,N_6877);
nand U7013 (N_7013,N_6795,N_6710);
nand U7014 (N_7014,N_6846,N_6953);
and U7015 (N_7015,N_6528,N_6538);
or U7016 (N_7016,N_6847,N_6602);
and U7017 (N_7017,N_6886,N_6726);
xor U7018 (N_7018,N_6956,N_6678);
and U7019 (N_7019,N_6585,N_6805);
xor U7020 (N_7020,N_6598,N_6774);
and U7021 (N_7021,N_6622,N_6771);
or U7022 (N_7022,N_6574,N_6888);
xor U7023 (N_7023,N_6611,N_6700);
nor U7024 (N_7024,N_6740,N_6934);
nand U7025 (N_7025,N_6746,N_6540);
nand U7026 (N_7026,N_6502,N_6850);
nor U7027 (N_7027,N_6989,N_6954);
xor U7028 (N_7028,N_6531,N_6750);
and U7029 (N_7029,N_6520,N_6546);
xnor U7030 (N_7030,N_6568,N_6960);
nor U7031 (N_7031,N_6842,N_6575);
and U7032 (N_7032,N_6809,N_6789);
xnor U7033 (N_7033,N_6524,N_6589);
or U7034 (N_7034,N_6702,N_6709);
nor U7035 (N_7035,N_6849,N_6858);
nand U7036 (N_7036,N_6892,N_6992);
nor U7037 (N_7037,N_6770,N_6659);
xnor U7038 (N_7038,N_6708,N_6747);
xor U7039 (N_7039,N_6984,N_6764);
or U7040 (N_7040,N_6566,N_6572);
and U7041 (N_7041,N_6844,N_6542);
or U7042 (N_7042,N_6517,N_6781);
or U7043 (N_7043,N_6973,N_6861);
nor U7044 (N_7044,N_6644,N_6612);
nor U7045 (N_7045,N_6620,N_6812);
xor U7046 (N_7046,N_6668,N_6558);
and U7047 (N_7047,N_6541,N_6997);
xor U7048 (N_7048,N_6995,N_6936);
nor U7049 (N_7049,N_6565,N_6964);
xor U7050 (N_7050,N_6500,N_6843);
nand U7051 (N_7051,N_6601,N_6868);
xor U7052 (N_7052,N_6706,N_6526);
or U7053 (N_7053,N_6518,N_6514);
nor U7054 (N_7054,N_6823,N_6730);
and U7055 (N_7055,N_6949,N_6641);
nor U7056 (N_7056,N_6825,N_6696);
and U7057 (N_7057,N_6511,N_6752);
and U7058 (N_7058,N_6910,N_6662);
nor U7059 (N_7059,N_6951,N_6894);
nor U7060 (N_7060,N_6667,N_6693);
and U7061 (N_7061,N_6615,N_6926);
and U7062 (N_7062,N_6833,N_6523);
xnor U7063 (N_7063,N_6939,N_6811);
xor U7064 (N_7064,N_6917,N_6688);
or U7065 (N_7065,N_6525,N_6830);
xnor U7066 (N_7066,N_6527,N_6906);
xor U7067 (N_7067,N_6503,N_6559);
nand U7068 (N_7068,N_6855,N_6676);
nor U7069 (N_7069,N_6636,N_6660);
nand U7070 (N_7070,N_6505,N_6506);
xor U7071 (N_7071,N_6535,N_6591);
and U7072 (N_7072,N_6785,N_6790);
or U7073 (N_7073,N_6651,N_6596);
xnor U7074 (N_7074,N_6647,N_6666);
and U7075 (N_7075,N_6670,N_6722);
nand U7076 (N_7076,N_6927,N_6777);
xor U7077 (N_7077,N_6915,N_6985);
and U7078 (N_7078,N_6533,N_6755);
nor U7079 (N_7079,N_6928,N_6691);
nor U7080 (N_7080,N_6779,N_6851);
nor U7081 (N_7081,N_6816,N_6796);
or U7082 (N_7082,N_6929,N_6852);
nor U7083 (N_7083,N_6875,N_6606);
and U7084 (N_7084,N_6878,N_6884);
nand U7085 (N_7085,N_6545,N_6768);
xnor U7086 (N_7086,N_6940,N_6705);
and U7087 (N_7087,N_6616,N_6595);
nor U7088 (N_7088,N_6946,N_6883);
xnor U7089 (N_7089,N_6663,N_6554);
or U7090 (N_7090,N_6610,N_6880);
xor U7091 (N_7091,N_6749,N_6639);
xnor U7092 (N_7092,N_6818,N_6899);
nor U7093 (N_7093,N_6994,N_6902);
xor U7094 (N_7094,N_6854,N_6549);
nor U7095 (N_7095,N_6599,N_6689);
or U7096 (N_7096,N_6724,N_6567);
xnor U7097 (N_7097,N_6557,N_6769);
or U7098 (N_7098,N_6707,N_6813);
xor U7099 (N_7099,N_6808,N_6810);
xnor U7100 (N_7100,N_6941,N_6675);
nor U7101 (N_7101,N_6970,N_6921);
nand U7102 (N_7102,N_6873,N_6773);
xor U7103 (N_7103,N_6890,N_6780);
nand U7104 (N_7104,N_6869,N_6962);
xor U7105 (N_7105,N_6632,N_6698);
xor U7106 (N_7106,N_6801,N_6658);
nor U7107 (N_7107,N_6551,N_6759);
xor U7108 (N_7108,N_6787,N_6590);
nand U7109 (N_7109,N_6573,N_6922);
and U7110 (N_7110,N_6694,N_6835);
nand U7111 (N_7111,N_6584,N_6864);
or U7112 (N_7112,N_6732,N_6501);
nor U7113 (N_7113,N_6553,N_6775);
or U7114 (N_7114,N_6959,N_6966);
xnor U7115 (N_7115,N_6544,N_6794);
nor U7116 (N_7116,N_6588,N_6652);
xor U7117 (N_7117,N_6762,N_6821);
nand U7118 (N_7118,N_6630,N_6640);
or U7119 (N_7119,N_6983,N_6729);
nor U7120 (N_7120,N_6912,N_6547);
or U7121 (N_7121,N_6839,N_6791);
and U7122 (N_7122,N_6581,N_6714);
or U7123 (N_7123,N_6712,N_6560);
and U7124 (N_7124,N_6674,N_6982);
or U7125 (N_7125,N_6998,N_6957);
and U7126 (N_7126,N_6733,N_6626);
and U7127 (N_7127,N_6753,N_6635);
nand U7128 (N_7128,N_6614,N_6720);
nor U7129 (N_7129,N_6745,N_6799);
nand U7130 (N_7130,N_6792,N_6905);
xnor U7131 (N_7131,N_6907,N_6664);
xnor U7132 (N_7132,N_6629,N_6945);
or U7133 (N_7133,N_6655,N_6911);
or U7134 (N_7134,N_6537,N_6761);
xnor U7135 (N_7135,N_6507,N_6695);
and U7136 (N_7136,N_6867,N_6742);
or U7137 (N_7137,N_6692,N_6932);
nand U7138 (N_7138,N_6803,N_6577);
or U7139 (N_7139,N_6600,N_6657);
xor U7140 (N_7140,N_6757,N_6918);
or U7141 (N_7141,N_6829,N_6550);
nand U7142 (N_7142,N_6690,N_6914);
and U7143 (N_7143,N_6786,N_6870);
nand U7144 (N_7144,N_6977,N_6993);
nor U7145 (N_7145,N_6944,N_6530);
and U7146 (N_7146,N_6646,N_6898);
nor U7147 (N_7147,N_6857,N_6815);
nand U7148 (N_7148,N_6580,N_6561);
nor U7149 (N_7149,N_6564,N_6685);
or U7150 (N_7150,N_6879,N_6671);
or U7151 (N_7151,N_6828,N_6570);
nor U7152 (N_7152,N_6807,N_6882);
and U7153 (N_7153,N_6605,N_6607);
or U7154 (N_7154,N_6797,N_6920);
and U7155 (N_7155,N_6721,N_6901);
nor U7156 (N_7156,N_6971,N_6521);
xor U7157 (N_7157,N_6991,N_6885);
nand U7158 (N_7158,N_6582,N_6648);
nand U7159 (N_7159,N_6723,N_6758);
nor U7160 (N_7160,N_6621,N_6738);
nor U7161 (N_7161,N_6856,N_6509);
and U7162 (N_7162,N_6824,N_6571);
nand U7163 (N_7163,N_6832,N_6543);
xnor U7164 (N_7164,N_6716,N_6725);
nor U7165 (N_7165,N_6597,N_6741);
xnor U7166 (N_7166,N_6638,N_6683);
and U7167 (N_7167,N_6961,N_6853);
and U7168 (N_7168,N_6778,N_6516);
nor U7169 (N_7169,N_6748,N_6765);
nand U7170 (N_7170,N_6760,N_6987);
nand U7171 (N_7171,N_6548,N_6996);
and U7172 (N_7172,N_6704,N_6968);
xnor U7173 (N_7173,N_6653,N_6974);
or U7174 (N_7174,N_6587,N_6603);
or U7175 (N_7175,N_6680,N_6699);
and U7176 (N_7176,N_6594,N_6562);
or U7177 (N_7177,N_6831,N_6665);
nor U7178 (N_7178,N_6776,N_6904);
xor U7179 (N_7179,N_6925,N_6931);
or U7180 (N_7180,N_6717,N_6754);
xnor U7181 (N_7181,N_6871,N_6913);
nand U7182 (N_7182,N_6837,N_6952);
or U7183 (N_7183,N_6623,N_6504);
or U7184 (N_7184,N_6814,N_6767);
xor U7185 (N_7185,N_6891,N_6728);
xnor U7186 (N_7186,N_6986,N_6739);
and U7187 (N_7187,N_6624,N_6889);
or U7188 (N_7188,N_6836,N_6645);
xor U7189 (N_7189,N_6903,N_6798);
xor U7190 (N_7190,N_6772,N_6512);
or U7191 (N_7191,N_6522,N_6617);
xor U7192 (N_7192,N_6744,N_6958);
and U7193 (N_7193,N_6919,N_6743);
xor U7194 (N_7194,N_6897,N_6872);
xor U7195 (N_7195,N_6822,N_6859);
xnor U7196 (N_7196,N_6800,N_6876);
xnor U7197 (N_7197,N_6763,N_6563);
xnor U7198 (N_7198,N_6938,N_6510);
nand U7199 (N_7199,N_6701,N_6736);
xor U7200 (N_7200,N_6838,N_6654);
nand U7201 (N_7201,N_6508,N_6916);
and U7202 (N_7202,N_6536,N_6593);
and U7203 (N_7203,N_6592,N_6649);
and U7204 (N_7204,N_6788,N_6988);
or U7205 (N_7205,N_6713,N_6784);
and U7206 (N_7206,N_6737,N_6924);
nor U7207 (N_7207,N_6981,N_6806);
nor U7208 (N_7208,N_6552,N_6999);
and U7209 (N_7209,N_6972,N_6866);
nor U7210 (N_7210,N_6673,N_6735);
or U7211 (N_7211,N_6529,N_6942);
and U7212 (N_7212,N_6845,N_6848);
and U7213 (N_7213,N_6711,N_6677);
nand U7214 (N_7214,N_6978,N_6895);
nor U7215 (N_7215,N_6609,N_6618);
or U7216 (N_7216,N_6513,N_6840);
or U7217 (N_7217,N_6756,N_6819);
and U7218 (N_7218,N_6697,N_6893);
and U7219 (N_7219,N_6863,N_6576);
and U7220 (N_7220,N_6860,N_6682);
or U7221 (N_7221,N_6976,N_6908);
or U7222 (N_7222,N_6804,N_6684);
and U7223 (N_7223,N_6556,N_6975);
nand U7224 (N_7224,N_6631,N_6783);
xor U7225 (N_7225,N_6943,N_6569);
and U7226 (N_7226,N_6619,N_6967);
xor U7227 (N_7227,N_6896,N_6669);
and U7228 (N_7228,N_6642,N_6608);
or U7229 (N_7229,N_6515,N_6656);
nand U7230 (N_7230,N_6633,N_6963);
nor U7231 (N_7231,N_6933,N_6613);
nor U7232 (N_7232,N_6782,N_6909);
nand U7233 (N_7233,N_6583,N_6793);
xnor U7234 (N_7234,N_6539,N_6628);
xnor U7235 (N_7235,N_6734,N_6923);
nor U7236 (N_7236,N_6604,N_6965);
xnor U7237 (N_7237,N_6900,N_6865);
xnor U7238 (N_7238,N_6718,N_6703);
and U7239 (N_7239,N_6862,N_6661);
xor U7240 (N_7240,N_6937,N_6727);
and U7241 (N_7241,N_6980,N_6826);
xor U7242 (N_7242,N_6719,N_6935);
nor U7243 (N_7243,N_6955,N_6643);
and U7244 (N_7244,N_6827,N_6751);
or U7245 (N_7245,N_6532,N_6841);
and U7246 (N_7246,N_6731,N_6834);
nor U7247 (N_7247,N_6679,N_6947);
and U7248 (N_7248,N_6817,N_6766);
or U7249 (N_7249,N_6979,N_6950);
and U7250 (N_7250,N_6857,N_6936);
nor U7251 (N_7251,N_6603,N_6500);
or U7252 (N_7252,N_6562,N_6797);
and U7253 (N_7253,N_6919,N_6778);
or U7254 (N_7254,N_6753,N_6545);
xor U7255 (N_7255,N_6619,N_6646);
nor U7256 (N_7256,N_6729,N_6835);
nor U7257 (N_7257,N_6889,N_6770);
xor U7258 (N_7258,N_6640,N_6744);
and U7259 (N_7259,N_6580,N_6782);
or U7260 (N_7260,N_6974,N_6581);
nand U7261 (N_7261,N_6699,N_6741);
nand U7262 (N_7262,N_6938,N_6635);
and U7263 (N_7263,N_6516,N_6594);
or U7264 (N_7264,N_6922,N_6826);
nand U7265 (N_7265,N_6803,N_6683);
xor U7266 (N_7266,N_6534,N_6550);
or U7267 (N_7267,N_6554,N_6687);
nor U7268 (N_7268,N_6975,N_6527);
nand U7269 (N_7269,N_6971,N_6585);
or U7270 (N_7270,N_6925,N_6956);
nand U7271 (N_7271,N_6879,N_6581);
xor U7272 (N_7272,N_6885,N_6895);
or U7273 (N_7273,N_6661,N_6529);
nand U7274 (N_7274,N_6965,N_6686);
nor U7275 (N_7275,N_6811,N_6878);
nand U7276 (N_7276,N_6784,N_6936);
xnor U7277 (N_7277,N_6638,N_6873);
nand U7278 (N_7278,N_6628,N_6513);
nand U7279 (N_7279,N_6776,N_6936);
xnor U7280 (N_7280,N_6949,N_6922);
nor U7281 (N_7281,N_6864,N_6950);
or U7282 (N_7282,N_6554,N_6916);
and U7283 (N_7283,N_6637,N_6540);
or U7284 (N_7284,N_6758,N_6989);
nor U7285 (N_7285,N_6965,N_6921);
or U7286 (N_7286,N_6870,N_6750);
or U7287 (N_7287,N_6519,N_6569);
xor U7288 (N_7288,N_6885,N_6644);
or U7289 (N_7289,N_6783,N_6674);
xor U7290 (N_7290,N_6798,N_6860);
nand U7291 (N_7291,N_6834,N_6613);
and U7292 (N_7292,N_6630,N_6841);
or U7293 (N_7293,N_6526,N_6695);
or U7294 (N_7294,N_6578,N_6982);
or U7295 (N_7295,N_6952,N_6949);
or U7296 (N_7296,N_6970,N_6999);
xnor U7297 (N_7297,N_6521,N_6694);
nor U7298 (N_7298,N_6830,N_6986);
nor U7299 (N_7299,N_6538,N_6859);
and U7300 (N_7300,N_6605,N_6948);
or U7301 (N_7301,N_6701,N_6855);
nand U7302 (N_7302,N_6989,N_6909);
nor U7303 (N_7303,N_6668,N_6655);
xnor U7304 (N_7304,N_6873,N_6840);
and U7305 (N_7305,N_6917,N_6962);
and U7306 (N_7306,N_6939,N_6713);
nand U7307 (N_7307,N_6966,N_6783);
or U7308 (N_7308,N_6982,N_6508);
nand U7309 (N_7309,N_6844,N_6612);
xor U7310 (N_7310,N_6821,N_6572);
nor U7311 (N_7311,N_6928,N_6986);
or U7312 (N_7312,N_6625,N_6953);
nor U7313 (N_7313,N_6840,N_6797);
or U7314 (N_7314,N_6656,N_6663);
nor U7315 (N_7315,N_6634,N_6545);
nor U7316 (N_7316,N_6836,N_6767);
nor U7317 (N_7317,N_6688,N_6954);
or U7318 (N_7318,N_6960,N_6583);
xor U7319 (N_7319,N_6896,N_6680);
nand U7320 (N_7320,N_6808,N_6689);
nor U7321 (N_7321,N_6786,N_6636);
or U7322 (N_7322,N_6502,N_6555);
nor U7323 (N_7323,N_6987,N_6899);
nor U7324 (N_7324,N_6894,N_6842);
xnor U7325 (N_7325,N_6932,N_6654);
nor U7326 (N_7326,N_6901,N_6849);
nand U7327 (N_7327,N_6520,N_6603);
nor U7328 (N_7328,N_6657,N_6973);
or U7329 (N_7329,N_6839,N_6820);
xor U7330 (N_7330,N_6803,N_6597);
and U7331 (N_7331,N_6537,N_6765);
nand U7332 (N_7332,N_6976,N_6623);
xnor U7333 (N_7333,N_6622,N_6889);
xnor U7334 (N_7334,N_6690,N_6607);
and U7335 (N_7335,N_6911,N_6916);
xor U7336 (N_7336,N_6583,N_6656);
and U7337 (N_7337,N_6939,N_6517);
or U7338 (N_7338,N_6639,N_6742);
or U7339 (N_7339,N_6798,N_6734);
xnor U7340 (N_7340,N_6773,N_6980);
nand U7341 (N_7341,N_6569,N_6609);
and U7342 (N_7342,N_6624,N_6713);
xor U7343 (N_7343,N_6801,N_6710);
nor U7344 (N_7344,N_6946,N_6613);
xor U7345 (N_7345,N_6625,N_6724);
xor U7346 (N_7346,N_6801,N_6725);
nor U7347 (N_7347,N_6796,N_6852);
or U7348 (N_7348,N_6622,N_6890);
nand U7349 (N_7349,N_6597,N_6710);
nand U7350 (N_7350,N_6810,N_6594);
and U7351 (N_7351,N_6782,N_6673);
or U7352 (N_7352,N_6661,N_6826);
xnor U7353 (N_7353,N_6696,N_6794);
nor U7354 (N_7354,N_6999,N_6671);
and U7355 (N_7355,N_6527,N_6552);
nand U7356 (N_7356,N_6986,N_6711);
nor U7357 (N_7357,N_6815,N_6902);
xor U7358 (N_7358,N_6885,N_6512);
or U7359 (N_7359,N_6789,N_6549);
and U7360 (N_7360,N_6916,N_6858);
nand U7361 (N_7361,N_6619,N_6763);
nand U7362 (N_7362,N_6670,N_6690);
xor U7363 (N_7363,N_6571,N_6792);
nand U7364 (N_7364,N_6792,N_6957);
nor U7365 (N_7365,N_6588,N_6518);
nor U7366 (N_7366,N_6543,N_6623);
or U7367 (N_7367,N_6864,N_6592);
or U7368 (N_7368,N_6859,N_6606);
nand U7369 (N_7369,N_6531,N_6867);
nor U7370 (N_7370,N_6768,N_6877);
and U7371 (N_7371,N_6634,N_6566);
or U7372 (N_7372,N_6708,N_6543);
nand U7373 (N_7373,N_6985,N_6550);
or U7374 (N_7374,N_6756,N_6749);
or U7375 (N_7375,N_6676,N_6517);
nor U7376 (N_7376,N_6688,N_6541);
xor U7377 (N_7377,N_6586,N_6965);
xnor U7378 (N_7378,N_6799,N_6893);
nand U7379 (N_7379,N_6849,N_6887);
nor U7380 (N_7380,N_6702,N_6968);
nand U7381 (N_7381,N_6760,N_6501);
and U7382 (N_7382,N_6709,N_6935);
and U7383 (N_7383,N_6613,N_6824);
or U7384 (N_7384,N_6517,N_6649);
nand U7385 (N_7385,N_6705,N_6613);
and U7386 (N_7386,N_6703,N_6859);
nor U7387 (N_7387,N_6635,N_6568);
xnor U7388 (N_7388,N_6695,N_6728);
nor U7389 (N_7389,N_6993,N_6814);
nor U7390 (N_7390,N_6721,N_6688);
or U7391 (N_7391,N_6896,N_6501);
or U7392 (N_7392,N_6919,N_6607);
xnor U7393 (N_7393,N_6750,N_6916);
nor U7394 (N_7394,N_6706,N_6765);
nand U7395 (N_7395,N_6564,N_6681);
nor U7396 (N_7396,N_6702,N_6884);
and U7397 (N_7397,N_6931,N_6848);
or U7398 (N_7398,N_6869,N_6674);
or U7399 (N_7399,N_6904,N_6562);
xor U7400 (N_7400,N_6813,N_6856);
nand U7401 (N_7401,N_6709,N_6758);
or U7402 (N_7402,N_6520,N_6944);
nand U7403 (N_7403,N_6973,N_6747);
or U7404 (N_7404,N_6732,N_6653);
nor U7405 (N_7405,N_6647,N_6539);
or U7406 (N_7406,N_6904,N_6577);
xor U7407 (N_7407,N_6705,N_6739);
and U7408 (N_7408,N_6849,N_6947);
and U7409 (N_7409,N_6897,N_6921);
or U7410 (N_7410,N_6934,N_6580);
and U7411 (N_7411,N_6693,N_6748);
xnor U7412 (N_7412,N_6606,N_6649);
xnor U7413 (N_7413,N_6624,N_6505);
nand U7414 (N_7414,N_6628,N_6537);
xnor U7415 (N_7415,N_6587,N_6988);
xor U7416 (N_7416,N_6923,N_6803);
nand U7417 (N_7417,N_6814,N_6830);
nand U7418 (N_7418,N_6771,N_6859);
nor U7419 (N_7419,N_6737,N_6726);
xor U7420 (N_7420,N_6549,N_6891);
nand U7421 (N_7421,N_6596,N_6969);
and U7422 (N_7422,N_6751,N_6857);
and U7423 (N_7423,N_6832,N_6707);
or U7424 (N_7424,N_6952,N_6918);
or U7425 (N_7425,N_6626,N_6819);
or U7426 (N_7426,N_6514,N_6819);
and U7427 (N_7427,N_6567,N_6808);
and U7428 (N_7428,N_6677,N_6681);
or U7429 (N_7429,N_6513,N_6557);
nand U7430 (N_7430,N_6970,N_6929);
nand U7431 (N_7431,N_6824,N_6735);
and U7432 (N_7432,N_6763,N_6588);
nor U7433 (N_7433,N_6844,N_6947);
xnor U7434 (N_7434,N_6794,N_6712);
and U7435 (N_7435,N_6933,N_6916);
and U7436 (N_7436,N_6981,N_6820);
nor U7437 (N_7437,N_6846,N_6500);
nor U7438 (N_7438,N_6860,N_6550);
and U7439 (N_7439,N_6747,N_6531);
and U7440 (N_7440,N_6958,N_6659);
or U7441 (N_7441,N_6945,N_6519);
or U7442 (N_7442,N_6513,N_6962);
or U7443 (N_7443,N_6821,N_6839);
and U7444 (N_7444,N_6910,N_6629);
or U7445 (N_7445,N_6570,N_6946);
xor U7446 (N_7446,N_6812,N_6946);
xor U7447 (N_7447,N_6828,N_6727);
nor U7448 (N_7448,N_6523,N_6934);
nor U7449 (N_7449,N_6831,N_6680);
nand U7450 (N_7450,N_6727,N_6955);
xnor U7451 (N_7451,N_6572,N_6790);
nand U7452 (N_7452,N_6942,N_6594);
xor U7453 (N_7453,N_6639,N_6614);
nor U7454 (N_7454,N_6804,N_6814);
xnor U7455 (N_7455,N_6610,N_6957);
xnor U7456 (N_7456,N_6842,N_6913);
and U7457 (N_7457,N_6559,N_6773);
or U7458 (N_7458,N_6516,N_6605);
or U7459 (N_7459,N_6704,N_6905);
nor U7460 (N_7460,N_6877,N_6741);
or U7461 (N_7461,N_6927,N_6928);
or U7462 (N_7462,N_6850,N_6736);
nand U7463 (N_7463,N_6818,N_6661);
or U7464 (N_7464,N_6542,N_6965);
nor U7465 (N_7465,N_6771,N_6543);
and U7466 (N_7466,N_6605,N_6985);
or U7467 (N_7467,N_6853,N_6894);
nand U7468 (N_7468,N_6620,N_6631);
nand U7469 (N_7469,N_6831,N_6548);
or U7470 (N_7470,N_6951,N_6608);
and U7471 (N_7471,N_6954,N_6617);
xnor U7472 (N_7472,N_6571,N_6679);
and U7473 (N_7473,N_6693,N_6539);
xor U7474 (N_7474,N_6598,N_6532);
or U7475 (N_7475,N_6631,N_6994);
nand U7476 (N_7476,N_6515,N_6665);
and U7477 (N_7477,N_6615,N_6727);
and U7478 (N_7478,N_6598,N_6561);
nand U7479 (N_7479,N_6723,N_6600);
nand U7480 (N_7480,N_6833,N_6539);
and U7481 (N_7481,N_6814,N_6900);
nand U7482 (N_7482,N_6627,N_6560);
or U7483 (N_7483,N_6558,N_6794);
nor U7484 (N_7484,N_6682,N_6775);
nor U7485 (N_7485,N_6931,N_6700);
nand U7486 (N_7486,N_6766,N_6758);
nor U7487 (N_7487,N_6965,N_6557);
nor U7488 (N_7488,N_6933,N_6720);
or U7489 (N_7489,N_6737,N_6936);
xnor U7490 (N_7490,N_6734,N_6791);
nand U7491 (N_7491,N_6936,N_6627);
nor U7492 (N_7492,N_6585,N_6602);
or U7493 (N_7493,N_6958,N_6916);
and U7494 (N_7494,N_6801,N_6620);
nor U7495 (N_7495,N_6885,N_6555);
nor U7496 (N_7496,N_6628,N_6871);
and U7497 (N_7497,N_6978,N_6697);
xnor U7498 (N_7498,N_6596,N_6999);
and U7499 (N_7499,N_6509,N_6885);
nand U7500 (N_7500,N_7340,N_7301);
xnor U7501 (N_7501,N_7469,N_7334);
nor U7502 (N_7502,N_7140,N_7431);
nand U7503 (N_7503,N_7433,N_7394);
or U7504 (N_7504,N_7008,N_7136);
nand U7505 (N_7505,N_7246,N_7261);
xor U7506 (N_7506,N_7476,N_7210);
xor U7507 (N_7507,N_7318,N_7275);
or U7508 (N_7508,N_7216,N_7420);
nand U7509 (N_7509,N_7101,N_7300);
xor U7510 (N_7510,N_7305,N_7422);
or U7511 (N_7511,N_7317,N_7247);
nand U7512 (N_7512,N_7360,N_7090);
nand U7513 (N_7513,N_7373,N_7039);
xnor U7514 (N_7514,N_7414,N_7458);
or U7515 (N_7515,N_7280,N_7480);
or U7516 (N_7516,N_7408,N_7111);
or U7517 (N_7517,N_7288,N_7016);
xor U7518 (N_7518,N_7400,N_7439);
and U7519 (N_7519,N_7377,N_7185);
xor U7520 (N_7520,N_7329,N_7260);
nand U7521 (N_7521,N_7000,N_7004);
or U7522 (N_7522,N_7158,N_7214);
xor U7523 (N_7523,N_7212,N_7355);
nor U7524 (N_7524,N_7027,N_7279);
and U7525 (N_7525,N_7201,N_7015);
nand U7526 (N_7526,N_7089,N_7436);
and U7527 (N_7527,N_7479,N_7134);
nor U7528 (N_7528,N_7467,N_7012);
or U7529 (N_7529,N_7445,N_7253);
nand U7530 (N_7530,N_7354,N_7105);
xnor U7531 (N_7531,N_7072,N_7009);
nand U7532 (N_7532,N_7374,N_7265);
or U7533 (N_7533,N_7311,N_7082);
xnor U7534 (N_7534,N_7276,N_7310);
nand U7535 (N_7535,N_7130,N_7125);
xor U7536 (N_7536,N_7452,N_7187);
or U7537 (N_7537,N_7338,N_7120);
and U7538 (N_7538,N_7497,N_7177);
xnor U7539 (N_7539,N_7309,N_7100);
xnor U7540 (N_7540,N_7383,N_7332);
xor U7541 (N_7541,N_7440,N_7196);
nand U7542 (N_7542,N_7413,N_7026);
or U7543 (N_7543,N_7407,N_7416);
xor U7544 (N_7544,N_7115,N_7245);
nor U7545 (N_7545,N_7093,N_7228);
nand U7546 (N_7546,N_7382,N_7496);
and U7547 (N_7547,N_7403,N_7449);
nand U7548 (N_7548,N_7432,N_7267);
nand U7549 (N_7549,N_7017,N_7257);
xor U7550 (N_7550,N_7242,N_7491);
xor U7551 (N_7551,N_7281,N_7024);
and U7552 (N_7552,N_7266,N_7258);
or U7553 (N_7553,N_7363,N_7038);
nor U7554 (N_7554,N_7337,N_7193);
nand U7555 (N_7555,N_7356,N_7369);
nand U7556 (N_7556,N_7492,N_7207);
nand U7557 (N_7557,N_7060,N_7028);
nand U7558 (N_7558,N_7031,N_7396);
or U7559 (N_7559,N_7078,N_7219);
nand U7560 (N_7560,N_7164,N_7002);
and U7561 (N_7561,N_7215,N_7083);
xor U7562 (N_7562,N_7325,N_7342);
or U7563 (N_7563,N_7316,N_7142);
or U7564 (N_7564,N_7298,N_7457);
nor U7565 (N_7565,N_7068,N_7121);
and U7566 (N_7566,N_7252,N_7293);
and U7567 (N_7567,N_7483,N_7468);
and U7568 (N_7568,N_7345,N_7154);
nand U7569 (N_7569,N_7314,N_7045);
or U7570 (N_7570,N_7451,N_7042);
or U7571 (N_7571,N_7152,N_7241);
nand U7572 (N_7572,N_7204,N_7071);
and U7573 (N_7573,N_7108,N_7447);
nand U7574 (N_7574,N_7430,N_7263);
or U7575 (N_7575,N_7268,N_7147);
nor U7576 (N_7576,N_7198,N_7390);
and U7577 (N_7577,N_7126,N_7073);
xnor U7578 (N_7578,N_7455,N_7194);
nor U7579 (N_7579,N_7323,N_7456);
xor U7580 (N_7580,N_7132,N_7106);
nand U7581 (N_7581,N_7076,N_7099);
and U7582 (N_7582,N_7064,N_7264);
xnor U7583 (N_7583,N_7434,N_7348);
xor U7584 (N_7584,N_7035,N_7402);
xnor U7585 (N_7585,N_7240,N_7249);
nand U7586 (N_7586,N_7146,N_7077);
and U7587 (N_7587,N_7143,N_7367);
nor U7588 (N_7588,N_7251,N_7096);
xnor U7589 (N_7589,N_7107,N_7159);
nor U7590 (N_7590,N_7368,N_7444);
xnor U7591 (N_7591,N_7395,N_7113);
nor U7592 (N_7592,N_7290,N_7224);
or U7593 (N_7593,N_7371,N_7389);
nor U7594 (N_7594,N_7061,N_7010);
or U7595 (N_7595,N_7464,N_7191);
or U7596 (N_7596,N_7427,N_7297);
xor U7597 (N_7597,N_7429,N_7322);
xor U7598 (N_7598,N_7361,N_7151);
nand U7599 (N_7599,N_7302,N_7087);
nand U7600 (N_7600,N_7284,N_7052);
and U7601 (N_7601,N_7353,N_7426);
or U7602 (N_7602,N_7192,N_7349);
nand U7603 (N_7603,N_7347,N_7172);
and U7604 (N_7604,N_7404,N_7285);
nor U7605 (N_7605,N_7482,N_7104);
xor U7606 (N_7606,N_7295,N_7123);
and U7607 (N_7607,N_7231,N_7425);
nand U7608 (N_7608,N_7428,N_7366);
or U7609 (N_7609,N_7448,N_7291);
nand U7610 (N_7610,N_7054,N_7047);
nand U7611 (N_7611,N_7270,N_7376);
and U7612 (N_7612,N_7161,N_7036);
nor U7613 (N_7613,N_7315,N_7379);
xnor U7614 (N_7614,N_7046,N_7238);
nand U7615 (N_7615,N_7109,N_7211);
nand U7616 (N_7616,N_7461,N_7074);
xor U7617 (N_7617,N_7135,N_7206);
or U7618 (N_7618,N_7237,N_7180);
nand U7619 (N_7619,N_7227,N_7163);
xor U7620 (N_7620,N_7014,N_7188);
nand U7621 (N_7621,N_7033,N_7179);
nand U7622 (N_7622,N_7048,N_7062);
and U7623 (N_7623,N_7313,N_7114);
or U7624 (N_7624,N_7223,N_7043);
and U7625 (N_7625,N_7375,N_7088);
nor U7626 (N_7626,N_7013,N_7319);
and U7627 (N_7627,N_7243,N_7272);
nor U7628 (N_7628,N_7475,N_7183);
nor U7629 (N_7629,N_7499,N_7058);
nor U7630 (N_7630,N_7128,N_7041);
nor U7631 (N_7631,N_7085,N_7443);
nand U7632 (N_7632,N_7029,N_7025);
xor U7633 (N_7633,N_7166,N_7195);
xor U7634 (N_7634,N_7330,N_7118);
xor U7635 (N_7635,N_7103,N_7442);
xnor U7636 (N_7636,N_7157,N_7358);
and U7637 (N_7637,N_7391,N_7040);
nand U7638 (N_7638,N_7001,N_7079);
nand U7639 (N_7639,N_7308,N_7067);
or U7640 (N_7640,N_7186,N_7484);
nand U7641 (N_7641,N_7486,N_7044);
xnor U7642 (N_7642,N_7156,N_7388);
and U7643 (N_7643,N_7006,N_7129);
nor U7644 (N_7644,N_7019,N_7303);
nand U7645 (N_7645,N_7450,N_7094);
or U7646 (N_7646,N_7144,N_7287);
or U7647 (N_7647,N_7435,N_7170);
and U7648 (N_7648,N_7080,N_7406);
nor U7649 (N_7649,N_7221,N_7057);
or U7650 (N_7650,N_7075,N_7490);
or U7651 (N_7651,N_7141,N_7454);
and U7652 (N_7652,N_7182,N_7133);
xor U7653 (N_7653,N_7437,N_7190);
xor U7654 (N_7654,N_7362,N_7419);
and U7655 (N_7655,N_7112,N_7155);
or U7656 (N_7656,N_7417,N_7149);
xnor U7657 (N_7657,N_7127,N_7131);
or U7658 (N_7658,N_7477,N_7021);
and U7659 (N_7659,N_7289,N_7091);
and U7660 (N_7660,N_7478,N_7160);
nor U7661 (N_7661,N_7065,N_7095);
nand U7662 (N_7662,N_7327,N_7222);
nor U7663 (N_7663,N_7271,N_7359);
xor U7664 (N_7664,N_7494,N_7066);
or U7665 (N_7665,N_7385,N_7168);
nand U7666 (N_7666,N_7466,N_7070);
and U7667 (N_7667,N_7259,N_7357);
xnor U7668 (N_7668,N_7336,N_7056);
and U7669 (N_7669,N_7411,N_7471);
nor U7670 (N_7670,N_7063,N_7324);
xor U7671 (N_7671,N_7339,N_7232);
xor U7672 (N_7672,N_7234,N_7392);
nand U7673 (N_7673,N_7165,N_7399);
nor U7674 (N_7674,N_7122,N_7370);
or U7675 (N_7675,N_7018,N_7364);
nor U7676 (N_7676,N_7269,N_7384);
nand U7677 (N_7677,N_7421,N_7493);
or U7678 (N_7678,N_7299,N_7333);
xnor U7679 (N_7679,N_7321,N_7032);
xnor U7680 (N_7680,N_7487,N_7199);
and U7681 (N_7681,N_7495,N_7352);
or U7682 (N_7682,N_7296,N_7007);
nor U7683 (N_7683,N_7472,N_7335);
and U7684 (N_7684,N_7346,N_7167);
or U7685 (N_7685,N_7460,N_7424);
nand U7686 (N_7686,N_7116,N_7277);
nor U7687 (N_7687,N_7173,N_7307);
xor U7688 (N_7688,N_7050,N_7169);
and U7689 (N_7689,N_7286,N_7244);
xor U7690 (N_7690,N_7453,N_7341);
and U7691 (N_7691,N_7378,N_7459);
nand U7692 (N_7692,N_7262,N_7412);
and U7693 (N_7693,N_7181,N_7003);
xor U7694 (N_7694,N_7176,N_7059);
and U7695 (N_7695,N_7441,N_7312);
or U7696 (N_7696,N_7320,N_7401);
xor U7697 (N_7697,N_7184,N_7485);
and U7698 (N_7698,N_7139,N_7150);
and U7699 (N_7699,N_7119,N_7055);
nor U7700 (N_7700,N_7235,N_7189);
xor U7701 (N_7701,N_7197,N_7473);
and U7702 (N_7702,N_7409,N_7034);
xor U7703 (N_7703,N_7023,N_7053);
xnor U7704 (N_7704,N_7248,N_7092);
and U7705 (N_7705,N_7381,N_7380);
nand U7706 (N_7706,N_7049,N_7153);
xor U7707 (N_7707,N_7350,N_7097);
or U7708 (N_7708,N_7331,N_7498);
nor U7709 (N_7709,N_7145,N_7202);
xor U7710 (N_7710,N_7306,N_7203);
nor U7711 (N_7711,N_7465,N_7229);
and U7712 (N_7712,N_7294,N_7171);
xnor U7713 (N_7713,N_7397,N_7239);
xor U7714 (N_7714,N_7069,N_7137);
xor U7715 (N_7715,N_7254,N_7225);
or U7716 (N_7716,N_7292,N_7446);
or U7717 (N_7717,N_7393,N_7274);
or U7718 (N_7718,N_7230,N_7423);
nor U7719 (N_7719,N_7213,N_7386);
or U7720 (N_7720,N_7005,N_7365);
or U7721 (N_7721,N_7304,N_7086);
or U7722 (N_7722,N_7328,N_7030);
xor U7723 (N_7723,N_7343,N_7351);
nand U7724 (N_7724,N_7084,N_7110);
and U7725 (N_7725,N_7326,N_7282);
xnor U7726 (N_7726,N_7037,N_7344);
and U7727 (N_7727,N_7418,N_7162);
and U7728 (N_7728,N_7148,N_7205);
nand U7729 (N_7729,N_7474,N_7481);
nor U7730 (N_7730,N_7174,N_7273);
nor U7731 (N_7731,N_7438,N_7138);
or U7732 (N_7732,N_7200,N_7102);
nor U7733 (N_7733,N_7278,N_7250);
nand U7734 (N_7734,N_7217,N_7081);
or U7735 (N_7735,N_7218,N_7209);
and U7736 (N_7736,N_7489,N_7462);
nor U7737 (N_7737,N_7226,N_7256);
nor U7738 (N_7738,N_7022,N_7233);
nor U7739 (N_7739,N_7051,N_7372);
and U7740 (N_7740,N_7470,N_7220);
xnor U7741 (N_7741,N_7488,N_7175);
xnor U7742 (N_7742,N_7405,N_7415);
nand U7743 (N_7743,N_7098,N_7398);
or U7744 (N_7744,N_7020,N_7178);
xor U7745 (N_7745,N_7011,N_7410);
and U7746 (N_7746,N_7208,N_7117);
xor U7747 (N_7747,N_7283,N_7463);
or U7748 (N_7748,N_7387,N_7255);
nor U7749 (N_7749,N_7124,N_7236);
nor U7750 (N_7750,N_7391,N_7192);
nor U7751 (N_7751,N_7490,N_7436);
and U7752 (N_7752,N_7174,N_7093);
nor U7753 (N_7753,N_7417,N_7352);
nor U7754 (N_7754,N_7014,N_7438);
and U7755 (N_7755,N_7132,N_7403);
nor U7756 (N_7756,N_7007,N_7158);
nand U7757 (N_7757,N_7318,N_7380);
nand U7758 (N_7758,N_7499,N_7459);
or U7759 (N_7759,N_7273,N_7324);
nor U7760 (N_7760,N_7023,N_7002);
xor U7761 (N_7761,N_7458,N_7184);
nand U7762 (N_7762,N_7021,N_7203);
nand U7763 (N_7763,N_7337,N_7446);
nand U7764 (N_7764,N_7132,N_7301);
nand U7765 (N_7765,N_7230,N_7210);
or U7766 (N_7766,N_7080,N_7027);
xor U7767 (N_7767,N_7143,N_7088);
nor U7768 (N_7768,N_7070,N_7468);
nand U7769 (N_7769,N_7070,N_7021);
and U7770 (N_7770,N_7111,N_7328);
and U7771 (N_7771,N_7021,N_7309);
nor U7772 (N_7772,N_7056,N_7061);
xor U7773 (N_7773,N_7170,N_7322);
nor U7774 (N_7774,N_7106,N_7060);
nor U7775 (N_7775,N_7447,N_7041);
nand U7776 (N_7776,N_7161,N_7325);
nor U7777 (N_7777,N_7264,N_7398);
nor U7778 (N_7778,N_7084,N_7329);
or U7779 (N_7779,N_7043,N_7167);
xnor U7780 (N_7780,N_7208,N_7090);
and U7781 (N_7781,N_7323,N_7340);
or U7782 (N_7782,N_7301,N_7449);
or U7783 (N_7783,N_7346,N_7128);
nand U7784 (N_7784,N_7430,N_7245);
nand U7785 (N_7785,N_7169,N_7285);
nand U7786 (N_7786,N_7094,N_7204);
nor U7787 (N_7787,N_7198,N_7190);
and U7788 (N_7788,N_7344,N_7361);
xnor U7789 (N_7789,N_7465,N_7400);
nand U7790 (N_7790,N_7185,N_7235);
nand U7791 (N_7791,N_7060,N_7146);
or U7792 (N_7792,N_7272,N_7033);
nor U7793 (N_7793,N_7039,N_7396);
nand U7794 (N_7794,N_7023,N_7017);
nor U7795 (N_7795,N_7351,N_7230);
or U7796 (N_7796,N_7401,N_7482);
nor U7797 (N_7797,N_7191,N_7083);
xnor U7798 (N_7798,N_7307,N_7252);
xor U7799 (N_7799,N_7334,N_7367);
or U7800 (N_7800,N_7476,N_7467);
xnor U7801 (N_7801,N_7105,N_7319);
xor U7802 (N_7802,N_7283,N_7280);
nor U7803 (N_7803,N_7094,N_7407);
and U7804 (N_7804,N_7286,N_7440);
or U7805 (N_7805,N_7437,N_7128);
nand U7806 (N_7806,N_7264,N_7214);
nand U7807 (N_7807,N_7333,N_7223);
nor U7808 (N_7808,N_7392,N_7376);
or U7809 (N_7809,N_7054,N_7150);
or U7810 (N_7810,N_7381,N_7155);
nor U7811 (N_7811,N_7430,N_7447);
or U7812 (N_7812,N_7212,N_7485);
xnor U7813 (N_7813,N_7348,N_7435);
nor U7814 (N_7814,N_7061,N_7206);
xor U7815 (N_7815,N_7093,N_7286);
xnor U7816 (N_7816,N_7405,N_7488);
xnor U7817 (N_7817,N_7436,N_7066);
nor U7818 (N_7818,N_7394,N_7189);
xor U7819 (N_7819,N_7368,N_7333);
nor U7820 (N_7820,N_7121,N_7078);
or U7821 (N_7821,N_7001,N_7322);
xor U7822 (N_7822,N_7229,N_7348);
or U7823 (N_7823,N_7017,N_7169);
and U7824 (N_7824,N_7309,N_7452);
nor U7825 (N_7825,N_7322,N_7171);
or U7826 (N_7826,N_7278,N_7149);
nor U7827 (N_7827,N_7341,N_7088);
xnor U7828 (N_7828,N_7409,N_7085);
or U7829 (N_7829,N_7213,N_7264);
and U7830 (N_7830,N_7385,N_7292);
nor U7831 (N_7831,N_7158,N_7168);
xnor U7832 (N_7832,N_7066,N_7119);
xor U7833 (N_7833,N_7033,N_7462);
xor U7834 (N_7834,N_7405,N_7329);
nand U7835 (N_7835,N_7174,N_7137);
and U7836 (N_7836,N_7129,N_7283);
nor U7837 (N_7837,N_7239,N_7472);
and U7838 (N_7838,N_7014,N_7142);
nand U7839 (N_7839,N_7308,N_7039);
nor U7840 (N_7840,N_7060,N_7351);
or U7841 (N_7841,N_7073,N_7146);
nor U7842 (N_7842,N_7490,N_7244);
or U7843 (N_7843,N_7238,N_7095);
or U7844 (N_7844,N_7421,N_7283);
and U7845 (N_7845,N_7464,N_7367);
and U7846 (N_7846,N_7035,N_7209);
and U7847 (N_7847,N_7158,N_7046);
and U7848 (N_7848,N_7449,N_7068);
nand U7849 (N_7849,N_7443,N_7051);
and U7850 (N_7850,N_7010,N_7392);
nand U7851 (N_7851,N_7441,N_7109);
nor U7852 (N_7852,N_7034,N_7386);
nor U7853 (N_7853,N_7472,N_7232);
xnor U7854 (N_7854,N_7488,N_7311);
nor U7855 (N_7855,N_7169,N_7316);
nor U7856 (N_7856,N_7297,N_7380);
xor U7857 (N_7857,N_7014,N_7123);
nand U7858 (N_7858,N_7188,N_7363);
or U7859 (N_7859,N_7224,N_7302);
xnor U7860 (N_7860,N_7389,N_7178);
and U7861 (N_7861,N_7482,N_7133);
or U7862 (N_7862,N_7390,N_7062);
nor U7863 (N_7863,N_7474,N_7103);
nand U7864 (N_7864,N_7238,N_7114);
or U7865 (N_7865,N_7274,N_7180);
or U7866 (N_7866,N_7116,N_7156);
xnor U7867 (N_7867,N_7041,N_7066);
xor U7868 (N_7868,N_7394,N_7003);
xnor U7869 (N_7869,N_7483,N_7424);
nor U7870 (N_7870,N_7421,N_7165);
and U7871 (N_7871,N_7164,N_7235);
or U7872 (N_7872,N_7100,N_7481);
nor U7873 (N_7873,N_7358,N_7418);
nor U7874 (N_7874,N_7231,N_7137);
nand U7875 (N_7875,N_7033,N_7231);
nor U7876 (N_7876,N_7226,N_7439);
nand U7877 (N_7877,N_7330,N_7235);
xor U7878 (N_7878,N_7480,N_7137);
nor U7879 (N_7879,N_7460,N_7148);
nand U7880 (N_7880,N_7031,N_7360);
xor U7881 (N_7881,N_7483,N_7498);
xor U7882 (N_7882,N_7466,N_7450);
nand U7883 (N_7883,N_7444,N_7489);
nor U7884 (N_7884,N_7039,N_7079);
or U7885 (N_7885,N_7127,N_7154);
or U7886 (N_7886,N_7426,N_7009);
nor U7887 (N_7887,N_7321,N_7402);
and U7888 (N_7888,N_7264,N_7083);
or U7889 (N_7889,N_7086,N_7294);
xor U7890 (N_7890,N_7275,N_7084);
xor U7891 (N_7891,N_7403,N_7304);
and U7892 (N_7892,N_7126,N_7432);
xor U7893 (N_7893,N_7190,N_7118);
or U7894 (N_7894,N_7005,N_7283);
or U7895 (N_7895,N_7204,N_7309);
xor U7896 (N_7896,N_7074,N_7316);
nor U7897 (N_7897,N_7185,N_7316);
or U7898 (N_7898,N_7228,N_7148);
xor U7899 (N_7899,N_7379,N_7365);
nand U7900 (N_7900,N_7255,N_7337);
or U7901 (N_7901,N_7209,N_7344);
and U7902 (N_7902,N_7378,N_7407);
nor U7903 (N_7903,N_7406,N_7089);
and U7904 (N_7904,N_7204,N_7108);
nand U7905 (N_7905,N_7223,N_7003);
nor U7906 (N_7906,N_7467,N_7426);
xnor U7907 (N_7907,N_7442,N_7401);
and U7908 (N_7908,N_7310,N_7213);
or U7909 (N_7909,N_7340,N_7471);
nor U7910 (N_7910,N_7435,N_7418);
or U7911 (N_7911,N_7130,N_7168);
and U7912 (N_7912,N_7423,N_7058);
xnor U7913 (N_7913,N_7435,N_7426);
nand U7914 (N_7914,N_7490,N_7089);
or U7915 (N_7915,N_7033,N_7411);
or U7916 (N_7916,N_7386,N_7345);
and U7917 (N_7917,N_7325,N_7389);
or U7918 (N_7918,N_7274,N_7203);
or U7919 (N_7919,N_7499,N_7337);
and U7920 (N_7920,N_7284,N_7340);
xnor U7921 (N_7921,N_7435,N_7161);
xor U7922 (N_7922,N_7065,N_7129);
nor U7923 (N_7923,N_7204,N_7442);
nor U7924 (N_7924,N_7253,N_7012);
and U7925 (N_7925,N_7224,N_7412);
and U7926 (N_7926,N_7012,N_7196);
xor U7927 (N_7927,N_7026,N_7258);
and U7928 (N_7928,N_7249,N_7287);
nor U7929 (N_7929,N_7434,N_7083);
and U7930 (N_7930,N_7267,N_7433);
xor U7931 (N_7931,N_7184,N_7464);
nand U7932 (N_7932,N_7461,N_7226);
nor U7933 (N_7933,N_7367,N_7429);
xor U7934 (N_7934,N_7484,N_7300);
or U7935 (N_7935,N_7307,N_7419);
or U7936 (N_7936,N_7488,N_7419);
and U7937 (N_7937,N_7137,N_7325);
nor U7938 (N_7938,N_7032,N_7148);
xnor U7939 (N_7939,N_7423,N_7460);
xor U7940 (N_7940,N_7494,N_7098);
nor U7941 (N_7941,N_7143,N_7140);
and U7942 (N_7942,N_7414,N_7383);
or U7943 (N_7943,N_7184,N_7476);
xor U7944 (N_7944,N_7456,N_7469);
xor U7945 (N_7945,N_7103,N_7382);
or U7946 (N_7946,N_7182,N_7170);
and U7947 (N_7947,N_7011,N_7017);
nand U7948 (N_7948,N_7103,N_7467);
nand U7949 (N_7949,N_7139,N_7433);
xnor U7950 (N_7950,N_7028,N_7391);
xor U7951 (N_7951,N_7082,N_7431);
xnor U7952 (N_7952,N_7156,N_7088);
nand U7953 (N_7953,N_7489,N_7384);
xnor U7954 (N_7954,N_7364,N_7281);
nor U7955 (N_7955,N_7333,N_7293);
and U7956 (N_7956,N_7159,N_7149);
and U7957 (N_7957,N_7038,N_7353);
and U7958 (N_7958,N_7498,N_7163);
nand U7959 (N_7959,N_7428,N_7342);
nand U7960 (N_7960,N_7290,N_7250);
nor U7961 (N_7961,N_7111,N_7373);
xnor U7962 (N_7962,N_7221,N_7069);
nand U7963 (N_7963,N_7218,N_7213);
or U7964 (N_7964,N_7262,N_7109);
and U7965 (N_7965,N_7223,N_7274);
xor U7966 (N_7966,N_7225,N_7213);
nor U7967 (N_7967,N_7234,N_7221);
nor U7968 (N_7968,N_7378,N_7105);
nand U7969 (N_7969,N_7128,N_7109);
and U7970 (N_7970,N_7246,N_7263);
or U7971 (N_7971,N_7075,N_7482);
and U7972 (N_7972,N_7254,N_7083);
and U7973 (N_7973,N_7396,N_7050);
xnor U7974 (N_7974,N_7210,N_7344);
nand U7975 (N_7975,N_7287,N_7283);
and U7976 (N_7976,N_7309,N_7130);
and U7977 (N_7977,N_7091,N_7272);
and U7978 (N_7978,N_7425,N_7012);
nand U7979 (N_7979,N_7189,N_7458);
nand U7980 (N_7980,N_7118,N_7408);
nand U7981 (N_7981,N_7139,N_7410);
nor U7982 (N_7982,N_7494,N_7192);
or U7983 (N_7983,N_7480,N_7471);
or U7984 (N_7984,N_7342,N_7131);
and U7985 (N_7985,N_7181,N_7479);
nand U7986 (N_7986,N_7362,N_7059);
or U7987 (N_7987,N_7356,N_7434);
nor U7988 (N_7988,N_7138,N_7261);
and U7989 (N_7989,N_7109,N_7298);
and U7990 (N_7990,N_7240,N_7459);
xor U7991 (N_7991,N_7237,N_7148);
nand U7992 (N_7992,N_7212,N_7326);
or U7993 (N_7993,N_7325,N_7397);
nor U7994 (N_7994,N_7425,N_7137);
and U7995 (N_7995,N_7351,N_7030);
nor U7996 (N_7996,N_7244,N_7264);
nand U7997 (N_7997,N_7233,N_7430);
or U7998 (N_7998,N_7179,N_7071);
and U7999 (N_7999,N_7105,N_7166);
and U8000 (N_8000,N_7840,N_7546);
xor U8001 (N_8001,N_7678,N_7581);
or U8002 (N_8002,N_7607,N_7574);
nand U8003 (N_8003,N_7972,N_7812);
or U8004 (N_8004,N_7951,N_7532);
and U8005 (N_8005,N_7758,N_7872);
nand U8006 (N_8006,N_7578,N_7770);
or U8007 (N_8007,N_7647,N_7804);
nor U8008 (N_8008,N_7708,N_7945);
and U8009 (N_8009,N_7886,N_7879);
xnor U8010 (N_8010,N_7825,N_7941);
and U8011 (N_8011,N_7746,N_7599);
or U8012 (N_8012,N_7779,N_7668);
and U8013 (N_8013,N_7997,N_7768);
nor U8014 (N_8014,N_7557,N_7965);
and U8015 (N_8015,N_7816,N_7631);
nand U8016 (N_8016,N_7595,N_7549);
xor U8017 (N_8017,N_7786,N_7508);
nor U8018 (N_8018,N_7521,N_7967);
xor U8019 (N_8019,N_7633,N_7792);
nor U8020 (N_8020,N_7656,N_7909);
or U8021 (N_8021,N_7822,N_7857);
nand U8022 (N_8022,N_7676,N_7712);
nor U8023 (N_8023,N_7893,N_7554);
xor U8024 (N_8024,N_7675,N_7700);
xnor U8025 (N_8025,N_7698,N_7918);
nand U8026 (N_8026,N_7826,N_7908);
xnor U8027 (N_8027,N_7805,N_7733);
nor U8028 (N_8028,N_7653,N_7960);
and U8029 (N_8029,N_7926,N_7902);
xor U8030 (N_8030,N_7524,N_7692);
or U8031 (N_8031,N_7571,N_7584);
or U8032 (N_8032,N_7637,N_7867);
or U8033 (N_8033,N_7568,N_7576);
or U8034 (N_8034,N_7685,N_7780);
and U8035 (N_8035,N_7741,N_7562);
xor U8036 (N_8036,N_7527,N_7869);
nand U8037 (N_8037,N_7836,N_7525);
nand U8038 (N_8038,N_7946,N_7710);
nor U8039 (N_8039,N_7709,N_7986);
or U8040 (N_8040,N_7962,N_7978);
and U8041 (N_8041,N_7817,N_7787);
nand U8042 (N_8042,N_7610,N_7624);
and U8043 (N_8043,N_7646,N_7850);
nor U8044 (N_8044,N_7801,N_7854);
and U8045 (N_8045,N_7809,N_7907);
nor U8046 (N_8046,N_7517,N_7531);
nand U8047 (N_8047,N_7636,N_7791);
nor U8048 (N_8048,N_7785,N_7775);
nor U8049 (N_8049,N_7652,N_7534);
or U8050 (N_8050,N_7659,N_7910);
and U8051 (N_8051,N_7838,N_7711);
and U8052 (N_8052,N_7703,N_7530);
nor U8053 (N_8053,N_7949,N_7832);
nor U8054 (N_8054,N_7940,N_7953);
nor U8055 (N_8055,N_7639,N_7990);
nor U8056 (N_8056,N_7665,N_7778);
or U8057 (N_8057,N_7669,N_7625);
and U8058 (N_8058,N_7740,N_7555);
xor U8059 (N_8059,N_7852,N_7769);
and U8060 (N_8060,N_7706,N_7980);
xor U8061 (N_8061,N_7617,N_7861);
nand U8062 (N_8062,N_7923,N_7842);
xnor U8063 (N_8063,N_7721,N_7514);
or U8064 (N_8064,N_7605,N_7833);
nand U8065 (N_8065,N_7702,N_7888);
xor U8066 (N_8066,N_7885,N_7681);
and U8067 (N_8067,N_7849,N_7900);
nor U8068 (N_8068,N_7690,N_7863);
nand U8069 (N_8069,N_7734,N_7696);
nor U8070 (N_8070,N_7701,N_7823);
or U8071 (N_8071,N_7616,N_7602);
or U8072 (N_8072,N_7829,N_7577);
and U8073 (N_8073,N_7723,N_7586);
xor U8074 (N_8074,N_7901,N_7819);
xnor U8075 (N_8075,N_7715,N_7757);
or U8076 (N_8076,N_7998,N_7632);
nand U8077 (N_8077,N_7540,N_7561);
or U8078 (N_8078,N_7841,N_7977);
xnor U8079 (N_8079,N_7516,N_7529);
nand U8080 (N_8080,N_7795,N_7635);
or U8081 (N_8081,N_7815,N_7657);
nand U8082 (N_8082,N_7880,N_7650);
and U8083 (N_8083,N_7731,N_7630);
xor U8084 (N_8084,N_7954,N_7982);
and U8085 (N_8085,N_7575,N_7619);
xor U8086 (N_8086,N_7883,N_7874);
or U8087 (N_8087,N_7512,N_7697);
nor U8088 (N_8088,N_7916,N_7970);
and U8089 (N_8089,N_7806,N_7627);
nor U8090 (N_8090,N_7594,N_7763);
and U8091 (N_8091,N_7856,N_7773);
nand U8092 (N_8092,N_7518,N_7713);
nor U8093 (N_8093,N_7543,N_7749);
nand U8094 (N_8094,N_7936,N_7563);
and U8095 (N_8095,N_7567,N_7913);
nand U8096 (N_8096,N_7547,N_7535);
and U8097 (N_8097,N_7590,N_7988);
nand U8098 (N_8098,N_7559,N_7727);
and U8099 (N_8099,N_7844,N_7660);
or U8100 (N_8100,N_7572,N_7608);
xnor U8101 (N_8101,N_7755,N_7771);
and U8102 (N_8102,N_7810,N_7903);
or U8103 (N_8103,N_7912,N_7649);
xor U8104 (N_8104,N_7742,N_7634);
nor U8105 (N_8105,N_7875,N_7767);
xnor U8106 (N_8106,N_7828,N_7975);
nor U8107 (N_8107,N_7588,N_7851);
xnor U8108 (N_8108,N_7609,N_7969);
and U8109 (N_8109,N_7745,N_7853);
nor U8110 (N_8110,N_7570,N_7762);
and U8111 (N_8111,N_7983,N_7550);
nor U8112 (N_8112,N_7612,N_7800);
or U8113 (N_8113,N_7515,N_7662);
or U8114 (N_8114,N_7878,N_7569);
or U8115 (N_8115,N_7759,N_7553);
and U8116 (N_8116,N_7580,N_7859);
and U8117 (N_8117,N_7994,N_7536);
nor U8118 (N_8118,N_7661,N_7989);
xor U8119 (N_8119,N_7579,N_7925);
or U8120 (N_8120,N_7987,N_7922);
nor U8121 (N_8121,N_7976,N_7620);
nand U8122 (N_8122,N_7958,N_7752);
nand U8123 (N_8123,N_7691,N_7519);
nor U8124 (N_8124,N_7682,N_7783);
or U8125 (N_8125,N_7939,N_7848);
xor U8126 (N_8126,N_7642,N_7993);
and U8127 (N_8127,N_7956,N_7931);
and U8128 (N_8128,N_7797,N_7917);
or U8129 (N_8129,N_7558,N_7716);
nor U8130 (N_8130,N_7585,N_7876);
or U8131 (N_8131,N_7793,N_7726);
nor U8132 (N_8132,N_7843,N_7655);
or U8133 (N_8133,N_7944,N_7808);
nor U8134 (N_8134,N_7729,N_7981);
and U8135 (N_8135,N_7618,N_7756);
nand U8136 (N_8136,N_7915,N_7807);
and U8137 (N_8137,N_7720,N_7603);
nand U8138 (N_8138,N_7587,N_7674);
or U8139 (N_8139,N_7928,N_7528);
xor U8140 (N_8140,N_7545,N_7526);
xnor U8141 (N_8141,N_7743,N_7704);
and U8142 (N_8142,N_7699,N_7613);
nor U8143 (N_8143,N_7796,N_7884);
xnor U8144 (N_8144,N_7537,N_7592);
xnor U8145 (N_8145,N_7739,N_7898);
and U8146 (N_8146,N_7513,N_7552);
or U8147 (N_8147,N_7934,N_7947);
and U8148 (N_8148,N_7604,N_7730);
or U8149 (N_8149,N_7952,N_7522);
nor U8150 (N_8150,N_7667,N_7628);
and U8151 (N_8151,N_7920,N_7979);
xor U8152 (N_8152,N_7641,N_7950);
and U8153 (N_8153,N_7764,N_7680);
nor U8154 (N_8154,N_7894,N_7629);
xnor U8155 (N_8155,N_7868,N_7695);
and U8156 (N_8156,N_7761,N_7736);
nor U8157 (N_8157,N_7506,N_7503);
nand U8158 (N_8158,N_7643,N_7666);
nand U8159 (N_8159,N_7974,N_7948);
and U8160 (N_8160,N_7935,N_7924);
or U8161 (N_8161,N_7672,N_7593);
and U8162 (N_8162,N_7626,N_7565);
nand U8163 (N_8163,N_7583,N_7985);
xor U8164 (N_8164,N_7664,N_7523);
xnor U8165 (N_8165,N_7638,N_7813);
nor U8166 (N_8166,N_7765,N_7510);
or U8167 (N_8167,N_7520,N_7718);
and U8168 (N_8168,N_7957,N_7648);
or U8169 (N_8169,N_7573,N_7799);
or U8170 (N_8170,N_7673,N_7644);
and U8171 (N_8171,N_7784,N_7938);
xor U8172 (N_8172,N_7564,N_7747);
nand U8173 (N_8173,N_7961,N_7847);
nor U8174 (N_8174,N_7866,N_7899);
xnor U8175 (N_8175,N_7919,N_7845);
nor U8176 (N_8176,N_7651,N_7670);
and U8177 (N_8177,N_7827,N_7995);
or U8178 (N_8178,N_7914,N_7622);
or U8179 (N_8179,N_7542,N_7694);
xnor U8180 (N_8180,N_7846,N_7904);
nand U8181 (N_8181,N_7548,N_7533);
xnor U8182 (N_8182,N_7890,N_7860);
and U8183 (N_8183,N_7640,N_7766);
nor U8184 (N_8184,N_7589,N_7927);
xnor U8185 (N_8185,N_7671,N_7679);
and U8186 (N_8186,N_7932,N_7556);
or U8187 (N_8187,N_7906,N_7751);
xnor U8188 (N_8188,N_7999,N_7889);
xor U8189 (N_8189,N_7933,N_7943);
or U8190 (N_8190,N_7887,N_7511);
nand U8191 (N_8191,N_7502,N_7966);
nand U8192 (N_8192,N_7737,N_7788);
or U8193 (N_8193,N_7873,N_7500);
nor U8194 (N_8194,N_7693,N_7782);
or U8195 (N_8195,N_7654,N_7501);
nand U8196 (N_8196,N_7539,N_7686);
nand U8197 (N_8197,N_7722,N_7621);
or U8198 (N_8198,N_7794,N_7677);
or U8199 (N_8199,N_7725,N_7753);
xor U8200 (N_8200,N_7858,N_7937);
nand U8201 (N_8201,N_7663,N_7790);
or U8202 (N_8202,N_7551,N_7748);
or U8203 (N_8203,N_7855,N_7688);
and U8204 (N_8204,N_7615,N_7831);
or U8205 (N_8205,N_7963,N_7871);
nand U8206 (N_8206,N_7566,N_7683);
and U8207 (N_8207,N_7802,N_7921);
xnor U8208 (N_8208,N_7882,N_7714);
or U8209 (N_8209,N_7968,N_7814);
and U8210 (N_8210,N_7964,N_7881);
or U8211 (N_8211,N_7509,N_7724);
and U8212 (N_8212,N_7774,N_7971);
and U8213 (N_8213,N_7892,N_7687);
and U8214 (N_8214,N_7835,N_7707);
and U8215 (N_8215,N_7839,N_7689);
xor U8216 (N_8216,N_7600,N_7623);
or U8217 (N_8217,N_7611,N_7973);
or U8218 (N_8218,N_7760,N_7705);
and U8219 (N_8219,N_7897,N_7959);
or U8220 (N_8220,N_7955,N_7591);
xnor U8221 (N_8221,N_7877,N_7834);
nand U8222 (N_8222,N_7830,N_7798);
nor U8223 (N_8223,N_7772,N_7821);
nand U8224 (N_8224,N_7837,N_7865);
xnor U8225 (N_8225,N_7744,N_7596);
and U8226 (N_8226,N_7811,N_7645);
or U8227 (N_8227,N_7597,N_7750);
nor U8228 (N_8228,N_7732,N_7606);
xnor U8229 (N_8229,N_7781,N_7684);
nor U8230 (N_8230,N_7717,N_7560);
nor U8231 (N_8231,N_7582,N_7992);
xnor U8232 (N_8232,N_7777,N_7864);
xor U8233 (N_8233,N_7789,N_7601);
and U8234 (N_8234,N_7614,N_7984);
or U8235 (N_8235,N_7991,N_7818);
or U8236 (N_8236,N_7862,N_7658);
or U8237 (N_8237,N_7544,N_7996);
nand U8238 (N_8238,N_7598,N_7824);
or U8239 (N_8239,N_7942,N_7719);
xor U8240 (N_8240,N_7541,N_7754);
nor U8241 (N_8241,N_7803,N_7738);
or U8242 (N_8242,N_7820,N_7905);
nor U8243 (N_8243,N_7870,N_7896);
or U8244 (N_8244,N_7507,N_7776);
nor U8245 (N_8245,N_7505,N_7728);
xor U8246 (N_8246,N_7930,N_7911);
or U8247 (N_8247,N_7895,N_7735);
nand U8248 (N_8248,N_7929,N_7891);
and U8249 (N_8249,N_7538,N_7504);
xor U8250 (N_8250,N_7753,N_7892);
or U8251 (N_8251,N_7622,N_7791);
or U8252 (N_8252,N_7788,N_7594);
xnor U8253 (N_8253,N_7881,N_7859);
xor U8254 (N_8254,N_7576,N_7987);
xnor U8255 (N_8255,N_7577,N_7755);
and U8256 (N_8256,N_7965,N_7841);
xnor U8257 (N_8257,N_7602,N_7896);
xor U8258 (N_8258,N_7896,N_7892);
xnor U8259 (N_8259,N_7982,N_7622);
xor U8260 (N_8260,N_7683,N_7922);
nand U8261 (N_8261,N_7510,N_7503);
nand U8262 (N_8262,N_7789,N_7550);
nand U8263 (N_8263,N_7578,N_7959);
nor U8264 (N_8264,N_7864,N_7841);
xnor U8265 (N_8265,N_7929,N_7616);
xnor U8266 (N_8266,N_7999,N_7766);
nor U8267 (N_8267,N_7652,N_7947);
nor U8268 (N_8268,N_7651,N_7513);
xnor U8269 (N_8269,N_7689,N_7545);
and U8270 (N_8270,N_7751,N_7698);
nor U8271 (N_8271,N_7639,N_7855);
and U8272 (N_8272,N_7747,N_7788);
nand U8273 (N_8273,N_7574,N_7610);
xnor U8274 (N_8274,N_7576,N_7526);
and U8275 (N_8275,N_7593,N_7834);
or U8276 (N_8276,N_7793,N_7694);
or U8277 (N_8277,N_7622,N_7585);
nor U8278 (N_8278,N_7697,N_7776);
or U8279 (N_8279,N_7734,N_7737);
or U8280 (N_8280,N_7980,N_7969);
or U8281 (N_8281,N_7882,N_7550);
xor U8282 (N_8282,N_7898,N_7793);
and U8283 (N_8283,N_7761,N_7962);
nor U8284 (N_8284,N_7978,N_7743);
or U8285 (N_8285,N_7818,N_7826);
nand U8286 (N_8286,N_7969,N_7882);
or U8287 (N_8287,N_7724,N_7848);
nand U8288 (N_8288,N_7853,N_7571);
nand U8289 (N_8289,N_7743,N_7961);
and U8290 (N_8290,N_7714,N_7754);
or U8291 (N_8291,N_7735,N_7630);
nor U8292 (N_8292,N_7662,N_7517);
and U8293 (N_8293,N_7701,N_7983);
xor U8294 (N_8294,N_7643,N_7798);
nand U8295 (N_8295,N_7757,N_7737);
nand U8296 (N_8296,N_7558,N_7889);
nor U8297 (N_8297,N_7981,N_7832);
xnor U8298 (N_8298,N_7921,N_7650);
nand U8299 (N_8299,N_7562,N_7566);
xnor U8300 (N_8300,N_7984,N_7659);
xor U8301 (N_8301,N_7528,N_7840);
nand U8302 (N_8302,N_7620,N_7717);
xor U8303 (N_8303,N_7763,N_7921);
or U8304 (N_8304,N_7601,N_7815);
nand U8305 (N_8305,N_7603,N_7633);
nor U8306 (N_8306,N_7748,N_7968);
nand U8307 (N_8307,N_7549,N_7750);
or U8308 (N_8308,N_7994,N_7651);
and U8309 (N_8309,N_7920,N_7710);
and U8310 (N_8310,N_7728,N_7563);
nand U8311 (N_8311,N_7713,N_7924);
nor U8312 (N_8312,N_7986,N_7853);
nand U8313 (N_8313,N_7524,N_7532);
xor U8314 (N_8314,N_7580,N_7670);
nor U8315 (N_8315,N_7749,N_7526);
nor U8316 (N_8316,N_7578,N_7916);
xor U8317 (N_8317,N_7654,N_7755);
xnor U8318 (N_8318,N_7845,N_7519);
nand U8319 (N_8319,N_7580,N_7949);
and U8320 (N_8320,N_7641,N_7503);
xor U8321 (N_8321,N_7854,N_7815);
nand U8322 (N_8322,N_7638,N_7723);
nor U8323 (N_8323,N_7561,N_7586);
or U8324 (N_8324,N_7844,N_7651);
nor U8325 (N_8325,N_7853,N_7827);
xnor U8326 (N_8326,N_7901,N_7556);
or U8327 (N_8327,N_7863,N_7930);
nand U8328 (N_8328,N_7727,N_7666);
nand U8329 (N_8329,N_7509,N_7881);
xnor U8330 (N_8330,N_7780,N_7706);
nor U8331 (N_8331,N_7500,N_7656);
nor U8332 (N_8332,N_7626,N_7839);
nand U8333 (N_8333,N_7611,N_7507);
nand U8334 (N_8334,N_7662,N_7911);
or U8335 (N_8335,N_7662,N_7648);
nor U8336 (N_8336,N_7785,N_7678);
nor U8337 (N_8337,N_7524,N_7823);
or U8338 (N_8338,N_7951,N_7866);
nor U8339 (N_8339,N_7567,N_7809);
nand U8340 (N_8340,N_7796,N_7785);
and U8341 (N_8341,N_7556,N_7842);
nor U8342 (N_8342,N_7770,N_7786);
or U8343 (N_8343,N_7778,N_7601);
and U8344 (N_8344,N_7628,N_7719);
nor U8345 (N_8345,N_7704,N_7674);
nor U8346 (N_8346,N_7886,N_7956);
or U8347 (N_8347,N_7770,N_7551);
nor U8348 (N_8348,N_7719,N_7899);
nor U8349 (N_8349,N_7791,N_7908);
nand U8350 (N_8350,N_7992,N_7599);
and U8351 (N_8351,N_7886,N_7983);
nand U8352 (N_8352,N_7942,N_7846);
nand U8353 (N_8353,N_7637,N_7852);
nor U8354 (N_8354,N_7507,N_7901);
xnor U8355 (N_8355,N_7953,N_7781);
xnor U8356 (N_8356,N_7637,N_7975);
nor U8357 (N_8357,N_7617,N_7905);
nor U8358 (N_8358,N_7611,N_7928);
xnor U8359 (N_8359,N_7823,N_7728);
and U8360 (N_8360,N_7704,N_7694);
and U8361 (N_8361,N_7923,N_7988);
xor U8362 (N_8362,N_7880,N_7789);
xnor U8363 (N_8363,N_7534,N_7989);
nand U8364 (N_8364,N_7893,N_7690);
or U8365 (N_8365,N_7528,N_7885);
xnor U8366 (N_8366,N_7855,N_7996);
nand U8367 (N_8367,N_7871,N_7773);
xor U8368 (N_8368,N_7841,N_7868);
xor U8369 (N_8369,N_7511,N_7972);
nor U8370 (N_8370,N_7884,N_7849);
nor U8371 (N_8371,N_7611,N_7503);
xor U8372 (N_8372,N_7793,N_7942);
xor U8373 (N_8373,N_7645,N_7692);
nor U8374 (N_8374,N_7991,N_7992);
nand U8375 (N_8375,N_7910,N_7936);
nor U8376 (N_8376,N_7852,N_7895);
nor U8377 (N_8377,N_7776,N_7584);
and U8378 (N_8378,N_7949,N_7850);
or U8379 (N_8379,N_7672,N_7871);
and U8380 (N_8380,N_7677,N_7783);
nand U8381 (N_8381,N_7961,N_7592);
or U8382 (N_8382,N_7692,N_7724);
or U8383 (N_8383,N_7609,N_7769);
and U8384 (N_8384,N_7879,N_7823);
nor U8385 (N_8385,N_7773,N_7569);
nor U8386 (N_8386,N_7611,N_7872);
and U8387 (N_8387,N_7988,N_7633);
and U8388 (N_8388,N_7752,N_7719);
nor U8389 (N_8389,N_7673,N_7982);
and U8390 (N_8390,N_7507,N_7909);
nor U8391 (N_8391,N_7517,N_7637);
and U8392 (N_8392,N_7639,N_7653);
nand U8393 (N_8393,N_7715,N_7635);
nand U8394 (N_8394,N_7791,N_7975);
or U8395 (N_8395,N_7810,N_7884);
nor U8396 (N_8396,N_7862,N_7619);
and U8397 (N_8397,N_7963,N_7674);
or U8398 (N_8398,N_7501,N_7918);
or U8399 (N_8399,N_7950,N_7846);
nand U8400 (N_8400,N_7759,N_7636);
or U8401 (N_8401,N_7998,N_7859);
nand U8402 (N_8402,N_7764,N_7644);
nand U8403 (N_8403,N_7618,N_7712);
or U8404 (N_8404,N_7834,N_7556);
or U8405 (N_8405,N_7727,N_7711);
xor U8406 (N_8406,N_7809,N_7954);
xnor U8407 (N_8407,N_7957,N_7744);
or U8408 (N_8408,N_7963,N_7544);
or U8409 (N_8409,N_7549,N_7963);
or U8410 (N_8410,N_7896,N_7840);
nand U8411 (N_8411,N_7569,N_7629);
xor U8412 (N_8412,N_7992,N_7921);
or U8413 (N_8413,N_7611,N_7952);
nor U8414 (N_8414,N_7616,N_7609);
nand U8415 (N_8415,N_7939,N_7860);
xnor U8416 (N_8416,N_7579,N_7875);
or U8417 (N_8417,N_7692,N_7893);
nand U8418 (N_8418,N_7821,N_7693);
nand U8419 (N_8419,N_7780,N_7953);
nor U8420 (N_8420,N_7757,N_7660);
and U8421 (N_8421,N_7593,N_7698);
or U8422 (N_8422,N_7780,N_7671);
or U8423 (N_8423,N_7754,N_7899);
or U8424 (N_8424,N_7776,N_7816);
nor U8425 (N_8425,N_7859,N_7937);
xor U8426 (N_8426,N_7620,N_7543);
and U8427 (N_8427,N_7816,N_7508);
or U8428 (N_8428,N_7651,N_7745);
nand U8429 (N_8429,N_7514,N_7798);
xor U8430 (N_8430,N_7925,N_7518);
and U8431 (N_8431,N_7690,N_7968);
nand U8432 (N_8432,N_7669,N_7968);
and U8433 (N_8433,N_7557,N_7713);
xnor U8434 (N_8434,N_7509,N_7612);
nor U8435 (N_8435,N_7980,N_7911);
nor U8436 (N_8436,N_7639,N_7816);
and U8437 (N_8437,N_7828,N_7866);
or U8438 (N_8438,N_7636,N_7523);
or U8439 (N_8439,N_7634,N_7838);
nand U8440 (N_8440,N_7604,N_7616);
nor U8441 (N_8441,N_7703,N_7908);
or U8442 (N_8442,N_7587,N_7629);
and U8443 (N_8443,N_7762,N_7531);
xor U8444 (N_8444,N_7614,N_7580);
nand U8445 (N_8445,N_7759,N_7938);
xor U8446 (N_8446,N_7551,N_7808);
or U8447 (N_8447,N_7635,N_7654);
and U8448 (N_8448,N_7655,N_7980);
or U8449 (N_8449,N_7531,N_7773);
and U8450 (N_8450,N_7623,N_7509);
xor U8451 (N_8451,N_7936,N_7554);
nand U8452 (N_8452,N_7641,N_7513);
nand U8453 (N_8453,N_7504,N_7523);
nor U8454 (N_8454,N_7609,N_7795);
nand U8455 (N_8455,N_7909,N_7623);
nor U8456 (N_8456,N_7973,N_7645);
nand U8457 (N_8457,N_7822,N_7584);
and U8458 (N_8458,N_7811,N_7543);
xnor U8459 (N_8459,N_7784,N_7747);
nor U8460 (N_8460,N_7954,N_7824);
and U8461 (N_8461,N_7900,N_7955);
and U8462 (N_8462,N_7532,N_7745);
xnor U8463 (N_8463,N_7704,N_7863);
nor U8464 (N_8464,N_7900,N_7551);
or U8465 (N_8465,N_7634,N_7948);
nand U8466 (N_8466,N_7863,N_7859);
or U8467 (N_8467,N_7831,N_7939);
or U8468 (N_8468,N_7715,N_7669);
nor U8469 (N_8469,N_7511,N_7994);
xor U8470 (N_8470,N_7663,N_7881);
and U8471 (N_8471,N_7952,N_7897);
or U8472 (N_8472,N_7687,N_7686);
nor U8473 (N_8473,N_7577,N_7695);
nand U8474 (N_8474,N_7515,N_7733);
or U8475 (N_8475,N_7877,N_7847);
and U8476 (N_8476,N_7739,N_7734);
or U8477 (N_8477,N_7722,N_7557);
and U8478 (N_8478,N_7833,N_7847);
nand U8479 (N_8479,N_7811,N_7846);
nand U8480 (N_8480,N_7620,N_7995);
and U8481 (N_8481,N_7754,N_7870);
xnor U8482 (N_8482,N_7861,N_7650);
xnor U8483 (N_8483,N_7954,N_7558);
nor U8484 (N_8484,N_7633,N_7646);
or U8485 (N_8485,N_7817,N_7626);
or U8486 (N_8486,N_7761,N_7517);
nor U8487 (N_8487,N_7743,N_7744);
nor U8488 (N_8488,N_7702,N_7911);
and U8489 (N_8489,N_7523,N_7826);
or U8490 (N_8490,N_7678,N_7526);
or U8491 (N_8491,N_7765,N_7551);
and U8492 (N_8492,N_7970,N_7875);
xnor U8493 (N_8493,N_7584,N_7696);
nor U8494 (N_8494,N_7943,N_7603);
or U8495 (N_8495,N_7602,N_7976);
xor U8496 (N_8496,N_7552,N_7832);
or U8497 (N_8497,N_7884,N_7823);
nor U8498 (N_8498,N_7636,N_7702);
or U8499 (N_8499,N_7993,N_7904);
or U8500 (N_8500,N_8096,N_8412);
nor U8501 (N_8501,N_8106,N_8281);
nand U8502 (N_8502,N_8304,N_8011);
nor U8503 (N_8503,N_8295,N_8424);
nand U8504 (N_8504,N_8449,N_8030);
and U8505 (N_8505,N_8349,N_8296);
xnor U8506 (N_8506,N_8398,N_8028);
nor U8507 (N_8507,N_8276,N_8239);
nor U8508 (N_8508,N_8159,N_8050);
nor U8509 (N_8509,N_8306,N_8075);
nor U8510 (N_8510,N_8454,N_8329);
nand U8511 (N_8511,N_8245,N_8175);
or U8512 (N_8512,N_8383,N_8390);
nor U8513 (N_8513,N_8382,N_8078);
xnor U8514 (N_8514,N_8014,N_8413);
nor U8515 (N_8515,N_8077,N_8148);
and U8516 (N_8516,N_8461,N_8475);
xnor U8517 (N_8517,N_8355,N_8287);
or U8518 (N_8518,N_8373,N_8026);
xnor U8519 (N_8519,N_8049,N_8019);
nor U8520 (N_8520,N_8309,N_8328);
or U8521 (N_8521,N_8481,N_8008);
xor U8522 (N_8522,N_8445,N_8226);
or U8523 (N_8523,N_8406,N_8060);
nor U8524 (N_8524,N_8240,N_8319);
xor U8525 (N_8525,N_8352,N_8083);
xnor U8526 (N_8526,N_8271,N_8336);
nor U8527 (N_8527,N_8236,N_8044);
nor U8528 (N_8528,N_8299,N_8260);
nand U8529 (N_8529,N_8080,N_8114);
xnor U8530 (N_8530,N_8135,N_8300);
nor U8531 (N_8531,N_8079,N_8171);
nand U8532 (N_8532,N_8187,N_8323);
nand U8533 (N_8533,N_8491,N_8418);
nor U8534 (N_8534,N_8032,N_8053);
nand U8535 (N_8535,N_8205,N_8298);
nand U8536 (N_8536,N_8376,N_8474);
nand U8537 (N_8537,N_8097,N_8331);
nand U8538 (N_8538,N_8003,N_8270);
and U8539 (N_8539,N_8433,N_8487);
nor U8540 (N_8540,N_8219,N_8371);
nor U8541 (N_8541,N_8178,N_8153);
nand U8542 (N_8542,N_8102,N_8291);
and U8543 (N_8543,N_8499,N_8472);
nand U8544 (N_8544,N_8016,N_8176);
nor U8545 (N_8545,N_8090,N_8456);
or U8546 (N_8546,N_8082,N_8410);
nand U8547 (N_8547,N_8092,N_8172);
and U8548 (N_8548,N_8058,N_8068);
xnor U8549 (N_8549,N_8112,N_8256);
nand U8550 (N_8550,N_8193,N_8460);
or U8551 (N_8551,N_8294,N_8031);
or U8552 (N_8552,N_8094,N_8126);
or U8553 (N_8553,N_8483,N_8490);
nor U8554 (N_8554,N_8129,N_8134);
nand U8555 (N_8555,N_8301,N_8190);
nand U8556 (N_8556,N_8415,N_8488);
nand U8557 (N_8557,N_8272,N_8332);
and U8558 (N_8558,N_8268,N_8285);
and U8559 (N_8559,N_8045,N_8013);
and U8560 (N_8560,N_8105,N_8066);
nand U8561 (N_8561,N_8109,N_8452);
and U8562 (N_8562,N_8217,N_8107);
nand U8563 (N_8563,N_8363,N_8467);
nor U8564 (N_8564,N_8160,N_8275);
and U8565 (N_8565,N_8036,N_8221);
nor U8566 (N_8566,N_8293,N_8391);
or U8567 (N_8567,N_8130,N_8432);
or U8568 (N_8568,N_8209,N_8196);
nand U8569 (N_8569,N_8279,N_8348);
xor U8570 (N_8570,N_8225,N_8142);
nor U8571 (N_8571,N_8115,N_8229);
or U8572 (N_8572,N_8419,N_8216);
or U8573 (N_8573,N_8441,N_8335);
nor U8574 (N_8574,N_8156,N_8211);
xor U8575 (N_8575,N_8318,N_8163);
nor U8576 (N_8576,N_8496,N_8386);
xor U8577 (N_8577,N_8143,N_8284);
and U8578 (N_8578,N_8034,N_8244);
nand U8579 (N_8579,N_8151,N_8429);
xnor U8580 (N_8580,N_8110,N_8223);
nor U8581 (N_8581,N_8040,N_8465);
nand U8582 (N_8582,N_8458,N_8098);
and U8583 (N_8583,N_8266,N_8379);
or U8584 (N_8584,N_8029,N_8360);
xnor U8585 (N_8585,N_8054,N_8063);
xnor U8586 (N_8586,N_8101,N_8227);
and U8587 (N_8587,N_8124,N_8241);
nand U8588 (N_8588,N_8056,N_8108);
and U8589 (N_8589,N_8263,N_8435);
nand U8590 (N_8590,N_8039,N_8141);
nand U8591 (N_8591,N_8322,N_8400);
nor U8592 (N_8592,N_8118,N_8315);
or U8593 (N_8593,N_8194,N_8428);
nor U8594 (N_8594,N_8234,N_8147);
or U8595 (N_8595,N_8354,N_8392);
and U8596 (N_8596,N_8302,N_8146);
xnor U8597 (N_8597,N_8128,N_8057);
nand U8598 (N_8598,N_8316,N_8208);
xor U8599 (N_8599,N_8283,N_8486);
nand U8600 (N_8600,N_8366,N_8069);
or U8601 (N_8601,N_8158,N_8277);
or U8602 (N_8602,N_8189,N_8334);
xnor U8603 (N_8603,N_8377,N_8005);
and U8604 (N_8604,N_8177,N_8342);
xor U8605 (N_8605,N_8414,N_8340);
nor U8606 (N_8606,N_8401,N_8485);
nor U8607 (N_8607,N_8230,N_8116);
and U8608 (N_8608,N_8367,N_8140);
and U8609 (N_8609,N_8427,N_8222);
and U8610 (N_8610,N_8002,N_8048);
and U8611 (N_8611,N_8059,N_8370);
nor U8612 (N_8612,N_8215,N_8369);
xor U8613 (N_8613,N_8085,N_8007);
nor U8614 (N_8614,N_8292,N_8289);
and U8615 (N_8615,N_8123,N_8182);
and U8616 (N_8616,N_8265,N_8165);
xor U8617 (N_8617,N_8183,N_8385);
and U8618 (N_8618,N_8333,N_8246);
and U8619 (N_8619,N_8337,N_8199);
and U8620 (N_8620,N_8339,N_8478);
nor U8621 (N_8621,N_8437,N_8250);
and U8622 (N_8622,N_8001,N_8430);
nor U8623 (N_8623,N_8210,N_8198);
nor U8624 (N_8624,N_8408,N_8168);
nand U8625 (N_8625,N_8440,N_8378);
nor U8626 (N_8626,N_8254,N_8242);
or U8627 (N_8627,N_8368,N_8020);
or U8628 (N_8628,N_8493,N_8046);
or U8629 (N_8629,N_8073,N_8061);
nand U8630 (N_8630,N_8055,N_8154);
xor U8631 (N_8631,N_8426,N_8494);
and U8632 (N_8632,N_8374,N_8338);
nand U8633 (N_8633,N_8303,N_8071);
nor U8634 (N_8634,N_8062,N_8010);
xor U8635 (N_8635,N_8004,N_8131);
nand U8636 (N_8636,N_8203,N_8249);
and U8637 (N_8637,N_8439,N_8072);
or U8638 (N_8638,N_8006,N_8346);
or U8639 (N_8639,N_8425,N_8384);
nand U8640 (N_8640,N_8233,N_8018);
nand U8641 (N_8641,N_8353,N_8009);
and U8642 (N_8642,N_8409,N_8074);
or U8643 (N_8643,N_8104,N_8280);
nor U8644 (N_8644,N_8396,N_8468);
and U8645 (N_8645,N_8081,N_8136);
and U8646 (N_8646,N_8269,N_8195);
or U8647 (N_8647,N_8420,N_8327);
nand U8648 (N_8648,N_8477,N_8479);
nor U8649 (N_8649,N_8325,N_8047);
nand U8650 (N_8650,N_8100,N_8162);
or U8651 (N_8651,N_8357,N_8207);
nor U8652 (N_8652,N_8457,N_8197);
or U8653 (N_8653,N_8464,N_8345);
and U8654 (N_8654,N_8381,N_8259);
nand U8655 (N_8655,N_8076,N_8372);
nand U8656 (N_8656,N_8286,N_8157);
xnor U8657 (N_8657,N_8305,N_8185);
nor U8658 (N_8658,N_8450,N_8117);
or U8659 (N_8659,N_8120,N_8365);
nor U8660 (N_8660,N_8489,N_8421);
or U8661 (N_8661,N_8111,N_8446);
or U8662 (N_8662,N_8297,N_8470);
nand U8663 (N_8663,N_8191,N_8466);
xnor U8664 (N_8664,N_8317,N_8150);
xor U8665 (N_8665,N_8231,N_8313);
or U8666 (N_8666,N_8051,N_8422);
nand U8667 (N_8667,N_8027,N_8404);
xnor U8668 (N_8668,N_8258,N_8037);
nand U8669 (N_8669,N_8288,N_8411);
nand U8670 (N_8670,N_8024,N_8038);
and U8671 (N_8671,N_8361,N_8350);
nand U8672 (N_8672,N_8164,N_8133);
or U8673 (N_8673,N_8393,N_8201);
nor U8674 (N_8674,N_8232,N_8235);
nand U8675 (N_8675,N_8389,N_8405);
or U8676 (N_8676,N_8138,N_8484);
nand U8677 (N_8677,N_8471,N_8200);
nand U8678 (N_8678,N_8498,N_8139);
or U8679 (N_8679,N_8169,N_8326);
nand U8680 (N_8680,N_8204,N_8495);
or U8681 (N_8681,N_8022,N_8341);
nor U8682 (N_8682,N_8149,N_8067);
and U8683 (N_8683,N_8359,N_8448);
and U8684 (N_8684,N_8202,N_8125);
or U8685 (N_8685,N_8407,N_8192);
nor U8686 (N_8686,N_8480,N_8463);
xor U8687 (N_8687,N_8442,N_8188);
and U8688 (N_8688,N_8251,N_8307);
nor U8689 (N_8689,N_8311,N_8206);
or U8690 (N_8690,N_8161,N_8255);
or U8691 (N_8691,N_8238,N_8145);
and U8692 (N_8692,N_8273,N_8091);
or U8693 (N_8693,N_8434,N_8086);
or U8694 (N_8694,N_8025,N_8438);
xnor U8695 (N_8695,N_8267,N_8375);
nand U8696 (N_8696,N_8423,N_8137);
nand U8697 (N_8697,N_8228,N_8213);
nor U8698 (N_8698,N_8274,N_8395);
nor U8699 (N_8699,N_8482,N_8462);
nand U8700 (N_8700,N_8212,N_8312);
nor U8701 (N_8701,N_8431,N_8416);
nand U8702 (N_8702,N_8113,N_8180);
nor U8703 (N_8703,N_8344,N_8132);
and U8704 (N_8704,N_8084,N_8358);
xnor U8705 (N_8705,N_8314,N_8394);
or U8706 (N_8706,N_8012,N_8173);
nor U8707 (N_8707,N_8473,N_8015);
xor U8708 (N_8708,N_8174,N_8184);
nor U8709 (N_8709,N_8388,N_8122);
or U8710 (N_8710,N_8093,N_8282);
or U8711 (N_8711,N_8237,N_8497);
or U8712 (N_8712,N_8000,N_8453);
xnor U8713 (N_8713,N_8099,N_8320);
nand U8714 (N_8714,N_8017,N_8476);
or U8715 (N_8715,N_8399,N_8033);
nor U8716 (N_8716,N_8127,N_8364);
nor U8717 (N_8717,N_8064,N_8351);
or U8718 (N_8718,N_8444,N_8065);
nor U8719 (N_8719,N_8347,N_8257);
and U8720 (N_8720,N_8021,N_8095);
xor U8721 (N_8721,N_8023,N_8459);
xor U8722 (N_8722,N_8121,N_8042);
nor U8723 (N_8723,N_8290,N_8417);
nand U8724 (N_8724,N_8089,N_8436);
and U8725 (N_8725,N_8043,N_8324);
nor U8726 (N_8726,N_8035,N_8451);
nand U8727 (N_8727,N_8343,N_8186);
nor U8728 (N_8728,N_8469,N_8310);
nand U8729 (N_8729,N_8166,N_8119);
or U8730 (N_8730,N_8321,N_8041);
and U8731 (N_8731,N_8087,N_8155);
nand U8732 (N_8732,N_8264,N_8403);
nand U8733 (N_8733,N_8170,N_8380);
nor U8734 (N_8734,N_8308,N_8088);
or U8735 (N_8735,N_8252,N_8214);
and U8736 (N_8736,N_8356,N_8248);
and U8737 (N_8737,N_8152,N_8455);
nor U8738 (N_8738,N_8492,N_8443);
and U8739 (N_8739,N_8220,N_8070);
nor U8740 (N_8740,N_8261,N_8387);
nor U8741 (N_8741,N_8262,N_8179);
nand U8742 (N_8742,N_8447,N_8167);
or U8743 (N_8743,N_8278,N_8330);
or U8744 (N_8744,N_8243,N_8253);
xnor U8745 (N_8745,N_8362,N_8402);
nor U8746 (N_8746,N_8181,N_8218);
and U8747 (N_8747,N_8224,N_8247);
nor U8748 (N_8748,N_8103,N_8144);
or U8749 (N_8749,N_8397,N_8052);
or U8750 (N_8750,N_8423,N_8139);
or U8751 (N_8751,N_8139,N_8056);
nand U8752 (N_8752,N_8252,N_8349);
or U8753 (N_8753,N_8237,N_8390);
xor U8754 (N_8754,N_8056,N_8329);
and U8755 (N_8755,N_8491,N_8052);
nor U8756 (N_8756,N_8339,N_8135);
xnor U8757 (N_8757,N_8317,N_8300);
nand U8758 (N_8758,N_8094,N_8103);
or U8759 (N_8759,N_8390,N_8377);
nand U8760 (N_8760,N_8424,N_8047);
and U8761 (N_8761,N_8210,N_8229);
nand U8762 (N_8762,N_8178,N_8449);
xnor U8763 (N_8763,N_8009,N_8267);
or U8764 (N_8764,N_8246,N_8358);
xor U8765 (N_8765,N_8357,N_8164);
nor U8766 (N_8766,N_8205,N_8348);
xnor U8767 (N_8767,N_8353,N_8284);
nor U8768 (N_8768,N_8451,N_8464);
xnor U8769 (N_8769,N_8214,N_8189);
nor U8770 (N_8770,N_8116,N_8421);
xor U8771 (N_8771,N_8441,N_8433);
nand U8772 (N_8772,N_8075,N_8465);
xor U8773 (N_8773,N_8316,N_8050);
nor U8774 (N_8774,N_8400,N_8002);
nor U8775 (N_8775,N_8364,N_8231);
xor U8776 (N_8776,N_8109,N_8089);
or U8777 (N_8777,N_8333,N_8128);
nor U8778 (N_8778,N_8131,N_8173);
nand U8779 (N_8779,N_8441,N_8345);
and U8780 (N_8780,N_8235,N_8086);
or U8781 (N_8781,N_8084,N_8396);
xor U8782 (N_8782,N_8369,N_8262);
and U8783 (N_8783,N_8127,N_8163);
nor U8784 (N_8784,N_8161,N_8488);
xnor U8785 (N_8785,N_8464,N_8378);
or U8786 (N_8786,N_8149,N_8211);
or U8787 (N_8787,N_8029,N_8200);
or U8788 (N_8788,N_8372,N_8114);
nand U8789 (N_8789,N_8098,N_8078);
xnor U8790 (N_8790,N_8114,N_8297);
nor U8791 (N_8791,N_8358,N_8365);
nor U8792 (N_8792,N_8251,N_8287);
nand U8793 (N_8793,N_8340,N_8326);
xor U8794 (N_8794,N_8150,N_8064);
and U8795 (N_8795,N_8239,N_8264);
nand U8796 (N_8796,N_8361,N_8476);
nor U8797 (N_8797,N_8319,N_8018);
nor U8798 (N_8798,N_8359,N_8442);
xnor U8799 (N_8799,N_8170,N_8262);
and U8800 (N_8800,N_8274,N_8230);
or U8801 (N_8801,N_8146,N_8223);
or U8802 (N_8802,N_8370,N_8408);
xnor U8803 (N_8803,N_8446,N_8481);
or U8804 (N_8804,N_8486,N_8179);
and U8805 (N_8805,N_8079,N_8096);
xor U8806 (N_8806,N_8380,N_8210);
nor U8807 (N_8807,N_8142,N_8358);
nand U8808 (N_8808,N_8297,N_8318);
and U8809 (N_8809,N_8375,N_8298);
and U8810 (N_8810,N_8280,N_8216);
xnor U8811 (N_8811,N_8273,N_8160);
or U8812 (N_8812,N_8287,N_8168);
nor U8813 (N_8813,N_8179,N_8243);
nand U8814 (N_8814,N_8227,N_8119);
xnor U8815 (N_8815,N_8301,N_8193);
nand U8816 (N_8816,N_8208,N_8249);
nand U8817 (N_8817,N_8330,N_8333);
nand U8818 (N_8818,N_8009,N_8145);
xnor U8819 (N_8819,N_8089,N_8125);
nand U8820 (N_8820,N_8097,N_8188);
or U8821 (N_8821,N_8380,N_8498);
nor U8822 (N_8822,N_8352,N_8379);
nand U8823 (N_8823,N_8446,N_8149);
or U8824 (N_8824,N_8294,N_8218);
and U8825 (N_8825,N_8190,N_8200);
nand U8826 (N_8826,N_8305,N_8453);
and U8827 (N_8827,N_8104,N_8478);
xnor U8828 (N_8828,N_8495,N_8297);
nand U8829 (N_8829,N_8390,N_8196);
or U8830 (N_8830,N_8042,N_8329);
xor U8831 (N_8831,N_8282,N_8394);
xnor U8832 (N_8832,N_8411,N_8184);
or U8833 (N_8833,N_8170,N_8317);
nand U8834 (N_8834,N_8017,N_8228);
nor U8835 (N_8835,N_8394,N_8321);
nand U8836 (N_8836,N_8152,N_8364);
xnor U8837 (N_8837,N_8492,N_8310);
nand U8838 (N_8838,N_8088,N_8057);
xnor U8839 (N_8839,N_8363,N_8425);
xnor U8840 (N_8840,N_8224,N_8327);
and U8841 (N_8841,N_8425,N_8204);
xor U8842 (N_8842,N_8295,N_8418);
xor U8843 (N_8843,N_8033,N_8138);
nor U8844 (N_8844,N_8315,N_8073);
nor U8845 (N_8845,N_8350,N_8258);
and U8846 (N_8846,N_8020,N_8124);
xor U8847 (N_8847,N_8185,N_8380);
nor U8848 (N_8848,N_8297,N_8240);
nand U8849 (N_8849,N_8243,N_8198);
xor U8850 (N_8850,N_8017,N_8026);
nor U8851 (N_8851,N_8209,N_8383);
xnor U8852 (N_8852,N_8154,N_8106);
and U8853 (N_8853,N_8081,N_8029);
nand U8854 (N_8854,N_8269,N_8375);
or U8855 (N_8855,N_8290,N_8344);
nor U8856 (N_8856,N_8133,N_8356);
xnor U8857 (N_8857,N_8118,N_8469);
xor U8858 (N_8858,N_8432,N_8345);
and U8859 (N_8859,N_8384,N_8465);
or U8860 (N_8860,N_8251,N_8076);
or U8861 (N_8861,N_8219,N_8423);
or U8862 (N_8862,N_8108,N_8459);
nor U8863 (N_8863,N_8477,N_8374);
or U8864 (N_8864,N_8296,N_8084);
nor U8865 (N_8865,N_8299,N_8315);
xor U8866 (N_8866,N_8231,N_8014);
and U8867 (N_8867,N_8068,N_8449);
nor U8868 (N_8868,N_8301,N_8434);
or U8869 (N_8869,N_8170,N_8193);
xnor U8870 (N_8870,N_8068,N_8217);
nand U8871 (N_8871,N_8450,N_8305);
nand U8872 (N_8872,N_8332,N_8000);
or U8873 (N_8873,N_8097,N_8026);
and U8874 (N_8874,N_8468,N_8010);
or U8875 (N_8875,N_8149,N_8389);
or U8876 (N_8876,N_8240,N_8029);
and U8877 (N_8877,N_8002,N_8376);
nor U8878 (N_8878,N_8475,N_8106);
xor U8879 (N_8879,N_8400,N_8075);
or U8880 (N_8880,N_8324,N_8335);
or U8881 (N_8881,N_8485,N_8283);
and U8882 (N_8882,N_8440,N_8194);
and U8883 (N_8883,N_8007,N_8376);
nor U8884 (N_8884,N_8377,N_8455);
nor U8885 (N_8885,N_8356,N_8448);
or U8886 (N_8886,N_8267,N_8482);
nand U8887 (N_8887,N_8042,N_8184);
or U8888 (N_8888,N_8462,N_8009);
xnor U8889 (N_8889,N_8438,N_8151);
or U8890 (N_8890,N_8236,N_8165);
or U8891 (N_8891,N_8216,N_8200);
or U8892 (N_8892,N_8201,N_8475);
nand U8893 (N_8893,N_8185,N_8383);
nor U8894 (N_8894,N_8327,N_8357);
and U8895 (N_8895,N_8419,N_8005);
and U8896 (N_8896,N_8060,N_8026);
or U8897 (N_8897,N_8485,N_8003);
or U8898 (N_8898,N_8221,N_8256);
xor U8899 (N_8899,N_8375,N_8364);
or U8900 (N_8900,N_8126,N_8342);
nand U8901 (N_8901,N_8344,N_8175);
or U8902 (N_8902,N_8273,N_8203);
xor U8903 (N_8903,N_8013,N_8318);
and U8904 (N_8904,N_8305,N_8430);
nand U8905 (N_8905,N_8170,N_8275);
or U8906 (N_8906,N_8348,N_8056);
nand U8907 (N_8907,N_8249,N_8420);
or U8908 (N_8908,N_8302,N_8448);
and U8909 (N_8909,N_8203,N_8491);
xnor U8910 (N_8910,N_8113,N_8069);
nand U8911 (N_8911,N_8337,N_8091);
nand U8912 (N_8912,N_8489,N_8459);
or U8913 (N_8913,N_8435,N_8115);
or U8914 (N_8914,N_8289,N_8312);
nor U8915 (N_8915,N_8022,N_8156);
and U8916 (N_8916,N_8298,N_8389);
nor U8917 (N_8917,N_8193,N_8185);
nor U8918 (N_8918,N_8135,N_8043);
nand U8919 (N_8919,N_8209,N_8393);
or U8920 (N_8920,N_8223,N_8359);
or U8921 (N_8921,N_8117,N_8457);
or U8922 (N_8922,N_8040,N_8097);
nor U8923 (N_8923,N_8184,N_8359);
nand U8924 (N_8924,N_8280,N_8461);
nand U8925 (N_8925,N_8301,N_8313);
nor U8926 (N_8926,N_8154,N_8443);
and U8927 (N_8927,N_8290,N_8474);
nor U8928 (N_8928,N_8435,N_8324);
xnor U8929 (N_8929,N_8245,N_8009);
or U8930 (N_8930,N_8472,N_8474);
and U8931 (N_8931,N_8348,N_8102);
nor U8932 (N_8932,N_8199,N_8245);
or U8933 (N_8933,N_8031,N_8203);
or U8934 (N_8934,N_8175,N_8024);
or U8935 (N_8935,N_8173,N_8036);
or U8936 (N_8936,N_8121,N_8207);
nand U8937 (N_8937,N_8373,N_8040);
xnor U8938 (N_8938,N_8178,N_8175);
nor U8939 (N_8939,N_8321,N_8305);
nand U8940 (N_8940,N_8110,N_8109);
nor U8941 (N_8941,N_8092,N_8004);
nand U8942 (N_8942,N_8312,N_8400);
nor U8943 (N_8943,N_8298,N_8021);
or U8944 (N_8944,N_8023,N_8384);
nor U8945 (N_8945,N_8498,N_8443);
nor U8946 (N_8946,N_8184,N_8185);
nand U8947 (N_8947,N_8199,N_8262);
xnor U8948 (N_8948,N_8031,N_8212);
xnor U8949 (N_8949,N_8087,N_8221);
xor U8950 (N_8950,N_8264,N_8023);
and U8951 (N_8951,N_8020,N_8418);
xnor U8952 (N_8952,N_8128,N_8405);
xnor U8953 (N_8953,N_8152,N_8234);
and U8954 (N_8954,N_8467,N_8147);
or U8955 (N_8955,N_8153,N_8381);
nand U8956 (N_8956,N_8340,N_8192);
nor U8957 (N_8957,N_8256,N_8137);
nand U8958 (N_8958,N_8470,N_8380);
nor U8959 (N_8959,N_8049,N_8283);
and U8960 (N_8960,N_8079,N_8062);
nor U8961 (N_8961,N_8206,N_8068);
nand U8962 (N_8962,N_8429,N_8025);
nor U8963 (N_8963,N_8034,N_8455);
nand U8964 (N_8964,N_8253,N_8276);
or U8965 (N_8965,N_8224,N_8049);
or U8966 (N_8966,N_8145,N_8342);
nand U8967 (N_8967,N_8205,N_8017);
nor U8968 (N_8968,N_8353,N_8023);
xor U8969 (N_8969,N_8381,N_8156);
nor U8970 (N_8970,N_8397,N_8445);
nor U8971 (N_8971,N_8110,N_8227);
and U8972 (N_8972,N_8169,N_8391);
nor U8973 (N_8973,N_8096,N_8162);
and U8974 (N_8974,N_8186,N_8423);
and U8975 (N_8975,N_8285,N_8314);
or U8976 (N_8976,N_8139,N_8226);
and U8977 (N_8977,N_8128,N_8248);
xor U8978 (N_8978,N_8189,N_8111);
nor U8979 (N_8979,N_8066,N_8259);
xor U8980 (N_8980,N_8370,N_8416);
nand U8981 (N_8981,N_8077,N_8042);
nor U8982 (N_8982,N_8187,N_8088);
or U8983 (N_8983,N_8335,N_8424);
xnor U8984 (N_8984,N_8053,N_8295);
and U8985 (N_8985,N_8135,N_8390);
and U8986 (N_8986,N_8350,N_8447);
nand U8987 (N_8987,N_8398,N_8242);
and U8988 (N_8988,N_8085,N_8301);
nor U8989 (N_8989,N_8388,N_8209);
nor U8990 (N_8990,N_8421,N_8106);
or U8991 (N_8991,N_8233,N_8072);
xor U8992 (N_8992,N_8264,N_8455);
and U8993 (N_8993,N_8340,N_8071);
nand U8994 (N_8994,N_8264,N_8359);
or U8995 (N_8995,N_8246,N_8008);
nor U8996 (N_8996,N_8380,N_8259);
nor U8997 (N_8997,N_8031,N_8326);
nand U8998 (N_8998,N_8152,N_8439);
or U8999 (N_8999,N_8149,N_8215);
nor U9000 (N_9000,N_8794,N_8502);
and U9001 (N_9001,N_8641,N_8587);
xor U9002 (N_9002,N_8554,N_8520);
or U9003 (N_9003,N_8533,N_8536);
or U9004 (N_9004,N_8698,N_8634);
nor U9005 (N_9005,N_8675,N_8732);
or U9006 (N_9006,N_8576,N_8983);
xnor U9007 (N_9007,N_8611,N_8510);
nor U9008 (N_9008,N_8774,N_8773);
nand U9009 (N_9009,N_8534,N_8710);
and U9010 (N_9010,N_8913,N_8936);
xnor U9011 (N_9011,N_8724,N_8876);
nor U9012 (N_9012,N_8821,N_8800);
xor U9013 (N_9013,N_8903,N_8809);
xor U9014 (N_9014,N_8963,N_8574);
nand U9015 (N_9015,N_8529,N_8575);
or U9016 (N_9016,N_8926,N_8530);
nand U9017 (N_9017,N_8967,N_8531);
nor U9018 (N_9018,N_8812,N_8814);
nor U9019 (N_9019,N_8831,N_8981);
xor U9020 (N_9020,N_8965,N_8894);
xnor U9021 (N_9021,N_8638,N_8598);
nand U9022 (N_9022,N_8793,N_8838);
nand U9023 (N_9023,N_8766,N_8852);
nand U9024 (N_9024,N_8892,N_8708);
and U9025 (N_9025,N_8617,N_8545);
and U9026 (N_9026,N_8860,N_8760);
xor U9027 (N_9027,N_8781,N_8777);
and U9028 (N_9028,N_8655,N_8986);
and U9029 (N_9029,N_8570,N_8900);
nand U9030 (N_9030,N_8719,N_8539);
or U9031 (N_9031,N_8842,N_8512);
nor U9032 (N_9032,N_8627,N_8779);
or U9033 (N_9033,N_8948,N_8807);
xnor U9034 (N_9034,N_8928,N_8863);
and U9035 (N_9035,N_8845,N_8820);
nor U9036 (N_9036,N_8739,N_8889);
nor U9037 (N_9037,N_8635,N_8680);
and U9038 (N_9038,N_8735,N_8717);
nand U9039 (N_9039,N_8548,N_8910);
and U9040 (N_9040,N_8853,N_8954);
nand U9041 (N_9041,N_8683,N_8591);
nor U9042 (N_9042,N_8718,N_8955);
nand U9043 (N_9043,N_8991,N_8897);
or U9044 (N_9044,N_8553,N_8677);
and U9045 (N_9045,N_8870,N_8504);
xnor U9046 (N_9046,N_8513,N_8972);
or U9047 (N_9047,N_8788,N_8790);
nor U9048 (N_9048,N_8632,N_8583);
or U9049 (N_9049,N_8526,N_8743);
or U9050 (N_9050,N_8841,N_8557);
or U9051 (N_9051,N_8979,N_8989);
nor U9052 (N_9052,N_8949,N_8924);
nand U9053 (N_9053,N_8857,N_8537);
xor U9054 (N_9054,N_8658,N_8975);
or U9055 (N_9055,N_8685,N_8668);
nor U9056 (N_9056,N_8599,N_8618);
nor U9057 (N_9057,N_8572,N_8604);
nor U9058 (N_9058,N_8856,N_8808);
nand U9059 (N_9059,N_8763,N_8843);
xnor U9060 (N_9060,N_8940,N_8945);
xnor U9061 (N_9061,N_8784,N_8912);
xor U9062 (N_9062,N_8996,N_8562);
xnor U9063 (N_9063,N_8902,N_8801);
nand U9064 (N_9064,N_8916,N_8561);
nor U9065 (N_9065,N_8911,N_8959);
or U9066 (N_9066,N_8585,N_8818);
nor U9067 (N_9067,N_8580,N_8589);
xnor U9068 (N_9068,N_8528,N_8799);
nor U9069 (N_9069,N_8721,N_8614);
and U9070 (N_9070,N_8725,N_8508);
or U9071 (N_9071,N_8559,N_8689);
nand U9072 (N_9072,N_8802,N_8759);
xnor U9073 (N_9073,N_8540,N_8934);
xnor U9074 (N_9074,N_8817,N_8563);
and U9075 (N_9075,N_8697,N_8824);
nor U9076 (N_9076,N_8908,N_8551);
and U9077 (N_9077,N_8958,N_8874);
or U9078 (N_9078,N_8560,N_8961);
or U9079 (N_9079,N_8659,N_8869);
nand U9080 (N_9080,N_8704,N_8726);
nor U9081 (N_9081,N_8693,N_8935);
xnor U9082 (N_9082,N_8883,N_8568);
and U9083 (N_9083,N_8806,N_8674);
xor U9084 (N_9084,N_8650,N_8640);
and U9085 (N_9085,N_8798,N_8645);
or U9086 (N_9086,N_8905,N_8501);
or U9087 (N_9087,N_8612,N_8714);
nand U9088 (N_9088,N_8858,N_8608);
or U9089 (N_9089,N_8519,N_8823);
nand U9090 (N_9090,N_8931,N_8851);
or U9091 (N_9091,N_8663,N_8613);
nand U9092 (N_9092,N_8930,N_8951);
or U9093 (N_9093,N_8847,N_8919);
xor U9094 (N_9094,N_8867,N_8648);
xnor U9095 (N_9095,N_8722,N_8741);
and U9096 (N_9096,N_8918,N_8630);
nand U9097 (N_9097,N_8923,N_8982);
nor U9098 (N_9098,N_8690,N_8767);
nand U9099 (N_9099,N_8571,N_8597);
xor U9100 (N_9100,N_8855,N_8768);
or U9101 (N_9101,N_8973,N_8866);
nor U9102 (N_9102,N_8652,N_8826);
nand U9103 (N_9103,N_8672,N_8624);
nand U9104 (N_9104,N_8661,N_8749);
or U9105 (N_9105,N_8832,N_8946);
nor U9106 (N_9106,N_8871,N_8816);
nor U9107 (N_9107,N_8771,N_8525);
nand U9108 (N_9108,N_8815,N_8976);
and U9109 (N_9109,N_8968,N_8854);
nor U9110 (N_9110,N_8915,N_8738);
xor U9111 (N_9111,N_8730,N_8873);
nand U9112 (N_9112,N_8601,N_8720);
nor U9113 (N_9113,N_8932,N_8657);
xor U9114 (N_9114,N_8836,N_8699);
or U9115 (N_9115,N_8558,N_8682);
or U9116 (N_9116,N_8942,N_8647);
xor U9117 (N_9117,N_8746,N_8977);
xor U9118 (N_9118,N_8628,N_8830);
xor U9119 (N_9119,N_8792,N_8791);
nand U9120 (N_9120,N_8990,N_8503);
or U9121 (N_9121,N_8745,N_8750);
nand U9122 (N_9122,N_8998,N_8547);
or U9123 (N_9123,N_8939,N_8925);
nand U9124 (N_9124,N_8765,N_8639);
xnor U9125 (N_9125,N_8950,N_8862);
and U9126 (N_9126,N_8868,N_8881);
or U9127 (N_9127,N_8783,N_8829);
nor U9128 (N_9128,N_8667,N_8596);
nor U9129 (N_9129,N_8888,N_8579);
or U9130 (N_9130,N_8654,N_8549);
nor U9131 (N_9131,N_8723,N_8676);
xor U9132 (N_9132,N_8679,N_8516);
or U9133 (N_9133,N_8715,N_8593);
or U9134 (N_9134,N_8891,N_8736);
nor U9135 (N_9135,N_8764,N_8899);
or U9136 (N_9136,N_8620,N_8625);
and U9137 (N_9137,N_8567,N_8956);
or U9138 (N_9138,N_8615,N_8651);
xor U9139 (N_9139,N_8947,N_8546);
nor U9140 (N_9140,N_8592,N_8692);
and U9141 (N_9141,N_8653,N_8671);
or U9142 (N_9142,N_8517,N_8872);
and U9143 (N_9143,N_8619,N_8805);
xnor U9144 (N_9144,N_8957,N_8590);
nor U9145 (N_9145,N_8769,N_8681);
nand U9146 (N_9146,N_8751,N_8636);
nand U9147 (N_9147,N_8929,N_8938);
or U9148 (N_9148,N_8544,N_8865);
nor U9149 (N_9149,N_8895,N_8952);
nand U9150 (N_9150,N_8688,N_8914);
nor U9151 (N_9151,N_8556,N_8626);
nor U9152 (N_9152,N_8787,N_8660);
nand U9153 (N_9153,N_8886,N_8518);
and U9154 (N_9154,N_8758,N_8532);
and U9155 (N_9155,N_8993,N_8974);
xor U9156 (N_9156,N_8844,N_8756);
or U9157 (N_9157,N_8696,N_8941);
nand U9158 (N_9158,N_8511,N_8964);
or U9159 (N_9159,N_8837,N_8581);
and U9160 (N_9160,N_8500,N_8670);
nand U9161 (N_9161,N_8971,N_8728);
xnor U9162 (N_9162,N_8775,N_8877);
and U9163 (N_9163,N_8541,N_8884);
and U9164 (N_9164,N_8762,N_8637);
xnor U9165 (N_9165,N_8827,N_8550);
nor U9166 (N_9166,N_8631,N_8804);
xor U9167 (N_9167,N_8789,N_8514);
xor U9168 (N_9168,N_8896,N_8780);
and U9169 (N_9169,N_8879,N_8864);
nand U9170 (N_9170,N_8524,N_8980);
nand U9171 (N_9171,N_8684,N_8582);
xnor U9172 (N_9172,N_8573,N_8810);
or U9173 (N_9173,N_8776,N_8995);
nor U9174 (N_9174,N_8729,N_8921);
xnor U9175 (N_9175,N_8621,N_8623);
nor U9176 (N_9176,N_8609,N_8709);
nor U9177 (N_9177,N_8778,N_8988);
xor U9178 (N_9178,N_8761,N_8564);
nand U9179 (N_9179,N_8909,N_8507);
xor U9180 (N_9180,N_8966,N_8822);
nand U9181 (N_9181,N_8882,N_8835);
nand U9182 (N_9182,N_8633,N_8937);
xnor U9183 (N_9183,N_8744,N_8848);
xor U9184 (N_9184,N_8523,N_8811);
xor U9185 (N_9185,N_8907,N_8713);
and U9186 (N_9186,N_8859,N_8849);
xnor U9187 (N_9187,N_8782,N_8694);
and U9188 (N_9188,N_8754,N_8839);
nand U9189 (N_9189,N_8642,N_8691);
and U9190 (N_9190,N_8953,N_8646);
or U9191 (N_9191,N_8880,N_8555);
nand U9192 (N_9192,N_8786,N_8616);
and U9193 (N_9193,N_8706,N_8994);
xor U9194 (N_9194,N_8662,N_8747);
nand U9195 (N_9195,N_8890,N_8740);
or U9196 (N_9196,N_8927,N_8875);
nor U9197 (N_9197,N_8878,N_8673);
and U9198 (N_9198,N_8584,N_8538);
nand U9199 (N_9199,N_8944,N_8701);
xor U9200 (N_9200,N_8960,N_8666);
or U9201 (N_9201,N_8695,N_8885);
or U9202 (N_9202,N_8622,N_8594);
xnor U9203 (N_9203,N_8700,N_8686);
and U9204 (N_9204,N_8610,N_8705);
or U9205 (N_9205,N_8734,N_8898);
and U9206 (N_9206,N_8906,N_8578);
nor U9207 (N_9207,N_8833,N_8987);
or U9208 (N_9208,N_8997,N_8606);
nor U9209 (N_9209,N_8552,N_8542);
nand U9210 (N_9210,N_8969,N_8569);
nor U9211 (N_9211,N_8737,N_8796);
and U9212 (N_9212,N_8985,N_8887);
nor U9213 (N_9213,N_8840,N_8703);
xor U9214 (N_9214,N_8566,N_8861);
and U9215 (N_9215,N_8772,N_8669);
or U9216 (N_9216,N_8819,N_8588);
xor U9217 (N_9217,N_8962,N_8521);
nor U9218 (N_9218,N_8595,N_8602);
or U9219 (N_9219,N_8515,N_8731);
nor U9220 (N_9220,N_8943,N_8505);
and U9221 (N_9221,N_8586,N_8733);
and U9222 (N_9222,N_8711,N_8753);
nor U9223 (N_9223,N_8978,N_8577);
xor U9224 (N_9224,N_8752,N_8607);
or U9225 (N_9225,N_8649,N_8797);
nor U9226 (N_9226,N_8527,N_8825);
nor U9227 (N_9227,N_8506,N_8970);
nor U9228 (N_9228,N_8678,N_8727);
and U9229 (N_9229,N_8893,N_8643);
and U9230 (N_9230,N_8846,N_8933);
and U9231 (N_9231,N_8702,N_8707);
and U9232 (N_9232,N_8665,N_8834);
nand U9233 (N_9233,N_8803,N_8644);
and U9234 (N_9234,N_8917,N_8664);
and U9235 (N_9235,N_8901,N_8656);
nand U9236 (N_9236,N_8687,N_8757);
and U9237 (N_9237,N_8795,N_8600);
and U9238 (N_9238,N_8565,N_8828);
xor U9239 (N_9239,N_8920,N_8850);
or U9240 (N_9240,N_8770,N_8712);
nor U9241 (N_9241,N_8629,N_8813);
nor U9242 (N_9242,N_8742,N_8785);
nor U9243 (N_9243,N_8999,N_8748);
and U9244 (N_9244,N_8605,N_8755);
nand U9245 (N_9245,N_8984,N_8543);
or U9246 (N_9246,N_8716,N_8509);
nor U9247 (N_9247,N_8522,N_8992);
nand U9248 (N_9248,N_8603,N_8535);
and U9249 (N_9249,N_8922,N_8904);
or U9250 (N_9250,N_8790,N_8669);
and U9251 (N_9251,N_8687,N_8565);
and U9252 (N_9252,N_8694,N_8675);
nor U9253 (N_9253,N_8563,N_8975);
xnor U9254 (N_9254,N_8912,N_8658);
xor U9255 (N_9255,N_8627,N_8889);
or U9256 (N_9256,N_8842,N_8850);
nor U9257 (N_9257,N_8801,N_8738);
nand U9258 (N_9258,N_8545,N_8793);
nand U9259 (N_9259,N_8641,N_8645);
xor U9260 (N_9260,N_8861,N_8839);
or U9261 (N_9261,N_8689,N_8510);
or U9262 (N_9262,N_8644,N_8606);
xnor U9263 (N_9263,N_8920,N_8977);
or U9264 (N_9264,N_8640,N_8878);
xor U9265 (N_9265,N_8667,N_8612);
and U9266 (N_9266,N_8617,N_8531);
or U9267 (N_9267,N_8552,N_8952);
nor U9268 (N_9268,N_8772,N_8558);
or U9269 (N_9269,N_8675,N_8585);
xnor U9270 (N_9270,N_8539,N_8632);
nor U9271 (N_9271,N_8875,N_8973);
xor U9272 (N_9272,N_8880,N_8965);
and U9273 (N_9273,N_8656,N_8882);
nor U9274 (N_9274,N_8757,N_8818);
nor U9275 (N_9275,N_8618,N_8600);
xnor U9276 (N_9276,N_8503,N_8917);
nor U9277 (N_9277,N_8917,N_8670);
and U9278 (N_9278,N_8555,N_8837);
nand U9279 (N_9279,N_8646,N_8805);
nor U9280 (N_9280,N_8921,N_8568);
xor U9281 (N_9281,N_8710,N_8623);
xor U9282 (N_9282,N_8569,N_8845);
xnor U9283 (N_9283,N_8614,N_8680);
and U9284 (N_9284,N_8720,N_8702);
nand U9285 (N_9285,N_8777,N_8713);
xor U9286 (N_9286,N_8818,N_8821);
nor U9287 (N_9287,N_8559,N_8757);
nor U9288 (N_9288,N_8704,N_8834);
or U9289 (N_9289,N_8793,N_8961);
nor U9290 (N_9290,N_8792,N_8732);
xnor U9291 (N_9291,N_8848,N_8835);
or U9292 (N_9292,N_8918,N_8859);
or U9293 (N_9293,N_8828,N_8714);
or U9294 (N_9294,N_8755,N_8668);
nor U9295 (N_9295,N_8994,N_8582);
nand U9296 (N_9296,N_8888,N_8690);
nand U9297 (N_9297,N_8917,N_8997);
nand U9298 (N_9298,N_8559,N_8657);
and U9299 (N_9299,N_8511,N_8794);
and U9300 (N_9300,N_8912,N_8621);
or U9301 (N_9301,N_8797,N_8688);
xor U9302 (N_9302,N_8587,N_8694);
nand U9303 (N_9303,N_8672,N_8539);
or U9304 (N_9304,N_8657,N_8508);
and U9305 (N_9305,N_8730,N_8968);
xor U9306 (N_9306,N_8979,N_8682);
nor U9307 (N_9307,N_8607,N_8768);
nor U9308 (N_9308,N_8828,N_8640);
or U9309 (N_9309,N_8796,N_8616);
or U9310 (N_9310,N_8583,N_8610);
or U9311 (N_9311,N_8905,N_8855);
or U9312 (N_9312,N_8691,N_8689);
or U9313 (N_9313,N_8587,N_8977);
xnor U9314 (N_9314,N_8999,N_8806);
and U9315 (N_9315,N_8618,N_8780);
xnor U9316 (N_9316,N_8938,N_8987);
or U9317 (N_9317,N_8589,N_8556);
nand U9318 (N_9318,N_8914,N_8901);
xnor U9319 (N_9319,N_8670,N_8962);
or U9320 (N_9320,N_8926,N_8844);
or U9321 (N_9321,N_8752,N_8969);
and U9322 (N_9322,N_8952,N_8863);
nand U9323 (N_9323,N_8823,N_8664);
xnor U9324 (N_9324,N_8737,N_8608);
and U9325 (N_9325,N_8822,N_8756);
or U9326 (N_9326,N_8966,N_8511);
nand U9327 (N_9327,N_8872,N_8637);
xnor U9328 (N_9328,N_8608,N_8968);
nor U9329 (N_9329,N_8971,N_8818);
and U9330 (N_9330,N_8820,N_8612);
xnor U9331 (N_9331,N_8954,N_8936);
nor U9332 (N_9332,N_8857,N_8601);
and U9333 (N_9333,N_8549,N_8797);
nand U9334 (N_9334,N_8645,N_8824);
xnor U9335 (N_9335,N_8707,N_8961);
and U9336 (N_9336,N_8795,N_8676);
nor U9337 (N_9337,N_8765,N_8940);
and U9338 (N_9338,N_8824,N_8794);
nand U9339 (N_9339,N_8992,N_8890);
nand U9340 (N_9340,N_8667,N_8740);
and U9341 (N_9341,N_8863,N_8718);
nand U9342 (N_9342,N_8511,N_8524);
nand U9343 (N_9343,N_8531,N_8748);
nor U9344 (N_9344,N_8918,N_8698);
and U9345 (N_9345,N_8521,N_8952);
and U9346 (N_9346,N_8730,N_8762);
nor U9347 (N_9347,N_8951,N_8603);
nand U9348 (N_9348,N_8581,N_8752);
xnor U9349 (N_9349,N_8890,N_8620);
xnor U9350 (N_9350,N_8929,N_8556);
xnor U9351 (N_9351,N_8693,N_8980);
and U9352 (N_9352,N_8836,N_8665);
xnor U9353 (N_9353,N_8763,N_8726);
nor U9354 (N_9354,N_8963,N_8906);
and U9355 (N_9355,N_8720,N_8963);
nor U9356 (N_9356,N_8921,N_8995);
and U9357 (N_9357,N_8689,N_8777);
and U9358 (N_9358,N_8500,N_8862);
xor U9359 (N_9359,N_8969,N_8502);
nand U9360 (N_9360,N_8599,N_8577);
nor U9361 (N_9361,N_8547,N_8508);
xnor U9362 (N_9362,N_8521,N_8981);
and U9363 (N_9363,N_8588,N_8711);
or U9364 (N_9364,N_8701,N_8886);
xor U9365 (N_9365,N_8833,N_8606);
nor U9366 (N_9366,N_8528,N_8514);
or U9367 (N_9367,N_8575,N_8634);
xnor U9368 (N_9368,N_8501,N_8929);
nand U9369 (N_9369,N_8798,N_8680);
or U9370 (N_9370,N_8562,N_8592);
or U9371 (N_9371,N_8515,N_8939);
or U9372 (N_9372,N_8654,N_8536);
nor U9373 (N_9373,N_8868,N_8912);
or U9374 (N_9374,N_8754,N_8971);
or U9375 (N_9375,N_8865,N_8853);
nand U9376 (N_9376,N_8920,N_8588);
nand U9377 (N_9377,N_8714,N_8699);
and U9378 (N_9378,N_8848,N_8906);
nand U9379 (N_9379,N_8866,N_8790);
nand U9380 (N_9380,N_8899,N_8689);
xnor U9381 (N_9381,N_8694,N_8684);
or U9382 (N_9382,N_8825,N_8998);
nor U9383 (N_9383,N_8603,N_8550);
nand U9384 (N_9384,N_8991,N_8600);
or U9385 (N_9385,N_8561,N_8674);
or U9386 (N_9386,N_8952,N_8584);
nand U9387 (N_9387,N_8844,N_8803);
and U9388 (N_9388,N_8646,N_8718);
xor U9389 (N_9389,N_8627,N_8600);
nor U9390 (N_9390,N_8755,N_8695);
or U9391 (N_9391,N_8710,N_8997);
xor U9392 (N_9392,N_8696,N_8781);
or U9393 (N_9393,N_8977,N_8763);
nor U9394 (N_9394,N_8550,N_8773);
nor U9395 (N_9395,N_8708,N_8823);
nand U9396 (N_9396,N_8766,N_8944);
nand U9397 (N_9397,N_8712,N_8644);
nor U9398 (N_9398,N_8714,N_8927);
xnor U9399 (N_9399,N_8728,N_8882);
or U9400 (N_9400,N_8722,N_8986);
or U9401 (N_9401,N_8590,N_8779);
nor U9402 (N_9402,N_8846,N_8740);
nor U9403 (N_9403,N_8786,N_8582);
xor U9404 (N_9404,N_8578,N_8800);
nor U9405 (N_9405,N_8534,N_8753);
nand U9406 (N_9406,N_8880,N_8755);
xor U9407 (N_9407,N_8880,N_8692);
nand U9408 (N_9408,N_8818,N_8884);
nor U9409 (N_9409,N_8519,N_8606);
nand U9410 (N_9410,N_8620,N_8904);
nand U9411 (N_9411,N_8827,N_8836);
xnor U9412 (N_9412,N_8739,N_8503);
nor U9413 (N_9413,N_8639,N_8619);
nand U9414 (N_9414,N_8891,N_8827);
and U9415 (N_9415,N_8628,N_8543);
xor U9416 (N_9416,N_8727,N_8625);
nor U9417 (N_9417,N_8989,N_8780);
xor U9418 (N_9418,N_8932,N_8586);
nand U9419 (N_9419,N_8642,N_8639);
nand U9420 (N_9420,N_8635,N_8911);
and U9421 (N_9421,N_8910,N_8526);
xnor U9422 (N_9422,N_8520,N_8936);
xor U9423 (N_9423,N_8660,N_8504);
xor U9424 (N_9424,N_8698,N_8898);
nor U9425 (N_9425,N_8796,N_8853);
and U9426 (N_9426,N_8962,N_8830);
and U9427 (N_9427,N_8631,N_8862);
and U9428 (N_9428,N_8580,N_8555);
xor U9429 (N_9429,N_8516,N_8511);
xnor U9430 (N_9430,N_8911,N_8971);
nand U9431 (N_9431,N_8882,N_8687);
nand U9432 (N_9432,N_8688,N_8751);
or U9433 (N_9433,N_8797,N_8884);
nor U9434 (N_9434,N_8851,N_8526);
or U9435 (N_9435,N_8517,N_8522);
or U9436 (N_9436,N_8812,N_8733);
or U9437 (N_9437,N_8834,N_8824);
or U9438 (N_9438,N_8816,N_8669);
nand U9439 (N_9439,N_8913,N_8874);
or U9440 (N_9440,N_8828,N_8755);
xor U9441 (N_9441,N_8717,N_8772);
or U9442 (N_9442,N_8582,N_8650);
nand U9443 (N_9443,N_8816,N_8847);
xnor U9444 (N_9444,N_8603,N_8753);
nor U9445 (N_9445,N_8978,N_8633);
and U9446 (N_9446,N_8912,N_8932);
xnor U9447 (N_9447,N_8865,N_8602);
and U9448 (N_9448,N_8915,N_8545);
or U9449 (N_9449,N_8970,N_8550);
or U9450 (N_9450,N_8906,N_8523);
xor U9451 (N_9451,N_8893,N_8724);
nand U9452 (N_9452,N_8627,N_8641);
nor U9453 (N_9453,N_8703,N_8566);
nand U9454 (N_9454,N_8861,N_8525);
xnor U9455 (N_9455,N_8709,N_8796);
nor U9456 (N_9456,N_8501,N_8970);
nor U9457 (N_9457,N_8824,N_8663);
or U9458 (N_9458,N_8947,N_8635);
nand U9459 (N_9459,N_8905,N_8749);
and U9460 (N_9460,N_8917,N_8930);
nor U9461 (N_9461,N_8685,N_8955);
and U9462 (N_9462,N_8957,N_8607);
and U9463 (N_9463,N_8667,N_8593);
nor U9464 (N_9464,N_8914,N_8609);
and U9465 (N_9465,N_8503,N_8784);
or U9466 (N_9466,N_8852,N_8512);
xnor U9467 (N_9467,N_8629,N_8751);
nor U9468 (N_9468,N_8979,N_8897);
and U9469 (N_9469,N_8930,N_8698);
xor U9470 (N_9470,N_8687,N_8999);
nor U9471 (N_9471,N_8692,N_8847);
or U9472 (N_9472,N_8553,N_8640);
and U9473 (N_9473,N_8780,N_8810);
and U9474 (N_9474,N_8786,N_8990);
xnor U9475 (N_9475,N_8811,N_8505);
nand U9476 (N_9476,N_8558,N_8746);
or U9477 (N_9477,N_8958,N_8776);
nand U9478 (N_9478,N_8855,N_8876);
nor U9479 (N_9479,N_8884,N_8849);
nand U9480 (N_9480,N_8708,N_8662);
nor U9481 (N_9481,N_8646,N_8959);
and U9482 (N_9482,N_8989,N_8575);
nand U9483 (N_9483,N_8878,N_8735);
nand U9484 (N_9484,N_8509,N_8512);
nand U9485 (N_9485,N_8747,N_8641);
or U9486 (N_9486,N_8915,N_8786);
and U9487 (N_9487,N_8865,N_8579);
nor U9488 (N_9488,N_8503,N_8508);
and U9489 (N_9489,N_8652,N_8947);
nand U9490 (N_9490,N_8981,N_8523);
xor U9491 (N_9491,N_8948,N_8920);
or U9492 (N_9492,N_8811,N_8851);
nand U9493 (N_9493,N_8737,N_8580);
nor U9494 (N_9494,N_8698,N_8645);
xnor U9495 (N_9495,N_8718,N_8501);
or U9496 (N_9496,N_8536,N_8977);
or U9497 (N_9497,N_8807,N_8622);
nor U9498 (N_9498,N_8818,N_8540);
and U9499 (N_9499,N_8669,N_8836);
nor U9500 (N_9500,N_9322,N_9463);
xor U9501 (N_9501,N_9013,N_9006);
and U9502 (N_9502,N_9487,N_9007);
xor U9503 (N_9503,N_9295,N_9077);
nor U9504 (N_9504,N_9204,N_9044);
nor U9505 (N_9505,N_9366,N_9473);
nand U9506 (N_9506,N_9241,N_9373);
nand U9507 (N_9507,N_9239,N_9298);
nor U9508 (N_9508,N_9047,N_9120);
and U9509 (N_9509,N_9059,N_9079);
and U9510 (N_9510,N_9187,N_9213);
nor U9511 (N_9511,N_9105,N_9174);
and U9512 (N_9512,N_9289,N_9001);
nor U9513 (N_9513,N_9210,N_9016);
and U9514 (N_9514,N_9107,N_9499);
nor U9515 (N_9515,N_9308,N_9029);
and U9516 (N_9516,N_9349,N_9458);
nand U9517 (N_9517,N_9165,N_9233);
nor U9518 (N_9518,N_9171,N_9246);
xnor U9519 (N_9519,N_9387,N_9113);
or U9520 (N_9520,N_9492,N_9043);
and U9521 (N_9521,N_9097,N_9066);
nor U9522 (N_9522,N_9136,N_9234);
and U9523 (N_9523,N_9443,N_9448);
xor U9524 (N_9524,N_9347,N_9130);
and U9525 (N_9525,N_9414,N_9276);
nor U9526 (N_9526,N_9074,N_9369);
xor U9527 (N_9527,N_9133,N_9202);
and U9528 (N_9528,N_9467,N_9312);
xnor U9529 (N_9529,N_9140,N_9109);
nor U9530 (N_9530,N_9098,N_9423);
or U9531 (N_9531,N_9309,N_9178);
nand U9532 (N_9532,N_9303,N_9407);
or U9533 (N_9533,N_9194,N_9403);
xnor U9534 (N_9534,N_9155,N_9485);
or U9535 (N_9535,N_9424,N_9033);
or U9536 (N_9536,N_9360,N_9015);
or U9537 (N_9537,N_9406,N_9383);
or U9538 (N_9538,N_9146,N_9264);
xnor U9539 (N_9539,N_9455,N_9083);
and U9540 (N_9540,N_9161,N_9252);
and U9541 (N_9541,N_9453,N_9248);
nor U9542 (N_9542,N_9129,N_9454);
xnor U9543 (N_9543,N_9353,N_9126);
xor U9544 (N_9544,N_9104,N_9476);
and U9545 (N_9545,N_9498,N_9311);
nor U9546 (N_9546,N_9219,N_9314);
or U9547 (N_9547,N_9346,N_9052);
nand U9548 (N_9548,N_9305,N_9231);
nand U9549 (N_9549,N_9223,N_9087);
nand U9550 (N_9550,N_9249,N_9188);
nand U9551 (N_9551,N_9474,N_9283);
nor U9552 (N_9552,N_9095,N_9090);
or U9553 (N_9553,N_9148,N_9002);
nand U9554 (N_9554,N_9365,N_9419);
xnor U9555 (N_9555,N_9153,N_9030);
or U9556 (N_9556,N_9464,N_9429);
or U9557 (N_9557,N_9340,N_9091);
xnor U9558 (N_9558,N_9193,N_9441);
nor U9559 (N_9559,N_9116,N_9280);
nand U9560 (N_9560,N_9056,N_9386);
and U9561 (N_9561,N_9118,N_9106);
nand U9562 (N_9562,N_9125,N_9151);
nor U9563 (N_9563,N_9137,N_9494);
nand U9564 (N_9564,N_9160,N_9124);
nor U9565 (N_9565,N_9380,N_9310);
nand U9566 (N_9566,N_9356,N_9232);
nor U9567 (N_9567,N_9082,N_9325);
and U9568 (N_9568,N_9085,N_9027);
or U9569 (N_9569,N_9479,N_9243);
xor U9570 (N_9570,N_9430,N_9497);
xnor U9571 (N_9571,N_9076,N_9335);
nor U9572 (N_9572,N_9245,N_9110);
xnor U9573 (N_9573,N_9446,N_9028);
xnor U9574 (N_9574,N_9049,N_9483);
and U9575 (N_9575,N_9230,N_9175);
nand U9576 (N_9576,N_9238,N_9435);
and U9577 (N_9577,N_9196,N_9010);
nor U9578 (N_9578,N_9149,N_9127);
nor U9579 (N_9579,N_9209,N_9332);
nor U9580 (N_9580,N_9361,N_9381);
or U9581 (N_9581,N_9061,N_9054);
xnor U9582 (N_9582,N_9117,N_9050);
nand U9583 (N_9583,N_9400,N_9447);
and U9584 (N_9584,N_9438,N_9046);
or U9585 (N_9585,N_9319,N_9168);
and U9586 (N_9586,N_9024,N_9431);
nor U9587 (N_9587,N_9269,N_9330);
and U9588 (N_9588,N_9073,N_9271);
and U9589 (N_9589,N_9362,N_9313);
nor U9590 (N_9590,N_9177,N_9031);
xnor U9591 (N_9591,N_9456,N_9432);
and U9592 (N_9592,N_9385,N_9329);
xor U9593 (N_9593,N_9358,N_9009);
nor U9594 (N_9594,N_9201,N_9156);
or U9595 (N_9595,N_9008,N_9382);
or U9596 (N_9596,N_9281,N_9062);
nor U9597 (N_9597,N_9328,N_9285);
nor U9598 (N_9598,N_9299,N_9375);
or U9599 (N_9599,N_9142,N_9203);
nand U9600 (N_9600,N_9162,N_9482);
xor U9601 (N_9601,N_9057,N_9401);
and U9602 (N_9602,N_9461,N_9226);
nor U9603 (N_9603,N_9191,N_9420);
nand U9604 (N_9604,N_9284,N_9014);
or U9605 (N_9605,N_9068,N_9434);
and U9606 (N_9606,N_9439,N_9197);
or U9607 (N_9607,N_9186,N_9063);
and U9608 (N_9608,N_9416,N_9247);
xnor U9609 (N_9609,N_9147,N_9268);
xnor U9610 (N_9610,N_9158,N_9290);
xnor U9611 (N_9611,N_9317,N_9286);
or U9612 (N_9612,N_9352,N_9261);
or U9613 (N_9613,N_9025,N_9108);
nand U9614 (N_9614,N_9145,N_9364);
nor U9615 (N_9615,N_9111,N_9170);
nand U9616 (N_9616,N_9055,N_9327);
and U9617 (N_9617,N_9410,N_9451);
and U9618 (N_9618,N_9023,N_9192);
and U9619 (N_9619,N_9300,N_9042);
nand U9620 (N_9620,N_9331,N_9215);
and U9621 (N_9621,N_9176,N_9377);
or U9622 (N_9622,N_9051,N_9307);
nor U9623 (N_9623,N_9277,N_9363);
or U9624 (N_9624,N_9379,N_9112);
xnor U9625 (N_9625,N_9172,N_9240);
nand U9626 (N_9626,N_9189,N_9397);
nor U9627 (N_9627,N_9152,N_9442);
or U9628 (N_9628,N_9368,N_9088);
or U9629 (N_9629,N_9121,N_9408);
nand U9630 (N_9630,N_9235,N_9257);
and U9631 (N_9631,N_9294,N_9093);
or U9632 (N_9632,N_9081,N_9086);
nor U9633 (N_9633,N_9478,N_9452);
and U9634 (N_9634,N_9418,N_9012);
xnor U9635 (N_9635,N_9341,N_9004);
or U9636 (N_9636,N_9164,N_9018);
or U9637 (N_9637,N_9396,N_9384);
xnor U9638 (N_9638,N_9065,N_9465);
and U9639 (N_9639,N_9200,N_9437);
nor U9640 (N_9640,N_9282,N_9242);
nor U9641 (N_9641,N_9302,N_9466);
nor U9642 (N_9642,N_9357,N_9251);
nand U9643 (N_9643,N_9236,N_9274);
xor U9644 (N_9644,N_9469,N_9490);
nor U9645 (N_9645,N_9391,N_9222);
or U9646 (N_9646,N_9496,N_9132);
nor U9647 (N_9647,N_9395,N_9011);
xnor U9648 (N_9648,N_9321,N_9278);
xor U9649 (N_9649,N_9260,N_9253);
nand U9650 (N_9650,N_9250,N_9019);
nor U9651 (N_9651,N_9224,N_9398);
and U9652 (N_9652,N_9344,N_9157);
or U9653 (N_9653,N_9199,N_9123);
nand U9654 (N_9654,N_9343,N_9181);
xnor U9655 (N_9655,N_9198,N_9316);
xnor U9656 (N_9656,N_9428,N_9338);
xnor U9657 (N_9657,N_9399,N_9275);
nand U9658 (N_9658,N_9184,N_9333);
nor U9659 (N_9659,N_9486,N_9037);
nand U9660 (N_9660,N_9342,N_9413);
nor U9661 (N_9661,N_9128,N_9064);
xor U9662 (N_9662,N_9425,N_9354);
or U9663 (N_9663,N_9227,N_9229);
nand U9664 (N_9664,N_9334,N_9388);
nand U9665 (N_9665,N_9339,N_9060);
nor U9666 (N_9666,N_9449,N_9103);
nor U9667 (N_9667,N_9460,N_9135);
nand U9668 (N_9668,N_9491,N_9134);
or U9669 (N_9669,N_9071,N_9070);
nand U9670 (N_9670,N_9468,N_9297);
or U9671 (N_9671,N_9211,N_9315);
nand U9672 (N_9672,N_9143,N_9237);
nand U9673 (N_9673,N_9348,N_9069);
xor U9674 (N_9674,N_9472,N_9003);
xnor U9675 (N_9675,N_9220,N_9345);
xnor U9676 (N_9676,N_9207,N_9167);
xor U9677 (N_9677,N_9034,N_9102);
xor U9678 (N_9678,N_9304,N_9411);
nor U9679 (N_9679,N_9350,N_9115);
or U9680 (N_9680,N_9444,N_9254);
xnor U9681 (N_9681,N_9475,N_9417);
and U9682 (N_9682,N_9067,N_9228);
or U9683 (N_9683,N_9150,N_9267);
xnor U9684 (N_9684,N_9038,N_9021);
nor U9685 (N_9685,N_9405,N_9216);
xor U9686 (N_9686,N_9263,N_9427);
xnor U9687 (N_9687,N_9041,N_9481);
or U9688 (N_9688,N_9206,N_9078);
xnor U9689 (N_9689,N_9218,N_9489);
nor U9690 (N_9690,N_9372,N_9119);
nand U9691 (N_9691,N_9470,N_9371);
or U9692 (N_9692,N_9291,N_9415);
nor U9693 (N_9693,N_9495,N_9017);
nor U9694 (N_9694,N_9421,N_9075);
or U9695 (N_9695,N_9306,N_9445);
xnor U9696 (N_9696,N_9180,N_9426);
nor U9697 (N_9697,N_9324,N_9390);
and U9698 (N_9698,N_9058,N_9273);
and U9699 (N_9699,N_9114,N_9040);
nand U9700 (N_9700,N_9412,N_9409);
nand U9701 (N_9701,N_9032,N_9138);
nor U9702 (N_9702,N_9378,N_9208);
nor U9703 (N_9703,N_9000,N_9096);
nor U9704 (N_9704,N_9488,N_9402);
xor U9705 (N_9705,N_9272,N_9089);
and U9706 (N_9706,N_9320,N_9053);
or U9707 (N_9707,N_9292,N_9100);
xnor U9708 (N_9708,N_9005,N_9185);
xor U9709 (N_9709,N_9287,N_9440);
or U9710 (N_9710,N_9163,N_9462);
xor U9711 (N_9711,N_9262,N_9326);
and U9712 (N_9712,N_9255,N_9159);
or U9713 (N_9713,N_9288,N_9144);
nand U9714 (N_9714,N_9036,N_9139);
xnor U9715 (N_9715,N_9190,N_9183);
xor U9716 (N_9716,N_9039,N_9020);
nand U9717 (N_9717,N_9480,N_9336);
and U9718 (N_9718,N_9045,N_9221);
and U9719 (N_9719,N_9394,N_9265);
xnor U9720 (N_9720,N_9154,N_9195);
nor U9721 (N_9721,N_9173,N_9022);
xnor U9722 (N_9722,N_9259,N_9099);
or U9723 (N_9723,N_9244,N_9182);
nand U9724 (N_9724,N_9084,N_9217);
nor U9725 (N_9725,N_9166,N_9393);
nand U9726 (N_9726,N_9459,N_9374);
nand U9727 (N_9727,N_9258,N_9072);
or U9728 (N_9728,N_9293,N_9131);
xor U9729 (N_9729,N_9389,N_9318);
and U9730 (N_9730,N_9323,N_9484);
nor U9731 (N_9731,N_9205,N_9080);
nor U9732 (N_9732,N_9094,N_9279);
nand U9733 (N_9733,N_9214,N_9048);
nor U9734 (N_9734,N_9337,N_9433);
xor U9735 (N_9735,N_9179,N_9392);
nand U9736 (N_9736,N_9471,N_9035);
and U9737 (N_9737,N_9404,N_9266);
or U9738 (N_9738,N_9301,N_9225);
nand U9739 (N_9739,N_9422,N_9457);
xnor U9740 (N_9740,N_9101,N_9141);
nand U9741 (N_9741,N_9355,N_9270);
or U9742 (N_9742,N_9256,N_9493);
nor U9743 (N_9743,N_9122,N_9296);
and U9744 (N_9744,N_9477,N_9367);
or U9745 (N_9745,N_9370,N_9092);
or U9746 (N_9746,N_9359,N_9376);
nor U9747 (N_9747,N_9026,N_9436);
nor U9748 (N_9748,N_9212,N_9351);
xnor U9749 (N_9749,N_9169,N_9450);
or U9750 (N_9750,N_9227,N_9048);
xnor U9751 (N_9751,N_9014,N_9228);
or U9752 (N_9752,N_9435,N_9377);
xnor U9753 (N_9753,N_9356,N_9442);
or U9754 (N_9754,N_9202,N_9027);
and U9755 (N_9755,N_9265,N_9335);
and U9756 (N_9756,N_9103,N_9346);
xor U9757 (N_9757,N_9195,N_9345);
and U9758 (N_9758,N_9168,N_9205);
nor U9759 (N_9759,N_9492,N_9112);
and U9760 (N_9760,N_9302,N_9132);
nand U9761 (N_9761,N_9142,N_9407);
and U9762 (N_9762,N_9177,N_9191);
nor U9763 (N_9763,N_9410,N_9114);
and U9764 (N_9764,N_9441,N_9057);
nor U9765 (N_9765,N_9483,N_9019);
xnor U9766 (N_9766,N_9458,N_9070);
or U9767 (N_9767,N_9397,N_9495);
nand U9768 (N_9768,N_9346,N_9199);
or U9769 (N_9769,N_9348,N_9409);
nand U9770 (N_9770,N_9346,N_9499);
and U9771 (N_9771,N_9227,N_9434);
xor U9772 (N_9772,N_9226,N_9312);
nand U9773 (N_9773,N_9114,N_9434);
or U9774 (N_9774,N_9150,N_9252);
nand U9775 (N_9775,N_9462,N_9123);
xor U9776 (N_9776,N_9418,N_9000);
and U9777 (N_9777,N_9149,N_9264);
xnor U9778 (N_9778,N_9203,N_9061);
nor U9779 (N_9779,N_9208,N_9045);
nand U9780 (N_9780,N_9274,N_9364);
or U9781 (N_9781,N_9318,N_9024);
xor U9782 (N_9782,N_9037,N_9341);
nand U9783 (N_9783,N_9126,N_9377);
or U9784 (N_9784,N_9312,N_9002);
and U9785 (N_9785,N_9349,N_9303);
xnor U9786 (N_9786,N_9229,N_9278);
nor U9787 (N_9787,N_9027,N_9054);
nor U9788 (N_9788,N_9132,N_9289);
or U9789 (N_9789,N_9458,N_9488);
xnor U9790 (N_9790,N_9433,N_9252);
nand U9791 (N_9791,N_9166,N_9461);
or U9792 (N_9792,N_9474,N_9429);
nand U9793 (N_9793,N_9134,N_9111);
xnor U9794 (N_9794,N_9252,N_9393);
nor U9795 (N_9795,N_9335,N_9107);
or U9796 (N_9796,N_9187,N_9259);
and U9797 (N_9797,N_9233,N_9113);
nand U9798 (N_9798,N_9206,N_9397);
nor U9799 (N_9799,N_9264,N_9094);
xor U9800 (N_9800,N_9448,N_9353);
nand U9801 (N_9801,N_9179,N_9344);
or U9802 (N_9802,N_9152,N_9433);
xnor U9803 (N_9803,N_9352,N_9495);
nor U9804 (N_9804,N_9143,N_9332);
or U9805 (N_9805,N_9217,N_9363);
and U9806 (N_9806,N_9135,N_9299);
xor U9807 (N_9807,N_9206,N_9283);
nor U9808 (N_9808,N_9271,N_9178);
xor U9809 (N_9809,N_9434,N_9158);
nand U9810 (N_9810,N_9345,N_9127);
nor U9811 (N_9811,N_9235,N_9271);
and U9812 (N_9812,N_9143,N_9185);
nor U9813 (N_9813,N_9059,N_9187);
nor U9814 (N_9814,N_9288,N_9228);
nor U9815 (N_9815,N_9339,N_9184);
or U9816 (N_9816,N_9421,N_9141);
and U9817 (N_9817,N_9126,N_9432);
xnor U9818 (N_9818,N_9320,N_9077);
nor U9819 (N_9819,N_9460,N_9267);
nor U9820 (N_9820,N_9353,N_9085);
or U9821 (N_9821,N_9249,N_9220);
xor U9822 (N_9822,N_9320,N_9252);
or U9823 (N_9823,N_9219,N_9347);
nor U9824 (N_9824,N_9059,N_9338);
and U9825 (N_9825,N_9276,N_9484);
nor U9826 (N_9826,N_9407,N_9069);
or U9827 (N_9827,N_9152,N_9217);
nand U9828 (N_9828,N_9432,N_9382);
nor U9829 (N_9829,N_9027,N_9310);
and U9830 (N_9830,N_9227,N_9185);
xnor U9831 (N_9831,N_9009,N_9428);
and U9832 (N_9832,N_9297,N_9017);
nand U9833 (N_9833,N_9350,N_9285);
nor U9834 (N_9834,N_9323,N_9274);
nand U9835 (N_9835,N_9057,N_9232);
nand U9836 (N_9836,N_9117,N_9090);
or U9837 (N_9837,N_9255,N_9198);
or U9838 (N_9838,N_9421,N_9403);
xnor U9839 (N_9839,N_9164,N_9231);
xor U9840 (N_9840,N_9454,N_9174);
nor U9841 (N_9841,N_9020,N_9422);
nor U9842 (N_9842,N_9111,N_9186);
nand U9843 (N_9843,N_9004,N_9168);
nand U9844 (N_9844,N_9052,N_9152);
nor U9845 (N_9845,N_9277,N_9237);
nor U9846 (N_9846,N_9357,N_9179);
or U9847 (N_9847,N_9217,N_9282);
and U9848 (N_9848,N_9082,N_9483);
and U9849 (N_9849,N_9199,N_9375);
xnor U9850 (N_9850,N_9083,N_9080);
xor U9851 (N_9851,N_9266,N_9323);
nor U9852 (N_9852,N_9020,N_9136);
xor U9853 (N_9853,N_9149,N_9104);
xor U9854 (N_9854,N_9160,N_9184);
and U9855 (N_9855,N_9497,N_9231);
xor U9856 (N_9856,N_9115,N_9474);
or U9857 (N_9857,N_9123,N_9198);
nand U9858 (N_9858,N_9459,N_9011);
nand U9859 (N_9859,N_9078,N_9115);
nor U9860 (N_9860,N_9291,N_9067);
nor U9861 (N_9861,N_9295,N_9399);
xor U9862 (N_9862,N_9353,N_9374);
nor U9863 (N_9863,N_9204,N_9103);
and U9864 (N_9864,N_9459,N_9406);
nor U9865 (N_9865,N_9229,N_9224);
nand U9866 (N_9866,N_9046,N_9462);
and U9867 (N_9867,N_9111,N_9363);
or U9868 (N_9868,N_9120,N_9062);
nor U9869 (N_9869,N_9149,N_9254);
or U9870 (N_9870,N_9183,N_9339);
xnor U9871 (N_9871,N_9013,N_9157);
xor U9872 (N_9872,N_9123,N_9281);
xnor U9873 (N_9873,N_9081,N_9326);
xnor U9874 (N_9874,N_9430,N_9452);
and U9875 (N_9875,N_9237,N_9093);
nor U9876 (N_9876,N_9268,N_9026);
nor U9877 (N_9877,N_9479,N_9132);
nand U9878 (N_9878,N_9326,N_9385);
nor U9879 (N_9879,N_9449,N_9391);
or U9880 (N_9880,N_9045,N_9212);
and U9881 (N_9881,N_9133,N_9099);
nor U9882 (N_9882,N_9379,N_9385);
or U9883 (N_9883,N_9266,N_9210);
nor U9884 (N_9884,N_9197,N_9413);
xnor U9885 (N_9885,N_9290,N_9016);
and U9886 (N_9886,N_9133,N_9154);
and U9887 (N_9887,N_9361,N_9269);
nor U9888 (N_9888,N_9359,N_9377);
or U9889 (N_9889,N_9275,N_9350);
nor U9890 (N_9890,N_9270,N_9384);
nand U9891 (N_9891,N_9408,N_9246);
nand U9892 (N_9892,N_9402,N_9168);
nand U9893 (N_9893,N_9062,N_9386);
nor U9894 (N_9894,N_9237,N_9128);
nand U9895 (N_9895,N_9244,N_9141);
xnor U9896 (N_9896,N_9267,N_9061);
nand U9897 (N_9897,N_9376,N_9026);
nor U9898 (N_9898,N_9435,N_9341);
nor U9899 (N_9899,N_9288,N_9486);
nand U9900 (N_9900,N_9361,N_9000);
xnor U9901 (N_9901,N_9157,N_9364);
nand U9902 (N_9902,N_9197,N_9171);
nor U9903 (N_9903,N_9308,N_9476);
xnor U9904 (N_9904,N_9454,N_9092);
xnor U9905 (N_9905,N_9486,N_9071);
nor U9906 (N_9906,N_9269,N_9121);
or U9907 (N_9907,N_9102,N_9298);
xnor U9908 (N_9908,N_9239,N_9122);
nand U9909 (N_9909,N_9192,N_9443);
nor U9910 (N_9910,N_9065,N_9212);
and U9911 (N_9911,N_9323,N_9242);
and U9912 (N_9912,N_9086,N_9393);
and U9913 (N_9913,N_9259,N_9060);
nand U9914 (N_9914,N_9066,N_9372);
and U9915 (N_9915,N_9181,N_9173);
nor U9916 (N_9916,N_9278,N_9203);
nor U9917 (N_9917,N_9031,N_9004);
and U9918 (N_9918,N_9362,N_9173);
xor U9919 (N_9919,N_9074,N_9193);
xnor U9920 (N_9920,N_9013,N_9281);
nand U9921 (N_9921,N_9185,N_9288);
nand U9922 (N_9922,N_9455,N_9177);
xor U9923 (N_9923,N_9315,N_9128);
and U9924 (N_9924,N_9031,N_9396);
and U9925 (N_9925,N_9296,N_9000);
nand U9926 (N_9926,N_9133,N_9185);
and U9927 (N_9927,N_9352,N_9311);
and U9928 (N_9928,N_9451,N_9474);
and U9929 (N_9929,N_9183,N_9304);
nand U9930 (N_9930,N_9167,N_9112);
nand U9931 (N_9931,N_9167,N_9124);
and U9932 (N_9932,N_9428,N_9191);
nand U9933 (N_9933,N_9370,N_9068);
and U9934 (N_9934,N_9241,N_9315);
or U9935 (N_9935,N_9268,N_9105);
or U9936 (N_9936,N_9012,N_9049);
and U9937 (N_9937,N_9198,N_9332);
xnor U9938 (N_9938,N_9135,N_9073);
or U9939 (N_9939,N_9446,N_9124);
and U9940 (N_9940,N_9469,N_9182);
nor U9941 (N_9941,N_9013,N_9341);
or U9942 (N_9942,N_9022,N_9446);
and U9943 (N_9943,N_9062,N_9127);
or U9944 (N_9944,N_9471,N_9194);
and U9945 (N_9945,N_9098,N_9374);
nand U9946 (N_9946,N_9253,N_9499);
nand U9947 (N_9947,N_9011,N_9102);
or U9948 (N_9948,N_9297,N_9400);
nor U9949 (N_9949,N_9481,N_9164);
and U9950 (N_9950,N_9125,N_9481);
and U9951 (N_9951,N_9456,N_9276);
xor U9952 (N_9952,N_9260,N_9147);
nand U9953 (N_9953,N_9375,N_9159);
and U9954 (N_9954,N_9155,N_9486);
nand U9955 (N_9955,N_9463,N_9253);
or U9956 (N_9956,N_9375,N_9222);
nor U9957 (N_9957,N_9458,N_9267);
and U9958 (N_9958,N_9222,N_9426);
nand U9959 (N_9959,N_9233,N_9130);
and U9960 (N_9960,N_9344,N_9089);
nand U9961 (N_9961,N_9379,N_9487);
and U9962 (N_9962,N_9404,N_9305);
nor U9963 (N_9963,N_9456,N_9484);
xnor U9964 (N_9964,N_9012,N_9263);
and U9965 (N_9965,N_9289,N_9308);
and U9966 (N_9966,N_9272,N_9017);
xor U9967 (N_9967,N_9113,N_9448);
nand U9968 (N_9968,N_9454,N_9109);
nand U9969 (N_9969,N_9438,N_9238);
nand U9970 (N_9970,N_9434,N_9028);
nand U9971 (N_9971,N_9433,N_9033);
nand U9972 (N_9972,N_9100,N_9494);
and U9973 (N_9973,N_9472,N_9284);
and U9974 (N_9974,N_9216,N_9331);
or U9975 (N_9975,N_9375,N_9351);
or U9976 (N_9976,N_9020,N_9052);
xor U9977 (N_9977,N_9174,N_9175);
xnor U9978 (N_9978,N_9285,N_9172);
and U9979 (N_9979,N_9223,N_9064);
nand U9980 (N_9980,N_9330,N_9074);
nand U9981 (N_9981,N_9116,N_9337);
and U9982 (N_9982,N_9295,N_9009);
and U9983 (N_9983,N_9191,N_9089);
xnor U9984 (N_9984,N_9460,N_9265);
nor U9985 (N_9985,N_9440,N_9197);
xnor U9986 (N_9986,N_9434,N_9177);
and U9987 (N_9987,N_9454,N_9031);
or U9988 (N_9988,N_9352,N_9295);
nor U9989 (N_9989,N_9123,N_9010);
or U9990 (N_9990,N_9173,N_9256);
and U9991 (N_9991,N_9451,N_9167);
nor U9992 (N_9992,N_9236,N_9164);
and U9993 (N_9993,N_9306,N_9308);
nor U9994 (N_9994,N_9025,N_9258);
xor U9995 (N_9995,N_9356,N_9039);
nor U9996 (N_9996,N_9172,N_9116);
xnor U9997 (N_9997,N_9099,N_9206);
nand U9998 (N_9998,N_9299,N_9234);
nor U9999 (N_9999,N_9143,N_9274);
or U10000 (N_10000,N_9505,N_9642);
nand U10001 (N_10001,N_9523,N_9992);
xor U10002 (N_10002,N_9987,N_9805);
and U10003 (N_10003,N_9792,N_9915);
and U10004 (N_10004,N_9968,N_9732);
or U10005 (N_10005,N_9519,N_9582);
nor U10006 (N_10006,N_9555,N_9541);
and U10007 (N_10007,N_9532,N_9881);
and U10008 (N_10008,N_9895,N_9695);
and U10009 (N_10009,N_9800,N_9727);
nand U10010 (N_10010,N_9528,N_9509);
nor U10011 (N_10011,N_9650,N_9852);
xnor U10012 (N_10012,N_9565,N_9859);
xor U10013 (N_10013,N_9539,N_9783);
and U10014 (N_10014,N_9659,N_9671);
nand U10015 (N_10015,N_9600,N_9752);
nor U10016 (N_10016,N_9696,N_9715);
nand U10017 (N_10017,N_9963,N_9922);
xnor U10018 (N_10018,N_9633,N_9973);
nand U10019 (N_10019,N_9798,N_9885);
xor U10020 (N_10020,N_9556,N_9807);
nand U10021 (N_10021,N_9803,N_9607);
xor U10022 (N_10022,N_9831,N_9662);
xnor U10023 (N_10023,N_9971,N_9668);
nor U10024 (N_10024,N_9572,N_9513);
nand U10025 (N_10025,N_9909,N_9744);
and U10026 (N_10026,N_9994,N_9848);
or U10027 (N_10027,N_9530,N_9670);
nor U10028 (N_10028,N_9873,N_9941);
and U10029 (N_10029,N_9967,N_9820);
nor U10030 (N_10030,N_9988,N_9746);
xnor U10031 (N_10031,N_9954,N_9797);
nand U10032 (N_10032,N_9969,N_9779);
xnor U10033 (N_10033,N_9767,N_9830);
xor U10034 (N_10034,N_9776,N_9773);
or U10035 (N_10035,N_9620,N_9894);
or U10036 (N_10036,N_9691,N_9764);
xor U10037 (N_10037,N_9561,N_9645);
nor U10038 (N_10038,N_9828,N_9960);
xnor U10039 (N_10039,N_9599,N_9958);
and U10040 (N_10040,N_9636,N_9566);
or U10041 (N_10041,N_9775,N_9839);
nor U10042 (N_10042,N_9931,N_9819);
xnor U10043 (N_10043,N_9726,N_9974);
or U10044 (N_10044,N_9921,N_9524);
nor U10045 (N_10045,N_9601,N_9578);
nor U10046 (N_10046,N_9900,N_9658);
and U10047 (N_10047,N_9758,N_9871);
or U10048 (N_10048,N_9625,N_9853);
xnor U10049 (N_10049,N_9869,N_9778);
nor U10050 (N_10050,N_9718,N_9863);
xnor U10051 (N_10051,N_9739,N_9694);
or U10052 (N_10052,N_9693,N_9680);
or U10053 (N_10053,N_9836,N_9711);
and U10054 (N_10054,N_9978,N_9554);
nand U10055 (N_10055,N_9510,N_9932);
and U10056 (N_10056,N_9849,N_9651);
and U10057 (N_10057,N_9784,N_9857);
or U10058 (N_10058,N_9868,N_9677);
or U10059 (N_10059,N_9598,N_9725);
xnor U10060 (N_10060,N_9708,N_9924);
or U10061 (N_10061,N_9794,N_9516);
nor U10062 (N_10062,N_9647,N_9602);
nor U10063 (N_10063,N_9957,N_9701);
nor U10064 (N_10064,N_9928,N_9705);
or U10065 (N_10065,N_9951,N_9989);
nand U10066 (N_10066,N_9638,N_9581);
nand U10067 (N_10067,N_9901,N_9750);
or U10068 (N_10068,N_9997,N_9891);
nand U10069 (N_10069,N_9765,N_9904);
xor U10070 (N_10070,N_9938,N_9747);
nand U10071 (N_10071,N_9802,N_9741);
nor U10072 (N_10072,N_9583,N_9856);
and U10073 (N_10073,N_9615,N_9772);
nor U10074 (N_10074,N_9824,N_9619);
nand U10075 (N_10075,N_9759,N_9501);
and U10076 (N_10076,N_9919,N_9858);
xnor U10077 (N_10077,N_9986,N_9793);
and U10078 (N_10078,N_9686,N_9811);
and U10079 (N_10079,N_9500,N_9514);
or U10080 (N_10080,N_9672,N_9875);
and U10081 (N_10081,N_9883,N_9712);
or U10082 (N_10082,N_9588,N_9506);
xnor U10083 (N_10083,N_9751,N_9704);
nand U10084 (N_10084,N_9795,N_9740);
nand U10085 (N_10085,N_9676,N_9801);
or U10086 (N_10086,N_9757,N_9503);
and U10087 (N_10087,N_9641,N_9903);
and U10088 (N_10088,N_9799,N_9700);
and U10089 (N_10089,N_9564,N_9804);
nor U10090 (N_10090,N_9590,N_9780);
and U10091 (N_10091,N_9735,N_9667);
nand U10092 (N_10092,N_9866,N_9923);
or U10093 (N_10093,N_9605,N_9716);
nor U10094 (N_10094,N_9550,N_9526);
or U10095 (N_10095,N_9635,N_9844);
xnor U10096 (N_10096,N_9766,N_9594);
or U10097 (N_10097,N_9703,N_9511);
or U10098 (N_10098,N_9892,N_9774);
nor U10099 (N_10099,N_9655,N_9610);
nor U10100 (N_10100,N_9925,N_9587);
and U10101 (N_10101,N_9535,N_9628);
xnor U10102 (N_10102,N_9557,N_9586);
nor U10103 (N_10103,N_9812,N_9936);
and U10104 (N_10104,N_9548,N_9674);
nor U10105 (N_10105,N_9684,N_9529);
and U10106 (N_10106,N_9991,N_9768);
xnor U10107 (N_10107,N_9675,N_9983);
nor U10108 (N_10108,N_9592,N_9567);
xnor U10109 (N_10109,N_9558,N_9930);
and U10110 (N_10110,N_9714,N_9818);
xnor U10111 (N_10111,N_9907,N_9884);
or U10112 (N_10112,N_9787,N_9770);
xnor U10113 (N_10113,N_9935,N_9872);
or U10114 (N_10114,N_9545,N_9597);
or U10115 (N_10115,N_9549,N_9748);
and U10116 (N_10116,N_9946,N_9851);
or U10117 (N_10117,N_9874,N_9916);
or U10118 (N_10118,N_9827,N_9710);
xor U10119 (N_10119,N_9737,N_9813);
and U10120 (N_10120,N_9707,N_9591);
xor U10121 (N_10121,N_9634,N_9660);
nand U10122 (N_10122,N_9666,N_9721);
nand U10123 (N_10123,N_9534,N_9860);
and U10124 (N_10124,N_9926,N_9604);
or U10125 (N_10125,N_9880,N_9664);
or U10126 (N_10126,N_9611,N_9882);
nor U10127 (N_10127,N_9966,N_9563);
xnor U10128 (N_10128,N_9639,N_9956);
xnor U10129 (N_10129,N_9728,N_9790);
or U10130 (N_10130,N_9908,N_9829);
and U10131 (N_10131,N_9842,N_9576);
or U10132 (N_10132,N_9621,N_9624);
nand U10133 (N_10133,N_9914,N_9981);
nand U10134 (N_10134,N_9669,N_9652);
nor U10135 (N_10135,N_9681,N_9911);
and U10136 (N_10136,N_9888,N_9878);
nor U10137 (N_10137,N_9846,N_9761);
nand U10138 (N_10138,N_9937,N_9618);
and U10139 (N_10139,N_9609,N_9833);
and U10140 (N_10140,N_9723,N_9940);
and U10141 (N_10141,N_9781,N_9815);
nor U10142 (N_10142,N_9569,N_9816);
nand U10143 (N_10143,N_9623,N_9673);
and U10144 (N_10144,N_9622,N_9870);
and U10145 (N_10145,N_9814,N_9709);
nor U10146 (N_10146,N_9985,N_9596);
nor U10147 (N_10147,N_9823,N_9947);
or U10148 (N_10148,N_9945,N_9975);
nor U10149 (N_10149,N_9791,N_9887);
xnor U10150 (N_10150,N_9905,N_9595);
xnor U10151 (N_10151,N_9754,N_9826);
xor U10152 (N_10152,N_9632,N_9537);
nor U10153 (N_10153,N_9729,N_9984);
and U10154 (N_10154,N_9962,N_9589);
nor U10155 (N_10155,N_9838,N_9612);
and U10156 (N_10156,N_9736,N_9522);
and U10157 (N_10157,N_9631,N_9899);
nand U10158 (N_10158,N_9690,N_9515);
nand U10159 (N_10159,N_9629,N_9982);
or U10160 (N_10160,N_9993,N_9553);
nand U10161 (N_10161,N_9998,N_9979);
or U10162 (N_10162,N_9850,N_9720);
nand U10163 (N_10163,N_9749,N_9538);
or U10164 (N_10164,N_9996,N_9646);
nand U10165 (N_10165,N_9689,N_9533);
xor U10166 (N_10166,N_9665,N_9810);
and U10167 (N_10167,N_9678,N_9719);
and U10168 (N_10168,N_9745,N_9679);
and U10169 (N_10169,N_9573,N_9755);
nand U10170 (N_10170,N_9656,N_9698);
and U10171 (N_10171,N_9939,N_9724);
nor U10172 (N_10172,N_9976,N_9855);
or U10173 (N_10173,N_9902,N_9661);
nand U10174 (N_10174,N_9950,N_9722);
or U10175 (N_10175,N_9806,N_9697);
and U10176 (N_10176,N_9593,N_9913);
nand U10177 (N_10177,N_9990,N_9699);
nand U10178 (N_10178,N_9644,N_9949);
xor U10179 (N_10179,N_9817,N_9942);
or U10180 (N_10180,N_9630,N_9585);
or U10181 (N_10181,N_9575,N_9972);
or U10182 (N_10182,N_9733,N_9648);
and U10183 (N_10183,N_9822,N_9753);
or U10184 (N_10184,N_9730,N_9626);
or U10185 (N_10185,N_9713,N_9959);
xor U10186 (N_10186,N_9613,N_9542);
nor U10187 (N_10187,N_9687,N_9692);
nand U10188 (N_10188,N_9889,N_9517);
or U10189 (N_10189,N_9837,N_9653);
or U10190 (N_10190,N_9518,N_9847);
nor U10191 (N_10191,N_9521,N_9546);
or U10192 (N_10192,N_9685,N_9527);
nand U10193 (N_10193,N_9504,N_9841);
and U10194 (N_10194,N_9877,N_9912);
nand U10195 (N_10195,N_9682,N_9965);
or U10196 (N_10196,N_9760,N_9608);
nor U10197 (N_10197,N_9890,N_9640);
nor U10198 (N_10198,N_9570,N_9865);
or U10199 (N_10199,N_9821,N_9977);
nand U10200 (N_10200,N_9657,N_9688);
nor U10201 (N_10201,N_9525,N_9577);
nand U10202 (N_10202,N_9502,N_9627);
nor U10203 (N_10203,N_9616,N_9603);
and U10204 (N_10204,N_9835,N_9559);
or U10205 (N_10205,N_9649,N_9920);
nand U10206 (N_10206,N_9756,N_9910);
xor U10207 (N_10207,N_9796,N_9832);
and U10208 (N_10208,N_9606,N_9785);
and U10209 (N_10209,N_9929,N_9825);
or U10210 (N_10210,N_9540,N_9717);
nand U10211 (N_10211,N_9584,N_9867);
and U10212 (N_10212,N_9614,N_9933);
nor U10213 (N_10213,N_9562,N_9543);
nor U10214 (N_10214,N_9637,N_9980);
or U10215 (N_10215,N_9560,N_9917);
nor U10216 (N_10216,N_9876,N_9777);
xnor U10217 (N_10217,N_9571,N_9970);
nor U10218 (N_10218,N_9843,N_9731);
or U10219 (N_10219,N_9568,N_9995);
or U10220 (N_10220,N_9654,N_9808);
or U10221 (N_10221,N_9771,N_9944);
and U10222 (N_10222,N_9961,N_9508);
xnor U10223 (N_10223,N_9788,N_9663);
or U10224 (N_10224,N_9918,N_9789);
or U10225 (N_10225,N_9617,N_9964);
and U10226 (N_10226,N_9955,N_9706);
xor U10227 (N_10227,N_9574,N_9782);
xnor U10228 (N_10228,N_9762,N_9531);
and U10229 (N_10229,N_9943,N_9734);
or U10230 (N_10230,N_9547,N_9551);
nand U10231 (N_10231,N_9906,N_9927);
nand U10232 (N_10232,N_9552,N_9742);
xor U10233 (N_10233,N_9854,N_9999);
and U10234 (N_10234,N_9769,N_9897);
xnor U10235 (N_10235,N_9738,N_9952);
or U10236 (N_10236,N_9896,N_9845);
xnor U10237 (N_10237,N_9763,N_9879);
nand U10238 (N_10238,N_9683,N_9743);
nand U10239 (N_10239,N_9507,N_9953);
nor U10240 (N_10240,N_9948,N_9536);
and U10241 (N_10241,N_9702,N_9580);
and U10242 (N_10242,N_9544,N_9643);
and U10243 (N_10243,N_9786,N_9934);
nand U10244 (N_10244,N_9579,N_9520);
and U10245 (N_10245,N_9893,N_9861);
nand U10246 (N_10246,N_9809,N_9834);
or U10247 (N_10247,N_9862,N_9840);
nand U10248 (N_10248,N_9512,N_9864);
and U10249 (N_10249,N_9886,N_9898);
xnor U10250 (N_10250,N_9836,N_9966);
and U10251 (N_10251,N_9863,N_9868);
xor U10252 (N_10252,N_9578,N_9706);
and U10253 (N_10253,N_9534,N_9577);
nor U10254 (N_10254,N_9525,N_9876);
and U10255 (N_10255,N_9668,N_9744);
or U10256 (N_10256,N_9948,N_9608);
nand U10257 (N_10257,N_9522,N_9833);
nor U10258 (N_10258,N_9889,N_9684);
nor U10259 (N_10259,N_9946,N_9938);
nand U10260 (N_10260,N_9651,N_9794);
xor U10261 (N_10261,N_9911,N_9762);
xnor U10262 (N_10262,N_9619,N_9572);
xnor U10263 (N_10263,N_9763,N_9622);
nand U10264 (N_10264,N_9783,N_9528);
or U10265 (N_10265,N_9623,N_9789);
xor U10266 (N_10266,N_9527,N_9808);
and U10267 (N_10267,N_9772,N_9544);
or U10268 (N_10268,N_9856,N_9670);
xor U10269 (N_10269,N_9560,N_9922);
or U10270 (N_10270,N_9564,N_9941);
and U10271 (N_10271,N_9956,N_9976);
xor U10272 (N_10272,N_9710,N_9711);
nand U10273 (N_10273,N_9669,N_9985);
or U10274 (N_10274,N_9529,N_9543);
xnor U10275 (N_10275,N_9699,N_9893);
nand U10276 (N_10276,N_9955,N_9931);
and U10277 (N_10277,N_9850,N_9597);
xnor U10278 (N_10278,N_9981,N_9705);
or U10279 (N_10279,N_9823,N_9613);
or U10280 (N_10280,N_9968,N_9784);
xnor U10281 (N_10281,N_9735,N_9865);
nand U10282 (N_10282,N_9786,N_9874);
xor U10283 (N_10283,N_9935,N_9808);
nor U10284 (N_10284,N_9830,N_9992);
nor U10285 (N_10285,N_9588,N_9873);
or U10286 (N_10286,N_9528,N_9919);
xnor U10287 (N_10287,N_9611,N_9517);
xor U10288 (N_10288,N_9911,N_9746);
or U10289 (N_10289,N_9981,N_9880);
nand U10290 (N_10290,N_9893,N_9609);
or U10291 (N_10291,N_9711,N_9865);
xor U10292 (N_10292,N_9788,N_9987);
nor U10293 (N_10293,N_9872,N_9645);
and U10294 (N_10294,N_9800,N_9606);
nand U10295 (N_10295,N_9873,N_9906);
and U10296 (N_10296,N_9818,N_9724);
or U10297 (N_10297,N_9798,N_9590);
nand U10298 (N_10298,N_9814,N_9589);
xnor U10299 (N_10299,N_9713,N_9655);
or U10300 (N_10300,N_9735,N_9599);
and U10301 (N_10301,N_9776,N_9598);
or U10302 (N_10302,N_9787,N_9861);
or U10303 (N_10303,N_9621,N_9550);
xnor U10304 (N_10304,N_9823,N_9688);
or U10305 (N_10305,N_9669,N_9806);
nand U10306 (N_10306,N_9562,N_9712);
xor U10307 (N_10307,N_9690,N_9736);
or U10308 (N_10308,N_9596,N_9707);
xnor U10309 (N_10309,N_9547,N_9590);
nor U10310 (N_10310,N_9602,N_9827);
xnor U10311 (N_10311,N_9706,N_9571);
xnor U10312 (N_10312,N_9801,N_9747);
and U10313 (N_10313,N_9609,N_9658);
or U10314 (N_10314,N_9813,N_9559);
xor U10315 (N_10315,N_9874,N_9979);
or U10316 (N_10316,N_9656,N_9940);
or U10317 (N_10317,N_9700,N_9958);
nand U10318 (N_10318,N_9938,N_9727);
and U10319 (N_10319,N_9984,N_9750);
xnor U10320 (N_10320,N_9658,N_9885);
or U10321 (N_10321,N_9564,N_9850);
or U10322 (N_10322,N_9759,N_9748);
xor U10323 (N_10323,N_9888,N_9640);
xnor U10324 (N_10324,N_9521,N_9646);
or U10325 (N_10325,N_9658,N_9551);
xnor U10326 (N_10326,N_9824,N_9685);
xnor U10327 (N_10327,N_9844,N_9849);
or U10328 (N_10328,N_9901,N_9587);
and U10329 (N_10329,N_9792,N_9647);
nor U10330 (N_10330,N_9590,N_9764);
nor U10331 (N_10331,N_9724,N_9990);
xnor U10332 (N_10332,N_9816,N_9792);
nand U10333 (N_10333,N_9649,N_9526);
nor U10334 (N_10334,N_9930,N_9800);
or U10335 (N_10335,N_9913,N_9654);
or U10336 (N_10336,N_9915,N_9910);
and U10337 (N_10337,N_9951,N_9903);
nor U10338 (N_10338,N_9865,N_9897);
xnor U10339 (N_10339,N_9941,N_9592);
nor U10340 (N_10340,N_9675,N_9945);
or U10341 (N_10341,N_9942,N_9911);
nor U10342 (N_10342,N_9637,N_9746);
xor U10343 (N_10343,N_9520,N_9612);
nor U10344 (N_10344,N_9558,N_9822);
or U10345 (N_10345,N_9784,N_9595);
or U10346 (N_10346,N_9555,N_9793);
nand U10347 (N_10347,N_9982,N_9903);
nor U10348 (N_10348,N_9799,N_9788);
nand U10349 (N_10349,N_9892,N_9745);
or U10350 (N_10350,N_9899,N_9593);
and U10351 (N_10351,N_9622,N_9984);
nor U10352 (N_10352,N_9948,N_9794);
or U10353 (N_10353,N_9816,N_9905);
nor U10354 (N_10354,N_9991,N_9910);
or U10355 (N_10355,N_9620,N_9720);
and U10356 (N_10356,N_9984,N_9500);
xor U10357 (N_10357,N_9952,N_9613);
nor U10358 (N_10358,N_9913,N_9918);
nand U10359 (N_10359,N_9837,N_9770);
and U10360 (N_10360,N_9794,N_9911);
nand U10361 (N_10361,N_9629,N_9875);
and U10362 (N_10362,N_9521,N_9691);
nand U10363 (N_10363,N_9853,N_9777);
or U10364 (N_10364,N_9982,N_9529);
and U10365 (N_10365,N_9948,N_9649);
xor U10366 (N_10366,N_9882,N_9877);
and U10367 (N_10367,N_9622,N_9790);
and U10368 (N_10368,N_9869,N_9754);
xnor U10369 (N_10369,N_9866,N_9511);
and U10370 (N_10370,N_9824,N_9960);
nand U10371 (N_10371,N_9689,N_9645);
and U10372 (N_10372,N_9512,N_9547);
or U10373 (N_10373,N_9909,N_9742);
and U10374 (N_10374,N_9805,N_9986);
or U10375 (N_10375,N_9574,N_9545);
nor U10376 (N_10376,N_9893,N_9762);
and U10377 (N_10377,N_9729,N_9752);
nand U10378 (N_10378,N_9988,N_9554);
and U10379 (N_10379,N_9895,N_9545);
or U10380 (N_10380,N_9876,N_9765);
xnor U10381 (N_10381,N_9743,N_9998);
and U10382 (N_10382,N_9634,N_9668);
and U10383 (N_10383,N_9743,N_9504);
or U10384 (N_10384,N_9585,N_9514);
nor U10385 (N_10385,N_9747,N_9827);
and U10386 (N_10386,N_9938,N_9608);
or U10387 (N_10387,N_9566,N_9706);
or U10388 (N_10388,N_9900,N_9672);
and U10389 (N_10389,N_9646,N_9904);
nand U10390 (N_10390,N_9762,N_9750);
and U10391 (N_10391,N_9594,N_9754);
or U10392 (N_10392,N_9673,N_9723);
xnor U10393 (N_10393,N_9614,N_9920);
nor U10394 (N_10394,N_9592,N_9985);
nor U10395 (N_10395,N_9870,N_9618);
nand U10396 (N_10396,N_9899,N_9847);
and U10397 (N_10397,N_9824,N_9856);
nor U10398 (N_10398,N_9805,N_9977);
or U10399 (N_10399,N_9884,N_9656);
nand U10400 (N_10400,N_9942,N_9639);
nand U10401 (N_10401,N_9946,N_9937);
xnor U10402 (N_10402,N_9893,N_9985);
nand U10403 (N_10403,N_9674,N_9735);
or U10404 (N_10404,N_9698,N_9943);
nand U10405 (N_10405,N_9753,N_9513);
and U10406 (N_10406,N_9813,N_9515);
xnor U10407 (N_10407,N_9552,N_9844);
xnor U10408 (N_10408,N_9554,N_9593);
nand U10409 (N_10409,N_9850,N_9718);
nand U10410 (N_10410,N_9635,N_9643);
or U10411 (N_10411,N_9891,N_9672);
xnor U10412 (N_10412,N_9961,N_9663);
or U10413 (N_10413,N_9953,N_9794);
nand U10414 (N_10414,N_9552,N_9598);
xor U10415 (N_10415,N_9913,N_9516);
or U10416 (N_10416,N_9814,N_9979);
nand U10417 (N_10417,N_9962,N_9675);
or U10418 (N_10418,N_9786,N_9673);
and U10419 (N_10419,N_9500,N_9862);
or U10420 (N_10420,N_9995,N_9864);
or U10421 (N_10421,N_9919,N_9579);
nand U10422 (N_10422,N_9724,N_9971);
or U10423 (N_10423,N_9636,N_9635);
nand U10424 (N_10424,N_9922,N_9793);
nor U10425 (N_10425,N_9954,N_9577);
nor U10426 (N_10426,N_9742,N_9736);
and U10427 (N_10427,N_9733,N_9527);
nand U10428 (N_10428,N_9846,N_9963);
nor U10429 (N_10429,N_9637,N_9979);
nand U10430 (N_10430,N_9533,N_9621);
or U10431 (N_10431,N_9698,N_9759);
or U10432 (N_10432,N_9504,N_9517);
nor U10433 (N_10433,N_9857,N_9903);
or U10434 (N_10434,N_9673,N_9950);
xor U10435 (N_10435,N_9740,N_9916);
nor U10436 (N_10436,N_9676,N_9531);
nand U10437 (N_10437,N_9535,N_9888);
xnor U10438 (N_10438,N_9650,N_9635);
xnor U10439 (N_10439,N_9532,N_9817);
nor U10440 (N_10440,N_9860,N_9629);
and U10441 (N_10441,N_9723,N_9582);
nand U10442 (N_10442,N_9945,N_9851);
or U10443 (N_10443,N_9756,N_9929);
or U10444 (N_10444,N_9978,N_9996);
and U10445 (N_10445,N_9547,N_9571);
nor U10446 (N_10446,N_9798,N_9874);
nor U10447 (N_10447,N_9618,N_9555);
or U10448 (N_10448,N_9882,N_9981);
or U10449 (N_10449,N_9984,N_9802);
nor U10450 (N_10450,N_9775,N_9891);
and U10451 (N_10451,N_9987,N_9835);
nand U10452 (N_10452,N_9704,N_9833);
nand U10453 (N_10453,N_9591,N_9600);
nor U10454 (N_10454,N_9829,N_9803);
xnor U10455 (N_10455,N_9895,N_9905);
nor U10456 (N_10456,N_9602,N_9726);
nor U10457 (N_10457,N_9573,N_9606);
nand U10458 (N_10458,N_9811,N_9678);
nor U10459 (N_10459,N_9848,N_9534);
nand U10460 (N_10460,N_9921,N_9500);
or U10461 (N_10461,N_9764,N_9619);
nand U10462 (N_10462,N_9548,N_9529);
nand U10463 (N_10463,N_9811,N_9963);
or U10464 (N_10464,N_9661,N_9758);
nor U10465 (N_10465,N_9951,N_9992);
nor U10466 (N_10466,N_9928,N_9790);
nand U10467 (N_10467,N_9793,N_9860);
or U10468 (N_10468,N_9928,N_9911);
and U10469 (N_10469,N_9571,N_9567);
nor U10470 (N_10470,N_9869,N_9717);
or U10471 (N_10471,N_9629,N_9798);
or U10472 (N_10472,N_9932,N_9648);
xor U10473 (N_10473,N_9761,N_9968);
nand U10474 (N_10474,N_9705,N_9535);
nand U10475 (N_10475,N_9634,N_9517);
or U10476 (N_10476,N_9751,N_9500);
or U10477 (N_10477,N_9658,N_9760);
and U10478 (N_10478,N_9876,N_9529);
xor U10479 (N_10479,N_9840,N_9970);
or U10480 (N_10480,N_9512,N_9673);
xor U10481 (N_10481,N_9637,N_9733);
nor U10482 (N_10482,N_9750,N_9817);
xor U10483 (N_10483,N_9537,N_9507);
nor U10484 (N_10484,N_9582,N_9860);
and U10485 (N_10485,N_9605,N_9671);
nor U10486 (N_10486,N_9666,N_9553);
xnor U10487 (N_10487,N_9788,N_9748);
nand U10488 (N_10488,N_9677,N_9636);
nand U10489 (N_10489,N_9806,N_9517);
nor U10490 (N_10490,N_9644,N_9978);
nor U10491 (N_10491,N_9993,N_9748);
and U10492 (N_10492,N_9712,N_9928);
xor U10493 (N_10493,N_9526,N_9787);
or U10494 (N_10494,N_9853,N_9837);
or U10495 (N_10495,N_9514,N_9796);
nor U10496 (N_10496,N_9689,N_9802);
nand U10497 (N_10497,N_9540,N_9903);
nand U10498 (N_10498,N_9839,N_9626);
nand U10499 (N_10499,N_9722,N_9511);
nand U10500 (N_10500,N_10242,N_10410);
and U10501 (N_10501,N_10011,N_10296);
nand U10502 (N_10502,N_10494,N_10070);
xor U10503 (N_10503,N_10367,N_10479);
or U10504 (N_10504,N_10475,N_10269);
or U10505 (N_10505,N_10031,N_10235);
nand U10506 (N_10506,N_10129,N_10039);
nor U10507 (N_10507,N_10270,N_10036);
nand U10508 (N_10508,N_10184,N_10227);
xnor U10509 (N_10509,N_10434,N_10286);
xnor U10510 (N_10510,N_10450,N_10195);
and U10511 (N_10511,N_10003,N_10153);
and U10512 (N_10512,N_10010,N_10412);
nor U10513 (N_10513,N_10355,N_10054);
xnor U10514 (N_10514,N_10482,N_10418);
xnor U10515 (N_10515,N_10188,N_10116);
nor U10516 (N_10516,N_10459,N_10488);
xnor U10517 (N_10517,N_10474,N_10277);
nor U10518 (N_10518,N_10272,N_10178);
xnor U10519 (N_10519,N_10215,N_10134);
xor U10520 (N_10520,N_10218,N_10170);
xor U10521 (N_10521,N_10231,N_10064);
xnor U10522 (N_10522,N_10008,N_10130);
or U10523 (N_10523,N_10062,N_10136);
and U10524 (N_10524,N_10457,N_10425);
nor U10525 (N_10525,N_10106,N_10347);
xor U10526 (N_10526,N_10169,N_10480);
and U10527 (N_10527,N_10144,N_10289);
and U10528 (N_10528,N_10373,N_10161);
and U10529 (N_10529,N_10377,N_10332);
nor U10530 (N_10530,N_10365,N_10466);
and U10531 (N_10531,N_10175,N_10496);
or U10532 (N_10532,N_10113,N_10283);
xnor U10533 (N_10533,N_10135,N_10461);
xor U10534 (N_10534,N_10453,N_10306);
or U10535 (N_10535,N_10383,N_10194);
nand U10536 (N_10536,N_10337,N_10088);
and U10537 (N_10537,N_10366,N_10239);
nor U10538 (N_10538,N_10469,N_10257);
xnor U10539 (N_10539,N_10291,N_10407);
nor U10540 (N_10540,N_10403,N_10063);
nand U10541 (N_10541,N_10455,N_10092);
nor U10542 (N_10542,N_10391,N_10172);
nor U10543 (N_10543,N_10154,N_10320);
or U10544 (N_10544,N_10348,N_10288);
nand U10545 (N_10545,N_10305,N_10318);
or U10546 (N_10546,N_10107,N_10380);
or U10547 (N_10547,N_10173,N_10430);
or U10548 (N_10548,N_10038,N_10137);
or U10549 (N_10549,N_10411,N_10302);
nor U10550 (N_10550,N_10171,N_10234);
nand U10551 (N_10551,N_10444,N_10275);
xor U10552 (N_10552,N_10284,N_10007);
nor U10553 (N_10553,N_10343,N_10065);
or U10554 (N_10554,N_10435,N_10233);
nand U10555 (N_10555,N_10265,N_10117);
and U10556 (N_10556,N_10341,N_10311);
nand U10557 (N_10557,N_10104,N_10087);
and U10558 (N_10558,N_10006,N_10022);
nor U10559 (N_10559,N_10440,N_10149);
xor U10560 (N_10560,N_10133,N_10359);
xnor U10561 (N_10561,N_10371,N_10191);
nor U10562 (N_10562,N_10078,N_10349);
nand U10563 (N_10563,N_10243,N_10351);
nor U10564 (N_10564,N_10478,N_10012);
nand U10565 (N_10565,N_10099,N_10246);
or U10566 (N_10566,N_10045,N_10122);
xor U10567 (N_10567,N_10294,N_10384);
nand U10568 (N_10568,N_10086,N_10448);
or U10569 (N_10569,N_10177,N_10433);
xnor U10570 (N_10570,N_10005,N_10477);
nand U10571 (N_10571,N_10163,N_10376);
and U10572 (N_10572,N_10364,N_10358);
nor U10573 (N_10573,N_10327,N_10160);
nor U10574 (N_10574,N_10100,N_10151);
and U10575 (N_10575,N_10271,N_10309);
and U10576 (N_10576,N_10350,N_10431);
or U10577 (N_10577,N_10324,N_10080);
and U10578 (N_10578,N_10285,N_10115);
nor U10579 (N_10579,N_10203,N_10382);
nor U10580 (N_10580,N_10489,N_10229);
nor U10581 (N_10581,N_10097,N_10110);
nand U10582 (N_10582,N_10046,N_10043);
nand U10583 (N_10583,N_10019,N_10325);
or U10584 (N_10584,N_10458,N_10491);
and U10585 (N_10585,N_10471,N_10408);
nand U10586 (N_10586,N_10159,N_10498);
and U10587 (N_10587,N_10150,N_10344);
or U10588 (N_10588,N_10297,N_10308);
and U10589 (N_10589,N_10386,N_10183);
nor U10590 (N_10590,N_10158,N_10143);
or U10591 (N_10591,N_10472,N_10476);
nand U10592 (N_10592,N_10274,N_10219);
nor U10593 (N_10593,N_10132,N_10220);
nand U10594 (N_10594,N_10211,N_10250);
nand U10595 (N_10595,N_10378,N_10241);
xnor U10596 (N_10596,N_10419,N_10361);
or U10597 (N_10597,N_10016,N_10244);
and U10598 (N_10598,N_10037,N_10413);
or U10599 (N_10599,N_10447,N_10147);
nor U10600 (N_10600,N_10093,N_10090);
xnor U10601 (N_10601,N_10009,N_10214);
and U10602 (N_10602,N_10180,N_10310);
or U10603 (N_10603,N_10298,N_10276);
or U10604 (N_10604,N_10199,N_10254);
nor U10605 (N_10605,N_10095,N_10481);
nor U10606 (N_10606,N_10404,N_10077);
nor U10607 (N_10607,N_10319,N_10048);
nor U10608 (N_10608,N_10345,N_10314);
nor U10609 (N_10609,N_10089,N_10105);
or U10610 (N_10610,N_10436,N_10432);
xor U10611 (N_10611,N_10317,N_10280);
and U10612 (N_10612,N_10399,N_10331);
xnor U10613 (N_10613,N_10210,N_10401);
xor U10614 (N_10614,N_10240,N_10426);
nor U10615 (N_10615,N_10190,N_10109);
xor U10616 (N_10616,N_10312,N_10394);
nand U10617 (N_10617,N_10279,N_10267);
or U10618 (N_10618,N_10222,N_10208);
nor U10619 (N_10619,N_10202,N_10050);
xor U10620 (N_10620,N_10439,N_10185);
or U10621 (N_10621,N_10492,N_10259);
nor U10622 (N_10622,N_10212,N_10186);
and U10623 (N_10623,N_10374,N_10262);
nand U10624 (N_10624,N_10084,N_10493);
and U10625 (N_10625,N_10200,N_10232);
xnor U10626 (N_10626,N_10142,N_10346);
xnor U10627 (N_10627,N_10363,N_10123);
nand U10628 (N_10628,N_10168,N_10072);
nand U10629 (N_10629,N_10193,N_10067);
nor U10630 (N_10630,N_10076,N_10181);
nand U10631 (N_10631,N_10096,N_10381);
nor U10632 (N_10632,N_10004,N_10253);
nor U10633 (N_10633,N_10301,N_10026);
or U10634 (N_10634,N_10372,N_10068);
xnor U10635 (N_10635,N_10463,N_10017);
xnor U10636 (N_10636,N_10035,N_10085);
and U10637 (N_10637,N_10354,N_10299);
xnor U10638 (N_10638,N_10238,N_10249);
xnor U10639 (N_10639,N_10353,N_10395);
xor U10640 (N_10640,N_10443,N_10146);
or U10641 (N_10641,N_10125,N_10082);
or U10642 (N_10642,N_10338,N_10230);
xor U10643 (N_10643,N_10176,N_10454);
nor U10644 (N_10644,N_10390,N_10449);
nand U10645 (N_10645,N_10464,N_10486);
or U10646 (N_10646,N_10487,N_10460);
nand U10647 (N_10647,N_10397,N_10424);
nor U10648 (N_10648,N_10307,N_10266);
or U10649 (N_10649,N_10405,N_10252);
or U10650 (N_10650,N_10442,N_10167);
and U10651 (N_10651,N_10393,N_10369);
or U10652 (N_10652,N_10189,N_10213);
or U10653 (N_10653,N_10079,N_10330);
or U10654 (N_10654,N_10042,N_10237);
nand U10655 (N_10655,N_10245,N_10485);
or U10656 (N_10656,N_10497,N_10462);
or U10657 (N_10657,N_10357,N_10192);
nor U10658 (N_10658,N_10256,N_10326);
xor U10659 (N_10659,N_10282,N_10295);
or U10660 (N_10660,N_10223,N_10131);
nand U10661 (N_10661,N_10198,N_10111);
xnor U10662 (N_10662,N_10217,N_10420);
nand U10663 (N_10663,N_10040,N_10293);
xor U10664 (N_10664,N_10114,N_10402);
or U10665 (N_10665,N_10015,N_10303);
nand U10666 (N_10666,N_10140,N_10335);
nand U10667 (N_10667,N_10069,N_10336);
xnor U10668 (N_10668,N_10162,N_10052);
or U10669 (N_10669,N_10207,N_10081);
or U10670 (N_10670,N_10422,N_10002);
nor U10671 (N_10671,N_10292,N_10101);
nand U10672 (N_10672,N_10251,N_10027);
xor U10673 (N_10673,N_10468,N_10416);
or U10674 (N_10674,N_10248,N_10138);
and U10675 (N_10675,N_10429,N_10427);
nand U10676 (N_10676,N_10152,N_10179);
nor U10677 (N_10677,N_10056,N_10128);
xnor U10678 (N_10678,N_10060,N_10127);
nor U10679 (N_10679,N_10197,N_10164);
nor U10680 (N_10680,N_10165,N_10273);
nor U10681 (N_10681,N_10118,N_10226);
nand U10682 (N_10682,N_10387,N_10228);
or U10683 (N_10683,N_10398,N_10261);
nand U10684 (N_10684,N_10333,N_10417);
xor U10685 (N_10685,N_10124,N_10339);
and U10686 (N_10686,N_10000,N_10368);
or U10687 (N_10687,N_10258,N_10061);
nor U10688 (N_10688,N_10421,N_10409);
nor U10689 (N_10689,N_10014,N_10495);
xnor U10690 (N_10690,N_10033,N_10316);
and U10691 (N_10691,N_10446,N_10224);
or U10692 (N_10692,N_10260,N_10247);
xor U10693 (N_10693,N_10322,N_10334);
or U10694 (N_10694,N_10470,N_10058);
xor U10695 (N_10695,N_10044,N_10406);
nand U10696 (N_10696,N_10073,N_10112);
nand U10697 (N_10697,N_10264,N_10313);
xor U10698 (N_10698,N_10018,N_10385);
nand U10699 (N_10699,N_10362,N_10290);
nor U10700 (N_10700,N_10216,N_10415);
nand U10701 (N_10701,N_10499,N_10196);
nor U10702 (N_10702,N_10389,N_10059);
xnor U10703 (N_10703,N_10323,N_10206);
and U10704 (N_10704,N_10483,N_10108);
nor U10705 (N_10705,N_10051,N_10021);
nand U10706 (N_10706,N_10187,N_10204);
nor U10707 (N_10707,N_10304,N_10379);
nor U10708 (N_10708,N_10263,N_10437);
or U10709 (N_10709,N_10157,N_10083);
and U10710 (N_10710,N_10278,N_10075);
nand U10711 (N_10711,N_10028,N_10091);
nand U10712 (N_10712,N_10360,N_10205);
nor U10713 (N_10713,N_10030,N_10428);
xnor U10714 (N_10714,N_10352,N_10209);
or U10715 (N_10715,N_10120,N_10055);
nor U10716 (N_10716,N_10414,N_10465);
or U10717 (N_10717,N_10236,N_10452);
or U10718 (N_10718,N_10047,N_10121);
nor U10719 (N_10719,N_10156,N_10456);
or U10720 (N_10720,N_10484,N_10102);
and U10721 (N_10721,N_10029,N_10451);
or U10722 (N_10722,N_10053,N_10438);
and U10723 (N_10723,N_10225,N_10141);
and U10724 (N_10724,N_10148,N_10315);
xor U10725 (N_10725,N_10342,N_10103);
xor U10726 (N_10726,N_10074,N_10356);
nand U10727 (N_10727,N_10281,N_10182);
or U10728 (N_10728,N_10032,N_10024);
and U10729 (N_10729,N_10119,N_10145);
nor U10730 (N_10730,N_10268,N_10155);
and U10731 (N_10731,N_10396,N_10066);
nor U10732 (N_10732,N_10287,N_10375);
nand U10733 (N_10733,N_10001,N_10392);
xor U10734 (N_10734,N_10139,N_10020);
xnor U10735 (N_10735,N_10423,N_10445);
nor U10736 (N_10736,N_10370,N_10400);
nor U10737 (N_10737,N_10388,N_10467);
xnor U10738 (N_10738,N_10328,N_10098);
or U10739 (N_10739,N_10490,N_10473);
xnor U10740 (N_10740,N_10057,N_10126);
xnor U10741 (N_10741,N_10201,N_10023);
nand U10742 (N_10742,N_10049,N_10174);
nor U10743 (N_10743,N_10329,N_10221);
or U10744 (N_10744,N_10300,N_10321);
and U10745 (N_10745,N_10034,N_10094);
nor U10746 (N_10746,N_10166,N_10340);
xor U10747 (N_10747,N_10441,N_10041);
nor U10748 (N_10748,N_10013,N_10255);
and U10749 (N_10749,N_10071,N_10025);
nor U10750 (N_10750,N_10359,N_10274);
nand U10751 (N_10751,N_10175,N_10350);
nor U10752 (N_10752,N_10356,N_10221);
xnor U10753 (N_10753,N_10227,N_10194);
and U10754 (N_10754,N_10350,N_10039);
or U10755 (N_10755,N_10365,N_10372);
xnor U10756 (N_10756,N_10084,N_10136);
nand U10757 (N_10757,N_10158,N_10027);
nand U10758 (N_10758,N_10168,N_10456);
xnor U10759 (N_10759,N_10320,N_10463);
nand U10760 (N_10760,N_10125,N_10269);
nor U10761 (N_10761,N_10267,N_10240);
or U10762 (N_10762,N_10358,N_10076);
or U10763 (N_10763,N_10449,N_10436);
nor U10764 (N_10764,N_10313,N_10345);
xor U10765 (N_10765,N_10261,N_10119);
or U10766 (N_10766,N_10153,N_10110);
nor U10767 (N_10767,N_10187,N_10104);
nand U10768 (N_10768,N_10464,N_10469);
nor U10769 (N_10769,N_10215,N_10271);
xor U10770 (N_10770,N_10088,N_10115);
nand U10771 (N_10771,N_10435,N_10090);
and U10772 (N_10772,N_10446,N_10057);
or U10773 (N_10773,N_10393,N_10454);
and U10774 (N_10774,N_10439,N_10155);
and U10775 (N_10775,N_10316,N_10172);
nand U10776 (N_10776,N_10270,N_10241);
nor U10777 (N_10777,N_10051,N_10273);
or U10778 (N_10778,N_10114,N_10417);
nor U10779 (N_10779,N_10121,N_10156);
nand U10780 (N_10780,N_10363,N_10120);
and U10781 (N_10781,N_10145,N_10202);
nor U10782 (N_10782,N_10111,N_10172);
xor U10783 (N_10783,N_10055,N_10292);
or U10784 (N_10784,N_10148,N_10209);
and U10785 (N_10785,N_10047,N_10309);
xor U10786 (N_10786,N_10328,N_10327);
xnor U10787 (N_10787,N_10254,N_10486);
xnor U10788 (N_10788,N_10018,N_10333);
or U10789 (N_10789,N_10433,N_10241);
xnor U10790 (N_10790,N_10204,N_10370);
xnor U10791 (N_10791,N_10306,N_10198);
and U10792 (N_10792,N_10463,N_10418);
xnor U10793 (N_10793,N_10257,N_10315);
and U10794 (N_10794,N_10093,N_10432);
nor U10795 (N_10795,N_10095,N_10213);
or U10796 (N_10796,N_10366,N_10181);
or U10797 (N_10797,N_10044,N_10288);
xor U10798 (N_10798,N_10480,N_10103);
nor U10799 (N_10799,N_10277,N_10468);
or U10800 (N_10800,N_10392,N_10059);
nor U10801 (N_10801,N_10109,N_10254);
xor U10802 (N_10802,N_10325,N_10335);
nor U10803 (N_10803,N_10219,N_10448);
or U10804 (N_10804,N_10217,N_10218);
nand U10805 (N_10805,N_10119,N_10368);
and U10806 (N_10806,N_10146,N_10401);
nor U10807 (N_10807,N_10485,N_10430);
and U10808 (N_10808,N_10061,N_10420);
and U10809 (N_10809,N_10109,N_10173);
xor U10810 (N_10810,N_10207,N_10479);
nand U10811 (N_10811,N_10409,N_10464);
nand U10812 (N_10812,N_10025,N_10045);
nor U10813 (N_10813,N_10461,N_10027);
nand U10814 (N_10814,N_10051,N_10430);
or U10815 (N_10815,N_10412,N_10192);
nand U10816 (N_10816,N_10034,N_10097);
and U10817 (N_10817,N_10001,N_10161);
nor U10818 (N_10818,N_10142,N_10151);
xor U10819 (N_10819,N_10392,N_10332);
nor U10820 (N_10820,N_10354,N_10028);
nor U10821 (N_10821,N_10397,N_10308);
or U10822 (N_10822,N_10471,N_10258);
nand U10823 (N_10823,N_10070,N_10225);
xor U10824 (N_10824,N_10278,N_10473);
xor U10825 (N_10825,N_10097,N_10430);
nor U10826 (N_10826,N_10173,N_10009);
nand U10827 (N_10827,N_10352,N_10309);
and U10828 (N_10828,N_10341,N_10190);
or U10829 (N_10829,N_10102,N_10354);
nand U10830 (N_10830,N_10227,N_10096);
xor U10831 (N_10831,N_10224,N_10075);
or U10832 (N_10832,N_10306,N_10401);
xor U10833 (N_10833,N_10422,N_10362);
nor U10834 (N_10834,N_10098,N_10059);
nor U10835 (N_10835,N_10080,N_10130);
nor U10836 (N_10836,N_10150,N_10351);
or U10837 (N_10837,N_10180,N_10144);
and U10838 (N_10838,N_10195,N_10405);
xnor U10839 (N_10839,N_10287,N_10249);
nor U10840 (N_10840,N_10106,N_10133);
xnor U10841 (N_10841,N_10023,N_10307);
and U10842 (N_10842,N_10223,N_10130);
and U10843 (N_10843,N_10346,N_10305);
xor U10844 (N_10844,N_10036,N_10275);
or U10845 (N_10845,N_10098,N_10442);
nor U10846 (N_10846,N_10067,N_10332);
and U10847 (N_10847,N_10337,N_10487);
and U10848 (N_10848,N_10434,N_10224);
xnor U10849 (N_10849,N_10305,N_10050);
and U10850 (N_10850,N_10302,N_10203);
nand U10851 (N_10851,N_10287,N_10153);
or U10852 (N_10852,N_10115,N_10260);
xor U10853 (N_10853,N_10073,N_10037);
or U10854 (N_10854,N_10125,N_10099);
and U10855 (N_10855,N_10306,N_10336);
xnor U10856 (N_10856,N_10303,N_10222);
or U10857 (N_10857,N_10116,N_10034);
xor U10858 (N_10858,N_10494,N_10295);
or U10859 (N_10859,N_10042,N_10472);
nor U10860 (N_10860,N_10197,N_10496);
and U10861 (N_10861,N_10140,N_10097);
xor U10862 (N_10862,N_10200,N_10060);
or U10863 (N_10863,N_10168,N_10410);
nor U10864 (N_10864,N_10455,N_10142);
nor U10865 (N_10865,N_10160,N_10203);
or U10866 (N_10866,N_10185,N_10492);
xnor U10867 (N_10867,N_10037,N_10494);
and U10868 (N_10868,N_10250,N_10478);
or U10869 (N_10869,N_10179,N_10286);
xnor U10870 (N_10870,N_10045,N_10158);
nor U10871 (N_10871,N_10369,N_10055);
or U10872 (N_10872,N_10076,N_10068);
xnor U10873 (N_10873,N_10312,N_10434);
xor U10874 (N_10874,N_10224,N_10049);
nor U10875 (N_10875,N_10469,N_10485);
nor U10876 (N_10876,N_10348,N_10226);
xnor U10877 (N_10877,N_10373,N_10163);
and U10878 (N_10878,N_10421,N_10111);
nand U10879 (N_10879,N_10232,N_10062);
and U10880 (N_10880,N_10140,N_10468);
nand U10881 (N_10881,N_10332,N_10312);
nand U10882 (N_10882,N_10171,N_10205);
xor U10883 (N_10883,N_10494,N_10169);
nand U10884 (N_10884,N_10207,N_10213);
and U10885 (N_10885,N_10478,N_10207);
nand U10886 (N_10886,N_10215,N_10476);
or U10887 (N_10887,N_10058,N_10292);
nand U10888 (N_10888,N_10171,N_10465);
and U10889 (N_10889,N_10177,N_10019);
nand U10890 (N_10890,N_10487,N_10491);
nand U10891 (N_10891,N_10424,N_10299);
nand U10892 (N_10892,N_10402,N_10196);
xor U10893 (N_10893,N_10050,N_10260);
and U10894 (N_10894,N_10488,N_10078);
nor U10895 (N_10895,N_10050,N_10437);
or U10896 (N_10896,N_10152,N_10203);
nand U10897 (N_10897,N_10356,N_10029);
nand U10898 (N_10898,N_10153,N_10034);
or U10899 (N_10899,N_10496,N_10491);
and U10900 (N_10900,N_10063,N_10433);
xnor U10901 (N_10901,N_10418,N_10284);
nand U10902 (N_10902,N_10075,N_10247);
nor U10903 (N_10903,N_10453,N_10007);
and U10904 (N_10904,N_10109,N_10365);
and U10905 (N_10905,N_10385,N_10491);
and U10906 (N_10906,N_10484,N_10418);
or U10907 (N_10907,N_10252,N_10422);
or U10908 (N_10908,N_10473,N_10290);
nand U10909 (N_10909,N_10330,N_10368);
nor U10910 (N_10910,N_10042,N_10107);
and U10911 (N_10911,N_10178,N_10075);
or U10912 (N_10912,N_10171,N_10252);
and U10913 (N_10913,N_10014,N_10099);
or U10914 (N_10914,N_10349,N_10471);
or U10915 (N_10915,N_10391,N_10388);
nor U10916 (N_10916,N_10099,N_10471);
or U10917 (N_10917,N_10178,N_10051);
xor U10918 (N_10918,N_10224,N_10368);
xor U10919 (N_10919,N_10408,N_10313);
xnor U10920 (N_10920,N_10179,N_10406);
xnor U10921 (N_10921,N_10006,N_10292);
or U10922 (N_10922,N_10095,N_10024);
or U10923 (N_10923,N_10331,N_10424);
nand U10924 (N_10924,N_10104,N_10335);
or U10925 (N_10925,N_10461,N_10118);
nor U10926 (N_10926,N_10215,N_10270);
or U10927 (N_10927,N_10202,N_10192);
xnor U10928 (N_10928,N_10307,N_10219);
and U10929 (N_10929,N_10240,N_10221);
and U10930 (N_10930,N_10112,N_10381);
nor U10931 (N_10931,N_10296,N_10446);
and U10932 (N_10932,N_10392,N_10298);
nor U10933 (N_10933,N_10274,N_10394);
nand U10934 (N_10934,N_10164,N_10256);
nand U10935 (N_10935,N_10119,N_10230);
nor U10936 (N_10936,N_10484,N_10450);
and U10937 (N_10937,N_10287,N_10130);
or U10938 (N_10938,N_10483,N_10303);
or U10939 (N_10939,N_10213,N_10306);
nor U10940 (N_10940,N_10374,N_10380);
or U10941 (N_10941,N_10111,N_10125);
or U10942 (N_10942,N_10149,N_10186);
or U10943 (N_10943,N_10481,N_10245);
nor U10944 (N_10944,N_10118,N_10267);
and U10945 (N_10945,N_10332,N_10379);
or U10946 (N_10946,N_10254,N_10197);
nor U10947 (N_10947,N_10431,N_10494);
or U10948 (N_10948,N_10474,N_10462);
xor U10949 (N_10949,N_10116,N_10272);
xor U10950 (N_10950,N_10422,N_10053);
or U10951 (N_10951,N_10339,N_10490);
nand U10952 (N_10952,N_10145,N_10208);
or U10953 (N_10953,N_10153,N_10215);
xor U10954 (N_10954,N_10025,N_10177);
nor U10955 (N_10955,N_10051,N_10023);
xor U10956 (N_10956,N_10045,N_10305);
nor U10957 (N_10957,N_10067,N_10331);
xnor U10958 (N_10958,N_10002,N_10341);
xnor U10959 (N_10959,N_10219,N_10157);
and U10960 (N_10960,N_10483,N_10007);
and U10961 (N_10961,N_10005,N_10366);
nand U10962 (N_10962,N_10354,N_10037);
nand U10963 (N_10963,N_10278,N_10290);
xor U10964 (N_10964,N_10311,N_10345);
nor U10965 (N_10965,N_10003,N_10093);
xor U10966 (N_10966,N_10161,N_10362);
and U10967 (N_10967,N_10194,N_10093);
nor U10968 (N_10968,N_10184,N_10017);
or U10969 (N_10969,N_10130,N_10254);
xor U10970 (N_10970,N_10234,N_10353);
and U10971 (N_10971,N_10443,N_10454);
or U10972 (N_10972,N_10469,N_10491);
xor U10973 (N_10973,N_10496,N_10183);
xor U10974 (N_10974,N_10045,N_10168);
and U10975 (N_10975,N_10495,N_10066);
xnor U10976 (N_10976,N_10154,N_10244);
and U10977 (N_10977,N_10322,N_10255);
or U10978 (N_10978,N_10230,N_10288);
xor U10979 (N_10979,N_10349,N_10088);
nor U10980 (N_10980,N_10240,N_10200);
nor U10981 (N_10981,N_10247,N_10040);
or U10982 (N_10982,N_10211,N_10002);
or U10983 (N_10983,N_10394,N_10292);
nand U10984 (N_10984,N_10223,N_10497);
nor U10985 (N_10985,N_10420,N_10175);
xnor U10986 (N_10986,N_10458,N_10250);
and U10987 (N_10987,N_10345,N_10202);
and U10988 (N_10988,N_10292,N_10363);
or U10989 (N_10989,N_10415,N_10425);
and U10990 (N_10990,N_10200,N_10447);
and U10991 (N_10991,N_10126,N_10110);
xor U10992 (N_10992,N_10128,N_10465);
nor U10993 (N_10993,N_10447,N_10297);
and U10994 (N_10994,N_10312,N_10110);
and U10995 (N_10995,N_10300,N_10259);
or U10996 (N_10996,N_10245,N_10218);
nor U10997 (N_10997,N_10315,N_10419);
nor U10998 (N_10998,N_10356,N_10237);
xor U10999 (N_10999,N_10059,N_10136);
and U11000 (N_11000,N_10999,N_10733);
nor U11001 (N_11001,N_10825,N_10796);
nor U11002 (N_11002,N_10522,N_10563);
and U11003 (N_11003,N_10828,N_10935);
xnor U11004 (N_11004,N_10583,N_10736);
xnor U11005 (N_11005,N_10647,N_10744);
nand U11006 (N_11006,N_10560,N_10766);
or U11007 (N_11007,N_10725,N_10639);
nand U11008 (N_11008,N_10957,N_10515);
nand U11009 (N_11009,N_10842,N_10875);
and U11010 (N_11010,N_10670,N_10595);
and U11011 (N_11011,N_10547,N_10973);
or U11012 (N_11012,N_10656,N_10518);
nor U11013 (N_11013,N_10528,N_10516);
nor U11014 (N_11014,N_10924,N_10531);
xor U11015 (N_11015,N_10952,N_10755);
nor U11016 (N_11016,N_10967,N_10513);
or U11017 (N_11017,N_10724,N_10554);
nor U11018 (N_11018,N_10698,N_10731);
nor U11019 (N_11019,N_10751,N_10584);
nand U11020 (N_11020,N_10809,N_10507);
nand U11021 (N_11021,N_10642,N_10675);
nor U11022 (N_11022,N_10890,N_10634);
and U11023 (N_11023,N_10839,N_10808);
nor U11024 (N_11024,N_10536,N_10974);
nand U11025 (N_11025,N_10549,N_10601);
or U11026 (N_11026,N_10718,N_10722);
or U11027 (N_11027,N_10691,N_10701);
and U11028 (N_11028,N_10623,N_10501);
nand U11029 (N_11029,N_10986,N_10747);
or U11030 (N_11030,N_10985,N_10785);
or U11031 (N_11031,N_10961,N_10877);
and U11032 (N_11032,N_10590,N_10616);
xnor U11033 (N_11033,N_10962,N_10772);
nand U11034 (N_11034,N_10754,N_10543);
nand U11035 (N_11035,N_10537,N_10844);
nor U11036 (N_11036,N_10867,N_10704);
and U11037 (N_11037,N_10949,N_10685);
nand U11038 (N_11038,N_10683,N_10887);
and U11039 (N_11039,N_10948,N_10661);
nand U11040 (N_11040,N_10566,N_10805);
xor U11041 (N_11041,N_10697,N_10599);
and U11042 (N_11042,N_10569,N_10795);
xor U11043 (N_11043,N_10835,N_10721);
nand U11044 (N_11044,N_10644,N_10810);
and U11045 (N_11045,N_10800,N_10770);
xnor U11046 (N_11046,N_10571,N_10862);
or U11047 (N_11047,N_10752,N_10971);
nor U11048 (N_11048,N_10976,N_10711);
nor U11049 (N_11049,N_10542,N_10960);
nand U11050 (N_11050,N_10928,N_10730);
nand U11051 (N_11051,N_10585,N_10719);
nand U11052 (N_11052,N_10605,N_10776);
or U11053 (N_11053,N_10598,N_10832);
xor U11054 (N_11054,N_10654,N_10758);
nand U11055 (N_11055,N_10622,N_10523);
or U11056 (N_11056,N_10527,N_10597);
nand U11057 (N_11057,N_10706,N_10911);
xor U11058 (N_11058,N_10658,N_10552);
or U11059 (N_11059,N_10743,N_10727);
nor U11060 (N_11060,N_10896,N_10612);
nor U11061 (N_11061,N_10892,N_10781);
or U11062 (N_11062,N_10633,N_10655);
nand U11063 (N_11063,N_10525,N_10607);
nor U11064 (N_11064,N_10717,N_10760);
or U11065 (N_11065,N_10780,N_10942);
nand U11066 (N_11066,N_10640,N_10530);
or U11067 (N_11067,N_10871,N_10915);
and U11068 (N_11068,N_10574,N_10749);
or U11069 (N_11069,N_10801,N_10845);
or U11070 (N_11070,N_10506,N_10895);
xnor U11071 (N_11071,N_10664,N_10782);
nand U11072 (N_11072,N_10550,N_10577);
xnor U11073 (N_11073,N_10994,N_10763);
and U11074 (N_11074,N_10826,N_10831);
xnor U11075 (N_11075,N_10578,N_10816);
nand U11076 (N_11076,N_10936,N_10557);
nand U11077 (N_11077,N_10676,N_10987);
nor U11078 (N_11078,N_10619,N_10672);
nor U11079 (N_11079,N_10740,N_10742);
and U11080 (N_11080,N_10545,N_10868);
and U11081 (N_11081,N_10524,N_10790);
or U11082 (N_11082,N_10723,N_10881);
or U11083 (N_11083,N_10645,N_10972);
nor U11084 (N_11084,N_10709,N_10561);
xnor U11085 (N_11085,N_10668,N_10682);
or U11086 (N_11086,N_10592,N_10850);
or U11087 (N_11087,N_10857,N_10600);
or U11088 (N_11088,N_10694,N_10880);
and U11089 (N_11089,N_10833,N_10716);
nand U11090 (N_11090,N_10617,N_10980);
and U11091 (N_11091,N_10753,N_10848);
nand U11092 (N_11092,N_10927,N_10837);
nand U11093 (N_11093,N_10579,N_10937);
nand U11094 (N_11094,N_10684,N_10686);
and U11095 (N_11095,N_10678,N_10765);
nor U11096 (N_11096,N_10629,N_10852);
nand U11097 (N_11097,N_10631,N_10863);
or U11098 (N_11098,N_10983,N_10945);
or U11099 (N_11099,N_10939,N_10720);
or U11100 (N_11100,N_10604,N_10514);
or U11101 (N_11101,N_10568,N_10856);
or U11102 (N_11102,N_10503,N_10541);
nor U11103 (N_11103,N_10659,N_10797);
or U11104 (N_11104,N_10827,N_10533);
xnor U11105 (N_11105,N_10933,N_10556);
or U11106 (N_11106,N_10705,N_10884);
or U11107 (N_11107,N_10990,N_10934);
and U11108 (N_11108,N_10912,N_10944);
and U11109 (N_11109,N_10943,N_10546);
and U11110 (N_11110,N_10692,N_10918);
or U11111 (N_11111,N_10728,N_10998);
nor U11112 (N_11112,N_10926,N_10914);
or U11113 (N_11113,N_10829,N_10677);
xor U11114 (N_11114,N_10648,N_10846);
xnor U11115 (N_11115,N_10535,N_10930);
nor U11116 (N_11116,N_10562,N_10786);
and U11117 (N_11117,N_10789,N_10570);
nand U11118 (N_11118,N_10575,N_10778);
nor U11119 (N_11119,N_10941,N_10613);
or U11120 (N_11120,N_10762,N_10874);
nand U11121 (N_11121,N_10687,N_10632);
nor U11122 (N_11122,N_10995,N_10872);
nor U11123 (N_11123,N_10788,N_10925);
xnor U11124 (N_11124,N_10910,N_10703);
or U11125 (N_11125,N_10602,N_10611);
nand U11126 (N_11126,N_10618,N_10919);
xor U11127 (N_11127,N_10699,N_10558);
xor U11128 (N_11128,N_10869,N_10965);
xnor U11129 (N_11129,N_10667,N_10768);
nand U11130 (N_11130,N_10851,N_10764);
or U11131 (N_11131,N_10759,N_10540);
nand U11132 (N_11132,N_10997,N_10932);
or U11133 (N_11133,N_10521,N_10643);
or U11134 (N_11134,N_10573,N_10886);
xor U11135 (N_11135,N_10773,N_10870);
and U11136 (N_11136,N_10970,N_10586);
nor U11137 (N_11137,N_10906,N_10984);
xnor U11138 (N_11138,N_10783,N_10534);
xnor U11139 (N_11139,N_10913,N_10861);
nor U11140 (N_11140,N_10843,N_10876);
nor U11141 (N_11141,N_10663,N_10609);
or U11142 (N_11142,N_10700,N_10806);
or U11143 (N_11143,N_10761,N_10958);
nand U11144 (N_11144,N_10505,N_10679);
and U11145 (N_11145,N_10581,N_10904);
xnor U11146 (N_11146,N_10779,N_10963);
nor U11147 (N_11147,N_10738,N_10903);
nor U11148 (N_11148,N_10898,N_10729);
nor U11149 (N_11149,N_10660,N_10813);
or U11150 (N_11150,N_10688,N_10519);
nand U11151 (N_11151,N_10538,N_10750);
and U11152 (N_11152,N_10854,N_10879);
nor U11153 (N_11153,N_10812,N_10500);
and U11154 (N_11154,N_10671,N_10565);
nand U11155 (N_11155,N_10741,N_10866);
or U11156 (N_11156,N_10964,N_10784);
and U11157 (N_11157,N_10849,N_10900);
or U11158 (N_11158,N_10793,N_10950);
xor U11159 (N_11159,N_10883,N_10951);
nor U11160 (N_11160,N_10799,N_10572);
and U11161 (N_11161,N_10509,N_10610);
or U11162 (N_11162,N_10502,N_10710);
nand U11163 (N_11163,N_10511,N_10504);
and U11164 (N_11164,N_10767,N_10836);
nor U11165 (N_11165,N_10931,N_10715);
nand U11166 (N_11166,N_10917,N_10582);
xor U11167 (N_11167,N_10596,N_10627);
nor U11168 (N_11168,N_10587,N_10746);
and U11169 (N_11169,N_10975,N_10737);
xor U11170 (N_11170,N_10508,N_10690);
xor U11171 (N_11171,N_10544,N_10641);
and U11172 (N_11172,N_10588,N_10916);
and U11173 (N_11173,N_10794,N_10966);
or U11174 (N_11174,N_10787,N_10988);
nor U11175 (N_11175,N_10593,N_10745);
and U11176 (N_11176,N_10920,N_10882);
nand U11177 (N_11177,N_10946,N_10662);
xnor U11178 (N_11178,N_10708,N_10955);
nor U11179 (N_11179,N_10996,N_10673);
or U11180 (N_11180,N_10624,N_10646);
and U11181 (N_11181,N_10638,N_10817);
nor U11182 (N_11182,N_10713,N_10732);
xnor U11183 (N_11183,N_10901,N_10769);
and U11184 (N_11184,N_10712,N_10815);
or U11185 (N_11185,N_10860,N_10714);
xnor U11186 (N_11186,N_10969,N_10968);
xnor U11187 (N_11187,N_10921,N_10680);
nor U11188 (N_11188,N_10665,N_10635);
nand U11189 (N_11189,N_10807,N_10991);
and U11190 (N_11190,N_10539,N_10978);
nor U11191 (N_11191,N_10636,N_10702);
or U11192 (N_11192,N_10657,N_10707);
or U11193 (N_11193,N_10567,N_10838);
xnor U11194 (N_11194,N_10865,N_10748);
and U11195 (N_11195,N_10981,N_10902);
and U11196 (N_11196,N_10532,N_10823);
xnor U11197 (N_11197,N_10814,N_10653);
nand U11198 (N_11198,N_10982,N_10989);
xnor U11199 (N_11199,N_10938,N_10628);
xor U11200 (N_11200,N_10953,N_10922);
nor U11201 (N_11201,N_10822,N_10517);
and U11202 (N_11202,N_10615,N_10847);
xnor U11203 (N_11203,N_10804,N_10821);
xor U11204 (N_11204,N_10603,N_10689);
nor U11205 (N_11205,N_10929,N_10757);
nor U11206 (N_11206,N_10548,N_10564);
nand U11207 (N_11207,N_10947,N_10651);
xnor U11208 (N_11208,N_10529,N_10859);
nor U11209 (N_11209,N_10853,N_10681);
nand U11210 (N_11210,N_10885,N_10803);
or U11211 (N_11211,N_10621,N_10551);
nand U11212 (N_11212,N_10591,N_10555);
and U11213 (N_11213,N_10907,N_10830);
nand U11214 (N_11214,N_10589,N_10889);
nor U11215 (N_11215,N_10693,N_10553);
xor U11216 (N_11216,N_10798,N_10802);
nor U11217 (N_11217,N_10649,N_10606);
and U11218 (N_11218,N_10739,N_10894);
nor U11219 (N_11219,N_10580,N_10735);
and U11220 (N_11220,N_10792,N_10510);
or U11221 (N_11221,N_10734,N_10630);
and U11222 (N_11222,N_10771,N_10669);
nor U11223 (N_11223,N_10841,N_10908);
nor U11224 (N_11224,N_10940,N_10992);
nor U11225 (N_11225,N_10559,N_10858);
and U11226 (N_11226,N_10626,N_10864);
nand U11227 (N_11227,N_10820,N_10625);
nand U11228 (N_11228,N_10909,N_10756);
nand U11229 (N_11229,N_10594,N_10614);
and U11230 (N_11230,N_10774,N_10993);
xnor U11231 (N_11231,N_10637,N_10840);
or U11232 (N_11232,N_10855,N_10650);
or U11233 (N_11233,N_10959,N_10791);
xnor U11234 (N_11234,N_10620,N_10512);
or U11235 (N_11235,N_10979,N_10775);
nor U11236 (N_11236,N_10526,N_10893);
nor U11237 (N_11237,N_10897,N_10666);
and U11238 (N_11238,N_10873,N_10777);
and U11239 (N_11239,N_10652,N_10819);
nor U11240 (N_11240,N_10899,N_10891);
nor U11241 (N_11241,N_10608,N_10811);
nor U11242 (N_11242,N_10905,N_10696);
xor U11243 (N_11243,N_10923,N_10956);
nor U11244 (N_11244,N_10576,N_10977);
or U11245 (N_11245,N_10954,N_10695);
and U11246 (N_11246,N_10674,N_10726);
xor U11247 (N_11247,N_10818,N_10878);
xnor U11248 (N_11248,N_10834,N_10520);
or U11249 (N_11249,N_10824,N_10888);
nand U11250 (N_11250,N_10788,N_10853);
nor U11251 (N_11251,N_10602,N_10858);
and U11252 (N_11252,N_10889,N_10811);
nand U11253 (N_11253,N_10961,N_10855);
or U11254 (N_11254,N_10505,N_10829);
nor U11255 (N_11255,N_10705,N_10751);
xnor U11256 (N_11256,N_10815,N_10692);
and U11257 (N_11257,N_10761,N_10821);
or U11258 (N_11258,N_10798,N_10980);
nor U11259 (N_11259,N_10816,N_10890);
nor U11260 (N_11260,N_10648,N_10886);
nor U11261 (N_11261,N_10614,N_10792);
nand U11262 (N_11262,N_10946,N_10560);
and U11263 (N_11263,N_10632,N_10676);
or U11264 (N_11264,N_10841,N_10818);
nand U11265 (N_11265,N_10535,N_10687);
or U11266 (N_11266,N_10761,N_10947);
nor U11267 (N_11267,N_10578,N_10746);
or U11268 (N_11268,N_10971,N_10620);
xor U11269 (N_11269,N_10671,N_10937);
or U11270 (N_11270,N_10795,N_10538);
and U11271 (N_11271,N_10930,N_10602);
and U11272 (N_11272,N_10703,N_10715);
nand U11273 (N_11273,N_10885,N_10893);
nand U11274 (N_11274,N_10798,N_10646);
xnor U11275 (N_11275,N_10543,N_10884);
xor U11276 (N_11276,N_10666,N_10539);
or U11277 (N_11277,N_10507,N_10901);
nor U11278 (N_11278,N_10902,N_10876);
xor U11279 (N_11279,N_10913,N_10698);
nor U11280 (N_11280,N_10846,N_10976);
xor U11281 (N_11281,N_10508,N_10731);
and U11282 (N_11282,N_10909,N_10874);
nand U11283 (N_11283,N_10988,N_10850);
nor U11284 (N_11284,N_10693,N_10640);
and U11285 (N_11285,N_10764,N_10510);
nor U11286 (N_11286,N_10906,N_10816);
or U11287 (N_11287,N_10844,N_10982);
or U11288 (N_11288,N_10830,N_10911);
xor U11289 (N_11289,N_10779,N_10737);
or U11290 (N_11290,N_10694,N_10871);
nand U11291 (N_11291,N_10526,N_10615);
or U11292 (N_11292,N_10521,N_10539);
xor U11293 (N_11293,N_10787,N_10987);
or U11294 (N_11294,N_10809,N_10755);
or U11295 (N_11295,N_10693,N_10634);
nand U11296 (N_11296,N_10662,N_10524);
or U11297 (N_11297,N_10672,N_10991);
nor U11298 (N_11298,N_10792,N_10936);
and U11299 (N_11299,N_10577,N_10943);
nand U11300 (N_11300,N_10630,N_10730);
nor U11301 (N_11301,N_10983,N_10766);
xor U11302 (N_11302,N_10907,N_10910);
or U11303 (N_11303,N_10915,N_10782);
xor U11304 (N_11304,N_10664,N_10515);
xnor U11305 (N_11305,N_10867,N_10894);
nand U11306 (N_11306,N_10673,N_10506);
and U11307 (N_11307,N_10626,N_10907);
nor U11308 (N_11308,N_10593,N_10840);
and U11309 (N_11309,N_10967,N_10609);
nand U11310 (N_11310,N_10580,N_10520);
nand U11311 (N_11311,N_10657,N_10599);
or U11312 (N_11312,N_10873,N_10632);
xor U11313 (N_11313,N_10711,N_10757);
nor U11314 (N_11314,N_10894,N_10614);
and U11315 (N_11315,N_10932,N_10860);
or U11316 (N_11316,N_10511,N_10918);
or U11317 (N_11317,N_10855,N_10608);
nand U11318 (N_11318,N_10563,N_10731);
xnor U11319 (N_11319,N_10541,N_10898);
or U11320 (N_11320,N_10723,N_10699);
nor U11321 (N_11321,N_10925,N_10915);
nor U11322 (N_11322,N_10889,N_10765);
nand U11323 (N_11323,N_10904,N_10845);
xor U11324 (N_11324,N_10856,N_10776);
and U11325 (N_11325,N_10674,N_10573);
or U11326 (N_11326,N_10595,N_10789);
and U11327 (N_11327,N_10719,N_10575);
or U11328 (N_11328,N_10638,N_10845);
or U11329 (N_11329,N_10863,N_10544);
xnor U11330 (N_11330,N_10791,N_10686);
or U11331 (N_11331,N_10626,N_10729);
xor U11332 (N_11332,N_10600,N_10647);
and U11333 (N_11333,N_10714,N_10897);
nor U11334 (N_11334,N_10987,N_10531);
and U11335 (N_11335,N_10509,N_10520);
nand U11336 (N_11336,N_10810,N_10816);
nor U11337 (N_11337,N_10677,N_10787);
or U11338 (N_11338,N_10588,N_10874);
or U11339 (N_11339,N_10803,N_10963);
xor U11340 (N_11340,N_10525,N_10592);
xnor U11341 (N_11341,N_10681,N_10627);
nor U11342 (N_11342,N_10519,N_10671);
nand U11343 (N_11343,N_10626,N_10676);
nor U11344 (N_11344,N_10749,N_10944);
nand U11345 (N_11345,N_10954,N_10514);
nand U11346 (N_11346,N_10967,N_10692);
nor U11347 (N_11347,N_10656,N_10538);
nor U11348 (N_11348,N_10960,N_10577);
nand U11349 (N_11349,N_10505,N_10807);
nand U11350 (N_11350,N_10787,N_10699);
xor U11351 (N_11351,N_10611,N_10516);
nor U11352 (N_11352,N_10881,N_10746);
nor U11353 (N_11353,N_10691,N_10955);
nor U11354 (N_11354,N_10993,N_10989);
xnor U11355 (N_11355,N_10655,N_10589);
or U11356 (N_11356,N_10528,N_10564);
and U11357 (N_11357,N_10901,N_10565);
xor U11358 (N_11358,N_10621,N_10833);
or U11359 (N_11359,N_10506,N_10887);
nor U11360 (N_11360,N_10899,N_10777);
xor U11361 (N_11361,N_10698,N_10931);
nand U11362 (N_11362,N_10981,N_10549);
nor U11363 (N_11363,N_10721,N_10967);
nor U11364 (N_11364,N_10984,N_10861);
nand U11365 (N_11365,N_10917,N_10768);
or U11366 (N_11366,N_10917,N_10993);
xnor U11367 (N_11367,N_10752,N_10755);
or U11368 (N_11368,N_10817,N_10834);
xor U11369 (N_11369,N_10896,N_10937);
nor U11370 (N_11370,N_10791,N_10665);
nand U11371 (N_11371,N_10978,N_10881);
nand U11372 (N_11372,N_10949,N_10925);
or U11373 (N_11373,N_10995,N_10655);
nor U11374 (N_11374,N_10688,N_10975);
nand U11375 (N_11375,N_10994,N_10897);
xor U11376 (N_11376,N_10661,N_10714);
xnor U11377 (N_11377,N_10704,N_10956);
nor U11378 (N_11378,N_10602,N_10950);
nand U11379 (N_11379,N_10983,N_10911);
or U11380 (N_11380,N_10859,N_10900);
or U11381 (N_11381,N_10803,N_10733);
or U11382 (N_11382,N_10687,N_10506);
nand U11383 (N_11383,N_10715,N_10687);
xnor U11384 (N_11384,N_10712,N_10802);
xnor U11385 (N_11385,N_10828,N_10778);
or U11386 (N_11386,N_10837,N_10632);
nor U11387 (N_11387,N_10953,N_10883);
or U11388 (N_11388,N_10964,N_10628);
xnor U11389 (N_11389,N_10748,N_10813);
xor U11390 (N_11390,N_10952,N_10658);
nor U11391 (N_11391,N_10896,N_10628);
nor U11392 (N_11392,N_10807,N_10814);
nand U11393 (N_11393,N_10913,N_10539);
nor U11394 (N_11394,N_10647,N_10751);
nor U11395 (N_11395,N_10827,N_10803);
and U11396 (N_11396,N_10854,N_10795);
nand U11397 (N_11397,N_10600,N_10549);
and U11398 (N_11398,N_10916,N_10532);
xor U11399 (N_11399,N_10884,N_10829);
nand U11400 (N_11400,N_10896,N_10996);
nand U11401 (N_11401,N_10924,N_10915);
xnor U11402 (N_11402,N_10815,N_10819);
or U11403 (N_11403,N_10518,N_10827);
or U11404 (N_11404,N_10672,N_10850);
nand U11405 (N_11405,N_10631,N_10816);
nor U11406 (N_11406,N_10793,N_10847);
nor U11407 (N_11407,N_10600,N_10899);
nor U11408 (N_11408,N_10886,N_10819);
and U11409 (N_11409,N_10998,N_10782);
nand U11410 (N_11410,N_10624,N_10741);
nor U11411 (N_11411,N_10813,N_10600);
and U11412 (N_11412,N_10868,N_10702);
and U11413 (N_11413,N_10987,N_10949);
xnor U11414 (N_11414,N_10637,N_10997);
xor U11415 (N_11415,N_10991,N_10838);
nand U11416 (N_11416,N_10768,N_10946);
nor U11417 (N_11417,N_10623,N_10542);
or U11418 (N_11418,N_10655,N_10616);
nor U11419 (N_11419,N_10910,N_10641);
nand U11420 (N_11420,N_10592,N_10821);
and U11421 (N_11421,N_10937,N_10818);
or U11422 (N_11422,N_10639,N_10592);
and U11423 (N_11423,N_10604,N_10735);
nor U11424 (N_11424,N_10641,N_10545);
nor U11425 (N_11425,N_10571,N_10918);
nand U11426 (N_11426,N_10512,N_10593);
or U11427 (N_11427,N_10967,N_10806);
and U11428 (N_11428,N_10599,N_10896);
nor U11429 (N_11429,N_10545,N_10644);
nor U11430 (N_11430,N_10926,N_10592);
and U11431 (N_11431,N_10995,N_10736);
nand U11432 (N_11432,N_10678,N_10741);
and U11433 (N_11433,N_10913,N_10880);
and U11434 (N_11434,N_10673,N_10601);
xor U11435 (N_11435,N_10510,N_10938);
nand U11436 (N_11436,N_10768,N_10658);
or U11437 (N_11437,N_10814,N_10576);
and U11438 (N_11438,N_10901,N_10509);
or U11439 (N_11439,N_10550,N_10524);
or U11440 (N_11440,N_10906,N_10913);
or U11441 (N_11441,N_10710,N_10818);
nor U11442 (N_11442,N_10600,N_10855);
or U11443 (N_11443,N_10948,N_10756);
or U11444 (N_11444,N_10701,N_10602);
and U11445 (N_11445,N_10704,N_10702);
nor U11446 (N_11446,N_10808,N_10621);
nand U11447 (N_11447,N_10830,N_10800);
and U11448 (N_11448,N_10788,N_10733);
or U11449 (N_11449,N_10906,N_10722);
nand U11450 (N_11450,N_10850,N_10856);
and U11451 (N_11451,N_10849,N_10725);
and U11452 (N_11452,N_10887,N_10576);
or U11453 (N_11453,N_10894,N_10522);
nand U11454 (N_11454,N_10843,N_10852);
or U11455 (N_11455,N_10564,N_10728);
nand U11456 (N_11456,N_10615,N_10661);
xnor U11457 (N_11457,N_10542,N_10582);
nand U11458 (N_11458,N_10819,N_10951);
xnor U11459 (N_11459,N_10841,N_10902);
and U11460 (N_11460,N_10795,N_10614);
or U11461 (N_11461,N_10696,N_10626);
nand U11462 (N_11462,N_10671,N_10817);
or U11463 (N_11463,N_10889,N_10629);
nand U11464 (N_11464,N_10730,N_10692);
and U11465 (N_11465,N_10942,N_10582);
nand U11466 (N_11466,N_10904,N_10771);
xor U11467 (N_11467,N_10888,N_10520);
nor U11468 (N_11468,N_10808,N_10698);
and U11469 (N_11469,N_10693,N_10958);
or U11470 (N_11470,N_10740,N_10652);
nand U11471 (N_11471,N_10542,N_10931);
and U11472 (N_11472,N_10982,N_10615);
nand U11473 (N_11473,N_10924,N_10512);
nand U11474 (N_11474,N_10508,N_10787);
nor U11475 (N_11475,N_10903,N_10823);
xor U11476 (N_11476,N_10884,N_10647);
xor U11477 (N_11477,N_10644,N_10957);
nand U11478 (N_11478,N_10567,N_10776);
nand U11479 (N_11479,N_10565,N_10948);
nor U11480 (N_11480,N_10640,N_10904);
xnor U11481 (N_11481,N_10960,N_10828);
and U11482 (N_11482,N_10898,N_10670);
xor U11483 (N_11483,N_10673,N_10990);
nand U11484 (N_11484,N_10802,N_10873);
nor U11485 (N_11485,N_10854,N_10522);
nor U11486 (N_11486,N_10980,N_10805);
xor U11487 (N_11487,N_10591,N_10685);
nor U11488 (N_11488,N_10607,N_10948);
and U11489 (N_11489,N_10698,N_10528);
nand U11490 (N_11490,N_10793,N_10869);
nand U11491 (N_11491,N_10670,N_10594);
or U11492 (N_11492,N_10615,N_10586);
nand U11493 (N_11493,N_10557,N_10751);
nand U11494 (N_11494,N_10900,N_10511);
or U11495 (N_11495,N_10784,N_10557);
nand U11496 (N_11496,N_10685,N_10916);
nand U11497 (N_11497,N_10553,N_10556);
and U11498 (N_11498,N_10936,N_10779);
nand U11499 (N_11499,N_10589,N_10573);
and U11500 (N_11500,N_11370,N_11111);
and U11501 (N_11501,N_11160,N_11498);
xor U11502 (N_11502,N_11438,N_11223);
nor U11503 (N_11503,N_11190,N_11271);
or U11504 (N_11504,N_11246,N_11466);
nand U11505 (N_11505,N_11492,N_11291);
or U11506 (N_11506,N_11331,N_11046);
and U11507 (N_11507,N_11432,N_11118);
xor U11508 (N_11508,N_11139,N_11040);
nand U11509 (N_11509,N_11250,N_11342);
or U11510 (N_11510,N_11390,N_11281);
and U11511 (N_11511,N_11032,N_11476);
or U11512 (N_11512,N_11109,N_11147);
nor U11513 (N_11513,N_11177,N_11297);
xnor U11514 (N_11514,N_11174,N_11430);
or U11515 (N_11515,N_11255,N_11140);
nand U11516 (N_11516,N_11361,N_11102);
xnor U11517 (N_11517,N_11153,N_11168);
nor U11518 (N_11518,N_11080,N_11386);
xor U11519 (N_11519,N_11487,N_11303);
nor U11520 (N_11520,N_11194,N_11106);
nor U11521 (N_11521,N_11004,N_11061);
xor U11522 (N_11522,N_11065,N_11403);
nor U11523 (N_11523,N_11346,N_11129);
xnor U11524 (N_11524,N_11339,N_11182);
or U11525 (N_11525,N_11460,N_11068);
xnor U11526 (N_11526,N_11031,N_11146);
nand U11527 (N_11527,N_11298,N_11284);
nor U11528 (N_11528,N_11204,N_11343);
or U11529 (N_11529,N_11202,N_11063);
nor U11530 (N_11530,N_11107,N_11021);
and U11531 (N_11531,N_11056,N_11469);
xnor U11532 (N_11532,N_11156,N_11385);
nor U11533 (N_11533,N_11286,N_11364);
or U11534 (N_11534,N_11208,N_11095);
and U11535 (N_11535,N_11071,N_11131);
xnor U11536 (N_11536,N_11406,N_11400);
nor U11537 (N_11537,N_11353,N_11167);
or U11538 (N_11538,N_11148,N_11435);
nor U11539 (N_11539,N_11277,N_11493);
and U11540 (N_11540,N_11285,N_11037);
nand U11541 (N_11541,N_11012,N_11072);
or U11542 (N_11542,N_11312,N_11247);
and U11543 (N_11543,N_11402,N_11424);
nor U11544 (N_11544,N_11011,N_11451);
nor U11545 (N_11545,N_11151,N_11366);
and U11546 (N_11546,N_11470,N_11007);
xor U11547 (N_11547,N_11444,N_11264);
and U11548 (N_11548,N_11067,N_11000);
nand U11549 (N_11549,N_11468,N_11422);
or U11550 (N_11550,N_11069,N_11409);
nand U11551 (N_11551,N_11036,N_11454);
or U11552 (N_11552,N_11041,N_11332);
and U11553 (N_11553,N_11196,N_11395);
and U11554 (N_11554,N_11333,N_11462);
nor U11555 (N_11555,N_11132,N_11251);
xor U11556 (N_11556,N_11209,N_11280);
nand U11557 (N_11557,N_11491,N_11391);
and U11558 (N_11558,N_11389,N_11175);
xor U11559 (N_11559,N_11099,N_11265);
and U11560 (N_11560,N_11016,N_11472);
nor U11561 (N_11561,N_11443,N_11098);
xnor U11562 (N_11562,N_11425,N_11112);
or U11563 (N_11563,N_11115,N_11218);
or U11564 (N_11564,N_11283,N_11412);
nand U11565 (N_11565,N_11038,N_11494);
nor U11566 (N_11566,N_11119,N_11445);
nor U11567 (N_11567,N_11481,N_11214);
xor U11568 (N_11568,N_11014,N_11378);
nor U11569 (N_11569,N_11211,N_11234);
xor U11570 (N_11570,N_11117,N_11348);
nand U11571 (N_11571,N_11164,N_11166);
or U11572 (N_11572,N_11024,N_11315);
and U11573 (N_11573,N_11242,N_11350);
nor U11574 (N_11574,N_11376,N_11496);
and U11575 (N_11575,N_11306,N_11133);
nand U11576 (N_11576,N_11467,N_11437);
or U11577 (N_11577,N_11192,N_11262);
xor U11578 (N_11578,N_11310,N_11354);
or U11579 (N_11579,N_11274,N_11159);
nand U11580 (N_11580,N_11313,N_11407);
xor U11581 (N_11581,N_11222,N_11050);
nor U11582 (N_11582,N_11236,N_11042);
nor U11583 (N_11583,N_11232,N_11455);
or U11584 (N_11584,N_11244,N_11170);
nor U11585 (N_11585,N_11157,N_11113);
nor U11586 (N_11586,N_11290,N_11154);
nor U11587 (N_11587,N_11052,N_11125);
nor U11588 (N_11588,N_11075,N_11230);
nor U11589 (N_11589,N_11296,N_11155);
and U11590 (N_11590,N_11377,N_11365);
xnor U11591 (N_11591,N_11076,N_11097);
nand U11592 (N_11592,N_11374,N_11039);
or U11593 (N_11593,N_11482,N_11198);
nand U11594 (N_11594,N_11427,N_11373);
xnor U11595 (N_11595,N_11461,N_11173);
xnor U11596 (N_11596,N_11272,N_11143);
nor U11597 (N_11597,N_11352,N_11187);
and U11598 (N_11598,N_11267,N_11420);
nor U11599 (N_11599,N_11404,N_11319);
or U11600 (N_11600,N_11320,N_11431);
or U11601 (N_11601,N_11300,N_11380);
or U11602 (N_11602,N_11200,N_11464);
xor U11603 (N_11603,N_11375,N_11077);
and U11604 (N_11604,N_11266,N_11417);
nand U11605 (N_11605,N_11261,N_11362);
or U11606 (N_11606,N_11488,N_11110);
and U11607 (N_11607,N_11446,N_11100);
or U11608 (N_11608,N_11135,N_11413);
and U11609 (N_11609,N_11235,N_11338);
and U11610 (N_11610,N_11340,N_11330);
xnor U11611 (N_11611,N_11189,N_11219);
or U11612 (N_11612,N_11321,N_11318);
nor U11613 (N_11613,N_11176,N_11322);
xor U11614 (N_11614,N_11458,N_11087);
nor U11615 (N_11615,N_11387,N_11185);
or U11616 (N_11616,N_11029,N_11019);
nand U11617 (N_11617,N_11171,N_11163);
and U11618 (N_11618,N_11142,N_11203);
or U11619 (N_11619,N_11263,N_11127);
nand U11620 (N_11620,N_11017,N_11270);
xnor U11621 (N_11621,N_11020,N_11399);
nor U11622 (N_11622,N_11256,N_11121);
xnor U11623 (N_11623,N_11079,N_11186);
and U11624 (N_11624,N_11311,N_11015);
xnor U11625 (N_11625,N_11237,N_11005);
nand U11626 (N_11626,N_11054,N_11055);
or U11627 (N_11627,N_11428,N_11368);
and U11628 (N_11628,N_11035,N_11258);
xor U11629 (N_11629,N_11439,N_11224);
xor U11630 (N_11630,N_11114,N_11228);
nand U11631 (N_11631,N_11144,N_11308);
xnor U11632 (N_11632,N_11452,N_11275);
and U11633 (N_11633,N_11216,N_11003);
and U11634 (N_11634,N_11442,N_11429);
nor U11635 (N_11635,N_11091,N_11447);
or U11636 (N_11636,N_11480,N_11257);
and U11637 (N_11637,N_11226,N_11134);
nor U11638 (N_11638,N_11199,N_11083);
and U11639 (N_11639,N_11128,N_11122);
nor U11640 (N_11640,N_11212,N_11317);
xor U11641 (N_11641,N_11411,N_11383);
nor U11642 (N_11642,N_11084,N_11233);
or U11643 (N_11643,N_11030,N_11025);
xor U11644 (N_11644,N_11096,N_11436);
nand U11645 (N_11645,N_11229,N_11410);
nor U11646 (N_11646,N_11108,N_11405);
xnor U11647 (N_11647,N_11201,N_11278);
nand U11648 (N_11648,N_11048,N_11355);
or U11649 (N_11649,N_11363,N_11490);
nand U11650 (N_11650,N_11090,N_11401);
or U11651 (N_11651,N_11162,N_11058);
xor U11652 (N_11652,N_11295,N_11206);
xnor U11653 (N_11653,N_11449,N_11066);
and U11654 (N_11654,N_11241,N_11240);
and U11655 (N_11655,N_11302,N_11423);
nor U11656 (N_11656,N_11273,N_11130);
and U11657 (N_11657,N_11334,N_11473);
xnor U11658 (N_11658,N_11184,N_11047);
xor U11659 (N_11659,N_11248,N_11381);
and U11660 (N_11660,N_11301,N_11254);
or U11661 (N_11661,N_11415,N_11382);
nor U11662 (N_11662,N_11215,N_11137);
or U11663 (N_11663,N_11351,N_11347);
nand U11664 (N_11664,N_11101,N_11045);
and U11665 (N_11665,N_11336,N_11252);
xnor U11666 (N_11666,N_11022,N_11120);
xor U11667 (N_11667,N_11323,N_11181);
or U11668 (N_11668,N_11471,N_11010);
nor U11669 (N_11669,N_11239,N_11051);
xor U11670 (N_11670,N_11392,N_11220);
nor U11671 (N_11671,N_11486,N_11026);
nor U11672 (N_11672,N_11499,N_11478);
nand U11673 (N_11673,N_11337,N_11064);
nor U11674 (N_11674,N_11357,N_11152);
nor U11675 (N_11675,N_11225,N_11178);
xor U11676 (N_11676,N_11335,N_11221);
nor U11677 (N_11677,N_11082,N_11292);
xnor U11678 (N_11678,N_11349,N_11172);
nand U11679 (N_11679,N_11002,N_11227);
xor U11680 (N_11680,N_11013,N_11018);
or U11681 (N_11681,N_11497,N_11314);
xnor U11682 (N_11682,N_11023,N_11456);
nor U11683 (N_11683,N_11104,N_11358);
or U11684 (N_11684,N_11495,N_11205);
and U11685 (N_11685,N_11356,N_11123);
and U11686 (N_11686,N_11165,N_11059);
or U11687 (N_11687,N_11393,N_11073);
xnor U11688 (N_11688,N_11078,N_11253);
nor U11689 (N_11689,N_11180,N_11197);
nor U11690 (N_11690,N_11419,N_11279);
or U11691 (N_11691,N_11360,N_11033);
or U11692 (N_11692,N_11094,N_11057);
nor U11693 (N_11693,N_11379,N_11440);
xor U11694 (N_11694,N_11367,N_11345);
nand U11695 (N_11695,N_11288,N_11243);
and U11696 (N_11696,N_11259,N_11138);
nor U11697 (N_11697,N_11421,N_11276);
xnor U11698 (N_11698,N_11433,N_11161);
nand U11699 (N_11699,N_11043,N_11008);
nor U11700 (N_11700,N_11136,N_11372);
nor U11701 (N_11701,N_11304,N_11158);
nor U11702 (N_11702,N_11062,N_11294);
nand U11703 (N_11703,N_11268,N_11105);
or U11704 (N_11704,N_11269,N_11369);
and U11705 (N_11705,N_11465,N_11028);
or U11706 (N_11706,N_11307,N_11074);
xor U11707 (N_11707,N_11169,N_11088);
nand U11708 (N_11708,N_11426,N_11441);
xor U11709 (N_11709,N_11213,N_11408);
nor U11710 (N_11710,N_11049,N_11149);
nor U11711 (N_11711,N_11489,N_11282);
nand U11712 (N_11712,N_11009,N_11341);
nand U11713 (N_11713,N_11093,N_11141);
and U11714 (N_11714,N_11316,N_11457);
nand U11715 (N_11715,N_11414,N_11289);
xor U11716 (N_11716,N_11418,N_11089);
or U11717 (N_11717,N_11124,N_11359);
nor U11718 (N_11718,N_11463,N_11305);
xnor U11719 (N_11719,N_11396,N_11448);
or U11720 (N_11720,N_11384,N_11053);
nor U11721 (N_11721,N_11260,N_11398);
nor U11722 (N_11722,N_11328,N_11484);
nand U11723 (N_11723,N_11183,N_11210);
nand U11724 (N_11724,N_11001,N_11453);
nor U11725 (N_11725,N_11006,N_11188);
and U11726 (N_11726,N_11475,N_11092);
nor U11727 (N_11727,N_11060,N_11070);
xor U11728 (N_11728,N_11249,N_11231);
or U11729 (N_11729,N_11324,N_11477);
or U11730 (N_11730,N_11459,N_11309);
nor U11731 (N_11731,N_11479,N_11299);
or U11732 (N_11732,N_11085,N_11195);
nand U11733 (N_11733,N_11238,N_11371);
or U11734 (N_11734,N_11081,N_11126);
and U11735 (N_11735,N_11326,N_11474);
nor U11736 (N_11736,N_11145,N_11193);
xor U11737 (N_11737,N_11217,N_11034);
or U11738 (N_11738,N_11450,N_11483);
and U11739 (N_11739,N_11394,N_11027);
and U11740 (N_11740,N_11329,N_11434);
and U11741 (N_11741,N_11397,N_11388);
nand U11742 (N_11742,N_11044,N_11150);
and U11743 (N_11743,N_11325,N_11245);
nand U11744 (N_11744,N_11103,N_11207);
and U11745 (N_11745,N_11086,N_11116);
nor U11746 (N_11746,N_11485,N_11344);
xor U11747 (N_11747,N_11287,N_11416);
or U11748 (N_11748,N_11179,N_11191);
nor U11749 (N_11749,N_11293,N_11327);
xor U11750 (N_11750,N_11118,N_11133);
nor U11751 (N_11751,N_11304,N_11143);
and U11752 (N_11752,N_11261,N_11121);
and U11753 (N_11753,N_11219,N_11234);
nor U11754 (N_11754,N_11209,N_11383);
or U11755 (N_11755,N_11028,N_11269);
and U11756 (N_11756,N_11265,N_11255);
nor U11757 (N_11757,N_11234,N_11205);
or U11758 (N_11758,N_11413,N_11014);
xor U11759 (N_11759,N_11296,N_11391);
xor U11760 (N_11760,N_11019,N_11416);
xor U11761 (N_11761,N_11232,N_11096);
nand U11762 (N_11762,N_11175,N_11478);
nor U11763 (N_11763,N_11183,N_11344);
or U11764 (N_11764,N_11186,N_11048);
or U11765 (N_11765,N_11063,N_11423);
xnor U11766 (N_11766,N_11416,N_11328);
and U11767 (N_11767,N_11086,N_11300);
xor U11768 (N_11768,N_11378,N_11097);
nor U11769 (N_11769,N_11198,N_11012);
nand U11770 (N_11770,N_11363,N_11163);
nand U11771 (N_11771,N_11328,N_11369);
nor U11772 (N_11772,N_11188,N_11397);
nand U11773 (N_11773,N_11230,N_11264);
nand U11774 (N_11774,N_11310,N_11264);
nor U11775 (N_11775,N_11436,N_11059);
or U11776 (N_11776,N_11381,N_11019);
and U11777 (N_11777,N_11392,N_11007);
nor U11778 (N_11778,N_11482,N_11264);
and U11779 (N_11779,N_11008,N_11200);
or U11780 (N_11780,N_11372,N_11144);
or U11781 (N_11781,N_11090,N_11446);
xor U11782 (N_11782,N_11361,N_11411);
and U11783 (N_11783,N_11103,N_11090);
and U11784 (N_11784,N_11410,N_11265);
and U11785 (N_11785,N_11283,N_11395);
or U11786 (N_11786,N_11136,N_11174);
and U11787 (N_11787,N_11450,N_11435);
nand U11788 (N_11788,N_11170,N_11180);
nor U11789 (N_11789,N_11241,N_11017);
nand U11790 (N_11790,N_11431,N_11382);
or U11791 (N_11791,N_11298,N_11302);
xnor U11792 (N_11792,N_11137,N_11329);
nor U11793 (N_11793,N_11097,N_11425);
or U11794 (N_11794,N_11034,N_11317);
xnor U11795 (N_11795,N_11418,N_11307);
xnor U11796 (N_11796,N_11197,N_11007);
and U11797 (N_11797,N_11484,N_11269);
nand U11798 (N_11798,N_11202,N_11360);
or U11799 (N_11799,N_11266,N_11497);
and U11800 (N_11800,N_11094,N_11409);
xor U11801 (N_11801,N_11384,N_11095);
nor U11802 (N_11802,N_11336,N_11300);
or U11803 (N_11803,N_11383,N_11351);
and U11804 (N_11804,N_11363,N_11432);
or U11805 (N_11805,N_11399,N_11235);
or U11806 (N_11806,N_11328,N_11112);
xnor U11807 (N_11807,N_11421,N_11140);
and U11808 (N_11808,N_11330,N_11110);
nor U11809 (N_11809,N_11309,N_11030);
or U11810 (N_11810,N_11144,N_11184);
or U11811 (N_11811,N_11429,N_11017);
nor U11812 (N_11812,N_11237,N_11387);
nor U11813 (N_11813,N_11331,N_11319);
nor U11814 (N_11814,N_11007,N_11491);
and U11815 (N_11815,N_11437,N_11066);
or U11816 (N_11816,N_11197,N_11216);
nor U11817 (N_11817,N_11154,N_11164);
or U11818 (N_11818,N_11318,N_11192);
and U11819 (N_11819,N_11422,N_11451);
nor U11820 (N_11820,N_11026,N_11189);
and U11821 (N_11821,N_11390,N_11308);
nor U11822 (N_11822,N_11116,N_11470);
and U11823 (N_11823,N_11200,N_11243);
xor U11824 (N_11824,N_11203,N_11079);
nor U11825 (N_11825,N_11066,N_11275);
nor U11826 (N_11826,N_11292,N_11233);
and U11827 (N_11827,N_11325,N_11470);
nand U11828 (N_11828,N_11202,N_11122);
nand U11829 (N_11829,N_11053,N_11157);
or U11830 (N_11830,N_11448,N_11379);
and U11831 (N_11831,N_11352,N_11463);
xnor U11832 (N_11832,N_11195,N_11377);
and U11833 (N_11833,N_11277,N_11291);
and U11834 (N_11834,N_11293,N_11128);
and U11835 (N_11835,N_11021,N_11154);
or U11836 (N_11836,N_11201,N_11269);
nand U11837 (N_11837,N_11155,N_11407);
and U11838 (N_11838,N_11210,N_11258);
and U11839 (N_11839,N_11087,N_11194);
xnor U11840 (N_11840,N_11341,N_11295);
or U11841 (N_11841,N_11327,N_11265);
or U11842 (N_11842,N_11356,N_11049);
nor U11843 (N_11843,N_11087,N_11133);
nor U11844 (N_11844,N_11350,N_11418);
nand U11845 (N_11845,N_11401,N_11012);
or U11846 (N_11846,N_11162,N_11271);
xor U11847 (N_11847,N_11156,N_11082);
or U11848 (N_11848,N_11366,N_11285);
or U11849 (N_11849,N_11368,N_11402);
nor U11850 (N_11850,N_11177,N_11155);
and U11851 (N_11851,N_11389,N_11252);
and U11852 (N_11852,N_11034,N_11146);
and U11853 (N_11853,N_11276,N_11241);
nor U11854 (N_11854,N_11312,N_11157);
or U11855 (N_11855,N_11470,N_11288);
or U11856 (N_11856,N_11178,N_11003);
or U11857 (N_11857,N_11103,N_11039);
and U11858 (N_11858,N_11038,N_11196);
and U11859 (N_11859,N_11247,N_11109);
nor U11860 (N_11860,N_11270,N_11317);
or U11861 (N_11861,N_11332,N_11030);
xnor U11862 (N_11862,N_11410,N_11444);
xor U11863 (N_11863,N_11225,N_11348);
and U11864 (N_11864,N_11192,N_11245);
xnor U11865 (N_11865,N_11025,N_11279);
xor U11866 (N_11866,N_11082,N_11190);
nor U11867 (N_11867,N_11068,N_11108);
nor U11868 (N_11868,N_11481,N_11151);
xnor U11869 (N_11869,N_11192,N_11025);
nor U11870 (N_11870,N_11342,N_11078);
or U11871 (N_11871,N_11327,N_11400);
or U11872 (N_11872,N_11231,N_11100);
xor U11873 (N_11873,N_11471,N_11110);
xor U11874 (N_11874,N_11436,N_11367);
xnor U11875 (N_11875,N_11496,N_11378);
or U11876 (N_11876,N_11271,N_11223);
or U11877 (N_11877,N_11311,N_11394);
and U11878 (N_11878,N_11082,N_11164);
and U11879 (N_11879,N_11483,N_11319);
nor U11880 (N_11880,N_11351,N_11152);
or U11881 (N_11881,N_11015,N_11370);
or U11882 (N_11882,N_11249,N_11206);
nor U11883 (N_11883,N_11167,N_11450);
nand U11884 (N_11884,N_11360,N_11209);
nor U11885 (N_11885,N_11004,N_11139);
nand U11886 (N_11886,N_11162,N_11188);
and U11887 (N_11887,N_11147,N_11199);
nand U11888 (N_11888,N_11311,N_11186);
nand U11889 (N_11889,N_11334,N_11204);
or U11890 (N_11890,N_11265,N_11067);
nand U11891 (N_11891,N_11090,N_11321);
xnor U11892 (N_11892,N_11489,N_11161);
nand U11893 (N_11893,N_11209,N_11314);
nor U11894 (N_11894,N_11417,N_11313);
or U11895 (N_11895,N_11208,N_11104);
and U11896 (N_11896,N_11268,N_11442);
nand U11897 (N_11897,N_11159,N_11234);
xor U11898 (N_11898,N_11479,N_11451);
nor U11899 (N_11899,N_11474,N_11252);
nand U11900 (N_11900,N_11044,N_11234);
or U11901 (N_11901,N_11384,N_11219);
or U11902 (N_11902,N_11486,N_11280);
and U11903 (N_11903,N_11018,N_11397);
or U11904 (N_11904,N_11331,N_11486);
nor U11905 (N_11905,N_11069,N_11208);
nor U11906 (N_11906,N_11244,N_11406);
nor U11907 (N_11907,N_11136,N_11166);
or U11908 (N_11908,N_11050,N_11060);
nand U11909 (N_11909,N_11269,N_11071);
nor U11910 (N_11910,N_11352,N_11314);
and U11911 (N_11911,N_11001,N_11421);
nand U11912 (N_11912,N_11302,N_11354);
nor U11913 (N_11913,N_11297,N_11331);
and U11914 (N_11914,N_11048,N_11011);
xor U11915 (N_11915,N_11415,N_11159);
nor U11916 (N_11916,N_11451,N_11285);
and U11917 (N_11917,N_11174,N_11365);
xor U11918 (N_11918,N_11040,N_11439);
nand U11919 (N_11919,N_11201,N_11429);
nor U11920 (N_11920,N_11293,N_11303);
nor U11921 (N_11921,N_11128,N_11147);
and U11922 (N_11922,N_11213,N_11067);
xor U11923 (N_11923,N_11154,N_11351);
nand U11924 (N_11924,N_11180,N_11255);
nor U11925 (N_11925,N_11183,N_11153);
or U11926 (N_11926,N_11471,N_11144);
or U11927 (N_11927,N_11479,N_11437);
or U11928 (N_11928,N_11418,N_11408);
or U11929 (N_11929,N_11335,N_11155);
nand U11930 (N_11930,N_11078,N_11252);
or U11931 (N_11931,N_11011,N_11151);
and U11932 (N_11932,N_11378,N_11067);
and U11933 (N_11933,N_11399,N_11492);
nand U11934 (N_11934,N_11353,N_11269);
nand U11935 (N_11935,N_11029,N_11083);
nand U11936 (N_11936,N_11364,N_11421);
and U11937 (N_11937,N_11012,N_11342);
xnor U11938 (N_11938,N_11317,N_11063);
and U11939 (N_11939,N_11404,N_11479);
xor U11940 (N_11940,N_11044,N_11304);
or U11941 (N_11941,N_11350,N_11495);
xor U11942 (N_11942,N_11417,N_11071);
or U11943 (N_11943,N_11283,N_11157);
and U11944 (N_11944,N_11466,N_11128);
and U11945 (N_11945,N_11028,N_11089);
or U11946 (N_11946,N_11334,N_11090);
or U11947 (N_11947,N_11089,N_11227);
nor U11948 (N_11948,N_11006,N_11068);
nand U11949 (N_11949,N_11410,N_11193);
and U11950 (N_11950,N_11423,N_11444);
nand U11951 (N_11951,N_11372,N_11220);
and U11952 (N_11952,N_11167,N_11334);
xnor U11953 (N_11953,N_11389,N_11430);
xnor U11954 (N_11954,N_11170,N_11042);
xnor U11955 (N_11955,N_11112,N_11393);
or U11956 (N_11956,N_11084,N_11046);
nand U11957 (N_11957,N_11437,N_11232);
and U11958 (N_11958,N_11026,N_11163);
xnor U11959 (N_11959,N_11198,N_11191);
nand U11960 (N_11960,N_11104,N_11350);
and U11961 (N_11961,N_11430,N_11147);
xnor U11962 (N_11962,N_11165,N_11452);
and U11963 (N_11963,N_11007,N_11358);
or U11964 (N_11964,N_11224,N_11009);
or U11965 (N_11965,N_11325,N_11182);
xor U11966 (N_11966,N_11106,N_11468);
or U11967 (N_11967,N_11387,N_11435);
nor U11968 (N_11968,N_11352,N_11304);
nor U11969 (N_11969,N_11011,N_11133);
nand U11970 (N_11970,N_11115,N_11029);
nor U11971 (N_11971,N_11391,N_11340);
nand U11972 (N_11972,N_11365,N_11139);
and U11973 (N_11973,N_11217,N_11419);
or U11974 (N_11974,N_11249,N_11280);
xnor U11975 (N_11975,N_11122,N_11198);
or U11976 (N_11976,N_11230,N_11392);
and U11977 (N_11977,N_11079,N_11053);
or U11978 (N_11978,N_11171,N_11466);
xor U11979 (N_11979,N_11308,N_11243);
or U11980 (N_11980,N_11050,N_11271);
nand U11981 (N_11981,N_11380,N_11399);
nand U11982 (N_11982,N_11380,N_11297);
and U11983 (N_11983,N_11408,N_11357);
xor U11984 (N_11984,N_11138,N_11460);
xor U11985 (N_11985,N_11052,N_11177);
or U11986 (N_11986,N_11447,N_11067);
nor U11987 (N_11987,N_11432,N_11392);
and U11988 (N_11988,N_11160,N_11190);
nand U11989 (N_11989,N_11493,N_11364);
nor U11990 (N_11990,N_11040,N_11207);
xor U11991 (N_11991,N_11214,N_11480);
or U11992 (N_11992,N_11491,N_11134);
nand U11993 (N_11993,N_11118,N_11221);
and U11994 (N_11994,N_11476,N_11432);
nor U11995 (N_11995,N_11440,N_11362);
xor U11996 (N_11996,N_11315,N_11317);
and U11997 (N_11997,N_11489,N_11313);
or U11998 (N_11998,N_11166,N_11301);
xor U11999 (N_11999,N_11252,N_11065);
nand U12000 (N_12000,N_11696,N_11649);
nor U12001 (N_12001,N_11887,N_11772);
nor U12002 (N_12002,N_11503,N_11642);
nor U12003 (N_12003,N_11656,N_11505);
xnor U12004 (N_12004,N_11980,N_11581);
nand U12005 (N_12005,N_11888,N_11645);
nor U12006 (N_12006,N_11660,N_11698);
nor U12007 (N_12007,N_11913,N_11557);
xor U12008 (N_12008,N_11543,N_11626);
nand U12009 (N_12009,N_11640,N_11765);
nor U12010 (N_12010,N_11542,N_11578);
and U12011 (N_12011,N_11742,N_11925);
and U12012 (N_12012,N_11554,N_11516);
nor U12013 (N_12013,N_11988,N_11868);
xnor U12014 (N_12014,N_11709,N_11527);
xor U12015 (N_12015,N_11630,N_11540);
and U12016 (N_12016,N_11504,N_11832);
or U12017 (N_12017,N_11892,N_11606);
or U12018 (N_12018,N_11890,N_11561);
and U12019 (N_12019,N_11762,N_11549);
and U12020 (N_12020,N_11811,N_11735);
and U12021 (N_12021,N_11781,N_11625);
xnor U12022 (N_12022,N_11595,N_11593);
and U12023 (N_12023,N_11634,N_11694);
nand U12024 (N_12024,N_11893,N_11759);
or U12025 (N_12025,N_11960,N_11512);
nor U12026 (N_12026,N_11619,N_11989);
nor U12027 (N_12027,N_11914,N_11760);
xor U12028 (N_12028,N_11835,N_11663);
and U12029 (N_12029,N_11718,N_11858);
and U12030 (N_12030,N_11929,N_11854);
or U12031 (N_12031,N_11629,N_11790);
xor U12032 (N_12032,N_11987,N_11917);
and U12033 (N_12033,N_11876,N_11627);
nor U12034 (N_12034,N_11921,N_11599);
xor U12035 (N_12035,N_11767,N_11721);
and U12036 (N_12036,N_11782,N_11970);
xor U12037 (N_12037,N_11613,N_11607);
xor U12038 (N_12038,N_11618,N_11550);
xnor U12039 (N_12039,N_11936,N_11776);
xnor U12040 (N_12040,N_11834,N_11779);
xor U12041 (N_12041,N_11555,N_11878);
nor U12042 (N_12042,N_11666,N_11730);
nor U12043 (N_12043,N_11902,N_11639);
nand U12044 (N_12044,N_11836,N_11553);
and U12045 (N_12045,N_11682,N_11792);
and U12046 (N_12046,N_11529,N_11611);
nand U12047 (N_12047,N_11753,N_11590);
nand U12048 (N_12048,N_11658,N_11506);
nand U12049 (N_12049,N_11954,N_11693);
nand U12050 (N_12050,N_11648,N_11756);
nor U12051 (N_12051,N_11522,N_11908);
or U12052 (N_12052,N_11563,N_11885);
nor U12053 (N_12053,N_11799,N_11794);
xnor U12054 (N_12054,N_11801,N_11855);
xnor U12055 (N_12055,N_11701,N_11712);
nand U12056 (N_12056,N_11728,N_11500);
and U12057 (N_12057,N_11707,N_11570);
or U12058 (N_12058,N_11872,N_11580);
or U12059 (N_12059,N_11907,N_11915);
nand U12060 (N_12060,N_11729,N_11999);
and U12061 (N_12061,N_11865,N_11846);
nand U12062 (N_12062,N_11797,N_11817);
or U12063 (N_12063,N_11830,N_11819);
or U12064 (N_12064,N_11995,N_11602);
and U12065 (N_12065,N_11699,N_11726);
or U12066 (N_12066,N_11866,N_11705);
or U12067 (N_12067,N_11652,N_11795);
nor U12068 (N_12068,N_11820,N_11669);
and U12069 (N_12069,N_11644,N_11831);
and U12070 (N_12070,N_11856,N_11654);
and U12071 (N_12071,N_11850,N_11774);
or U12072 (N_12072,N_11918,N_11558);
or U12073 (N_12073,N_11508,N_11899);
nor U12074 (N_12074,N_11556,N_11873);
nor U12075 (N_12075,N_11968,N_11577);
xnor U12076 (N_12076,N_11814,N_11998);
xor U12077 (N_12077,N_11862,N_11604);
nand U12078 (N_12078,N_11686,N_11646);
nand U12079 (N_12079,N_11881,N_11897);
nand U12080 (N_12080,N_11965,N_11572);
nand U12081 (N_12081,N_11547,N_11631);
xnor U12082 (N_12082,N_11871,N_11636);
xnor U12083 (N_12083,N_11879,N_11976);
and U12084 (N_12084,N_11757,N_11904);
nor U12085 (N_12085,N_11743,N_11773);
nor U12086 (N_12086,N_11544,N_11708);
xnor U12087 (N_12087,N_11853,N_11906);
and U12088 (N_12088,N_11661,N_11741);
nand U12089 (N_12089,N_11972,N_11905);
and U12090 (N_12090,N_11867,N_11538);
or U12091 (N_12091,N_11518,N_11515);
or U12092 (N_12092,N_11677,N_11585);
or U12093 (N_12093,N_11755,N_11937);
or U12094 (N_12094,N_11628,N_11901);
nand U12095 (N_12095,N_11588,N_11943);
xnor U12096 (N_12096,N_11884,N_11513);
and U12097 (N_12097,N_11732,N_11610);
or U12098 (N_12098,N_11821,N_11617);
xnor U12099 (N_12099,N_11812,N_11993);
xnor U12100 (N_12100,N_11546,N_11584);
nand U12101 (N_12101,N_11796,N_11637);
or U12102 (N_12102,N_11818,N_11775);
or U12103 (N_12103,N_11545,N_11829);
and U12104 (N_12104,N_11955,N_11752);
xor U12105 (N_12105,N_11502,N_11785);
xnor U12106 (N_12106,N_11870,N_11891);
nor U12107 (N_12107,N_11573,N_11882);
nor U12108 (N_12108,N_11739,N_11662);
xor U12109 (N_12109,N_11964,N_11690);
and U12110 (N_12110,N_11715,N_11851);
and U12111 (N_12111,N_11804,N_11719);
nand U12112 (N_12112,N_11982,N_11950);
nand U12113 (N_12113,N_11717,N_11938);
or U12114 (N_12114,N_11751,N_11519);
nand U12115 (N_12115,N_11525,N_11569);
or U12116 (N_12116,N_11837,N_11736);
or U12117 (N_12117,N_11843,N_11744);
nor U12118 (N_12118,N_11521,N_11911);
nor U12119 (N_12119,N_11552,N_11576);
nand U12120 (N_12120,N_11511,N_11841);
or U12121 (N_12121,N_11994,N_11940);
nand U12122 (N_12122,N_11621,N_11520);
or U12123 (N_12123,N_11746,N_11874);
nor U12124 (N_12124,N_11671,N_11838);
or U12125 (N_12125,N_11716,N_11849);
nor U12126 (N_12126,N_11952,N_11883);
or U12127 (N_12127,N_11860,N_11798);
and U12128 (N_12128,N_11605,N_11623);
or U12129 (N_12129,N_11608,N_11571);
nand U12130 (N_12130,N_11591,N_11784);
nor U12131 (N_12131,N_11771,N_11963);
and U12132 (N_12132,N_11909,N_11979);
nand U12133 (N_12133,N_11526,N_11926);
or U12134 (N_12134,N_11806,N_11560);
xor U12135 (N_12135,N_11803,N_11778);
nand U12136 (N_12136,N_11749,N_11859);
xnor U12137 (N_12137,N_11780,N_11766);
and U12138 (N_12138,N_11761,N_11704);
nand U12139 (N_12139,N_11793,N_11548);
xor U12140 (N_12140,N_11676,N_11802);
and U12141 (N_12141,N_11714,N_11864);
nor U12142 (N_12142,N_11598,N_11592);
or U12143 (N_12143,N_11533,N_11655);
nor U12144 (N_12144,N_11847,N_11641);
nand U12145 (N_12145,N_11857,N_11895);
nand U12146 (N_12146,N_11532,N_11510);
or U12147 (N_12147,N_11653,N_11934);
and U12148 (N_12148,N_11680,N_11931);
xnor U12149 (N_12149,N_11981,N_11703);
xnor U12150 (N_12150,N_11638,N_11966);
or U12151 (N_12151,N_11758,N_11537);
or U12152 (N_12152,N_11842,N_11531);
or U12153 (N_12153,N_11800,N_11973);
and U12154 (N_12154,N_11528,N_11657);
and U12155 (N_12155,N_11582,N_11863);
or U12156 (N_12156,N_11562,N_11579);
or U12157 (N_12157,N_11957,N_11996);
nand U12158 (N_12158,N_11684,N_11622);
nand U12159 (N_12159,N_11689,N_11947);
and U12160 (N_12160,N_11674,N_11787);
xor U12161 (N_12161,N_11647,N_11861);
or U12162 (N_12162,N_11928,N_11738);
or U12163 (N_12163,N_11589,N_11734);
xor U12164 (N_12164,N_11668,N_11534);
and U12165 (N_12165,N_11675,N_11783);
and U12166 (N_12166,N_11731,N_11889);
and U12167 (N_12167,N_11535,N_11935);
and U12168 (N_12168,N_11609,N_11808);
xor U12169 (N_12169,N_11985,N_11961);
nor U12170 (N_12170,N_11737,N_11596);
and U12171 (N_12171,N_11975,N_11825);
or U12172 (N_12172,N_11810,N_11681);
or U12173 (N_12173,N_11791,N_11769);
xor U12174 (N_12174,N_11650,N_11962);
or U12175 (N_12175,N_11706,N_11969);
and U12176 (N_12176,N_11786,N_11939);
nor U12177 (N_12177,N_11710,N_11594);
nand U12178 (N_12178,N_11539,N_11824);
xor U12179 (N_12179,N_11956,N_11984);
or U12180 (N_12180,N_11501,N_11815);
nor U12181 (N_12181,N_11740,N_11659);
xor U12182 (N_12182,N_11635,N_11840);
nor U12183 (N_12183,N_11691,N_11685);
xor U12184 (N_12184,N_11983,N_11932);
nor U12185 (N_12185,N_11930,N_11839);
nand U12186 (N_12186,N_11551,N_11945);
or U12187 (N_12187,N_11789,N_11823);
xor U12188 (N_12188,N_11978,N_11898);
nor U12189 (N_12189,N_11614,N_11844);
xnor U12190 (N_12190,N_11875,N_11764);
nand U12191 (N_12191,N_11967,N_11651);
nor U12192 (N_12192,N_11949,N_11948);
xnor U12193 (N_12193,N_11941,N_11700);
nand U12194 (N_12194,N_11683,N_11670);
xnor U12195 (N_12195,N_11679,N_11927);
and U12196 (N_12196,N_11992,N_11828);
and U12197 (N_12197,N_11869,N_11687);
xnor U12198 (N_12198,N_11807,N_11903);
nor U12199 (N_12199,N_11665,N_11568);
nand U12200 (N_12200,N_11991,N_11722);
and U12201 (N_12201,N_11564,N_11946);
nor U12202 (N_12202,N_11507,N_11620);
nand U12203 (N_12203,N_11974,N_11959);
nor U12204 (N_12204,N_11697,N_11541);
nand U12205 (N_12205,N_11986,N_11951);
and U12206 (N_12206,N_11920,N_11845);
nor U12207 (N_12207,N_11509,N_11664);
nor U12208 (N_12208,N_11816,N_11750);
or U12209 (N_12209,N_11805,N_11944);
nand U12210 (N_12210,N_11612,N_11536);
nor U12211 (N_12211,N_11530,N_11601);
nand U12212 (N_12212,N_11667,N_11997);
nand U12213 (N_12213,N_11673,N_11809);
or U12214 (N_12214,N_11632,N_11894);
xnor U12215 (N_12215,N_11942,N_11748);
nand U12216 (N_12216,N_11692,N_11924);
xor U12217 (N_12217,N_11616,N_11788);
nor U12218 (N_12218,N_11745,N_11559);
xor U12219 (N_12219,N_11770,N_11713);
nand U12220 (N_12220,N_11923,N_11896);
or U12221 (N_12221,N_11754,N_11886);
and U12222 (N_12222,N_11524,N_11910);
nand U12223 (N_12223,N_11724,N_11565);
xor U12224 (N_12224,N_11615,N_11678);
and U12225 (N_12225,N_11597,N_11723);
nand U12226 (N_12226,N_11953,N_11912);
or U12227 (N_12227,N_11768,N_11826);
or U12228 (N_12228,N_11747,N_11958);
and U12229 (N_12229,N_11725,N_11933);
and U12230 (N_12230,N_11971,N_11633);
and U12231 (N_12231,N_11813,N_11586);
or U12232 (N_12232,N_11575,N_11695);
xor U12233 (N_12233,N_11566,N_11574);
and U12234 (N_12234,N_11733,N_11643);
xor U12235 (N_12235,N_11514,N_11624);
nand U12236 (N_12236,N_11977,N_11777);
nor U12237 (N_12237,N_11833,N_11900);
or U12238 (N_12238,N_11711,N_11916);
xor U12239 (N_12239,N_11567,N_11827);
xor U12240 (N_12240,N_11600,N_11852);
and U12241 (N_12241,N_11583,N_11702);
xnor U12242 (N_12242,N_11688,N_11523);
xnor U12243 (N_12243,N_11672,N_11877);
and U12244 (N_12244,N_11720,N_11880);
nor U12245 (N_12245,N_11848,N_11517);
nand U12246 (N_12246,N_11822,N_11763);
nor U12247 (N_12247,N_11727,N_11587);
nor U12248 (N_12248,N_11990,N_11919);
and U12249 (N_12249,N_11922,N_11603);
or U12250 (N_12250,N_11627,N_11817);
nand U12251 (N_12251,N_11500,N_11914);
nor U12252 (N_12252,N_11834,N_11520);
and U12253 (N_12253,N_11750,N_11721);
nor U12254 (N_12254,N_11610,N_11523);
xor U12255 (N_12255,N_11567,N_11786);
or U12256 (N_12256,N_11714,N_11870);
or U12257 (N_12257,N_11672,N_11821);
nor U12258 (N_12258,N_11667,N_11628);
nand U12259 (N_12259,N_11542,N_11777);
xor U12260 (N_12260,N_11571,N_11536);
nor U12261 (N_12261,N_11880,N_11746);
nor U12262 (N_12262,N_11768,N_11510);
and U12263 (N_12263,N_11627,N_11795);
xor U12264 (N_12264,N_11882,N_11618);
or U12265 (N_12265,N_11548,N_11926);
nand U12266 (N_12266,N_11568,N_11907);
nor U12267 (N_12267,N_11855,N_11790);
and U12268 (N_12268,N_11657,N_11712);
nor U12269 (N_12269,N_11612,N_11945);
and U12270 (N_12270,N_11519,N_11587);
or U12271 (N_12271,N_11761,N_11532);
and U12272 (N_12272,N_11752,N_11725);
xor U12273 (N_12273,N_11817,N_11578);
or U12274 (N_12274,N_11884,N_11846);
or U12275 (N_12275,N_11995,N_11920);
nor U12276 (N_12276,N_11728,N_11710);
and U12277 (N_12277,N_11879,N_11627);
or U12278 (N_12278,N_11917,N_11587);
or U12279 (N_12279,N_11643,N_11587);
xor U12280 (N_12280,N_11931,N_11956);
or U12281 (N_12281,N_11808,N_11945);
nor U12282 (N_12282,N_11896,N_11726);
xnor U12283 (N_12283,N_11615,N_11670);
nand U12284 (N_12284,N_11582,N_11638);
and U12285 (N_12285,N_11748,N_11596);
or U12286 (N_12286,N_11991,N_11807);
or U12287 (N_12287,N_11623,N_11782);
or U12288 (N_12288,N_11626,N_11852);
or U12289 (N_12289,N_11898,N_11897);
or U12290 (N_12290,N_11967,N_11902);
nand U12291 (N_12291,N_11846,N_11526);
or U12292 (N_12292,N_11814,N_11586);
or U12293 (N_12293,N_11561,N_11875);
nand U12294 (N_12294,N_11673,N_11589);
nor U12295 (N_12295,N_11659,N_11705);
xnor U12296 (N_12296,N_11555,N_11551);
xor U12297 (N_12297,N_11674,N_11796);
nand U12298 (N_12298,N_11833,N_11915);
xnor U12299 (N_12299,N_11976,N_11573);
or U12300 (N_12300,N_11911,N_11509);
or U12301 (N_12301,N_11681,N_11927);
nor U12302 (N_12302,N_11812,N_11645);
or U12303 (N_12303,N_11592,N_11532);
or U12304 (N_12304,N_11787,N_11981);
and U12305 (N_12305,N_11549,N_11996);
nand U12306 (N_12306,N_11541,N_11512);
nor U12307 (N_12307,N_11868,N_11929);
or U12308 (N_12308,N_11710,N_11522);
nand U12309 (N_12309,N_11501,N_11579);
or U12310 (N_12310,N_11930,N_11953);
nor U12311 (N_12311,N_11588,N_11549);
and U12312 (N_12312,N_11847,N_11592);
xnor U12313 (N_12313,N_11821,N_11759);
or U12314 (N_12314,N_11651,N_11598);
nand U12315 (N_12315,N_11772,N_11706);
and U12316 (N_12316,N_11766,N_11806);
or U12317 (N_12317,N_11986,N_11689);
or U12318 (N_12318,N_11513,N_11960);
and U12319 (N_12319,N_11604,N_11772);
xor U12320 (N_12320,N_11954,N_11845);
nor U12321 (N_12321,N_11528,N_11904);
nand U12322 (N_12322,N_11897,N_11757);
xor U12323 (N_12323,N_11521,N_11919);
xor U12324 (N_12324,N_11988,N_11995);
xor U12325 (N_12325,N_11614,N_11981);
xor U12326 (N_12326,N_11646,N_11609);
or U12327 (N_12327,N_11890,N_11705);
nand U12328 (N_12328,N_11882,N_11802);
and U12329 (N_12329,N_11537,N_11769);
xnor U12330 (N_12330,N_11607,N_11647);
and U12331 (N_12331,N_11787,N_11501);
or U12332 (N_12332,N_11568,N_11633);
and U12333 (N_12333,N_11833,N_11599);
and U12334 (N_12334,N_11829,N_11704);
and U12335 (N_12335,N_11871,N_11534);
xor U12336 (N_12336,N_11760,N_11593);
and U12337 (N_12337,N_11884,N_11768);
and U12338 (N_12338,N_11882,N_11863);
xor U12339 (N_12339,N_11574,N_11970);
xor U12340 (N_12340,N_11676,N_11539);
and U12341 (N_12341,N_11614,N_11698);
nor U12342 (N_12342,N_11865,N_11520);
and U12343 (N_12343,N_11717,N_11909);
nand U12344 (N_12344,N_11705,N_11581);
xnor U12345 (N_12345,N_11939,N_11985);
and U12346 (N_12346,N_11535,N_11889);
or U12347 (N_12347,N_11634,N_11861);
xnor U12348 (N_12348,N_11690,N_11925);
and U12349 (N_12349,N_11702,N_11691);
nor U12350 (N_12350,N_11972,N_11881);
nor U12351 (N_12351,N_11748,N_11743);
nor U12352 (N_12352,N_11573,N_11829);
xnor U12353 (N_12353,N_11663,N_11526);
nand U12354 (N_12354,N_11764,N_11530);
and U12355 (N_12355,N_11648,N_11527);
and U12356 (N_12356,N_11739,N_11525);
or U12357 (N_12357,N_11727,N_11757);
and U12358 (N_12358,N_11938,N_11798);
nand U12359 (N_12359,N_11734,N_11890);
and U12360 (N_12360,N_11700,N_11534);
nand U12361 (N_12361,N_11660,N_11725);
or U12362 (N_12362,N_11668,N_11505);
nand U12363 (N_12363,N_11661,N_11521);
nand U12364 (N_12364,N_11583,N_11621);
or U12365 (N_12365,N_11927,N_11719);
or U12366 (N_12366,N_11692,N_11898);
xnor U12367 (N_12367,N_11697,N_11826);
nor U12368 (N_12368,N_11577,N_11928);
xnor U12369 (N_12369,N_11662,N_11944);
nand U12370 (N_12370,N_11930,N_11518);
nand U12371 (N_12371,N_11563,N_11782);
nand U12372 (N_12372,N_11720,N_11914);
or U12373 (N_12373,N_11704,N_11673);
nand U12374 (N_12374,N_11950,N_11717);
nand U12375 (N_12375,N_11871,N_11751);
or U12376 (N_12376,N_11754,N_11820);
xor U12377 (N_12377,N_11872,N_11676);
nand U12378 (N_12378,N_11796,N_11987);
nand U12379 (N_12379,N_11506,N_11992);
nor U12380 (N_12380,N_11793,N_11816);
nor U12381 (N_12381,N_11902,N_11781);
or U12382 (N_12382,N_11712,N_11634);
nor U12383 (N_12383,N_11868,N_11524);
and U12384 (N_12384,N_11590,N_11622);
or U12385 (N_12385,N_11743,N_11851);
nor U12386 (N_12386,N_11808,N_11982);
nor U12387 (N_12387,N_11685,N_11611);
nor U12388 (N_12388,N_11674,N_11818);
nand U12389 (N_12389,N_11644,N_11502);
nor U12390 (N_12390,N_11706,N_11580);
nor U12391 (N_12391,N_11666,N_11769);
nand U12392 (N_12392,N_11547,N_11764);
nor U12393 (N_12393,N_11912,N_11588);
and U12394 (N_12394,N_11931,N_11520);
xor U12395 (N_12395,N_11901,N_11510);
or U12396 (N_12396,N_11714,N_11576);
xnor U12397 (N_12397,N_11875,N_11820);
and U12398 (N_12398,N_11929,N_11746);
or U12399 (N_12399,N_11669,N_11612);
nor U12400 (N_12400,N_11958,N_11691);
and U12401 (N_12401,N_11510,N_11897);
xnor U12402 (N_12402,N_11683,N_11625);
nand U12403 (N_12403,N_11639,N_11624);
nor U12404 (N_12404,N_11617,N_11532);
nand U12405 (N_12405,N_11976,N_11996);
nand U12406 (N_12406,N_11555,N_11884);
nand U12407 (N_12407,N_11689,N_11736);
nand U12408 (N_12408,N_11581,N_11656);
and U12409 (N_12409,N_11831,N_11916);
nand U12410 (N_12410,N_11924,N_11703);
xor U12411 (N_12411,N_11683,N_11781);
nand U12412 (N_12412,N_11688,N_11805);
nand U12413 (N_12413,N_11514,N_11950);
nand U12414 (N_12414,N_11822,N_11592);
xor U12415 (N_12415,N_11796,N_11550);
nor U12416 (N_12416,N_11616,N_11726);
or U12417 (N_12417,N_11856,N_11977);
nor U12418 (N_12418,N_11541,N_11945);
and U12419 (N_12419,N_11770,N_11873);
nand U12420 (N_12420,N_11828,N_11576);
or U12421 (N_12421,N_11631,N_11912);
and U12422 (N_12422,N_11761,N_11833);
xor U12423 (N_12423,N_11553,N_11920);
nor U12424 (N_12424,N_11547,N_11758);
nand U12425 (N_12425,N_11507,N_11773);
and U12426 (N_12426,N_11522,N_11672);
or U12427 (N_12427,N_11643,N_11922);
nand U12428 (N_12428,N_11732,N_11797);
or U12429 (N_12429,N_11532,N_11681);
xor U12430 (N_12430,N_11538,N_11593);
nor U12431 (N_12431,N_11819,N_11799);
xor U12432 (N_12432,N_11649,N_11820);
xor U12433 (N_12433,N_11726,N_11859);
nor U12434 (N_12434,N_11759,N_11854);
and U12435 (N_12435,N_11568,N_11515);
xnor U12436 (N_12436,N_11739,N_11522);
xor U12437 (N_12437,N_11571,N_11678);
or U12438 (N_12438,N_11685,N_11853);
nor U12439 (N_12439,N_11842,N_11736);
xnor U12440 (N_12440,N_11818,N_11710);
or U12441 (N_12441,N_11578,N_11678);
or U12442 (N_12442,N_11715,N_11886);
xnor U12443 (N_12443,N_11638,N_11613);
nor U12444 (N_12444,N_11707,N_11562);
nand U12445 (N_12445,N_11605,N_11652);
nor U12446 (N_12446,N_11671,N_11628);
nor U12447 (N_12447,N_11800,N_11779);
nor U12448 (N_12448,N_11742,N_11744);
or U12449 (N_12449,N_11990,N_11868);
or U12450 (N_12450,N_11842,N_11652);
xnor U12451 (N_12451,N_11504,N_11956);
nand U12452 (N_12452,N_11958,N_11671);
and U12453 (N_12453,N_11925,N_11824);
xor U12454 (N_12454,N_11568,N_11816);
and U12455 (N_12455,N_11587,N_11918);
and U12456 (N_12456,N_11691,N_11746);
nand U12457 (N_12457,N_11522,N_11944);
nand U12458 (N_12458,N_11743,N_11758);
nor U12459 (N_12459,N_11613,N_11976);
nor U12460 (N_12460,N_11500,N_11602);
nand U12461 (N_12461,N_11762,N_11802);
and U12462 (N_12462,N_11939,N_11922);
nand U12463 (N_12463,N_11728,N_11785);
nand U12464 (N_12464,N_11817,N_11505);
and U12465 (N_12465,N_11669,N_11519);
and U12466 (N_12466,N_11510,N_11669);
nand U12467 (N_12467,N_11600,N_11885);
or U12468 (N_12468,N_11748,N_11719);
or U12469 (N_12469,N_11783,N_11916);
nand U12470 (N_12470,N_11770,N_11749);
or U12471 (N_12471,N_11940,N_11910);
and U12472 (N_12472,N_11614,N_11760);
xor U12473 (N_12473,N_11844,N_11838);
nand U12474 (N_12474,N_11969,N_11525);
xor U12475 (N_12475,N_11635,N_11762);
nand U12476 (N_12476,N_11911,N_11506);
nor U12477 (N_12477,N_11951,N_11665);
nor U12478 (N_12478,N_11728,N_11667);
xor U12479 (N_12479,N_11888,N_11752);
and U12480 (N_12480,N_11921,N_11535);
and U12481 (N_12481,N_11548,N_11929);
xor U12482 (N_12482,N_11762,N_11818);
xor U12483 (N_12483,N_11724,N_11658);
xor U12484 (N_12484,N_11596,N_11584);
nor U12485 (N_12485,N_11571,N_11638);
or U12486 (N_12486,N_11671,N_11797);
nand U12487 (N_12487,N_11984,N_11842);
or U12488 (N_12488,N_11601,N_11783);
and U12489 (N_12489,N_11622,N_11730);
xor U12490 (N_12490,N_11893,N_11701);
nor U12491 (N_12491,N_11829,N_11607);
and U12492 (N_12492,N_11760,N_11823);
or U12493 (N_12493,N_11689,N_11822);
xor U12494 (N_12494,N_11594,N_11598);
or U12495 (N_12495,N_11642,N_11920);
nor U12496 (N_12496,N_11882,N_11973);
nand U12497 (N_12497,N_11831,N_11973);
nand U12498 (N_12498,N_11625,N_11568);
xor U12499 (N_12499,N_11786,N_11823);
nand U12500 (N_12500,N_12310,N_12008);
xor U12501 (N_12501,N_12375,N_12267);
nor U12502 (N_12502,N_12296,N_12161);
nor U12503 (N_12503,N_12291,N_12016);
xnor U12504 (N_12504,N_12341,N_12305);
and U12505 (N_12505,N_12404,N_12303);
nor U12506 (N_12506,N_12211,N_12055);
or U12507 (N_12507,N_12402,N_12293);
and U12508 (N_12508,N_12027,N_12236);
or U12509 (N_12509,N_12198,N_12365);
or U12510 (N_12510,N_12227,N_12197);
or U12511 (N_12511,N_12485,N_12014);
nor U12512 (N_12512,N_12112,N_12141);
and U12513 (N_12513,N_12186,N_12472);
nand U12514 (N_12514,N_12177,N_12041);
nand U12515 (N_12515,N_12244,N_12328);
or U12516 (N_12516,N_12152,N_12459);
xor U12517 (N_12517,N_12462,N_12194);
and U12518 (N_12518,N_12460,N_12321);
xnor U12519 (N_12519,N_12376,N_12201);
or U12520 (N_12520,N_12160,N_12077);
or U12521 (N_12521,N_12486,N_12349);
nand U12522 (N_12522,N_12277,N_12458);
and U12523 (N_12523,N_12325,N_12348);
or U12524 (N_12524,N_12115,N_12171);
xor U12525 (N_12525,N_12276,N_12097);
or U12526 (N_12526,N_12265,N_12421);
xnor U12527 (N_12527,N_12024,N_12213);
xor U12528 (N_12528,N_12253,N_12260);
nand U12529 (N_12529,N_12364,N_12167);
nand U12530 (N_12530,N_12354,N_12423);
or U12531 (N_12531,N_12337,N_12367);
or U12532 (N_12532,N_12436,N_12250);
nand U12533 (N_12533,N_12398,N_12051);
nor U12534 (N_12534,N_12268,N_12382);
nor U12535 (N_12535,N_12129,N_12195);
xnor U12536 (N_12536,N_12280,N_12451);
or U12537 (N_12537,N_12353,N_12079);
nor U12538 (N_12538,N_12053,N_12358);
nand U12539 (N_12539,N_12146,N_12220);
and U12540 (N_12540,N_12448,N_12380);
xor U12541 (N_12541,N_12180,N_12271);
nand U12542 (N_12542,N_12003,N_12093);
and U12543 (N_12543,N_12062,N_12431);
and U12544 (N_12544,N_12206,N_12479);
or U12545 (N_12545,N_12158,N_12435);
and U12546 (N_12546,N_12470,N_12287);
xnor U12547 (N_12547,N_12307,N_12111);
nor U12548 (N_12548,N_12099,N_12314);
nor U12549 (N_12549,N_12105,N_12281);
or U12550 (N_12550,N_12335,N_12480);
and U12551 (N_12551,N_12336,N_12165);
nand U12552 (N_12552,N_12103,N_12481);
or U12553 (N_12553,N_12425,N_12025);
or U12554 (N_12554,N_12350,N_12407);
nand U12555 (N_12555,N_12187,N_12444);
nor U12556 (N_12556,N_12173,N_12301);
or U12557 (N_12557,N_12339,N_12015);
xor U12558 (N_12558,N_12330,N_12441);
xor U12559 (N_12559,N_12168,N_12096);
nor U12560 (N_12560,N_12128,N_12032);
or U12561 (N_12561,N_12484,N_12315);
nand U12562 (N_12562,N_12332,N_12379);
nand U12563 (N_12563,N_12148,N_12216);
nand U12564 (N_12564,N_12355,N_12020);
xor U12565 (N_12565,N_12333,N_12429);
xnor U12566 (N_12566,N_12151,N_12499);
and U12567 (N_12567,N_12316,N_12174);
xnor U12568 (N_12568,N_12179,N_12474);
or U12569 (N_12569,N_12278,N_12043);
nand U12570 (N_12570,N_12106,N_12284);
or U12571 (N_12571,N_12400,N_12469);
and U12572 (N_12572,N_12192,N_12150);
or U12573 (N_12573,N_12114,N_12292);
nor U12574 (N_12574,N_12210,N_12492);
nand U12575 (N_12575,N_12411,N_12274);
xor U12576 (N_12576,N_12401,N_12455);
or U12577 (N_12577,N_12313,N_12413);
xnor U12578 (N_12578,N_12231,N_12100);
or U12579 (N_12579,N_12011,N_12362);
and U12580 (N_12580,N_12245,N_12306);
or U12581 (N_12581,N_12243,N_12422);
nor U12582 (N_12582,N_12496,N_12266);
xor U12583 (N_12583,N_12030,N_12075);
and U12584 (N_12584,N_12002,N_12416);
xor U12585 (N_12585,N_12230,N_12110);
nor U12586 (N_12586,N_12054,N_12483);
or U12587 (N_12587,N_12338,N_12312);
nand U12588 (N_12588,N_12098,N_12249);
or U12589 (N_12589,N_12345,N_12252);
or U12590 (N_12590,N_12371,N_12241);
nor U12591 (N_12591,N_12139,N_12369);
xnor U12592 (N_12592,N_12395,N_12482);
or U12593 (N_12593,N_12162,N_12092);
or U12594 (N_12594,N_12246,N_12392);
nor U12595 (N_12595,N_12304,N_12351);
and U12596 (N_12596,N_12359,N_12127);
and U12597 (N_12597,N_12466,N_12327);
nand U12598 (N_12598,N_12397,N_12142);
nand U12599 (N_12599,N_12428,N_12120);
xnor U12600 (N_12600,N_12403,N_12270);
xnor U12601 (N_12601,N_12282,N_12056);
or U12602 (N_12602,N_12089,N_12399);
xnor U12603 (N_12603,N_12119,N_12334);
nor U12604 (N_12604,N_12134,N_12001);
nand U12605 (N_12605,N_12294,N_12144);
xnor U12606 (N_12606,N_12193,N_12045);
nor U12607 (N_12607,N_12132,N_12487);
xnor U12608 (N_12608,N_12452,N_12035);
or U12609 (N_12609,N_12137,N_12476);
nor U12610 (N_12610,N_12248,N_12450);
nor U12611 (N_12611,N_12417,N_12176);
nand U12612 (N_12612,N_12122,N_12237);
xnor U12613 (N_12613,N_12497,N_12059);
xnor U12614 (N_12614,N_12238,N_12084);
xnor U12615 (N_12615,N_12409,N_12021);
nor U12616 (N_12616,N_12204,N_12317);
nand U12617 (N_12617,N_12135,N_12078);
nand U12618 (N_12618,N_12205,N_12124);
xnor U12619 (N_12619,N_12288,N_12060);
xor U12620 (N_12620,N_12360,N_12390);
and U12621 (N_12621,N_12036,N_12082);
and U12622 (N_12622,N_12473,N_12368);
nand U12623 (N_12623,N_12214,N_12387);
or U12624 (N_12624,N_12117,N_12298);
xnor U12625 (N_12625,N_12088,N_12071);
or U12626 (N_12626,N_12415,N_12203);
and U12627 (N_12627,N_12494,N_12275);
and U12628 (N_12628,N_12131,N_12223);
or U12629 (N_12629,N_12070,N_12440);
nand U12630 (N_12630,N_12269,N_12190);
or U12631 (N_12631,N_12004,N_12263);
nor U12632 (N_12632,N_12290,N_12286);
and U12633 (N_12633,N_12229,N_12430);
xnor U12634 (N_12634,N_12145,N_12361);
nor U12635 (N_12635,N_12199,N_12342);
or U12636 (N_12636,N_12189,N_12121);
or U12637 (N_12637,N_12136,N_12491);
nand U12638 (N_12638,N_12299,N_12068);
or U12639 (N_12639,N_12493,N_12057);
or U12640 (N_12640,N_12373,N_12490);
and U12641 (N_12641,N_12226,N_12295);
or U12642 (N_12642,N_12356,N_12069);
or U12643 (N_12643,N_12309,N_12258);
xor U12644 (N_12644,N_12381,N_12104);
xnor U12645 (N_12645,N_12155,N_12076);
or U12646 (N_12646,N_12495,N_12156);
nand U12647 (N_12647,N_12118,N_12443);
nor U12648 (N_12648,N_12394,N_12219);
nor U12649 (N_12649,N_12464,N_12461);
nand U12650 (N_12650,N_12026,N_12233);
nand U12651 (N_12651,N_12363,N_12023);
nand U12652 (N_12652,N_12209,N_12101);
or U12653 (N_12653,N_12251,N_12391);
and U12654 (N_12654,N_12357,N_12449);
or U12655 (N_12655,N_12018,N_12273);
xnor U12656 (N_12656,N_12346,N_12157);
nor U12657 (N_12657,N_12169,N_12300);
xnor U12658 (N_12658,N_12065,N_12182);
nor U12659 (N_12659,N_12159,N_12225);
nor U12660 (N_12660,N_12326,N_12329);
nand U12661 (N_12661,N_12471,N_12467);
xnor U12662 (N_12662,N_12366,N_12447);
nand U12663 (N_12663,N_12384,N_12164);
nand U12664 (N_12664,N_12324,N_12412);
or U12665 (N_12665,N_12090,N_12038);
nand U12666 (N_12666,N_12012,N_12072);
nor U12667 (N_12667,N_12283,N_12005);
and U12668 (N_12668,N_12279,N_12039);
xnor U12669 (N_12669,N_12109,N_12130);
or U12670 (N_12670,N_12427,N_12311);
or U12671 (N_12671,N_12224,N_12228);
xor U12672 (N_12672,N_12261,N_12445);
xor U12673 (N_12673,N_12116,N_12302);
nor U12674 (N_12674,N_12297,N_12221);
and U12675 (N_12675,N_12419,N_12331);
xor U12676 (N_12676,N_12029,N_12086);
nor U12677 (N_12677,N_12031,N_12347);
or U12678 (N_12678,N_12143,N_12457);
nor U12679 (N_12679,N_12085,N_12138);
or U12680 (N_12680,N_12439,N_12405);
xor U12681 (N_12681,N_12212,N_12061);
and U12682 (N_12682,N_12170,N_12377);
xnor U12683 (N_12683,N_12048,N_12126);
xor U12684 (N_12684,N_12178,N_12388);
xnor U12685 (N_12685,N_12442,N_12000);
or U12686 (N_12686,N_12235,N_12185);
nor U12687 (N_12687,N_12166,N_12477);
nand U12688 (N_12688,N_12083,N_12149);
nor U12689 (N_12689,N_12172,N_12108);
and U12690 (N_12690,N_12344,N_12247);
and U12691 (N_12691,N_12370,N_12389);
xor U12692 (N_12692,N_12222,N_12010);
and U12693 (N_12693,N_12208,N_12022);
or U12694 (N_12694,N_12123,N_12322);
nand U12695 (N_12695,N_12113,N_12285);
and U12696 (N_12696,N_12107,N_12013);
nor U12697 (N_12697,N_12232,N_12259);
nor U12698 (N_12698,N_12207,N_12067);
nor U12699 (N_12699,N_12262,N_12468);
xnor U12700 (N_12700,N_12396,N_12319);
nor U12701 (N_12701,N_12308,N_12033);
nand U12702 (N_12702,N_12006,N_12087);
nor U12703 (N_12703,N_12385,N_12181);
xnor U12704 (N_12704,N_12017,N_12153);
nor U12705 (N_12705,N_12408,N_12218);
and U12706 (N_12706,N_12386,N_12066);
and U12707 (N_12707,N_12410,N_12133);
and U12708 (N_12708,N_12047,N_12264);
nand U12709 (N_12709,N_12343,N_12091);
xnor U12710 (N_12710,N_12256,N_12372);
or U12711 (N_12711,N_12163,N_12257);
or U12712 (N_12712,N_12489,N_12465);
nor U12713 (N_12713,N_12034,N_12406);
xor U12714 (N_12714,N_12046,N_12196);
nor U12715 (N_12715,N_12217,N_12378);
nand U12716 (N_12716,N_12463,N_12432);
and U12717 (N_12717,N_12074,N_12175);
or U12718 (N_12718,N_12318,N_12255);
nand U12719 (N_12719,N_12140,N_12456);
xnor U12720 (N_12720,N_12289,N_12446);
nand U12721 (N_12721,N_12239,N_12191);
xor U12722 (N_12722,N_12094,N_12374);
and U12723 (N_12723,N_12147,N_12475);
nand U12724 (N_12724,N_12414,N_12418);
nor U12725 (N_12725,N_12454,N_12340);
or U12726 (N_12726,N_12040,N_12202);
xnor U12727 (N_12727,N_12437,N_12073);
or U12728 (N_12728,N_12050,N_12352);
or U12729 (N_12729,N_12028,N_12080);
nor U12730 (N_12730,N_12007,N_12063);
nand U12731 (N_12731,N_12240,N_12323);
and U12732 (N_12732,N_12234,N_12052);
nand U12733 (N_12733,N_12393,N_12044);
or U12734 (N_12734,N_12037,N_12426);
xor U12735 (N_12735,N_12242,N_12188);
nand U12736 (N_12736,N_12058,N_12042);
xor U12737 (N_12737,N_12183,N_12498);
nor U12738 (N_12738,N_12009,N_12434);
nor U12739 (N_12739,N_12424,N_12081);
or U12740 (N_12740,N_12200,N_12272);
nor U12741 (N_12741,N_12019,N_12478);
or U12742 (N_12742,N_12095,N_12184);
and U12743 (N_12743,N_12453,N_12064);
and U12744 (N_12744,N_12154,N_12102);
nor U12745 (N_12745,N_12254,N_12420);
nand U12746 (N_12746,N_12320,N_12215);
xor U12747 (N_12747,N_12125,N_12438);
nand U12748 (N_12748,N_12049,N_12433);
nand U12749 (N_12749,N_12383,N_12488);
and U12750 (N_12750,N_12010,N_12430);
xor U12751 (N_12751,N_12230,N_12472);
xor U12752 (N_12752,N_12173,N_12029);
xor U12753 (N_12753,N_12085,N_12257);
nand U12754 (N_12754,N_12043,N_12145);
nand U12755 (N_12755,N_12277,N_12058);
and U12756 (N_12756,N_12329,N_12159);
xor U12757 (N_12757,N_12268,N_12331);
or U12758 (N_12758,N_12102,N_12376);
and U12759 (N_12759,N_12231,N_12395);
or U12760 (N_12760,N_12075,N_12231);
nor U12761 (N_12761,N_12104,N_12286);
nor U12762 (N_12762,N_12370,N_12441);
or U12763 (N_12763,N_12303,N_12372);
xnor U12764 (N_12764,N_12228,N_12443);
or U12765 (N_12765,N_12479,N_12414);
nor U12766 (N_12766,N_12269,N_12439);
nor U12767 (N_12767,N_12193,N_12088);
or U12768 (N_12768,N_12180,N_12479);
nand U12769 (N_12769,N_12042,N_12320);
or U12770 (N_12770,N_12184,N_12303);
xnor U12771 (N_12771,N_12125,N_12087);
xor U12772 (N_12772,N_12429,N_12205);
or U12773 (N_12773,N_12313,N_12266);
or U12774 (N_12774,N_12318,N_12333);
xnor U12775 (N_12775,N_12268,N_12313);
nand U12776 (N_12776,N_12427,N_12315);
xnor U12777 (N_12777,N_12447,N_12251);
xnor U12778 (N_12778,N_12468,N_12493);
nor U12779 (N_12779,N_12206,N_12055);
or U12780 (N_12780,N_12069,N_12154);
or U12781 (N_12781,N_12353,N_12311);
nand U12782 (N_12782,N_12326,N_12035);
or U12783 (N_12783,N_12200,N_12228);
or U12784 (N_12784,N_12186,N_12102);
xnor U12785 (N_12785,N_12354,N_12199);
nand U12786 (N_12786,N_12072,N_12041);
nand U12787 (N_12787,N_12395,N_12097);
and U12788 (N_12788,N_12364,N_12061);
or U12789 (N_12789,N_12169,N_12438);
nor U12790 (N_12790,N_12378,N_12233);
nor U12791 (N_12791,N_12120,N_12261);
and U12792 (N_12792,N_12001,N_12383);
and U12793 (N_12793,N_12017,N_12369);
nand U12794 (N_12794,N_12467,N_12233);
xor U12795 (N_12795,N_12170,N_12057);
nor U12796 (N_12796,N_12452,N_12374);
and U12797 (N_12797,N_12062,N_12301);
nand U12798 (N_12798,N_12408,N_12018);
and U12799 (N_12799,N_12266,N_12037);
nor U12800 (N_12800,N_12415,N_12206);
nor U12801 (N_12801,N_12170,N_12195);
and U12802 (N_12802,N_12443,N_12355);
and U12803 (N_12803,N_12009,N_12471);
nor U12804 (N_12804,N_12263,N_12459);
xnor U12805 (N_12805,N_12446,N_12154);
xnor U12806 (N_12806,N_12131,N_12370);
nor U12807 (N_12807,N_12163,N_12141);
xnor U12808 (N_12808,N_12083,N_12028);
nor U12809 (N_12809,N_12219,N_12326);
nand U12810 (N_12810,N_12395,N_12474);
nand U12811 (N_12811,N_12425,N_12109);
nand U12812 (N_12812,N_12170,N_12139);
nand U12813 (N_12813,N_12162,N_12179);
xor U12814 (N_12814,N_12086,N_12251);
nand U12815 (N_12815,N_12211,N_12121);
and U12816 (N_12816,N_12090,N_12374);
and U12817 (N_12817,N_12062,N_12245);
nor U12818 (N_12818,N_12477,N_12247);
or U12819 (N_12819,N_12019,N_12203);
nor U12820 (N_12820,N_12147,N_12195);
and U12821 (N_12821,N_12442,N_12365);
xnor U12822 (N_12822,N_12379,N_12292);
nor U12823 (N_12823,N_12004,N_12202);
or U12824 (N_12824,N_12402,N_12317);
or U12825 (N_12825,N_12451,N_12389);
nor U12826 (N_12826,N_12064,N_12363);
or U12827 (N_12827,N_12426,N_12188);
and U12828 (N_12828,N_12120,N_12156);
or U12829 (N_12829,N_12444,N_12163);
nor U12830 (N_12830,N_12011,N_12320);
nor U12831 (N_12831,N_12376,N_12342);
or U12832 (N_12832,N_12340,N_12220);
nand U12833 (N_12833,N_12080,N_12289);
xor U12834 (N_12834,N_12205,N_12110);
xnor U12835 (N_12835,N_12198,N_12488);
xnor U12836 (N_12836,N_12136,N_12193);
xnor U12837 (N_12837,N_12229,N_12471);
and U12838 (N_12838,N_12180,N_12203);
xor U12839 (N_12839,N_12300,N_12066);
xor U12840 (N_12840,N_12408,N_12280);
or U12841 (N_12841,N_12302,N_12076);
or U12842 (N_12842,N_12001,N_12253);
and U12843 (N_12843,N_12328,N_12174);
nor U12844 (N_12844,N_12334,N_12133);
or U12845 (N_12845,N_12134,N_12038);
or U12846 (N_12846,N_12005,N_12111);
and U12847 (N_12847,N_12416,N_12087);
xnor U12848 (N_12848,N_12163,N_12342);
nand U12849 (N_12849,N_12112,N_12437);
xnor U12850 (N_12850,N_12336,N_12004);
xor U12851 (N_12851,N_12386,N_12024);
nand U12852 (N_12852,N_12109,N_12245);
xor U12853 (N_12853,N_12327,N_12214);
or U12854 (N_12854,N_12344,N_12271);
xor U12855 (N_12855,N_12391,N_12355);
nand U12856 (N_12856,N_12237,N_12056);
or U12857 (N_12857,N_12304,N_12064);
and U12858 (N_12858,N_12250,N_12274);
and U12859 (N_12859,N_12389,N_12484);
nor U12860 (N_12860,N_12116,N_12414);
nand U12861 (N_12861,N_12081,N_12281);
or U12862 (N_12862,N_12402,N_12254);
xnor U12863 (N_12863,N_12341,N_12259);
xnor U12864 (N_12864,N_12469,N_12436);
nor U12865 (N_12865,N_12163,N_12279);
xnor U12866 (N_12866,N_12141,N_12197);
nor U12867 (N_12867,N_12249,N_12167);
xor U12868 (N_12868,N_12383,N_12164);
nand U12869 (N_12869,N_12304,N_12111);
nor U12870 (N_12870,N_12061,N_12021);
nand U12871 (N_12871,N_12281,N_12195);
and U12872 (N_12872,N_12440,N_12408);
nor U12873 (N_12873,N_12000,N_12327);
xor U12874 (N_12874,N_12110,N_12347);
or U12875 (N_12875,N_12250,N_12327);
or U12876 (N_12876,N_12322,N_12494);
or U12877 (N_12877,N_12092,N_12009);
xor U12878 (N_12878,N_12303,N_12223);
nand U12879 (N_12879,N_12123,N_12146);
or U12880 (N_12880,N_12115,N_12421);
nand U12881 (N_12881,N_12202,N_12368);
and U12882 (N_12882,N_12181,N_12361);
nand U12883 (N_12883,N_12488,N_12155);
nand U12884 (N_12884,N_12017,N_12024);
xnor U12885 (N_12885,N_12488,N_12058);
nand U12886 (N_12886,N_12450,N_12162);
and U12887 (N_12887,N_12330,N_12421);
or U12888 (N_12888,N_12459,N_12082);
or U12889 (N_12889,N_12301,N_12119);
xor U12890 (N_12890,N_12008,N_12082);
nor U12891 (N_12891,N_12410,N_12083);
and U12892 (N_12892,N_12022,N_12395);
nand U12893 (N_12893,N_12116,N_12383);
nor U12894 (N_12894,N_12471,N_12079);
xnor U12895 (N_12895,N_12180,N_12372);
nor U12896 (N_12896,N_12342,N_12330);
xnor U12897 (N_12897,N_12463,N_12429);
nand U12898 (N_12898,N_12181,N_12407);
or U12899 (N_12899,N_12480,N_12448);
nand U12900 (N_12900,N_12154,N_12245);
nand U12901 (N_12901,N_12399,N_12484);
xnor U12902 (N_12902,N_12479,N_12300);
or U12903 (N_12903,N_12458,N_12016);
xnor U12904 (N_12904,N_12221,N_12239);
and U12905 (N_12905,N_12281,N_12385);
nand U12906 (N_12906,N_12393,N_12333);
xor U12907 (N_12907,N_12221,N_12436);
xnor U12908 (N_12908,N_12275,N_12288);
nor U12909 (N_12909,N_12168,N_12106);
nor U12910 (N_12910,N_12370,N_12082);
or U12911 (N_12911,N_12010,N_12323);
or U12912 (N_12912,N_12417,N_12108);
or U12913 (N_12913,N_12439,N_12222);
nand U12914 (N_12914,N_12287,N_12154);
or U12915 (N_12915,N_12250,N_12106);
xnor U12916 (N_12916,N_12361,N_12285);
and U12917 (N_12917,N_12072,N_12255);
and U12918 (N_12918,N_12049,N_12228);
nor U12919 (N_12919,N_12195,N_12051);
nand U12920 (N_12920,N_12351,N_12346);
nand U12921 (N_12921,N_12424,N_12202);
xnor U12922 (N_12922,N_12318,N_12079);
xor U12923 (N_12923,N_12028,N_12134);
nor U12924 (N_12924,N_12133,N_12037);
and U12925 (N_12925,N_12398,N_12322);
nand U12926 (N_12926,N_12151,N_12200);
xor U12927 (N_12927,N_12388,N_12229);
xnor U12928 (N_12928,N_12359,N_12344);
nand U12929 (N_12929,N_12437,N_12247);
nor U12930 (N_12930,N_12469,N_12113);
nor U12931 (N_12931,N_12082,N_12278);
or U12932 (N_12932,N_12198,N_12122);
or U12933 (N_12933,N_12498,N_12115);
and U12934 (N_12934,N_12449,N_12284);
and U12935 (N_12935,N_12275,N_12255);
nor U12936 (N_12936,N_12099,N_12119);
nand U12937 (N_12937,N_12049,N_12414);
nor U12938 (N_12938,N_12049,N_12051);
xor U12939 (N_12939,N_12384,N_12114);
and U12940 (N_12940,N_12442,N_12450);
nand U12941 (N_12941,N_12120,N_12031);
and U12942 (N_12942,N_12145,N_12161);
or U12943 (N_12943,N_12116,N_12270);
nand U12944 (N_12944,N_12060,N_12180);
or U12945 (N_12945,N_12391,N_12328);
xor U12946 (N_12946,N_12392,N_12081);
and U12947 (N_12947,N_12020,N_12011);
and U12948 (N_12948,N_12134,N_12224);
nand U12949 (N_12949,N_12374,N_12407);
nand U12950 (N_12950,N_12245,N_12114);
nand U12951 (N_12951,N_12076,N_12147);
xnor U12952 (N_12952,N_12062,N_12261);
nor U12953 (N_12953,N_12340,N_12183);
nor U12954 (N_12954,N_12339,N_12470);
xor U12955 (N_12955,N_12049,N_12352);
xnor U12956 (N_12956,N_12280,N_12351);
and U12957 (N_12957,N_12004,N_12354);
nand U12958 (N_12958,N_12391,N_12439);
or U12959 (N_12959,N_12180,N_12127);
and U12960 (N_12960,N_12031,N_12221);
xor U12961 (N_12961,N_12200,N_12291);
or U12962 (N_12962,N_12285,N_12247);
nand U12963 (N_12963,N_12317,N_12357);
and U12964 (N_12964,N_12423,N_12230);
or U12965 (N_12965,N_12205,N_12023);
xor U12966 (N_12966,N_12012,N_12340);
and U12967 (N_12967,N_12360,N_12447);
nand U12968 (N_12968,N_12125,N_12029);
nor U12969 (N_12969,N_12383,N_12020);
and U12970 (N_12970,N_12216,N_12060);
xnor U12971 (N_12971,N_12049,N_12156);
nor U12972 (N_12972,N_12355,N_12070);
nand U12973 (N_12973,N_12437,N_12225);
or U12974 (N_12974,N_12179,N_12290);
and U12975 (N_12975,N_12344,N_12222);
nor U12976 (N_12976,N_12052,N_12360);
and U12977 (N_12977,N_12146,N_12200);
or U12978 (N_12978,N_12212,N_12284);
xor U12979 (N_12979,N_12275,N_12294);
xor U12980 (N_12980,N_12463,N_12471);
nor U12981 (N_12981,N_12121,N_12481);
xor U12982 (N_12982,N_12039,N_12145);
nor U12983 (N_12983,N_12499,N_12177);
and U12984 (N_12984,N_12264,N_12461);
nor U12985 (N_12985,N_12394,N_12171);
nor U12986 (N_12986,N_12456,N_12062);
xor U12987 (N_12987,N_12140,N_12417);
nand U12988 (N_12988,N_12449,N_12341);
nor U12989 (N_12989,N_12101,N_12276);
nor U12990 (N_12990,N_12372,N_12022);
nor U12991 (N_12991,N_12214,N_12242);
and U12992 (N_12992,N_12482,N_12102);
and U12993 (N_12993,N_12093,N_12182);
and U12994 (N_12994,N_12067,N_12076);
and U12995 (N_12995,N_12155,N_12337);
nor U12996 (N_12996,N_12288,N_12382);
nor U12997 (N_12997,N_12267,N_12131);
or U12998 (N_12998,N_12247,N_12240);
or U12999 (N_12999,N_12245,N_12061);
and U13000 (N_13000,N_12959,N_12525);
and U13001 (N_13001,N_12947,N_12572);
nor U13002 (N_13002,N_12526,N_12948);
xor U13003 (N_13003,N_12570,N_12528);
nand U13004 (N_13004,N_12730,N_12835);
nor U13005 (N_13005,N_12882,N_12825);
nand U13006 (N_13006,N_12575,N_12551);
or U13007 (N_13007,N_12544,N_12993);
and U13008 (N_13008,N_12776,N_12591);
nand U13009 (N_13009,N_12890,N_12650);
nand U13010 (N_13010,N_12606,N_12777);
xor U13011 (N_13011,N_12695,N_12571);
xor U13012 (N_13012,N_12949,N_12703);
nor U13013 (N_13013,N_12712,N_12964);
or U13014 (N_13014,N_12660,N_12589);
and U13015 (N_13015,N_12880,N_12532);
xor U13016 (N_13016,N_12738,N_12837);
or U13017 (N_13017,N_12663,N_12578);
and U13018 (N_13018,N_12697,N_12809);
xor U13019 (N_13019,N_12594,N_12597);
xnor U13020 (N_13020,N_12855,N_12656);
nor U13021 (N_13021,N_12966,N_12520);
nand U13022 (N_13022,N_12917,N_12553);
nor U13023 (N_13023,N_12740,N_12834);
and U13024 (N_13024,N_12931,N_12613);
and U13025 (N_13025,N_12951,N_12543);
or U13026 (N_13026,N_12652,N_12793);
xnor U13027 (N_13027,N_12794,N_12599);
nor U13028 (N_13028,N_12512,N_12534);
nand U13029 (N_13029,N_12554,N_12546);
or U13030 (N_13030,N_12506,N_12886);
or U13031 (N_13031,N_12742,N_12724);
xnor U13032 (N_13032,N_12896,N_12617);
xnor U13033 (N_13033,N_12582,N_12604);
and U13034 (N_13034,N_12971,N_12874);
and U13035 (N_13035,N_12782,N_12845);
nor U13036 (N_13036,N_12826,N_12545);
and U13037 (N_13037,N_12561,N_12997);
and U13038 (N_13038,N_12502,N_12622);
and U13039 (N_13039,N_12875,N_12945);
nor U13040 (N_13040,N_12692,N_12583);
nor U13041 (N_13041,N_12722,N_12979);
or U13042 (N_13042,N_12668,N_12511);
xnor U13043 (N_13043,N_12610,N_12967);
nor U13044 (N_13044,N_12999,N_12641);
nor U13045 (N_13045,N_12555,N_12704);
nor U13046 (N_13046,N_12649,N_12535);
nor U13047 (N_13047,N_12976,N_12864);
nand U13048 (N_13048,N_12667,N_12500);
xor U13049 (N_13049,N_12625,N_12743);
nor U13050 (N_13050,N_12521,N_12923);
nand U13051 (N_13051,N_12892,N_12618);
nor U13052 (N_13052,N_12548,N_12974);
nand U13053 (N_13053,N_12932,N_12728);
or U13054 (N_13054,N_12560,N_12763);
xor U13055 (N_13055,N_12564,N_12600);
xnor U13056 (N_13056,N_12795,N_12889);
nor U13057 (N_13057,N_12566,N_12920);
and U13058 (N_13058,N_12647,N_12779);
or U13059 (N_13059,N_12873,N_12860);
nand U13060 (N_13060,N_12662,N_12879);
nor U13061 (N_13061,N_12760,N_12579);
and U13062 (N_13062,N_12638,N_12508);
xnor U13063 (N_13063,N_12933,N_12877);
nor U13064 (N_13064,N_12513,N_12585);
and U13065 (N_13065,N_12669,N_12861);
and U13066 (N_13066,N_12928,N_12624);
xor U13067 (N_13067,N_12698,N_12772);
or U13068 (N_13068,N_12659,N_12941);
xnor U13069 (N_13069,N_12858,N_12620);
nand U13070 (N_13070,N_12637,N_12567);
xor U13071 (N_13071,N_12986,N_12792);
nor U13072 (N_13072,N_12975,N_12628);
nor U13073 (N_13073,N_12727,N_12876);
nor U13074 (N_13074,N_12770,N_12745);
and U13075 (N_13075,N_12842,N_12717);
nand U13076 (N_13076,N_12934,N_12644);
and U13077 (N_13077,N_12693,N_12725);
and U13078 (N_13078,N_12800,N_12953);
xnor U13079 (N_13079,N_12501,N_12994);
nor U13080 (N_13080,N_12574,N_12987);
nor U13081 (N_13081,N_12847,N_12655);
and U13082 (N_13082,N_12653,N_12819);
xor U13083 (N_13083,N_12988,N_12853);
nor U13084 (N_13084,N_12666,N_12801);
xor U13085 (N_13085,N_12780,N_12516);
nand U13086 (N_13086,N_12630,N_12689);
nor U13087 (N_13087,N_12831,N_12903);
xor U13088 (N_13088,N_12510,N_12705);
xnor U13089 (N_13089,N_12621,N_12899);
or U13090 (N_13090,N_12626,N_12642);
nor U13091 (N_13091,N_12867,N_12900);
nor U13092 (N_13092,N_12552,N_12542);
nor U13093 (N_13093,N_12752,N_12539);
nand U13094 (N_13094,N_12588,N_12865);
or U13095 (N_13095,N_12901,N_12957);
xnor U13096 (N_13096,N_12848,N_12814);
nand U13097 (N_13097,N_12887,N_12691);
xnor U13098 (N_13098,N_12563,N_12716);
and U13099 (N_13099,N_12584,N_12758);
xor U13100 (N_13100,N_12962,N_12774);
nand U13101 (N_13101,N_12911,N_12746);
and U13102 (N_13102,N_12768,N_12839);
nand U13103 (N_13103,N_12737,N_12784);
nand U13104 (N_13104,N_12682,N_12507);
and U13105 (N_13105,N_12816,N_12576);
nor U13106 (N_13106,N_12778,N_12913);
and U13107 (N_13107,N_12658,N_12843);
xnor U13108 (N_13108,N_12970,N_12872);
nand U13109 (N_13109,N_12568,N_12519);
nor U13110 (N_13110,N_12905,N_12940);
or U13111 (N_13111,N_12771,N_12714);
or U13112 (N_13112,N_12824,N_12925);
and U13113 (N_13113,N_12851,N_12690);
nand U13114 (N_13114,N_12969,N_12830);
nand U13115 (N_13115,N_12844,N_12643);
or U13116 (N_13116,N_12919,N_12651);
xor U13117 (N_13117,N_12537,N_12696);
nor U13118 (N_13118,N_12836,N_12587);
nand U13119 (N_13119,N_12893,N_12744);
and U13120 (N_13120,N_12881,N_12805);
nor U13121 (N_13121,N_12687,N_12927);
or U13122 (N_13122,N_12884,N_12912);
and U13123 (N_13123,N_12736,N_12810);
or U13124 (N_13124,N_12870,N_12577);
nand U13125 (N_13125,N_12765,N_12751);
and U13126 (N_13126,N_12973,N_12895);
nor U13127 (N_13127,N_12918,N_12868);
nand U13128 (N_13128,N_12812,N_12661);
and U13129 (N_13129,N_12950,N_12926);
or U13130 (N_13130,N_12846,N_12711);
or U13131 (N_13131,N_12929,N_12935);
nor U13132 (N_13132,N_12632,N_12798);
and U13133 (N_13133,N_12531,N_12883);
or U13134 (N_13134,N_12503,N_12955);
and U13135 (N_13135,N_12657,N_12761);
and U13136 (N_13136,N_12715,N_12517);
and U13137 (N_13137,N_12985,N_12978);
xnor U13138 (N_13138,N_12700,N_12523);
and U13139 (N_13139,N_12827,N_12963);
nor U13140 (N_13140,N_12720,N_12958);
nand U13141 (N_13141,N_12527,N_12766);
nor U13142 (N_13142,N_12791,N_12592);
or U13143 (N_13143,N_12671,N_12995);
and U13144 (N_13144,N_12541,N_12665);
xor U13145 (N_13145,N_12909,N_12767);
nand U13146 (N_13146,N_12598,N_12707);
and U13147 (N_13147,N_12802,N_12863);
or U13148 (N_13148,N_12673,N_12747);
or U13149 (N_13149,N_12869,N_12732);
and U13150 (N_13150,N_12960,N_12939);
xor U13151 (N_13151,N_12936,N_12965);
nand U13152 (N_13152,N_12908,N_12759);
and U13153 (N_13153,N_12675,N_12547);
nand U13154 (N_13154,N_12590,N_12762);
nor U13155 (N_13155,N_12756,N_12701);
and U13156 (N_13156,N_12862,N_12924);
nor U13157 (N_13157,N_12937,N_12674);
xnor U13158 (N_13158,N_12734,N_12664);
and U13159 (N_13159,N_12823,N_12757);
nor U13160 (N_13160,N_12921,N_12954);
and U13161 (N_13161,N_12529,N_12681);
and U13162 (N_13162,N_12533,N_12788);
xor U13163 (N_13163,N_12914,N_12731);
and U13164 (N_13164,N_12946,N_12938);
xor U13165 (N_13165,N_12719,N_12898);
nand U13166 (N_13166,N_12559,N_12748);
xor U13167 (N_13167,N_12557,N_12634);
nand U13168 (N_13168,N_12708,N_12565);
and U13169 (N_13169,N_12619,N_12904);
nand U13170 (N_13170,N_12885,N_12808);
or U13171 (N_13171,N_12854,N_12556);
and U13172 (N_13172,N_12749,N_12850);
and U13173 (N_13173,N_12683,N_12857);
nor U13174 (N_13174,N_12549,N_12741);
nor U13175 (N_13175,N_12968,N_12943);
nor U13176 (N_13176,N_12721,N_12633);
and U13177 (N_13177,N_12755,N_12670);
and U13178 (N_13178,N_12787,N_12573);
nand U13179 (N_13179,N_12856,N_12569);
nor U13180 (N_13180,N_12645,N_12789);
and U13181 (N_13181,N_12723,N_12612);
xor U13182 (N_13182,N_12739,N_12609);
nor U13183 (N_13183,N_12676,N_12803);
or U13184 (N_13184,N_12894,N_12790);
nand U13185 (N_13185,N_12849,N_12603);
nor U13186 (N_13186,N_12694,N_12991);
nand U13187 (N_13187,N_12735,N_12733);
and U13188 (N_13188,N_12804,N_12605);
xor U13189 (N_13189,N_12518,N_12709);
nand U13190 (N_13190,N_12829,N_12684);
and U13191 (N_13191,N_12702,N_12891);
nor U13192 (N_13192,N_12828,N_12852);
nand U13193 (N_13193,N_12706,N_12718);
and U13194 (N_13194,N_12635,N_12907);
xnor U13195 (N_13195,N_12593,N_12930);
nor U13196 (N_13196,N_12504,N_12984);
xnor U13197 (N_13197,N_12640,N_12980);
nand U13198 (N_13198,N_12538,N_12942);
nand U13199 (N_13199,N_12944,N_12977);
or U13200 (N_13200,N_12841,N_12639);
xor U13201 (N_13201,N_12781,N_12678);
and U13202 (N_13202,N_12813,N_12614);
nand U13203 (N_13203,N_12595,N_12818);
nor U13204 (N_13204,N_12680,N_12688);
xor U13205 (N_13205,N_12611,N_12580);
nor U13206 (N_13206,N_12998,N_12910);
xnor U13207 (N_13207,N_12710,N_12769);
or U13208 (N_13208,N_12811,N_12602);
xor U13209 (N_13209,N_12726,N_12775);
nand U13210 (N_13210,N_12536,N_12822);
or U13211 (N_13211,N_12956,N_12820);
nor U13212 (N_13212,N_12996,N_12509);
xnor U13213 (N_13213,N_12952,N_12888);
and U13214 (N_13214,N_12972,N_12562);
or U13215 (N_13215,N_12922,N_12785);
or U13216 (N_13216,N_12897,N_12783);
nand U13217 (N_13217,N_12729,N_12859);
or U13218 (N_13218,N_12679,N_12550);
and U13219 (N_13219,N_12832,N_12514);
or U13220 (N_13220,N_12807,N_12608);
nor U13221 (N_13221,N_12821,N_12631);
or U13222 (N_13222,N_12586,N_12636);
nand U13223 (N_13223,N_12815,N_12754);
nor U13224 (N_13224,N_12786,N_12982);
nor U13225 (N_13225,N_12629,N_12685);
nor U13226 (N_13226,N_12581,N_12866);
and U13227 (N_13227,N_12558,N_12796);
nor U13228 (N_13228,N_12764,N_12833);
or U13229 (N_13229,N_12992,N_12990);
and U13230 (N_13230,N_12961,N_12648);
nand U13231 (N_13231,N_12915,N_12983);
xnor U13232 (N_13232,N_12524,N_12878);
and U13233 (N_13233,N_12750,N_12615);
or U13234 (N_13234,N_12989,N_12817);
and U13235 (N_13235,N_12686,N_12773);
nand U13236 (N_13236,N_12838,N_12505);
or U13237 (N_13237,N_12753,N_12806);
or U13238 (N_13238,N_12797,N_12515);
xnor U13239 (N_13239,N_12616,N_12902);
nor U13240 (N_13240,N_12713,N_12906);
or U13241 (N_13241,N_12646,N_12699);
nand U13242 (N_13242,N_12596,N_12623);
xnor U13243 (N_13243,N_12522,N_12871);
or U13244 (N_13244,N_12540,N_12607);
xor U13245 (N_13245,N_12530,N_12601);
nand U13246 (N_13246,N_12677,N_12840);
and U13247 (N_13247,N_12799,N_12981);
nor U13248 (N_13248,N_12654,N_12672);
and U13249 (N_13249,N_12916,N_12627);
xor U13250 (N_13250,N_12841,N_12500);
or U13251 (N_13251,N_12712,N_12769);
and U13252 (N_13252,N_12804,N_12617);
nand U13253 (N_13253,N_12837,N_12562);
xnor U13254 (N_13254,N_12686,N_12835);
xor U13255 (N_13255,N_12503,N_12651);
nand U13256 (N_13256,N_12787,N_12880);
nand U13257 (N_13257,N_12877,N_12815);
nand U13258 (N_13258,N_12606,N_12729);
nand U13259 (N_13259,N_12971,N_12898);
and U13260 (N_13260,N_12636,N_12976);
and U13261 (N_13261,N_12826,N_12867);
or U13262 (N_13262,N_12763,N_12713);
xnor U13263 (N_13263,N_12680,N_12610);
nand U13264 (N_13264,N_12580,N_12731);
nand U13265 (N_13265,N_12975,N_12631);
and U13266 (N_13266,N_12858,N_12791);
nor U13267 (N_13267,N_12503,N_12558);
xor U13268 (N_13268,N_12923,N_12591);
nand U13269 (N_13269,N_12506,N_12643);
xor U13270 (N_13270,N_12528,N_12630);
and U13271 (N_13271,N_12676,N_12555);
or U13272 (N_13272,N_12607,N_12992);
or U13273 (N_13273,N_12526,N_12714);
nand U13274 (N_13274,N_12542,N_12540);
and U13275 (N_13275,N_12697,N_12581);
and U13276 (N_13276,N_12959,N_12681);
or U13277 (N_13277,N_12817,N_12778);
xnor U13278 (N_13278,N_12773,N_12872);
nand U13279 (N_13279,N_12692,N_12615);
xnor U13280 (N_13280,N_12975,N_12724);
nor U13281 (N_13281,N_12656,N_12517);
or U13282 (N_13282,N_12983,N_12638);
nand U13283 (N_13283,N_12729,N_12810);
or U13284 (N_13284,N_12938,N_12830);
and U13285 (N_13285,N_12880,N_12640);
nor U13286 (N_13286,N_12949,N_12866);
xnor U13287 (N_13287,N_12726,N_12661);
xnor U13288 (N_13288,N_12727,N_12893);
or U13289 (N_13289,N_12590,N_12644);
xnor U13290 (N_13290,N_12757,N_12982);
nand U13291 (N_13291,N_12662,N_12922);
or U13292 (N_13292,N_12998,N_12911);
nand U13293 (N_13293,N_12537,N_12517);
nor U13294 (N_13294,N_12558,N_12852);
xnor U13295 (N_13295,N_12639,N_12947);
nor U13296 (N_13296,N_12594,N_12651);
or U13297 (N_13297,N_12986,N_12869);
nor U13298 (N_13298,N_12737,N_12736);
nand U13299 (N_13299,N_12966,N_12726);
nor U13300 (N_13300,N_12618,N_12624);
or U13301 (N_13301,N_12815,N_12896);
nor U13302 (N_13302,N_12601,N_12764);
xor U13303 (N_13303,N_12563,N_12639);
xor U13304 (N_13304,N_12799,N_12989);
nor U13305 (N_13305,N_12924,N_12726);
xor U13306 (N_13306,N_12529,N_12823);
xor U13307 (N_13307,N_12857,N_12684);
nand U13308 (N_13308,N_12618,N_12860);
and U13309 (N_13309,N_12796,N_12953);
and U13310 (N_13310,N_12758,N_12950);
nor U13311 (N_13311,N_12774,N_12655);
or U13312 (N_13312,N_12666,N_12998);
and U13313 (N_13313,N_12560,N_12590);
and U13314 (N_13314,N_12835,N_12692);
and U13315 (N_13315,N_12534,N_12747);
nor U13316 (N_13316,N_12909,N_12735);
or U13317 (N_13317,N_12934,N_12801);
xor U13318 (N_13318,N_12960,N_12879);
or U13319 (N_13319,N_12959,N_12647);
nand U13320 (N_13320,N_12730,N_12715);
nor U13321 (N_13321,N_12519,N_12952);
and U13322 (N_13322,N_12621,N_12912);
xor U13323 (N_13323,N_12608,N_12906);
and U13324 (N_13324,N_12760,N_12890);
xnor U13325 (N_13325,N_12521,N_12544);
xor U13326 (N_13326,N_12898,N_12894);
nand U13327 (N_13327,N_12820,N_12578);
xor U13328 (N_13328,N_12792,N_12817);
xor U13329 (N_13329,N_12565,N_12638);
nor U13330 (N_13330,N_12956,N_12682);
or U13331 (N_13331,N_12788,N_12827);
nand U13332 (N_13332,N_12992,N_12914);
nand U13333 (N_13333,N_12517,N_12669);
xor U13334 (N_13334,N_12725,N_12572);
nand U13335 (N_13335,N_12983,N_12694);
or U13336 (N_13336,N_12534,N_12879);
nand U13337 (N_13337,N_12849,N_12852);
and U13338 (N_13338,N_12941,N_12787);
or U13339 (N_13339,N_12651,N_12720);
nand U13340 (N_13340,N_12773,N_12771);
nor U13341 (N_13341,N_12663,N_12756);
xnor U13342 (N_13342,N_12929,N_12907);
or U13343 (N_13343,N_12790,N_12518);
xor U13344 (N_13344,N_12956,N_12522);
and U13345 (N_13345,N_12834,N_12510);
nor U13346 (N_13346,N_12782,N_12621);
xor U13347 (N_13347,N_12957,N_12932);
nand U13348 (N_13348,N_12935,N_12900);
or U13349 (N_13349,N_12920,N_12514);
and U13350 (N_13350,N_12529,N_12714);
nand U13351 (N_13351,N_12917,N_12590);
or U13352 (N_13352,N_12968,N_12748);
xor U13353 (N_13353,N_12575,N_12824);
nor U13354 (N_13354,N_12591,N_12507);
and U13355 (N_13355,N_12806,N_12634);
xor U13356 (N_13356,N_12748,N_12838);
and U13357 (N_13357,N_12850,N_12729);
and U13358 (N_13358,N_12877,N_12862);
or U13359 (N_13359,N_12856,N_12836);
nand U13360 (N_13360,N_12703,N_12535);
or U13361 (N_13361,N_12903,N_12600);
xnor U13362 (N_13362,N_12940,N_12875);
xnor U13363 (N_13363,N_12565,N_12639);
or U13364 (N_13364,N_12844,N_12854);
and U13365 (N_13365,N_12578,N_12685);
xor U13366 (N_13366,N_12979,N_12737);
and U13367 (N_13367,N_12750,N_12806);
or U13368 (N_13368,N_12844,N_12950);
nand U13369 (N_13369,N_12543,N_12849);
and U13370 (N_13370,N_12751,N_12863);
nor U13371 (N_13371,N_12550,N_12978);
and U13372 (N_13372,N_12984,N_12832);
and U13373 (N_13373,N_12782,N_12745);
or U13374 (N_13374,N_12771,N_12550);
and U13375 (N_13375,N_12784,N_12686);
or U13376 (N_13376,N_12998,N_12869);
nor U13377 (N_13377,N_12689,N_12881);
xnor U13378 (N_13378,N_12761,N_12562);
or U13379 (N_13379,N_12654,N_12534);
xnor U13380 (N_13380,N_12738,N_12999);
nor U13381 (N_13381,N_12935,N_12707);
or U13382 (N_13382,N_12853,N_12899);
nand U13383 (N_13383,N_12806,N_12606);
nand U13384 (N_13384,N_12737,N_12777);
nor U13385 (N_13385,N_12834,N_12588);
and U13386 (N_13386,N_12702,N_12902);
and U13387 (N_13387,N_12520,N_12846);
nand U13388 (N_13388,N_12825,N_12865);
nand U13389 (N_13389,N_12709,N_12567);
or U13390 (N_13390,N_12522,N_12873);
or U13391 (N_13391,N_12653,N_12886);
nor U13392 (N_13392,N_12689,N_12548);
or U13393 (N_13393,N_12832,N_12978);
xor U13394 (N_13394,N_12685,N_12897);
nand U13395 (N_13395,N_12970,N_12983);
nor U13396 (N_13396,N_12736,N_12742);
and U13397 (N_13397,N_12764,N_12712);
nor U13398 (N_13398,N_12584,N_12754);
or U13399 (N_13399,N_12642,N_12775);
and U13400 (N_13400,N_12526,N_12633);
xnor U13401 (N_13401,N_12839,N_12892);
nand U13402 (N_13402,N_12500,N_12818);
nand U13403 (N_13403,N_12963,N_12783);
nor U13404 (N_13404,N_12503,N_12770);
xor U13405 (N_13405,N_12735,N_12985);
nor U13406 (N_13406,N_12535,N_12626);
or U13407 (N_13407,N_12834,N_12953);
nand U13408 (N_13408,N_12577,N_12500);
xnor U13409 (N_13409,N_12832,N_12605);
nand U13410 (N_13410,N_12692,N_12519);
xnor U13411 (N_13411,N_12532,N_12772);
and U13412 (N_13412,N_12664,N_12701);
nand U13413 (N_13413,N_12925,N_12596);
or U13414 (N_13414,N_12629,N_12850);
or U13415 (N_13415,N_12889,N_12862);
nand U13416 (N_13416,N_12683,N_12693);
nand U13417 (N_13417,N_12915,N_12846);
or U13418 (N_13418,N_12505,N_12573);
xor U13419 (N_13419,N_12952,N_12853);
and U13420 (N_13420,N_12776,N_12683);
or U13421 (N_13421,N_12675,N_12699);
nand U13422 (N_13422,N_12822,N_12914);
xor U13423 (N_13423,N_12629,N_12596);
and U13424 (N_13424,N_12649,N_12504);
and U13425 (N_13425,N_12926,N_12775);
nand U13426 (N_13426,N_12799,N_12532);
xor U13427 (N_13427,N_12851,N_12541);
xnor U13428 (N_13428,N_12627,N_12716);
nand U13429 (N_13429,N_12608,N_12916);
and U13430 (N_13430,N_12960,N_12849);
xnor U13431 (N_13431,N_12588,N_12913);
and U13432 (N_13432,N_12926,N_12996);
and U13433 (N_13433,N_12933,N_12718);
nand U13434 (N_13434,N_12558,N_12579);
and U13435 (N_13435,N_12713,N_12680);
or U13436 (N_13436,N_12648,N_12922);
nor U13437 (N_13437,N_12617,N_12589);
or U13438 (N_13438,N_12737,N_12778);
xnor U13439 (N_13439,N_12794,N_12502);
nor U13440 (N_13440,N_12739,N_12726);
xor U13441 (N_13441,N_12980,N_12867);
nand U13442 (N_13442,N_12543,N_12672);
nor U13443 (N_13443,N_12671,N_12682);
or U13444 (N_13444,N_12865,N_12856);
and U13445 (N_13445,N_12502,N_12526);
and U13446 (N_13446,N_12661,N_12610);
nor U13447 (N_13447,N_12864,N_12704);
or U13448 (N_13448,N_12504,N_12617);
nor U13449 (N_13449,N_12679,N_12894);
nand U13450 (N_13450,N_12662,N_12984);
nor U13451 (N_13451,N_12526,N_12646);
nor U13452 (N_13452,N_12767,N_12819);
or U13453 (N_13453,N_12666,N_12553);
xnor U13454 (N_13454,N_12980,N_12582);
nor U13455 (N_13455,N_12953,N_12867);
and U13456 (N_13456,N_12969,N_12615);
nor U13457 (N_13457,N_12830,N_12581);
xnor U13458 (N_13458,N_12627,N_12994);
nor U13459 (N_13459,N_12692,N_12949);
xnor U13460 (N_13460,N_12701,N_12757);
xnor U13461 (N_13461,N_12573,N_12809);
nand U13462 (N_13462,N_12589,N_12844);
xor U13463 (N_13463,N_12781,N_12517);
nand U13464 (N_13464,N_12744,N_12725);
nand U13465 (N_13465,N_12889,N_12664);
nand U13466 (N_13466,N_12613,N_12718);
and U13467 (N_13467,N_12713,N_12972);
and U13468 (N_13468,N_12778,N_12544);
xor U13469 (N_13469,N_12845,N_12746);
or U13470 (N_13470,N_12703,N_12744);
and U13471 (N_13471,N_12602,N_12815);
nand U13472 (N_13472,N_12619,N_12730);
nand U13473 (N_13473,N_12766,N_12969);
and U13474 (N_13474,N_12796,N_12532);
nand U13475 (N_13475,N_12762,N_12740);
nor U13476 (N_13476,N_12745,N_12646);
and U13477 (N_13477,N_12871,N_12571);
xnor U13478 (N_13478,N_12735,N_12938);
nor U13479 (N_13479,N_12579,N_12929);
or U13480 (N_13480,N_12823,N_12961);
xor U13481 (N_13481,N_12566,N_12725);
or U13482 (N_13482,N_12737,N_12983);
and U13483 (N_13483,N_12963,N_12604);
and U13484 (N_13484,N_12861,N_12631);
nor U13485 (N_13485,N_12550,N_12925);
xnor U13486 (N_13486,N_12960,N_12950);
and U13487 (N_13487,N_12987,N_12678);
nand U13488 (N_13488,N_12755,N_12941);
nor U13489 (N_13489,N_12560,N_12669);
nand U13490 (N_13490,N_12843,N_12992);
or U13491 (N_13491,N_12987,N_12524);
and U13492 (N_13492,N_12833,N_12984);
xnor U13493 (N_13493,N_12932,N_12952);
xor U13494 (N_13494,N_12895,N_12855);
and U13495 (N_13495,N_12750,N_12584);
or U13496 (N_13496,N_12758,N_12839);
xor U13497 (N_13497,N_12672,N_12697);
nor U13498 (N_13498,N_12731,N_12670);
or U13499 (N_13499,N_12766,N_12851);
nor U13500 (N_13500,N_13096,N_13264);
and U13501 (N_13501,N_13399,N_13404);
nor U13502 (N_13502,N_13110,N_13260);
xor U13503 (N_13503,N_13358,N_13158);
and U13504 (N_13504,N_13302,N_13215);
nor U13505 (N_13505,N_13006,N_13197);
xor U13506 (N_13506,N_13168,N_13130);
or U13507 (N_13507,N_13427,N_13193);
nand U13508 (N_13508,N_13083,N_13199);
nor U13509 (N_13509,N_13224,N_13471);
nor U13510 (N_13510,N_13415,N_13336);
nand U13511 (N_13511,N_13346,N_13277);
or U13512 (N_13512,N_13405,N_13155);
nor U13513 (N_13513,N_13079,N_13126);
and U13514 (N_13514,N_13340,N_13452);
nor U13515 (N_13515,N_13437,N_13312);
xnor U13516 (N_13516,N_13383,N_13227);
nand U13517 (N_13517,N_13107,N_13357);
xnor U13518 (N_13518,N_13234,N_13065);
xnor U13519 (N_13519,N_13271,N_13254);
and U13520 (N_13520,N_13183,N_13046);
xor U13521 (N_13521,N_13474,N_13174);
nor U13522 (N_13522,N_13294,N_13338);
and U13523 (N_13523,N_13318,N_13253);
xor U13524 (N_13524,N_13024,N_13327);
nand U13525 (N_13525,N_13282,N_13274);
xor U13526 (N_13526,N_13162,N_13468);
xnor U13527 (N_13527,N_13036,N_13093);
or U13528 (N_13528,N_13388,N_13186);
and U13529 (N_13529,N_13394,N_13479);
nand U13530 (N_13530,N_13444,N_13090);
or U13531 (N_13531,N_13418,N_13494);
and U13532 (N_13532,N_13379,N_13409);
xor U13533 (N_13533,N_13495,N_13167);
nor U13534 (N_13534,N_13116,N_13015);
or U13535 (N_13535,N_13011,N_13221);
xnor U13536 (N_13536,N_13456,N_13066);
and U13537 (N_13537,N_13101,N_13176);
nand U13538 (N_13538,N_13434,N_13124);
and U13539 (N_13539,N_13021,N_13099);
and U13540 (N_13540,N_13283,N_13304);
or U13541 (N_13541,N_13053,N_13122);
nor U13542 (N_13542,N_13117,N_13425);
nor U13543 (N_13543,N_13332,N_13345);
and U13544 (N_13544,N_13477,N_13407);
xnor U13545 (N_13545,N_13300,N_13320);
nor U13546 (N_13546,N_13134,N_13056);
or U13547 (N_13547,N_13104,N_13014);
and U13548 (N_13548,N_13373,N_13401);
and U13549 (N_13549,N_13200,N_13400);
and U13550 (N_13550,N_13424,N_13050);
nand U13551 (N_13551,N_13291,N_13261);
and U13552 (N_13552,N_13348,N_13395);
xnor U13553 (N_13553,N_13089,N_13371);
nor U13554 (N_13554,N_13272,N_13125);
xor U13555 (N_13555,N_13423,N_13275);
xor U13556 (N_13556,N_13005,N_13040);
and U13557 (N_13557,N_13390,N_13019);
nor U13558 (N_13558,N_13301,N_13218);
xor U13559 (N_13559,N_13372,N_13329);
or U13560 (N_13560,N_13073,N_13003);
and U13561 (N_13561,N_13041,N_13240);
or U13562 (N_13562,N_13440,N_13088);
or U13563 (N_13563,N_13285,N_13097);
xor U13564 (N_13564,N_13105,N_13368);
nand U13565 (N_13565,N_13069,N_13182);
nand U13566 (N_13566,N_13378,N_13054);
nor U13567 (N_13567,N_13127,N_13025);
xnor U13568 (N_13568,N_13386,N_13201);
and U13569 (N_13569,N_13194,N_13326);
or U13570 (N_13570,N_13287,N_13236);
and U13571 (N_13571,N_13463,N_13075);
and U13572 (N_13572,N_13493,N_13012);
or U13573 (N_13573,N_13419,N_13141);
xor U13574 (N_13574,N_13316,N_13289);
and U13575 (N_13575,N_13026,N_13109);
and U13576 (N_13576,N_13487,N_13288);
nor U13577 (N_13577,N_13462,N_13255);
nand U13578 (N_13578,N_13132,N_13049);
and U13579 (N_13579,N_13363,N_13350);
nor U13580 (N_13580,N_13068,N_13273);
xor U13581 (N_13581,N_13061,N_13481);
nand U13582 (N_13582,N_13233,N_13016);
xnor U13583 (N_13583,N_13185,N_13108);
nand U13584 (N_13584,N_13499,N_13343);
or U13585 (N_13585,N_13210,N_13416);
and U13586 (N_13586,N_13489,N_13439);
xnor U13587 (N_13587,N_13145,N_13370);
nand U13588 (N_13588,N_13428,N_13038);
nand U13589 (N_13589,N_13391,N_13147);
and U13590 (N_13590,N_13223,N_13196);
and U13591 (N_13591,N_13173,N_13103);
or U13592 (N_13592,N_13458,N_13131);
and U13593 (N_13593,N_13151,N_13453);
nand U13594 (N_13594,N_13118,N_13002);
nor U13595 (N_13595,N_13295,N_13460);
xor U13596 (N_13596,N_13498,N_13094);
and U13597 (N_13597,N_13192,N_13031);
nor U13598 (N_13598,N_13010,N_13359);
and U13599 (N_13599,N_13270,N_13319);
nor U13600 (N_13600,N_13208,N_13483);
and U13601 (N_13601,N_13365,N_13081);
nor U13602 (N_13602,N_13137,N_13204);
xor U13603 (N_13603,N_13202,N_13485);
nor U13604 (N_13604,N_13252,N_13190);
xnor U13605 (N_13605,N_13374,N_13263);
or U13606 (N_13606,N_13058,N_13142);
nor U13607 (N_13607,N_13175,N_13461);
and U13608 (N_13608,N_13445,N_13450);
or U13609 (N_13609,N_13059,N_13308);
and U13610 (N_13610,N_13091,N_13375);
nor U13611 (N_13611,N_13044,N_13212);
xnor U13612 (N_13612,N_13143,N_13140);
and U13613 (N_13613,N_13403,N_13051);
nand U13614 (N_13614,N_13331,N_13412);
nand U13615 (N_13615,N_13009,N_13228);
nand U13616 (N_13616,N_13478,N_13426);
nand U13617 (N_13617,N_13177,N_13298);
or U13618 (N_13618,N_13045,N_13238);
or U13619 (N_13619,N_13465,N_13259);
or U13620 (N_13620,N_13153,N_13303);
and U13621 (N_13621,N_13013,N_13203);
and U13622 (N_13622,N_13070,N_13353);
nand U13623 (N_13623,N_13451,N_13286);
and U13624 (N_13624,N_13347,N_13023);
xnor U13625 (N_13625,N_13420,N_13156);
and U13626 (N_13626,N_13048,N_13382);
nand U13627 (N_13627,N_13361,N_13213);
nor U13628 (N_13628,N_13310,N_13402);
or U13629 (N_13629,N_13328,N_13008);
or U13630 (N_13630,N_13028,N_13446);
or U13631 (N_13631,N_13047,N_13480);
nand U13632 (N_13632,N_13442,N_13082);
xnor U13633 (N_13633,N_13064,N_13406);
or U13634 (N_13634,N_13466,N_13018);
or U13635 (N_13635,N_13095,N_13473);
nand U13636 (N_13636,N_13146,N_13242);
xor U13637 (N_13637,N_13100,N_13389);
or U13638 (N_13638,N_13413,N_13317);
nor U13639 (N_13639,N_13396,N_13102);
and U13640 (N_13640,N_13311,N_13219);
nor U13641 (N_13641,N_13237,N_13033);
nor U13642 (N_13642,N_13341,N_13339);
or U13643 (N_13643,N_13266,N_13032);
and U13644 (N_13644,N_13376,N_13217);
and U13645 (N_13645,N_13188,N_13290);
or U13646 (N_13646,N_13251,N_13349);
or U13647 (N_13647,N_13246,N_13464);
or U13648 (N_13648,N_13454,N_13144);
nand U13649 (N_13649,N_13037,N_13457);
nand U13650 (N_13650,N_13092,N_13292);
nor U13651 (N_13651,N_13136,N_13245);
or U13652 (N_13652,N_13157,N_13152);
nand U13653 (N_13653,N_13247,N_13179);
nor U13654 (N_13654,N_13472,N_13355);
xnor U13655 (N_13655,N_13241,N_13080);
and U13656 (N_13656,N_13232,N_13313);
nor U13657 (N_13657,N_13414,N_13138);
nor U13658 (N_13658,N_13377,N_13169);
xnor U13659 (N_13659,N_13225,N_13393);
nor U13660 (N_13660,N_13262,N_13170);
and U13661 (N_13661,N_13189,N_13397);
nand U13662 (N_13662,N_13482,N_13344);
nor U13663 (N_13663,N_13380,N_13307);
nand U13664 (N_13664,N_13447,N_13408);
xor U13665 (N_13665,N_13384,N_13244);
and U13666 (N_13666,N_13432,N_13239);
nand U13667 (N_13667,N_13085,N_13161);
and U13668 (N_13668,N_13211,N_13330);
nand U13669 (N_13669,N_13488,N_13306);
or U13670 (N_13670,N_13035,N_13430);
and U13671 (N_13671,N_13150,N_13367);
nand U13672 (N_13672,N_13258,N_13475);
and U13673 (N_13673,N_13029,N_13476);
nand U13674 (N_13674,N_13159,N_13184);
or U13675 (N_13675,N_13323,N_13265);
nand U13676 (N_13676,N_13165,N_13305);
nor U13677 (N_13677,N_13062,N_13268);
nor U13678 (N_13678,N_13497,N_13180);
or U13679 (N_13679,N_13207,N_13063);
and U13680 (N_13680,N_13269,N_13490);
xor U13681 (N_13681,N_13352,N_13387);
nand U13682 (N_13682,N_13071,N_13337);
nor U13683 (N_13683,N_13148,N_13076);
nand U13684 (N_13684,N_13334,N_13030);
nor U13685 (N_13685,N_13429,N_13496);
and U13686 (N_13686,N_13164,N_13216);
nand U13687 (N_13687,N_13448,N_13299);
xor U13688 (N_13688,N_13280,N_13243);
and U13689 (N_13689,N_13369,N_13149);
or U13690 (N_13690,N_13250,N_13276);
nand U13691 (N_13691,N_13057,N_13314);
and U13692 (N_13692,N_13086,N_13354);
or U13693 (N_13693,N_13226,N_13017);
nor U13694 (N_13694,N_13467,N_13004);
and U13695 (N_13695,N_13325,N_13360);
xnor U13696 (N_13696,N_13135,N_13139);
nand U13697 (N_13697,N_13333,N_13106);
or U13698 (N_13698,N_13043,N_13385);
nand U13699 (N_13699,N_13441,N_13195);
xor U13700 (N_13700,N_13364,N_13222);
or U13701 (N_13701,N_13322,N_13257);
or U13702 (N_13702,N_13181,N_13392);
or U13703 (N_13703,N_13335,N_13133);
nand U13704 (N_13704,N_13455,N_13160);
and U13705 (N_13705,N_13220,N_13027);
nand U13706 (N_13706,N_13410,N_13074);
xnor U13707 (N_13707,N_13055,N_13205);
nor U13708 (N_13708,N_13324,N_13438);
nor U13709 (N_13709,N_13492,N_13214);
xnor U13710 (N_13710,N_13112,N_13128);
or U13711 (N_13711,N_13039,N_13171);
nor U13712 (N_13712,N_13278,N_13443);
nor U13713 (N_13713,N_13431,N_13491);
and U13714 (N_13714,N_13209,N_13235);
and U13715 (N_13715,N_13435,N_13230);
and U13716 (N_13716,N_13470,N_13114);
nor U13717 (N_13717,N_13020,N_13293);
and U13718 (N_13718,N_13007,N_13000);
nor U13719 (N_13719,N_13297,N_13469);
nand U13720 (N_13720,N_13119,N_13433);
and U13721 (N_13721,N_13087,N_13198);
xor U13722 (N_13722,N_13123,N_13256);
or U13723 (N_13723,N_13052,N_13022);
and U13724 (N_13724,N_13284,N_13484);
nand U13725 (N_13725,N_13206,N_13411);
nor U13726 (N_13726,N_13060,N_13486);
xor U13727 (N_13727,N_13321,N_13078);
xor U13728 (N_13728,N_13267,N_13084);
xnor U13729 (N_13729,N_13309,N_13417);
nand U13730 (N_13730,N_13229,N_13067);
nor U13731 (N_13731,N_13342,N_13249);
xor U13732 (N_13732,N_13042,N_13398);
nor U13733 (N_13733,N_13166,N_13356);
xnor U13734 (N_13734,N_13449,N_13001);
or U13735 (N_13735,N_13163,N_13072);
nor U13736 (N_13736,N_13421,N_13191);
nand U13737 (N_13737,N_13281,N_13121);
nor U13738 (N_13738,N_13366,N_13120);
nand U13739 (N_13739,N_13178,N_13154);
or U13740 (N_13740,N_13113,N_13111);
and U13741 (N_13741,N_13296,N_13248);
nor U13742 (N_13742,N_13115,N_13034);
xnor U13743 (N_13743,N_13172,N_13362);
nor U13744 (N_13744,N_13436,N_13381);
xnor U13745 (N_13745,N_13187,N_13098);
nand U13746 (N_13746,N_13315,N_13231);
nand U13747 (N_13747,N_13077,N_13129);
and U13748 (N_13748,N_13279,N_13459);
nor U13749 (N_13749,N_13422,N_13351);
nor U13750 (N_13750,N_13412,N_13438);
xor U13751 (N_13751,N_13254,N_13491);
nand U13752 (N_13752,N_13092,N_13021);
xnor U13753 (N_13753,N_13183,N_13093);
or U13754 (N_13754,N_13137,N_13488);
xnor U13755 (N_13755,N_13458,N_13495);
and U13756 (N_13756,N_13255,N_13066);
xnor U13757 (N_13757,N_13352,N_13122);
xor U13758 (N_13758,N_13063,N_13261);
and U13759 (N_13759,N_13204,N_13064);
and U13760 (N_13760,N_13172,N_13063);
xor U13761 (N_13761,N_13314,N_13316);
and U13762 (N_13762,N_13130,N_13145);
nand U13763 (N_13763,N_13331,N_13039);
and U13764 (N_13764,N_13279,N_13053);
nor U13765 (N_13765,N_13427,N_13498);
or U13766 (N_13766,N_13232,N_13298);
and U13767 (N_13767,N_13118,N_13346);
or U13768 (N_13768,N_13476,N_13147);
nand U13769 (N_13769,N_13353,N_13419);
nand U13770 (N_13770,N_13254,N_13138);
or U13771 (N_13771,N_13416,N_13026);
nor U13772 (N_13772,N_13131,N_13238);
or U13773 (N_13773,N_13244,N_13122);
nor U13774 (N_13774,N_13143,N_13438);
nand U13775 (N_13775,N_13279,N_13060);
nor U13776 (N_13776,N_13292,N_13391);
nor U13777 (N_13777,N_13195,N_13034);
or U13778 (N_13778,N_13110,N_13230);
xor U13779 (N_13779,N_13011,N_13441);
nor U13780 (N_13780,N_13205,N_13422);
nand U13781 (N_13781,N_13392,N_13481);
nand U13782 (N_13782,N_13243,N_13228);
or U13783 (N_13783,N_13287,N_13299);
nand U13784 (N_13784,N_13435,N_13109);
nor U13785 (N_13785,N_13133,N_13001);
or U13786 (N_13786,N_13487,N_13254);
nand U13787 (N_13787,N_13140,N_13261);
xnor U13788 (N_13788,N_13144,N_13112);
or U13789 (N_13789,N_13101,N_13389);
and U13790 (N_13790,N_13040,N_13172);
or U13791 (N_13791,N_13086,N_13387);
or U13792 (N_13792,N_13357,N_13493);
xor U13793 (N_13793,N_13320,N_13087);
and U13794 (N_13794,N_13262,N_13461);
or U13795 (N_13795,N_13235,N_13060);
or U13796 (N_13796,N_13466,N_13399);
nor U13797 (N_13797,N_13095,N_13189);
and U13798 (N_13798,N_13042,N_13393);
and U13799 (N_13799,N_13470,N_13360);
nor U13800 (N_13800,N_13194,N_13193);
nor U13801 (N_13801,N_13174,N_13048);
nand U13802 (N_13802,N_13415,N_13189);
and U13803 (N_13803,N_13462,N_13382);
nand U13804 (N_13804,N_13334,N_13462);
and U13805 (N_13805,N_13131,N_13270);
nor U13806 (N_13806,N_13103,N_13489);
xor U13807 (N_13807,N_13139,N_13469);
or U13808 (N_13808,N_13128,N_13167);
and U13809 (N_13809,N_13430,N_13191);
or U13810 (N_13810,N_13480,N_13407);
and U13811 (N_13811,N_13233,N_13385);
nand U13812 (N_13812,N_13288,N_13422);
or U13813 (N_13813,N_13374,N_13251);
or U13814 (N_13814,N_13449,N_13421);
nand U13815 (N_13815,N_13423,N_13276);
or U13816 (N_13816,N_13102,N_13457);
xnor U13817 (N_13817,N_13448,N_13159);
and U13818 (N_13818,N_13226,N_13061);
and U13819 (N_13819,N_13455,N_13310);
and U13820 (N_13820,N_13307,N_13433);
and U13821 (N_13821,N_13323,N_13154);
and U13822 (N_13822,N_13470,N_13434);
xnor U13823 (N_13823,N_13293,N_13488);
and U13824 (N_13824,N_13222,N_13153);
and U13825 (N_13825,N_13139,N_13310);
nand U13826 (N_13826,N_13308,N_13325);
nand U13827 (N_13827,N_13404,N_13469);
or U13828 (N_13828,N_13081,N_13065);
nor U13829 (N_13829,N_13096,N_13320);
xnor U13830 (N_13830,N_13127,N_13402);
and U13831 (N_13831,N_13016,N_13139);
nor U13832 (N_13832,N_13114,N_13460);
nor U13833 (N_13833,N_13078,N_13178);
or U13834 (N_13834,N_13059,N_13198);
and U13835 (N_13835,N_13231,N_13459);
nand U13836 (N_13836,N_13021,N_13225);
nor U13837 (N_13837,N_13191,N_13014);
nand U13838 (N_13838,N_13403,N_13173);
and U13839 (N_13839,N_13245,N_13242);
nor U13840 (N_13840,N_13364,N_13249);
or U13841 (N_13841,N_13457,N_13035);
nand U13842 (N_13842,N_13160,N_13161);
nor U13843 (N_13843,N_13040,N_13340);
nand U13844 (N_13844,N_13028,N_13406);
and U13845 (N_13845,N_13426,N_13174);
or U13846 (N_13846,N_13207,N_13472);
or U13847 (N_13847,N_13144,N_13047);
nand U13848 (N_13848,N_13423,N_13368);
nand U13849 (N_13849,N_13316,N_13220);
xor U13850 (N_13850,N_13324,N_13165);
nor U13851 (N_13851,N_13472,N_13129);
xnor U13852 (N_13852,N_13126,N_13037);
or U13853 (N_13853,N_13197,N_13428);
nor U13854 (N_13854,N_13451,N_13257);
nor U13855 (N_13855,N_13087,N_13243);
nor U13856 (N_13856,N_13048,N_13074);
xnor U13857 (N_13857,N_13231,N_13107);
and U13858 (N_13858,N_13246,N_13232);
xnor U13859 (N_13859,N_13488,N_13366);
xor U13860 (N_13860,N_13220,N_13307);
nand U13861 (N_13861,N_13017,N_13326);
xnor U13862 (N_13862,N_13475,N_13045);
or U13863 (N_13863,N_13173,N_13227);
nand U13864 (N_13864,N_13435,N_13267);
nand U13865 (N_13865,N_13137,N_13431);
nand U13866 (N_13866,N_13122,N_13435);
and U13867 (N_13867,N_13169,N_13120);
nand U13868 (N_13868,N_13318,N_13219);
xnor U13869 (N_13869,N_13471,N_13210);
nand U13870 (N_13870,N_13090,N_13003);
or U13871 (N_13871,N_13400,N_13294);
or U13872 (N_13872,N_13327,N_13190);
nor U13873 (N_13873,N_13212,N_13230);
xor U13874 (N_13874,N_13349,N_13047);
nor U13875 (N_13875,N_13239,N_13431);
nor U13876 (N_13876,N_13147,N_13370);
nand U13877 (N_13877,N_13352,N_13043);
or U13878 (N_13878,N_13142,N_13010);
nand U13879 (N_13879,N_13424,N_13296);
or U13880 (N_13880,N_13308,N_13476);
nand U13881 (N_13881,N_13258,N_13329);
and U13882 (N_13882,N_13440,N_13171);
nand U13883 (N_13883,N_13058,N_13458);
nor U13884 (N_13884,N_13264,N_13260);
xnor U13885 (N_13885,N_13340,N_13466);
and U13886 (N_13886,N_13200,N_13458);
nand U13887 (N_13887,N_13173,N_13410);
and U13888 (N_13888,N_13025,N_13257);
nor U13889 (N_13889,N_13396,N_13132);
nand U13890 (N_13890,N_13178,N_13269);
nand U13891 (N_13891,N_13215,N_13121);
nand U13892 (N_13892,N_13310,N_13132);
and U13893 (N_13893,N_13175,N_13222);
nand U13894 (N_13894,N_13126,N_13370);
and U13895 (N_13895,N_13039,N_13257);
and U13896 (N_13896,N_13011,N_13451);
nor U13897 (N_13897,N_13349,N_13168);
or U13898 (N_13898,N_13172,N_13038);
xnor U13899 (N_13899,N_13096,N_13180);
or U13900 (N_13900,N_13393,N_13163);
nor U13901 (N_13901,N_13345,N_13280);
nor U13902 (N_13902,N_13005,N_13403);
nor U13903 (N_13903,N_13427,N_13351);
nand U13904 (N_13904,N_13275,N_13366);
nand U13905 (N_13905,N_13229,N_13006);
xor U13906 (N_13906,N_13004,N_13334);
or U13907 (N_13907,N_13012,N_13127);
and U13908 (N_13908,N_13483,N_13060);
nand U13909 (N_13909,N_13068,N_13391);
xnor U13910 (N_13910,N_13270,N_13019);
or U13911 (N_13911,N_13130,N_13142);
or U13912 (N_13912,N_13422,N_13349);
nand U13913 (N_13913,N_13119,N_13442);
nand U13914 (N_13914,N_13433,N_13356);
nand U13915 (N_13915,N_13178,N_13122);
nor U13916 (N_13916,N_13028,N_13357);
nor U13917 (N_13917,N_13304,N_13495);
nor U13918 (N_13918,N_13364,N_13097);
and U13919 (N_13919,N_13102,N_13137);
nor U13920 (N_13920,N_13096,N_13275);
nor U13921 (N_13921,N_13244,N_13104);
nor U13922 (N_13922,N_13164,N_13217);
xor U13923 (N_13923,N_13200,N_13218);
or U13924 (N_13924,N_13240,N_13070);
or U13925 (N_13925,N_13334,N_13101);
xnor U13926 (N_13926,N_13069,N_13305);
xor U13927 (N_13927,N_13371,N_13343);
or U13928 (N_13928,N_13318,N_13167);
and U13929 (N_13929,N_13151,N_13310);
nand U13930 (N_13930,N_13000,N_13099);
nand U13931 (N_13931,N_13076,N_13122);
nor U13932 (N_13932,N_13068,N_13213);
nor U13933 (N_13933,N_13326,N_13395);
and U13934 (N_13934,N_13035,N_13412);
or U13935 (N_13935,N_13245,N_13209);
nor U13936 (N_13936,N_13385,N_13088);
and U13937 (N_13937,N_13059,N_13102);
xnor U13938 (N_13938,N_13136,N_13266);
nor U13939 (N_13939,N_13180,N_13487);
or U13940 (N_13940,N_13265,N_13234);
and U13941 (N_13941,N_13447,N_13307);
nor U13942 (N_13942,N_13376,N_13318);
nand U13943 (N_13943,N_13269,N_13121);
nor U13944 (N_13944,N_13286,N_13456);
and U13945 (N_13945,N_13367,N_13000);
and U13946 (N_13946,N_13266,N_13084);
nor U13947 (N_13947,N_13079,N_13065);
nand U13948 (N_13948,N_13199,N_13063);
or U13949 (N_13949,N_13227,N_13338);
nand U13950 (N_13950,N_13192,N_13369);
nand U13951 (N_13951,N_13362,N_13049);
or U13952 (N_13952,N_13137,N_13268);
or U13953 (N_13953,N_13211,N_13386);
xnor U13954 (N_13954,N_13131,N_13229);
or U13955 (N_13955,N_13364,N_13192);
nor U13956 (N_13956,N_13199,N_13197);
nand U13957 (N_13957,N_13388,N_13098);
and U13958 (N_13958,N_13413,N_13429);
and U13959 (N_13959,N_13106,N_13360);
nor U13960 (N_13960,N_13131,N_13269);
nor U13961 (N_13961,N_13342,N_13432);
nor U13962 (N_13962,N_13193,N_13457);
nor U13963 (N_13963,N_13269,N_13158);
and U13964 (N_13964,N_13336,N_13107);
nand U13965 (N_13965,N_13312,N_13109);
and U13966 (N_13966,N_13023,N_13110);
xnor U13967 (N_13967,N_13101,N_13280);
or U13968 (N_13968,N_13175,N_13347);
or U13969 (N_13969,N_13300,N_13228);
or U13970 (N_13970,N_13184,N_13210);
xor U13971 (N_13971,N_13387,N_13497);
nand U13972 (N_13972,N_13180,N_13319);
nand U13973 (N_13973,N_13281,N_13440);
or U13974 (N_13974,N_13069,N_13196);
or U13975 (N_13975,N_13189,N_13492);
or U13976 (N_13976,N_13076,N_13010);
or U13977 (N_13977,N_13239,N_13471);
and U13978 (N_13978,N_13185,N_13013);
xnor U13979 (N_13979,N_13382,N_13099);
or U13980 (N_13980,N_13497,N_13411);
xnor U13981 (N_13981,N_13113,N_13398);
nand U13982 (N_13982,N_13487,N_13223);
or U13983 (N_13983,N_13230,N_13114);
xnor U13984 (N_13984,N_13080,N_13274);
xnor U13985 (N_13985,N_13012,N_13044);
nor U13986 (N_13986,N_13289,N_13066);
xor U13987 (N_13987,N_13135,N_13398);
and U13988 (N_13988,N_13062,N_13192);
xnor U13989 (N_13989,N_13172,N_13016);
nand U13990 (N_13990,N_13468,N_13202);
or U13991 (N_13991,N_13169,N_13108);
and U13992 (N_13992,N_13008,N_13396);
nand U13993 (N_13993,N_13220,N_13036);
nand U13994 (N_13994,N_13110,N_13024);
nor U13995 (N_13995,N_13458,N_13232);
nor U13996 (N_13996,N_13297,N_13206);
nand U13997 (N_13997,N_13308,N_13343);
xnor U13998 (N_13998,N_13329,N_13138);
and U13999 (N_13999,N_13031,N_13100);
and U14000 (N_14000,N_13722,N_13715);
nor U14001 (N_14001,N_13746,N_13896);
xor U14002 (N_14002,N_13576,N_13712);
nor U14003 (N_14003,N_13514,N_13950);
xnor U14004 (N_14004,N_13974,N_13721);
nand U14005 (N_14005,N_13582,N_13506);
or U14006 (N_14006,N_13937,N_13566);
xnor U14007 (N_14007,N_13917,N_13604);
and U14008 (N_14008,N_13623,N_13588);
and U14009 (N_14009,N_13541,N_13994);
or U14010 (N_14010,N_13959,N_13631);
and U14011 (N_14011,N_13632,N_13798);
or U14012 (N_14012,N_13502,N_13810);
or U14013 (N_14013,N_13790,N_13861);
nand U14014 (N_14014,N_13530,N_13688);
nand U14015 (N_14015,N_13880,N_13649);
and U14016 (N_14016,N_13613,N_13955);
and U14017 (N_14017,N_13516,N_13823);
and U14018 (N_14018,N_13922,N_13628);
or U14019 (N_14019,N_13510,N_13953);
nand U14020 (N_14020,N_13513,N_13816);
and U14021 (N_14021,N_13923,N_13667);
xor U14022 (N_14022,N_13946,N_13756);
xnor U14023 (N_14023,N_13822,N_13949);
nand U14024 (N_14024,N_13711,N_13504);
nand U14025 (N_14025,N_13802,N_13735);
or U14026 (N_14026,N_13903,N_13993);
xnor U14027 (N_14027,N_13617,N_13651);
and U14028 (N_14028,N_13501,N_13720);
and U14029 (N_14029,N_13945,N_13518);
xnor U14030 (N_14030,N_13723,N_13719);
and U14031 (N_14031,N_13612,N_13886);
xnor U14032 (N_14032,N_13505,N_13771);
nand U14033 (N_14033,N_13834,N_13879);
and U14034 (N_14034,N_13882,N_13671);
xnor U14035 (N_14035,N_13813,N_13767);
nand U14036 (N_14036,N_13564,N_13643);
and U14037 (N_14037,N_13654,N_13806);
and U14038 (N_14038,N_13619,N_13768);
nor U14039 (N_14039,N_13796,N_13567);
and U14040 (N_14040,N_13833,N_13738);
and U14041 (N_14041,N_13681,N_13553);
and U14042 (N_14042,N_13672,N_13557);
xnor U14043 (N_14043,N_13965,N_13826);
nand U14044 (N_14044,N_13935,N_13578);
or U14045 (N_14045,N_13842,N_13921);
or U14046 (N_14046,N_13990,N_13758);
or U14047 (N_14047,N_13988,N_13661);
nand U14048 (N_14048,N_13542,N_13512);
and U14049 (N_14049,N_13890,N_13815);
nand U14050 (N_14050,N_13701,N_13753);
xor U14051 (N_14051,N_13547,N_13799);
nor U14052 (N_14052,N_13726,N_13770);
and U14053 (N_14053,N_13583,N_13962);
xnor U14054 (N_14054,N_13774,N_13634);
or U14055 (N_14055,N_13591,N_13640);
nand U14056 (N_14056,N_13734,N_13779);
or U14057 (N_14057,N_13677,N_13876);
and U14058 (N_14058,N_13836,N_13772);
and U14059 (N_14059,N_13916,N_13893);
and U14060 (N_14060,N_13718,N_13811);
or U14061 (N_14061,N_13626,N_13532);
nor U14062 (N_14062,N_13891,N_13705);
nand U14063 (N_14063,N_13989,N_13752);
nor U14064 (N_14064,N_13691,N_13874);
nor U14065 (N_14065,N_13603,N_13878);
xnor U14066 (N_14066,N_13618,N_13936);
nand U14067 (N_14067,N_13702,N_13663);
and U14068 (N_14068,N_13630,N_13957);
nand U14069 (N_14069,N_13572,N_13706);
or U14070 (N_14070,N_13650,N_13938);
or U14071 (N_14071,N_13870,N_13868);
xnor U14072 (N_14072,N_13956,N_13728);
or U14073 (N_14073,N_13717,N_13764);
xnor U14074 (N_14074,N_13739,N_13551);
and U14075 (N_14075,N_13637,N_13847);
nor U14076 (N_14076,N_13692,N_13855);
and U14077 (N_14077,N_13508,N_13844);
and U14078 (N_14078,N_13670,N_13927);
nor U14079 (N_14079,N_13827,N_13967);
and U14080 (N_14080,N_13975,N_13549);
nand U14081 (N_14081,N_13933,N_13581);
and U14082 (N_14082,N_13625,N_13821);
and U14083 (N_14083,N_13812,N_13574);
nand U14084 (N_14084,N_13761,N_13570);
or U14085 (N_14085,N_13795,N_13697);
xnor U14086 (N_14086,N_13981,N_13809);
nor U14087 (N_14087,N_13608,N_13787);
nor U14088 (N_14088,N_13976,N_13596);
and U14089 (N_14089,N_13524,N_13569);
xnor U14090 (N_14090,N_13624,N_13777);
nor U14091 (N_14091,N_13716,N_13900);
and U14092 (N_14092,N_13980,N_13869);
or U14093 (N_14093,N_13710,N_13776);
and U14094 (N_14094,N_13559,N_13881);
nand U14095 (N_14095,N_13912,N_13820);
nor U14096 (N_14096,N_13932,N_13808);
and U14097 (N_14097,N_13794,N_13598);
and U14098 (N_14098,N_13839,N_13859);
or U14099 (N_14099,N_13966,N_13843);
and U14100 (N_14100,N_13611,N_13755);
nand U14101 (N_14101,N_13775,N_13732);
nand U14102 (N_14102,N_13902,N_13620);
nor U14103 (N_14103,N_13856,N_13646);
xnor U14104 (N_14104,N_13904,N_13676);
nand U14105 (N_14105,N_13866,N_13920);
xor U14106 (N_14106,N_13595,N_13780);
or U14107 (N_14107,N_13848,N_13985);
nand U14108 (N_14108,N_13525,N_13766);
nor U14109 (N_14109,N_13942,N_13644);
nand U14110 (N_14110,N_13642,N_13838);
or U14111 (N_14111,N_13754,N_13805);
nand U14112 (N_14112,N_13519,N_13892);
xor U14113 (N_14113,N_13851,N_13875);
nor U14114 (N_14114,N_13606,N_13968);
nand U14115 (N_14115,N_13684,N_13995);
nand U14116 (N_14116,N_13500,N_13763);
nor U14117 (N_14117,N_13854,N_13602);
nand U14118 (N_14118,N_13931,N_13915);
nand U14119 (N_14119,N_13698,N_13907);
or U14120 (N_14120,N_13585,N_13592);
nor U14121 (N_14121,N_13709,N_13977);
xnor U14122 (N_14122,N_13759,N_13972);
or U14123 (N_14123,N_13521,N_13694);
xnor U14124 (N_14124,N_13647,N_13944);
nor U14125 (N_14125,N_13948,N_13703);
and U14126 (N_14126,N_13546,N_13837);
nor U14127 (N_14127,N_13538,N_13607);
xor U14128 (N_14128,N_13693,N_13835);
or U14129 (N_14129,N_13616,N_13829);
nor U14130 (N_14130,N_13793,N_13889);
and U14131 (N_14131,N_13913,N_13971);
nor U14132 (N_14132,N_13939,N_13713);
xnor U14133 (N_14133,N_13653,N_13533);
nor U14134 (N_14134,N_13887,N_13695);
nand U14135 (N_14135,N_13573,N_13511);
xnor U14136 (N_14136,N_13791,N_13601);
xor U14137 (N_14137,N_13800,N_13804);
or U14138 (N_14138,N_13803,N_13509);
or U14139 (N_14139,N_13924,N_13638);
xor U14140 (N_14140,N_13888,N_13930);
nor U14141 (N_14141,N_13914,N_13778);
or U14142 (N_14142,N_13584,N_13841);
xor U14143 (N_14143,N_13529,N_13978);
or U14144 (N_14144,N_13825,N_13568);
nor U14145 (N_14145,N_13633,N_13742);
and U14146 (N_14146,N_13901,N_13765);
xor U14147 (N_14147,N_13554,N_13526);
xnor U14148 (N_14148,N_13683,N_13690);
and U14149 (N_14149,N_13655,N_13828);
nand U14150 (N_14150,N_13947,N_13750);
nor U14151 (N_14151,N_13873,N_13792);
or U14152 (N_14152,N_13961,N_13749);
xor U14153 (N_14153,N_13852,N_13964);
xor U14154 (N_14154,N_13958,N_13898);
xnor U14155 (N_14155,N_13507,N_13555);
nor U14156 (N_14156,N_13534,N_13515);
nor U14157 (N_14157,N_13575,N_13659);
or U14158 (N_14158,N_13540,N_13700);
nor U14159 (N_14159,N_13560,N_13665);
nor U14160 (N_14160,N_13982,N_13909);
or U14161 (N_14161,N_13589,N_13562);
nor U14162 (N_14162,N_13729,N_13788);
xor U14163 (N_14163,N_13737,N_13940);
nand U14164 (N_14164,N_13556,N_13819);
or U14165 (N_14165,N_13867,N_13733);
and U14166 (N_14166,N_13877,N_13668);
nor U14167 (N_14167,N_13979,N_13991);
nand U14168 (N_14168,N_13741,N_13905);
or U14169 (N_14169,N_13528,N_13605);
xor U14170 (N_14170,N_13571,N_13531);
or U14171 (N_14171,N_13831,N_13731);
nand U14172 (N_14172,N_13622,N_13801);
nand U14173 (N_14173,N_13662,N_13747);
nor U14174 (N_14174,N_13656,N_13884);
and U14175 (N_14175,N_13600,N_13593);
nand U14176 (N_14176,N_13745,N_13941);
nand U14177 (N_14177,N_13997,N_13645);
or U14178 (N_14178,N_13621,N_13535);
and U14179 (N_14179,N_13864,N_13707);
and U14180 (N_14180,N_13725,N_13925);
and U14181 (N_14181,N_13635,N_13908);
or U14182 (N_14182,N_13641,N_13951);
nand U14183 (N_14183,N_13675,N_13952);
nor U14184 (N_14184,N_13609,N_13918);
nand U14185 (N_14185,N_13579,N_13565);
or U14186 (N_14186,N_13669,N_13830);
or U14187 (N_14187,N_13523,N_13860);
nor U14188 (N_14188,N_13687,N_13679);
xnor U14189 (N_14189,N_13773,N_13615);
or U14190 (N_14190,N_13666,N_13818);
or U14191 (N_14191,N_13517,N_13730);
or U14192 (N_14192,N_13680,N_13587);
or U14193 (N_14193,N_13963,N_13863);
nand U14194 (N_14194,N_13883,N_13699);
and U14195 (N_14195,N_13545,N_13911);
nor U14196 (N_14196,N_13597,N_13561);
and U14197 (N_14197,N_13973,N_13894);
or U14198 (N_14198,N_13689,N_13599);
xor U14199 (N_14199,N_13996,N_13845);
and U14200 (N_14200,N_13849,N_13648);
and U14201 (N_14201,N_13782,N_13674);
or U14202 (N_14202,N_13897,N_13544);
or U14203 (N_14203,N_13885,N_13577);
and U14204 (N_14204,N_13899,N_13850);
nor U14205 (N_14205,N_13832,N_13895);
nor U14206 (N_14206,N_13743,N_13539);
and U14207 (N_14207,N_13906,N_13954);
or U14208 (N_14208,N_13594,N_13580);
nand U14209 (N_14209,N_13682,N_13748);
nand U14210 (N_14210,N_13708,N_13926);
nand U14211 (N_14211,N_13757,N_13871);
nand U14212 (N_14212,N_13744,N_13543);
nand U14213 (N_14213,N_13769,N_13736);
xnor U14214 (N_14214,N_13696,N_13724);
xor U14215 (N_14215,N_13807,N_13987);
or U14216 (N_14216,N_13727,N_13960);
xnor U14217 (N_14217,N_13783,N_13639);
nand U14218 (N_14218,N_13784,N_13558);
nand U14219 (N_14219,N_13527,N_13919);
or U14220 (N_14220,N_13969,N_13824);
nand U14221 (N_14221,N_13627,N_13934);
nand U14222 (N_14222,N_13928,N_13522);
or U14223 (N_14223,N_13664,N_13636);
nand U14224 (N_14224,N_13614,N_13872);
and U14225 (N_14225,N_13781,N_13610);
nand U14226 (N_14226,N_13943,N_13983);
xnor U14227 (N_14227,N_13590,N_13817);
xor U14228 (N_14228,N_13992,N_13865);
or U14229 (N_14229,N_13846,N_13840);
and U14230 (N_14230,N_13814,N_13786);
or U14231 (N_14231,N_13658,N_13537);
nand U14232 (N_14232,N_13785,N_13586);
nor U14233 (N_14233,N_13685,N_13999);
nand U14234 (N_14234,N_13714,N_13548);
or U14235 (N_14235,N_13552,N_13652);
or U14236 (N_14236,N_13673,N_13862);
and U14237 (N_14237,N_13986,N_13550);
nor U14238 (N_14238,N_13789,N_13660);
and U14239 (N_14239,N_13857,N_13760);
xor U14240 (N_14240,N_13858,N_13740);
nand U14241 (N_14241,N_13797,N_13929);
nand U14242 (N_14242,N_13853,N_13657);
nor U14243 (N_14243,N_13686,N_13910);
nor U14244 (N_14244,N_13970,N_13563);
nand U14245 (N_14245,N_13520,N_13751);
xnor U14246 (N_14246,N_13704,N_13998);
and U14247 (N_14247,N_13678,N_13629);
nor U14248 (N_14248,N_13536,N_13984);
xor U14249 (N_14249,N_13503,N_13762);
nand U14250 (N_14250,N_13825,N_13895);
and U14251 (N_14251,N_13841,N_13613);
xor U14252 (N_14252,N_13846,N_13731);
nor U14253 (N_14253,N_13989,N_13933);
or U14254 (N_14254,N_13874,N_13781);
xor U14255 (N_14255,N_13937,N_13615);
nor U14256 (N_14256,N_13726,N_13532);
nand U14257 (N_14257,N_13924,N_13561);
and U14258 (N_14258,N_13709,N_13892);
nor U14259 (N_14259,N_13598,N_13997);
nor U14260 (N_14260,N_13754,N_13968);
nand U14261 (N_14261,N_13953,N_13866);
or U14262 (N_14262,N_13555,N_13530);
or U14263 (N_14263,N_13959,N_13935);
and U14264 (N_14264,N_13672,N_13683);
and U14265 (N_14265,N_13680,N_13673);
and U14266 (N_14266,N_13922,N_13941);
nand U14267 (N_14267,N_13743,N_13753);
nand U14268 (N_14268,N_13642,N_13887);
xor U14269 (N_14269,N_13964,N_13781);
or U14270 (N_14270,N_13685,N_13865);
xor U14271 (N_14271,N_13623,N_13726);
and U14272 (N_14272,N_13511,N_13545);
and U14273 (N_14273,N_13671,N_13516);
nand U14274 (N_14274,N_13691,N_13962);
and U14275 (N_14275,N_13840,N_13753);
and U14276 (N_14276,N_13522,N_13542);
or U14277 (N_14277,N_13539,N_13681);
nor U14278 (N_14278,N_13909,N_13555);
or U14279 (N_14279,N_13537,N_13547);
xnor U14280 (N_14280,N_13989,N_13996);
and U14281 (N_14281,N_13780,N_13639);
or U14282 (N_14282,N_13719,N_13631);
nor U14283 (N_14283,N_13652,N_13986);
xnor U14284 (N_14284,N_13518,N_13632);
nand U14285 (N_14285,N_13703,N_13722);
xor U14286 (N_14286,N_13793,N_13803);
or U14287 (N_14287,N_13853,N_13910);
or U14288 (N_14288,N_13889,N_13635);
nor U14289 (N_14289,N_13775,N_13777);
xor U14290 (N_14290,N_13773,N_13863);
nand U14291 (N_14291,N_13753,N_13615);
xor U14292 (N_14292,N_13705,N_13623);
nor U14293 (N_14293,N_13989,N_13675);
xnor U14294 (N_14294,N_13533,N_13836);
xor U14295 (N_14295,N_13531,N_13691);
and U14296 (N_14296,N_13989,N_13822);
and U14297 (N_14297,N_13830,N_13731);
or U14298 (N_14298,N_13625,N_13747);
and U14299 (N_14299,N_13705,N_13711);
xor U14300 (N_14300,N_13660,N_13805);
nor U14301 (N_14301,N_13963,N_13760);
xnor U14302 (N_14302,N_13601,N_13645);
xor U14303 (N_14303,N_13893,N_13504);
and U14304 (N_14304,N_13798,N_13622);
and U14305 (N_14305,N_13519,N_13764);
or U14306 (N_14306,N_13676,N_13980);
xor U14307 (N_14307,N_13654,N_13665);
nor U14308 (N_14308,N_13999,N_13605);
nor U14309 (N_14309,N_13913,N_13625);
xor U14310 (N_14310,N_13726,N_13888);
xnor U14311 (N_14311,N_13997,N_13879);
nand U14312 (N_14312,N_13648,N_13704);
xnor U14313 (N_14313,N_13721,N_13814);
nand U14314 (N_14314,N_13767,N_13750);
nand U14315 (N_14315,N_13654,N_13614);
or U14316 (N_14316,N_13720,N_13741);
and U14317 (N_14317,N_13548,N_13882);
and U14318 (N_14318,N_13873,N_13883);
or U14319 (N_14319,N_13816,N_13546);
xor U14320 (N_14320,N_13596,N_13959);
xnor U14321 (N_14321,N_13535,N_13649);
nand U14322 (N_14322,N_13853,N_13570);
nand U14323 (N_14323,N_13519,N_13916);
xnor U14324 (N_14324,N_13783,N_13748);
xor U14325 (N_14325,N_13551,N_13541);
nor U14326 (N_14326,N_13671,N_13894);
and U14327 (N_14327,N_13536,N_13616);
nand U14328 (N_14328,N_13724,N_13882);
xnor U14329 (N_14329,N_13872,N_13797);
and U14330 (N_14330,N_13762,N_13678);
nor U14331 (N_14331,N_13860,N_13698);
or U14332 (N_14332,N_13974,N_13719);
nand U14333 (N_14333,N_13638,N_13987);
xnor U14334 (N_14334,N_13568,N_13875);
or U14335 (N_14335,N_13509,N_13557);
xor U14336 (N_14336,N_13785,N_13854);
nand U14337 (N_14337,N_13609,N_13990);
and U14338 (N_14338,N_13705,N_13739);
nand U14339 (N_14339,N_13989,N_13565);
nand U14340 (N_14340,N_13597,N_13540);
nor U14341 (N_14341,N_13802,N_13750);
and U14342 (N_14342,N_13893,N_13737);
nand U14343 (N_14343,N_13754,N_13901);
and U14344 (N_14344,N_13852,N_13593);
and U14345 (N_14345,N_13771,N_13564);
and U14346 (N_14346,N_13600,N_13869);
nor U14347 (N_14347,N_13947,N_13839);
nor U14348 (N_14348,N_13619,N_13787);
and U14349 (N_14349,N_13776,N_13535);
and U14350 (N_14350,N_13984,N_13740);
or U14351 (N_14351,N_13781,N_13506);
nand U14352 (N_14352,N_13874,N_13617);
nor U14353 (N_14353,N_13674,N_13999);
or U14354 (N_14354,N_13645,N_13657);
xnor U14355 (N_14355,N_13518,N_13954);
xor U14356 (N_14356,N_13809,N_13773);
and U14357 (N_14357,N_13969,N_13802);
nand U14358 (N_14358,N_13832,N_13818);
nor U14359 (N_14359,N_13557,N_13943);
and U14360 (N_14360,N_13523,N_13906);
nand U14361 (N_14361,N_13980,N_13639);
or U14362 (N_14362,N_13935,N_13672);
and U14363 (N_14363,N_13640,N_13912);
xor U14364 (N_14364,N_13660,N_13875);
nand U14365 (N_14365,N_13599,N_13844);
nand U14366 (N_14366,N_13900,N_13781);
xor U14367 (N_14367,N_13557,N_13977);
nor U14368 (N_14368,N_13664,N_13717);
and U14369 (N_14369,N_13870,N_13928);
xnor U14370 (N_14370,N_13832,N_13535);
nor U14371 (N_14371,N_13799,N_13792);
nor U14372 (N_14372,N_13944,N_13551);
nand U14373 (N_14373,N_13877,N_13943);
xor U14374 (N_14374,N_13628,N_13615);
or U14375 (N_14375,N_13561,N_13607);
xor U14376 (N_14376,N_13647,N_13910);
or U14377 (N_14377,N_13670,N_13920);
nor U14378 (N_14378,N_13975,N_13880);
nand U14379 (N_14379,N_13820,N_13712);
nand U14380 (N_14380,N_13527,N_13582);
xnor U14381 (N_14381,N_13570,N_13716);
nand U14382 (N_14382,N_13513,N_13893);
or U14383 (N_14383,N_13994,N_13551);
nand U14384 (N_14384,N_13782,N_13651);
or U14385 (N_14385,N_13805,N_13920);
or U14386 (N_14386,N_13719,N_13529);
nor U14387 (N_14387,N_13904,N_13783);
or U14388 (N_14388,N_13602,N_13539);
xor U14389 (N_14389,N_13671,N_13500);
and U14390 (N_14390,N_13913,N_13954);
nor U14391 (N_14391,N_13994,N_13658);
and U14392 (N_14392,N_13912,N_13884);
or U14393 (N_14393,N_13557,N_13844);
nor U14394 (N_14394,N_13972,N_13863);
and U14395 (N_14395,N_13515,N_13955);
nor U14396 (N_14396,N_13563,N_13826);
nor U14397 (N_14397,N_13668,N_13541);
nor U14398 (N_14398,N_13924,N_13672);
and U14399 (N_14399,N_13546,N_13564);
nand U14400 (N_14400,N_13640,N_13779);
nand U14401 (N_14401,N_13542,N_13653);
nand U14402 (N_14402,N_13975,N_13877);
nand U14403 (N_14403,N_13891,N_13915);
or U14404 (N_14404,N_13784,N_13598);
xnor U14405 (N_14405,N_13772,N_13843);
and U14406 (N_14406,N_13567,N_13747);
nor U14407 (N_14407,N_13752,N_13689);
or U14408 (N_14408,N_13769,N_13555);
nand U14409 (N_14409,N_13663,N_13748);
nand U14410 (N_14410,N_13802,N_13982);
nand U14411 (N_14411,N_13904,N_13897);
xnor U14412 (N_14412,N_13803,N_13998);
xnor U14413 (N_14413,N_13980,N_13775);
or U14414 (N_14414,N_13994,N_13535);
and U14415 (N_14415,N_13581,N_13918);
or U14416 (N_14416,N_13991,N_13517);
and U14417 (N_14417,N_13704,N_13715);
nand U14418 (N_14418,N_13844,N_13819);
nand U14419 (N_14419,N_13625,N_13543);
and U14420 (N_14420,N_13829,N_13666);
xnor U14421 (N_14421,N_13843,N_13616);
nand U14422 (N_14422,N_13766,N_13991);
and U14423 (N_14423,N_13994,N_13679);
and U14424 (N_14424,N_13506,N_13528);
xor U14425 (N_14425,N_13690,N_13741);
xnor U14426 (N_14426,N_13773,N_13607);
nor U14427 (N_14427,N_13970,N_13694);
and U14428 (N_14428,N_13648,N_13522);
and U14429 (N_14429,N_13620,N_13856);
xor U14430 (N_14430,N_13673,N_13608);
xnor U14431 (N_14431,N_13618,N_13544);
xnor U14432 (N_14432,N_13791,N_13690);
or U14433 (N_14433,N_13656,N_13724);
xnor U14434 (N_14434,N_13790,N_13949);
or U14435 (N_14435,N_13661,N_13719);
xnor U14436 (N_14436,N_13965,N_13672);
xor U14437 (N_14437,N_13622,N_13755);
nor U14438 (N_14438,N_13735,N_13584);
and U14439 (N_14439,N_13702,N_13738);
nand U14440 (N_14440,N_13562,N_13866);
and U14441 (N_14441,N_13859,N_13864);
xor U14442 (N_14442,N_13588,N_13528);
xnor U14443 (N_14443,N_13738,N_13931);
and U14444 (N_14444,N_13770,N_13937);
or U14445 (N_14445,N_13814,N_13670);
or U14446 (N_14446,N_13952,N_13863);
or U14447 (N_14447,N_13546,N_13554);
or U14448 (N_14448,N_13876,N_13697);
and U14449 (N_14449,N_13759,N_13527);
xor U14450 (N_14450,N_13651,N_13691);
or U14451 (N_14451,N_13808,N_13526);
xnor U14452 (N_14452,N_13683,N_13746);
nand U14453 (N_14453,N_13552,N_13933);
nor U14454 (N_14454,N_13907,N_13665);
nor U14455 (N_14455,N_13799,N_13964);
nand U14456 (N_14456,N_13697,N_13710);
nand U14457 (N_14457,N_13904,N_13843);
and U14458 (N_14458,N_13503,N_13796);
nor U14459 (N_14459,N_13546,N_13714);
nand U14460 (N_14460,N_13547,N_13687);
nor U14461 (N_14461,N_13714,N_13699);
nor U14462 (N_14462,N_13542,N_13874);
nor U14463 (N_14463,N_13895,N_13598);
nand U14464 (N_14464,N_13630,N_13724);
or U14465 (N_14465,N_13720,N_13542);
xnor U14466 (N_14466,N_13927,N_13958);
nor U14467 (N_14467,N_13548,N_13628);
and U14468 (N_14468,N_13622,N_13728);
or U14469 (N_14469,N_13893,N_13755);
nor U14470 (N_14470,N_13733,N_13634);
and U14471 (N_14471,N_13595,N_13825);
nand U14472 (N_14472,N_13630,N_13558);
xnor U14473 (N_14473,N_13893,N_13706);
and U14474 (N_14474,N_13643,N_13570);
or U14475 (N_14475,N_13810,N_13915);
and U14476 (N_14476,N_13587,N_13525);
xor U14477 (N_14477,N_13937,N_13745);
xor U14478 (N_14478,N_13730,N_13813);
nor U14479 (N_14479,N_13727,N_13874);
xor U14480 (N_14480,N_13868,N_13665);
nand U14481 (N_14481,N_13915,N_13790);
or U14482 (N_14482,N_13611,N_13802);
or U14483 (N_14483,N_13988,N_13781);
xor U14484 (N_14484,N_13742,N_13898);
and U14485 (N_14485,N_13864,N_13602);
nand U14486 (N_14486,N_13987,N_13742);
and U14487 (N_14487,N_13834,N_13878);
nand U14488 (N_14488,N_13855,N_13848);
or U14489 (N_14489,N_13810,N_13643);
nand U14490 (N_14490,N_13977,N_13538);
nor U14491 (N_14491,N_13959,N_13966);
and U14492 (N_14492,N_13843,N_13902);
and U14493 (N_14493,N_13974,N_13660);
or U14494 (N_14494,N_13814,N_13544);
and U14495 (N_14495,N_13520,N_13607);
or U14496 (N_14496,N_13937,N_13966);
or U14497 (N_14497,N_13540,N_13873);
or U14498 (N_14498,N_13943,N_13739);
and U14499 (N_14499,N_13687,N_13514);
xor U14500 (N_14500,N_14466,N_14087);
nor U14501 (N_14501,N_14454,N_14113);
nor U14502 (N_14502,N_14024,N_14203);
and U14503 (N_14503,N_14261,N_14047);
or U14504 (N_14504,N_14268,N_14478);
nor U14505 (N_14505,N_14145,N_14419);
nand U14506 (N_14506,N_14151,N_14218);
and U14507 (N_14507,N_14140,N_14273);
nand U14508 (N_14508,N_14306,N_14220);
nand U14509 (N_14509,N_14107,N_14102);
or U14510 (N_14510,N_14452,N_14252);
nand U14511 (N_14511,N_14115,N_14118);
and U14512 (N_14512,N_14355,N_14235);
and U14513 (N_14513,N_14396,N_14223);
nor U14514 (N_14514,N_14176,N_14077);
nand U14515 (N_14515,N_14373,N_14301);
and U14516 (N_14516,N_14324,N_14479);
and U14517 (N_14517,N_14021,N_14084);
and U14518 (N_14518,N_14428,N_14397);
and U14519 (N_14519,N_14362,N_14269);
nor U14520 (N_14520,N_14376,N_14061);
nor U14521 (N_14521,N_14097,N_14048);
nand U14522 (N_14522,N_14039,N_14333);
xor U14523 (N_14523,N_14049,N_14193);
or U14524 (N_14524,N_14357,N_14144);
nor U14525 (N_14525,N_14210,N_14133);
nand U14526 (N_14526,N_14074,N_14109);
nor U14527 (N_14527,N_14225,N_14310);
or U14528 (N_14528,N_14425,N_14316);
nand U14529 (N_14529,N_14449,N_14286);
or U14530 (N_14530,N_14023,N_14068);
or U14531 (N_14531,N_14209,N_14386);
xnor U14532 (N_14532,N_14058,N_14293);
nor U14533 (N_14533,N_14250,N_14228);
nor U14534 (N_14534,N_14100,N_14358);
or U14535 (N_14535,N_14050,N_14407);
or U14536 (N_14536,N_14240,N_14089);
xnor U14537 (N_14537,N_14244,N_14088);
and U14538 (N_14538,N_14305,N_14142);
or U14539 (N_14539,N_14206,N_14067);
xor U14540 (N_14540,N_14405,N_14290);
nand U14541 (N_14541,N_14062,N_14344);
nor U14542 (N_14542,N_14483,N_14046);
or U14543 (N_14543,N_14326,N_14359);
nand U14544 (N_14544,N_14274,N_14494);
nor U14545 (N_14545,N_14280,N_14124);
or U14546 (N_14546,N_14146,N_14270);
nand U14547 (N_14547,N_14410,N_14330);
nor U14548 (N_14548,N_14338,N_14471);
nand U14549 (N_14549,N_14229,N_14092);
nor U14550 (N_14550,N_14308,N_14367);
nand U14551 (N_14551,N_14042,N_14184);
nor U14552 (N_14552,N_14003,N_14219);
nand U14553 (N_14553,N_14304,N_14159);
or U14554 (N_14554,N_14031,N_14093);
and U14555 (N_14555,N_14251,N_14423);
and U14556 (N_14556,N_14297,N_14319);
or U14557 (N_14557,N_14231,N_14400);
xor U14558 (N_14558,N_14444,N_14379);
nor U14559 (N_14559,N_14139,N_14360);
or U14560 (N_14560,N_14439,N_14365);
xnor U14561 (N_14561,N_14421,N_14096);
nor U14562 (N_14562,N_14129,N_14177);
xnor U14563 (N_14563,N_14034,N_14447);
and U14564 (N_14564,N_14432,N_14291);
xor U14565 (N_14565,N_14288,N_14493);
xor U14566 (N_14566,N_14180,N_14117);
nor U14567 (N_14567,N_14311,N_14472);
nand U14568 (N_14568,N_14434,N_14295);
or U14569 (N_14569,N_14267,N_14227);
and U14570 (N_14570,N_14128,N_14166);
nor U14571 (N_14571,N_14005,N_14320);
or U14572 (N_14572,N_14491,N_14266);
nor U14573 (N_14573,N_14299,N_14429);
or U14574 (N_14574,N_14053,N_14202);
nand U14575 (N_14575,N_14325,N_14236);
nand U14576 (N_14576,N_14336,N_14382);
nor U14577 (N_14577,N_14232,N_14181);
nor U14578 (N_14578,N_14294,N_14450);
nor U14579 (N_14579,N_14322,N_14374);
nor U14580 (N_14580,N_14329,N_14403);
xnor U14581 (N_14581,N_14019,N_14127);
nand U14582 (N_14582,N_14198,N_14340);
or U14583 (N_14583,N_14343,N_14287);
or U14584 (N_14584,N_14247,N_14368);
nor U14585 (N_14585,N_14207,N_14440);
xor U14586 (N_14586,N_14060,N_14038);
or U14587 (N_14587,N_14073,N_14285);
or U14588 (N_14588,N_14474,N_14378);
nor U14589 (N_14589,N_14197,N_14243);
xnor U14590 (N_14590,N_14221,N_14485);
nor U14591 (N_14591,N_14189,N_14211);
or U14592 (N_14592,N_14204,N_14347);
nor U14593 (N_14593,N_14424,N_14114);
and U14594 (N_14594,N_14462,N_14131);
and U14595 (N_14595,N_14433,N_14278);
xor U14596 (N_14596,N_14385,N_14111);
xnor U14597 (N_14597,N_14409,N_14103);
xnor U14598 (N_14598,N_14352,N_14191);
nand U14599 (N_14599,N_14249,N_14464);
or U14600 (N_14600,N_14354,N_14026);
nor U14601 (N_14601,N_14253,N_14040);
nand U14602 (N_14602,N_14430,N_14482);
nand U14603 (N_14603,N_14081,N_14143);
nand U14604 (N_14604,N_14190,N_14417);
nor U14605 (N_14605,N_14392,N_14296);
and U14606 (N_14606,N_14463,N_14028);
nor U14607 (N_14607,N_14468,N_14427);
nor U14608 (N_14608,N_14486,N_14036);
xnor U14609 (N_14609,N_14363,N_14342);
xnor U14610 (N_14610,N_14254,N_14230);
nand U14611 (N_14611,N_14130,N_14317);
and U14612 (N_14612,N_14256,N_14004);
and U14613 (N_14613,N_14125,N_14484);
nand U14614 (N_14614,N_14281,N_14263);
nor U14615 (N_14615,N_14199,N_14361);
and U14616 (N_14616,N_14442,N_14276);
xnor U14617 (N_14617,N_14303,N_14105);
nand U14618 (N_14618,N_14056,N_14262);
and U14619 (N_14619,N_14033,N_14018);
and U14620 (N_14620,N_14108,N_14496);
and U14621 (N_14621,N_14346,N_14436);
and U14622 (N_14622,N_14137,N_14331);
or U14623 (N_14623,N_14315,N_14161);
or U14624 (N_14624,N_14116,N_14149);
or U14625 (N_14625,N_14134,N_14371);
and U14626 (N_14626,N_14110,N_14214);
nor U14627 (N_14627,N_14292,N_14313);
nand U14628 (N_14628,N_14298,N_14183);
xor U14629 (N_14629,N_14422,N_14160);
or U14630 (N_14630,N_14171,N_14489);
nor U14631 (N_14631,N_14233,N_14123);
nor U14632 (N_14632,N_14101,N_14328);
nand U14633 (N_14633,N_14196,N_14321);
nand U14634 (N_14634,N_14339,N_14453);
nor U14635 (N_14635,N_14488,N_14394);
or U14636 (N_14636,N_14009,N_14165);
xnor U14637 (N_14637,N_14175,N_14408);
or U14638 (N_14638,N_14002,N_14112);
nor U14639 (N_14639,N_14476,N_14029);
xor U14640 (N_14640,N_14337,N_14045);
nor U14641 (N_14641,N_14446,N_14217);
or U14642 (N_14642,N_14390,N_14154);
or U14643 (N_14643,N_14099,N_14226);
nor U14644 (N_14644,N_14282,N_14356);
and U14645 (N_14645,N_14377,N_14495);
nor U14646 (N_14646,N_14451,N_14467);
nand U14647 (N_14647,N_14259,N_14415);
nand U14648 (N_14648,N_14272,N_14212);
xor U14649 (N_14649,N_14201,N_14258);
nor U14650 (N_14650,N_14079,N_14375);
xnor U14651 (N_14651,N_14312,N_14348);
and U14652 (N_14652,N_14063,N_14426);
nor U14653 (N_14653,N_14260,N_14025);
and U14654 (N_14654,N_14470,N_14119);
xor U14655 (N_14655,N_14148,N_14309);
xnor U14656 (N_14656,N_14186,N_14072);
nor U14657 (N_14657,N_14401,N_14323);
nor U14658 (N_14658,N_14008,N_14492);
nor U14659 (N_14659,N_14384,N_14168);
or U14660 (N_14660,N_14413,N_14064);
nor U14661 (N_14661,N_14445,N_14086);
or U14662 (N_14662,N_14490,N_14037);
nand U14663 (N_14663,N_14366,N_14167);
nand U14664 (N_14664,N_14138,N_14469);
and U14665 (N_14665,N_14411,N_14153);
nand U14666 (N_14666,N_14314,N_14477);
or U14667 (N_14667,N_14136,N_14279);
xnor U14668 (N_14668,N_14017,N_14182);
nand U14669 (N_14669,N_14289,N_14091);
xnor U14670 (N_14670,N_14006,N_14497);
xor U14671 (N_14671,N_14398,N_14179);
xor U14672 (N_14672,N_14126,N_14054);
or U14673 (N_14673,N_14481,N_14032);
or U14674 (N_14674,N_14345,N_14335);
or U14675 (N_14675,N_14275,N_14458);
nand U14676 (N_14676,N_14157,N_14412);
xnor U14677 (N_14677,N_14195,N_14265);
nor U14678 (N_14678,N_14465,N_14349);
xor U14679 (N_14679,N_14106,N_14395);
and U14680 (N_14680,N_14372,N_14135);
and U14681 (N_14681,N_14420,N_14381);
or U14682 (N_14682,N_14155,N_14069);
nor U14683 (N_14683,N_14030,N_14461);
nand U14684 (N_14684,N_14076,N_14192);
xnor U14685 (N_14685,N_14122,N_14011);
nor U14686 (N_14686,N_14150,N_14334);
and U14687 (N_14687,N_14383,N_14431);
xnor U14688 (N_14688,N_14010,N_14443);
nand U14689 (N_14689,N_14215,N_14070);
or U14690 (N_14690,N_14041,N_14255);
nand U14691 (N_14691,N_14350,N_14205);
xnor U14692 (N_14692,N_14438,N_14075);
nand U14693 (N_14693,N_14237,N_14059);
and U14694 (N_14694,N_14162,N_14082);
nor U14695 (N_14695,N_14104,N_14185);
xor U14696 (N_14696,N_14012,N_14277);
nand U14697 (N_14697,N_14085,N_14245);
nand U14698 (N_14698,N_14460,N_14393);
xnor U14699 (N_14699,N_14456,N_14035);
xnor U14700 (N_14700,N_14257,N_14441);
nand U14701 (N_14701,N_14013,N_14007);
xor U14702 (N_14702,N_14455,N_14351);
xor U14703 (N_14703,N_14459,N_14200);
nand U14704 (N_14704,N_14057,N_14271);
nor U14705 (N_14705,N_14475,N_14078);
and U14706 (N_14706,N_14435,N_14353);
and U14707 (N_14707,N_14173,N_14234);
nand U14708 (N_14708,N_14389,N_14147);
nor U14709 (N_14709,N_14132,N_14065);
xnor U14710 (N_14710,N_14283,N_14238);
or U14711 (N_14711,N_14187,N_14169);
xor U14712 (N_14712,N_14498,N_14055);
nor U14713 (N_14713,N_14341,N_14208);
xor U14714 (N_14714,N_14188,N_14364);
and U14715 (N_14715,N_14152,N_14213);
and U14716 (N_14716,N_14307,N_14080);
nand U14717 (N_14717,N_14216,N_14222);
nand U14718 (N_14718,N_14332,N_14090);
xnor U14719 (N_14719,N_14248,N_14418);
xor U14720 (N_14720,N_14020,N_14302);
nand U14721 (N_14721,N_14300,N_14380);
and U14722 (N_14722,N_14014,N_14448);
xor U14723 (N_14723,N_14000,N_14094);
or U14724 (N_14724,N_14242,N_14178);
and U14725 (N_14725,N_14416,N_14194);
xor U14726 (N_14726,N_14241,N_14327);
nor U14727 (N_14727,N_14120,N_14391);
and U14728 (N_14728,N_14387,N_14095);
nor U14729 (N_14729,N_14174,N_14499);
and U14730 (N_14730,N_14121,N_14246);
nand U14731 (N_14731,N_14370,N_14027);
or U14732 (N_14732,N_14052,N_14043);
nor U14733 (N_14733,N_14016,N_14480);
nand U14734 (N_14734,N_14156,N_14071);
nand U14735 (N_14735,N_14158,N_14284);
or U14736 (N_14736,N_14164,N_14264);
and U14737 (N_14737,N_14404,N_14015);
or U14738 (N_14738,N_14044,N_14141);
xor U14739 (N_14739,N_14239,N_14163);
or U14740 (N_14740,N_14437,N_14487);
and U14741 (N_14741,N_14172,N_14414);
or U14742 (N_14742,N_14399,N_14406);
xor U14743 (N_14743,N_14001,N_14318);
xor U14744 (N_14744,N_14457,N_14369);
xnor U14745 (N_14745,N_14170,N_14224);
and U14746 (N_14746,N_14066,N_14388);
or U14747 (N_14747,N_14473,N_14022);
nand U14748 (N_14748,N_14402,N_14083);
and U14749 (N_14749,N_14051,N_14098);
nand U14750 (N_14750,N_14284,N_14018);
and U14751 (N_14751,N_14427,N_14356);
or U14752 (N_14752,N_14481,N_14219);
or U14753 (N_14753,N_14303,N_14092);
xor U14754 (N_14754,N_14284,N_14473);
xor U14755 (N_14755,N_14060,N_14483);
xnor U14756 (N_14756,N_14187,N_14477);
or U14757 (N_14757,N_14008,N_14078);
xor U14758 (N_14758,N_14097,N_14211);
xnor U14759 (N_14759,N_14290,N_14384);
xor U14760 (N_14760,N_14281,N_14321);
xnor U14761 (N_14761,N_14409,N_14347);
nand U14762 (N_14762,N_14186,N_14384);
or U14763 (N_14763,N_14057,N_14021);
and U14764 (N_14764,N_14098,N_14386);
xor U14765 (N_14765,N_14216,N_14226);
xor U14766 (N_14766,N_14076,N_14405);
and U14767 (N_14767,N_14088,N_14157);
or U14768 (N_14768,N_14157,N_14211);
and U14769 (N_14769,N_14006,N_14262);
xnor U14770 (N_14770,N_14169,N_14271);
nand U14771 (N_14771,N_14148,N_14361);
xnor U14772 (N_14772,N_14299,N_14160);
nand U14773 (N_14773,N_14179,N_14450);
nor U14774 (N_14774,N_14382,N_14030);
or U14775 (N_14775,N_14015,N_14135);
or U14776 (N_14776,N_14054,N_14110);
nor U14777 (N_14777,N_14441,N_14159);
and U14778 (N_14778,N_14218,N_14109);
nor U14779 (N_14779,N_14074,N_14041);
xor U14780 (N_14780,N_14268,N_14290);
nand U14781 (N_14781,N_14283,N_14378);
nand U14782 (N_14782,N_14400,N_14132);
or U14783 (N_14783,N_14121,N_14241);
nor U14784 (N_14784,N_14268,N_14087);
xor U14785 (N_14785,N_14155,N_14435);
nor U14786 (N_14786,N_14431,N_14445);
xnor U14787 (N_14787,N_14017,N_14085);
nand U14788 (N_14788,N_14065,N_14210);
nor U14789 (N_14789,N_14122,N_14085);
and U14790 (N_14790,N_14379,N_14325);
or U14791 (N_14791,N_14266,N_14195);
or U14792 (N_14792,N_14189,N_14282);
xnor U14793 (N_14793,N_14190,N_14175);
nand U14794 (N_14794,N_14384,N_14077);
xor U14795 (N_14795,N_14083,N_14043);
nor U14796 (N_14796,N_14486,N_14481);
nor U14797 (N_14797,N_14361,N_14287);
xnor U14798 (N_14798,N_14277,N_14371);
nand U14799 (N_14799,N_14349,N_14470);
and U14800 (N_14800,N_14158,N_14011);
nor U14801 (N_14801,N_14485,N_14450);
nor U14802 (N_14802,N_14073,N_14386);
and U14803 (N_14803,N_14071,N_14321);
xnor U14804 (N_14804,N_14392,N_14234);
nor U14805 (N_14805,N_14409,N_14183);
or U14806 (N_14806,N_14350,N_14326);
nor U14807 (N_14807,N_14386,N_14035);
or U14808 (N_14808,N_14364,N_14142);
and U14809 (N_14809,N_14019,N_14291);
xnor U14810 (N_14810,N_14426,N_14056);
nor U14811 (N_14811,N_14446,N_14466);
nor U14812 (N_14812,N_14354,N_14395);
xor U14813 (N_14813,N_14269,N_14129);
or U14814 (N_14814,N_14005,N_14314);
xnor U14815 (N_14815,N_14448,N_14156);
or U14816 (N_14816,N_14238,N_14379);
xnor U14817 (N_14817,N_14077,N_14227);
nor U14818 (N_14818,N_14273,N_14475);
or U14819 (N_14819,N_14347,N_14486);
xnor U14820 (N_14820,N_14086,N_14120);
and U14821 (N_14821,N_14244,N_14351);
nand U14822 (N_14822,N_14484,N_14463);
and U14823 (N_14823,N_14019,N_14002);
nor U14824 (N_14824,N_14089,N_14482);
nor U14825 (N_14825,N_14217,N_14389);
nand U14826 (N_14826,N_14344,N_14197);
xnor U14827 (N_14827,N_14420,N_14436);
nand U14828 (N_14828,N_14073,N_14343);
or U14829 (N_14829,N_14451,N_14135);
nand U14830 (N_14830,N_14321,N_14013);
and U14831 (N_14831,N_14080,N_14264);
or U14832 (N_14832,N_14439,N_14065);
nand U14833 (N_14833,N_14366,N_14009);
and U14834 (N_14834,N_14028,N_14054);
xnor U14835 (N_14835,N_14095,N_14090);
nand U14836 (N_14836,N_14493,N_14190);
nand U14837 (N_14837,N_14429,N_14267);
and U14838 (N_14838,N_14215,N_14467);
xor U14839 (N_14839,N_14372,N_14085);
and U14840 (N_14840,N_14154,N_14356);
nand U14841 (N_14841,N_14196,N_14345);
and U14842 (N_14842,N_14162,N_14006);
and U14843 (N_14843,N_14080,N_14210);
nand U14844 (N_14844,N_14441,N_14107);
or U14845 (N_14845,N_14311,N_14404);
xnor U14846 (N_14846,N_14422,N_14015);
and U14847 (N_14847,N_14448,N_14457);
nand U14848 (N_14848,N_14329,N_14472);
and U14849 (N_14849,N_14418,N_14490);
and U14850 (N_14850,N_14132,N_14242);
nor U14851 (N_14851,N_14010,N_14228);
nor U14852 (N_14852,N_14016,N_14433);
xor U14853 (N_14853,N_14262,N_14304);
nor U14854 (N_14854,N_14046,N_14202);
or U14855 (N_14855,N_14184,N_14286);
nor U14856 (N_14856,N_14116,N_14135);
nor U14857 (N_14857,N_14131,N_14085);
or U14858 (N_14858,N_14236,N_14277);
and U14859 (N_14859,N_14371,N_14175);
xor U14860 (N_14860,N_14274,N_14237);
and U14861 (N_14861,N_14431,N_14059);
nor U14862 (N_14862,N_14289,N_14224);
or U14863 (N_14863,N_14374,N_14488);
nand U14864 (N_14864,N_14328,N_14409);
and U14865 (N_14865,N_14241,N_14038);
xor U14866 (N_14866,N_14144,N_14139);
xnor U14867 (N_14867,N_14317,N_14323);
nor U14868 (N_14868,N_14143,N_14301);
xnor U14869 (N_14869,N_14164,N_14292);
and U14870 (N_14870,N_14416,N_14003);
nand U14871 (N_14871,N_14453,N_14395);
nor U14872 (N_14872,N_14439,N_14421);
nand U14873 (N_14873,N_14188,N_14252);
nor U14874 (N_14874,N_14388,N_14376);
xor U14875 (N_14875,N_14206,N_14285);
and U14876 (N_14876,N_14330,N_14067);
nand U14877 (N_14877,N_14075,N_14193);
and U14878 (N_14878,N_14054,N_14362);
nand U14879 (N_14879,N_14309,N_14393);
xor U14880 (N_14880,N_14117,N_14213);
or U14881 (N_14881,N_14225,N_14133);
xnor U14882 (N_14882,N_14074,N_14321);
nand U14883 (N_14883,N_14096,N_14139);
nor U14884 (N_14884,N_14141,N_14465);
nand U14885 (N_14885,N_14422,N_14227);
or U14886 (N_14886,N_14147,N_14304);
or U14887 (N_14887,N_14296,N_14088);
and U14888 (N_14888,N_14058,N_14483);
nand U14889 (N_14889,N_14326,N_14118);
or U14890 (N_14890,N_14026,N_14235);
xor U14891 (N_14891,N_14197,N_14162);
or U14892 (N_14892,N_14045,N_14368);
xor U14893 (N_14893,N_14125,N_14323);
or U14894 (N_14894,N_14346,N_14108);
nor U14895 (N_14895,N_14055,N_14409);
nand U14896 (N_14896,N_14223,N_14016);
and U14897 (N_14897,N_14286,N_14252);
nand U14898 (N_14898,N_14100,N_14041);
xnor U14899 (N_14899,N_14379,N_14194);
xnor U14900 (N_14900,N_14463,N_14398);
and U14901 (N_14901,N_14311,N_14206);
xor U14902 (N_14902,N_14279,N_14395);
and U14903 (N_14903,N_14208,N_14048);
xor U14904 (N_14904,N_14039,N_14452);
or U14905 (N_14905,N_14430,N_14235);
nor U14906 (N_14906,N_14419,N_14147);
and U14907 (N_14907,N_14450,N_14380);
xor U14908 (N_14908,N_14425,N_14191);
and U14909 (N_14909,N_14448,N_14052);
nor U14910 (N_14910,N_14446,N_14334);
and U14911 (N_14911,N_14196,N_14135);
nor U14912 (N_14912,N_14284,N_14343);
xnor U14913 (N_14913,N_14292,N_14472);
nor U14914 (N_14914,N_14223,N_14170);
nand U14915 (N_14915,N_14375,N_14303);
nor U14916 (N_14916,N_14052,N_14153);
nand U14917 (N_14917,N_14377,N_14405);
nor U14918 (N_14918,N_14030,N_14100);
and U14919 (N_14919,N_14468,N_14262);
nor U14920 (N_14920,N_14340,N_14350);
nor U14921 (N_14921,N_14000,N_14246);
nor U14922 (N_14922,N_14348,N_14373);
or U14923 (N_14923,N_14008,N_14067);
nand U14924 (N_14924,N_14315,N_14326);
nor U14925 (N_14925,N_14083,N_14483);
xnor U14926 (N_14926,N_14246,N_14152);
nor U14927 (N_14927,N_14495,N_14402);
or U14928 (N_14928,N_14256,N_14321);
xor U14929 (N_14929,N_14238,N_14284);
nor U14930 (N_14930,N_14401,N_14397);
or U14931 (N_14931,N_14414,N_14011);
xnor U14932 (N_14932,N_14133,N_14136);
nor U14933 (N_14933,N_14007,N_14252);
nor U14934 (N_14934,N_14130,N_14263);
or U14935 (N_14935,N_14002,N_14051);
nand U14936 (N_14936,N_14021,N_14460);
nor U14937 (N_14937,N_14396,N_14058);
xor U14938 (N_14938,N_14062,N_14072);
nor U14939 (N_14939,N_14185,N_14168);
or U14940 (N_14940,N_14472,N_14460);
or U14941 (N_14941,N_14253,N_14459);
nand U14942 (N_14942,N_14207,N_14270);
xor U14943 (N_14943,N_14083,N_14448);
and U14944 (N_14944,N_14426,N_14235);
xor U14945 (N_14945,N_14068,N_14266);
xnor U14946 (N_14946,N_14329,N_14391);
and U14947 (N_14947,N_14353,N_14180);
nand U14948 (N_14948,N_14498,N_14245);
xor U14949 (N_14949,N_14296,N_14150);
or U14950 (N_14950,N_14497,N_14458);
nor U14951 (N_14951,N_14169,N_14308);
nand U14952 (N_14952,N_14480,N_14040);
and U14953 (N_14953,N_14106,N_14123);
xor U14954 (N_14954,N_14374,N_14444);
nand U14955 (N_14955,N_14029,N_14465);
nor U14956 (N_14956,N_14135,N_14055);
and U14957 (N_14957,N_14076,N_14114);
nand U14958 (N_14958,N_14201,N_14065);
and U14959 (N_14959,N_14468,N_14181);
nand U14960 (N_14960,N_14154,N_14060);
nand U14961 (N_14961,N_14105,N_14200);
or U14962 (N_14962,N_14325,N_14138);
xor U14963 (N_14963,N_14295,N_14416);
nor U14964 (N_14964,N_14243,N_14360);
or U14965 (N_14965,N_14342,N_14422);
or U14966 (N_14966,N_14171,N_14005);
nand U14967 (N_14967,N_14361,N_14465);
nand U14968 (N_14968,N_14098,N_14413);
or U14969 (N_14969,N_14479,N_14457);
nor U14970 (N_14970,N_14141,N_14457);
nor U14971 (N_14971,N_14440,N_14186);
and U14972 (N_14972,N_14437,N_14068);
nor U14973 (N_14973,N_14429,N_14189);
xor U14974 (N_14974,N_14063,N_14015);
and U14975 (N_14975,N_14199,N_14031);
and U14976 (N_14976,N_14135,N_14141);
nand U14977 (N_14977,N_14438,N_14294);
or U14978 (N_14978,N_14302,N_14247);
xnor U14979 (N_14979,N_14368,N_14331);
xnor U14980 (N_14980,N_14015,N_14012);
and U14981 (N_14981,N_14167,N_14146);
nand U14982 (N_14982,N_14274,N_14395);
nor U14983 (N_14983,N_14099,N_14351);
xor U14984 (N_14984,N_14457,N_14331);
and U14985 (N_14985,N_14312,N_14395);
nand U14986 (N_14986,N_14493,N_14379);
nor U14987 (N_14987,N_14492,N_14012);
nor U14988 (N_14988,N_14158,N_14315);
and U14989 (N_14989,N_14188,N_14047);
or U14990 (N_14990,N_14354,N_14258);
or U14991 (N_14991,N_14101,N_14369);
nand U14992 (N_14992,N_14476,N_14223);
xor U14993 (N_14993,N_14020,N_14015);
xor U14994 (N_14994,N_14477,N_14488);
nand U14995 (N_14995,N_14022,N_14191);
or U14996 (N_14996,N_14021,N_14441);
nor U14997 (N_14997,N_14284,N_14222);
nand U14998 (N_14998,N_14434,N_14142);
xor U14999 (N_14999,N_14308,N_14266);
nor U15000 (N_15000,N_14643,N_14952);
xor U15001 (N_15001,N_14743,N_14505);
nor U15002 (N_15002,N_14798,N_14636);
nor U15003 (N_15003,N_14672,N_14913);
and U15004 (N_15004,N_14546,N_14508);
or U15005 (N_15005,N_14825,N_14610);
and U15006 (N_15006,N_14565,N_14753);
and U15007 (N_15007,N_14554,N_14662);
or U15008 (N_15008,N_14593,N_14831);
or U15009 (N_15009,N_14755,N_14735);
and U15010 (N_15010,N_14917,N_14980);
nor U15011 (N_15011,N_14993,N_14550);
or U15012 (N_15012,N_14630,N_14804);
and U15013 (N_15013,N_14608,N_14632);
nor U15014 (N_15014,N_14561,N_14797);
and U15015 (N_15015,N_14674,N_14939);
nand U15016 (N_15016,N_14585,N_14663);
and U15017 (N_15017,N_14745,N_14951);
xor U15018 (N_15018,N_14877,N_14789);
xor U15019 (N_15019,N_14973,N_14620);
or U15020 (N_15020,N_14599,N_14527);
and U15021 (N_15021,N_14556,N_14640);
nand U15022 (N_15022,N_14580,N_14639);
and U15023 (N_15023,N_14734,N_14953);
nor U15024 (N_15024,N_14905,N_14901);
nor U15025 (N_15025,N_14757,N_14523);
or U15026 (N_15026,N_14704,N_14719);
and U15027 (N_15027,N_14591,N_14826);
nor U15028 (N_15028,N_14827,N_14821);
xnor U15029 (N_15029,N_14881,N_14856);
nor U15030 (N_15030,N_14794,N_14967);
xor U15031 (N_15031,N_14616,N_14852);
xnor U15032 (N_15032,N_14851,N_14687);
and U15033 (N_15033,N_14812,N_14539);
nor U15034 (N_15034,N_14989,N_14916);
and U15035 (N_15035,N_14680,N_14511);
or U15036 (N_15036,N_14850,N_14665);
and U15037 (N_15037,N_14892,N_14834);
and U15038 (N_15038,N_14518,N_14691);
xor U15039 (N_15039,N_14992,N_14818);
and U15040 (N_15040,N_14710,N_14517);
xor U15041 (N_15041,N_14525,N_14840);
and U15042 (N_15042,N_14654,N_14646);
nor U15043 (N_15043,N_14739,N_14957);
and U15044 (N_15044,N_14693,N_14996);
xnor U15045 (N_15045,N_14648,N_14614);
or U15046 (N_15046,N_14664,N_14965);
and U15047 (N_15047,N_14833,N_14857);
or U15048 (N_15048,N_14716,N_14947);
and U15049 (N_15049,N_14775,N_14863);
and U15050 (N_15050,N_14923,N_14893);
nor U15051 (N_15051,N_14751,N_14962);
nand U15052 (N_15052,N_14650,N_14873);
xnor U15053 (N_15053,N_14995,N_14990);
nand U15054 (N_15054,N_14669,N_14619);
xnor U15055 (N_15055,N_14549,N_14964);
and U15056 (N_15056,N_14657,N_14879);
nand U15057 (N_15057,N_14933,N_14559);
xnor U15058 (N_15058,N_14586,N_14595);
nand U15059 (N_15059,N_14543,N_14786);
xor U15060 (N_15060,N_14661,N_14617);
or U15061 (N_15061,N_14538,N_14972);
nor U15062 (N_15062,N_14724,N_14911);
nand U15063 (N_15063,N_14584,N_14869);
or U15064 (N_15064,N_14747,N_14988);
nand U15065 (N_15065,N_14723,N_14532);
or U15066 (N_15066,N_14545,N_14820);
and U15067 (N_15067,N_14981,N_14612);
xnor U15068 (N_15068,N_14712,N_14598);
or U15069 (N_15069,N_14813,N_14829);
nor U15070 (N_15070,N_14501,N_14768);
nand U15071 (N_15071,N_14793,N_14887);
or U15072 (N_15072,N_14603,N_14621);
nand U15073 (N_15073,N_14854,N_14656);
and U15074 (N_15074,N_14777,N_14866);
and U15075 (N_15075,N_14961,N_14782);
and U15076 (N_15076,N_14645,N_14823);
xnor U15077 (N_15077,N_14513,N_14909);
nor U15078 (N_15078,N_14781,N_14904);
or U15079 (N_15079,N_14932,N_14903);
or U15080 (N_15080,N_14531,N_14582);
or U15081 (N_15081,N_14875,N_14861);
xnor U15082 (N_15082,N_14708,N_14884);
nor U15083 (N_15083,N_14600,N_14711);
xnor U15084 (N_15084,N_14537,N_14948);
and U15085 (N_15085,N_14890,N_14926);
xnor U15086 (N_15086,N_14722,N_14690);
or U15087 (N_15087,N_14713,N_14737);
xor U15088 (N_15088,N_14516,N_14571);
xor U15089 (N_15089,N_14970,N_14845);
and U15090 (N_15090,N_14795,N_14928);
or U15091 (N_15091,N_14900,N_14925);
nand U15092 (N_15092,N_14730,N_14566);
xor U15093 (N_15093,N_14849,N_14929);
xnor U15094 (N_15094,N_14945,N_14898);
or U15095 (N_15095,N_14936,N_14882);
xnor U15096 (N_15096,N_14971,N_14703);
xor U15097 (N_15097,N_14935,N_14968);
xnor U15098 (N_15098,N_14848,N_14897);
and U15099 (N_15099,N_14579,N_14644);
and U15100 (N_15100,N_14689,N_14668);
nor U15101 (N_15101,N_14853,N_14696);
xnor U15102 (N_15102,N_14637,N_14752);
nor U15103 (N_15103,N_14540,N_14805);
xor U15104 (N_15104,N_14569,N_14670);
nand U15105 (N_15105,N_14756,N_14528);
nor U15106 (N_15106,N_14762,N_14800);
nor U15107 (N_15107,N_14914,N_14938);
or U15108 (N_15108,N_14548,N_14717);
nor U15109 (N_15109,N_14628,N_14767);
nor U15110 (N_15110,N_14623,N_14727);
xnor U15111 (N_15111,N_14783,N_14512);
xnor U15112 (N_15112,N_14846,N_14758);
and U15113 (N_15113,N_14924,N_14822);
xor U15114 (N_15114,N_14847,N_14570);
xnor U15115 (N_15115,N_14740,N_14977);
or U15116 (N_15116,N_14720,N_14799);
nand U15117 (N_15117,N_14682,N_14659);
xnor U15118 (N_15118,N_14551,N_14563);
xnor U15119 (N_15119,N_14785,N_14955);
nand U15120 (N_15120,N_14660,N_14694);
or U15121 (N_15121,N_14838,N_14702);
nand U15122 (N_15122,N_14746,N_14934);
xnor U15123 (N_15123,N_14773,N_14560);
and U15124 (N_15124,N_14521,N_14606);
and U15125 (N_15125,N_14792,N_14918);
nand U15126 (N_15126,N_14759,N_14842);
nand U15127 (N_15127,N_14986,N_14906);
or U15128 (N_15128,N_14984,N_14673);
nand U15129 (N_15129,N_14994,N_14985);
or U15130 (N_15130,N_14524,N_14862);
and U15131 (N_15131,N_14679,N_14557);
nor U15132 (N_15132,N_14567,N_14983);
xnor U15133 (N_15133,N_14878,N_14611);
nor U15134 (N_15134,N_14533,N_14754);
and U15135 (N_15135,N_14681,N_14987);
and U15136 (N_15136,N_14509,N_14613);
nor U15137 (N_15137,N_14707,N_14627);
nand U15138 (N_15138,N_14806,N_14975);
nor U15139 (N_15139,N_14819,N_14676);
nand U15140 (N_15140,N_14653,N_14808);
or U15141 (N_15141,N_14715,N_14809);
xor U15142 (N_15142,N_14535,N_14705);
and U15143 (N_15143,N_14652,N_14578);
nand U15144 (N_15144,N_14562,N_14700);
nor U15145 (N_15145,N_14868,N_14576);
and U15146 (N_15146,N_14506,N_14976);
nor U15147 (N_15147,N_14859,N_14675);
or U15148 (N_15148,N_14718,N_14891);
or U15149 (N_15149,N_14649,N_14536);
nand U15150 (N_15150,N_14922,N_14733);
xor U15151 (N_15151,N_14515,N_14769);
nand U15152 (N_15152,N_14592,N_14688);
nand U15153 (N_15153,N_14966,N_14625);
or U15154 (N_15154,N_14522,N_14507);
xor U15155 (N_15155,N_14896,N_14695);
nor U15156 (N_15156,N_14858,N_14774);
or U15157 (N_15157,N_14692,N_14589);
nand U15158 (N_15158,N_14500,N_14763);
nand U15159 (N_15159,N_14969,N_14633);
nand U15160 (N_15160,N_14779,N_14944);
xor U15161 (N_15161,N_14658,N_14997);
nor U15162 (N_15162,N_14738,N_14915);
xor U15163 (N_15163,N_14889,N_14817);
and U15164 (N_15164,N_14635,N_14671);
and U15165 (N_15165,N_14504,N_14602);
nor U15166 (N_15166,N_14796,N_14736);
xnor U15167 (N_15167,N_14729,N_14583);
or U15168 (N_15168,N_14942,N_14553);
and U15169 (N_15169,N_14855,N_14828);
nor U15170 (N_15170,N_14655,N_14830);
or U15171 (N_15171,N_14581,N_14765);
or U15172 (N_15172,N_14860,N_14555);
and U15173 (N_15173,N_14921,N_14954);
or U15174 (N_15174,N_14683,N_14941);
nand U15175 (N_15175,N_14638,N_14502);
and U15176 (N_15176,N_14697,N_14801);
nor U15177 (N_15177,N_14999,N_14959);
nor U15178 (N_15178,N_14963,N_14514);
nand U15179 (N_15179,N_14641,N_14815);
xor U15180 (N_15180,N_14824,N_14931);
or U15181 (N_15181,N_14686,N_14749);
nor U15182 (N_15182,N_14547,N_14764);
or U15183 (N_15183,N_14605,N_14978);
or U15184 (N_15184,N_14766,N_14910);
or U15185 (N_15185,N_14940,N_14698);
or U15186 (N_15186,N_14744,N_14872);
nand U15187 (N_15187,N_14902,N_14564);
nand U15188 (N_15188,N_14802,N_14886);
and U15189 (N_15189,N_14732,N_14750);
or U15190 (N_15190,N_14885,N_14776);
or U15191 (N_15191,N_14642,N_14832);
nor U15192 (N_15192,N_14958,N_14721);
nand U15193 (N_15193,N_14597,N_14526);
and U15194 (N_15194,N_14519,N_14907);
xnor U15195 (N_15195,N_14510,N_14651);
nand U15196 (N_15196,N_14725,N_14596);
xor U15197 (N_15197,N_14574,N_14974);
nor U15198 (N_15198,N_14629,N_14647);
nand U15199 (N_15199,N_14667,N_14634);
nor U15200 (N_15200,N_14920,N_14544);
xor U15201 (N_15201,N_14979,N_14709);
and U15202 (N_15202,N_14714,N_14899);
or U15203 (N_15203,N_14677,N_14876);
nor U15204 (N_15204,N_14631,N_14609);
nor U15205 (N_15205,N_14760,N_14844);
nand U15206 (N_15206,N_14573,N_14741);
or U15207 (N_15207,N_14731,N_14807);
or U15208 (N_15208,N_14685,N_14864);
nand U15209 (N_15209,N_14810,N_14699);
xor U15210 (N_15210,N_14927,N_14624);
or U15211 (N_15211,N_14706,N_14865);
or U15212 (N_15212,N_14874,N_14930);
nor U15213 (N_15213,N_14787,N_14894);
or U15214 (N_15214,N_14888,N_14542);
nor U15215 (N_15215,N_14895,N_14520);
or U15216 (N_15216,N_14960,N_14761);
nand U15217 (N_15217,N_14814,N_14778);
and U15218 (N_15218,N_14836,N_14588);
nor U15219 (N_15219,N_14982,N_14587);
nand U15220 (N_15220,N_14788,N_14530);
and U15221 (N_15221,N_14558,N_14771);
xnor U15222 (N_15222,N_14784,N_14811);
nand U15223 (N_15223,N_14912,N_14883);
and U15224 (N_15224,N_14956,N_14835);
and U15225 (N_15225,N_14577,N_14837);
xor U15226 (N_15226,N_14791,N_14946);
nand U15227 (N_15227,N_14880,N_14622);
nand U15228 (N_15228,N_14803,N_14568);
or U15229 (N_15229,N_14594,N_14839);
xnor U15230 (N_15230,N_14678,N_14728);
xnor U15231 (N_15231,N_14503,N_14618);
xor U15232 (N_15232,N_14534,N_14816);
and U15233 (N_15233,N_14943,N_14867);
nand U15234 (N_15234,N_14601,N_14572);
or U15235 (N_15235,N_14748,N_14772);
and U15236 (N_15236,N_14529,N_14991);
nand U15237 (N_15237,N_14908,N_14841);
nand U15238 (N_15238,N_14871,N_14870);
or U15239 (N_15239,N_14949,N_14950);
and U15240 (N_15240,N_14998,N_14552);
nor U15241 (N_15241,N_14937,N_14726);
and U15242 (N_15242,N_14607,N_14541);
and U15243 (N_15243,N_14590,N_14742);
xor U15244 (N_15244,N_14701,N_14790);
and U15245 (N_15245,N_14843,N_14684);
and U15246 (N_15246,N_14780,N_14666);
nor U15247 (N_15247,N_14615,N_14626);
nor U15248 (N_15248,N_14919,N_14575);
and U15249 (N_15249,N_14604,N_14770);
nor U15250 (N_15250,N_14893,N_14859);
or U15251 (N_15251,N_14696,N_14597);
nand U15252 (N_15252,N_14870,N_14883);
xor U15253 (N_15253,N_14597,N_14515);
and U15254 (N_15254,N_14562,N_14648);
and U15255 (N_15255,N_14924,N_14548);
and U15256 (N_15256,N_14608,N_14950);
nor U15257 (N_15257,N_14714,N_14716);
xnor U15258 (N_15258,N_14599,N_14672);
and U15259 (N_15259,N_14880,N_14593);
xnor U15260 (N_15260,N_14707,N_14569);
or U15261 (N_15261,N_14737,N_14680);
nor U15262 (N_15262,N_14980,N_14652);
or U15263 (N_15263,N_14513,N_14769);
xnor U15264 (N_15264,N_14770,N_14759);
nand U15265 (N_15265,N_14631,N_14983);
xnor U15266 (N_15266,N_14692,N_14687);
and U15267 (N_15267,N_14573,N_14760);
or U15268 (N_15268,N_14833,N_14746);
xor U15269 (N_15269,N_14986,N_14577);
or U15270 (N_15270,N_14654,N_14576);
and U15271 (N_15271,N_14854,N_14825);
nor U15272 (N_15272,N_14990,N_14774);
nand U15273 (N_15273,N_14972,N_14881);
nor U15274 (N_15274,N_14992,N_14581);
and U15275 (N_15275,N_14828,N_14856);
nand U15276 (N_15276,N_14843,N_14705);
nand U15277 (N_15277,N_14504,N_14895);
nand U15278 (N_15278,N_14520,N_14805);
nand U15279 (N_15279,N_14996,N_14839);
and U15280 (N_15280,N_14693,N_14969);
nor U15281 (N_15281,N_14673,N_14765);
nand U15282 (N_15282,N_14778,N_14969);
or U15283 (N_15283,N_14730,N_14704);
xor U15284 (N_15284,N_14940,N_14664);
nand U15285 (N_15285,N_14782,N_14705);
or U15286 (N_15286,N_14588,N_14553);
nor U15287 (N_15287,N_14656,N_14628);
xor U15288 (N_15288,N_14729,N_14843);
xor U15289 (N_15289,N_14724,N_14795);
xor U15290 (N_15290,N_14980,N_14787);
nand U15291 (N_15291,N_14561,N_14535);
or U15292 (N_15292,N_14793,N_14619);
nand U15293 (N_15293,N_14535,N_14860);
or U15294 (N_15294,N_14853,N_14594);
nor U15295 (N_15295,N_14787,N_14713);
xor U15296 (N_15296,N_14940,N_14841);
or U15297 (N_15297,N_14826,N_14869);
and U15298 (N_15298,N_14635,N_14979);
and U15299 (N_15299,N_14615,N_14600);
or U15300 (N_15300,N_14898,N_14943);
xnor U15301 (N_15301,N_14603,N_14696);
nand U15302 (N_15302,N_14854,N_14871);
nor U15303 (N_15303,N_14653,N_14638);
nor U15304 (N_15304,N_14799,N_14764);
nand U15305 (N_15305,N_14525,N_14586);
nor U15306 (N_15306,N_14740,N_14709);
nand U15307 (N_15307,N_14934,N_14702);
nand U15308 (N_15308,N_14547,N_14563);
nand U15309 (N_15309,N_14860,N_14738);
nand U15310 (N_15310,N_14619,N_14713);
nand U15311 (N_15311,N_14591,N_14694);
nand U15312 (N_15312,N_14994,N_14751);
xor U15313 (N_15313,N_14605,N_14682);
nand U15314 (N_15314,N_14619,N_14749);
xnor U15315 (N_15315,N_14546,N_14789);
nor U15316 (N_15316,N_14872,N_14665);
xnor U15317 (N_15317,N_14837,N_14836);
nor U15318 (N_15318,N_14722,N_14718);
xnor U15319 (N_15319,N_14542,N_14949);
nand U15320 (N_15320,N_14709,N_14752);
nand U15321 (N_15321,N_14559,N_14751);
nor U15322 (N_15322,N_14563,N_14983);
and U15323 (N_15323,N_14756,N_14567);
xnor U15324 (N_15324,N_14582,N_14529);
nand U15325 (N_15325,N_14857,N_14516);
or U15326 (N_15326,N_14824,N_14749);
nor U15327 (N_15327,N_14996,N_14924);
and U15328 (N_15328,N_14684,N_14890);
or U15329 (N_15329,N_14536,N_14763);
or U15330 (N_15330,N_14660,N_14620);
nor U15331 (N_15331,N_14769,N_14994);
nor U15332 (N_15332,N_14548,N_14734);
and U15333 (N_15333,N_14610,N_14939);
xnor U15334 (N_15334,N_14641,N_14760);
nor U15335 (N_15335,N_14625,N_14616);
and U15336 (N_15336,N_14958,N_14828);
or U15337 (N_15337,N_14644,N_14915);
and U15338 (N_15338,N_14785,N_14819);
xnor U15339 (N_15339,N_14677,N_14514);
or U15340 (N_15340,N_14580,N_14964);
or U15341 (N_15341,N_14944,N_14699);
and U15342 (N_15342,N_14638,N_14892);
nand U15343 (N_15343,N_14893,N_14579);
or U15344 (N_15344,N_14829,N_14879);
nand U15345 (N_15345,N_14516,N_14705);
nand U15346 (N_15346,N_14771,N_14867);
nand U15347 (N_15347,N_14608,N_14904);
and U15348 (N_15348,N_14521,N_14604);
or U15349 (N_15349,N_14958,N_14634);
xor U15350 (N_15350,N_14685,N_14664);
nand U15351 (N_15351,N_14978,N_14762);
or U15352 (N_15352,N_14971,N_14581);
xnor U15353 (N_15353,N_14663,N_14825);
nand U15354 (N_15354,N_14821,N_14735);
xnor U15355 (N_15355,N_14711,N_14562);
or U15356 (N_15356,N_14578,N_14748);
xnor U15357 (N_15357,N_14999,N_14560);
nand U15358 (N_15358,N_14992,N_14815);
nor U15359 (N_15359,N_14692,N_14578);
nor U15360 (N_15360,N_14605,N_14937);
or U15361 (N_15361,N_14695,N_14790);
xnor U15362 (N_15362,N_14606,N_14504);
or U15363 (N_15363,N_14810,N_14533);
nand U15364 (N_15364,N_14666,N_14734);
or U15365 (N_15365,N_14669,N_14544);
nor U15366 (N_15366,N_14889,N_14609);
xnor U15367 (N_15367,N_14914,N_14847);
nor U15368 (N_15368,N_14895,N_14872);
and U15369 (N_15369,N_14613,N_14846);
or U15370 (N_15370,N_14692,N_14786);
and U15371 (N_15371,N_14513,N_14825);
or U15372 (N_15372,N_14978,N_14886);
xnor U15373 (N_15373,N_14692,N_14597);
nor U15374 (N_15374,N_14839,N_14620);
or U15375 (N_15375,N_14753,N_14883);
and U15376 (N_15376,N_14983,N_14595);
nor U15377 (N_15377,N_14909,N_14797);
and U15378 (N_15378,N_14608,N_14922);
and U15379 (N_15379,N_14791,N_14519);
nand U15380 (N_15380,N_14521,N_14753);
and U15381 (N_15381,N_14620,N_14915);
nor U15382 (N_15382,N_14877,N_14824);
and U15383 (N_15383,N_14671,N_14925);
nand U15384 (N_15384,N_14656,N_14706);
and U15385 (N_15385,N_14624,N_14803);
or U15386 (N_15386,N_14687,N_14781);
and U15387 (N_15387,N_14890,N_14840);
nand U15388 (N_15388,N_14819,N_14886);
xor U15389 (N_15389,N_14991,N_14748);
and U15390 (N_15390,N_14824,N_14514);
or U15391 (N_15391,N_14796,N_14541);
and U15392 (N_15392,N_14578,N_14706);
and U15393 (N_15393,N_14862,N_14929);
or U15394 (N_15394,N_14679,N_14843);
or U15395 (N_15395,N_14701,N_14717);
and U15396 (N_15396,N_14621,N_14588);
nor U15397 (N_15397,N_14942,N_14889);
nor U15398 (N_15398,N_14691,N_14807);
xnor U15399 (N_15399,N_14797,N_14957);
and U15400 (N_15400,N_14855,N_14587);
and U15401 (N_15401,N_14872,N_14966);
nor U15402 (N_15402,N_14741,N_14910);
xnor U15403 (N_15403,N_14613,N_14805);
xnor U15404 (N_15404,N_14978,N_14529);
xnor U15405 (N_15405,N_14955,N_14985);
and U15406 (N_15406,N_14684,N_14927);
nor U15407 (N_15407,N_14889,N_14800);
nand U15408 (N_15408,N_14831,N_14787);
or U15409 (N_15409,N_14572,N_14610);
or U15410 (N_15410,N_14734,N_14836);
and U15411 (N_15411,N_14922,N_14974);
xnor U15412 (N_15412,N_14877,N_14647);
or U15413 (N_15413,N_14660,N_14662);
nand U15414 (N_15414,N_14799,N_14696);
nor U15415 (N_15415,N_14922,N_14609);
and U15416 (N_15416,N_14810,N_14724);
and U15417 (N_15417,N_14648,N_14956);
and U15418 (N_15418,N_14923,N_14922);
nor U15419 (N_15419,N_14638,N_14718);
nor U15420 (N_15420,N_14528,N_14822);
nor U15421 (N_15421,N_14581,N_14567);
nor U15422 (N_15422,N_14567,N_14778);
or U15423 (N_15423,N_14630,N_14528);
or U15424 (N_15424,N_14621,N_14668);
and U15425 (N_15425,N_14594,N_14663);
or U15426 (N_15426,N_14624,N_14611);
xnor U15427 (N_15427,N_14523,N_14646);
or U15428 (N_15428,N_14939,N_14822);
nor U15429 (N_15429,N_14753,N_14701);
nor U15430 (N_15430,N_14981,N_14931);
nor U15431 (N_15431,N_14690,N_14799);
or U15432 (N_15432,N_14632,N_14691);
and U15433 (N_15433,N_14622,N_14654);
and U15434 (N_15434,N_14585,N_14782);
xor U15435 (N_15435,N_14679,N_14704);
xor U15436 (N_15436,N_14841,N_14721);
nor U15437 (N_15437,N_14685,N_14583);
nor U15438 (N_15438,N_14985,N_14863);
nand U15439 (N_15439,N_14591,N_14853);
or U15440 (N_15440,N_14991,N_14585);
and U15441 (N_15441,N_14510,N_14617);
and U15442 (N_15442,N_14930,N_14790);
and U15443 (N_15443,N_14568,N_14740);
xnor U15444 (N_15444,N_14932,N_14865);
and U15445 (N_15445,N_14598,N_14979);
nand U15446 (N_15446,N_14634,N_14791);
nand U15447 (N_15447,N_14876,N_14834);
nand U15448 (N_15448,N_14650,N_14722);
nand U15449 (N_15449,N_14905,N_14990);
and U15450 (N_15450,N_14895,N_14644);
nor U15451 (N_15451,N_14984,N_14924);
nor U15452 (N_15452,N_14732,N_14967);
nand U15453 (N_15453,N_14622,N_14750);
or U15454 (N_15454,N_14691,N_14845);
and U15455 (N_15455,N_14906,N_14606);
and U15456 (N_15456,N_14923,N_14885);
nor U15457 (N_15457,N_14949,N_14825);
or U15458 (N_15458,N_14732,N_14881);
nand U15459 (N_15459,N_14720,N_14861);
xor U15460 (N_15460,N_14712,N_14876);
nor U15461 (N_15461,N_14903,N_14875);
nand U15462 (N_15462,N_14642,N_14577);
nor U15463 (N_15463,N_14764,N_14947);
and U15464 (N_15464,N_14557,N_14522);
and U15465 (N_15465,N_14518,N_14566);
or U15466 (N_15466,N_14967,N_14572);
nand U15467 (N_15467,N_14949,N_14844);
or U15468 (N_15468,N_14504,N_14917);
nor U15469 (N_15469,N_14937,N_14679);
nand U15470 (N_15470,N_14998,N_14624);
xor U15471 (N_15471,N_14581,N_14923);
nor U15472 (N_15472,N_14584,N_14746);
and U15473 (N_15473,N_14780,N_14680);
or U15474 (N_15474,N_14757,N_14867);
and U15475 (N_15475,N_14540,N_14647);
nor U15476 (N_15476,N_14834,N_14601);
and U15477 (N_15477,N_14653,N_14561);
xor U15478 (N_15478,N_14666,N_14811);
nor U15479 (N_15479,N_14729,N_14721);
and U15480 (N_15480,N_14773,N_14825);
nand U15481 (N_15481,N_14934,N_14929);
xor U15482 (N_15482,N_14824,N_14778);
or U15483 (N_15483,N_14810,N_14725);
or U15484 (N_15484,N_14564,N_14695);
nand U15485 (N_15485,N_14554,N_14877);
nand U15486 (N_15486,N_14825,N_14682);
and U15487 (N_15487,N_14686,N_14739);
and U15488 (N_15488,N_14628,N_14654);
and U15489 (N_15489,N_14830,N_14759);
or U15490 (N_15490,N_14794,N_14741);
nor U15491 (N_15491,N_14700,N_14638);
or U15492 (N_15492,N_14977,N_14590);
nand U15493 (N_15493,N_14832,N_14675);
and U15494 (N_15494,N_14948,N_14950);
xnor U15495 (N_15495,N_14814,N_14921);
and U15496 (N_15496,N_14869,N_14608);
nand U15497 (N_15497,N_14520,N_14987);
and U15498 (N_15498,N_14632,N_14576);
and U15499 (N_15499,N_14694,N_14722);
and U15500 (N_15500,N_15433,N_15292);
nand U15501 (N_15501,N_15461,N_15259);
nor U15502 (N_15502,N_15148,N_15435);
nor U15503 (N_15503,N_15418,N_15086);
nor U15504 (N_15504,N_15049,N_15192);
and U15505 (N_15505,N_15145,N_15225);
and U15506 (N_15506,N_15173,N_15368);
nor U15507 (N_15507,N_15409,N_15016);
or U15508 (N_15508,N_15458,N_15208);
or U15509 (N_15509,N_15098,N_15227);
and U15510 (N_15510,N_15226,N_15353);
xor U15511 (N_15511,N_15338,N_15046);
nand U15512 (N_15512,N_15447,N_15381);
and U15513 (N_15513,N_15413,N_15432);
nand U15514 (N_15514,N_15481,N_15161);
and U15515 (N_15515,N_15350,N_15289);
or U15516 (N_15516,N_15277,N_15396);
xnor U15517 (N_15517,N_15464,N_15121);
nand U15518 (N_15518,N_15356,N_15184);
or U15519 (N_15519,N_15067,N_15278);
xor U15520 (N_15520,N_15238,N_15188);
nand U15521 (N_15521,N_15220,N_15203);
nor U15522 (N_15522,N_15460,N_15168);
nor U15523 (N_15523,N_15013,N_15354);
or U15524 (N_15524,N_15109,N_15079);
nor U15525 (N_15525,N_15267,N_15189);
nor U15526 (N_15526,N_15398,N_15101);
xnor U15527 (N_15527,N_15299,N_15175);
nand U15528 (N_15528,N_15323,N_15474);
xor U15529 (N_15529,N_15361,N_15296);
or U15530 (N_15530,N_15229,N_15454);
xor U15531 (N_15531,N_15139,N_15159);
nor U15532 (N_15532,N_15248,N_15141);
and U15533 (N_15533,N_15097,N_15253);
and U15534 (N_15534,N_15310,N_15463);
and U15535 (N_15535,N_15283,N_15151);
nor U15536 (N_15536,N_15216,N_15477);
xor U15537 (N_15537,N_15233,N_15077);
and U15538 (N_15538,N_15219,N_15024);
or U15539 (N_15539,N_15252,N_15450);
or U15540 (N_15540,N_15397,N_15230);
nand U15541 (N_15541,N_15351,N_15152);
nor U15542 (N_15542,N_15471,N_15130);
nand U15543 (N_15543,N_15053,N_15140);
or U15544 (N_15544,N_15105,N_15214);
and U15545 (N_15545,N_15282,N_15102);
or U15546 (N_15546,N_15254,N_15185);
nor U15547 (N_15547,N_15115,N_15123);
xnor U15548 (N_15548,N_15199,N_15134);
nor U15549 (N_15549,N_15399,N_15076);
and U15550 (N_15550,N_15269,N_15228);
and U15551 (N_15551,N_15059,N_15487);
nand U15552 (N_15552,N_15126,N_15094);
xnor U15553 (N_15553,N_15304,N_15411);
xnor U15554 (N_15554,N_15436,N_15057);
or U15555 (N_15555,N_15155,N_15324);
and U15556 (N_15556,N_15256,N_15172);
xor U15557 (N_15557,N_15313,N_15038);
nand U15558 (N_15558,N_15288,N_15273);
xor U15559 (N_15559,N_15497,N_15030);
or U15560 (N_15560,N_15430,N_15206);
nand U15561 (N_15561,N_15298,N_15062);
and U15562 (N_15562,N_15265,N_15111);
nor U15563 (N_15563,N_15327,N_15459);
or U15564 (N_15564,N_15328,N_15190);
xor U15565 (N_15565,N_15000,N_15349);
and U15566 (N_15566,N_15387,N_15498);
xnor U15567 (N_15567,N_15455,N_15096);
xnor U15568 (N_15568,N_15378,N_15008);
nor U15569 (N_15569,N_15309,N_15321);
xor U15570 (N_15570,N_15440,N_15001);
nor U15571 (N_15571,N_15007,N_15394);
xnor U15572 (N_15572,N_15065,N_15330);
or U15573 (N_15573,N_15493,N_15462);
and U15574 (N_15574,N_15197,N_15210);
xnor U15575 (N_15575,N_15372,N_15176);
nor U15576 (N_15576,N_15438,N_15090);
nor U15577 (N_15577,N_15043,N_15488);
xnor U15578 (N_15578,N_15293,N_15095);
nand U15579 (N_15579,N_15495,N_15202);
xnor U15580 (N_15580,N_15445,N_15177);
nand U15581 (N_15581,N_15200,N_15414);
or U15582 (N_15582,N_15364,N_15028);
nor U15583 (N_15583,N_15376,N_15224);
or U15584 (N_15584,N_15171,N_15118);
nand U15585 (N_15585,N_15110,N_15068);
nor U15586 (N_15586,N_15251,N_15261);
xnor U15587 (N_15587,N_15250,N_15431);
nand U15588 (N_15588,N_15335,N_15033);
nand U15589 (N_15589,N_15093,N_15205);
xor U15590 (N_15590,N_15017,N_15422);
and U15591 (N_15591,N_15476,N_15294);
nor U15592 (N_15592,N_15421,N_15204);
nand U15593 (N_15593,N_15044,N_15469);
or U15594 (N_15594,N_15083,N_15039);
and U15595 (N_15595,N_15218,N_15237);
xor U15596 (N_15596,N_15131,N_15339);
xnor U15597 (N_15597,N_15342,N_15272);
xor U15598 (N_15598,N_15449,N_15318);
nor U15599 (N_15599,N_15395,N_15085);
and U15600 (N_15600,N_15291,N_15164);
and U15601 (N_15601,N_15198,N_15280);
or U15602 (N_15602,N_15315,N_15078);
nand U15603 (N_15603,N_15392,N_15332);
nor U15604 (N_15604,N_15362,N_15036);
nand U15605 (N_15605,N_15325,N_15149);
nor U15606 (N_15606,N_15012,N_15014);
and U15607 (N_15607,N_15467,N_15120);
or U15608 (N_15608,N_15195,N_15169);
xor U15609 (N_15609,N_15334,N_15047);
and U15610 (N_15610,N_15271,N_15307);
and U15611 (N_15611,N_15371,N_15162);
xor U15612 (N_15612,N_15061,N_15147);
and U15613 (N_15613,N_15496,N_15041);
or U15614 (N_15614,N_15018,N_15236);
xnor U15615 (N_15615,N_15344,N_15346);
nor U15616 (N_15616,N_15006,N_15170);
nor U15617 (N_15617,N_15179,N_15402);
nor U15618 (N_15618,N_15405,N_15150);
xnor U15619 (N_15619,N_15404,N_15249);
xnor U15620 (N_15620,N_15287,N_15066);
nor U15621 (N_15621,N_15478,N_15015);
and U15622 (N_15622,N_15032,N_15329);
xnor U15623 (N_15623,N_15004,N_15138);
nor U15624 (N_15624,N_15305,N_15285);
nor U15625 (N_15625,N_15439,N_15358);
or U15626 (N_15626,N_15382,N_15040);
nand U15627 (N_15627,N_15196,N_15117);
or U15628 (N_15628,N_15391,N_15490);
nand U15629 (N_15629,N_15167,N_15146);
and U15630 (N_15630,N_15457,N_15142);
nor U15631 (N_15631,N_15181,N_15011);
nor U15632 (N_15632,N_15035,N_15133);
and U15633 (N_15633,N_15025,N_15367);
nor U15634 (N_15634,N_15489,N_15499);
nand U15635 (N_15635,N_15153,N_15400);
nor U15636 (N_15636,N_15240,N_15255);
nor U15637 (N_15637,N_15055,N_15160);
xnor U15638 (N_15638,N_15124,N_15482);
xor U15639 (N_15639,N_15108,N_15320);
nand U15640 (N_15640,N_15021,N_15451);
or U15641 (N_15641,N_15491,N_15116);
or U15642 (N_15642,N_15263,N_15388);
xnor U15643 (N_15643,N_15215,N_15485);
nor U15644 (N_15644,N_15275,N_15375);
nor U15645 (N_15645,N_15360,N_15026);
or U15646 (N_15646,N_15075,N_15416);
nor U15647 (N_15647,N_15379,N_15157);
and U15648 (N_15648,N_15027,N_15104);
nand U15649 (N_15649,N_15494,N_15366);
xor U15650 (N_15650,N_15089,N_15410);
or U15651 (N_15651,N_15442,N_15020);
nand U15652 (N_15652,N_15473,N_15306);
or U15653 (N_15653,N_15002,N_15034);
nand U15654 (N_15654,N_15322,N_15235);
xnor U15655 (N_15655,N_15303,N_15377);
xnor U15656 (N_15656,N_15088,N_15453);
or U15657 (N_15657,N_15401,N_15308);
and U15658 (N_15658,N_15212,N_15099);
xor U15659 (N_15659,N_15319,N_15174);
nand U15660 (N_15660,N_15073,N_15386);
and U15661 (N_15661,N_15279,N_15343);
nand U15662 (N_15662,N_15340,N_15191);
nor U15663 (N_15663,N_15213,N_15163);
nor U15664 (N_15664,N_15052,N_15129);
nor U15665 (N_15665,N_15486,N_15480);
and U15666 (N_15666,N_15128,N_15245);
or U15667 (N_15667,N_15448,N_15125);
nand U15668 (N_15668,N_15403,N_15302);
xnor U15669 (N_15669,N_15019,N_15470);
nand U15670 (N_15670,N_15472,N_15048);
or U15671 (N_15671,N_15426,N_15363);
and U15672 (N_15672,N_15301,N_15333);
xor U15673 (N_15673,N_15223,N_15080);
xnor U15674 (N_15674,N_15058,N_15003);
nand U15675 (N_15675,N_15187,N_15446);
nand U15676 (N_15676,N_15260,N_15370);
xor U15677 (N_15677,N_15060,N_15316);
xnor U15678 (N_15678,N_15234,N_15347);
nand U15679 (N_15679,N_15374,N_15064);
or U15680 (N_15680,N_15070,N_15087);
nand U15681 (N_15681,N_15326,N_15389);
nor U15682 (N_15682,N_15317,N_15465);
nor U15683 (N_15683,N_15373,N_15217);
and U15684 (N_15684,N_15297,N_15479);
and U15685 (N_15685,N_15434,N_15331);
and U15686 (N_15686,N_15425,N_15166);
nand U15687 (N_15687,N_15183,N_15010);
nand U15688 (N_15688,N_15103,N_15247);
and U15689 (N_15689,N_15136,N_15071);
or U15690 (N_15690,N_15452,N_15258);
nor U15691 (N_15691,N_15408,N_15132);
or U15692 (N_15692,N_15483,N_15050);
nand U15693 (N_15693,N_15295,N_15051);
nand U15694 (N_15694,N_15284,N_15312);
or U15695 (N_15695,N_15268,N_15031);
nand U15696 (N_15696,N_15385,N_15286);
xor U15697 (N_15697,N_15221,N_15201);
nor U15698 (N_15698,N_15009,N_15042);
or U15699 (N_15699,N_15054,N_15407);
nand U15700 (N_15700,N_15456,N_15154);
xor U15701 (N_15701,N_15074,N_15429);
xnor U15702 (N_15702,N_15135,N_15165);
xnor U15703 (N_15703,N_15415,N_15262);
nand U15704 (N_15704,N_15112,N_15243);
and U15705 (N_15705,N_15420,N_15137);
or U15706 (N_15706,N_15056,N_15266);
or U15707 (N_15707,N_15106,N_15127);
and U15708 (N_15708,N_15390,N_15100);
nand U15709 (N_15709,N_15383,N_15357);
nor U15710 (N_15710,N_15239,N_15029);
or U15711 (N_15711,N_15443,N_15264);
nor U15712 (N_15712,N_15311,N_15393);
or U15713 (N_15713,N_15182,N_15072);
xor U15714 (N_15714,N_15122,N_15257);
nand U15715 (N_15715,N_15276,N_15037);
nor U15716 (N_15716,N_15424,N_15437);
nand U15717 (N_15717,N_15492,N_15113);
xnor U15718 (N_15718,N_15186,N_15355);
nor U15719 (N_15719,N_15180,N_15144);
and U15720 (N_15720,N_15092,N_15069);
and U15721 (N_15721,N_15084,N_15337);
nand U15722 (N_15722,N_15081,N_15369);
or U15723 (N_15723,N_15352,N_15345);
or U15724 (N_15724,N_15246,N_15419);
or U15725 (N_15725,N_15441,N_15178);
nand U15726 (N_15726,N_15336,N_15468);
nor U15727 (N_15727,N_15274,N_15359);
nand U15728 (N_15728,N_15412,N_15005);
and U15729 (N_15729,N_15193,N_15091);
nand U15730 (N_15730,N_15444,N_15270);
nand U15731 (N_15731,N_15232,N_15143);
nand U15732 (N_15732,N_15281,N_15380);
and U15733 (N_15733,N_15475,N_15290);
nor U15734 (N_15734,N_15466,N_15207);
or U15735 (N_15735,N_15427,N_15314);
xor U15736 (N_15736,N_15022,N_15211);
xnor U15737 (N_15737,N_15023,N_15423);
and U15738 (N_15738,N_15158,N_15156);
nor U15739 (N_15739,N_15045,N_15300);
or U15740 (N_15740,N_15222,N_15242);
nor U15741 (N_15741,N_15063,N_15406);
nor U15742 (N_15742,N_15417,N_15365);
xnor U15743 (N_15743,N_15428,N_15384);
and U15744 (N_15744,N_15114,N_15082);
and U15745 (N_15745,N_15119,N_15231);
xnor U15746 (N_15746,N_15194,N_15209);
and U15747 (N_15747,N_15341,N_15107);
xor U15748 (N_15748,N_15484,N_15348);
nor U15749 (N_15749,N_15241,N_15244);
and U15750 (N_15750,N_15306,N_15497);
xor U15751 (N_15751,N_15312,N_15490);
nand U15752 (N_15752,N_15143,N_15060);
or U15753 (N_15753,N_15278,N_15162);
and U15754 (N_15754,N_15149,N_15038);
xor U15755 (N_15755,N_15089,N_15085);
or U15756 (N_15756,N_15189,N_15367);
and U15757 (N_15757,N_15238,N_15222);
nor U15758 (N_15758,N_15429,N_15428);
nor U15759 (N_15759,N_15195,N_15335);
xor U15760 (N_15760,N_15498,N_15306);
nand U15761 (N_15761,N_15112,N_15042);
nor U15762 (N_15762,N_15456,N_15146);
or U15763 (N_15763,N_15329,N_15409);
and U15764 (N_15764,N_15477,N_15443);
nor U15765 (N_15765,N_15405,N_15040);
xor U15766 (N_15766,N_15152,N_15136);
nand U15767 (N_15767,N_15251,N_15265);
or U15768 (N_15768,N_15123,N_15462);
nor U15769 (N_15769,N_15479,N_15095);
and U15770 (N_15770,N_15135,N_15108);
and U15771 (N_15771,N_15002,N_15475);
nor U15772 (N_15772,N_15070,N_15072);
nor U15773 (N_15773,N_15323,N_15183);
nor U15774 (N_15774,N_15065,N_15344);
or U15775 (N_15775,N_15027,N_15494);
and U15776 (N_15776,N_15336,N_15302);
and U15777 (N_15777,N_15144,N_15312);
and U15778 (N_15778,N_15291,N_15253);
nand U15779 (N_15779,N_15149,N_15121);
nor U15780 (N_15780,N_15274,N_15432);
nor U15781 (N_15781,N_15229,N_15257);
nand U15782 (N_15782,N_15412,N_15193);
nor U15783 (N_15783,N_15099,N_15240);
xor U15784 (N_15784,N_15414,N_15198);
and U15785 (N_15785,N_15009,N_15439);
xnor U15786 (N_15786,N_15231,N_15460);
xnor U15787 (N_15787,N_15229,N_15039);
nand U15788 (N_15788,N_15133,N_15041);
nand U15789 (N_15789,N_15424,N_15284);
xnor U15790 (N_15790,N_15381,N_15399);
or U15791 (N_15791,N_15261,N_15144);
nor U15792 (N_15792,N_15109,N_15179);
or U15793 (N_15793,N_15224,N_15131);
or U15794 (N_15794,N_15333,N_15270);
xnor U15795 (N_15795,N_15349,N_15453);
nand U15796 (N_15796,N_15415,N_15196);
nand U15797 (N_15797,N_15020,N_15469);
and U15798 (N_15798,N_15046,N_15195);
and U15799 (N_15799,N_15148,N_15429);
xor U15800 (N_15800,N_15158,N_15321);
xor U15801 (N_15801,N_15408,N_15218);
xor U15802 (N_15802,N_15127,N_15416);
or U15803 (N_15803,N_15352,N_15198);
and U15804 (N_15804,N_15229,N_15206);
xor U15805 (N_15805,N_15179,N_15349);
and U15806 (N_15806,N_15015,N_15433);
nor U15807 (N_15807,N_15399,N_15227);
and U15808 (N_15808,N_15396,N_15414);
xor U15809 (N_15809,N_15354,N_15136);
nor U15810 (N_15810,N_15198,N_15373);
or U15811 (N_15811,N_15280,N_15458);
nand U15812 (N_15812,N_15320,N_15303);
nand U15813 (N_15813,N_15020,N_15035);
nand U15814 (N_15814,N_15117,N_15235);
xnor U15815 (N_15815,N_15293,N_15295);
and U15816 (N_15816,N_15219,N_15084);
nand U15817 (N_15817,N_15199,N_15193);
nand U15818 (N_15818,N_15452,N_15416);
or U15819 (N_15819,N_15432,N_15097);
xor U15820 (N_15820,N_15481,N_15444);
nand U15821 (N_15821,N_15128,N_15445);
and U15822 (N_15822,N_15367,N_15425);
and U15823 (N_15823,N_15441,N_15485);
or U15824 (N_15824,N_15130,N_15436);
or U15825 (N_15825,N_15041,N_15095);
xnor U15826 (N_15826,N_15032,N_15043);
and U15827 (N_15827,N_15365,N_15043);
or U15828 (N_15828,N_15353,N_15061);
nor U15829 (N_15829,N_15041,N_15061);
xnor U15830 (N_15830,N_15243,N_15042);
nand U15831 (N_15831,N_15221,N_15159);
xnor U15832 (N_15832,N_15473,N_15124);
nor U15833 (N_15833,N_15240,N_15077);
and U15834 (N_15834,N_15260,N_15381);
or U15835 (N_15835,N_15173,N_15349);
and U15836 (N_15836,N_15285,N_15105);
and U15837 (N_15837,N_15296,N_15010);
or U15838 (N_15838,N_15447,N_15304);
or U15839 (N_15839,N_15020,N_15376);
nor U15840 (N_15840,N_15200,N_15279);
nor U15841 (N_15841,N_15449,N_15079);
and U15842 (N_15842,N_15328,N_15484);
nand U15843 (N_15843,N_15365,N_15153);
or U15844 (N_15844,N_15380,N_15267);
xor U15845 (N_15845,N_15154,N_15072);
or U15846 (N_15846,N_15101,N_15318);
nand U15847 (N_15847,N_15452,N_15175);
xnor U15848 (N_15848,N_15199,N_15316);
nor U15849 (N_15849,N_15191,N_15483);
xnor U15850 (N_15850,N_15024,N_15285);
and U15851 (N_15851,N_15166,N_15040);
or U15852 (N_15852,N_15010,N_15306);
or U15853 (N_15853,N_15422,N_15007);
or U15854 (N_15854,N_15006,N_15127);
or U15855 (N_15855,N_15470,N_15120);
and U15856 (N_15856,N_15367,N_15365);
nand U15857 (N_15857,N_15403,N_15358);
and U15858 (N_15858,N_15445,N_15327);
and U15859 (N_15859,N_15425,N_15313);
nor U15860 (N_15860,N_15046,N_15141);
nand U15861 (N_15861,N_15324,N_15358);
nor U15862 (N_15862,N_15249,N_15495);
or U15863 (N_15863,N_15070,N_15157);
xor U15864 (N_15864,N_15278,N_15263);
or U15865 (N_15865,N_15280,N_15150);
and U15866 (N_15866,N_15353,N_15128);
nor U15867 (N_15867,N_15140,N_15306);
or U15868 (N_15868,N_15356,N_15248);
and U15869 (N_15869,N_15427,N_15240);
and U15870 (N_15870,N_15342,N_15455);
or U15871 (N_15871,N_15422,N_15187);
nand U15872 (N_15872,N_15031,N_15475);
nor U15873 (N_15873,N_15143,N_15442);
or U15874 (N_15874,N_15371,N_15089);
or U15875 (N_15875,N_15020,N_15425);
nand U15876 (N_15876,N_15383,N_15156);
nand U15877 (N_15877,N_15109,N_15090);
nand U15878 (N_15878,N_15467,N_15319);
nand U15879 (N_15879,N_15091,N_15430);
and U15880 (N_15880,N_15387,N_15389);
nor U15881 (N_15881,N_15170,N_15362);
nor U15882 (N_15882,N_15384,N_15025);
and U15883 (N_15883,N_15495,N_15487);
and U15884 (N_15884,N_15466,N_15120);
or U15885 (N_15885,N_15193,N_15102);
and U15886 (N_15886,N_15076,N_15491);
or U15887 (N_15887,N_15050,N_15462);
nand U15888 (N_15888,N_15397,N_15062);
nor U15889 (N_15889,N_15188,N_15113);
nand U15890 (N_15890,N_15266,N_15173);
and U15891 (N_15891,N_15236,N_15414);
nand U15892 (N_15892,N_15392,N_15415);
xnor U15893 (N_15893,N_15302,N_15399);
or U15894 (N_15894,N_15321,N_15120);
or U15895 (N_15895,N_15046,N_15121);
or U15896 (N_15896,N_15470,N_15465);
and U15897 (N_15897,N_15223,N_15388);
and U15898 (N_15898,N_15229,N_15239);
nand U15899 (N_15899,N_15305,N_15268);
xor U15900 (N_15900,N_15355,N_15282);
xnor U15901 (N_15901,N_15425,N_15465);
nor U15902 (N_15902,N_15032,N_15197);
or U15903 (N_15903,N_15232,N_15382);
and U15904 (N_15904,N_15338,N_15099);
and U15905 (N_15905,N_15041,N_15336);
or U15906 (N_15906,N_15306,N_15407);
xor U15907 (N_15907,N_15437,N_15102);
nor U15908 (N_15908,N_15285,N_15373);
and U15909 (N_15909,N_15100,N_15143);
nor U15910 (N_15910,N_15474,N_15046);
or U15911 (N_15911,N_15206,N_15193);
or U15912 (N_15912,N_15082,N_15125);
and U15913 (N_15913,N_15225,N_15324);
xor U15914 (N_15914,N_15212,N_15033);
and U15915 (N_15915,N_15334,N_15328);
nor U15916 (N_15916,N_15365,N_15095);
xor U15917 (N_15917,N_15058,N_15133);
and U15918 (N_15918,N_15280,N_15356);
or U15919 (N_15919,N_15224,N_15439);
nor U15920 (N_15920,N_15259,N_15158);
nor U15921 (N_15921,N_15375,N_15448);
and U15922 (N_15922,N_15325,N_15492);
xor U15923 (N_15923,N_15499,N_15119);
or U15924 (N_15924,N_15032,N_15362);
nor U15925 (N_15925,N_15238,N_15358);
and U15926 (N_15926,N_15431,N_15264);
nor U15927 (N_15927,N_15121,N_15402);
xnor U15928 (N_15928,N_15348,N_15485);
or U15929 (N_15929,N_15115,N_15015);
and U15930 (N_15930,N_15344,N_15187);
nor U15931 (N_15931,N_15038,N_15081);
nor U15932 (N_15932,N_15173,N_15189);
nor U15933 (N_15933,N_15081,N_15395);
nand U15934 (N_15934,N_15398,N_15143);
or U15935 (N_15935,N_15275,N_15046);
nand U15936 (N_15936,N_15199,N_15400);
nor U15937 (N_15937,N_15245,N_15112);
or U15938 (N_15938,N_15258,N_15467);
or U15939 (N_15939,N_15005,N_15346);
nor U15940 (N_15940,N_15160,N_15490);
xnor U15941 (N_15941,N_15077,N_15441);
xnor U15942 (N_15942,N_15316,N_15217);
and U15943 (N_15943,N_15035,N_15013);
or U15944 (N_15944,N_15113,N_15327);
nand U15945 (N_15945,N_15363,N_15199);
xor U15946 (N_15946,N_15392,N_15237);
and U15947 (N_15947,N_15084,N_15077);
nor U15948 (N_15948,N_15218,N_15003);
or U15949 (N_15949,N_15413,N_15077);
or U15950 (N_15950,N_15325,N_15343);
xor U15951 (N_15951,N_15046,N_15233);
and U15952 (N_15952,N_15471,N_15008);
nand U15953 (N_15953,N_15477,N_15436);
xnor U15954 (N_15954,N_15467,N_15075);
nor U15955 (N_15955,N_15363,N_15319);
nor U15956 (N_15956,N_15480,N_15409);
nor U15957 (N_15957,N_15021,N_15117);
and U15958 (N_15958,N_15307,N_15093);
nor U15959 (N_15959,N_15220,N_15127);
nand U15960 (N_15960,N_15186,N_15087);
xor U15961 (N_15961,N_15475,N_15162);
nand U15962 (N_15962,N_15384,N_15206);
and U15963 (N_15963,N_15029,N_15130);
nand U15964 (N_15964,N_15294,N_15065);
nor U15965 (N_15965,N_15139,N_15281);
and U15966 (N_15966,N_15265,N_15012);
or U15967 (N_15967,N_15434,N_15490);
and U15968 (N_15968,N_15096,N_15229);
and U15969 (N_15969,N_15025,N_15327);
and U15970 (N_15970,N_15326,N_15139);
nand U15971 (N_15971,N_15463,N_15407);
and U15972 (N_15972,N_15346,N_15076);
nand U15973 (N_15973,N_15453,N_15332);
and U15974 (N_15974,N_15466,N_15094);
nand U15975 (N_15975,N_15281,N_15043);
and U15976 (N_15976,N_15296,N_15091);
nor U15977 (N_15977,N_15186,N_15032);
or U15978 (N_15978,N_15399,N_15409);
and U15979 (N_15979,N_15281,N_15409);
nor U15980 (N_15980,N_15262,N_15282);
xor U15981 (N_15981,N_15226,N_15010);
nor U15982 (N_15982,N_15381,N_15463);
nand U15983 (N_15983,N_15075,N_15151);
or U15984 (N_15984,N_15438,N_15445);
xor U15985 (N_15985,N_15218,N_15187);
xor U15986 (N_15986,N_15346,N_15430);
xnor U15987 (N_15987,N_15247,N_15256);
nor U15988 (N_15988,N_15102,N_15485);
or U15989 (N_15989,N_15351,N_15179);
and U15990 (N_15990,N_15480,N_15068);
or U15991 (N_15991,N_15163,N_15345);
nor U15992 (N_15992,N_15242,N_15381);
or U15993 (N_15993,N_15364,N_15245);
nor U15994 (N_15994,N_15061,N_15355);
and U15995 (N_15995,N_15136,N_15275);
and U15996 (N_15996,N_15413,N_15264);
nand U15997 (N_15997,N_15052,N_15304);
or U15998 (N_15998,N_15485,N_15451);
nor U15999 (N_15999,N_15394,N_15252);
or U16000 (N_16000,N_15638,N_15960);
nor U16001 (N_16001,N_15889,N_15553);
or U16002 (N_16002,N_15745,N_15757);
nand U16003 (N_16003,N_15985,N_15844);
xnor U16004 (N_16004,N_15552,N_15743);
nor U16005 (N_16005,N_15565,N_15878);
or U16006 (N_16006,N_15645,N_15585);
nand U16007 (N_16007,N_15504,N_15627);
xnor U16008 (N_16008,N_15704,N_15673);
or U16009 (N_16009,N_15635,N_15934);
xor U16010 (N_16010,N_15534,N_15539);
nor U16011 (N_16011,N_15897,N_15803);
nand U16012 (N_16012,N_15954,N_15778);
or U16013 (N_16013,N_15596,N_15707);
or U16014 (N_16014,N_15579,N_15871);
xor U16015 (N_16015,N_15508,N_15996);
nand U16016 (N_16016,N_15722,N_15516);
xor U16017 (N_16017,N_15631,N_15678);
or U16018 (N_16018,N_15905,N_15920);
nor U16019 (N_16019,N_15687,N_15930);
or U16020 (N_16020,N_15626,N_15587);
xnor U16021 (N_16021,N_15706,N_15511);
xor U16022 (N_16022,N_15894,N_15616);
or U16023 (N_16023,N_15559,N_15509);
nand U16024 (N_16024,N_15952,N_15606);
nand U16025 (N_16025,N_15829,N_15946);
nor U16026 (N_16026,N_15927,N_15551);
and U16027 (N_16027,N_15970,N_15835);
or U16028 (N_16028,N_15978,N_15964);
nor U16029 (N_16029,N_15681,N_15977);
xnor U16030 (N_16030,N_15953,N_15938);
nor U16031 (N_16031,N_15791,N_15965);
or U16032 (N_16032,N_15529,N_15676);
xnor U16033 (N_16033,N_15799,N_15562);
nand U16034 (N_16034,N_15518,N_15981);
nor U16035 (N_16035,N_15610,N_15522);
and U16036 (N_16036,N_15919,N_15991);
nor U16037 (N_16037,N_15775,N_15832);
or U16038 (N_16038,N_15726,N_15852);
nand U16039 (N_16039,N_15926,N_15860);
or U16040 (N_16040,N_15865,N_15692);
nor U16041 (N_16041,N_15914,N_15805);
nor U16042 (N_16042,N_15634,N_15575);
nor U16043 (N_16043,N_15910,N_15891);
xor U16044 (N_16044,N_15502,N_15881);
and U16045 (N_16045,N_15794,N_15724);
nor U16046 (N_16046,N_15694,N_15998);
and U16047 (N_16047,N_15615,N_15619);
nor U16048 (N_16048,N_15750,N_15813);
nand U16049 (N_16049,N_15679,N_15856);
or U16050 (N_16050,N_15877,N_15543);
and U16051 (N_16051,N_15641,N_15668);
xor U16052 (N_16052,N_15594,N_15849);
and U16053 (N_16053,N_15702,N_15963);
and U16054 (N_16054,N_15556,N_15672);
or U16055 (N_16055,N_15830,N_15741);
xnor U16056 (N_16056,N_15975,N_15931);
and U16057 (N_16057,N_15990,N_15908);
nand U16058 (N_16058,N_15736,N_15994);
and U16059 (N_16059,N_15503,N_15686);
and U16060 (N_16060,N_15505,N_15734);
xor U16061 (N_16061,N_15727,N_15818);
nand U16062 (N_16062,N_15958,N_15658);
or U16063 (N_16063,N_15842,N_15876);
or U16064 (N_16064,N_15657,N_15933);
xor U16065 (N_16065,N_15582,N_15886);
xnor U16066 (N_16066,N_15854,N_15797);
and U16067 (N_16067,N_15642,N_15697);
or U16068 (N_16068,N_15628,N_15513);
nor U16069 (N_16069,N_15901,N_15680);
nand U16070 (N_16070,N_15776,N_15535);
or U16071 (N_16071,N_15997,N_15721);
and U16072 (N_16072,N_15725,N_15753);
nand U16073 (N_16073,N_15758,N_15624);
nand U16074 (N_16074,N_15833,N_15730);
nand U16075 (N_16075,N_15817,N_15590);
or U16076 (N_16076,N_15760,N_15550);
nand U16077 (N_16077,N_15701,N_15523);
nand U16078 (N_16078,N_15524,N_15688);
nand U16079 (N_16079,N_15816,N_15696);
and U16080 (N_16080,N_15683,N_15782);
xor U16081 (N_16081,N_15913,N_15583);
and U16082 (N_16082,N_15731,N_15633);
nand U16083 (N_16083,N_15851,N_15577);
or U16084 (N_16084,N_15510,N_15995);
xnor U16085 (N_16085,N_15517,N_15784);
xnor U16086 (N_16086,N_15820,N_15671);
and U16087 (N_16087,N_15532,N_15549);
nor U16088 (N_16088,N_15564,N_15506);
nand U16089 (N_16089,N_15873,N_15648);
or U16090 (N_16090,N_15588,N_15838);
nand U16091 (N_16091,N_15869,N_15989);
and U16092 (N_16092,N_15917,N_15733);
nor U16093 (N_16093,N_15780,N_15774);
nor U16094 (N_16094,N_15858,N_15501);
and U16095 (N_16095,N_15685,N_15547);
and U16096 (N_16096,N_15812,N_15520);
nand U16097 (N_16097,N_15662,N_15793);
nor U16098 (N_16098,N_15567,N_15973);
nor U16099 (N_16099,N_15622,N_15800);
nand U16100 (N_16100,N_15868,N_15592);
or U16101 (N_16101,N_15738,N_15664);
or U16102 (N_16102,N_15767,N_15530);
and U16103 (N_16103,N_15762,N_15531);
xnor U16104 (N_16104,N_15843,N_15935);
nand U16105 (N_16105,N_15789,N_15841);
xor U16106 (N_16106,N_15831,N_15756);
and U16107 (N_16107,N_15863,N_15602);
xor U16108 (N_16108,N_15909,N_15732);
xor U16109 (N_16109,N_15893,N_15859);
nand U16110 (N_16110,N_15554,N_15608);
or U16111 (N_16111,N_15944,N_15809);
nor U16112 (N_16112,N_15742,N_15884);
nand U16113 (N_16113,N_15880,N_15751);
nand U16114 (N_16114,N_15922,N_15512);
nor U16115 (N_16115,N_15507,N_15866);
or U16116 (N_16116,N_15514,N_15705);
nand U16117 (N_16117,N_15693,N_15669);
and U16118 (N_16118,N_15650,N_15739);
nor U16119 (N_16119,N_15703,N_15867);
xor U16120 (N_16120,N_15644,N_15824);
or U16121 (N_16121,N_15661,N_15666);
nand U16122 (N_16122,N_15874,N_15923);
or U16123 (N_16123,N_15718,N_15617);
and U16124 (N_16124,N_15747,N_15620);
nand U16125 (N_16125,N_15828,N_15848);
and U16126 (N_16126,N_15546,N_15654);
or U16127 (N_16127,N_15561,N_15987);
nor U16128 (N_16128,N_15754,N_15779);
nor U16129 (N_16129,N_15538,N_15663);
xor U16130 (N_16130,N_15821,N_15968);
nand U16131 (N_16131,N_15875,N_15837);
or U16132 (N_16132,N_15630,N_15749);
nor U16133 (N_16133,N_15993,N_15898);
nor U16134 (N_16134,N_15639,N_15541);
nor U16135 (N_16135,N_15940,N_15864);
nand U16136 (N_16136,N_15568,N_15961);
and U16137 (N_16137,N_15887,N_15771);
and U16138 (N_16138,N_15902,N_15788);
or U16139 (N_16139,N_15607,N_15536);
and U16140 (N_16140,N_15971,N_15801);
nor U16141 (N_16141,N_15979,N_15907);
nand U16142 (N_16142,N_15895,N_15651);
nand U16143 (N_16143,N_15655,N_15807);
or U16144 (N_16144,N_15915,N_15573);
and U16145 (N_16145,N_15684,N_15647);
xor U16146 (N_16146,N_15956,N_15586);
nor U16147 (N_16147,N_15798,N_15951);
nand U16148 (N_16148,N_15834,N_15665);
xnor U16149 (N_16149,N_15735,N_15840);
and U16150 (N_16150,N_15815,N_15737);
or U16151 (N_16151,N_15636,N_15521);
or U16152 (N_16152,N_15770,N_15921);
or U16153 (N_16153,N_15755,N_15823);
xor U16154 (N_16154,N_15792,N_15597);
nand U16155 (N_16155,N_15611,N_15729);
xnor U16156 (N_16156,N_15677,N_15937);
nor U16157 (N_16157,N_15984,N_15584);
and U16158 (N_16158,N_15795,N_15716);
and U16159 (N_16159,N_15836,N_15717);
xor U16160 (N_16160,N_15912,N_15855);
nand U16161 (N_16161,N_15939,N_15572);
and U16162 (N_16162,N_15786,N_15708);
and U16163 (N_16163,N_15846,N_15896);
nand U16164 (N_16164,N_15527,N_15980);
xor U16165 (N_16165,N_15720,N_15787);
nand U16166 (N_16166,N_15746,N_15580);
nand U16167 (N_16167,N_15605,N_15571);
xnor U16168 (N_16168,N_15783,N_15764);
xnor U16169 (N_16169,N_15695,N_15728);
or U16170 (N_16170,N_15906,N_15804);
or U16171 (N_16171,N_15916,N_15942);
nand U16172 (N_16172,N_15675,N_15698);
and U16173 (N_16173,N_15621,N_15766);
xor U16174 (N_16174,N_15500,N_15777);
nor U16175 (N_16175,N_15637,N_15557);
and U16176 (N_16176,N_15936,N_15932);
xnor U16177 (N_16177,N_15850,N_15808);
and U16178 (N_16178,N_15781,N_15558);
nand U16179 (N_16179,N_15581,N_15542);
and U16180 (N_16180,N_15966,N_15814);
nand U16181 (N_16181,N_15623,N_15924);
or U16182 (N_16182,N_15879,N_15544);
nand U16183 (N_16183,N_15526,N_15691);
and U16184 (N_16184,N_15862,N_15853);
and U16185 (N_16185,N_15948,N_15670);
or U16186 (N_16186,N_15811,N_15659);
nand U16187 (N_16187,N_15759,N_15613);
or U16188 (N_16188,N_15545,N_15763);
nor U16189 (N_16189,N_15983,N_15992);
or U16190 (N_16190,N_15537,N_15822);
and U16191 (N_16191,N_15769,N_15819);
nor U16192 (N_16192,N_15892,N_15653);
nand U16193 (N_16193,N_15719,N_15682);
nor U16194 (N_16194,N_15625,N_15612);
and U16195 (N_16195,N_15962,N_15748);
and U16196 (N_16196,N_15576,N_15976);
nand U16197 (N_16197,N_15674,N_15882);
nor U16198 (N_16198,N_15941,N_15929);
nor U16199 (N_16199,N_15555,N_15918);
nor U16200 (N_16200,N_15861,N_15569);
or U16201 (N_16201,N_15699,N_15723);
nand U16202 (N_16202,N_15986,N_15982);
or U16203 (N_16203,N_15945,N_15604);
nand U16204 (N_16204,N_15827,N_15714);
or U16205 (N_16205,N_15548,N_15563);
xnor U16206 (N_16206,N_15525,N_15652);
xor U16207 (N_16207,N_15646,N_15643);
xnor U16208 (N_16208,N_15601,N_15629);
and U16209 (N_16209,N_15640,N_15911);
or U16210 (N_16210,N_15712,N_15614);
nand U16211 (N_16211,N_15802,N_15761);
nor U16212 (N_16212,N_15632,N_15772);
nor U16213 (N_16213,N_15595,N_15904);
xnor U16214 (N_16214,N_15603,N_15900);
and U16215 (N_16215,N_15885,N_15825);
nor U16216 (N_16216,N_15752,N_15689);
or U16217 (N_16217,N_15574,N_15660);
nor U16218 (N_16218,N_15711,N_15618);
xor U16219 (N_16219,N_15806,N_15826);
and U16220 (N_16220,N_15949,N_15649);
xor U16221 (N_16221,N_15709,N_15667);
or U16222 (N_16222,N_15857,N_15888);
or U16223 (N_16223,N_15899,N_15890);
xor U16224 (N_16224,N_15810,N_15519);
nor U16225 (N_16225,N_15600,N_15967);
and U16226 (N_16226,N_15999,N_15785);
and U16227 (N_16227,N_15773,N_15925);
and U16228 (N_16228,N_15591,N_15959);
and U16229 (N_16229,N_15589,N_15656);
or U16230 (N_16230,N_15790,N_15768);
xnor U16231 (N_16231,N_15528,N_15566);
nor U16232 (N_16232,N_15765,N_15957);
and U16233 (N_16233,N_15883,N_15950);
nand U16234 (N_16234,N_15943,N_15974);
or U16235 (N_16235,N_15710,N_15515);
nor U16236 (N_16236,N_15969,N_15955);
xnor U16237 (N_16237,N_15570,N_15700);
nor U16238 (N_16238,N_15560,N_15903);
or U16239 (N_16239,N_15740,N_15845);
nor U16240 (N_16240,N_15540,N_15744);
or U16241 (N_16241,N_15598,N_15796);
xnor U16242 (N_16242,N_15988,N_15870);
nand U16243 (N_16243,N_15533,N_15609);
or U16244 (N_16244,N_15839,N_15947);
nor U16245 (N_16245,N_15872,N_15928);
xnor U16246 (N_16246,N_15578,N_15715);
nor U16247 (N_16247,N_15972,N_15847);
and U16248 (N_16248,N_15690,N_15593);
or U16249 (N_16249,N_15599,N_15713);
or U16250 (N_16250,N_15980,N_15806);
xnor U16251 (N_16251,N_15690,N_15644);
nand U16252 (N_16252,N_15712,N_15576);
and U16253 (N_16253,N_15516,N_15802);
xor U16254 (N_16254,N_15512,N_15806);
nor U16255 (N_16255,N_15552,N_15647);
and U16256 (N_16256,N_15533,N_15564);
or U16257 (N_16257,N_15966,N_15658);
or U16258 (N_16258,N_15534,N_15527);
and U16259 (N_16259,N_15867,N_15851);
xnor U16260 (N_16260,N_15991,N_15509);
xnor U16261 (N_16261,N_15766,N_15732);
nand U16262 (N_16262,N_15531,N_15985);
or U16263 (N_16263,N_15649,N_15913);
nor U16264 (N_16264,N_15613,N_15998);
and U16265 (N_16265,N_15842,N_15746);
nand U16266 (N_16266,N_15882,N_15898);
and U16267 (N_16267,N_15942,N_15561);
or U16268 (N_16268,N_15641,N_15615);
nor U16269 (N_16269,N_15929,N_15834);
nor U16270 (N_16270,N_15700,N_15699);
xnor U16271 (N_16271,N_15947,N_15863);
nand U16272 (N_16272,N_15553,N_15696);
nand U16273 (N_16273,N_15940,N_15559);
or U16274 (N_16274,N_15584,N_15926);
nor U16275 (N_16275,N_15703,N_15837);
nor U16276 (N_16276,N_15555,N_15512);
nor U16277 (N_16277,N_15554,N_15925);
or U16278 (N_16278,N_15772,N_15860);
or U16279 (N_16279,N_15702,N_15892);
or U16280 (N_16280,N_15634,N_15560);
and U16281 (N_16281,N_15962,N_15579);
nand U16282 (N_16282,N_15608,N_15577);
xor U16283 (N_16283,N_15610,N_15857);
or U16284 (N_16284,N_15572,N_15936);
and U16285 (N_16285,N_15917,N_15544);
and U16286 (N_16286,N_15558,N_15940);
nor U16287 (N_16287,N_15798,N_15597);
nor U16288 (N_16288,N_15704,N_15836);
and U16289 (N_16289,N_15708,N_15892);
or U16290 (N_16290,N_15757,N_15781);
nand U16291 (N_16291,N_15987,N_15597);
nor U16292 (N_16292,N_15556,N_15512);
nand U16293 (N_16293,N_15526,N_15575);
or U16294 (N_16294,N_15737,N_15968);
and U16295 (N_16295,N_15718,N_15761);
or U16296 (N_16296,N_15956,N_15895);
or U16297 (N_16297,N_15922,N_15652);
nand U16298 (N_16298,N_15579,N_15593);
xnor U16299 (N_16299,N_15805,N_15696);
and U16300 (N_16300,N_15571,N_15607);
or U16301 (N_16301,N_15581,N_15915);
and U16302 (N_16302,N_15955,N_15838);
nand U16303 (N_16303,N_15736,N_15788);
or U16304 (N_16304,N_15865,N_15890);
xor U16305 (N_16305,N_15845,N_15603);
or U16306 (N_16306,N_15550,N_15607);
and U16307 (N_16307,N_15618,N_15825);
nor U16308 (N_16308,N_15706,N_15596);
nand U16309 (N_16309,N_15811,N_15625);
nor U16310 (N_16310,N_15893,N_15819);
or U16311 (N_16311,N_15991,N_15865);
nor U16312 (N_16312,N_15825,N_15522);
or U16313 (N_16313,N_15776,N_15623);
or U16314 (N_16314,N_15676,N_15855);
or U16315 (N_16315,N_15676,N_15656);
nor U16316 (N_16316,N_15797,N_15612);
nand U16317 (N_16317,N_15906,N_15970);
xor U16318 (N_16318,N_15598,N_15828);
xnor U16319 (N_16319,N_15828,N_15638);
and U16320 (N_16320,N_15702,N_15827);
xnor U16321 (N_16321,N_15529,N_15835);
or U16322 (N_16322,N_15712,N_15952);
and U16323 (N_16323,N_15526,N_15959);
or U16324 (N_16324,N_15872,N_15509);
xnor U16325 (N_16325,N_15963,N_15829);
nand U16326 (N_16326,N_15850,N_15596);
nand U16327 (N_16327,N_15898,N_15552);
nand U16328 (N_16328,N_15788,N_15924);
xnor U16329 (N_16329,N_15527,N_15894);
or U16330 (N_16330,N_15786,N_15789);
nand U16331 (N_16331,N_15734,N_15883);
nor U16332 (N_16332,N_15700,N_15840);
nand U16333 (N_16333,N_15639,N_15636);
and U16334 (N_16334,N_15858,N_15866);
nor U16335 (N_16335,N_15609,N_15972);
and U16336 (N_16336,N_15764,N_15571);
or U16337 (N_16337,N_15541,N_15815);
xnor U16338 (N_16338,N_15714,N_15707);
nor U16339 (N_16339,N_15677,N_15744);
nor U16340 (N_16340,N_15510,N_15656);
xnor U16341 (N_16341,N_15892,N_15864);
or U16342 (N_16342,N_15546,N_15543);
or U16343 (N_16343,N_15976,N_15865);
and U16344 (N_16344,N_15514,N_15715);
nor U16345 (N_16345,N_15970,N_15674);
or U16346 (N_16346,N_15574,N_15873);
nand U16347 (N_16347,N_15998,N_15626);
xor U16348 (N_16348,N_15942,N_15573);
or U16349 (N_16349,N_15940,N_15694);
nand U16350 (N_16350,N_15771,N_15502);
or U16351 (N_16351,N_15904,N_15827);
nor U16352 (N_16352,N_15629,N_15606);
xnor U16353 (N_16353,N_15524,N_15939);
nand U16354 (N_16354,N_15797,N_15853);
xnor U16355 (N_16355,N_15774,N_15558);
nor U16356 (N_16356,N_15870,N_15758);
xnor U16357 (N_16357,N_15866,N_15932);
nand U16358 (N_16358,N_15530,N_15507);
xnor U16359 (N_16359,N_15678,N_15946);
xnor U16360 (N_16360,N_15534,N_15971);
and U16361 (N_16361,N_15946,N_15814);
nor U16362 (N_16362,N_15972,N_15829);
nand U16363 (N_16363,N_15590,N_15856);
and U16364 (N_16364,N_15719,N_15623);
or U16365 (N_16365,N_15758,N_15920);
and U16366 (N_16366,N_15846,N_15587);
xnor U16367 (N_16367,N_15517,N_15582);
xnor U16368 (N_16368,N_15707,N_15758);
nor U16369 (N_16369,N_15872,N_15773);
and U16370 (N_16370,N_15726,N_15921);
and U16371 (N_16371,N_15787,N_15526);
nor U16372 (N_16372,N_15552,N_15685);
nor U16373 (N_16373,N_15731,N_15600);
nor U16374 (N_16374,N_15811,N_15500);
or U16375 (N_16375,N_15817,N_15922);
nand U16376 (N_16376,N_15599,N_15524);
and U16377 (N_16377,N_15611,N_15642);
or U16378 (N_16378,N_15716,N_15842);
nor U16379 (N_16379,N_15972,N_15983);
or U16380 (N_16380,N_15716,N_15719);
nand U16381 (N_16381,N_15577,N_15591);
or U16382 (N_16382,N_15610,N_15784);
nor U16383 (N_16383,N_15564,N_15617);
and U16384 (N_16384,N_15756,N_15880);
nand U16385 (N_16385,N_15675,N_15893);
and U16386 (N_16386,N_15697,N_15704);
xnor U16387 (N_16387,N_15852,N_15513);
nor U16388 (N_16388,N_15740,N_15971);
and U16389 (N_16389,N_15988,N_15972);
nor U16390 (N_16390,N_15975,N_15658);
nand U16391 (N_16391,N_15970,N_15859);
nand U16392 (N_16392,N_15739,N_15623);
xnor U16393 (N_16393,N_15733,N_15969);
nand U16394 (N_16394,N_15644,N_15927);
or U16395 (N_16395,N_15979,N_15980);
or U16396 (N_16396,N_15599,N_15831);
nand U16397 (N_16397,N_15767,N_15757);
and U16398 (N_16398,N_15754,N_15636);
nand U16399 (N_16399,N_15764,N_15572);
or U16400 (N_16400,N_15784,N_15792);
and U16401 (N_16401,N_15653,N_15570);
xor U16402 (N_16402,N_15826,N_15975);
and U16403 (N_16403,N_15965,N_15669);
and U16404 (N_16404,N_15520,N_15784);
nor U16405 (N_16405,N_15844,N_15624);
nand U16406 (N_16406,N_15922,N_15782);
xnor U16407 (N_16407,N_15789,N_15670);
xnor U16408 (N_16408,N_15882,N_15639);
and U16409 (N_16409,N_15880,N_15636);
xor U16410 (N_16410,N_15861,N_15631);
nand U16411 (N_16411,N_15625,N_15972);
or U16412 (N_16412,N_15557,N_15726);
and U16413 (N_16413,N_15577,N_15927);
nor U16414 (N_16414,N_15957,N_15833);
and U16415 (N_16415,N_15557,N_15875);
xor U16416 (N_16416,N_15563,N_15891);
nand U16417 (N_16417,N_15853,N_15951);
and U16418 (N_16418,N_15863,N_15697);
and U16419 (N_16419,N_15832,N_15519);
nand U16420 (N_16420,N_15566,N_15979);
nor U16421 (N_16421,N_15992,N_15567);
or U16422 (N_16422,N_15573,N_15519);
nand U16423 (N_16423,N_15871,N_15649);
or U16424 (N_16424,N_15854,N_15577);
nand U16425 (N_16425,N_15902,N_15713);
xor U16426 (N_16426,N_15823,N_15814);
nand U16427 (N_16427,N_15671,N_15792);
or U16428 (N_16428,N_15727,N_15598);
xnor U16429 (N_16429,N_15567,N_15841);
xor U16430 (N_16430,N_15826,N_15702);
xor U16431 (N_16431,N_15789,N_15825);
nand U16432 (N_16432,N_15554,N_15724);
nor U16433 (N_16433,N_15911,N_15575);
and U16434 (N_16434,N_15563,N_15935);
nor U16435 (N_16435,N_15861,N_15692);
xnor U16436 (N_16436,N_15695,N_15726);
or U16437 (N_16437,N_15917,N_15913);
and U16438 (N_16438,N_15873,N_15852);
nor U16439 (N_16439,N_15975,N_15733);
or U16440 (N_16440,N_15978,N_15983);
nand U16441 (N_16441,N_15701,N_15865);
nor U16442 (N_16442,N_15652,N_15722);
xor U16443 (N_16443,N_15805,N_15816);
xnor U16444 (N_16444,N_15550,N_15711);
nor U16445 (N_16445,N_15616,N_15786);
xnor U16446 (N_16446,N_15858,N_15698);
xor U16447 (N_16447,N_15632,N_15591);
or U16448 (N_16448,N_15856,N_15647);
nor U16449 (N_16449,N_15731,N_15946);
or U16450 (N_16450,N_15978,N_15946);
xnor U16451 (N_16451,N_15703,N_15653);
and U16452 (N_16452,N_15900,N_15631);
and U16453 (N_16453,N_15866,N_15887);
nand U16454 (N_16454,N_15890,N_15946);
xor U16455 (N_16455,N_15785,N_15932);
xnor U16456 (N_16456,N_15777,N_15802);
xor U16457 (N_16457,N_15941,N_15505);
nor U16458 (N_16458,N_15990,N_15960);
or U16459 (N_16459,N_15939,N_15699);
xor U16460 (N_16460,N_15840,N_15821);
nand U16461 (N_16461,N_15747,N_15701);
nand U16462 (N_16462,N_15654,N_15946);
nor U16463 (N_16463,N_15978,N_15573);
or U16464 (N_16464,N_15633,N_15990);
nor U16465 (N_16465,N_15984,N_15625);
xor U16466 (N_16466,N_15565,N_15866);
nand U16467 (N_16467,N_15971,N_15957);
nand U16468 (N_16468,N_15722,N_15606);
or U16469 (N_16469,N_15502,N_15505);
or U16470 (N_16470,N_15990,N_15930);
and U16471 (N_16471,N_15809,N_15661);
nor U16472 (N_16472,N_15709,N_15594);
nor U16473 (N_16473,N_15539,N_15626);
xnor U16474 (N_16474,N_15770,N_15986);
or U16475 (N_16475,N_15522,N_15543);
and U16476 (N_16476,N_15685,N_15667);
nor U16477 (N_16477,N_15831,N_15527);
xnor U16478 (N_16478,N_15534,N_15995);
xnor U16479 (N_16479,N_15780,N_15544);
nand U16480 (N_16480,N_15599,N_15815);
nand U16481 (N_16481,N_15827,N_15777);
nand U16482 (N_16482,N_15933,N_15598);
nor U16483 (N_16483,N_15743,N_15853);
nor U16484 (N_16484,N_15842,N_15875);
or U16485 (N_16485,N_15964,N_15523);
nor U16486 (N_16486,N_15506,N_15810);
nand U16487 (N_16487,N_15670,N_15604);
nand U16488 (N_16488,N_15557,N_15759);
nor U16489 (N_16489,N_15941,N_15916);
xor U16490 (N_16490,N_15738,N_15736);
and U16491 (N_16491,N_15926,N_15943);
nor U16492 (N_16492,N_15784,N_15671);
and U16493 (N_16493,N_15789,N_15869);
nand U16494 (N_16494,N_15645,N_15627);
or U16495 (N_16495,N_15668,N_15992);
and U16496 (N_16496,N_15695,N_15972);
nand U16497 (N_16497,N_15520,N_15649);
nor U16498 (N_16498,N_15511,N_15757);
xnor U16499 (N_16499,N_15636,N_15516);
xor U16500 (N_16500,N_16145,N_16315);
or U16501 (N_16501,N_16235,N_16057);
and U16502 (N_16502,N_16259,N_16285);
or U16503 (N_16503,N_16483,N_16308);
nor U16504 (N_16504,N_16365,N_16256);
or U16505 (N_16505,N_16381,N_16043);
nand U16506 (N_16506,N_16296,N_16229);
or U16507 (N_16507,N_16210,N_16112);
xnor U16508 (N_16508,N_16358,N_16261);
or U16509 (N_16509,N_16138,N_16175);
nand U16510 (N_16510,N_16083,N_16001);
xor U16511 (N_16511,N_16497,N_16306);
nand U16512 (N_16512,N_16300,N_16196);
and U16513 (N_16513,N_16238,N_16234);
nand U16514 (N_16514,N_16343,N_16474);
nand U16515 (N_16515,N_16061,N_16445);
nor U16516 (N_16516,N_16101,N_16137);
and U16517 (N_16517,N_16327,N_16218);
nor U16518 (N_16518,N_16357,N_16128);
nand U16519 (N_16519,N_16289,N_16363);
and U16520 (N_16520,N_16331,N_16035);
and U16521 (N_16521,N_16075,N_16416);
nor U16522 (N_16522,N_16286,N_16313);
nand U16523 (N_16523,N_16385,N_16265);
xnor U16524 (N_16524,N_16487,N_16183);
nand U16525 (N_16525,N_16338,N_16231);
and U16526 (N_16526,N_16236,N_16320);
xor U16527 (N_16527,N_16147,N_16168);
or U16528 (N_16528,N_16355,N_16018);
or U16529 (N_16529,N_16213,N_16202);
xnor U16530 (N_16530,N_16100,N_16014);
and U16531 (N_16531,N_16373,N_16311);
nand U16532 (N_16532,N_16444,N_16475);
or U16533 (N_16533,N_16485,N_16178);
or U16534 (N_16534,N_16378,N_16098);
and U16535 (N_16535,N_16245,N_16181);
nand U16536 (N_16536,N_16465,N_16203);
and U16537 (N_16537,N_16103,N_16070);
and U16538 (N_16538,N_16151,N_16194);
nand U16539 (N_16539,N_16033,N_16076);
xnor U16540 (N_16540,N_16339,N_16490);
or U16541 (N_16541,N_16477,N_16127);
xnor U16542 (N_16542,N_16433,N_16443);
xnor U16543 (N_16543,N_16163,N_16152);
and U16544 (N_16544,N_16116,N_16460);
or U16545 (N_16545,N_16251,N_16262);
xnor U16546 (N_16546,N_16362,N_16044);
xor U16547 (N_16547,N_16169,N_16491);
or U16548 (N_16548,N_16392,N_16117);
xor U16549 (N_16549,N_16106,N_16020);
xnor U16550 (N_16550,N_16185,N_16224);
xnor U16551 (N_16551,N_16370,N_16166);
and U16552 (N_16552,N_16063,N_16375);
nand U16553 (N_16553,N_16240,N_16431);
and U16554 (N_16554,N_16427,N_16393);
nand U16555 (N_16555,N_16060,N_16144);
nand U16556 (N_16556,N_16182,N_16412);
xnor U16557 (N_16557,N_16442,N_16454);
xnor U16558 (N_16558,N_16102,N_16160);
or U16559 (N_16559,N_16078,N_16471);
or U16560 (N_16560,N_16092,N_16071);
and U16561 (N_16561,N_16226,N_16028);
nand U16562 (N_16562,N_16420,N_16464);
xnor U16563 (N_16563,N_16439,N_16067);
xnor U16564 (N_16564,N_16223,N_16006);
or U16565 (N_16565,N_16013,N_16212);
nor U16566 (N_16566,N_16250,N_16222);
nor U16567 (N_16567,N_16409,N_16207);
and U16568 (N_16568,N_16039,N_16190);
and U16569 (N_16569,N_16255,N_16332);
xor U16570 (N_16570,N_16188,N_16453);
nor U16571 (N_16571,N_16211,N_16371);
or U16572 (N_16572,N_16022,N_16012);
or U16573 (N_16573,N_16323,N_16346);
nand U16574 (N_16574,N_16288,N_16488);
or U16575 (N_16575,N_16221,N_16027);
nand U16576 (N_16576,N_16056,N_16047);
nor U16577 (N_16577,N_16459,N_16026);
nor U16578 (N_16578,N_16037,N_16333);
and U16579 (N_16579,N_16199,N_16165);
xnor U16580 (N_16580,N_16372,N_16081);
xnor U16581 (N_16581,N_16398,N_16205);
and U16582 (N_16582,N_16390,N_16336);
nor U16583 (N_16583,N_16032,N_16282);
and U16584 (N_16584,N_16316,N_16239);
xor U16585 (N_16585,N_16177,N_16384);
nor U16586 (N_16586,N_16353,N_16271);
or U16587 (N_16587,N_16120,N_16426);
nor U16588 (N_16588,N_16318,N_16179);
or U16589 (N_16589,N_16146,N_16200);
or U16590 (N_16590,N_16085,N_16499);
and U16591 (N_16591,N_16024,N_16228);
nor U16592 (N_16592,N_16297,N_16309);
or U16593 (N_16593,N_16325,N_16480);
or U16594 (N_16594,N_16495,N_16298);
and U16595 (N_16595,N_16268,N_16023);
nand U16596 (N_16596,N_16302,N_16246);
xnor U16597 (N_16597,N_16415,N_16161);
and U16598 (N_16598,N_16432,N_16054);
nor U16599 (N_16599,N_16281,N_16304);
xnor U16600 (N_16600,N_16425,N_16414);
and U16601 (N_16601,N_16278,N_16424);
nand U16602 (N_16602,N_16277,N_16025);
nand U16603 (N_16603,N_16466,N_16258);
or U16604 (N_16604,N_16348,N_16312);
nor U16605 (N_16605,N_16118,N_16294);
or U16606 (N_16606,N_16328,N_16419);
xnor U16607 (N_16607,N_16260,N_16142);
nor U16608 (N_16608,N_16461,N_16321);
nor U16609 (N_16609,N_16301,N_16052);
or U16610 (N_16610,N_16051,N_16011);
or U16611 (N_16611,N_16383,N_16215);
or U16612 (N_16612,N_16064,N_16386);
nand U16613 (N_16613,N_16247,N_16208);
or U16614 (N_16614,N_16493,N_16233);
and U16615 (N_16615,N_16340,N_16449);
and U16616 (N_16616,N_16150,N_16330);
and U16617 (N_16617,N_16269,N_16379);
or U16618 (N_16618,N_16072,N_16481);
xnor U16619 (N_16619,N_16389,N_16482);
xnor U16620 (N_16620,N_16458,N_16069);
or U16621 (N_16621,N_16141,N_16124);
and U16622 (N_16622,N_16397,N_16295);
nand U16623 (N_16623,N_16374,N_16176);
nor U16624 (N_16624,N_16492,N_16053);
nor U16625 (N_16625,N_16391,N_16396);
xor U16626 (N_16626,N_16167,N_16337);
xor U16627 (N_16627,N_16248,N_16402);
nor U16628 (N_16628,N_16287,N_16430);
nand U16629 (N_16629,N_16496,N_16342);
or U16630 (N_16630,N_16280,N_16017);
nand U16631 (N_16631,N_16068,N_16084);
and U16632 (N_16632,N_16319,N_16180);
nand U16633 (N_16633,N_16048,N_16403);
or U16634 (N_16634,N_16317,N_16031);
or U16635 (N_16635,N_16010,N_16091);
or U16636 (N_16636,N_16154,N_16029);
nor U16637 (N_16637,N_16111,N_16354);
and U16638 (N_16638,N_16034,N_16015);
or U16639 (N_16639,N_16299,N_16105);
or U16640 (N_16640,N_16108,N_16476);
nand U16641 (N_16641,N_16195,N_16438);
and U16642 (N_16642,N_16356,N_16377);
or U16643 (N_16643,N_16401,N_16036);
or U16644 (N_16644,N_16095,N_16447);
xnor U16645 (N_16645,N_16267,N_16349);
nor U16646 (N_16646,N_16206,N_16109);
nand U16647 (N_16647,N_16382,N_16451);
nor U16648 (N_16648,N_16292,N_16156);
nand U16649 (N_16649,N_16115,N_16040);
nor U16650 (N_16650,N_16473,N_16408);
or U16651 (N_16651,N_16434,N_16204);
nor U16652 (N_16652,N_16273,N_16073);
xor U16653 (N_16653,N_16227,N_16411);
and U16654 (N_16654,N_16314,N_16489);
or U16655 (N_16655,N_16395,N_16388);
nand U16656 (N_16656,N_16284,N_16113);
nand U16657 (N_16657,N_16394,N_16359);
and U16658 (N_16658,N_16086,N_16237);
xnor U16659 (N_16659,N_16276,N_16254);
xnor U16660 (N_16660,N_16189,N_16122);
nor U16661 (N_16661,N_16217,N_16209);
nor U16662 (N_16662,N_16417,N_16042);
xnor U16663 (N_16663,N_16253,N_16066);
nand U16664 (N_16664,N_16136,N_16470);
nand U16665 (N_16665,N_16479,N_16159);
or U16666 (N_16666,N_16087,N_16279);
xor U16667 (N_16667,N_16041,N_16274);
xnor U16668 (N_16668,N_16399,N_16422);
or U16669 (N_16669,N_16158,N_16324);
or U16670 (N_16670,N_16360,N_16114);
or U16671 (N_16671,N_16155,N_16050);
nor U16672 (N_16672,N_16450,N_16405);
nand U16673 (N_16673,N_16005,N_16429);
nand U16674 (N_16674,N_16437,N_16310);
nand U16675 (N_16675,N_16074,N_16478);
or U16676 (N_16676,N_16457,N_16361);
and U16677 (N_16677,N_16404,N_16088);
nand U16678 (N_16678,N_16368,N_16019);
nand U16679 (N_16679,N_16406,N_16149);
or U16680 (N_16680,N_16139,N_16170);
xor U16681 (N_16681,N_16272,N_16003);
nand U16682 (N_16682,N_16187,N_16110);
nand U16683 (N_16683,N_16462,N_16134);
nand U16684 (N_16684,N_16376,N_16143);
or U16685 (N_16685,N_16077,N_16446);
or U16686 (N_16686,N_16004,N_16172);
and U16687 (N_16687,N_16219,N_16441);
nand U16688 (N_16688,N_16303,N_16249);
xnor U16689 (N_16689,N_16387,N_16232);
xor U16690 (N_16690,N_16225,N_16440);
nor U16691 (N_16691,N_16468,N_16484);
and U16692 (N_16692,N_16428,N_16242);
and U16693 (N_16693,N_16171,N_16096);
xor U16694 (N_16694,N_16448,N_16089);
and U16695 (N_16695,N_16038,N_16174);
or U16696 (N_16696,N_16059,N_16264);
nor U16697 (N_16697,N_16350,N_16090);
nor U16698 (N_16698,N_16494,N_16364);
xnor U16699 (N_16699,N_16198,N_16410);
nand U16700 (N_16700,N_16000,N_16099);
and U16701 (N_16701,N_16126,N_16119);
nand U16702 (N_16702,N_16079,N_16230);
nand U16703 (N_16703,N_16243,N_16472);
xor U16704 (N_16704,N_16162,N_16421);
and U16705 (N_16705,N_16293,N_16283);
nand U16706 (N_16706,N_16341,N_16007);
and U16707 (N_16707,N_16266,N_16030);
nand U16708 (N_16708,N_16148,N_16418);
or U16709 (N_16709,N_16352,N_16455);
or U16710 (N_16710,N_16322,N_16486);
nand U16711 (N_16711,N_16367,N_16125);
and U16712 (N_16712,N_16065,N_16400);
or U16713 (N_16713,N_16214,N_16351);
and U16714 (N_16714,N_16435,N_16080);
and U16715 (N_16715,N_16062,N_16345);
nand U16716 (N_16716,N_16244,N_16216);
nand U16717 (N_16717,N_16307,N_16407);
and U16718 (N_16718,N_16192,N_16157);
or U16719 (N_16719,N_16263,N_16423);
and U16720 (N_16720,N_16173,N_16498);
or U16721 (N_16721,N_16082,N_16413);
nand U16722 (N_16722,N_16369,N_16133);
nand U16723 (N_16723,N_16121,N_16049);
or U16724 (N_16724,N_16008,N_16193);
and U16725 (N_16725,N_16380,N_16002);
nor U16726 (N_16726,N_16009,N_16104);
and U16727 (N_16727,N_16366,N_16456);
and U16728 (N_16728,N_16436,N_16326);
or U16729 (N_16729,N_16290,N_16335);
nand U16730 (N_16730,N_16220,N_16463);
and U16731 (N_16731,N_16469,N_16184);
nand U16732 (N_16732,N_16270,N_16093);
nor U16733 (N_16733,N_16045,N_16135);
or U16734 (N_16734,N_16055,N_16123);
xnor U16735 (N_16735,N_16094,N_16329);
xor U16736 (N_16736,N_16046,N_16107);
or U16737 (N_16737,N_16058,N_16164);
or U16738 (N_16738,N_16467,N_16257);
and U16739 (N_16739,N_16201,N_16197);
or U16740 (N_16740,N_16241,N_16130);
xor U16741 (N_16741,N_16452,N_16131);
nand U16742 (N_16742,N_16291,N_16132);
nor U16743 (N_16743,N_16097,N_16016);
or U16744 (N_16744,N_16191,N_16140);
and U16745 (N_16745,N_16186,N_16252);
or U16746 (N_16746,N_16153,N_16334);
nor U16747 (N_16747,N_16129,N_16344);
and U16748 (N_16748,N_16305,N_16347);
xor U16749 (N_16749,N_16021,N_16275);
nand U16750 (N_16750,N_16067,N_16317);
nor U16751 (N_16751,N_16205,N_16461);
nand U16752 (N_16752,N_16475,N_16015);
nor U16753 (N_16753,N_16128,N_16078);
and U16754 (N_16754,N_16413,N_16340);
xor U16755 (N_16755,N_16171,N_16226);
or U16756 (N_16756,N_16064,N_16052);
xor U16757 (N_16757,N_16271,N_16087);
or U16758 (N_16758,N_16460,N_16270);
nor U16759 (N_16759,N_16104,N_16455);
xor U16760 (N_16760,N_16126,N_16319);
nor U16761 (N_16761,N_16496,N_16058);
nor U16762 (N_16762,N_16332,N_16059);
and U16763 (N_16763,N_16132,N_16370);
and U16764 (N_16764,N_16044,N_16423);
or U16765 (N_16765,N_16479,N_16253);
nand U16766 (N_16766,N_16281,N_16074);
nand U16767 (N_16767,N_16403,N_16073);
or U16768 (N_16768,N_16271,N_16418);
or U16769 (N_16769,N_16350,N_16460);
nand U16770 (N_16770,N_16138,N_16393);
and U16771 (N_16771,N_16096,N_16158);
and U16772 (N_16772,N_16155,N_16492);
xor U16773 (N_16773,N_16260,N_16254);
or U16774 (N_16774,N_16469,N_16248);
nor U16775 (N_16775,N_16405,N_16311);
nor U16776 (N_16776,N_16379,N_16451);
or U16777 (N_16777,N_16012,N_16312);
nand U16778 (N_16778,N_16407,N_16464);
nand U16779 (N_16779,N_16274,N_16089);
nand U16780 (N_16780,N_16057,N_16098);
or U16781 (N_16781,N_16217,N_16408);
or U16782 (N_16782,N_16466,N_16467);
and U16783 (N_16783,N_16458,N_16400);
xor U16784 (N_16784,N_16166,N_16297);
or U16785 (N_16785,N_16382,N_16413);
and U16786 (N_16786,N_16211,N_16414);
and U16787 (N_16787,N_16447,N_16231);
nand U16788 (N_16788,N_16402,N_16381);
or U16789 (N_16789,N_16286,N_16180);
nand U16790 (N_16790,N_16365,N_16425);
nand U16791 (N_16791,N_16482,N_16191);
nand U16792 (N_16792,N_16138,N_16090);
nor U16793 (N_16793,N_16147,N_16233);
or U16794 (N_16794,N_16177,N_16249);
and U16795 (N_16795,N_16103,N_16176);
nor U16796 (N_16796,N_16095,N_16242);
nand U16797 (N_16797,N_16292,N_16024);
nand U16798 (N_16798,N_16321,N_16464);
xnor U16799 (N_16799,N_16426,N_16143);
and U16800 (N_16800,N_16440,N_16385);
xor U16801 (N_16801,N_16336,N_16146);
nand U16802 (N_16802,N_16024,N_16493);
nand U16803 (N_16803,N_16001,N_16096);
and U16804 (N_16804,N_16069,N_16373);
xor U16805 (N_16805,N_16494,N_16086);
and U16806 (N_16806,N_16367,N_16429);
or U16807 (N_16807,N_16133,N_16053);
or U16808 (N_16808,N_16259,N_16144);
or U16809 (N_16809,N_16138,N_16024);
xnor U16810 (N_16810,N_16045,N_16127);
nor U16811 (N_16811,N_16109,N_16447);
or U16812 (N_16812,N_16493,N_16019);
nand U16813 (N_16813,N_16454,N_16419);
or U16814 (N_16814,N_16073,N_16318);
nand U16815 (N_16815,N_16111,N_16364);
or U16816 (N_16816,N_16047,N_16088);
and U16817 (N_16817,N_16180,N_16355);
or U16818 (N_16818,N_16187,N_16296);
or U16819 (N_16819,N_16213,N_16142);
nand U16820 (N_16820,N_16067,N_16165);
nand U16821 (N_16821,N_16434,N_16238);
xnor U16822 (N_16822,N_16126,N_16068);
xnor U16823 (N_16823,N_16051,N_16361);
xor U16824 (N_16824,N_16413,N_16132);
or U16825 (N_16825,N_16417,N_16139);
and U16826 (N_16826,N_16371,N_16075);
nor U16827 (N_16827,N_16105,N_16036);
or U16828 (N_16828,N_16442,N_16317);
and U16829 (N_16829,N_16320,N_16471);
and U16830 (N_16830,N_16100,N_16146);
and U16831 (N_16831,N_16348,N_16468);
xnor U16832 (N_16832,N_16205,N_16146);
xnor U16833 (N_16833,N_16437,N_16362);
xnor U16834 (N_16834,N_16303,N_16102);
nor U16835 (N_16835,N_16496,N_16138);
nor U16836 (N_16836,N_16180,N_16161);
or U16837 (N_16837,N_16317,N_16361);
and U16838 (N_16838,N_16069,N_16140);
and U16839 (N_16839,N_16086,N_16028);
xor U16840 (N_16840,N_16179,N_16378);
or U16841 (N_16841,N_16241,N_16290);
nand U16842 (N_16842,N_16124,N_16381);
nor U16843 (N_16843,N_16427,N_16125);
or U16844 (N_16844,N_16460,N_16131);
nor U16845 (N_16845,N_16333,N_16211);
nand U16846 (N_16846,N_16203,N_16091);
xnor U16847 (N_16847,N_16165,N_16351);
nor U16848 (N_16848,N_16416,N_16040);
and U16849 (N_16849,N_16133,N_16324);
nor U16850 (N_16850,N_16299,N_16040);
nor U16851 (N_16851,N_16043,N_16284);
and U16852 (N_16852,N_16114,N_16039);
nand U16853 (N_16853,N_16003,N_16078);
xor U16854 (N_16854,N_16196,N_16158);
nand U16855 (N_16855,N_16217,N_16437);
or U16856 (N_16856,N_16158,N_16142);
and U16857 (N_16857,N_16275,N_16339);
nor U16858 (N_16858,N_16369,N_16378);
nand U16859 (N_16859,N_16301,N_16251);
xor U16860 (N_16860,N_16127,N_16028);
and U16861 (N_16861,N_16124,N_16302);
and U16862 (N_16862,N_16464,N_16470);
nor U16863 (N_16863,N_16310,N_16036);
and U16864 (N_16864,N_16445,N_16008);
and U16865 (N_16865,N_16477,N_16372);
and U16866 (N_16866,N_16101,N_16197);
nand U16867 (N_16867,N_16053,N_16284);
xnor U16868 (N_16868,N_16107,N_16181);
xor U16869 (N_16869,N_16150,N_16174);
nand U16870 (N_16870,N_16191,N_16208);
nor U16871 (N_16871,N_16016,N_16256);
or U16872 (N_16872,N_16247,N_16246);
nor U16873 (N_16873,N_16113,N_16175);
and U16874 (N_16874,N_16430,N_16456);
nand U16875 (N_16875,N_16291,N_16063);
or U16876 (N_16876,N_16100,N_16445);
or U16877 (N_16877,N_16465,N_16479);
nand U16878 (N_16878,N_16411,N_16159);
nand U16879 (N_16879,N_16220,N_16384);
nand U16880 (N_16880,N_16220,N_16060);
and U16881 (N_16881,N_16081,N_16326);
nor U16882 (N_16882,N_16435,N_16318);
nand U16883 (N_16883,N_16395,N_16053);
xor U16884 (N_16884,N_16025,N_16457);
xor U16885 (N_16885,N_16177,N_16378);
or U16886 (N_16886,N_16114,N_16206);
xor U16887 (N_16887,N_16056,N_16220);
nor U16888 (N_16888,N_16109,N_16469);
nor U16889 (N_16889,N_16437,N_16337);
xnor U16890 (N_16890,N_16023,N_16266);
xor U16891 (N_16891,N_16190,N_16198);
xor U16892 (N_16892,N_16359,N_16349);
xor U16893 (N_16893,N_16203,N_16410);
nand U16894 (N_16894,N_16069,N_16452);
or U16895 (N_16895,N_16131,N_16497);
or U16896 (N_16896,N_16379,N_16033);
and U16897 (N_16897,N_16083,N_16023);
or U16898 (N_16898,N_16452,N_16097);
and U16899 (N_16899,N_16339,N_16297);
and U16900 (N_16900,N_16320,N_16188);
or U16901 (N_16901,N_16100,N_16127);
or U16902 (N_16902,N_16030,N_16360);
or U16903 (N_16903,N_16343,N_16459);
nor U16904 (N_16904,N_16209,N_16354);
and U16905 (N_16905,N_16220,N_16390);
xor U16906 (N_16906,N_16401,N_16082);
nand U16907 (N_16907,N_16194,N_16221);
nand U16908 (N_16908,N_16227,N_16118);
xor U16909 (N_16909,N_16222,N_16060);
and U16910 (N_16910,N_16287,N_16238);
nand U16911 (N_16911,N_16305,N_16434);
nor U16912 (N_16912,N_16167,N_16365);
or U16913 (N_16913,N_16355,N_16114);
xor U16914 (N_16914,N_16205,N_16286);
nor U16915 (N_16915,N_16108,N_16174);
or U16916 (N_16916,N_16347,N_16059);
nand U16917 (N_16917,N_16109,N_16159);
nor U16918 (N_16918,N_16067,N_16413);
nor U16919 (N_16919,N_16098,N_16240);
xor U16920 (N_16920,N_16313,N_16248);
xor U16921 (N_16921,N_16383,N_16223);
nand U16922 (N_16922,N_16390,N_16489);
and U16923 (N_16923,N_16499,N_16476);
nand U16924 (N_16924,N_16302,N_16204);
nand U16925 (N_16925,N_16268,N_16281);
nor U16926 (N_16926,N_16255,N_16278);
and U16927 (N_16927,N_16066,N_16009);
nand U16928 (N_16928,N_16427,N_16319);
nand U16929 (N_16929,N_16085,N_16043);
nand U16930 (N_16930,N_16016,N_16209);
xor U16931 (N_16931,N_16218,N_16472);
nor U16932 (N_16932,N_16143,N_16054);
xor U16933 (N_16933,N_16281,N_16297);
nor U16934 (N_16934,N_16069,N_16025);
nor U16935 (N_16935,N_16110,N_16103);
nor U16936 (N_16936,N_16157,N_16080);
xnor U16937 (N_16937,N_16371,N_16067);
xor U16938 (N_16938,N_16410,N_16262);
and U16939 (N_16939,N_16353,N_16482);
nor U16940 (N_16940,N_16462,N_16482);
nor U16941 (N_16941,N_16298,N_16283);
and U16942 (N_16942,N_16163,N_16467);
nor U16943 (N_16943,N_16157,N_16252);
xnor U16944 (N_16944,N_16334,N_16082);
nand U16945 (N_16945,N_16356,N_16480);
xor U16946 (N_16946,N_16497,N_16438);
nor U16947 (N_16947,N_16319,N_16098);
and U16948 (N_16948,N_16169,N_16417);
xor U16949 (N_16949,N_16046,N_16441);
nand U16950 (N_16950,N_16010,N_16461);
xnor U16951 (N_16951,N_16366,N_16045);
or U16952 (N_16952,N_16304,N_16193);
or U16953 (N_16953,N_16438,N_16336);
nand U16954 (N_16954,N_16008,N_16367);
or U16955 (N_16955,N_16424,N_16266);
nor U16956 (N_16956,N_16117,N_16077);
and U16957 (N_16957,N_16408,N_16053);
nor U16958 (N_16958,N_16267,N_16165);
xnor U16959 (N_16959,N_16146,N_16182);
nand U16960 (N_16960,N_16233,N_16210);
nand U16961 (N_16961,N_16069,N_16057);
or U16962 (N_16962,N_16460,N_16031);
nand U16963 (N_16963,N_16048,N_16023);
xnor U16964 (N_16964,N_16284,N_16148);
and U16965 (N_16965,N_16232,N_16383);
xor U16966 (N_16966,N_16101,N_16004);
nand U16967 (N_16967,N_16365,N_16026);
and U16968 (N_16968,N_16107,N_16367);
or U16969 (N_16969,N_16044,N_16136);
nand U16970 (N_16970,N_16109,N_16012);
nor U16971 (N_16971,N_16211,N_16434);
and U16972 (N_16972,N_16008,N_16473);
nor U16973 (N_16973,N_16461,N_16370);
xnor U16974 (N_16974,N_16381,N_16050);
nor U16975 (N_16975,N_16320,N_16178);
and U16976 (N_16976,N_16258,N_16349);
and U16977 (N_16977,N_16109,N_16132);
and U16978 (N_16978,N_16339,N_16218);
nand U16979 (N_16979,N_16438,N_16069);
nor U16980 (N_16980,N_16466,N_16005);
xnor U16981 (N_16981,N_16002,N_16042);
nor U16982 (N_16982,N_16349,N_16317);
nor U16983 (N_16983,N_16014,N_16317);
nand U16984 (N_16984,N_16177,N_16451);
or U16985 (N_16985,N_16359,N_16357);
nand U16986 (N_16986,N_16492,N_16266);
nand U16987 (N_16987,N_16198,N_16273);
and U16988 (N_16988,N_16383,N_16472);
xor U16989 (N_16989,N_16245,N_16354);
or U16990 (N_16990,N_16349,N_16050);
nand U16991 (N_16991,N_16132,N_16377);
nand U16992 (N_16992,N_16298,N_16496);
or U16993 (N_16993,N_16131,N_16070);
and U16994 (N_16994,N_16487,N_16326);
nand U16995 (N_16995,N_16076,N_16243);
nor U16996 (N_16996,N_16323,N_16008);
or U16997 (N_16997,N_16229,N_16446);
and U16998 (N_16998,N_16010,N_16007);
or U16999 (N_16999,N_16272,N_16300);
xor U17000 (N_17000,N_16934,N_16933);
nand U17001 (N_17001,N_16893,N_16729);
nor U17002 (N_17002,N_16593,N_16651);
or U17003 (N_17003,N_16615,N_16877);
nand U17004 (N_17004,N_16709,N_16944);
nor U17005 (N_17005,N_16853,N_16627);
or U17006 (N_17006,N_16866,N_16769);
and U17007 (N_17007,N_16661,N_16976);
or U17008 (N_17008,N_16561,N_16842);
nor U17009 (N_17009,N_16935,N_16808);
xor U17010 (N_17010,N_16584,N_16822);
or U17011 (N_17011,N_16927,N_16677);
xor U17012 (N_17012,N_16660,N_16872);
nor U17013 (N_17013,N_16868,N_16685);
and U17014 (N_17014,N_16666,N_16992);
nand U17015 (N_17015,N_16936,N_16713);
nand U17016 (N_17016,N_16977,N_16884);
nand U17017 (N_17017,N_16688,N_16676);
and U17018 (N_17018,N_16879,N_16840);
nor U17019 (N_17019,N_16728,N_16587);
xnor U17020 (N_17020,N_16532,N_16925);
and U17021 (N_17021,N_16781,N_16815);
nand U17022 (N_17022,N_16520,N_16556);
nor U17023 (N_17023,N_16574,N_16572);
nand U17024 (N_17024,N_16784,N_16723);
nor U17025 (N_17025,N_16550,N_16777);
nor U17026 (N_17026,N_16670,N_16653);
xor U17027 (N_17027,N_16617,N_16507);
and U17028 (N_17028,N_16748,N_16775);
nand U17029 (N_17029,N_16797,N_16898);
nand U17030 (N_17030,N_16869,N_16521);
xnor U17031 (N_17031,N_16938,N_16758);
and U17032 (N_17032,N_16715,N_16985);
or U17033 (N_17033,N_16900,N_16701);
xor U17034 (N_17034,N_16943,N_16503);
nor U17035 (N_17035,N_16500,N_16776);
nand U17036 (N_17036,N_16622,N_16778);
or U17037 (N_17037,N_16523,N_16553);
or U17038 (N_17038,N_16821,N_16870);
or U17039 (N_17039,N_16980,N_16964);
or U17040 (N_17040,N_16659,N_16923);
or U17041 (N_17041,N_16754,N_16696);
nand U17042 (N_17042,N_16512,N_16803);
or U17043 (N_17043,N_16832,N_16626);
nor U17044 (N_17044,N_16551,N_16562);
xor U17045 (N_17045,N_16811,N_16699);
nand U17046 (N_17046,N_16639,N_16989);
nor U17047 (N_17047,N_16759,N_16890);
nor U17048 (N_17048,N_16575,N_16929);
xor U17049 (N_17049,N_16823,N_16590);
and U17050 (N_17050,N_16851,N_16711);
or U17051 (N_17051,N_16644,N_16638);
and U17052 (N_17052,N_16692,N_16645);
and U17053 (N_17053,N_16524,N_16668);
or U17054 (N_17054,N_16613,N_16860);
xnor U17055 (N_17055,N_16721,N_16907);
xor U17056 (N_17056,N_16886,N_16541);
and U17057 (N_17057,N_16779,N_16588);
xnor U17058 (N_17058,N_16988,N_16513);
and U17059 (N_17059,N_16831,N_16979);
and U17060 (N_17060,N_16838,N_16554);
xor U17061 (N_17061,N_16675,N_16747);
xor U17062 (N_17062,N_16843,N_16634);
and U17063 (N_17063,N_16643,N_16571);
nand U17064 (N_17064,N_16874,N_16847);
xnor U17065 (N_17065,N_16941,N_16631);
xnor U17066 (N_17066,N_16540,N_16946);
nor U17067 (N_17067,N_16891,N_16586);
nor U17068 (N_17068,N_16609,N_16973);
xor U17069 (N_17069,N_16607,N_16739);
nor U17070 (N_17070,N_16705,N_16732);
xnor U17071 (N_17071,N_16928,N_16509);
xor U17072 (N_17072,N_16612,N_16919);
xor U17073 (N_17073,N_16700,N_16972);
nor U17074 (N_17074,N_16859,N_16885);
and U17075 (N_17075,N_16955,N_16640);
nand U17076 (N_17076,N_16516,N_16930);
xnor U17077 (N_17077,N_16506,N_16873);
xnor U17078 (N_17078,N_16818,N_16763);
nand U17079 (N_17079,N_16826,N_16816);
nand U17080 (N_17080,N_16642,N_16599);
and U17081 (N_17081,N_16570,N_16647);
nor U17082 (N_17082,N_16883,N_16616);
nand U17083 (N_17083,N_16620,N_16915);
or U17084 (N_17084,N_16585,N_16981);
nor U17085 (N_17085,N_16504,N_16792);
xor U17086 (N_17086,N_16549,N_16555);
xor U17087 (N_17087,N_16531,N_16880);
xnor U17088 (N_17088,N_16908,N_16809);
or U17089 (N_17089,N_16737,N_16761);
and U17090 (N_17090,N_16892,N_16529);
or U17091 (N_17091,N_16546,N_16750);
xor U17092 (N_17092,N_16602,N_16780);
xor U17093 (N_17093,N_16606,N_16583);
or U17094 (N_17094,N_16994,N_16578);
and U17095 (N_17095,N_16738,N_16846);
xor U17096 (N_17096,N_16845,N_16910);
nand U17097 (N_17097,N_16827,N_16543);
nor U17098 (N_17098,N_16694,N_16533);
and U17099 (N_17099,N_16905,N_16514);
nor U17100 (N_17100,N_16537,N_16863);
or U17101 (N_17101,N_16906,N_16970);
or U17102 (N_17102,N_16684,N_16760);
nor U17103 (N_17103,N_16962,N_16594);
nand U17104 (N_17104,N_16901,N_16918);
and U17105 (N_17105,N_16968,N_16913);
and U17106 (N_17106,N_16722,N_16530);
xnor U17107 (N_17107,N_16702,N_16741);
nor U17108 (N_17108,N_16600,N_16596);
xnor U17109 (N_17109,N_16878,N_16959);
nor U17110 (N_17110,N_16736,N_16791);
nand U17111 (N_17111,N_16745,N_16652);
and U17112 (N_17112,N_16681,N_16814);
nor U17113 (N_17113,N_16717,N_16689);
nor U17114 (N_17114,N_16757,N_16719);
nor U17115 (N_17115,N_16559,N_16577);
and U17116 (N_17116,N_16591,N_16558);
xor U17117 (N_17117,N_16857,N_16767);
or U17118 (N_17118,N_16753,N_16786);
nor U17119 (N_17119,N_16864,N_16508);
xor U17120 (N_17120,N_16637,N_16982);
and U17121 (N_17121,N_16614,N_16836);
or U17122 (N_17122,N_16686,N_16862);
and U17123 (N_17123,N_16665,N_16682);
xor U17124 (N_17124,N_16518,N_16904);
xor U17125 (N_17125,N_16691,N_16641);
xor U17126 (N_17126,N_16727,N_16894);
or U17127 (N_17127,N_16993,N_16855);
or U17128 (N_17128,N_16597,N_16733);
or U17129 (N_17129,N_16505,N_16770);
nor U17130 (N_17130,N_16807,N_16932);
or U17131 (N_17131,N_16751,N_16920);
or U17132 (N_17132,N_16517,N_16548);
and U17133 (N_17133,N_16744,N_16848);
xnor U17134 (N_17134,N_16630,N_16534);
or U17135 (N_17135,N_16695,N_16697);
nor U17136 (N_17136,N_16867,N_16755);
xor U17137 (N_17137,N_16710,N_16997);
nand U17138 (N_17138,N_16984,N_16511);
xor U17139 (N_17139,N_16954,N_16568);
xor U17140 (N_17140,N_16967,N_16895);
nand U17141 (N_17141,N_16693,N_16662);
xor U17142 (N_17142,N_16817,N_16714);
nand U17143 (N_17143,N_16734,N_16795);
or U17144 (N_17144,N_16844,N_16909);
nand U17145 (N_17145,N_16810,N_16731);
and U17146 (N_17146,N_16628,N_16706);
nand U17147 (N_17147,N_16765,N_16749);
or U17148 (N_17148,N_16704,N_16703);
nor U17149 (N_17149,N_16610,N_16636);
or U17150 (N_17150,N_16942,N_16538);
and U17151 (N_17151,N_16672,N_16772);
and U17152 (N_17152,N_16798,N_16592);
nor U17153 (N_17153,N_16820,N_16718);
nand U17154 (N_17154,N_16528,N_16812);
nand U17155 (N_17155,N_16806,N_16576);
xnor U17156 (N_17156,N_16899,N_16957);
nor U17157 (N_17157,N_16604,N_16945);
xor U17158 (N_17158,N_16996,N_16793);
and U17159 (N_17159,N_16589,N_16605);
nand U17160 (N_17160,N_16567,N_16849);
xnor U17161 (N_17161,N_16657,N_16563);
nor U17162 (N_17162,N_16850,N_16678);
nor U17163 (N_17163,N_16743,N_16830);
nand U17164 (N_17164,N_16952,N_16535);
and U17165 (N_17165,N_16951,N_16648);
nand U17166 (N_17166,N_16773,N_16888);
nand U17167 (N_17167,N_16544,N_16931);
and U17168 (N_17168,N_16834,N_16601);
or U17169 (N_17169,N_16825,N_16632);
and U17170 (N_17170,N_16624,N_16582);
xor U17171 (N_17171,N_16947,N_16712);
or U17172 (N_17172,N_16991,N_16673);
nand U17173 (N_17173,N_16725,N_16939);
nand U17174 (N_17174,N_16547,N_16565);
nor U17175 (N_17175,N_16545,N_16999);
or U17176 (N_17176,N_16986,N_16958);
nor U17177 (N_17177,N_16948,N_16740);
and U17178 (N_17178,N_16618,N_16841);
and U17179 (N_17179,N_16526,N_16771);
xnor U17180 (N_17180,N_16680,N_16861);
xnor U17181 (N_17181,N_16966,N_16813);
or U17182 (N_17182,N_16829,N_16802);
nand U17183 (N_17183,N_16995,N_16876);
nor U17184 (N_17184,N_16635,N_16510);
xnor U17185 (N_17185,N_16756,N_16730);
nor U17186 (N_17186,N_16698,N_16961);
nor U17187 (N_17187,N_16573,N_16949);
xor U17188 (N_17188,N_16683,N_16804);
nor U17189 (N_17189,N_16914,N_16839);
or U17190 (N_17190,N_16794,N_16819);
nor U17191 (N_17191,N_16724,N_16858);
or U17192 (N_17192,N_16542,N_16983);
xnor U17193 (N_17193,N_16735,N_16940);
or U17194 (N_17194,N_16619,N_16746);
nand U17195 (N_17195,N_16679,N_16824);
nor U17196 (N_17196,N_16950,N_16921);
xnor U17197 (N_17197,N_16865,N_16536);
or U17198 (N_17198,N_16965,N_16887);
and U17199 (N_17199,N_16953,N_16581);
xnor U17200 (N_17200,N_16766,N_16963);
nand U17201 (N_17201,N_16787,N_16937);
nor U17202 (N_17202,N_16911,N_16790);
xor U17203 (N_17203,N_16882,N_16805);
nand U17204 (N_17204,N_16990,N_16629);
and U17205 (N_17205,N_16595,N_16854);
or U17206 (N_17206,N_16716,N_16603);
nand U17207 (N_17207,N_16852,N_16902);
and U17208 (N_17208,N_16833,N_16598);
and U17209 (N_17209,N_16564,N_16881);
xor U17210 (N_17210,N_16871,N_16789);
or U17211 (N_17211,N_16956,N_16687);
xnor U17212 (N_17212,N_16916,N_16960);
xor U17213 (N_17213,N_16525,N_16522);
or U17214 (N_17214,N_16654,N_16742);
or U17215 (N_17215,N_16782,N_16608);
nor U17216 (N_17216,N_16922,N_16527);
or U17217 (N_17217,N_16690,N_16975);
and U17218 (N_17218,N_16667,N_16764);
nor U17219 (N_17219,N_16669,N_16978);
or U17220 (N_17220,N_16552,N_16835);
nor U17221 (N_17221,N_16912,N_16579);
and U17222 (N_17222,N_16774,N_16658);
nor U17223 (N_17223,N_16566,N_16971);
nand U17224 (N_17224,N_16663,N_16875);
or U17225 (N_17225,N_16674,N_16896);
or U17226 (N_17226,N_16664,N_16560);
nand U17227 (N_17227,N_16557,N_16569);
and U17228 (N_17228,N_16646,N_16987);
nand U17229 (N_17229,N_16924,N_16917);
nor U17230 (N_17230,N_16633,N_16720);
and U17231 (N_17231,N_16752,N_16519);
nand U17232 (N_17232,N_16799,N_16856);
nand U17233 (N_17233,N_16708,N_16897);
or U17234 (N_17234,N_16501,N_16800);
and U17235 (N_17235,N_16998,N_16649);
and U17236 (N_17236,N_16788,N_16889);
and U17237 (N_17237,N_16796,N_16926);
nor U17238 (N_17238,N_16580,N_16623);
nor U17239 (N_17239,N_16768,N_16783);
nor U17240 (N_17240,N_16625,N_16903);
nor U17241 (N_17241,N_16974,N_16671);
or U17242 (N_17242,N_16656,N_16650);
nor U17243 (N_17243,N_16539,N_16502);
nand U17244 (N_17244,N_16621,N_16611);
nand U17245 (N_17245,N_16515,N_16762);
xor U17246 (N_17246,N_16969,N_16655);
nor U17247 (N_17247,N_16828,N_16837);
nor U17248 (N_17248,N_16785,N_16801);
or U17249 (N_17249,N_16707,N_16726);
nor U17250 (N_17250,N_16586,N_16764);
nor U17251 (N_17251,N_16904,N_16708);
xor U17252 (N_17252,N_16925,N_16689);
xnor U17253 (N_17253,N_16890,N_16861);
and U17254 (N_17254,N_16795,N_16904);
or U17255 (N_17255,N_16815,N_16804);
nor U17256 (N_17256,N_16512,N_16625);
nand U17257 (N_17257,N_16936,N_16950);
nor U17258 (N_17258,N_16748,N_16791);
nor U17259 (N_17259,N_16793,N_16688);
and U17260 (N_17260,N_16535,N_16730);
nand U17261 (N_17261,N_16978,N_16886);
or U17262 (N_17262,N_16597,N_16870);
and U17263 (N_17263,N_16597,N_16988);
and U17264 (N_17264,N_16803,N_16722);
xnor U17265 (N_17265,N_16979,N_16929);
or U17266 (N_17266,N_16593,N_16560);
nand U17267 (N_17267,N_16721,N_16895);
nor U17268 (N_17268,N_16638,N_16919);
nand U17269 (N_17269,N_16937,N_16860);
or U17270 (N_17270,N_16717,N_16992);
and U17271 (N_17271,N_16608,N_16552);
or U17272 (N_17272,N_16704,N_16689);
and U17273 (N_17273,N_16815,N_16825);
xnor U17274 (N_17274,N_16653,N_16829);
or U17275 (N_17275,N_16762,N_16781);
nor U17276 (N_17276,N_16937,N_16975);
xnor U17277 (N_17277,N_16708,N_16870);
nor U17278 (N_17278,N_16913,N_16950);
nand U17279 (N_17279,N_16697,N_16853);
nor U17280 (N_17280,N_16949,N_16602);
xnor U17281 (N_17281,N_16513,N_16825);
nand U17282 (N_17282,N_16734,N_16815);
or U17283 (N_17283,N_16740,N_16949);
and U17284 (N_17284,N_16790,N_16978);
xnor U17285 (N_17285,N_16561,N_16803);
or U17286 (N_17286,N_16572,N_16557);
and U17287 (N_17287,N_16855,N_16599);
nand U17288 (N_17288,N_16950,N_16682);
nand U17289 (N_17289,N_16663,N_16890);
or U17290 (N_17290,N_16609,N_16848);
xnor U17291 (N_17291,N_16578,N_16896);
and U17292 (N_17292,N_16655,N_16621);
nand U17293 (N_17293,N_16946,N_16644);
and U17294 (N_17294,N_16614,N_16772);
nor U17295 (N_17295,N_16988,N_16539);
and U17296 (N_17296,N_16891,N_16720);
nand U17297 (N_17297,N_16716,N_16506);
nand U17298 (N_17298,N_16818,N_16838);
or U17299 (N_17299,N_16801,N_16744);
xor U17300 (N_17300,N_16942,N_16982);
and U17301 (N_17301,N_16936,N_16832);
xnor U17302 (N_17302,N_16949,N_16662);
nor U17303 (N_17303,N_16598,N_16677);
or U17304 (N_17304,N_16786,N_16717);
and U17305 (N_17305,N_16679,N_16608);
nor U17306 (N_17306,N_16862,N_16584);
xnor U17307 (N_17307,N_16809,N_16621);
nor U17308 (N_17308,N_16694,N_16713);
nor U17309 (N_17309,N_16865,N_16824);
xor U17310 (N_17310,N_16903,N_16987);
and U17311 (N_17311,N_16934,N_16999);
xor U17312 (N_17312,N_16917,N_16778);
or U17313 (N_17313,N_16527,N_16718);
xnor U17314 (N_17314,N_16812,N_16933);
xor U17315 (N_17315,N_16824,N_16966);
or U17316 (N_17316,N_16898,N_16824);
or U17317 (N_17317,N_16978,N_16821);
and U17318 (N_17318,N_16823,N_16677);
or U17319 (N_17319,N_16881,N_16804);
nand U17320 (N_17320,N_16627,N_16919);
xnor U17321 (N_17321,N_16565,N_16894);
nand U17322 (N_17322,N_16617,N_16977);
nor U17323 (N_17323,N_16516,N_16772);
nand U17324 (N_17324,N_16912,N_16974);
nor U17325 (N_17325,N_16634,N_16708);
nor U17326 (N_17326,N_16757,N_16892);
or U17327 (N_17327,N_16780,N_16677);
nand U17328 (N_17328,N_16709,N_16570);
nor U17329 (N_17329,N_16627,N_16773);
xnor U17330 (N_17330,N_16918,N_16855);
and U17331 (N_17331,N_16889,N_16771);
or U17332 (N_17332,N_16884,N_16969);
and U17333 (N_17333,N_16985,N_16853);
xor U17334 (N_17334,N_16762,N_16861);
xor U17335 (N_17335,N_16824,N_16626);
nor U17336 (N_17336,N_16693,N_16810);
nor U17337 (N_17337,N_16803,N_16887);
and U17338 (N_17338,N_16873,N_16813);
xor U17339 (N_17339,N_16922,N_16528);
nor U17340 (N_17340,N_16593,N_16707);
and U17341 (N_17341,N_16781,N_16623);
nor U17342 (N_17342,N_16756,N_16737);
xnor U17343 (N_17343,N_16573,N_16884);
xor U17344 (N_17344,N_16990,N_16832);
and U17345 (N_17345,N_16901,N_16729);
nand U17346 (N_17346,N_16965,N_16955);
nor U17347 (N_17347,N_16693,N_16738);
nand U17348 (N_17348,N_16645,N_16546);
and U17349 (N_17349,N_16624,N_16961);
xnor U17350 (N_17350,N_16972,N_16916);
and U17351 (N_17351,N_16917,N_16789);
xnor U17352 (N_17352,N_16914,N_16953);
xor U17353 (N_17353,N_16725,N_16750);
nand U17354 (N_17354,N_16518,N_16970);
nor U17355 (N_17355,N_16907,N_16943);
and U17356 (N_17356,N_16606,N_16623);
nand U17357 (N_17357,N_16734,N_16524);
xor U17358 (N_17358,N_16619,N_16830);
nand U17359 (N_17359,N_16721,N_16711);
nor U17360 (N_17360,N_16762,N_16621);
and U17361 (N_17361,N_16779,N_16998);
nand U17362 (N_17362,N_16516,N_16627);
and U17363 (N_17363,N_16637,N_16786);
nor U17364 (N_17364,N_16504,N_16697);
nand U17365 (N_17365,N_16634,N_16893);
nand U17366 (N_17366,N_16825,N_16921);
nand U17367 (N_17367,N_16790,N_16759);
nand U17368 (N_17368,N_16534,N_16831);
or U17369 (N_17369,N_16756,N_16800);
and U17370 (N_17370,N_16834,N_16534);
and U17371 (N_17371,N_16788,N_16830);
nand U17372 (N_17372,N_16913,N_16694);
nand U17373 (N_17373,N_16893,N_16504);
nor U17374 (N_17374,N_16852,N_16502);
nand U17375 (N_17375,N_16587,N_16520);
nand U17376 (N_17376,N_16731,N_16943);
nor U17377 (N_17377,N_16845,N_16514);
xor U17378 (N_17378,N_16976,N_16635);
and U17379 (N_17379,N_16852,N_16998);
or U17380 (N_17380,N_16525,N_16788);
nand U17381 (N_17381,N_16686,N_16524);
and U17382 (N_17382,N_16606,N_16819);
and U17383 (N_17383,N_16616,N_16571);
xor U17384 (N_17384,N_16500,N_16515);
and U17385 (N_17385,N_16946,N_16610);
or U17386 (N_17386,N_16563,N_16709);
xor U17387 (N_17387,N_16855,N_16771);
nor U17388 (N_17388,N_16715,N_16558);
and U17389 (N_17389,N_16844,N_16940);
nor U17390 (N_17390,N_16538,N_16661);
nand U17391 (N_17391,N_16712,N_16614);
or U17392 (N_17392,N_16555,N_16930);
nor U17393 (N_17393,N_16664,N_16976);
nand U17394 (N_17394,N_16760,N_16895);
nor U17395 (N_17395,N_16725,N_16608);
nand U17396 (N_17396,N_16612,N_16722);
or U17397 (N_17397,N_16877,N_16554);
nor U17398 (N_17398,N_16629,N_16529);
or U17399 (N_17399,N_16699,N_16512);
or U17400 (N_17400,N_16869,N_16754);
and U17401 (N_17401,N_16701,N_16991);
nand U17402 (N_17402,N_16973,N_16693);
nand U17403 (N_17403,N_16911,N_16983);
xnor U17404 (N_17404,N_16759,N_16996);
xor U17405 (N_17405,N_16573,N_16601);
xor U17406 (N_17406,N_16597,N_16945);
or U17407 (N_17407,N_16919,N_16587);
nand U17408 (N_17408,N_16714,N_16921);
xnor U17409 (N_17409,N_16885,N_16567);
and U17410 (N_17410,N_16908,N_16647);
nor U17411 (N_17411,N_16850,N_16556);
nand U17412 (N_17412,N_16668,N_16734);
xnor U17413 (N_17413,N_16611,N_16845);
and U17414 (N_17414,N_16938,N_16881);
or U17415 (N_17415,N_16553,N_16709);
xor U17416 (N_17416,N_16788,N_16699);
and U17417 (N_17417,N_16912,N_16743);
and U17418 (N_17418,N_16789,N_16902);
nor U17419 (N_17419,N_16699,N_16960);
xor U17420 (N_17420,N_16993,N_16652);
and U17421 (N_17421,N_16730,N_16512);
nand U17422 (N_17422,N_16977,N_16788);
xor U17423 (N_17423,N_16930,N_16651);
or U17424 (N_17424,N_16511,N_16769);
and U17425 (N_17425,N_16995,N_16689);
and U17426 (N_17426,N_16801,N_16773);
and U17427 (N_17427,N_16796,N_16951);
and U17428 (N_17428,N_16659,N_16916);
and U17429 (N_17429,N_16712,N_16804);
nor U17430 (N_17430,N_16792,N_16798);
xor U17431 (N_17431,N_16734,N_16519);
nand U17432 (N_17432,N_16714,N_16749);
nand U17433 (N_17433,N_16573,N_16635);
and U17434 (N_17434,N_16635,N_16747);
or U17435 (N_17435,N_16824,N_16831);
or U17436 (N_17436,N_16652,N_16538);
and U17437 (N_17437,N_16519,N_16599);
xnor U17438 (N_17438,N_16849,N_16761);
nor U17439 (N_17439,N_16780,N_16651);
or U17440 (N_17440,N_16721,N_16627);
nand U17441 (N_17441,N_16799,N_16752);
and U17442 (N_17442,N_16990,N_16939);
nor U17443 (N_17443,N_16680,N_16679);
nor U17444 (N_17444,N_16778,N_16504);
or U17445 (N_17445,N_16608,N_16558);
and U17446 (N_17446,N_16845,N_16527);
or U17447 (N_17447,N_16545,N_16852);
and U17448 (N_17448,N_16913,N_16533);
nand U17449 (N_17449,N_16654,N_16570);
or U17450 (N_17450,N_16589,N_16619);
xor U17451 (N_17451,N_16542,N_16520);
or U17452 (N_17452,N_16824,N_16691);
nand U17453 (N_17453,N_16728,N_16708);
nor U17454 (N_17454,N_16952,N_16553);
xor U17455 (N_17455,N_16584,N_16952);
and U17456 (N_17456,N_16691,N_16639);
nand U17457 (N_17457,N_16794,N_16987);
nand U17458 (N_17458,N_16722,N_16729);
nand U17459 (N_17459,N_16795,N_16577);
nor U17460 (N_17460,N_16810,N_16803);
nor U17461 (N_17461,N_16987,N_16532);
and U17462 (N_17462,N_16875,N_16706);
nor U17463 (N_17463,N_16553,N_16802);
xnor U17464 (N_17464,N_16849,N_16814);
and U17465 (N_17465,N_16541,N_16533);
or U17466 (N_17466,N_16550,N_16865);
nor U17467 (N_17467,N_16763,N_16912);
or U17468 (N_17468,N_16871,N_16957);
or U17469 (N_17469,N_16630,N_16575);
xor U17470 (N_17470,N_16701,N_16725);
and U17471 (N_17471,N_16921,N_16717);
xnor U17472 (N_17472,N_16567,N_16992);
nand U17473 (N_17473,N_16566,N_16705);
xnor U17474 (N_17474,N_16579,N_16932);
xor U17475 (N_17475,N_16722,N_16558);
and U17476 (N_17476,N_16739,N_16748);
nor U17477 (N_17477,N_16634,N_16560);
xor U17478 (N_17478,N_16520,N_16582);
xnor U17479 (N_17479,N_16708,N_16594);
or U17480 (N_17480,N_16654,N_16996);
or U17481 (N_17481,N_16699,N_16563);
nor U17482 (N_17482,N_16738,N_16783);
nor U17483 (N_17483,N_16840,N_16708);
nor U17484 (N_17484,N_16657,N_16854);
nor U17485 (N_17485,N_16542,N_16527);
and U17486 (N_17486,N_16786,N_16613);
nand U17487 (N_17487,N_16516,N_16957);
nor U17488 (N_17488,N_16695,N_16839);
nand U17489 (N_17489,N_16818,N_16613);
and U17490 (N_17490,N_16738,N_16986);
nor U17491 (N_17491,N_16516,N_16555);
nor U17492 (N_17492,N_16580,N_16864);
or U17493 (N_17493,N_16549,N_16673);
and U17494 (N_17494,N_16545,N_16610);
nor U17495 (N_17495,N_16737,N_16577);
nor U17496 (N_17496,N_16837,N_16859);
or U17497 (N_17497,N_16903,N_16506);
and U17498 (N_17498,N_16887,N_16643);
nand U17499 (N_17499,N_16617,N_16651);
and U17500 (N_17500,N_17356,N_17099);
or U17501 (N_17501,N_17471,N_17262);
nand U17502 (N_17502,N_17268,N_17265);
nand U17503 (N_17503,N_17093,N_17428);
nand U17504 (N_17504,N_17088,N_17073);
xor U17505 (N_17505,N_17245,N_17174);
xnor U17506 (N_17506,N_17000,N_17486);
nand U17507 (N_17507,N_17059,N_17061);
nor U17508 (N_17508,N_17327,N_17082);
nor U17509 (N_17509,N_17032,N_17341);
or U17510 (N_17510,N_17065,N_17201);
or U17511 (N_17511,N_17170,N_17117);
xor U17512 (N_17512,N_17068,N_17041);
or U17513 (N_17513,N_17326,N_17134);
nand U17514 (N_17514,N_17028,N_17141);
and U17515 (N_17515,N_17179,N_17296);
or U17516 (N_17516,N_17148,N_17317);
xor U17517 (N_17517,N_17476,N_17285);
nor U17518 (N_17518,N_17136,N_17217);
and U17519 (N_17519,N_17015,N_17302);
nor U17520 (N_17520,N_17127,N_17399);
and U17521 (N_17521,N_17490,N_17482);
nand U17522 (N_17522,N_17376,N_17043);
xor U17523 (N_17523,N_17485,N_17350);
and U17524 (N_17524,N_17018,N_17135);
xnor U17525 (N_17525,N_17044,N_17091);
nor U17526 (N_17526,N_17299,N_17131);
nor U17527 (N_17527,N_17488,N_17063);
and U17528 (N_17528,N_17125,N_17241);
and U17529 (N_17529,N_17142,N_17126);
nor U17530 (N_17530,N_17338,N_17054);
or U17531 (N_17531,N_17042,N_17367);
and U17532 (N_17532,N_17449,N_17260);
or U17533 (N_17533,N_17240,N_17055);
nor U17534 (N_17534,N_17416,N_17069);
and U17535 (N_17535,N_17047,N_17422);
nor U17536 (N_17536,N_17297,N_17253);
nor U17537 (N_17537,N_17194,N_17329);
or U17538 (N_17538,N_17316,N_17491);
nor U17539 (N_17539,N_17120,N_17357);
or U17540 (N_17540,N_17288,N_17076);
or U17541 (N_17541,N_17244,N_17252);
and U17542 (N_17542,N_17344,N_17430);
nand U17543 (N_17543,N_17331,N_17007);
nand U17544 (N_17544,N_17366,N_17480);
xnor U17545 (N_17545,N_17365,N_17492);
nor U17546 (N_17546,N_17242,N_17175);
xor U17547 (N_17547,N_17300,N_17128);
xnor U17548 (N_17548,N_17332,N_17005);
nor U17549 (N_17549,N_17226,N_17154);
or U17550 (N_17550,N_17308,N_17204);
xor U17551 (N_17551,N_17418,N_17410);
and U17552 (N_17552,N_17133,N_17320);
nor U17553 (N_17553,N_17411,N_17023);
nand U17554 (N_17554,N_17130,N_17465);
or U17555 (N_17555,N_17423,N_17340);
nor U17556 (N_17556,N_17248,N_17377);
nand U17557 (N_17557,N_17261,N_17477);
nand U17558 (N_17558,N_17186,N_17178);
nor U17559 (N_17559,N_17163,N_17314);
nor U17560 (N_17560,N_17239,N_17284);
nand U17561 (N_17561,N_17461,N_17029);
nand U17562 (N_17562,N_17474,N_17279);
and U17563 (N_17563,N_17305,N_17336);
nor U17564 (N_17564,N_17192,N_17439);
nand U17565 (N_17565,N_17092,N_17315);
or U17566 (N_17566,N_17074,N_17427);
or U17567 (N_17567,N_17034,N_17359);
nand U17568 (N_17568,N_17420,N_17400);
and U17569 (N_17569,N_17026,N_17387);
and U17570 (N_17570,N_17251,N_17049);
and U17571 (N_17571,N_17100,N_17149);
nor U17572 (N_17572,N_17066,N_17493);
xnor U17573 (N_17573,N_17460,N_17182);
and U17574 (N_17574,N_17275,N_17045);
nand U17575 (N_17575,N_17421,N_17335);
xor U17576 (N_17576,N_17382,N_17196);
and U17577 (N_17577,N_17095,N_17379);
or U17578 (N_17578,N_17013,N_17072);
nand U17579 (N_17579,N_17447,N_17020);
and U17580 (N_17580,N_17216,N_17152);
xor U17581 (N_17581,N_17184,N_17349);
and U17582 (N_17582,N_17323,N_17115);
nor U17583 (N_17583,N_17090,N_17052);
xor U17584 (N_17584,N_17027,N_17236);
nor U17585 (N_17585,N_17031,N_17304);
xnor U17586 (N_17586,N_17348,N_17098);
or U17587 (N_17587,N_17259,N_17443);
or U17588 (N_17588,N_17437,N_17232);
and U17589 (N_17589,N_17272,N_17002);
nor U17590 (N_17590,N_17203,N_17106);
xnor U17591 (N_17591,N_17499,N_17140);
nand U17592 (N_17592,N_17156,N_17413);
nand U17593 (N_17593,N_17190,N_17124);
nor U17594 (N_17594,N_17173,N_17187);
or U17595 (N_17595,N_17455,N_17132);
xor U17596 (N_17596,N_17224,N_17024);
xor U17597 (N_17597,N_17278,N_17456);
or U17598 (N_17598,N_17303,N_17330);
nor U17599 (N_17599,N_17385,N_17064);
xnor U17600 (N_17600,N_17398,N_17159);
nand U17601 (N_17601,N_17221,N_17138);
nand U17602 (N_17602,N_17038,N_17151);
nor U17603 (N_17603,N_17352,N_17109);
xnor U17604 (N_17604,N_17466,N_17172);
xor U17605 (N_17605,N_17424,N_17371);
nand U17606 (N_17606,N_17351,N_17155);
and U17607 (N_17607,N_17249,N_17322);
nand U17608 (N_17608,N_17393,N_17150);
nor U17609 (N_17609,N_17033,N_17019);
and U17610 (N_17610,N_17458,N_17408);
nor U17611 (N_17611,N_17429,N_17078);
and U17612 (N_17612,N_17210,N_17145);
nand U17613 (N_17613,N_17062,N_17267);
nand U17614 (N_17614,N_17266,N_17467);
xor U17615 (N_17615,N_17280,N_17016);
xor U17616 (N_17616,N_17185,N_17358);
nand U17617 (N_17617,N_17484,N_17030);
or U17618 (N_17618,N_17328,N_17269);
nand U17619 (N_17619,N_17318,N_17257);
and U17620 (N_17620,N_17227,N_17215);
xor U17621 (N_17621,N_17058,N_17395);
nand U17622 (N_17622,N_17089,N_17081);
nand U17623 (N_17623,N_17487,N_17139);
and U17624 (N_17624,N_17289,N_17293);
xor U17625 (N_17625,N_17111,N_17229);
and U17626 (N_17626,N_17080,N_17071);
xor U17627 (N_17627,N_17198,N_17085);
and U17628 (N_17628,N_17067,N_17056);
and U17629 (N_17629,N_17189,N_17405);
nand U17630 (N_17630,N_17219,N_17223);
or U17631 (N_17631,N_17372,N_17258);
and U17632 (N_17632,N_17457,N_17087);
and U17633 (N_17633,N_17495,N_17220);
nand U17634 (N_17634,N_17050,N_17380);
nand U17635 (N_17635,N_17277,N_17401);
and U17636 (N_17636,N_17337,N_17364);
nand U17637 (N_17637,N_17419,N_17397);
nor U17638 (N_17638,N_17452,N_17137);
and U17639 (N_17639,N_17426,N_17103);
nand U17640 (N_17640,N_17473,N_17402);
or U17641 (N_17641,N_17209,N_17346);
xnor U17642 (N_17642,N_17247,N_17008);
and U17643 (N_17643,N_17324,N_17414);
and U17644 (N_17644,N_17006,N_17406);
nand U17645 (N_17645,N_17070,N_17368);
and U17646 (N_17646,N_17121,N_17205);
or U17647 (N_17647,N_17213,N_17407);
nand U17648 (N_17648,N_17048,N_17388);
or U17649 (N_17649,N_17483,N_17037);
xor U17650 (N_17650,N_17214,N_17325);
or U17651 (N_17651,N_17361,N_17309);
nand U17652 (N_17652,N_17004,N_17113);
nand U17653 (N_17653,N_17207,N_17310);
nand U17654 (N_17654,N_17475,N_17355);
nand U17655 (N_17655,N_17176,N_17146);
nand U17656 (N_17656,N_17237,N_17234);
xnor U17657 (N_17657,N_17129,N_17231);
nor U17658 (N_17658,N_17193,N_17206);
nand U17659 (N_17659,N_17157,N_17147);
nand U17660 (N_17660,N_17464,N_17225);
xor U17661 (N_17661,N_17311,N_17290);
and U17662 (N_17662,N_17208,N_17010);
and U17663 (N_17663,N_17021,N_17191);
nor U17664 (N_17664,N_17102,N_17084);
or U17665 (N_17665,N_17250,N_17270);
xor U17666 (N_17666,N_17412,N_17025);
nand U17667 (N_17667,N_17255,N_17306);
nor U17668 (N_17668,N_17230,N_17169);
and U17669 (N_17669,N_17212,N_17286);
and U17670 (N_17670,N_17403,N_17183);
xnor U17671 (N_17671,N_17321,N_17431);
xnor U17672 (N_17672,N_17307,N_17039);
and U17673 (N_17673,N_17360,N_17294);
nor U17674 (N_17674,N_17478,N_17362);
and U17675 (N_17675,N_17375,N_17389);
and U17676 (N_17676,N_17391,N_17075);
xor U17677 (N_17677,N_17101,N_17404);
or U17678 (N_17678,N_17470,N_17451);
xor U17679 (N_17679,N_17392,N_17112);
nor U17680 (N_17680,N_17009,N_17435);
nor U17681 (N_17681,N_17003,N_17425);
and U17682 (N_17682,N_17445,N_17394);
or U17683 (N_17683,N_17011,N_17434);
and U17684 (N_17684,N_17166,N_17256);
and U17685 (N_17685,N_17343,N_17243);
nand U17686 (N_17686,N_17313,N_17086);
and U17687 (N_17687,N_17441,N_17162);
and U17688 (N_17688,N_17040,N_17276);
xnor U17689 (N_17689,N_17195,N_17433);
xnor U17690 (N_17690,N_17295,N_17264);
or U17691 (N_17691,N_17188,N_17180);
and U17692 (N_17692,N_17334,N_17060);
nand U17693 (N_17693,N_17444,N_17468);
xnor U17694 (N_17694,N_17238,N_17096);
nand U17695 (N_17695,N_17202,N_17373);
xor U17696 (N_17696,N_17218,N_17228);
nor U17697 (N_17697,N_17051,N_17012);
nor U17698 (N_17698,N_17415,N_17200);
and U17699 (N_17699,N_17469,N_17354);
nand U17700 (N_17700,N_17353,N_17287);
nand U17701 (N_17701,N_17118,N_17254);
nor U17702 (N_17702,N_17235,N_17035);
or U17703 (N_17703,N_17298,N_17097);
xnor U17704 (N_17704,N_17263,N_17440);
and U17705 (N_17705,N_17446,N_17384);
or U17706 (N_17706,N_17442,N_17436);
and U17707 (N_17707,N_17274,N_17312);
or U17708 (N_17708,N_17378,N_17481);
nand U17709 (N_17709,N_17083,N_17417);
xnor U17710 (N_17710,N_17158,N_17496);
nand U17711 (N_17711,N_17161,N_17104);
nor U17712 (N_17712,N_17114,N_17022);
or U17713 (N_17713,N_17199,N_17119);
nand U17714 (N_17714,N_17438,N_17036);
or U17715 (N_17715,N_17246,N_17222);
nor U17716 (N_17716,N_17453,N_17291);
or U17717 (N_17717,N_17181,N_17472);
nand U17718 (N_17718,N_17396,N_17374);
nand U17719 (N_17719,N_17001,N_17165);
nand U17720 (N_17720,N_17177,N_17370);
nand U17721 (N_17721,N_17171,N_17057);
xnor U17722 (N_17722,N_17211,N_17116);
nor U17723 (N_17723,N_17462,N_17342);
and U17724 (N_17724,N_17369,N_17463);
nor U17725 (N_17725,N_17164,N_17292);
or U17726 (N_17726,N_17108,N_17077);
or U17727 (N_17727,N_17110,N_17273);
nand U17728 (N_17728,N_17143,N_17107);
nand U17729 (N_17729,N_17123,N_17459);
or U17730 (N_17730,N_17301,N_17319);
xor U17731 (N_17731,N_17390,N_17333);
nor U17732 (N_17732,N_17168,N_17383);
or U17733 (N_17733,N_17498,N_17105);
xnor U17734 (N_17734,N_17448,N_17432);
nor U17735 (N_17735,N_17497,N_17079);
or U17736 (N_17736,N_17153,N_17014);
and U17737 (N_17737,N_17494,N_17386);
nand U17738 (N_17738,N_17283,N_17167);
xor U17739 (N_17739,N_17094,N_17454);
or U17740 (N_17740,N_17339,N_17450);
xnor U17741 (N_17741,N_17233,N_17345);
and U17742 (N_17742,N_17347,N_17046);
xnor U17743 (N_17743,N_17271,N_17479);
or U17744 (N_17744,N_17122,N_17381);
nor U17745 (N_17745,N_17197,N_17281);
xnor U17746 (N_17746,N_17144,N_17282);
nor U17747 (N_17747,N_17409,N_17053);
xnor U17748 (N_17748,N_17017,N_17489);
nor U17749 (N_17749,N_17363,N_17160);
and U17750 (N_17750,N_17191,N_17114);
nor U17751 (N_17751,N_17353,N_17309);
and U17752 (N_17752,N_17202,N_17342);
or U17753 (N_17753,N_17437,N_17480);
nand U17754 (N_17754,N_17103,N_17006);
or U17755 (N_17755,N_17042,N_17145);
xor U17756 (N_17756,N_17321,N_17390);
and U17757 (N_17757,N_17262,N_17480);
nor U17758 (N_17758,N_17071,N_17242);
or U17759 (N_17759,N_17300,N_17112);
nor U17760 (N_17760,N_17289,N_17283);
xor U17761 (N_17761,N_17241,N_17482);
nand U17762 (N_17762,N_17023,N_17187);
nand U17763 (N_17763,N_17175,N_17270);
nand U17764 (N_17764,N_17121,N_17198);
nor U17765 (N_17765,N_17048,N_17489);
and U17766 (N_17766,N_17086,N_17219);
xnor U17767 (N_17767,N_17452,N_17223);
nand U17768 (N_17768,N_17206,N_17414);
and U17769 (N_17769,N_17109,N_17247);
nand U17770 (N_17770,N_17173,N_17087);
or U17771 (N_17771,N_17029,N_17275);
xor U17772 (N_17772,N_17114,N_17495);
xor U17773 (N_17773,N_17169,N_17458);
or U17774 (N_17774,N_17056,N_17017);
xnor U17775 (N_17775,N_17066,N_17327);
or U17776 (N_17776,N_17324,N_17435);
nor U17777 (N_17777,N_17221,N_17282);
nand U17778 (N_17778,N_17398,N_17219);
or U17779 (N_17779,N_17054,N_17017);
and U17780 (N_17780,N_17272,N_17053);
nand U17781 (N_17781,N_17018,N_17391);
xnor U17782 (N_17782,N_17259,N_17334);
or U17783 (N_17783,N_17330,N_17257);
and U17784 (N_17784,N_17394,N_17405);
nor U17785 (N_17785,N_17413,N_17143);
nor U17786 (N_17786,N_17010,N_17017);
nand U17787 (N_17787,N_17310,N_17103);
or U17788 (N_17788,N_17212,N_17348);
and U17789 (N_17789,N_17478,N_17140);
and U17790 (N_17790,N_17410,N_17478);
or U17791 (N_17791,N_17448,N_17456);
and U17792 (N_17792,N_17312,N_17177);
and U17793 (N_17793,N_17059,N_17442);
and U17794 (N_17794,N_17110,N_17080);
or U17795 (N_17795,N_17456,N_17256);
or U17796 (N_17796,N_17316,N_17193);
nand U17797 (N_17797,N_17408,N_17252);
nor U17798 (N_17798,N_17409,N_17345);
xor U17799 (N_17799,N_17326,N_17265);
xnor U17800 (N_17800,N_17051,N_17377);
nand U17801 (N_17801,N_17209,N_17089);
nor U17802 (N_17802,N_17405,N_17007);
and U17803 (N_17803,N_17456,N_17130);
xor U17804 (N_17804,N_17304,N_17093);
nand U17805 (N_17805,N_17192,N_17252);
or U17806 (N_17806,N_17132,N_17373);
or U17807 (N_17807,N_17480,N_17096);
nor U17808 (N_17808,N_17328,N_17137);
nand U17809 (N_17809,N_17298,N_17265);
xnor U17810 (N_17810,N_17179,N_17241);
or U17811 (N_17811,N_17052,N_17298);
or U17812 (N_17812,N_17424,N_17115);
and U17813 (N_17813,N_17025,N_17135);
nor U17814 (N_17814,N_17017,N_17485);
nor U17815 (N_17815,N_17114,N_17487);
and U17816 (N_17816,N_17062,N_17255);
or U17817 (N_17817,N_17047,N_17337);
nor U17818 (N_17818,N_17476,N_17261);
nand U17819 (N_17819,N_17196,N_17108);
and U17820 (N_17820,N_17095,N_17406);
or U17821 (N_17821,N_17116,N_17314);
or U17822 (N_17822,N_17267,N_17274);
nor U17823 (N_17823,N_17457,N_17340);
and U17824 (N_17824,N_17396,N_17269);
nor U17825 (N_17825,N_17106,N_17393);
nand U17826 (N_17826,N_17299,N_17070);
and U17827 (N_17827,N_17330,N_17046);
nand U17828 (N_17828,N_17117,N_17196);
and U17829 (N_17829,N_17397,N_17364);
or U17830 (N_17830,N_17266,N_17407);
and U17831 (N_17831,N_17119,N_17016);
xor U17832 (N_17832,N_17283,N_17369);
and U17833 (N_17833,N_17441,N_17269);
nor U17834 (N_17834,N_17153,N_17183);
nand U17835 (N_17835,N_17100,N_17421);
nand U17836 (N_17836,N_17057,N_17382);
and U17837 (N_17837,N_17496,N_17203);
xor U17838 (N_17838,N_17270,N_17464);
nand U17839 (N_17839,N_17335,N_17454);
nor U17840 (N_17840,N_17327,N_17349);
and U17841 (N_17841,N_17107,N_17426);
nand U17842 (N_17842,N_17170,N_17253);
nand U17843 (N_17843,N_17152,N_17250);
and U17844 (N_17844,N_17420,N_17236);
xor U17845 (N_17845,N_17225,N_17222);
and U17846 (N_17846,N_17085,N_17336);
nor U17847 (N_17847,N_17498,N_17008);
nor U17848 (N_17848,N_17346,N_17407);
xnor U17849 (N_17849,N_17443,N_17158);
nor U17850 (N_17850,N_17472,N_17247);
and U17851 (N_17851,N_17206,N_17406);
or U17852 (N_17852,N_17193,N_17052);
nand U17853 (N_17853,N_17293,N_17007);
xor U17854 (N_17854,N_17249,N_17331);
or U17855 (N_17855,N_17283,N_17443);
or U17856 (N_17856,N_17469,N_17207);
xnor U17857 (N_17857,N_17027,N_17287);
nand U17858 (N_17858,N_17433,N_17232);
nor U17859 (N_17859,N_17077,N_17369);
nand U17860 (N_17860,N_17134,N_17252);
nor U17861 (N_17861,N_17156,N_17235);
xnor U17862 (N_17862,N_17489,N_17295);
and U17863 (N_17863,N_17205,N_17342);
nand U17864 (N_17864,N_17196,N_17069);
or U17865 (N_17865,N_17194,N_17140);
xnor U17866 (N_17866,N_17273,N_17285);
nor U17867 (N_17867,N_17406,N_17021);
xor U17868 (N_17868,N_17124,N_17146);
and U17869 (N_17869,N_17074,N_17493);
or U17870 (N_17870,N_17356,N_17005);
nand U17871 (N_17871,N_17309,N_17279);
or U17872 (N_17872,N_17364,N_17152);
nand U17873 (N_17873,N_17096,N_17467);
or U17874 (N_17874,N_17250,N_17383);
and U17875 (N_17875,N_17312,N_17215);
xnor U17876 (N_17876,N_17419,N_17364);
nand U17877 (N_17877,N_17245,N_17000);
and U17878 (N_17878,N_17363,N_17474);
or U17879 (N_17879,N_17069,N_17385);
or U17880 (N_17880,N_17358,N_17365);
nand U17881 (N_17881,N_17250,N_17241);
nand U17882 (N_17882,N_17350,N_17291);
nand U17883 (N_17883,N_17425,N_17265);
nand U17884 (N_17884,N_17149,N_17356);
or U17885 (N_17885,N_17320,N_17333);
or U17886 (N_17886,N_17042,N_17332);
nor U17887 (N_17887,N_17298,N_17358);
and U17888 (N_17888,N_17221,N_17293);
or U17889 (N_17889,N_17100,N_17040);
and U17890 (N_17890,N_17269,N_17420);
or U17891 (N_17891,N_17188,N_17012);
or U17892 (N_17892,N_17275,N_17331);
or U17893 (N_17893,N_17106,N_17068);
or U17894 (N_17894,N_17185,N_17336);
and U17895 (N_17895,N_17104,N_17139);
nand U17896 (N_17896,N_17171,N_17011);
nand U17897 (N_17897,N_17193,N_17108);
nor U17898 (N_17898,N_17124,N_17264);
and U17899 (N_17899,N_17048,N_17080);
or U17900 (N_17900,N_17334,N_17044);
and U17901 (N_17901,N_17081,N_17195);
nand U17902 (N_17902,N_17480,N_17309);
xnor U17903 (N_17903,N_17188,N_17228);
nor U17904 (N_17904,N_17472,N_17375);
xnor U17905 (N_17905,N_17042,N_17410);
nand U17906 (N_17906,N_17356,N_17451);
and U17907 (N_17907,N_17178,N_17074);
nand U17908 (N_17908,N_17151,N_17341);
nor U17909 (N_17909,N_17474,N_17053);
and U17910 (N_17910,N_17059,N_17066);
xor U17911 (N_17911,N_17447,N_17486);
xor U17912 (N_17912,N_17317,N_17428);
and U17913 (N_17913,N_17359,N_17109);
and U17914 (N_17914,N_17296,N_17313);
xnor U17915 (N_17915,N_17293,N_17349);
and U17916 (N_17916,N_17075,N_17053);
xnor U17917 (N_17917,N_17397,N_17223);
nand U17918 (N_17918,N_17318,N_17211);
nor U17919 (N_17919,N_17458,N_17158);
or U17920 (N_17920,N_17381,N_17166);
nand U17921 (N_17921,N_17041,N_17418);
and U17922 (N_17922,N_17310,N_17288);
or U17923 (N_17923,N_17315,N_17494);
and U17924 (N_17924,N_17323,N_17259);
nor U17925 (N_17925,N_17074,N_17212);
or U17926 (N_17926,N_17486,N_17198);
nand U17927 (N_17927,N_17014,N_17176);
nor U17928 (N_17928,N_17131,N_17198);
xor U17929 (N_17929,N_17451,N_17415);
nor U17930 (N_17930,N_17203,N_17089);
nand U17931 (N_17931,N_17392,N_17110);
xor U17932 (N_17932,N_17095,N_17157);
and U17933 (N_17933,N_17147,N_17172);
or U17934 (N_17934,N_17148,N_17393);
nand U17935 (N_17935,N_17456,N_17459);
nor U17936 (N_17936,N_17268,N_17455);
nor U17937 (N_17937,N_17199,N_17024);
nand U17938 (N_17938,N_17001,N_17407);
xor U17939 (N_17939,N_17300,N_17482);
nor U17940 (N_17940,N_17428,N_17496);
nand U17941 (N_17941,N_17394,N_17396);
or U17942 (N_17942,N_17229,N_17374);
or U17943 (N_17943,N_17118,N_17469);
or U17944 (N_17944,N_17387,N_17242);
nor U17945 (N_17945,N_17312,N_17061);
xnor U17946 (N_17946,N_17267,N_17496);
or U17947 (N_17947,N_17326,N_17261);
nand U17948 (N_17948,N_17277,N_17049);
xor U17949 (N_17949,N_17343,N_17472);
nor U17950 (N_17950,N_17200,N_17172);
xor U17951 (N_17951,N_17189,N_17378);
xnor U17952 (N_17952,N_17215,N_17381);
and U17953 (N_17953,N_17114,N_17344);
nand U17954 (N_17954,N_17046,N_17387);
xnor U17955 (N_17955,N_17315,N_17300);
xor U17956 (N_17956,N_17127,N_17312);
nand U17957 (N_17957,N_17226,N_17311);
nand U17958 (N_17958,N_17432,N_17390);
or U17959 (N_17959,N_17145,N_17394);
nand U17960 (N_17960,N_17366,N_17075);
nor U17961 (N_17961,N_17480,N_17124);
nand U17962 (N_17962,N_17075,N_17264);
or U17963 (N_17963,N_17306,N_17352);
or U17964 (N_17964,N_17249,N_17420);
and U17965 (N_17965,N_17410,N_17116);
nor U17966 (N_17966,N_17280,N_17458);
or U17967 (N_17967,N_17498,N_17040);
nor U17968 (N_17968,N_17133,N_17346);
or U17969 (N_17969,N_17346,N_17193);
nor U17970 (N_17970,N_17494,N_17365);
nand U17971 (N_17971,N_17264,N_17196);
nand U17972 (N_17972,N_17322,N_17206);
nand U17973 (N_17973,N_17423,N_17338);
xnor U17974 (N_17974,N_17004,N_17172);
xnor U17975 (N_17975,N_17237,N_17029);
xor U17976 (N_17976,N_17089,N_17323);
and U17977 (N_17977,N_17366,N_17104);
xor U17978 (N_17978,N_17072,N_17276);
or U17979 (N_17979,N_17177,N_17119);
and U17980 (N_17980,N_17232,N_17235);
nand U17981 (N_17981,N_17493,N_17445);
or U17982 (N_17982,N_17185,N_17042);
or U17983 (N_17983,N_17197,N_17179);
nor U17984 (N_17984,N_17185,N_17093);
xor U17985 (N_17985,N_17279,N_17247);
xnor U17986 (N_17986,N_17205,N_17106);
nor U17987 (N_17987,N_17462,N_17410);
xnor U17988 (N_17988,N_17185,N_17159);
nor U17989 (N_17989,N_17370,N_17125);
xnor U17990 (N_17990,N_17357,N_17006);
xnor U17991 (N_17991,N_17418,N_17457);
nand U17992 (N_17992,N_17002,N_17005);
and U17993 (N_17993,N_17444,N_17418);
xor U17994 (N_17994,N_17071,N_17485);
nor U17995 (N_17995,N_17207,N_17009);
nand U17996 (N_17996,N_17213,N_17082);
nand U17997 (N_17997,N_17159,N_17281);
nor U17998 (N_17998,N_17021,N_17347);
and U17999 (N_17999,N_17412,N_17226);
or U18000 (N_18000,N_17676,N_17814);
or U18001 (N_18001,N_17725,N_17955);
and U18002 (N_18002,N_17980,N_17897);
nand U18003 (N_18003,N_17697,N_17618);
nor U18004 (N_18004,N_17742,N_17642);
xnor U18005 (N_18005,N_17906,N_17520);
or U18006 (N_18006,N_17616,N_17869);
or U18007 (N_18007,N_17913,N_17889);
or U18008 (N_18008,N_17579,N_17507);
nand U18009 (N_18009,N_17510,N_17943);
xor U18010 (N_18010,N_17599,N_17515);
xnor U18011 (N_18011,N_17838,N_17924);
nor U18012 (N_18012,N_17753,N_17537);
and U18013 (N_18013,N_17681,N_17509);
xnor U18014 (N_18014,N_17790,N_17713);
and U18015 (N_18015,N_17904,N_17653);
and U18016 (N_18016,N_17680,N_17709);
nor U18017 (N_18017,N_17857,N_17893);
xnor U18018 (N_18018,N_17929,N_17634);
nand U18019 (N_18019,N_17885,N_17744);
nand U18020 (N_18020,N_17862,N_17819);
xor U18021 (N_18021,N_17738,N_17733);
xor U18022 (N_18022,N_17915,N_17908);
nand U18023 (N_18023,N_17772,N_17797);
and U18024 (N_18024,N_17582,N_17925);
or U18025 (N_18025,N_17597,N_17584);
and U18026 (N_18026,N_17881,N_17916);
nand U18027 (N_18027,N_17707,N_17962);
nor U18028 (N_18028,N_17820,N_17502);
nand U18029 (N_18029,N_17706,N_17677);
xor U18030 (N_18030,N_17778,N_17636);
and U18031 (N_18031,N_17831,N_17546);
and U18032 (N_18032,N_17934,N_17526);
nand U18033 (N_18033,N_17909,N_17567);
and U18034 (N_18034,N_17570,N_17566);
or U18035 (N_18035,N_17796,N_17606);
nor U18036 (N_18036,N_17583,N_17506);
nand U18037 (N_18037,N_17734,N_17754);
xor U18038 (N_18038,N_17817,N_17731);
or U18039 (N_18039,N_17821,N_17740);
nand U18040 (N_18040,N_17755,N_17927);
nand U18041 (N_18041,N_17612,N_17837);
and U18042 (N_18042,N_17504,N_17780);
and U18043 (N_18043,N_17699,N_17628);
nor U18044 (N_18044,N_17545,N_17611);
nand U18045 (N_18045,N_17593,N_17947);
xor U18046 (N_18046,N_17933,N_17688);
xor U18047 (N_18047,N_17708,N_17660);
and U18048 (N_18048,N_17842,N_17890);
and U18049 (N_18049,N_17967,N_17860);
nand U18050 (N_18050,N_17609,N_17964);
nor U18051 (N_18051,N_17861,N_17696);
or U18052 (N_18052,N_17539,N_17730);
or U18053 (N_18053,N_17850,N_17588);
nand U18054 (N_18054,N_17601,N_17878);
or U18055 (N_18055,N_17843,N_17750);
xnor U18056 (N_18056,N_17716,N_17759);
or U18057 (N_18057,N_17525,N_17595);
nand U18058 (N_18058,N_17517,N_17991);
xnor U18059 (N_18059,N_17942,N_17719);
or U18060 (N_18060,N_17779,N_17970);
xor U18061 (N_18061,N_17631,N_17559);
or U18062 (N_18062,N_17587,N_17528);
and U18063 (N_18063,N_17959,N_17690);
and U18064 (N_18064,N_17990,N_17605);
nand U18065 (N_18065,N_17912,N_17640);
nor U18066 (N_18066,N_17589,N_17701);
and U18067 (N_18067,N_17996,N_17921);
and U18068 (N_18068,N_17864,N_17918);
or U18069 (N_18069,N_17939,N_17807);
and U18070 (N_18070,N_17580,N_17718);
or U18071 (N_18071,N_17795,N_17729);
nor U18072 (N_18072,N_17594,N_17532);
or U18073 (N_18073,N_17765,N_17988);
and U18074 (N_18074,N_17997,N_17931);
nand U18075 (N_18075,N_17669,N_17743);
nand U18076 (N_18076,N_17500,N_17828);
nand U18077 (N_18077,N_17674,N_17639);
xor U18078 (N_18078,N_17766,N_17882);
nor U18079 (N_18079,N_17949,N_17829);
nor U18080 (N_18080,N_17935,N_17863);
nor U18081 (N_18081,N_17784,N_17622);
and U18082 (N_18082,N_17787,N_17717);
nor U18083 (N_18083,N_17815,N_17608);
or U18084 (N_18084,N_17875,N_17969);
nor U18085 (N_18085,N_17656,N_17793);
nor U18086 (N_18086,N_17961,N_17705);
nor U18087 (N_18087,N_17663,N_17693);
or U18088 (N_18088,N_17675,N_17826);
or U18089 (N_18089,N_17768,N_17569);
nand U18090 (N_18090,N_17662,N_17521);
or U18091 (N_18091,N_17541,N_17548);
nor U18092 (N_18092,N_17971,N_17945);
xnor U18093 (N_18093,N_17602,N_17886);
xor U18094 (N_18094,N_17505,N_17747);
or U18095 (N_18095,N_17694,N_17848);
or U18096 (N_18096,N_17518,N_17535);
and U18097 (N_18097,N_17776,N_17799);
or U18098 (N_18098,N_17975,N_17757);
nor U18099 (N_18099,N_17648,N_17655);
and U18100 (N_18100,N_17892,N_17626);
or U18101 (N_18101,N_17806,N_17667);
and U18102 (N_18102,N_17972,N_17572);
or U18103 (N_18103,N_17880,N_17625);
nand U18104 (N_18104,N_17930,N_17522);
nand U18105 (N_18105,N_17685,N_17534);
xnor U18106 (N_18106,N_17888,N_17564);
nand U18107 (N_18107,N_17581,N_17809);
nand U18108 (N_18108,N_17649,N_17651);
or U18109 (N_18109,N_17513,N_17901);
and U18110 (N_18110,N_17610,N_17760);
and U18111 (N_18111,N_17773,N_17987);
nor U18112 (N_18112,N_17849,N_17858);
nand U18113 (N_18113,N_17902,N_17657);
and U18114 (N_18114,N_17907,N_17756);
xnor U18115 (N_18115,N_17895,N_17551);
nand U18116 (N_18116,N_17898,N_17578);
and U18117 (N_18117,N_17683,N_17547);
xor U18118 (N_18118,N_17607,N_17571);
and U18119 (N_18119,N_17562,N_17963);
nor U18120 (N_18120,N_17968,N_17726);
and U18121 (N_18121,N_17977,N_17804);
or U18122 (N_18122,N_17833,N_17560);
nor U18123 (N_18123,N_17698,N_17865);
xnor U18124 (N_18124,N_17900,N_17769);
or U18125 (N_18125,N_17712,N_17512);
nand U18126 (N_18126,N_17650,N_17788);
and U18127 (N_18127,N_17574,N_17585);
or U18128 (N_18128,N_17830,N_17550);
nand U18129 (N_18129,N_17966,N_17956);
xnor U18130 (N_18130,N_17923,N_17710);
and U18131 (N_18131,N_17573,N_17812);
xor U18132 (N_18132,N_17877,N_17530);
and U18133 (N_18133,N_17922,N_17883);
or U18134 (N_18134,N_17714,N_17617);
nand U18135 (N_18135,N_17627,N_17727);
or U18136 (N_18136,N_17533,N_17735);
or U18137 (N_18137,N_17832,N_17552);
and U18138 (N_18138,N_17957,N_17944);
nor U18139 (N_18139,N_17974,N_17576);
and U18140 (N_18140,N_17720,N_17543);
nor U18141 (N_18141,N_17604,N_17700);
nand U18142 (N_18142,N_17846,N_17781);
nor U18143 (N_18143,N_17643,N_17978);
xor U18144 (N_18144,N_17800,N_17982);
nor U18145 (N_18145,N_17686,N_17767);
xor U18146 (N_18146,N_17563,N_17575);
nor U18147 (N_18147,N_17704,N_17758);
nor U18148 (N_18148,N_17917,N_17941);
nor U18149 (N_18149,N_17808,N_17702);
nor U18150 (N_18150,N_17603,N_17899);
xnor U18151 (N_18151,N_17855,N_17866);
nand U18152 (N_18152,N_17994,N_17845);
nor U18153 (N_18153,N_17695,N_17554);
or U18154 (N_18154,N_17501,N_17928);
or U18155 (N_18155,N_17728,N_17519);
nand U18156 (N_18156,N_17981,N_17937);
nand U18157 (N_18157,N_17839,N_17687);
nand U18158 (N_18158,N_17984,N_17771);
and U18159 (N_18159,N_17998,N_17762);
and U18160 (N_18160,N_17868,N_17958);
nand U18161 (N_18161,N_17798,N_17553);
nand U18162 (N_18162,N_17615,N_17508);
xor U18163 (N_18163,N_17646,N_17932);
xnor U18164 (N_18164,N_17973,N_17976);
and U18165 (N_18165,N_17666,N_17884);
xnor U18166 (N_18166,N_17835,N_17722);
nor U18167 (N_18167,N_17891,N_17561);
and U18168 (N_18168,N_17684,N_17825);
and U18169 (N_18169,N_17876,N_17903);
nor U18170 (N_18170,N_17668,N_17527);
nand U18171 (N_18171,N_17624,N_17841);
nand U18172 (N_18172,N_17647,N_17985);
nor U18173 (N_18173,N_17802,N_17993);
or U18174 (N_18174,N_17544,N_17524);
or U18175 (N_18175,N_17568,N_17936);
or U18176 (N_18176,N_17911,N_17818);
or U18177 (N_18177,N_17986,N_17516);
xor U18178 (N_18178,N_17805,N_17785);
xor U18179 (N_18179,N_17590,N_17542);
nand U18180 (N_18180,N_17940,N_17689);
nand U18181 (N_18181,N_17873,N_17792);
xor U18182 (N_18182,N_17816,N_17920);
nor U18183 (N_18183,N_17774,N_17598);
xnor U18184 (N_18184,N_17786,N_17586);
nand U18185 (N_18185,N_17960,N_17999);
nor U18186 (N_18186,N_17775,N_17670);
nor U18187 (N_18187,N_17810,N_17619);
nor U18188 (N_18188,N_17514,N_17761);
xor U18189 (N_18189,N_17844,N_17659);
nor U18190 (N_18190,N_17748,N_17894);
nand U18191 (N_18191,N_17803,N_17919);
xnor U18192 (N_18192,N_17638,N_17853);
nand U18193 (N_18193,N_17989,N_17953);
xor U18194 (N_18194,N_17664,N_17672);
nor U18195 (N_18195,N_17867,N_17874);
nor U18196 (N_18196,N_17538,N_17813);
xor U18197 (N_18197,N_17910,N_17665);
nand U18198 (N_18198,N_17896,N_17637);
nor U18199 (N_18199,N_17801,N_17952);
or U18200 (N_18200,N_17536,N_17852);
and U18201 (N_18201,N_17954,N_17549);
and U18202 (N_18202,N_17946,N_17951);
and U18203 (N_18203,N_17591,N_17763);
and U18204 (N_18204,N_17879,N_17870);
nor U18205 (N_18205,N_17887,N_17556);
and U18206 (N_18206,N_17979,N_17711);
and U18207 (N_18207,N_17926,N_17523);
nand U18208 (N_18208,N_17691,N_17678);
nand U18209 (N_18209,N_17623,N_17789);
xnor U18210 (N_18210,N_17948,N_17600);
nand U18211 (N_18211,N_17840,N_17851);
or U18212 (N_18212,N_17577,N_17746);
xnor U18213 (N_18213,N_17950,N_17682);
nor U18214 (N_18214,N_17692,N_17558);
xor U18215 (N_18215,N_17992,N_17741);
and U18216 (N_18216,N_17724,N_17938);
xor U18217 (N_18217,N_17629,N_17751);
nor U18218 (N_18218,N_17641,N_17965);
and U18219 (N_18219,N_17811,N_17540);
nand U18220 (N_18220,N_17596,N_17827);
xor U18221 (N_18221,N_17592,N_17503);
and U18222 (N_18222,N_17732,N_17633);
nor U18223 (N_18223,N_17652,N_17620);
nor U18224 (N_18224,N_17847,N_17770);
or U18225 (N_18225,N_17983,N_17645);
nor U18226 (N_18226,N_17854,N_17673);
nor U18227 (N_18227,N_17752,N_17679);
and U18228 (N_18228,N_17531,N_17671);
xor U18229 (N_18229,N_17630,N_17822);
nand U18230 (N_18230,N_17621,N_17632);
xor U18231 (N_18231,N_17715,N_17703);
xor U18232 (N_18232,N_17723,N_17859);
nand U18233 (N_18233,N_17872,N_17644);
nor U18234 (N_18234,N_17783,N_17658);
and U18235 (N_18235,N_17836,N_17834);
nor U18236 (N_18236,N_17823,N_17791);
xor U18237 (N_18237,N_17613,N_17871);
and U18238 (N_18238,N_17905,N_17654);
nor U18239 (N_18239,N_17661,N_17736);
nor U18240 (N_18240,N_17856,N_17739);
xnor U18241 (N_18241,N_17565,N_17555);
nor U18242 (N_18242,N_17995,N_17721);
nor U18243 (N_18243,N_17635,N_17777);
xor U18244 (N_18244,N_17794,N_17824);
and U18245 (N_18245,N_17764,N_17745);
nand U18246 (N_18246,N_17749,N_17782);
nor U18247 (N_18247,N_17557,N_17614);
or U18248 (N_18248,N_17529,N_17511);
nand U18249 (N_18249,N_17737,N_17914);
or U18250 (N_18250,N_17811,N_17646);
or U18251 (N_18251,N_17634,N_17784);
and U18252 (N_18252,N_17762,N_17513);
and U18253 (N_18253,N_17771,N_17588);
xnor U18254 (N_18254,N_17957,N_17521);
or U18255 (N_18255,N_17502,N_17646);
xor U18256 (N_18256,N_17927,N_17799);
xor U18257 (N_18257,N_17892,N_17596);
and U18258 (N_18258,N_17993,N_17931);
or U18259 (N_18259,N_17692,N_17852);
or U18260 (N_18260,N_17803,N_17786);
xor U18261 (N_18261,N_17727,N_17918);
or U18262 (N_18262,N_17543,N_17952);
and U18263 (N_18263,N_17839,N_17604);
nand U18264 (N_18264,N_17774,N_17547);
or U18265 (N_18265,N_17622,N_17935);
and U18266 (N_18266,N_17788,N_17751);
xnor U18267 (N_18267,N_17722,N_17733);
nor U18268 (N_18268,N_17543,N_17844);
xor U18269 (N_18269,N_17686,N_17984);
nor U18270 (N_18270,N_17999,N_17666);
nand U18271 (N_18271,N_17964,N_17541);
or U18272 (N_18272,N_17554,N_17528);
and U18273 (N_18273,N_17614,N_17523);
xor U18274 (N_18274,N_17595,N_17667);
and U18275 (N_18275,N_17525,N_17984);
and U18276 (N_18276,N_17687,N_17563);
xnor U18277 (N_18277,N_17674,N_17522);
nor U18278 (N_18278,N_17595,N_17917);
nor U18279 (N_18279,N_17739,N_17968);
nor U18280 (N_18280,N_17649,N_17766);
nand U18281 (N_18281,N_17855,N_17995);
nand U18282 (N_18282,N_17583,N_17739);
or U18283 (N_18283,N_17845,N_17719);
nor U18284 (N_18284,N_17932,N_17805);
xnor U18285 (N_18285,N_17979,N_17912);
nand U18286 (N_18286,N_17890,N_17761);
nor U18287 (N_18287,N_17968,N_17651);
nand U18288 (N_18288,N_17818,N_17981);
nor U18289 (N_18289,N_17630,N_17918);
or U18290 (N_18290,N_17659,N_17529);
or U18291 (N_18291,N_17977,N_17983);
nand U18292 (N_18292,N_17695,N_17876);
and U18293 (N_18293,N_17717,N_17955);
xnor U18294 (N_18294,N_17661,N_17741);
nor U18295 (N_18295,N_17746,N_17981);
nor U18296 (N_18296,N_17708,N_17621);
and U18297 (N_18297,N_17929,N_17610);
nor U18298 (N_18298,N_17793,N_17871);
nand U18299 (N_18299,N_17555,N_17794);
or U18300 (N_18300,N_17979,N_17978);
xor U18301 (N_18301,N_17756,N_17554);
xnor U18302 (N_18302,N_17735,N_17787);
nor U18303 (N_18303,N_17938,N_17516);
or U18304 (N_18304,N_17517,N_17766);
xor U18305 (N_18305,N_17515,N_17792);
xnor U18306 (N_18306,N_17752,N_17943);
nor U18307 (N_18307,N_17992,N_17977);
or U18308 (N_18308,N_17733,N_17746);
and U18309 (N_18309,N_17946,N_17935);
nand U18310 (N_18310,N_17848,N_17601);
or U18311 (N_18311,N_17552,N_17526);
and U18312 (N_18312,N_17590,N_17978);
nand U18313 (N_18313,N_17566,N_17665);
and U18314 (N_18314,N_17522,N_17981);
or U18315 (N_18315,N_17529,N_17588);
and U18316 (N_18316,N_17589,N_17677);
xor U18317 (N_18317,N_17679,N_17537);
and U18318 (N_18318,N_17643,N_17687);
nor U18319 (N_18319,N_17935,N_17714);
nand U18320 (N_18320,N_17526,N_17645);
and U18321 (N_18321,N_17754,N_17790);
nand U18322 (N_18322,N_17529,N_17578);
and U18323 (N_18323,N_17914,N_17713);
and U18324 (N_18324,N_17998,N_17637);
and U18325 (N_18325,N_17958,N_17573);
or U18326 (N_18326,N_17650,N_17880);
xor U18327 (N_18327,N_17851,N_17846);
nand U18328 (N_18328,N_17841,N_17824);
and U18329 (N_18329,N_17782,N_17512);
xor U18330 (N_18330,N_17988,N_17721);
nor U18331 (N_18331,N_17762,N_17739);
nor U18332 (N_18332,N_17768,N_17630);
nor U18333 (N_18333,N_17647,N_17743);
nand U18334 (N_18334,N_17860,N_17785);
nand U18335 (N_18335,N_17951,N_17762);
and U18336 (N_18336,N_17753,N_17644);
or U18337 (N_18337,N_17913,N_17677);
or U18338 (N_18338,N_17632,N_17985);
or U18339 (N_18339,N_17727,N_17742);
and U18340 (N_18340,N_17935,N_17835);
nand U18341 (N_18341,N_17952,N_17786);
and U18342 (N_18342,N_17800,N_17835);
xnor U18343 (N_18343,N_17620,N_17763);
or U18344 (N_18344,N_17519,N_17744);
nor U18345 (N_18345,N_17809,N_17918);
and U18346 (N_18346,N_17686,N_17854);
xnor U18347 (N_18347,N_17646,N_17756);
nand U18348 (N_18348,N_17917,N_17681);
nor U18349 (N_18349,N_17706,N_17792);
xor U18350 (N_18350,N_17596,N_17691);
or U18351 (N_18351,N_17559,N_17562);
nor U18352 (N_18352,N_17776,N_17567);
and U18353 (N_18353,N_17564,N_17996);
or U18354 (N_18354,N_17712,N_17811);
nor U18355 (N_18355,N_17575,N_17822);
xor U18356 (N_18356,N_17624,N_17764);
nor U18357 (N_18357,N_17638,N_17760);
xnor U18358 (N_18358,N_17993,N_17962);
and U18359 (N_18359,N_17524,N_17939);
nand U18360 (N_18360,N_17979,N_17559);
or U18361 (N_18361,N_17944,N_17510);
nor U18362 (N_18362,N_17883,N_17655);
or U18363 (N_18363,N_17831,N_17633);
nor U18364 (N_18364,N_17818,N_17739);
nor U18365 (N_18365,N_17778,N_17764);
nand U18366 (N_18366,N_17784,N_17707);
and U18367 (N_18367,N_17569,N_17976);
and U18368 (N_18368,N_17528,N_17512);
nor U18369 (N_18369,N_17674,N_17888);
or U18370 (N_18370,N_17690,N_17809);
and U18371 (N_18371,N_17967,N_17673);
or U18372 (N_18372,N_17610,N_17876);
nand U18373 (N_18373,N_17947,N_17962);
xnor U18374 (N_18374,N_17732,N_17929);
and U18375 (N_18375,N_17748,N_17809);
xor U18376 (N_18376,N_17565,N_17521);
nand U18377 (N_18377,N_17885,N_17785);
and U18378 (N_18378,N_17874,N_17681);
nor U18379 (N_18379,N_17787,N_17655);
or U18380 (N_18380,N_17928,N_17626);
xnor U18381 (N_18381,N_17881,N_17582);
xor U18382 (N_18382,N_17707,N_17884);
nand U18383 (N_18383,N_17803,N_17669);
nand U18384 (N_18384,N_17889,N_17523);
xnor U18385 (N_18385,N_17604,N_17828);
nor U18386 (N_18386,N_17675,N_17762);
or U18387 (N_18387,N_17809,N_17620);
or U18388 (N_18388,N_17640,N_17777);
nand U18389 (N_18389,N_17518,N_17734);
xnor U18390 (N_18390,N_17509,N_17893);
xnor U18391 (N_18391,N_17643,N_17694);
xor U18392 (N_18392,N_17942,N_17956);
nor U18393 (N_18393,N_17691,N_17639);
xor U18394 (N_18394,N_17586,N_17661);
and U18395 (N_18395,N_17765,N_17681);
nand U18396 (N_18396,N_17861,N_17816);
and U18397 (N_18397,N_17577,N_17825);
nor U18398 (N_18398,N_17562,N_17776);
nand U18399 (N_18399,N_17679,N_17710);
and U18400 (N_18400,N_17679,N_17869);
nand U18401 (N_18401,N_17953,N_17530);
and U18402 (N_18402,N_17729,N_17823);
or U18403 (N_18403,N_17901,N_17963);
nor U18404 (N_18404,N_17593,N_17873);
xnor U18405 (N_18405,N_17782,N_17784);
nor U18406 (N_18406,N_17934,N_17529);
or U18407 (N_18407,N_17761,N_17568);
xnor U18408 (N_18408,N_17904,N_17543);
and U18409 (N_18409,N_17962,N_17734);
or U18410 (N_18410,N_17549,N_17700);
or U18411 (N_18411,N_17764,N_17581);
and U18412 (N_18412,N_17920,N_17810);
or U18413 (N_18413,N_17915,N_17678);
or U18414 (N_18414,N_17951,N_17770);
and U18415 (N_18415,N_17905,N_17560);
xnor U18416 (N_18416,N_17544,N_17653);
or U18417 (N_18417,N_17610,N_17593);
or U18418 (N_18418,N_17908,N_17669);
or U18419 (N_18419,N_17841,N_17954);
xor U18420 (N_18420,N_17853,N_17837);
nand U18421 (N_18421,N_17797,N_17742);
or U18422 (N_18422,N_17703,N_17793);
and U18423 (N_18423,N_17991,N_17778);
nand U18424 (N_18424,N_17949,N_17815);
or U18425 (N_18425,N_17891,N_17603);
or U18426 (N_18426,N_17791,N_17580);
nand U18427 (N_18427,N_17665,N_17609);
or U18428 (N_18428,N_17572,N_17685);
or U18429 (N_18429,N_17854,N_17962);
nand U18430 (N_18430,N_17955,N_17928);
or U18431 (N_18431,N_17932,N_17501);
or U18432 (N_18432,N_17855,N_17569);
nand U18433 (N_18433,N_17739,N_17923);
and U18434 (N_18434,N_17675,N_17986);
or U18435 (N_18435,N_17568,N_17506);
nor U18436 (N_18436,N_17503,N_17516);
and U18437 (N_18437,N_17848,N_17776);
and U18438 (N_18438,N_17595,N_17970);
nand U18439 (N_18439,N_17773,N_17907);
nand U18440 (N_18440,N_17851,N_17557);
or U18441 (N_18441,N_17806,N_17526);
and U18442 (N_18442,N_17798,N_17742);
nor U18443 (N_18443,N_17557,N_17803);
xnor U18444 (N_18444,N_17692,N_17637);
xnor U18445 (N_18445,N_17682,N_17993);
nor U18446 (N_18446,N_17575,N_17537);
and U18447 (N_18447,N_17577,N_17927);
nand U18448 (N_18448,N_17681,N_17545);
or U18449 (N_18449,N_17976,N_17683);
nor U18450 (N_18450,N_17830,N_17859);
nor U18451 (N_18451,N_17614,N_17602);
nor U18452 (N_18452,N_17775,N_17872);
xor U18453 (N_18453,N_17937,N_17925);
or U18454 (N_18454,N_17852,N_17746);
xnor U18455 (N_18455,N_17549,N_17841);
or U18456 (N_18456,N_17947,N_17731);
and U18457 (N_18457,N_17713,N_17653);
nor U18458 (N_18458,N_17814,N_17786);
or U18459 (N_18459,N_17864,N_17697);
nand U18460 (N_18460,N_17640,N_17740);
nor U18461 (N_18461,N_17942,N_17823);
and U18462 (N_18462,N_17903,N_17628);
and U18463 (N_18463,N_17981,N_17616);
xor U18464 (N_18464,N_17631,N_17675);
xor U18465 (N_18465,N_17617,N_17917);
nor U18466 (N_18466,N_17765,N_17806);
or U18467 (N_18467,N_17907,N_17941);
xnor U18468 (N_18468,N_17768,N_17539);
nand U18469 (N_18469,N_17597,N_17606);
nor U18470 (N_18470,N_17596,N_17712);
nor U18471 (N_18471,N_17822,N_17591);
xnor U18472 (N_18472,N_17728,N_17808);
or U18473 (N_18473,N_17656,N_17909);
nand U18474 (N_18474,N_17864,N_17740);
or U18475 (N_18475,N_17580,N_17982);
xor U18476 (N_18476,N_17968,N_17888);
xor U18477 (N_18477,N_17922,N_17500);
and U18478 (N_18478,N_17973,N_17829);
nor U18479 (N_18479,N_17695,N_17935);
xnor U18480 (N_18480,N_17532,N_17945);
nand U18481 (N_18481,N_17707,N_17759);
xor U18482 (N_18482,N_17882,N_17625);
nand U18483 (N_18483,N_17837,N_17545);
and U18484 (N_18484,N_17729,N_17698);
and U18485 (N_18485,N_17502,N_17612);
and U18486 (N_18486,N_17754,N_17963);
or U18487 (N_18487,N_17926,N_17533);
xnor U18488 (N_18488,N_17864,N_17981);
and U18489 (N_18489,N_17592,N_17807);
and U18490 (N_18490,N_17599,N_17918);
xnor U18491 (N_18491,N_17704,N_17759);
nor U18492 (N_18492,N_17616,N_17906);
and U18493 (N_18493,N_17554,N_17937);
or U18494 (N_18494,N_17994,N_17592);
or U18495 (N_18495,N_17803,N_17857);
and U18496 (N_18496,N_17796,N_17808);
and U18497 (N_18497,N_17742,N_17941);
or U18498 (N_18498,N_17548,N_17868);
nor U18499 (N_18499,N_17592,N_17625);
and U18500 (N_18500,N_18497,N_18123);
nand U18501 (N_18501,N_18414,N_18312);
xnor U18502 (N_18502,N_18023,N_18150);
or U18503 (N_18503,N_18305,N_18470);
xor U18504 (N_18504,N_18263,N_18232);
nand U18505 (N_18505,N_18499,N_18046);
and U18506 (N_18506,N_18304,N_18446);
xor U18507 (N_18507,N_18119,N_18400);
and U18508 (N_18508,N_18125,N_18282);
nor U18509 (N_18509,N_18262,N_18469);
and U18510 (N_18510,N_18315,N_18195);
xor U18511 (N_18511,N_18049,N_18277);
and U18512 (N_18512,N_18308,N_18116);
and U18513 (N_18513,N_18172,N_18454);
xnor U18514 (N_18514,N_18124,N_18292);
xnor U18515 (N_18515,N_18090,N_18412);
or U18516 (N_18516,N_18081,N_18160);
or U18517 (N_18517,N_18214,N_18426);
or U18518 (N_18518,N_18145,N_18171);
nand U18519 (N_18519,N_18130,N_18323);
nand U18520 (N_18520,N_18228,N_18436);
nand U18521 (N_18521,N_18389,N_18102);
xor U18522 (N_18522,N_18005,N_18168);
nand U18523 (N_18523,N_18182,N_18121);
nor U18524 (N_18524,N_18202,N_18492);
nor U18525 (N_18525,N_18165,N_18151);
or U18526 (N_18526,N_18293,N_18169);
or U18527 (N_18527,N_18427,N_18137);
nand U18528 (N_18528,N_18474,N_18087);
nor U18529 (N_18529,N_18114,N_18284);
and U18530 (N_18530,N_18348,N_18043);
xor U18531 (N_18531,N_18140,N_18144);
nand U18532 (N_18532,N_18268,N_18175);
and U18533 (N_18533,N_18158,N_18237);
nand U18534 (N_18534,N_18111,N_18489);
or U18535 (N_18535,N_18203,N_18281);
and U18536 (N_18536,N_18373,N_18011);
xnor U18537 (N_18537,N_18340,N_18099);
or U18538 (N_18538,N_18328,N_18456);
xor U18539 (N_18539,N_18197,N_18425);
and U18540 (N_18540,N_18135,N_18227);
nor U18541 (N_18541,N_18076,N_18048);
nand U18542 (N_18542,N_18013,N_18423);
nand U18543 (N_18543,N_18355,N_18117);
xor U18544 (N_18544,N_18342,N_18288);
nor U18545 (N_18545,N_18176,N_18068);
nor U18546 (N_18546,N_18139,N_18387);
xnor U18547 (N_18547,N_18213,N_18255);
nand U18548 (N_18548,N_18283,N_18394);
nor U18549 (N_18549,N_18363,N_18115);
nor U18550 (N_18550,N_18154,N_18494);
or U18551 (N_18551,N_18084,N_18375);
xnor U18552 (N_18552,N_18325,N_18364);
or U18553 (N_18553,N_18476,N_18209);
xor U18554 (N_18554,N_18174,N_18337);
and U18555 (N_18555,N_18485,N_18257);
or U18556 (N_18556,N_18444,N_18194);
nor U18557 (N_18557,N_18067,N_18314);
and U18558 (N_18558,N_18461,N_18396);
and U18559 (N_18559,N_18062,N_18368);
and U18560 (N_18560,N_18391,N_18138);
xor U18561 (N_18561,N_18256,N_18153);
nor U18562 (N_18562,N_18180,N_18251);
and U18563 (N_18563,N_18215,N_18261);
xnor U18564 (N_18564,N_18190,N_18411);
xnor U18565 (N_18565,N_18258,N_18351);
or U18566 (N_18566,N_18462,N_18073);
or U18567 (N_18567,N_18422,N_18302);
and U18568 (N_18568,N_18059,N_18108);
xnor U18569 (N_18569,N_18430,N_18272);
nand U18570 (N_18570,N_18353,N_18134);
xnor U18571 (N_18571,N_18047,N_18061);
nand U18572 (N_18572,N_18109,N_18239);
and U18573 (N_18573,N_18481,N_18352);
or U18574 (N_18574,N_18279,N_18206);
nand U18575 (N_18575,N_18432,N_18393);
xor U18576 (N_18576,N_18045,N_18086);
nor U18577 (N_18577,N_18468,N_18088);
nand U18578 (N_18578,N_18035,N_18357);
and U18579 (N_18579,N_18185,N_18001);
nand U18580 (N_18580,N_18204,N_18475);
xnor U18581 (N_18581,N_18424,N_18056);
and U18582 (N_18582,N_18147,N_18242);
nand U18583 (N_18583,N_18041,N_18372);
or U18584 (N_18584,N_18007,N_18397);
or U18585 (N_18585,N_18163,N_18004);
and U18586 (N_18586,N_18224,N_18126);
nor U18587 (N_18587,N_18120,N_18069);
nand U18588 (N_18588,N_18344,N_18039);
nand U18589 (N_18589,N_18338,N_18085);
or U18590 (N_18590,N_18455,N_18271);
or U18591 (N_18591,N_18026,N_18266);
or U18592 (N_18592,N_18198,N_18409);
or U18593 (N_18593,N_18162,N_18399);
or U18594 (N_18594,N_18188,N_18301);
and U18595 (N_18595,N_18128,N_18415);
xor U18596 (N_18596,N_18094,N_18066);
nor U18597 (N_18597,N_18038,N_18447);
and U18598 (N_18598,N_18365,N_18441);
xnor U18599 (N_18599,N_18452,N_18332);
nand U18600 (N_18600,N_18486,N_18463);
and U18601 (N_18601,N_18296,N_18410);
xor U18602 (N_18602,N_18434,N_18129);
nand U18603 (N_18603,N_18419,N_18278);
xor U18604 (N_18604,N_18071,N_18220);
xnor U18605 (N_18605,N_18280,N_18478);
xor U18606 (N_18606,N_18244,N_18466);
nor U18607 (N_18607,N_18063,N_18388);
nand U18608 (N_18608,N_18386,N_18498);
xnor U18609 (N_18609,N_18378,N_18127);
and U18610 (N_18610,N_18101,N_18330);
xnor U18611 (N_18611,N_18217,N_18420);
and U18612 (N_18612,N_18253,N_18407);
nand U18613 (N_18613,N_18313,N_18226);
nor U18614 (N_18614,N_18054,N_18377);
and U18615 (N_18615,N_18300,N_18491);
nor U18616 (N_18616,N_18095,N_18448);
or U18617 (N_18617,N_18369,N_18082);
xor U18618 (N_18618,N_18183,N_18181);
xnor U18619 (N_18619,N_18376,N_18210);
nor U18620 (N_18620,N_18029,N_18297);
or U18621 (N_18621,N_18083,N_18316);
and U18622 (N_18622,N_18383,N_18488);
nand U18623 (N_18623,N_18006,N_18319);
xor U18624 (N_18624,N_18052,N_18247);
or U18625 (N_18625,N_18453,N_18092);
nor U18626 (N_18626,N_18070,N_18398);
nor U18627 (N_18627,N_18199,N_18339);
xor U18628 (N_18628,N_18072,N_18496);
and U18629 (N_18629,N_18347,N_18274);
and U18630 (N_18630,N_18152,N_18093);
xnor U18631 (N_18631,N_18249,N_18350);
or U18632 (N_18632,N_18349,N_18042);
xnor U18633 (N_18633,N_18290,N_18177);
and U18634 (N_18634,N_18345,N_18459);
or U18635 (N_18635,N_18166,N_18473);
nand U18636 (N_18636,N_18077,N_18421);
xor U18637 (N_18637,N_18022,N_18104);
xor U18638 (N_18638,N_18472,N_18103);
nor U18639 (N_18639,N_18318,N_18065);
or U18640 (N_18640,N_18431,N_18053);
or U18641 (N_18641,N_18034,N_18259);
nor U18642 (N_18642,N_18321,N_18136);
or U18643 (N_18643,N_18324,N_18219);
nand U18644 (N_18644,N_18385,N_18458);
xnor U18645 (N_18645,N_18435,N_18367);
xnor U18646 (N_18646,N_18406,N_18200);
or U18647 (N_18647,N_18016,N_18250);
and U18648 (N_18648,N_18078,N_18055);
nand U18649 (N_18649,N_18295,N_18429);
or U18650 (N_18650,N_18019,N_18142);
nand U18651 (N_18651,N_18225,N_18107);
or U18652 (N_18652,N_18012,N_18014);
nor U18653 (N_18653,N_18311,N_18418);
or U18654 (N_18654,N_18359,N_18403);
nor U18655 (N_18655,N_18408,N_18428);
xnor U18656 (N_18656,N_18231,N_18405);
nand U18657 (N_18657,N_18031,N_18437);
and U18658 (N_18658,N_18112,N_18075);
and U18659 (N_18659,N_18471,N_18003);
nand U18660 (N_18660,N_18449,N_18482);
nor U18661 (N_18661,N_18370,N_18156);
or U18662 (N_18662,N_18159,N_18229);
nor U18663 (N_18663,N_18241,N_18265);
nand U18664 (N_18664,N_18433,N_18036);
nand U18665 (N_18665,N_18341,N_18015);
nor U18666 (N_18666,N_18098,N_18218);
and U18667 (N_18667,N_18100,N_18211);
and U18668 (N_18668,N_18221,N_18331);
xor U18669 (N_18669,N_18322,N_18192);
nor U18670 (N_18670,N_18000,N_18273);
nor U18671 (N_18671,N_18057,N_18133);
nor U18672 (N_18672,N_18243,N_18392);
and U18673 (N_18673,N_18382,N_18484);
nor U18674 (N_18674,N_18413,N_18050);
and U18675 (N_18675,N_18254,N_18208);
nand U18676 (N_18676,N_18490,N_18487);
nand U18677 (N_18677,N_18106,N_18021);
xor U18678 (N_18678,N_18270,N_18167);
and U18679 (N_18679,N_18234,N_18445);
or U18680 (N_18680,N_18064,N_18384);
and U18681 (N_18681,N_18381,N_18390);
or U18682 (N_18682,N_18223,N_18189);
xnor U18683 (N_18683,N_18450,N_18310);
or U18684 (N_18684,N_18245,N_18196);
xor U18685 (N_18685,N_18289,N_18010);
xor U18686 (N_18686,N_18178,N_18326);
or U18687 (N_18687,N_18457,N_18366);
and U18688 (N_18688,N_18089,N_18033);
xnor U18689 (N_18689,N_18264,N_18236);
and U18690 (N_18690,N_18334,N_18122);
nand U18691 (N_18691,N_18360,N_18132);
nand U18692 (N_18692,N_18027,N_18238);
or U18693 (N_18693,N_18193,N_18028);
nand U18694 (N_18694,N_18191,N_18358);
and U18695 (N_18695,N_18287,N_18024);
or U18696 (N_18696,N_18002,N_18020);
or U18697 (N_18697,N_18155,N_18483);
nor U18698 (N_18698,N_18044,N_18161);
or U18699 (N_18699,N_18074,N_18495);
xnor U18700 (N_18700,N_18205,N_18096);
nand U18701 (N_18701,N_18320,N_18164);
or U18702 (N_18702,N_18118,N_18395);
xor U18703 (N_18703,N_18333,N_18252);
and U18704 (N_18704,N_18317,N_18362);
nor U18705 (N_18705,N_18299,N_18025);
and U18706 (N_18706,N_18404,N_18346);
nor U18707 (N_18707,N_18079,N_18184);
nor U18708 (N_18708,N_18212,N_18148);
nor U18709 (N_18709,N_18294,N_18187);
and U18710 (N_18710,N_18438,N_18131);
xnor U18711 (N_18711,N_18240,N_18285);
xor U18712 (N_18712,N_18105,N_18008);
and U18713 (N_18713,N_18451,N_18248);
nor U18714 (N_18714,N_18402,N_18467);
nor U18715 (N_18715,N_18361,N_18207);
or U18716 (N_18716,N_18267,N_18329);
xnor U18717 (N_18717,N_18298,N_18309);
nor U18718 (N_18718,N_18216,N_18439);
or U18719 (N_18719,N_18246,N_18335);
nand U18720 (N_18720,N_18009,N_18380);
nor U18721 (N_18721,N_18379,N_18143);
and U18722 (N_18722,N_18222,N_18465);
xnor U18723 (N_18723,N_18032,N_18186);
nor U18724 (N_18724,N_18051,N_18442);
or U18725 (N_18725,N_18201,N_18037);
or U18726 (N_18726,N_18030,N_18480);
nor U18727 (N_18727,N_18286,N_18230);
and U18728 (N_18728,N_18443,N_18276);
nor U18729 (N_18729,N_18091,N_18356);
xor U18730 (N_18730,N_18113,N_18464);
xor U18731 (N_18731,N_18018,N_18269);
and U18732 (N_18732,N_18440,N_18275);
nor U18733 (N_18733,N_18291,N_18170);
nor U18734 (N_18734,N_18110,N_18371);
nor U18735 (N_18735,N_18336,N_18060);
nor U18736 (N_18736,N_18479,N_18460);
xnor U18737 (N_18737,N_18040,N_18307);
nor U18738 (N_18738,N_18149,N_18260);
or U18739 (N_18739,N_18401,N_18097);
or U18740 (N_18740,N_18233,N_18179);
nand U18741 (N_18741,N_18173,N_18157);
or U18742 (N_18742,N_18306,N_18058);
nand U18743 (N_18743,N_18017,N_18354);
or U18744 (N_18744,N_18417,N_18235);
nand U18745 (N_18745,N_18303,N_18080);
and U18746 (N_18746,N_18146,N_18416);
nand U18747 (N_18747,N_18141,N_18374);
xnor U18748 (N_18748,N_18343,N_18493);
nor U18749 (N_18749,N_18477,N_18327);
and U18750 (N_18750,N_18003,N_18027);
nor U18751 (N_18751,N_18005,N_18466);
or U18752 (N_18752,N_18249,N_18255);
nor U18753 (N_18753,N_18062,N_18143);
nor U18754 (N_18754,N_18030,N_18024);
nor U18755 (N_18755,N_18403,N_18067);
or U18756 (N_18756,N_18404,N_18417);
xor U18757 (N_18757,N_18228,N_18426);
or U18758 (N_18758,N_18474,N_18079);
xor U18759 (N_18759,N_18180,N_18377);
nor U18760 (N_18760,N_18119,N_18201);
and U18761 (N_18761,N_18099,N_18407);
or U18762 (N_18762,N_18379,N_18124);
and U18763 (N_18763,N_18027,N_18006);
and U18764 (N_18764,N_18398,N_18053);
and U18765 (N_18765,N_18493,N_18366);
or U18766 (N_18766,N_18384,N_18197);
or U18767 (N_18767,N_18035,N_18140);
and U18768 (N_18768,N_18023,N_18498);
nand U18769 (N_18769,N_18307,N_18240);
xor U18770 (N_18770,N_18267,N_18202);
or U18771 (N_18771,N_18022,N_18204);
or U18772 (N_18772,N_18144,N_18104);
nand U18773 (N_18773,N_18261,N_18064);
nand U18774 (N_18774,N_18308,N_18010);
nand U18775 (N_18775,N_18350,N_18463);
and U18776 (N_18776,N_18435,N_18358);
and U18777 (N_18777,N_18253,N_18154);
or U18778 (N_18778,N_18064,N_18151);
nand U18779 (N_18779,N_18171,N_18044);
and U18780 (N_18780,N_18165,N_18175);
and U18781 (N_18781,N_18297,N_18376);
or U18782 (N_18782,N_18323,N_18229);
xnor U18783 (N_18783,N_18233,N_18062);
and U18784 (N_18784,N_18297,N_18097);
nand U18785 (N_18785,N_18231,N_18225);
nand U18786 (N_18786,N_18011,N_18263);
nor U18787 (N_18787,N_18216,N_18311);
xnor U18788 (N_18788,N_18019,N_18040);
xor U18789 (N_18789,N_18061,N_18360);
or U18790 (N_18790,N_18376,N_18007);
xor U18791 (N_18791,N_18444,N_18410);
nor U18792 (N_18792,N_18106,N_18015);
xor U18793 (N_18793,N_18250,N_18422);
or U18794 (N_18794,N_18131,N_18251);
xnor U18795 (N_18795,N_18019,N_18202);
or U18796 (N_18796,N_18103,N_18169);
and U18797 (N_18797,N_18469,N_18320);
nor U18798 (N_18798,N_18221,N_18351);
or U18799 (N_18799,N_18088,N_18191);
or U18800 (N_18800,N_18232,N_18247);
and U18801 (N_18801,N_18252,N_18394);
or U18802 (N_18802,N_18360,N_18397);
and U18803 (N_18803,N_18458,N_18114);
and U18804 (N_18804,N_18253,N_18278);
nand U18805 (N_18805,N_18208,N_18169);
xnor U18806 (N_18806,N_18304,N_18358);
xor U18807 (N_18807,N_18232,N_18259);
nand U18808 (N_18808,N_18084,N_18443);
nand U18809 (N_18809,N_18135,N_18389);
and U18810 (N_18810,N_18178,N_18474);
or U18811 (N_18811,N_18051,N_18274);
nand U18812 (N_18812,N_18009,N_18029);
or U18813 (N_18813,N_18046,N_18251);
and U18814 (N_18814,N_18468,N_18327);
nand U18815 (N_18815,N_18136,N_18023);
nor U18816 (N_18816,N_18003,N_18372);
and U18817 (N_18817,N_18459,N_18196);
nor U18818 (N_18818,N_18095,N_18149);
or U18819 (N_18819,N_18044,N_18442);
xnor U18820 (N_18820,N_18360,N_18246);
nor U18821 (N_18821,N_18137,N_18245);
nor U18822 (N_18822,N_18494,N_18401);
nor U18823 (N_18823,N_18428,N_18322);
nor U18824 (N_18824,N_18048,N_18363);
xnor U18825 (N_18825,N_18432,N_18016);
or U18826 (N_18826,N_18146,N_18279);
or U18827 (N_18827,N_18195,N_18240);
and U18828 (N_18828,N_18041,N_18342);
or U18829 (N_18829,N_18329,N_18035);
nand U18830 (N_18830,N_18408,N_18377);
nand U18831 (N_18831,N_18469,N_18493);
nand U18832 (N_18832,N_18030,N_18407);
or U18833 (N_18833,N_18150,N_18282);
and U18834 (N_18834,N_18291,N_18087);
xor U18835 (N_18835,N_18053,N_18478);
nor U18836 (N_18836,N_18228,N_18449);
or U18837 (N_18837,N_18257,N_18436);
xor U18838 (N_18838,N_18035,N_18067);
nor U18839 (N_18839,N_18483,N_18344);
nor U18840 (N_18840,N_18402,N_18224);
nand U18841 (N_18841,N_18426,N_18241);
nor U18842 (N_18842,N_18448,N_18382);
or U18843 (N_18843,N_18170,N_18340);
or U18844 (N_18844,N_18316,N_18405);
xnor U18845 (N_18845,N_18242,N_18171);
and U18846 (N_18846,N_18327,N_18349);
and U18847 (N_18847,N_18265,N_18059);
and U18848 (N_18848,N_18317,N_18370);
or U18849 (N_18849,N_18023,N_18416);
nor U18850 (N_18850,N_18025,N_18022);
or U18851 (N_18851,N_18095,N_18121);
and U18852 (N_18852,N_18030,N_18100);
nand U18853 (N_18853,N_18154,N_18260);
xor U18854 (N_18854,N_18331,N_18118);
and U18855 (N_18855,N_18395,N_18073);
nor U18856 (N_18856,N_18362,N_18484);
nand U18857 (N_18857,N_18415,N_18098);
nor U18858 (N_18858,N_18412,N_18351);
nor U18859 (N_18859,N_18061,N_18443);
nand U18860 (N_18860,N_18254,N_18418);
nor U18861 (N_18861,N_18135,N_18295);
nor U18862 (N_18862,N_18079,N_18202);
xor U18863 (N_18863,N_18240,N_18383);
and U18864 (N_18864,N_18150,N_18200);
and U18865 (N_18865,N_18437,N_18158);
or U18866 (N_18866,N_18434,N_18127);
nor U18867 (N_18867,N_18356,N_18171);
or U18868 (N_18868,N_18365,N_18422);
or U18869 (N_18869,N_18097,N_18105);
and U18870 (N_18870,N_18229,N_18332);
or U18871 (N_18871,N_18129,N_18185);
nand U18872 (N_18872,N_18435,N_18372);
xor U18873 (N_18873,N_18175,N_18018);
nor U18874 (N_18874,N_18406,N_18095);
nor U18875 (N_18875,N_18234,N_18140);
or U18876 (N_18876,N_18489,N_18270);
and U18877 (N_18877,N_18301,N_18494);
nor U18878 (N_18878,N_18248,N_18078);
and U18879 (N_18879,N_18007,N_18005);
or U18880 (N_18880,N_18259,N_18056);
or U18881 (N_18881,N_18358,N_18070);
or U18882 (N_18882,N_18008,N_18107);
nand U18883 (N_18883,N_18215,N_18270);
or U18884 (N_18884,N_18404,N_18199);
and U18885 (N_18885,N_18399,N_18336);
and U18886 (N_18886,N_18158,N_18266);
nor U18887 (N_18887,N_18212,N_18006);
or U18888 (N_18888,N_18432,N_18416);
xor U18889 (N_18889,N_18028,N_18009);
or U18890 (N_18890,N_18141,N_18013);
nor U18891 (N_18891,N_18225,N_18249);
nand U18892 (N_18892,N_18442,N_18447);
xnor U18893 (N_18893,N_18383,N_18335);
nand U18894 (N_18894,N_18383,N_18088);
or U18895 (N_18895,N_18009,N_18330);
xor U18896 (N_18896,N_18221,N_18340);
nor U18897 (N_18897,N_18444,N_18060);
nand U18898 (N_18898,N_18367,N_18094);
nor U18899 (N_18899,N_18268,N_18192);
nand U18900 (N_18900,N_18173,N_18456);
nand U18901 (N_18901,N_18079,N_18025);
and U18902 (N_18902,N_18244,N_18377);
or U18903 (N_18903,N_18396,N_18381);
or U18904 (N_18904,N_18218,N_18274);
nor U18905 (N_18905,N_18265,N_18025);
xnor U18906 (N_18906,N_18426,N_18384);
and U18907 (N_18907,N_18130,N_18138);
xnor U18908 (N_18908,N_18397,N_18404);
nor U18909 (N_18909,N_18184,N_18245);
or U18910 (N_18910,N_18030,N_18019);
or U18911 (N_18911,N_18323,N_18026);
nor U18912 (N_18912,N_18407,N_18266);
xnor U18913 (N_18913,N_18402,N_18093);
xnor U18914 (N_18914,N_18458,N_18419);
nor U18915 (N_18915,N_18171,N_18260);
nor U18916 (N_18916,N_18064,N_18341);
xor U18917 (N_18917,N_18316,N_18469);
and U18918 (N_18918,N_18238,N_18147);
nand U18919 (N_18919,N_18103,N_18495);
nor U18920 (N_18920,N_18312,N_18455);
or U18921 (N_18921,N_18244,N_18359);
or U18922 (N_18922,N_18429,N_18091);
and U18923 (N_18923,N_18336,N_18417);
xnor U18924 (N_18924,N_18124,N_18203);
xnor U18925 (N_18925,N_18403,N_18113);
xnor U18926 (N_18926,N_18122,N_18479);
or U18927 (N_18927,N_18088,N_18338);
or U18928 (N_18928,N_18270,N_18100);
and U18929 (N_18929,N_18313,N_18170);
or U18930 (N_18930,N_18034,N_18448);
and U18931 (N_18931,N_18493,N_18068);
nand U18932 (N_18932,N_18104,N_18024);
nand U18933 (N_18933,N_18409,N_18382);
nand U18934 (N_18934,N_18297,N_18083);
nor U18935 (N_18935,N_18450,N_18372);
nand U18936 (N_18936,N_18014,N_18399);
xor U18937 (N_18937,N_18430,N_18209);
nor U18938 (N_18938,N_18159,N_18422);
nand U18939 (N_18939,N_18364,N_18175);
or U18940 (N_18940,N_18150,N_18490);
xor U18941 (N_18941,N_18436,N_18258);
nand U18942 (N_18942,N_18431,N_18179);
or U18943 (N_18943,N_18210,N_18395);
or U18944 (N_18944,N_18185,N_18253);
nor U18945 (N_18945,N_18295,N_18268);
nand U18946 (N_18946,N_18342,N_18159);
nor U18947 (N_18947,N_18149,N_18442);
nor U18948 (N_18948,N_18474,N_18363);
xor U18949 (N_18949,N_18259,N_18061);
nor U18950 (N_18950,N_18133,N_18366);
and U18951 (N_18951,N_18054,N_18355);
xnor U18952 (N_18952,N_18385,N_18325);
or U18953 (N_18953,N_18331,N_18251);
and U18954 (N_18954,N_18192,N_18022);
nand U18955 (N_18955,N_18156,N_18298);
or U18956 (N_18956,N_18117,N_18245);
nand U18957 (N_18957,N_18063,N_18395);
xnor U18958 (N_18958,N_18490,N_18338);
or U18959 (N_18959,N_18095,N_18421);
and U18960 (N_18960,N_18124,N_18343);
xnor U18961 (N_18961,N_18407,N_18267);
and U18962 (N_18962,N_18200,N_18004);
or U18963 (N_18963,N_18093,N_18052);
xnor U18964 (N_18964,N_18469,N_18198);
nand U18965 (N_18965,N_18205,N_18355);
xor U18966 (N_18966,N_18463,N_18442);
or U18967 (N_18967,N_18304,N_18453);
nand U18968 (N_18968,N_18250,N_18161);
or U18969 (N_18969,N_18203,N_18370);
or U18970 (N_18970,N_18437,N_18397);
xor U18971 (N_18971,N_18114,N_18347);
nand U18972 (N_18972,N_18055,N_18283);
nor U18973 (N_18973,N_18430,N_18402);
and U18974 (N_18974,N_18168,N_18085);
and U18975 (N_18975,N_18462,N_18154);
and U18976 (N_18976,N_18464,N_18428);
nand U18977 (N_18977,N_18129,N_18277);
xor U18978 (N_18978,N_18185,N_18417);
nor U18979 (N_18979,N_18488,N_18277);
nor U18980 (N_18980,N_18142,N_18055);
and U18981 (N_18981,N_18474,N_18307);
and U18982 (N_18982,N_18300,N_18206);
nor U18983 (N_18983,N_18037,N_18311);
and U18984 (N_18984,N_18234,N_18448);
nor U18985 (N_18985,N_18499,N_18168);
nor U18986 (N_18986,N_18054,N_18242);
xor U18987 (N_18987,N_18356,N_18129);
nor U18988 (N_18988,N_18403,N_18064);
or U18989 (N_18989,N_18194,N_18081);
nand U18990 (N_18990,N_18061,N_18458);
xor U18991 (N_18991,N_18121,N_18093);
or U18992 (N_18992,N_18176,N_18093);
and U18993 (N_18993,N_18389,N_18005);
nand U18994 (N_18994,N_18181,N_18417);
nand U18995 (N_18995,N_18259,N_18008);
nor U18996 (N_18996,N_18393,N_18408);
and U18997 (N_18997,N_18282,N_18319);
nor U18998 (N_18998,N_18130,N_18093);
nor U18999 (N_18999,N_18435,N_18280);
and U19000 (N_19000,N_18546,N_18797);
nand U19001 (N_19001,N_18556,N_18937);
nand U19002 (N_19002,N_18817,N_18846);
nor U19003 (N_19003,N_18988,N_18998);
and U19004 (N_19004,N_18993,N_18819);
and U19005 (N_19005,N_18512,N_18767);
or U19006 (N_19006,N_18590,N_18867);
xnor U19007 (N_19007,N_18895,N_18650);
or U19008 (N_19008,N_18707,N_18602);
nand U19009 (N_19009,N_18757,N_18515);
nor U19010 (N_19010,N_18584,N_18604);
or U19011 (N_19011,N_18997,N_18785);
xnor U19012 (N_19012,N_18522,N_18923);
xor U19013 (N_19013,N_18743,N_18925);
xor U19014 (N_19014,N_18886,N_18645);
and U19015 (N_19015,N_18878,N_18622);
or U19016 (N_19016,N_18549,N_18681);
and U19017 (N_19017,N_18762,N_18862);
or U19018 (N_19018,N_18657,N_18698);
nor U19019 (N_19019,N_18874,N_18502);
and U19020 (N_19020,N_18559,N_18986);
and U19021 (N_19021,N_18844,N_18848);
nand U19022 (N_19022,N_18588,N_18688);
nand U19023 (N_19023,N_18721,N_18784);
nor U19024 (N_19024,N_18894,N_18802);
or U19025 (N_19025,N_18795,N_18551);
nand U19026 (N_19026,N_18912,N_18732);
nand U19027 (N_19027,N_18741,N_18620);
nor U19028 (N_19028,N_18542,N_18643);
or U19029 (N_19029,N_18617,N_18913);
xor U19030 (N_19030,N_18513,N_18979);
nand U19031 (N_19031,N_18634,N_18823);
and U19032 (N_19032,N_18699,N_18853);
or U19033 (N_19033,N_18856,N_18568);
nand U19034 (N_19034,N_18888,N_18609);
nor U19035 (N_19035,N_18552,N_18964);
or U19036 (N_19036,N_18768,N_18991);
nor U19037 (N_19037,N_18800,N_18563);
nor U19038 (N_19038,N_18576,N_18995);
xnor U19039 (N_19039,N_18745,N_18765);
nand U19040 (N_19040,N_18796,N_18591);
xnor U19041 (N_19041,N_18854,N_18792);
nor U19042 (N_19042,N_18934,N_18504);
and U19043 (N_19043,N_18731,N_18756);
nand U19044 (N_19044,N_18526,N_18729);
nor U19045 (N_19045,N_18957,N_18706);
nor U19046 (N_19046,N_18916,N_18586);
and U19047 (N_19047,N_18763,N_18749);
nor U19048 (N_19048,N_18907,N_18766);
or U19049 (N_19049,N_18971,N_18808);
or U19050 (N_19050,N_18892,N_18703);
or U19051 (N_19051,N_18603,N_18669);
xnor U19052 (N_19052,N_18655,N_18921);
and U19053 (N_19053,N_18781,N_18932);
or U19054 (N_19054,N_18735,N_18810);
xnor U19055 (N_19055,N_18582,N_18638);
xnor U19056 (N_19056,N_18969,N_18677);
and U19057 (N_19057,N_18651,N_18889);
xnor U19058 (N_19058,N_18573,N_18543);
or U19059 (N_19059,N_18564,N_18898);
nand U19060 (N_19060,N_18996,N_18697);
or U19061 (N_19061,N_18989,N_18942);
or U19062 (N_19062,N_18560,N_18639);
nand U19063 (N_19063,N_18960,N_18740);
and U19064 (N_19064,N_18812,N_18659);
nor U19065 (N_19065,N_18536,N_18637);
nand U19066 (N_19066,N_18919,N_18652);
nor U19067 (N_19067,N_18719,N_18668);
xor U19068 (N_19068,N_18829,N_18963);
or U19069 (N_19069,N_18857,N_18860);
and U19070 (N_19070,N_18834,N_18570);
xnor U19071 (N_19071,N_18608,N_18647);
nor U19072 (N_19072,N_18877,N_18720);
nor U19073 (N_19073,N_18793,N_18641);
or U19074 (N_19074,N_18709,N_18929);
or U19075 (N_19075,N_18999,N_18572);
xnor U19076 (N_19076,N_18881,N_18702);
and U19077 (N_19077,N_18832,N_18596);
or U19078 (N_19078,N_18683,N_18836);
or U19079 (N_19079,N_18558,N_18565);
nand U19080 (N_19080,N_18672,N_18935);
and U19081 (N_19081,N_18852,N_18624);
nand U19082 (N_19082,N_18820,N_18945);
nor U19083 (N_19083,N_18890,N_18733);
or U19084 (N_19084,N_18712,N_18744);
xnor U19085 (N_19085,N_18725,N_18805);
xor U19086 (N_19086,N_18972,N_18845);
xor U19087 (N_19087,N_18673,N_18701);
nand U19088 (N_19088,N_18789,N_18761);
or U19089 (N_19089,N_18534,N_18627);
nand U19090 (N_19090,N_18692,N_18578);
nor U19091 (N_19091,N_18629,N_18946);
xor U19092 (N_19092,N_18553,N_18633);
nand U19093 (N_19093,N_18779,N_18961);
nand U19094 (N_19094,N_18686,N_18980);
xor U19095 (N_19095,N_18727,N_18966);
xnor U19096 (N_19096,N_18640,N_18505);
nor U19097 (N_19097,N_18911,N_18598);
nand U19098 (N_19098,N_18632,N_18994);
xnor U19099 (N_19099,N_18787,N_18926);
or U19100 (N_19100,N_18630,N_18518);
nor U19101 (N_19101,N_18685,N_18806);
nor U19102 (N_19102,N_18790,N_18694);
nand U19103 (N_19103,N_18696,N_18944);
nand U19104 (N_19104,N_18544,N_18503);
xor U19105 (N_19105,N_18649,N_18855);
nand U19106 (N_19106,N_18516,N_18959);
or U19107 (N_19107,N_18918,N_18597);
and U19108 (N_19108,N_18506,N_18667);
nand U19109 (N_19109,N_18555,N_18962);
and U19110 (N_19110,N_18835,N_18660);
nand U19111 (N_19111,N_18742,N_18747);
and U19112 (N_19112,N_18987,N_18571);
xor U19113 (N_19113,N_18566,N_18753);
xor U19114 (N_19114,N_18953,N_18864);
and U19115 (N_19115,N_18924,N_18983);
xor U19116 (N_19116,N_18738,N_18887);
nor U19117 (N_19117,N_18865,N_18992);
xor U19118 (N_19118,N_18769,N_18858);
nand U19119 (N_19119,N_18548,N_18896);
and U19120 (N_19120,N_18663,N_18816);
xnor U19121 (N_19121,N_18956,N_18521);
nand U19122 (N_19122,N_18607,N_18523);
nand U19123 (N_19123,N_18850,N_18826);
nor U19124 (N_19124,N_18818,N_18517);
xor U19125 (N_19125,N_18938,N_18869);
or U19126 (N_19126,N_18658,N_18990);
xor U19127 (N_19127,N_18827,N_18905);
nand U19128 (N_19128,N_18859,N_18734);
or U19129 (N_19129,N_18567,N_18876);
or U19130 (N_19130,N_18939,N_18958);
nor U19131 (N_19131,N_18847,N_18750);
or U19132 (N_19132,N_18884,N_18705);
nor U19133 (N_19133,N_18626,N_18977);
xnor U19134 (N_19134,N_18581,N_18809);
xor U19135 (N_19135,N_18759,N_18840);
nor U19136 (N_19136,N_18531,N_18868);
nand U19137 (N_19137,N_18751,N_18982);
nor U19138 (N_19138,N_18941,N_18654);
and U19139 (N_19139,N_18838,N_18891);
xor U19140 (N_19140,N_18967,N_18936);
and U19141 (N_19141,N_18691,N_18830);
and U19142 (N_19142,N_18601,N_18822);
nor U19143 (N_19143,N_18955,N_18613);
nand U19144 (N_19144,N_18695,N_18831);
nor U19145 (N_19145,N_18550,N_18915);
or U19146 (N_19146,N_18870,N_18863);
and U19147 (N_19147,N_18533,N_18511);
xnor U19148 (N_19148,N_18737,N_18801);
or U19149 (N_19149,N_18611,N_18680);
nor U19150 (N_19150,N_18748,N_18930);
nor U19151 (N_19151,N_18661,N_18928);
nand U19152 (N_19152,N_18833,N_18773);
nand U19153 (N_19153,N_18786,N_18646);
nor U19154 (N_19154,N_18529,N_18580);
nor U19155 (N_19155,N_18662,N_18537);
nor U19156 (N_19156,N_18507,N_18689);
nor U19157 (N_19157,N_18722,N_18614);
nor U19158 (N_19158,N_18981,N_18807);
nor U19159 (N_19159,N_18885,N_18524);
nor U19160 (N_19160,N_18616,N_18950);
nor U19161 (N_19161,N_18909,N_18778);
xor U19162 (N_19162,N_18758,N_18628);
nand U19163 (N_19163,N_18927,N_18554);
and U19164 (N_19164,N_18837,N_18951);
nand U19165 (N_19165,N_18535,N_18714);
nand U19166 (N_19166,N_18538,N_18906);
xnor U19167 (N_19167,N_18562,N_18690);
or U19168 (N_19168,N_18824,N_18711);
nand U19169 (N_19169,N_18772,N_18754);
xor U19170 (N_19170,N_18561,N_18799);
nand U19171 (N_19171,N_18540,N_18775);
or U19172 (N_19172,N_18783,N_18674);
or U19173 (N_19173,N_18900,N_18931);
xnor U19174 (N_19174,N_18615,N_18873);
nor U19175 (N_19175,N_18794,N_18973);
xor U19176 (N_19176,N_18730,N_18700);
and U19177 (N_19177,N_18539,N_18975);
nand U19178 (N_19178,N_18569,N_18501);
xnor U19179 (N_19179,N_18618,N_18849);
or U19180 (N_19180,N_18693,N_18716);
nand U19181 (N_19181,N_18606,N_18713);
xor U19182 (N_19182,N_18947,N_18500);
or U19183 (N_19183,N_18541,N_18592);
and U19184 (N_19184,N_18600,N_18527);
xnor U19185 (N_19185,N_18861,N_18587);
and U19186 (N_19186,N_18871,N_18623);
nand U19187 (N_19187,N_18612,N_18708);
xnor U19188 (N_19188,N_18679,N_18514);
xor U19189 (N_19189,N_18676,N_18520);
and U19190 (N_19190,N_18519,N_18755);
xor U19191 (N_19191,N_18726,N_18682);
nand U19192 (N_19192,N_18509,N_18704);
or U19193 (N_19193,N_18717,N_18595);
nor U19194 (N_19194,N_18771,N_18678);
nand U19195 (N_19195,N_18557,N_18776);
or U19196 (N_19196,N_18510,N_18718);
or U19197 (N_19197,N_18920,N_18798);
nand U19198 (N_19198,N_18901,N_18904);
or U19199 (N_19199,N_18736,N_18943);
and U19200 (N_19200,N_18985,N_18788);
and U19201 (N_19201,N_18724,N_18914);
or U19202 (N_19202,N_18804,N_18665);
nand U19203 (N_19203,N_18774,N_18644);
nand U19204 (N_19204,N_18978,N_18897);
or U19205 (N_19205,N_18948,N_18828);
xor U19206 (N_19206,N_18619,N_18508);
and U19207 (N_19207,N_18675,N_18687);
nand U19208 (N_19208,N_18965,N_18666);
nand U19209 (N_19209,N_18670,N_18528);
nand U19210 (N_19210,N_18764,N_18922);
nor U19211 (N_19211,N_18814,N_18605);
nor U19212 (N_19212,N_18879,N_18594);
or U19213 (N_19213,N_18976,N_18968);
xnor U19214 (N_19214,N_18974,N_18671);
and U19215 (N_19215,N_18899,N_18984);
nand U19216 (N_19216,N_18882,N_18770);
nor U19217 (N_19217,N_18777,N_18545);
or U19218 (N_19218,N_18903,N_18780);
and U19219 (N_19219,N_18530,N_18625);
nand U19220 (N_19220,N_18585,N_18746);
xnor U19221 (N_19221,N_18813,N_18839);
nor U19222 (N_19222,N_18684,N_18811);
xnor U19223 (N_19223,N_18970,N_18575);
or U19224 (N_19224,N_18952,N_18910);
nand U19225 (N_19225,N_18866,N_18574);
xor U19226 (N_19226,N_18893,N_18841);
nand U19227 (N_19227,N_18883,N_18610);
and U19228 (N_19228,N_18599,N_18902);
xnor U19229 (N_19229,N_18949,N_18954);
and U19230 (N_19230,N_18815,N_18656);
xor U19231 (N_19231,N_18715,N_18843);
xnor U19232 (N_19232,N_18739,N_18583);
or U19233 (N_19233,N_18803,N_18917);
nor U19234 (N_19234,N_18579,N_18825);
or U19235 (N_19235,N_18875,N_18940);
and U19236 (N_19236,N_18547,N_18908);
xnor U19237 (N_19237,N_18842,N_18821);
nand U19238 (N_19238,N_18880,N_18593);
nand U19239 (N_19239,N_18782,N_18851);
nand U19240 (N_19240,N_18653,N_18933);
xor U19241 (N_19241,N_18791,N_18577);
xnor U19242 (N_19242,N_18631,N_18532);
nor U19243 (N_19243,N_18710,N_18636);
nand U19244 (N_19244,N_18642,N_18621);
or U19245 (N_19245,N_18635,N_18648);
or U19246 (N_19246,N_18525,N_18723);
and U19247 (N_19247,N_18664,N_18752);
nor U19248 (N_19248,N_18589,N_18872);
or U19249 (N_19249,N_18760,N_18728);
nand U19250 (N_19250,N_18592,N_18744);
nor U19251 (N_19251,N_18676,N_18693);
or U19252 (N_19252,N_18554,N_18906);
and U19253 (N_19253,N_18940,N_18979);
nand U19254 (N_19254,N_18955,N_18681);
or U19255 (N_19255,N_18626,N_18621);
nor U19256 (N_19256,N_18986,N_18690);
nand U19257 (N_19257,N_18725,N_18849);
xor U19258 (N_19258,N_18570,N_18849);
xnor U19259 (N_19259,N_18850,N_18617);
nor U19260 (N_19260,N_18965,N_18798);
and U19261 (N_19261,N_18664,N_18642);
and U19262 (N_19262,N_18940,N_18975);
nor U19263 (N_19263,N_18781,N_18668);
nor U19264 (N_19264,N_18705,N_18821);
nor U19265 (N_19265,N_18548,N_18816);
xnor U19266 (N_19266,N_18582,N_18944);
and U19267 (N_19267,N_18938,N_18644);
xor U19268 (N_19268,N_18556,N_18895);
or U19269 (N_19269,N_18584,N_18537);
nand U19270 (N_19270,N_18740,N_18803);
or U19271 (N_19271,N_18753,N_18914);
or U19272 (N_19272,N_18867,N_18798);
xor U19273 (N_19273,N_18698,N_18906);
xnor U19274 (N_19274,N_18911,N_18579);
nand U19275 (N_19275,N_18974,N_18941);
and U19276 (N_19276,N_18926,N_18708);
or U19277 (N_19277,N_18680,N_18511);
nand U19278 (N_19278,N_18945,N_18720);
nor U19279 (N_19279,N_18617,N_18633);
nand U19280 (N_19280,N_18870,N_18696);
nor U19281 (N_19281,N_18665,N_18508);
xor U19282 (N_19282,N_18731,N_18832);
or U19283 (N_19283,N_18591,N_18669);
or U19284 (N_19284,N_18543,N_18954);
or U19285 (N_19285,N_18697,N_18664);
and U19286 (N_19286,N_18816,N_18733);
xor U19287 (N_19287,N_18753,N_18608);
nand U19288 (N_19288,N_18575,N_18860);
nand U19289 (N_19289,N_18724,N_18630);
and U19290 (N_19290,N_18839,N_18526);
nor U19291 (N_19291,N_18714,N_18531);
and U19292 (N_19292,N_18503,N_18898);
xor U19293 (N_19293,N_18566,N_18735);
nor U19294 (N_19294,N_18767,N_18759);
xnor U19295 (N_19295,N_18894,N_18779);
or U19296 (N_19296,N_18586,N_18898);
nor U19297 (N_19297,N_18674,N_18509);
nor U19298 (N_19298,N_18500,N_18964);
xor U19299 (N_19299,N_18939,N_18529);
or U19300 (N_19300,N_18791,N_18982);
or U19301 (N_19301,N_18574,N_18549);
xor U19302 (N_19302,N_18744,N_18854);
and U19303 (N_19303,N_18522,N_18978);
xnor U19304 (N_19304,N_18567,N_18563);
or U19305 (N_19305,N_18928,N_18876);
or U19306 (N_19306,N_18914,N_18973);
nor U19307 (N_19307,N_18618,N_18828);
and U19308 (N_19308,N_18699,N_18920);
or U19309 (N_19309,N_18845,N_18507);
nor U19310 (N_19310,N_18794,N_18987);
and U19311 (N_19311,N_18982,N_18528);
xor U19312 (N_19312,N_18930,N_18548);
or U19313 (N_19313,N_18552,N_18564);
xnor U19314 (N_19314,N_18534,N_18642);
xnor U19315 (N_19315,N_18896,N_18973);
and U19316 (N_19316,N_18987,N_18753);
or U19317 (N_19317,N_18733,N_18962);
nor U19318 (N_19318,N_18588,N_18718);
and U19319 (N_19319,N_18576,N_18645);
or U19320 (N_19320,N_18744,N_18821);
and U19321 (N_19321,N_18932,N_18632);
nand U19322 (N_19322,N_18939,N_18564);
or U19323 (N_19323,N_18862,N_18686);
nor U19324 (N_19324,N_18553,N_18632);
xor U19325 (N_19325,N_18514,N_18651);
xor U19326 (N_19326,N_18855,N_18682);
or U19327 (N_19327,N_18833,N_18898);
or U19328 (N_19328,N_18959,N_18749);
nand U19329 (N_19329,N_18958,N_18843);
nand U19330 (N_19330,N_18887,N_18846);
or U19331 (N_19331,N_18615,N_18849);
nor U19332 (N_19332,N_18557,N_18723);
xor U19333 (N_19333,N_18894,N_18897);
and U19334 (N_19334,N_18757,N_18821);
nor U19335 (N_19335,N_18517,N_18612);
xor U19336 (N_19336,N_18822,N_18832);
nor U19337 (N_19337,N_18737,N_18769);
xor U19338 (N_19338,N_18941,N_18712);
nand U19339 (N_19339,N_18764,N_18620);
and U19340 (N_19340,N_18805,N_18554);
xnor U19341 (N_19341,N_18635,N_18766);
or U19342 (N_19342,N_18781,N_18890);
nand U19343 (N_19343,N_18563,N_18604);
nor U19344 (N_19344,N_18775,N_18875);
nand U19345 (N_19345,N_18549,N_18557);
xnor U19346 (N_19346,N_18835,N_18688);
nand U19347 (N_19347,N_18626,N_18615);
and U19348 (N_19348,N_18764,N_18518);
nor U19349 (N_19349,N_18851,N_18793);
xor U19350 (N_19350,N_18552,N_18952);
and U19351 (N_19351,N_18774,N_18805);
and U19352 (N_19352,N_18565,N_18654);
nor U19353 (N_19353,N_18714,N_18680);
or U19354 (N_19354,N_18921,N_18730);
or U19355 (N_19355,N_18817,N_18546);
nand U19356 (N_19356,N_18758,N_18874);
nand U19357 (N_19357,N_18542,N_18947);
nand U19358 (N_19358,N_18705,N_18615);
or U19359 (N_19359,N_18980,N_18702);
or U19360 (N_19360,N_18898,N_18627);
nand U19361 (N_19361,N_18551,N_18649);
nor U19362 (N_19362,N_18840,N_18647);
or U19363 (N_19363,N_18687,N_18637);
or U19364 (N_19364,N_18811,N_18669);
or U19365 (N_19365,N_18720,N_18808);
nand U19366 (N_19366,N_18780,N_18544);
nor U19367 (N_19367,N_18519,N_18500);
nor U19368 (N_19368,N_18567,N_18536);
nor U19369 (N_19369,N_18711,N_18790);
and U19370 (N_19370,N_18706,N_18830);
and U19371 (N_19371,N_18512,N_18747);
nand U19372 (N_19372,N_18976,N_18994);
xor U19373 (N_19373,N_18993,N_18940);
nand U19374 (N_19374,N_18731,N_18796);
and U19375 (N_19375,N_18522,N_18711);
or U19376 (N_19376,N_18914,N_18751);
nand U19377 (N_19377,N_18558,N_18931);
nor U19378 (N_19378,N_18959,N_18521);
nor U19379 (N_19379,N_18865,N_18952);
nand U19380 (N_19380,N_18914,N_18555);
xor U19381 (N_19381,N_18612,N_18521);
or U19382 (N_19382,N_18727,N_18672);
nand U19383 (N_19383,N_18773,N_18679);
and U19384 (N_19384,N_18856,N_18878);
nor U19385 (N_19385,N_18714,N_18702);
nor U19386 (N_19386,N_18680,N_18958);
xor U19387 (N_19387,N_18648,N_18580);
or U19388 (N_19388,N_18829,N_18686);
nor U19389 (N_19389,N_18690,N_18863);
nand U19390 (N_19390,N_18767,N_18617);
nand U19391 (N_19391,N_18556,N_18609);
xnor U19392 (N_19392,N_18606,N_18853);
nand U19393 (N_19393,N_18647,N_18641);
or U19394 (N_19394,N_18848,N_18812);
xor U19395 (N_19395,N_18500,N_18763);
nor U19396 (N_19396,N_18663,N_18680);
xnor U19397 (N_19397,N_18734,N_18727);
nand U19398 (N_19398,N_18844,N_18831);
or U19399 (N_19399,N_18523,N_18783);
and U19400 (N_19400,N_18735,N_18614);
nor U19401 (N_19401,N_18869,N_18622);
and U19402 (N_19402,N_18832,N_18993);
and U19403 (N_19403,N_18811,N_18602);
and U19404 (N_19404,N_18553,N_18945);
or U19405 (N_19405,N_18814,N_18712);
nand U19406 (N_19406,N_18973,N_18833);
xor U19407 (N_19407,N_18739,N_18924);
nand U19408 (N_19408,N_18844,N_18502);
nand U19409 (N_19409,N_18980,N_18666);
xnor U19410 (N_19410,N_18670,N_18803);
and U19411 (N_19411,N_18745,N_18711);
nor U19412 (N_19412,N_18946,N_18530);
and U19413 (N_19413,N_18700,N_18823);
nand U19414 (N_19414,N_18705,N_18953);
nand U19415 (N_19415,N_18700,N_18783);
nand U19416 (N_19416,N_18745,N_18614);
nor U19417 (N_19417,N_18666,N_18827);
nand U19418 (N_19418,N_18865,N_18520);
nand U19419 (N_19419,N_18744,N_18723);
and U19420 (N_19420,N_18636,N_18841);
or U19421 (N_19421,N_18879,N_18682);
or U19422 (N_19422,N_18759,N_18890);
xnor U19423 (N_19423,N_18539,N_18899);
xor U19424 (N_19424,N_18932,N_18981);
nand U19425 (N_19425,N_18836,N_18763);
or U19426 (N_19426,N_18643,N_18772);
nand U19427 (N_19427,N_18679,N_18937);
nor U19428 (N_19428,N_18571,N_18790);
or U19429 (N_19429,N_18970,N_18882);
nor U19430 (N_19430,N_18605,N_18637);
and U19431 (N_19431,N_18610,N_18721);
nand U19432 (N_19432,N_18662,N_18512);
or U19433 (N_19433,N_18995,N_18815);
xor U19434 (N_19434,N_18933,N_18859);
and U19435 (N_19435,N_18785,N_18950);
xnor U19436 (N_19436,N_18822,N_18606);
nand U19437 (N_19437,N_18577,N_18882);
or U19438 (N_19438,N_18807,N_18576);
xor U19439 (N_19439,N_18612,N_18504);
and U19440 (N_19440,N_18635,N_18589);
and U19441 (N_19441,N_18535,N_18920);
or U19442 (N_19442,N_18959,N_18823);
nor U19443 (N_19443,N_18771,N_18844);
nor U19444 (N_19444,N_18563,N_18742);
xor U19445 (N_19445,N_18665,N_18575);
nand U19446 (N_19446,N_18544,N_18781);
nand U19447 (N_19447,N_18821,N_18998);
nor U19448 (N_19448,N_18836,N_18975);
xnor U19449 (N_19449,N_18543,N_18944);
nand U19450 (N_19450,N_18946,N_18555);
and U19451 (N_19451,N_18666,N_18741);
and U19452 (N_19452,N_18696,N_18860);
xor U19453 (N_19453,N_18991,N_18548);
nand U19454 (N_19454,N_18734,N_18774);
nor U19455 (N_19455,N_18681,N_18896);
xor U19456 (N_19456,N_18563,N_18684);
xor U19457 (N_19457,N_18795,N_18804);
nand U19458 (N_19458,N_18942,N_18627);
nor U19459 (N_19459,N_18854,N_18906);
nand U19460 (N_19460,N_18749,N_18608);
nand U19461 (N_19461,N_18753,N_18916);
nand U19462 (N_19462,N_18863,N_18638);
or U19463 (N_19463,N_18640,N_18735);
nand U19464 (N_19464,N_18595,N_18574);
xnor U19465 (N_19465,N_18762,N_18508);
and U19466 (N_19466,N_18503,N_18932);
or U19467 (N_19467,N_18968,N_18701);
xor U19468 (N_19468,N_18604,N_18993);
xnor U19469 (N_19469,N_18987,N_18921);
and U19470 (N_19470,N_18817,N_18505);
nand U19471 (N_19471,N_18528,N_18976);
or U19472 (N_19472,N_18552,N_18709);
nor U19473 (N_19473,N_18639,N_18909);
and U19474 (N_19474,N_18555,N_18747);
or U19475 (N_19475,N_18807,N_18789);
nor U19476 (N_19476,N_18901,N_18647);
nand U19477 (N_19477,N_18945,N_18855);
and U19478 (N_19478,N_18524,N_18600);
and U19479 (N_19479,N_18578,N_18894);
xor U19480 (N_19480,N_18967,N_18665);
nand U19481 (N_19481,N_18849,N_18663);
and U19482 (N_19482,N_18911,N_18685);
nand U19483 (N_19483,N_18643,N_18783);
nand U19484 (N_19484,N_18587,N_18849);
nor U19485 (N_19485,N_18900,N_18893);
or U19486 (N_19486,N_18828,N_18514);
nor U19487 (N_19487,N_18726,N_18786);
nor U19488 (N_19488,N_18842,N_18726);
xor U19489 (N_19489,N_18762,N_18716);
and U19490 (N_19490,N_18569,N_18574);
or U19491 (N_19491,N_18802,N_18501);
nor U19492 (N_19492,N_18730,N_18508);
or U19493 (N_19493,N_18647,N_18738);
nand U19494 (N_19494,N_18634,N_18980);
xnor U19495 (N_19495,N_18552,N_18534);
nor U19496 (N_19496,N_18571,N_18883);
and U19497 (N_19497,N_18737,N_18705);
nor U19498 (N_19498,N_18999,N_18585);
nor U19499 (N_19499,N_18834,N_18774);
or U19500 (N_19500,N_19448,N_19268);
and U19501 (N_19501,N_19497,N_19366);
and U19502 (N_19502,N_19278,N_19145);
nor U19503 (N_19503,N_19462,N_19177);
or U19504 (N_19504,N_19126,N_19224);
or U19505 (N_19505,N_19281,N_19276);
nand U19506 (N_19506,N_19430,N_19110);
and U19507 (N_19507,N_19104,N_19128);
or U19508 (N_19508,N_19286,N_19309);
nor U19509 (N_19509,N_19021,N_19130);
or U19510 (N_19510,N_19258,N_19213);
nor U19511 (N_19511,N_19489,N_19208);
nand U19512 (N_19512,N_19407,N_19354);
nand U19513 (N_19513,N_19120,N_19211);
xor U19514 (N_19514,N_19101,N_19075);
nand U19515 (N_19515,N_19191,N_19297);
or U19516 (N_19516,N_19364,N_19294);
nand U19517 (N_19517,N_19272,N_19105);
and U19518 (N_19518,N_19081,N_19000);
nand U19519 (N_19519,N_19236,N_19209);
xor U19520 (N_19520,N_19119,N_19311);
nor U19521 (N_19521,N_19051,N_19320);
nor U19522 (N_19522,N_19025,N_19280);
nand U19523 (N_19523,N_19234,N_19322);
and U19524 (N_19524,N_19262,N_19499);
or U19525 (N_19525,N_19222,N_19386);
xnor U19526 (N_19526,N_19240,N_19457);
or U19527 (N_19527,N_19397,N_19217);
or U19528 (N_19528,N_19091,N_19377);
xnor U19529 (N_19529,N_19346,N_19432);
nand U19530 (N_19530,N_19201,N_19429);
nor U19531 (N_19531,N_19406,N_19413);
nor U19532 (N_19532,N_19047,N_19405);
nand U19533 (N_19533,N_19328,N_19469);
and U19534 (N_19534,N_19308,N_19060);
xnor U19535 (N_19535,N_19492,N_19160);
and U19536 (N_19536,N_19050,N_19334);
nor U19537 (N_19537,N_19159,N_19395);
and U19538 (N_19538,N_19345,N_19073);
xnor U19539 (N_19539,N_19185,N_19052);
nand U19540 (N_19540,N_19292,N_19284);
xor U19541 (N_19541,N_19491,N_19495);
nand U19542 (N_19542,N_19192,N_19028);
xor U19543 (N_19543,N_19347,N_19404);
or U19544 (N_19544,N_19383,N_19478);
nor U19545 (N_19545,N_19436,N_19166);
nor U19546 (N_19546,N_19238,N_19336);
or U19547 (N_19547,N_19488,N_19199);
or U19548 (N_19548,N_19312,N_19136);
nor U19549 (N_19549,N_19232,N_19250);
xnor U19550 (N_19550,N_19040,N_19034);
nand U19551 (N_19551,N_19269,N_19233);
nor U19552 (N_19552,N_19423,N_19067);
and U19553 (N_19553,N_19323,N_19303);
xor U19554 (N_19554,N_19493,N_19024);
xnor U19555 (N_19555,N_19049,N_19480);
nand U19556 (N_19556,N_19156,N_19263);
nor U19557 (N_19557,N_19291,N_19006);
nand U19558 (N_19558,N_19335,N_19100);
or U19559 (N_19559,N_19113,N_19279);
and U19560 (N_19560,N_19146,N_19450);
nor U19561 (N_19561,N_19362,N_19390);
xnor U19562 (N_19562,N_19064,N_19498);
nor U19563 (N_19563,N_19402,N_19237);
nand U19564 (N_19564,N_19273,N_19307);
or U19565 (N_19565,N_19058,N_19243);
nor U19566 (N_19566,N_19031,N_19443);
and U19567 (N_19567,N_19037,N_19435);
and U19568 (N_19568,N_19274,N_19020);
xor U19569 (N_19569,N_19079,N_19108);
nor U19570 (N_19570,N_19340,N_19218);
nand U19571 (N_19571,N_19415,N_19385);
nor U19572 (N_19572,N_19041,N_19214);
and U19573 (N_19573,N_19044,N_19332);
nand U19574 (N_19574,N_19396,N_19341);
and U19575 (N_19575,N_19143,N_19361);
nand U19576 (N_19576,N_19463,N_19369);
and U19577 (N_19577,N_19056,N_19382);
xnor U19578 (N_19578,N_19427,N_19220);
nor U19579 (N_19579,N_19121,N_19077);
xor U19580 (N_19580,N_19223,N_19168);
xor U19581 (N_19581,N_19378,N_19225);
or U19582 (N_19582,N_19392,N_19318);
nand U19583 (N_19583,N_19290,N_19442);
nor U19584 (N_19584,N_19389,N_19090);
nand U19585 (N_19585,N_19331,N_19017);
and U19586 (N_19586,N_19296,N_19210);
xor U19587 (N_19587,N_19084,N_19476);
or U19588 (N_19588,N_19411,N_19189);
and U19589 (N_19589,N_19456,N_19271);
and U19590 (N_19590,N_19245,N_19251);
or U19591 (N_19591,N_19445,N_19475);
nor U19592 (N_19592,N_19188,N_19381);
nor U19593 (N_19593,N_19097,N_19319);
nand U19594 (N_19594,N_19474,N_19365);
or U19595 (N_19595,N_19471,N_19200);
nand U19596 (N_19596,N_19418,N_19124);
nor U19597 (N_19597,N_19115,N_19012);
and U19598 (N_19598,N_19326,N_19370);
xnor U19599 (N_19599,N_19255,N_19433);
and U19600 (N_19600,N_19198,N_19248);
and U19601 (N_19601,N_19473,N_19464);
nor U19602 (N_19602,N_19419,N_19148);
xor U19603 (N_19603,N_19116,N_19219);
nor U19604 (N_19604,N_19408,N_19235);
nand U19605 (N_19605,N_19313,N_19132);
or U19606 (N_19606,N_19440,N_19015);
or U19607 (N_19607,N_19003,N_19078);
xnor U19608 (N_19608,N_19039,N_19468);
or U19609 (N_19609,N_19428,N_19131);
or U19610 (N_19610,N_19086,N_19212);
nand U19611 (N_19611,N_19324,N_19453);
or U19612 (N_19612,N_19344,N_19002);
nand U19613 (N_19613,N_19122,N_19123);
and U19614 (N_19614,N_19070,N_19111);
or U19615 (N_19615,N_19016,N_19410);
or U19616 (N_19616,N_19302,N_19173);
nor U19617 (N_19617,N_19425,N_19196);
xor U19618 (N_19618,N_19172,N_19096);
nand U19619 (N_19619,N_19246,N_19190);
nand U19620 (N_19620,N_19141,N_19106);
and U19621 (N_19621,N_19005,N_19316);
and U19622 (N_19622,N_19162,N_19367);
and U19623 (N_19623,N_19071,N_19289);
xnor U19624 (N_19624,N_19117,N_19349);
nand U19625 (N_19625,N_19242,N_19048);
xnor U19626 (N_19626,N_19158,N_19061);
nor U19627 (N_19627,N_19252,N_19043);
or U19628 (N_19628,N_19373,N_19348);
xnor U19629 (N_19629,N_19195,N_19342);
nand U19630 (N_19630,N_19446,N_19472);
and U19631 (N_19631,N_19253,N_19151);
xor U19632 (N_19632,N_19321,N_19149);
nor U19633 (N_19633,N_19317,N_19076);
nand U19634 (N_19634,N_19357,N_19412);
nor U19635 (N_19635,N_19065,N_19023);
xor U19636 (N_19636,N_19496,N_19301);
and U19637 (N_19637,N_19103,N_19169);
nor U19638 (N_19638,N_19063,N_19197);
xnor U19639 (N_19639,N_19282,N_19259);
nor U19640 (N_19640,N_19451,N_19387);
nand U19641 (N_19641,N_19186,N_19352);
xor U19642 (N_19642,N_19444,N_19363);
or U19643 (N_19643,N_19339,N_19114);
or U19644 (N_19644,N_19266,N_19306);
and U19645 (N_19645,N_19055,N_19351);
nor U19646 (N_19646,N_19487,N_19455);
xnor U19647 (N_19647,N_19304,N_19482);
xor U19648 (N_19648,N_19007,N_19376);
nor U19649 (N_19649,N_19494,N_19265);
nand U19650 (N_19650,N_19431,N_19356);
or U19651 (N_19651,N_19033,N_19414);
nand U19652 (N_19652,N_19439,N_19082);
or U19653 (N_19653,N_19098,N_19270);
nor U19654 (N_19654,N_19193,N_19062);
and U19655 (N_19655,N_19022,N_19372);
xnor U19656 (N_19656,N_19032,N_19194);
nand U19657 (N_19657,N_19176,N_19484);
nor U19658 (N_19658,N_19138,N_19118);
nor U19659 (N_19659,N_19379,N_19264);
or U19660 (N_19660,N_19483,N_19393);
nand U19661 (N_19661,N_19010,N_19434);
nor U19662 (N_19662,N_19305,N_19355);
nor U19663 (N_19663,N_19204,N_19422);
xnor U19664 (N_19664,N_19454,N_19421);
xnor U19665 (N_19665,N_19458,N_19459);
nand U19666 (N_19666,N_19069,N_19129);
and U19667 (N_19667,N_19202,N_19298);
and U19668 (N_19668,N_19161,N_19452);
and U19669 (N_19669,N_19283,N_19142);
and U19670 (N_19670,N_19150,N_19447);
nor U19671 (N_19671,N_19094,N_19013);
or U19672 (N_19672,N_19384,N_19371);
nor U19673 (N_19673,N_19239,N_19035);
or U19674 (N_19674,N_19267,N_19299);
or U19675 (N_19675,N_19178,N_19368);
nor U19676 (N_19676,N_19315,N_19490);
nand U19677 (N_19677,N_19004,N_19054);
and U19678 (N_19678,N_19231,N_19001);
nor U19679 (N_19679,N_19018,N_19256);
and U19680 (N_19680,N_19045,N_19449);
xnor U19681 (N_19681,N_19438,N_19260);
or U19682 (N_19682,N_19042,N_19477);
and U19683 (N_19683,N_19140,N_19359);
or U19684 (N_19684,N_19295,N_19470);
nor U19685 (N_19685,N_19059,N_19154);
xor U19686 (N_19686,N_19074,N_19241);
nor U19687 (N_19687,N_19329,N_19133);
and U19688 (N_19688,N_19247,N_19107);
or U19689 (N_19689,N_19481,N_19337);
nand U19690 (N_19690,N_19338,N_19226);
or U19691 (N_19691,N_19380,N_19230);
nor U19692 (N_19692,N_19360,N_19424);
nand U19693 (N_19693,N_19403,N_19398);
nand U19694 (N_19694,N_19157,N_19112);
and U19695 (N_19695,N_19011,N_19175);
nor U19696 (N_19696,N_19257,N_19275);
xor U19697 (N_19697,N_19353,N_19485);
nand U19698 (N_19698,N_19479,N_19486);
nand U19699 (N_19699,N_19228,N_19394);
nor U19700 (N_19700,N_19099,N_19019);
or U19701 (N_19701,N_19087,N_19437);
nor U19702 (N_19702,N_19182,N_19467);
and U19703 (N_19703,N_19027,N_19203);
xnor U19704 (N_19704,N_19008,N_19036);
or U19705 (N_19705,N_19314,N_19109);
and U19706 (N_19706,N_19327,N_19333);
or U19707 (N_19707,N_19125,N_19388);
nand U19708 (N_19708,N_19152,N_19441);
nor U19709 (N_19709,N_19134,N_19088);
nor U19710 (N_19710,N_19287,N_19089);
and U19711 (N_19711,N_19288,N_19416);
and U19712 (N_19712,N_19080,N_19300);
xnor U19713 (N_19713,N_19399,N_19068);
xor U19714 (N_19714,N_19009,N_19187);
nand U19715 (N_19715,N_19029,N_19277);
xnor U19716 (N_19716,N_19207,N_19249);
xnor U19717 (N_19717,N_19460,N_19215);
or U19718 (N_19718,N_19310,N_19343);
and U19719 (N_19719,N_19164,N_19053);
xnor U19720 (N_19720,N_19183,N_19466);
xnor U19721 (N_19721,N_19144,N_19391);
xnor U19722 (N_19722,N_19420,N_19254);
and U19723 (N_19723,N_19374,N_19426);
xnor U19724 (N_19724,N_19181,N_19135);
nor U19725 (N_19725,N_19170,N_19375);
or U19726 (N_19726,N_19293,N_19285);
xnor U19727 (N_19727,N_19401,N_19153);
nand U19728 (N_19728,N_19057,N_19330);
and U19729 (N_19729,N_19046,N_19102);
nor U19730 (N_19730,N_19167,N_19066);
nand U19731 (N_19731,N_19092,N_19093);
nor U19732 (N_19732,N_19417,N_19216);
xor U19733 (N_19733,N_19072,N_19038);
or U19734 (N_19734,N_19206,N_19165);
or U19735 (N_19735,N_19137,N_19400);
or U19736 (N_19736,N_19163,N_19147);
nor U19737 (N_19737,N_19221,N_19014);
nor U19738 (N_19738,N_19174,N_19465);
or U19739 (N_19739,N_19325,N_19139);
nand U19740 (N_19740,N_19026,N_19127);
nor U19741 (N_19741,N_19085,N_19350);
nor U19742 (N_19742,N_19171,N_19358);
nor U19743 (N_19743,N_19180,N_19095);
and U19744 (N_19744,N_19155,N_19179);
nand U19745 (N_19745,N_19409,N_19227);
nor U19746 (N_19746,N_19030,N_19229);
nor U19747 (N_19747,N_19083,N_19184);
or U19748 (N_19748,N_19461,N_19205);
xnor U19749 (N_19749,N_19261,N_19244);
xnor U19750 (N_19750,N_19001,N_19050);
nand U19751 (N_19751,N_19052,N_19257);
nor U19752 (N_19752,N_19439,N_19244);
or U19753 (N_19753,N_19499,N_19408);
or U19754 (N_19754,N_19246,N_19224);
nor U19755 (N_19755,N_19337,N_19232);
and U19756 (N_19756,N_19019,N_19150);
xor U19757 (N_19757,N_19263,N_19053);
nand U19758 (N_19758,N_19275,N_19107);
and U19759 (N_19759,N_19113,N_19469);
or U19760 (N_19760,N_19237,N_19155);
and U19761 (N_19761,N_19154,N_19382);
and U19762 (N_19762,N_19255,N_19343);
nor U19763 (N_19763,N_19061,N_19210);
nand U19764 (N_19764,N_19009,N_19201);
or U19765 (N_19765,N_19427,N_19059);
nand U19766 (N_19766,N_19359,N_19042);
and U19767 (N_19767,N_19032,N_19317);
and U19768 (N_19768,N_19382,N_19445);
xor U19769 (N_19769,N_19444,N_19259);
nand U19770 (N_19770,N_19003,N_19400);
nor U19771 (N_19771,N_19405,N_19156);
and U19772 (N_19772,N_19189,N_19353);
nand U19773 (N_19773,N_19169,N_19476);
or U19774 (N_19774,N_19437,N_19177);
and U19775 (N_19775,N_19032,N_19389);
xor U19776 (N_19776,N_19308,N_19417);
or U19777 (N_19777,N_19434,N_19169);
or U19778 (N_19778,N_19061,N_19105);
nor U19779 (N_19779,N_19188,N_19140);
nand U19780 (N_19780,N_19225,N_19498);
and U19781 (N_19781,N_19016,N_19013);
or U19782 (N_19782,N_19024,N_19032);
and U19783 (N_19783,N_19470,N_19337);
nand U19784 (N_19784,N_19418,N_19483);
and U19785 (N_19785,N_19003,N_19402);
nor U19786 (N_19786,N_19488,N_19238);
xnor U19787 (N_19787,N_19381,N_19495);
or U19788 (N_19788,N_19269,N_19055);
xor U19789 (N_19789,N_19114,N_19151);
nor U19790 (N_19790,N_19284,N_19138);
or U19791 (N_19791,N_19125,N_19110);
and U19792 (N_19792,N_19026,N_19447);
and U19793 (N_19793,N_19264,N_19224);
and U19794 (N_19794,N_19383,N_19028);
nand U19795 (N_19795,N_19076,N_19466);
or U19796 (N_19796,N_19030,N_19488);
and U19797 (N_19797,N_19027,N_19081);
and U19798 (N_19798,N_19047,N_19308);
or U19799 (N_19799,N_19217,N_19141);
or U19800 (N_19800,N_19274,N_19223);
xor U19801 (N_19801,N_19354,N_19400);
nand U19802 (N_19802,N_19236,N_19208);
and U19803 (N_19803,N_19418,N_19354);
nor U19804 (N_19804,N_19070,N_19363);
xnor U19805 (N_19805,N_19052,N_19481);
nand U19806 (N_19806,N_19200,N_19183);
nand U19807 (N_19807,N_19107,N_19353);
nor U19808 (N_19808,N_19428,N_19265);
or U19809 (N_19809,N_19132,N_19155);
nor U19810 (N_19810,N_19406,N_19153);
xnor U19811 (N_19811,N_19306,N_19037);
nor U19812 (N_19812,N_19071,N_19146);
or U19813 (N_19813,N_19209,N_19273);
nor U19814 (N_19814,N_19347,N_19363);
and U19815 (N_19815,N_19386,N_19380);
xnor U19816 (N_19816,N_19038,N_19332);
or U19817 (N_19817,N_19094,N_19146);
or U19818 (N_19818,N_19366,N_19118);
nand U19819 (N_19819,N_19337,N_19149);
and U19820 (N_19820,N_19377,N_19197);
nand U19821 (N_19821,N_19157,N_19438);
xor U19822 (N_19822,N_19207,N_19268);
or U19823 (N_19823,N_19489,N_19194);
nand U19824 (N_19824,N_19218,N_19028);
xnor U19825 (N_19825,N_19034,N_19361);
xor U19826 (N_19826,N_19460,N_19082);
or U19827 (N_19827,N_19479,N_19437);
nand U19828 (N_19828,N_19053,N_19319);
or U19829 (N_19829,N_19027,N_19127);
or U19830 (N_19830,N_19236,N_19150);
and U19831 (N_19831,N_19198,N_19452);
or U19832 (N_19832,N_19196,N_19167);
xor U19833 (N_19833,N_19042,N_19002);
or U19834 (N_19834,N_19037,N_19336);
and U19835 (N_19835,N_19093,N_19195);
or U19836 (N_19836,N_19220,N_19122);
or U19837 (N_19837,N_19142,N_19207);
and U19838 (N_19838,N_19225,N_19376);
xor U19839 (N_19839,N_19042,N_19459);
nand U19840 (N_19840,N_19115,N_19026);
xor U19841 (N_19841,N_19053,N_19450);
nor U19842 (N_19842,N_19353,N_19052);
and U19843 (N_19843,N_19446,N_19006);
or U19844 (N_19844,N_19214,N_19180);
nor U19845 (N_19845,N_19460,N_19064);
or U19846 (N_19846,N_19022,N_19299);
xor U19847 (N_19847,N_19238,N_19043);
xor U19848 (N_19848,N_19209,N_19280);
nand U19849 (N_19849,N_19297,N_19176);
xnor U19850 (N_19850,N_19219,N_19285);
nor U19851 (N_19851,N_19198,N_19419);
nand U19852 (N_19852,N_19030,N_19259);
nand U19853 (N_19853,N_19010,N_19148);
xnor U19854 (N_19854,N_19480,N_19224);
nor U19855 (N_19855,N_19446,N_19022);
nand U19856 (N_19856,N_19448,N_19380);
nand U19857 (N_19857,N_19422,N_19162);
xnor U19858 (N_19858,N_19346,N_19023);
and U19859 (N_19859,N_19285,N_19443);
nor U19860 (N_19860,N_19315,N_19475);
xnor U19861 (N_19861,N_19170,N_19113);
or U19862 (N_19862,N_19276,N_19361);
or U19863 (N_19863,N_19217,N_19354);
and U19864 (N_19864,N_19398,N_19400);
nor U19865 (N_19865,N_19292,N_19240);
nand U19866 (N_19866,N_19365,N_19265);
and U19867 (N_19867,N_19010,N_19422);
nor U19868 (N_19868,N_19426,N_19267);
xor U19869 (N_19869,N_19418,N_19448);
nor U19870 (N_19870,N_19053,N_19497);
or U19871 (N_19871,N_19357,N_19130);
or U19872 (N_19872,N_19031,N_19089);
nor U19873 (N_19873,N_19282,N_19116);
nand U19874 (N_19874,N_19170,N_19339);
or U19875 (N_19875,N_19459,N_19361);
nand U19876 (N_19876,N_19089,N_19200);
or U19877 (N_19877,N_19315,N_19419);
nor U19878 (N_19878,N_19238,N_19175);
xnor U19879 (N_19879,N_19163,N_19215);
and U19880 (N_19880,N_19261,N_19273);
nand U19881 (N_19881,N_19343,N_19464);
xnor U19882 (N_19882,N_19129,N_19292);
or U19883 (N_19883,N_19369,N_19065);
and U19884 (N_19884,N_19116,N_19112);
xnor U19885 (N_19885,N_19293,N_19457);
or U19886 (N_19886,N_19258,N_19328);
and U19887 (N_19887,N_19401,N_19110);
nor U19888 (N_19888,N_19088,N_19035);
xnor U19889 (N_19889,N_19455,N_19328);
or U19890 (N_19890,N_19181,N_19114);
xnor U19891 (N_19891,N_19403,N_19270);
or U19892 (N_19892,N_19188,N_19076);
and U19893 (N_19893,N_19466,N_19396);
or U19894 (N_19894,N_19132,N_19396);
or U19895 (N_19895,N_19443,N_19024);
nor U19896 (N_19896,N_19350,N_19458);
nor U19897 (N_19897,N_19398,N_19324);
nand U19898 (N_19898,N_19493,N_19131);
and U19899 (N_19899,N_19023,N_19292);
nor U19900 (N_19900,N_19193,N_19122);
nand U19901 (N_19901,N_19458,N_19266);
and U19902 (N_19902,N_19090,N_19328);
xnor U19903 (N_19903,N_19179,N_19072);
nand U19904 (N_19904,N_19028,N_19149);
xor U19905 (N_19905,N_19198,N_19179);
and U19906 (N_19906,N_19166,N_19073);
and U19907 (N_19907,N_19077,N_19239);
nand U19908 (N_19908,N_19371,N_19407);
xor U19909 (N_19909,N_19387,N_19034);
and U19910 (N_19910,N_19030,N_19418);
nand U19911 (N_19911,N_19335,N_19068);
nand U19912 (N_19912,N_19198,N_19080);
nor U19913 (N_19913,N_19103,N_19354);
nor U19914 (N_19914,N_19003,N_19460);
nand U19915 (N_19915,N_19031,N_19365);
xor U19916 (N_19916,N_19236,N_19333);
nor U19917 (N_19917,N_19022,N_19031);
xor U19918 (N_19918,N_19440,N_19299);
and U19919 (N_19919,N_19208,N_19258);
nor U19920 (N_19920,N_19070,N_19285);
nor U19921 (N_19921,N_19181,N_19165);
or U19922 (N_19922,N_19101,N_19265);
xnor U19923 (N_19923,N_19001,N_19070);
nand U19924 (N_19924,N_19041,N_19450);
nand U19925 (N_19925,N_19089,N_19469);
xor U19926 (N_19926,N_19102,N_19165);
nand U19927 (N_19927,N_19365,N_19221);
nor U19928 (N_19928,N_19093,N_19237);
or U19929 (N_19929,N_19413,N_19443);
and U19930 (N_19930,N_19162,N_19188);
xnor U19931 (N_19931,N_19022,N_19214);
nor U19932 (N_19932,N_19071,N_19485);
or U19933 (N_19933,N_19136,N_19000);
or U19934 (N_19934,N_19130,N_19140);
nand U19935 (N_19935,N_19109,N_19431);
xor U19936 (N_19936,N_19084,N_19390);
nand U19937 (N_19937,N_19464,N_19291);
nor U19938 (N_19938,N_19219,N_19247);
or U19939 (N_19939,N_19368,N_19439);
xnor U19940 (N_19940,N_19466,N_19417);
and U19941 (N_19941,N_19226,N_19434);
xor U19942 (N_19942,N_19326,N_19158);
xnor U19943 (N_19943,N_19228,N_19221);
xnor U19944 (N_19944,N_19277,N_19013);
xnor U19945 (N_19945,N_19052,N_19378);
nand U19946 (N_19946,N_19170,N_19048);
nand U19947 (N_19947,N_19015,N_19178);
nand U19948 (N_19948,N_19439,N_19250);
xor U19949 (N_19949,N_19333,N_19225);
and U19950 (N_19950,N_19027,N_19309);
or U19951 (N_19951,N_19101,N_19358);
nand U19952 (N_19952,N_19049,N_19348);
nor U19953 (N_19953,N_19072,N_19104);
nand U19954 (N_19954,N_19164,N_19325);
nor U19955 (N_19955,N_19008,N_19491);
nand U19956 (N_19956,N_19455,N_19102);
xnor U19957 (N_19957,N_19050,N_19378);
nand U19958 (N_19958,N_19069,N_19448);
xnor U19959 (N_19959,N_19311,N_19403);
or U19960 (N_19960,N_19373,N_19078);
nand U19961 (N_19961,N_19152,N_19494);
nor U19962 (N_19962,N_19310,N_19116);
nand U19963 (N_19963,N_19317,N_19078);
nor U19964 (N_19964,N_19011,N_19161);
nor U19965 (N_19965,N_19304,N_19227);
xor U19966 (N_19966,N_19363,N_19417);
nor U19967 (N_19967,N_19378,N_19145);
nor U19968 (N_19968,N_19381,N_19328);
nand U19969 (N_19969,N_19262,N_19396);
and U19970 (N_19970,N_19480,N_19262);
or U19971 (N_19971,N_19020,N_19423);
or U19972 (N_19972,N_19116,N_19485);
or U19973 (N_19973,N_19026,N_19492);
or U19974 (N_19974,N_19441,N_19045);
nor U19975 (N_19975,N_19485,N_19306);
nand U19976 (N_19976,N_19061,N_19157);
or U19977 (N_19977,N_19420,N_19498);
xor U19978 (N_19978,N_19415,N_19356);
and U19979 (N_19979,N_19349,N_19461);
nor U19980 (N_19980,N_19178,N_19348);
xor U19981 (N_19981,N_19268,N_19121);
and U19982 (N_19982,N_19168,N_19437);
nor U19983 (N_19983,N_19388,N_19122);
and U19984 (N_19984,N_19366,N_19363);
or U19985 (N_19985,N_19012,N_19227);
and U19986 (N_19986,N_19012,N_19345);
or U19987 (N_19987,N_19319,N_19244);
nor U19988 (N_19988,N_19398,N_19375);
nand U19989 (N_19989,N_19376,N_19265);
and U19990 (N_19990,N_19144,N_19184);
or U19991 (N_19991,N_19169,N_19100);
nor U19992 (N_19992,N_19438,N_19046);
or U19993 (N_19993,N_19180,N_19414);
nand U19994 (N_19994,N_19322,N_19422);
nand U19995 (N_19995,N_19010,N_19289);
nand U19996 (N_19996,N_19364,N_19432);
nor U19997 (N_19997,N_19099,N_19344);
nor U19998 (N_19998,N_19464,N_19084);
or U19999 (N_19999,N_19136,N_19061);
nor UO_0 (O_0,N_19738,N_19612);
or UO_1 (O_1,N_19630,N_19861);
nand UO_2 (O_2,N_19645,N_19769);
and UO_3 (O_3,N_19625,N_19588);
and UO_4 (O_4,N_19619,N_19954);
or UO_5 (O_5,N_19979,N_19787);
xnor UO_6 (O_6,N_19981,N_19910);
nor UO_7 (O_7,N_19566,N_19605);
or UO_8 (O_8,N_19674,N_19830);
xor UO_9 (O_9,N_19644,N_19632);
nor UO_10 (O_10,N_19646,N_19693);
nor UO_11 (O_11,N_19567,N_19937);
and UO_12 (O_12,N_19851,N_19871);
nor UO_13 (O_13,N_19989,N_19565);
and UO_14 (O_14,N_19501,N_19660);
or UO_15 (O_15,N_19839,N_19731);
xnor UO_16 (O_16,N_19542,N_19992);
xor UO_17 (O_17,N_19572,N_19672);
nor UO_18 (O_18,N_19704,N_19600);
nor UO_19 (O_19,N_19698,N_19783);
nand UO_20 (O_20,N_19975,N_19626);
or UO_21 (O_21,N_19855,N_19754);
or UO_22 (O_22,N_19797,N_19734);
nand UO_23 (O_23,N_19701,N_19916);
and UO_24 (O_24,N_19997,N_19924);
nor UO_25 (O_25,N_19950,N_19640);
nor UO_26 (O_26,N_19815,N_19750);
xor UO_27 (O_27,N_19584,N_19943);
or UO_28 (O_28,N_19928,N_19993);
and UO_29 (O_29,N_19994,N_19827);
nor UO_30 (O_30,N_19513,N_19836);
or UO_31 (O_31,N_19893,N_19617);
or UO_32 (O_32,N_19814,N_19613);
nor UO_33 (O_33,N_19706,N_19531);
xor UO_34 (O_34,N_19803,N_19875);
nand UO_35 (O_35,N_19877,N_19892);
and UO_36 (O_36,N_19543,N_19708);
or UO_37 (O_37,N_19684,N_19932);
and UO_38 (O_38,N_19604,N_19691);
or UO_39 (O_39,N_19810,N_19707);
or UO_40 (O_40,N_19547,N_19872);
and UO_41 (O_41,N_19823,N_19649);
nor UO_42 (O_42,N_19665,N_19558);
nand UO_43 (O_43,N_19907,N_19801);
xnor UO_44 (O_44,N_19550,N_19618);
or UO_45 (O_45,N_19570,N_19526);
nand UO_46 (O_46,N_19533,N_19862);
xor UO_47 (O_47,N_19522,N_19776);
and UO_48 (O_48,N_19867,N_19723);
nor UO_49 (O_49,N_19843,N_19675);
and UO_50 (O_50,N_19812,N_19933);
xnor UO_51 (O_51,N_19802,N_19510);
nor UO_52 (O_52,N_19695,N_19524);
or UO_53 (O_53,N_19796,N_19821);
xor UO_54 (O_54,N_19541,N_19727);
nor UO_55 (O_55,N_19743,N_19599);
xnor UO_56 (O_56,N_19784,N_19966);
or UO_57 (O_57,N_19809,N_19906);
and UO_58 (O_58,N_19897,N_19752);
and UO_59 (O_59,N_19656,N_19974);
and UO_60 (O_60,N_19895,N_19564);
nand UO_61 (O_61,N_19820,N_19788);
or UO_62 (O_62,N_19987,N_19965);
and UO_63 (O_63,N_19940,N_19984);
and UO_64 (O_64,N_19991,N_19960);
or UO_65 (O_65,N_19887,N_19833);
nor UO_66 (O_66,N_19739,N_19745);
and UO_67 (O_67,N_19848,N_19702);
nor UO_68 (O_68,N_19770,N_19726);
nor UO_69 (O_69,N_19722,N_19751);
and UO_70 (O_70,N_19973,N_19583);
nor UO_71 (O_71,N_19760,N_19904);
xnor UO_72 (O_72,N_19516,N_19792);
nand UO_73 (O_73,N_19900,N_19534);
nand UO_74 (O_74,N_19602,N_19849);
and UO_75 (O_75,N_19757,N_19507);
nor UO_76 (O_76,N_19798,N_19868);
xor UO_77 (O_77,N_19782,N_19901);
nand UO_78 (O_78,N_19712,N_19753);
or UO_79 (O_79,N_19648,N_19955);
and UO_80 (O_80,N_19627,N_19818);
nand UO_81 (O_81,N_19537,N_19999);
xor UO_82 (O_82,N_19768,N_19985);
xnor UO_83 (O_83,N_19554,N_19610);
nand UO_84 (O_84,N_19664,N_19641);
or UO_85 (O_85,N_19905,N_19676);
xor UO_86 (O_86,N_19607,N_19549);
or UO_87 (O_87,N_19864,N_19689);
xor UO_88 (O_88,N_19976,N_19678);
nand UO_89 (O_89,N_19719,N_19765);
nand UO_90 (O_90,N_19755,N_19616);
xor UO_91 (O_91,N_19759,N_19587);
xor UO_92 (O_92,N_19568,N_19594);
nand UO_93 (O_93,N_19687,N_19529);
or UO_94 (O_94,N_19835,N_19655);
and UO_95 (O_95,N_19988,N_19666);
nand UO_96 (O_96,N_19761,N_19560);
or UO_97 (O_97,N_19720,N_19683);
and UO_98 (O_98,N_19575,N_19902);
or UO_99 (O_99,N_19539,N_19934);
nand UO_100 (O_100,N_19585,N_19736);
xnor UO_101 (O_101,N_19786,N_19692);
or UO_102 (O_102,N_19685,N_19576);
nor UO_103 (O_103,N_19816,N_19899);
xnor UO_104 (O_104,N_19650,N_19847);
and UO_105 (O_105,N_19733,N_19525);
nor UO_106 (O_106,N_19824,N_19885);
and UO_107 (O_107,N_19995,N_19948);
nand UO_108 (O_108,N_19742,N_19746);
nor UO_109 (O_109,N_19508,N_19996);
nand UO_110 (O_110,N_19548,N_19914);
and UO_111 (O_111,N_19896,N_19611);
and UO_112 (O_112,N_19747,N_19653);
and UO_113 (O_113,N_19555,N_19980);
nand UO_114 (O_114,N_19832,N_19579);
or UO_115 (O_115,N_19623,N_19710);
nor UO_116 (O_116,N_19777,N_19521);
nor UO_117 (O_117,N_19732,N_19890);
and UO_118 (O_118,N_19961,N_19963);
or UO_119 (O_119,N_19941,N_19721);
nand UO_120 (O_120,N_19898,N_19639);
and UO_121 (O_121,N_19773,N_19523);
and UO_122 (O_122,N_19952,N_19737);
or UO_123 (O_123,N_19962,N_19971);
and UO_124 (O_124,N_19858,N_19629);
or UO_125 (O_125,N_19926,N_19582);
or UO_126 (O_126,N_19621,N_19959);
nand UO_127 (O_127,N_19574,N_19935);
or UO_128 (O_128,N_19735,N_19696);
nor UO_129 (O_129,N_19819,N_19883);
or UO_130 (O_130,N_19859,N_19923);
xor UO_131 (O_131,N_19790,N_19552);
nor UO_132 (O_132,N_19657,N_19535);
or UO_133 (O_133,N_19998,N_19799);
and UO_134 (O_134,N_19822,N_19800);
xor UO_135 (O_135,N_19778,N_19571);
xnor UO_136 (O_136,N_19882,N_19785);
xor UO_137 (O_137,N_19563,N_19667);
or UO_138 (O_138,N_19592,N_19964);
nand UO_139 (O_139,N_19580,N_19551);
nor UO_140 (O_140,N_19581,N_19635);
xnor UO_141 (O_141,N_19519,N_19586);
and UO_142 (O_142,N_19857,N_19945);
or UO_143 (O_143,N_19593,N_19825);
or UO_144 (O_144,N_19595,N_19879);
xnor UO_145 (O_145,N_19694,N_19863);
xor UO_146 (O_146,N_19968,N_19977);
or UO_147 (O_147,N_19917,N_19876);
xnor UO_148 (O_148,N_19669,N_19953);
nand UO_149 (O_149,N_19884,N_19502);
nor UO_150 (O_150,N_19682,N_19506);
xnor UO_151 (O_151,N_19969,N_19775);
or UO_152 (O_152,N_19763,N_19614);
nor UO_153 (O_153,N_19615,N_19844);
or UO_154 (O_154,N_19756,N_19918);
or UO_155 (O_155,N_19651,N_19697);
nor UO_156 (O_156,N_19517,N_19578);
xor UO_157 (O_157,N_19659,N_19972);
nand UO_158 (O_158,N_19511,N_19663);
nand UO_159 (O_159,N_19700,N_19573);
and UO_160 (O_160,N_19781,N_19869);
xnor UO_161 (O_161,N_19530,N_19562);
nor UO_162 (O_162,N_19559,N_19894);
and UO_163 (O_163,N_19624,N_19677);
and UO_164 (O_164,N_19789,N_19637);
and UO_165 (O_165,N_19505,N_19540);
nor UO_166 (O_166,N_19717,N_19634);
or UO_167 (O_167,N_19919,N_19725);
and UO_168 (O_168,N_19628,N_19946);
or UO_169 (O_169,N_19598,N_19670);
or UO_170 (O_170,N_19744,N_19638);
or UO_171 (O_171,N_19764,N_19647);
nor UO_172 (O_172,N_19956,N_19873);
or UO_173 (O_173,N_19703,N_19779);
xor UO_174 (O_174,N_19866,N_19709);
or UO_175 (O_175,N_19852,N_19921);
xnor UO_176 (O_176,N_19658,N_19514);
and UO_177 (O_177,N_19741,N_19716);
nor UO_178 (O_178,N_19681,N_19606);
or UO_179 (O_179,N_19589,N_19699);
and UO_180 (O_180,N_19982,N_19990);
xor UO_181 (O_181,N_19880,N_19569);
xnor UO_182 (O_182,N_19730,N_19806);
and UO_183 (O_183,N_19967,N_19553);
nand UO_184 (O_184,N_19661,N_19913);
or UO_185 (O_185,N_19874,N_19556);
xnor UO_186 (O_186,N_19561,N_19983);
nand UO_187 (O_187,N_19544,N_19688);
nand UO_188 (O_188,N_19949,N_19620);
or UO_189 (O_189,N_19633,N_19690);
or UO_190 (O_190,N_19642,N_19938);
nor UO_191 (O_191,N_19856,N_19622);
nand UO_192 (O_192,N_19795,N_19608);
nor UO_193 (O_193,N_19829,N_19673);
and UO_194 (O_194,N_19915,N_19854);
xor UO_195 (O_195,N_19837,N_19780);
nand UO_196 (O_196,N_19597,N_19654);
and UO_197 (O_197,N_19532,N_19886);
xor UO_198 (O_198,N_19958,N_19504);
nor UO_199 (O_199,N_19828,N_19889);
or UO_200 (O_200,N_19500,N_19601);
nor UO_201 (O_201,N_19845,N_19729);
and UO_202 (O_202,N_19546,N_19536);
or UO_203 (O_203,N_19772,N_19986);
xnor UO_204 (O_204,N_19936,N_19939);
or UO_205 (O_205,N_19891,N_19631);
or UO_206 (O_206,N_19603,N_19748);
and UO_207 (O_207,N_19805,N_19860);
nand UO_208 (O_208,N_19774,N_19912);
nand UO_209 (O_209,N_19590,N_19643);
nand UO_210 (O_210,N_19545,N_19881);
and UO_211 (O_211,N_19853,N_19609);
nand UO_212 (O_212,N_19927,N_19662);
nand UO_213 (O_213,N_19515,N_19518);
xnor UO_214 (O_214,N_19817,N_19679);
xnor UO_215 (O_215,N_19686,N_19978);
nand UO_216 (O_216,N_19509,N_19925);
xnor UO_217 (O_217,N_19512,N_19527);
xor UO_218 (O_218,N_19636,N_19911);
nor UO_219 (O_219,N_19711,N_19841);
and UO_220 (O_220,N_19846,N_19930);
nor UO_221 (O_221,N_19842,N_19791);
xnor UO_222 (O_222,N_19850,N_19947);
nor UO_223 (O_223,N_19718,N_19596);
xnor UO_224 (O_224,N_19807,N_19762);
nor UO_225 (O_225,N_19831,N_19528);
or UO_226 (O_226,N_19834,N_19652);
xor UO_227 (O_227,N_19794,N_19808);
or UO_228 (O_228,N_19908,N_19903);
or UO_229 (O_229,N_19970,N_19557);
xnor UO_230 (O_230,N_19671,N_19520);
xnor UO_231 (O_231,N_19714,N_19713);
nand UO_232 (O_232,N_19813,N_19888);
and UO_233 (O_233,N_19957,N_19680);
or UO_234 (O_234,N_19826,N_19804);
nor UO_235 (O_235,N_19740,N_19705);
and UO_236 (O_236,N_19878,N_19811);
or UO_237 (O_237,N_19870,N_19503);
nor UO_238 (O_238,N_19749,N_19538);
and UO_239 (O_239,N_19942,N_19840);
and UO_240 (O_240,N_19766,N_19758);
nor UO_241 (O_241,N_19591,N_19951);
nand UO_242 (O_242,N_19944,N_19767);
and UO_243 (O_243,N_19865,N_19909);
and UO_244 (O_244,N_19838,N_19922);
and UO_245 (O_245,N_19715,N_19728);
or UO_246 (O_246,N_19771,N_19929);
nand UO_247 (O_247,N_19793,N_19931);
nor UO_248 (O_248,N_19920,N_19577);
and UO_249 (O_249,N_19724,N_19668);
xnor UO_250 (O_250,N_19928,N_19768);
nor UO_251 (O_251,N_19731,N_19722);
xnor UO_252 (O_252,N_19771,N_19913);
nor UO_253 (O_253,N_19851,N_19716);
or UO_254 (O_254,N_19503,N_19536);
xnor UO_255 (O_255,N_19912,N_19858);
or UO_256 (O_256,N_19900,N_19894);
nand UO_257 (O_257,N_19522,N_19962);
nand UO_258 (O_258,N_19664,N_19600);
and UO_259 (O_259,N_19600,N_19766);
nand UO_260 (O_260,N_19518,N_19663);
nand UO_261 (O_261,N_19965,N_19573);
xnor UO_262 (O_262,N_19729,N_19640);
nand UO_263 (O_263,N_19580,N_19790);
nand UO_264 (O_264,N_19984,N_19850);
nand UO_265 (O_265,N_19783,N_19619);
xor UO_266 (O_266,N_19771,N_19720);
and UO_267 (O_267,N_19571,N_19583);
or UO_268 (O_268,N_19806,N_19982);
nor UO_269 (O_269,N_19684,N_19650);
xor UO_270 (O_270,N_19615,N_19743);
or UO_271 (O_271,N_19508,N_19890);
and UO_272 (O_272,N_19763,N_19925);
xor UO_273 (O_273,N_19772,N_19989);
nor UO_274 (O_274,N_19641,N_19787);
xnor UO_275 (O_275,N_19710,N_19946);
and UO_276 (O_276,N_19962,N_19577);
nand UO_277 (O_277,N_19587,N_19811);
or UO_278 (O_278,N_19562,N_19715);
or UO_279 (O_279,N_19900,N_19946);
and UO_280 (O_280,N_19857,N_19697);
and UO_281 (O_281,N_19528,N_19766);
nor UO_282 (O_282,N_19869,N_19672);
nor UO_283 (O_283,N_19989,N_19508);
and UO_284 (O_284,N_19572,N_19791);
nor UO_285 (O_285,N_19905,N_19511);
xor UO_286 (O_286,N_19907,N_19525);
xor UO_287 (O_287,N_19582,N_19913);
nor UO_288 (O_288,N_19703,N_19885);
nand UO_289 (O_289,N_19975,N_19857);
nand UO_290 (O_290,N_19694,N_19722);
nor UO_291 (O_291,N_19992,N_19758);
and UO_292 (O_292,N_19687,N_19637);
nor UO_293 (O_293,N_19723,N_19946);
or UO_294 (O_294,N_19940,N_19915);
and UO_295 (O_295,N_19898,N_19682);
nand UO_296 (O_296,N_19609,N_19767);
xor UO_297 (O_297,N_19853,N_19780);
nor UO_298 (O_298,N_19911,N_19881);
nor UO_299 (O_299,N_19894,N_19687);
nor UO_300 (O_300,N_19549,N_19781);
or UO_301 (O_301,N_19931,N_19687);
or UO_302 (O_302,N_19637,N_19832);
nand UO_303 (O_303,N_19575,N_19798);
xor UO_304 (O_304,N_19729,N_19746);
xor UO_305 (O_305,N_19786,N_19817);
xnor UO_306 (O_306,N_19544,N_19902);
or UO_307 (O_307,N_19666,N_19738);
nor UO_308 (O_308,N_19649,N_19926);
or UO_309 (O_309,N_19612,N_19587);
nand UO_310 (O_310,N_19886,N_19602);
nand UO_311 (O_311,N_19673,N_19868);
nand UO_312 (O_312,N_19511,N_19753);
xor UO_313 (O_313,N_19657,N_19929);
xnor UO_314 (O_314,N_19604,N_19911);
xnor UO_315 (O_315,N_19775,N_19705);
nand UO_316 (O_316,N_19837,N_19644);
and UO_317 (O_317,N_19913,N_19961);
and UO_318 (O_318,N_19845,N_19963);
xor UO_319 (O_319,N_19820,N_19668);
or UO_320 (O_320,N_19941,N_19628);
nand UO_321 (O_321,N_19993,N_19889);
nor UO_322 (O_322,N_19517,N_19804);
xor UO_323 (O_323,N_19633,N_19931);
or UO_324 (O_324,N_19908,N_19886);
nand UO_325 (O_325,N_19562,N_19819);
or UO_326 (O_326,N_19724,N_19680);
xnor UO_327 (O_327,N_19989,N_19688);
nor UO_328 (O_328,N_19857,N_19894);
nor UO_329 (O_329,N_19696,N_19963);
nand UO_330 (O_330,N_19965,N_19741);
or UO_331 (O_331,N_19703,N_19556);
nand UO_332 (O_332,N_19993,N_19673);
nor UO_333 (O_333,N_19751,N_19843);
nand UO_334 (O_334,N_19712,N_19608);
nand UO_335 (O_335,N_19882,N_19905);
nor UO_336 (O_336,N_19866,N_19996);
xnor UO_337 (O_337,N_19983,N_19940);
nand UO_338 (O_338,N_19546,N_19871);
nand UO_339 (O_339,N_19631,N_19920);
or UO_340 (O_340,N_19658,N_19569);
xnor UO_341 (O_341,N_19865,N_19720);
xnor UO_342 (O_342,N_19803,N_19741);
xnor UO_343 (O_343,N_19549,N_19773);
or UO_344 (O_344,N_19595,N_19913);
nand UO_345 (O_345,N_19757,N_19866);
and UO_346 (O_346,N_19876,N_19996);
nand UO_347 (O_347,N_19747,N_19816);
and UO_348 (O_348,N_19520,N_19867);
nand UO_349 (O_349,N_19923,N_19936);
or UO_350 (O_350,N_19921,N_19527);
nand UO_351 (O_351,N_19901,N_19614);
or UO_352 (O_352,N_19574,N_19791);
nor UO_353 (O_353,N_19572,N_19948);
and UO_354 (O_354,N_19862,N_19750);
nand UO_355 (O_355,N_19809,N_19548);
nor UO_356 (O_356,N_19939,N_19910);
and UO_357 (O_357,N_19852,N_19607);
xor UO_358 (O_358,N_19557,N_19968);
and UO_359 (O_359,N_19515,N_19826);
or UO_360 (O_360,N_19838,N_19790);
nand UO_361 (O_361,N_19661,N_19649);
or UO_362 (O_362,N_19787,N_19749);
xnor UO_363 (O_363,N_19800,N_19883);
xor UO_364 (O_364,N_19666,N_19764);
nand UO_365 (O_365,N_19962,N_19940);
xor UO_366 (O_366,N_19982,N_19857);
xor UO_367 (O_367,N_19614,N_19981);
nand UO_368 (O_368,N_19806,N_19516);
xor UO_369 (O_369,N_19999,N_19977);
xor UO_370 (O_370,N_19818,N_19848);
nand UO_371 (O_371,N_19878,N_19567);
and UO_372 (O_372,N_19641,N_19881);
xor UO_373 (O_373,N_19936,N_19867);
xor UO_374 (O_374,N_19556,N_19667);
xnor UO_375 (O_375,N_19955,N_19873);
nand UO_376 (O_376,N_19730,N_19989);
nor UO_377 (O_377,N_19638,N_19842);
and UO_378 (O_378,N_19552,N_19676);
or UO_379 (O_379,N_19571,N_19537);
nand UO_380 (O_380,N_19651,N_19566);
xnor UO_381 (O_381,N_19861,N_19768);
or UO_382 (O_382,N_19578,N_19799);
xor UO_383 (O_383,N_19814,N_19847);
nand UO_384 (O_384,N_19617,N_19894);
nand UO_385 (O_385,N_19553,N_19900);
or UO_386 (O_386,N_19508,N_19799);
nand UO_387 (O_387,N_19756,N_19612);
or UO_388 (O_388,N_19962,N_19750);
nor UO_389 (O_389,N_19803,N_19975);
nand UO_390 (O_390,N_19630,N_19922);
and UO_391 (O_391,N_19875,N_19986);
xor UO_392 (O_392,N_19546,N_19658);
nand UO_393 (O_393,N_19676,N_19530);
nor UO_394 (O_394,N_19757,N_19802);
or UO_395 (O_395,N_19953,N_19782);
nor UO_396 (O_396,N_19649,N_19556);
nand UO_397 (O_397,N_19683,N_19513);
and UO_398 (O_398,N_19862,N_19626);
xnor UO_399 (O_399,N_19556,N_19946);
or UO_400 (O_400,N_19887,N_19912);
nand UO_401 (O_401,N_19712,N_19619);
nand UO_402 (O_402,N_19518,N_19994);
nor UO_403 (O_403,N_19950,N_19969);
nor UO_404 (O_404,N_19985,N_19797);
nor UO_405 (O_405,N_19756,N_19549);
nor UO_406 (O_406,N_19950,N_19667);
nor UO_407 (O_407,N_19695,N_19939);
or UO_408 (O_408,N_19827,N_19882);
or UO_409 (O_409,N_19766,N_19686);
nand UO_410 (O_410,N_19520,N_19827);
nand UO_411 (O_411,N_19735,N_19536);
nand UO_412 (O_412,N_19721,N_19910);
xnor UO_413 (O_413,N_19966,N_19524);
nand UO_414 (O_414,N_19585,N_19569);
and UO_415 (O_415,N_19756,N_19770);
nand UO_416 (O_416,N_19592,N_19780);
nor UO_417 (O_417,N_19788,N_19790);
xnor UO_418 (O_418,N_19631,N_19957);
nand UO_419 (O_419,N_19680,N_19747);
nor UO_420 (O_420,N_19784,N_19788);
xor UO_421 (O_421,N_19858,N_19811);
nor UO_422 (O_422,N_19729,N_19942);
nand UO_423 (O_423,N_19545,N_19918);
nand UO_424 (O_424,N_19665,N_19683);
xor UO_425 (O_425,N_19723,N_19601);
nand UO_426 (O_426,N_19522,N_19722);
xor UO_427 (O_427,N_19855,N_19910);
xor UO_428 (O_428,N_19999,N_19908);
and UO_429 (O_429,N_19936,N_19518);
nand UO_430 (O_430,N_19794,N_19978);
and UO_431 (O_431,N_19736,N_19796);
xnor UO_432 (O_432,N_19663,N_19539);
xor UO_433 (O_433,N_19677,N_19939);
xor UO_434 (O_434,N_19508,N_19999);
nor UO_435 (O_435,N_19961,N_19734);
or UO_436 (O_436,N_19733,N_19656);
or UO_437 (O_437,N_19761,N_19731);
or UO_438 (O_438,N_19744,N_19554);
nor UO_439 (O_439,N_19904,N_19724);
or UO_440 (O_440,N_19644,N_19876);
and UO_441 (O_441,N_19680,N_19734);
xnor UO_442 (O_442,N_19613,N_19788);
nor UO_443 (O_443,N_19949,N_19673);
xnor UO_444 (O_444,N_19734,N_19606);
and UO_445 (O_445,N_19526,N_19939);
nand UO_446 (O_446,N_19941,N_19972);
nor UO_447 (O_447,N_19575,N_19659);
nor UO_448 (O_448,N_19819,N_19768);
nor UO_449 (O_449,N_19743,N_19719);
xor UO_450 (O_450,N_19685,N_19977);
xnor UO_451 (O_451,N_19937,N_19839);
or UO_452 (O_452,N_19503,N_19710);
and UO_453 (O_453,N_19829,N_19657);
or UO_454 (O_454,N_19959,N_19560);
and UO_455 (O_455,N_19797,N_19546);
nor UO_456 (O_456,N_19774,N_19624);
xnor UO_457 (O_457,N_19685,N_19761);
and UO_458 (O_458,N_19835,N_19708);
or UO_459 (O_459,N_19661,N_19998);
and UO_460 (O_460,N_19692,N_19736);
or UO_461 (O_461,N_19758,N_19977);
nor UO_462 (O_462,N_19791,N_19726);
or UO_463 (O_463,N_19857,N_19511);
and UO_464 (O_464,N_19977,N_19768);
xnor UO_465 (O_465,N_19818,N_19744);
nor UO_466 (O_466,N_19554,N_19658);
and UO_467 (O_467,N_19770,N_19745);
nor UO_468 (O_468,N_19705,N_19642);
nor UO_469 (O_469,N_19987,N_19797);
nand UO_470 (O_470,N_19762,N_19579);
or UO_471 (O_471,N_19928,N_19715);
or UO_472 (O_472,N_19963,N_19901);
xor UO_473 (O_473,N_19536,N_19528);
xor UO_474 (O_474,N_19934,N_19600);
nor UO_475 (O_475,N_19656,N_19884);
or UO_476 (O_476,N_19951,N_19688);
or UO_477 (O_477,N_19501,N_19546);
and UO_478 (O_478,N_19762,N_19745);
or UO_479 (O_479,N_19739,N_19836);
nand UO_480 (O_480,N_19932,N_19896);
and UO_481 (O_481,N_19877,N_19917);
or UO_482 (O_482,N_19593,N_19535);
nand UO_483 (O_483,N_19632,N_19795);
nor UO_484 (O_484,N_19799,N_19830);
xnor UO_485 (O_485,N_19875,N_19621);
and UO_486 (O_486,N_19620,N_19933);
or UO_487 (O_487,N_19983,N_19749);
nor UO_488 (O_488,N_19880,N_19749);
xor UO_489 (O_489,N_19564,N_19598);
and UO_490 (O_490,N_19561,N_19874);
or UO_491 (O_491,N_19521,N_19702);
xor UO_492 (O_492,N_19905,N_19791);
xor UO_493 (O_493,N_19847,N_19779);
and UO_494 (O_494,N_19891,N_19740);
xor UO_495 (O_495,N_19691,N_19938);
nand UO_496 (O_496,N_19737,N_19587);
nand UO_497 (O_497,N_19889,N_19573);
nand UO_498 (O_498,N_19955,N_19934);
xnor UO_499 (O_499,N_19793,N_19884);
nor UO_500 (O_500,N_19597,N_19839);
or UO_501 (O_501,N_19963,N_19640);
nand UO_502 (O_502,N_19935,N_19763);
nand UO_503 (O_503,N_19636,N_19985);
or UO_504 (O_504,N_19708,N_19867);
nand UO_505 (O_505,N_19782,N_19564);
nor UO_506 (O_506,N_19509,N_19762);
or UO_507 (O_507,N_19588,N_19913);
nand UO_508 (O_508,N_19535,N_19629);
xor UO_509 (O_509,N_19650,N_19821);
nor UO_510 (O_510,N_19747,N_19858);
xnor UO_511 (O_511,N_19675,N_19584);
and UO_512 (O_512,N_19586,N_19919);
xor UO_513 (O_513,N_19721,N_19926);
nor UO_514 (O_514,N_19937,N_19996);
nand UO_515 (O_515,N_19778,N_19797);
and UO_516 (O_516,N_19948,N_19917);
nand UO_517 (O_517,N_19952,N_19794);
nand UO_518 (O_518,N_19948,N_19509);
xnor UO_519 (O_519,N_19866,N_19666);
or UO_520 (O_520,N_19620,N_19564);
or UO_521 (O_521,N_19985,N_19556);
xnor UO_522 (O_522,N_19707,N_19616);
nor UO_523 (O_523,N_19800,N_19905);
xnor UO_524 (O_524,N_19749,N_19607);
xor UO_525 (O_525,N_19597,N_19999);
nand UO_526 (O_526,N_19549,N_19501);
xnor UO_527 (O_527,N_19653,N_19929);
nand UO_528 (O_528,N_19907,N_19809);
or UO_529 (O_529,N_19710,N_19938);
or UO_530 (O_530,N_19573,N_19803);
and UO_531 (O_531,N_19591,N_19608);
nand UO_532 (O_532,N_19914,N_19866);
xnor UO_533 (O_533,N_19697,N_19610);
xor UO_534 (O_534,N_19754,N_19839);
or UO_535 (O_535,N_19999,N_19814);
nor UO_536 (O_536,N_19827,N_19616);
nand UO_537 (O_537,N_19837,N_19586);
nand UO_538 (O_538,N_19922,N_19852);
nor UO_539 (O_539,N_19878,N_19932);
nand UO_540 (O_540,N_19737,N_19947);
xnor UO_541 (O_541,N_19558,N_19764);
nand UO_542 (O_542,N_19826,N_19843);
and UO_543 (O_543,N_19934,N_19662);
nor UO_544 (O_544,N_19929,N_19529);
xnor UO_545 (O_545,N_19635,N_19887);
or UO_546 (O_546,N_19980,N_19877);
xor UO_547 (O_547,N_19660,N_19825);
nand UO_548 (O_548,N_19755,N_19905);
or UO_549 (O_549,N_19533,N_19831);
and UO_550 (O_550,N_19979,N_19990);
xor UO_551 (O_551,N_19653,N_19639);
or UO_552 (O_552,N_19626,N_19621);
or UO_553 (O_553,N_19986,N_19823);
xnor UO_554 (O_554,N_19734,N_19743);
and UO_555 (O_555,N_19549,N_19771);
xor UO_556 (O_556,N_19579,N_19765);
and UO_557 (O_557,N_19835,N_19666);
nor UO_558 (O_558,N_19816,N_19960);
xor UO_559 (O_559,N_19794,N_19573);
nor UO_560 (O_560,N_19912,N_19869);
nor UO_561 (O_561,N_19628,N_19653);
nand UO_562 (O_562,N_19697,N_19974);
and UO_563 (O_563,N_19683,N_19666);
nor UO_564 (O_564,N_19986,N_19919);
and UO_565 (O_565,N_19659,N_19712);
nand UO_566 (O_566,N_19961,N_19931);
nor UO_567 (O_567,N_19663,N_19531);
and UO_568 (O_568,N_19715,N_19669);
and UO_569 (O_569,N_19980,N_19616);
and UO_570 (O_570,N_19845,N_19663);
and UO_571 (O_571,N_19623,N_19713);
nand UO_572 (O_572,N_19588,N_19934);
nand UO_573 (O_573,N_19973,N_19572);
and UO_574 (O_574,N_19554,N_19661);
and UO_575 (O_575,N_19907,N_19979);
nor UO_576 (O_576,N_19965,N_19933);
and UO_577 (O_577,N_19877,N_19710);
xor UO_578 (O_578,N_19543,N_19621);
and UO_579 (O_579,N_19988,N_19906);
nor UO_580 (O_580,N_19558,N_19897);
or UO_581 (O_581,N_19640,N_19628);
nor UO_582 (O_582,N_19801,N_19687);
and UO_583 (O_583,N_19890,N_19710);
and UO_584 (O_584,N_19698,N_19639);
nand UO_585 (O_585,N_19896,N_19929);
nor UO_586 (O_586,N_19946,N_19644);
and UO_587 (O_587,N_19730,N_19521);
nand UO_588 (O_588,N_19881,N_19850);
nand UO_589 (O_589,N_19941,N_19581);
and UO_590 (O_590,N_19668,N_19718);
and UO_591 (O_591,N_19742,N_19997);
or UO_592 (O_592,N_19542,N_19514);
or UO_593 (O_593,N_19908,N_19835);
and UO_594 (O_594,N_19521,N_19667);
nor UO_595 (O_595,N_19628,N_19684);
xnor UO_596 (O_596,N_19959,N_19966);
or UO_597 (O_597,N_19557,N_19519);
or UO_598 (O_598,N_19522,N_19730);
nand UO_599 (O_599,N_19575,N_19569);
and UO_600 (O_600,N_19865,N_19619);
nand UO_601 (O_601,N_19924,N_19510);
or UO_602 (O_602,N_19989,N_19888);
or UO_603 (O_603,N_19941,N_19752);
nor UO_604 (O_604,N_19897,N_19839);
and UO_605 (O_605,N_19984,N_19638);
xnor UO_606 (O_606,N_19709,N_19968);
nor UO_607 (O_607,N_19829,N_19579);
nand UO_608 (O_608,N_19843,N_19615);
nand UO_609 (O_609,N_19711,N_19897);
and UO_610 (O_610,N_19557,N_19937);
and UO_611 (O_611,N_19580,N_19650);
nor UO_612 (O_612,N_19778,N_19894);
nand UO_613 (O_613,N_19566,N_19753);
nor UO_614 (O_614,N_19706,N_19840);
or UO_615 (O_615,N_19703,N_19719);
or UO_616 (O_616,N_19819,N_19685);
nor UO_617 (O_617,N_19793,N_19920);
nand UO_618 (O_618,N_19978,N_19879);
nor UO_619 (O_619,N_19928,N_19523);
and UO_620 (O_620,N_19714,N_19914);
or UO_621 (O_621,N_19552,N_19986);
xor UO_622 (O_622,N_19567,N_19867);
xnor UO_623 (O_623,N_19787,N_19616);
nand UO_624 (O_624,N_19954,N_19903);
nor UO_625 (O_625,N_19945,N_19515);
or UO_626 (O_626,N_19683,N_19714);
nor UO_627 (O_627,N_19680,N_19508);
xnor UO_628 (O_628,N_19771,N_19551);
xnor UO_629 (O_629,N_19996,N_19739);
nand UO_630 (O_630,N_19518,N_19513);
xor UO_631 (O_631,N_19897,N_19886);
and UO_632 (O_632,N_19996,N_19754);
nor UO_633 (O_633,N_19664,N_19913);
nor UO_634 (O_634,N_19916,N_19524);
and UO_635 (O_635,N_19729,N_19733);
nor UO_636 (O_636,N_19593,N_19720);
nor UO_637 (O_637,N_19605,N_19741);
nand UO_638 (O_638,N_19687,N_19551);
nor UO_639 (O_639,N_19900,N_19693);
and UO_640 (O_640,N_19689,N_19613);
and UO_641 (O_641,N_19708,N_19992);
and UO_642 (O_642,N_19794,N_19839);
xor UO_643 (O_643,N_19672,N_19678);
nand UO_644 (O_644,N_19642,N_19671);
nand UO_645 (O_645,N_19853,N_19998);
xnor UO_646 (O_646,N_19875,N_19810);
nor UO_647 (O_647,N_19847,N_19981);
nand UO_648 (O_648,N_19658,N_19856);
or UO_649 (O_649,N_19733,N_19731);
xnor UO_650 (O_650,N_19682,N_19915);
nand UO_651 (O_651,N_19546,N_19518);
and UO_652 (O_652,N_19675,N_19945);
xor UO_653 (O_653,N_19790,N_19950);
nand UO_654 (O_654,N_19728,N_19581);
or UO_655 (O_655,N_19507,N_19597);
nor UO_656 (O_656,N_19501,N_19694);
or UO_657 (O_657,N_19873,N_19875);
nor UO_658 (O_658,N_19954,N_19823);
xnor UO_659 (O_659,N_19607,N_19841);
xnor UO_660 (O_660,N_19979,N_19626);
and UO_661 (O_661,N_19974,N_19729);
and UO_662 (O_662,N_19959,N_19854);
nor UO_663 (O_663,N_19834,N_19942);
and UO_664 (O_664,N_19645,N_19687);
xor UO_665 (O_665,N_19772,N_19848);
nor UO_666 (O_666,N_19604,N_19678);
nor UO_667 (O_667,N_19596,N_19573);
or UO_668 (O_668,N_19753,N_19952);
xor UO_669 (O_669,N_19534,N_19636);
and UO_670 (O_670,N_19865,N_19732);
xnor UO_671 (O_671,N_19806,N_19923);
nor UO_672 (O_672,N_19788,N_19899);
nor UO_673 (O_673,N_19689,N_19647);
nor UO_674 (O_674,N_19888,N_19599);
and UO_675 (O_675,N_19704,N_19998);
or UO_676 (O_676,N_19782,N_19722);
xor UO_677 (O_677,N_19865,N_19920);
or UO_678 (O_678,N_19904,N_19680);
nor UO_679 (O_679,N_19579,N_19664);
nand UO_680 (O_680,N_19709,N_19764);
or UO_681 (O_681,N_19529,N_19915);
nand UO_682 (O_682,N_19679,N_19858);
nand UO_683 (O_683,N_19753,N_19831);
and UO_684 (O_684,N_19933,N_19660);
nor UO_685 (O_685,N_19647,N_19922);
or UO_686 (O_686,N_19994,N_19608);
nor UO_687 (O_687,N_19670,N_19638);
or UO_688 (O_688,N_19730,N_19578);
xnor UO_689 (O_689,N_19875,N_19706);
or UO_690 (O_690,N_19808,N_19976);
nand UO_691 (O_691,N_19898,N_19848);
or UO_692 (O_692,N_19676,N_19775);
nor UO_693 (O_693,N_19900,N_19919);
nor UO_694 (O_694,N_19513,N_19865);
and UO_695 (O_695,N_19860,N_19560);
xor UO_696 (O_696,N_19895,N_19945);
xor UO_697 (O_697,N_19730,N_19620);
xor UO_698 (O_698,N_19616,N_19779);
nor UO_699 (O_699,N_19754,N_19593);
nor UO_700 (O_700,N_19909,N_19578);
nor UO_701 (O_701,N_19634,N_19787);
or UO_702 (O_702,N_19996,N_19975);
nand UO_703 (O_703,N_19720,N_19950);
nand UO_704 (O_704,N_19652,N_19535);
nand UO_705 (O_705,N_19906,N_19843);
nor UO_706 (O_706,N_19881,N_19778);
nor UO_707 (O_707,N_19697,N_19814);
nor UO_708 (O_708,N_19702,N_19739);
xnor UO_709 (O_709,N_19566,N_19598);
or UO_710 (O_710,N_19920,N_19524);
nor UO_711 (O_711,N_19998,N_19931);
and UO_712 (O_712,N_19819,N_19907);
xnor UO_713 (O_713,N_19855,N_19514);
xor UO_714 (O_714,N_19757,N_19981);
xor UO_715 (O_715,N_19853,N_19714);
xor UO_716 (O_716,N_19658,N_19820);
xor UO_717 (O_717,N_19983,N_19618);
nand UO_718 (O_718,N_19759,N_19721);
nor UO_719 (O_719,N_19990,N_19746);
and UO_720 (O_720,N_19685,N_19727);
nor UO_721 (O_721,N_19769,N_19759);
or UO_722 (O_722,N_19594,N_19697);
or UO_723 (O_723,N_19967,N_19885);
nor UO_724 (O_724,N_19988,N_19907);
nor UO_725 (O_725,N_19632,N_19527);
or UO_726 (O_726,N_19512,N_19905);
and UO_727 (O_727,N_19725,N_19649);
nor UO_728 (O_728,N_19534,N_19646);
nand UO_729 (O_729,N_19925,N_19641);
and UO_730 (O_730,N_19650,N_19748);
nand UO_731 (O_731,N_19749,N_19544);
or UO_732 (O_732,N_19903,N_19727);
and UO_733 (O_733,N_19635,N_19698);
nand UO_734 (O_734,N_19954,N_19867);
nor UO_735 (O_735,N_19921,N_19748);
nand UO_736 (O_736,N_19646,N_19852);
and UO_737 (O_737,N_19553,N_19721);
nor UO_738 (O_738,N_19971,N_19583);
nand UO_739 (O_739,N_19832,N_19827);
or UO_740 (O_740,N_19639,N_19757);
xnor UO_741 (O_741,N_19525,N_19694);
nand UO_742 (O_742,N_19949,N_19951);
xnor UO_743 (O_743,N_19756,N_19734);
nor UO_744 (O_744,N_19694,N_19743);
and UO_745 (O_745,N_19609,N_19914);
xor UO_746 (O_746,N_19855,N_19812);
or UO_747 (O_747,N_19947,N_19990);
xor UO_748 (O_748,N_19641,N_19612);
nor UO_749 (O_749,N_19581,N_19792);
nor UO_750 (O_750,N_19693,N_19628);
or UO_751 (O_751,N_19630,N_19860);
and UO_752 (O_752,N_19995,N_19834);
and UO_753 (O_753,N_19923,N_19653);
nand UO_754 (O_754,N_19813,N_19666);
and UO_755 (O_755,N_19736,N_19562);
and UO_756 (O_756,N_19730,N_19836);
or UO_757 (O_757,N_19632,N_19780);
xor UO_758 (O_758,N_19883,N_19690);
nand UO_759 (O_759,N_19580,N_19577);
or UO_760 (O_760,N_19883,N_19912);
xnor UO_761 (O_761,N_19735,N_19632);
and UO_762 (O_762,N_19543,N_19525);
nor UO_763 (O_763,N_19640,N_19611);
xnor UO_764 (O_764,N_19766,N_19927);
xor UO_765 (O_765,N_19715,N_19758);
xor UO_766 (O_766,N_19549,N_19923);
and UO_767 (O_767,N_19627,N_19965);
xor UO_768 (O_768,N_19948,N_19533);
or UO_769 (O_769,N_19806,N_19600);
or UO_770 (O_770,N_19864,N_19511);
nor UO_771 (O_771,N_19835,N_19967);
or UO_772 (O_772,N_19638,N_19716);
and UO_773 (O_773,N_19864,N_19952);
nor UO_774 (O_774,N_19560,N_19983);
or UO_775 (O_775,N_19551,N_19987);
nor UO_776 (O_776,N_19648,N_19826);
xnor UO_777 (O_777,N_19695,N_19804);
or UO_778 (O_778,N_19813,N_19896);
nand UO_779 (O_779,N_19577,N_19732);
or UO_780 (O_780,N_19535,N_19613);
xor UO_781 (O_781,N_19564,N_19636);
nor UO_782 (O_782,N_19869,N_19618);
nor UO_783 (O_783,N_19595,N_19600);
and UO_784 (O_784,N_19892,N_19870);
or UO_785 (O_785,N_19875,N_19772);
or UO_786 (O_786,N_19545,N_19944);
nand UO_787 (O_787,N_19766,N_19663);
xor UO_788 (O_788,N_19719,N_19705);
xnor UO_789 (O_789,N_19716,N_19721);
or UO_790 (O_790,N_19661,N_19908);
or UO_791 (O_791,N_19519,N_19845);
nor UO_792 (O_792,N_19999,N_19891);
or UO_793 (O_793,N_19838,N_19956);
and UO_794 (O_794,N_19544,N_19527);
or UO_795 (O_795,N_19513,N_19863);
and UO_796 (O_796,N_19582,N_19675);
nand UO_797 (O_797,N_19842,N_19585);
nor UO_798 (O_798,N_19947,N_19741);
nor UO_799 (O_799,N_19975,N_19575);
nor UO_800 (O_800,N_19503,N_19809);
xnor UO_801 (O_801,N_19578,N_19553);
nor UO_802 (O_802,N_19932,N_19752);
or UO_803 (O_803,N_19696,N_19877);
nor UO_804 (O_804,N_19642,N_19646);
nand UO_805 (O_805,N_19767,N_19763);
xnor UO_806 (O_806,N_19896,N_19532);
nor UO_807 (O_807,N_19521,N_19756);
nand UO_808 (O_808,N_19638,N_19522);
and UO_809 (O_809,N_19895,N_19961);
xor UO_810 (O_810,N_19544,N_19682);
xor UO_811 (O_811,N_19590,N_19514);
or UO_812 (O_812,N_19583,N_19578);
or UO_813 (O_813,N_19617,N_19793);
xnor UO_814 (O_814,N_19911,N_19539);
nand UO_815 (O_815,N_19567,N_19758);
and UO_816 (O_816,N_19512,N_19712);
nand UO_817 (O_817,N_19719,N_19529);
or UO_818 (O_818,N_19863,N_19976);
nand UO_819 (O_819,N_19778,N_19702);
or UO_820 (O_820,N_19595,N_19789);
nor UO_821 (O_821,N_19627,N_19873);
nor UO_822 (O_822,N_19572,N_19780);
or UO_823 (O_823,N_19994,N_19961);
xnor UO_824 (O_824,N_19876,N_19739);
nand UO_825 (O_825,N_19717,N_19600);
xnor UO_826 (O_826,N_19870,N_19615);
nor UO_827 (O_827,N_19700,N_19713);
or UO_828 (O_828,N_19687,N_19875);
xnor UO_829 (O_829,N_19977,N_19604);
nor UO_830 (O_830,N_19889,N_19702);
nand UO_831 (O_831,N_19688,N_19764);
and UO_832 (O_832,N_19697,N_19542);
or UO_833 (O_833,N_19679,N_19693);
nand UO_834 (O_834,N_19569,N_19662);
xnor UO_835 (O_835,N_19908,N_19560);
nand UO_836 (O_836,N_19837,N_19960);
or UO_837 (O_837,N_19790,N_19994);
xor UO_838 (O_838,N_19735,N_19700);
xor UO_839 (O_839,N_19909,N_19518);
or UO_840 (O_840,N_19671,N_19570);
nand UO_841 (O_841,N_19519,N_19572);
nand UO_842 (O_842,N_19763,N_19908);
nand UO_843 (O_843,N_19933,N_19905);
nor UO_844 (O_844,N_19720,N_19981);
xor UO_845 (O_845,N_19707,N_19569);
and UO_846 (O_846,N_19696,N_19516);
or UO_847 (O_847,N_19663,N_19728);
or UO_848 (O_848,N_19717,N_19880);
or UO_849 (O_849,N_19713,N_19894);
nor UO_850 (O_850,N_19926,N_19955);
and UO_851 (O_851,N_19697,N_19739);
and UO_852 (O_852,N_19988,N_19664);
or UO_853 (O_853,N_19850,N_19646);
xor UO_854 (O_854,N_19954,N_19984);
and UO_855 (O_855,N_19714,N_19934);
and UO_856 (O_856,N_19748,N_19974);
nand UO_857 (O_857,N_19805,N_19598);
nand UO_858 (O_858,N_19793,N_19953);
nor UO_859 (O_859,N_19955,N_19742);
nand UO_860 (O_860,N_19525,N_19635);
xnor UO_861 (O_861,N_19580,N_19570);
or UO_862 (O_862,N_19931,N_19500);
nand UO_863 (O_863,N_19649,N_19637);
xnor UO_864 (O_864,N_19978,N_19557);
or UO_865 (O_865,N_19941,N_19537);
and UO_866 (O_866,N_19791,N_19771);
xor UO_867 (O_867,N_19759,N_19541);
nand UO_868 (O_868,N_19573,N_19648);
nor UO_869 (O_869,N_19502,N_19726);
nor UO_870 (O_870,N_19700,N_19696);
xnor UO_871 (O_871,N_19867,N_19982);
and UO_872 (O_872,N_19506,N_19520);
nor UO_873 (O_873,N_19650,N_19953);
nand UO_874 (O_874,N_19737,N_19790);
or UO_875 (O_875,N_19689,N_19850);
xnor UO_876 (O_876,N_19914,N_19861);
nor UO_877 (O_877,N_19727,N_19680);
xnor UO_878 (O_878,N_19854,N_19980);
xor UO_879 (O_879,N_19641,N_19950);
nor UO_880 (O_880,N_19703,N_19623);
and UO_881 (O_881,N_19781,N_19966);
nand UO_882 (O_882,N_19748,N_19882);
nor UO_883 (O_883,N_19794,N_19948);
xnor UO_884 (O_884,N_19506,N_19641);
and UO_885 (O_885,N_19538,N_19790);
xor UO_886 (O_886,N_19765,N_19834);
nor UO_887 (O_887,N_19581,N_19922);
or UO_888 (O_888,N_19506,N_19976);
nand UO_889 (O_889,N_19777,N_19956);
nand UO_890 (O_890,N_19706,N_19611);
or UO_891 (O_891,N_19636,N_19921);
or UO_892 (O_892,N_19803,N_19911);
nor UO_893 (O_893,N_19766,N_19515);
nand UO_894 (O_894,N_19680,N_19520);
or UO_895 (O_895,N_19600,N_19753);
xor UO_896 (O_896,N_19771,N_19807);
xnor UO_897 (O_897,N_19600,N_19864);
xnor UO_898 (O_898,N_19975,N_19771);
nor UO_899 (O_899,N_19831,N_19986);
or UO_900 (O_900,N_19717,N_19921);
and UO_901 (O_901,N_19706,N_19854);
or UO_902 (O_902,N_19803,N_19560);
nand UO_903 (O_903,N_19567,N_19917);
or UO_904 (O_904,N_19507,N_19741);
and UO_905 (O_905,N_19824,N_19869);
and UO_906 (O_906,N_19631,N_19701);
and UO_907 (O_907,N_19766,N_19920);
xnor UO_908 (O_908,N_19681,N_19992);
nand UO_909 (O_909,N_19909,N_19690);
nor UO_910 (O_910,N_19973,N_19555);
or UO_911 (O_911,N_19900,N_19760);
and UO_912 (O_912,N_19696,N_19749);
xor UO_913 (O_913,N_19885,N_19602);
nand UO_914 (O_914,N_19905,N_19505);
or UO_915 (O_915,N_19826,N_19751);
and UO_916 (O_916,N_19969,N_19977);
nand UO_917 (O_917,N_19762,N_19515);
or UO_918 (O_918,N_19912,N_19659);
nand UO_919 (O_919,N_19978,N_19913);
nor UO_920 (O_920,N_19760,N_19812);
and UO_921 (O_921,N_19624,N_19884);
and UO_922 (O_922,N_19931,N_19617);
nand UO_923 (O_923,N_19739,N_19880);
xnor UO_924 (O_924,N_19902,N_19503);
xnor UO_925 (O_925,N_19966,N_19915);
or UO_926 (O_926,N_19966,N_19542);
nand UO_927 (O_927,N_19841,N_19571);
nand UO_928 (O_928,N_19652,N_19997);
or UO_929 (O_929,N_19712,N_19686);
and UO_930 (O_930,N_19807,N_19539);
nand UO_931 (O_931,N_19613,N_19849);
nand UO_932 (O_932,N_19845,N_19501);
or UO_933 (O_933,N_19609,N_19756);
or UO_934 (O_934,N_19597,N_19941);
nand UO_935 (O_935,N_19618,N_19834);
and UO_936 (O_936,N_19830,N_19649);
and UO_937 (O_937,N_19586,N_19876);
nand UO_938 (O_938,N_19858,N_19886);
nor UO_939 (O_939,N_19612,N_19583);
and UO_940 (O_940,N_19854,N_19539);
nor UO_941 (O_941,N_19557,N_19529);
nor UO_942 (O_942,N_19622,N_19640);
or UO_943 (O_943,N_19848,N_19512);
nor UO_944 (O_944,N_19776,N_19654);
nor UO_945 (O_945,N_19687,N_19993);
and UO_946 (O_946,N_19676,N_19975);
and UO_947 (O_947,N_19511,N_19924);
and UO_948 (O_948,N_19606,N_19885);
xor UO_949 (O_949,N_19592,N_19570);
and UO_950 (O_950,N_19759,N_19963);
nand UO_951 (O_951,N_19916,N_19879);
nor UO_952 (O_952,N_19649,N_19693);
or UO_953 (O_953,N_19938,N_19887);
and UO_954 (O_954,N_19633,N_19754);
xor UO_955 (O_955,N_19755,N_19822);
nor UO_956 (O_956,N_19906,N_19935);
nand UO_957 (O_957,N_19903,N_19634);
nor UO_958 (O_958,N_19512,N_19772);
nand UO_959 (O_959,N_19564,N_19714);
nand UO_960 (O_960,N_19510,N_19823);
and UO_961 (O_961,N_19916,N_19527);
or UO_962 (O_962,N_19683,N_19687);
or UO_963 (O_963,N_19609,N_19545);
nor UO_964 (O_964,N_19979,N_19727);
and UO_965 (O_965,N_19572,N_19646);
xor UO_966 (O_966,N_19599,N_19648);
nand UO_967 (O_967,N_19674,N_19819);
nor UO_968 (O_968,N_19728,N_19686);
nand UO_969 (O_969,N_19592,N_19668);
nor UO_970 (O_970,N_19778,N_19606);
or UO_971 (O_971,N_19819,N_19663);
xnor UO_972 (O_972,N_19896,N_19663);
or UO_973 (O_973,N_19767,N_19606);
xnor UO_974 (O_974,N_19968,N_19849);
nand UO_975 (O_975,N_19526,N_19780);
nand UO_976 (O_976,N_19783,N_19621);
nor UO_977 (O_977,N_19649,N_19647);
and UO_978 (O_978,N_19726,N_19910);
and UO_979 (O_979,N_19958,N_19869);
xor UO_980 (O_980,N_19964,N_19947);
nor UO_981 (O_981,N_19515,N_19658);
or UO_982 (O_982,N_19756,N_19670);
and UO_983 (O_983,N_19911,N_19591);
xnor UO_984 (O_984,N_19962,N_19647);
nand UO_985 (O_985,N_19934,N_19959);
nor UO_986 (O_986,N_19511,N_19968);
nand UO_987 (O_987,N_19906,N_19889);
nor UO_988 (O_988,N_19761,N_19957);
xor UO_989 (O_989,N_19754,N_19946);
and UO_990 (O_990,N_19670,N_19803);
and UO_991 (O_991,N_19999,N_19922);
nor UO_992 (O_992,N_19941,N_19693);
nand UO_993 (O_993,N_19753,N_19784);
or UO_994 (O_994,N_19538,N_19512);
nand UO_995 (O_995,N_19607,N_19844);
or UO_996 (O_996,N_19889,N_19752);
nor UO_997 (O_997,N_19881,N_19849);
or UO_998 (O_998,N_19749,N_19971);
xnor UO_999 (O_999,N_19612,N_19579);
nand UO_1000 (O_1000,N_19680,N_19777);
xnor UO_1001 (O_1001,N_19629,N_19878);
or UO_1002 (O_1002,N_19947,N_19968);
or UO_1003 (O_1003,N_19825,N_19979);
and UO_1004 (O_1004,N_19879,N_19701);
xor UO_1005 (O_1005,N_19656,N_19641);
nand UO_1006 (O_1006,N_19916,N_19815);
nor UO_1007 (O_1007,N_19733,N_19950);
xor UO_1008 (O_1008,N_19830,N_19841);
xnor UO_1009 (O_1009,N_19729,N_19819);
xnor UO_1010 (O_1010,N_19700,N_19928);
or UO_1011 (O_1011,N_19705,N_19641);
and UO_1012 (O_1012,N_19778,N_19777);
xor UO_1013 (O_1013,N_19502,N_19844);
or UO_1014 (O_1014,N_19729,N_19568);
nand UO_1015 (O_1015,N_19538,N_19839);
nand UO_1016 (O_1016,N_19605,N_19676);
xnor UO_1017 (O_1017,N_19597,N_19620);
nand UO_1018 (O_1018,N_19646,N_19614);
and UO_1019 (O_1019,N_19769,N_19624);
xnor UO_1020 (O_1020,N_19824,N_19690);
nand UO_1021 (O_1021,N_19523,N_19637);
nand UO_1022 (O_1022,N_19861,N_19837);
nand UO_1023 (O_1023,N_19868,N_19874);
and UO_1024 (O_1024,N_19522,N_19731);
and UO_1025 (O_1025,N_19671,N_19853);
xor UO_1026 (O_1026,N_19887,N_19899);
nand UO_1027 (O_1027,N_19500,N_19907);
or UO_1028 (O_1028,N_19818,N_19672);
nor UO_1029 (O_1029,N_19768,N_19602);
xnor UO_1030 (O_1030,N_19995,N_19962);
xor UO_1031 (O_1031,N_19690,N_19924);
nand UO_1032 (O_1032,N_19781,N_19922);
or UO_1033 (O_1033,N_19712,N_19794);
or UO_1034 (O_1034,N_19762,N_19777);
nor UO_1035 (O_1035,N_19703,N_19816);
nor UO_1036 (O_1036,N_19885,N_19654);
and UO_1037 (O_1037,N_19767,N_19783);
xor UO_1038 (O_1038,N_19647,N_19751);
xnor UO_1039 (O_1039,N_19835,N_19644);
nor UO_1040 (O_1040,N_19538,N_19885);
nand UO_1041 (O_1041,N_19590,N_19861);
xor UO_1042 (O_1042,N_19532,N_19831);
nand UO_1043 (O_1043,N_19831,N_19630);
or UO_1044 (O_1044,N_19775,N_19947);
nor UO_1045 (O_1045,N_19539,N_19502);
or UO_1046 (O_1046,N_19684,N_19936);
and UO_1047 (O_1047,N_19870,N_19710);
nand UO_1048 (O_1048,N_19508,N_19864);
nor UO_1049 (O_1049,N_19961,N_19628);
xnor UO_1050 (O_1050,N_19658,N_19831);
or UO_1051 (O_1051,N_19859,N_19664);
or UO_1052 (O_1052,N_19834,N_19593);
xor UO_1053 (O_1053,N_19530,N_19872);
xnor UO_1054 (O_1054,N_19762,N_19854);
or UO_1055 (O_1055,N_19676,N_19979);
xor UO_1056 (O_1056,N_19736,N_19628);
nand UO_1057 (O_1057,N_19641,N_19638);
nor UO_1058 (O_1058,N_19864,N_19545);
xor UO_1059 (O_1059,N_19982,N_19713);
nand UO_1060 (O_1060,N_19995,N_19617);
nor UO_1061 (O_1061,N_19867,N_19967);
and UO_1062 (O_1062,N_19831,N_19713);
or UO_1063 (O_1063,N_19603,N_19545);
nor UO_1064 (O_1064,N_19750,N_19864);
nand UO_1065 (O_1065,N_19780,N_19861);
nor UO_1066 (O_1066,N_19984,N_19756);
or UO_1067 (O_1067,N_19903,N_19722);
nor UO_1068 (O_1068,N_19632,N_19869);
nand UO_1069 (O_1069,N_19751,N_19878);
xnor UO_1070 (O_1070,N_19789,N_19929);
nand UO_1071 (O_1071,N_19745,N_19815);
and UO_1072 (O_1072,N_19603,N_19799);
xor UO_1073 (O_1073,N_19986,N_19689);
and UO_1074 (O_1074,N_19755,N_19789);
nor UO_1075 (O_1075,N_19812,N_19520);
and UO_1076 (O_1076,N_19734,N_19771);
xor UO_1077 (O_1077,N_19578,N_19726);
nand UO_1078 (O_1078,N_19618,N_19698);
and UO_1079 (O_1079,N_19966,N_19639);
nand UO_1080 (O_1080,N_19603,N_19544);
xnor UO_1081 (O_1081,N_19985,N_19834);
nand UO_1082 (O_1082,N_19801,N_19932);
nor UO_1083 (O_1083,N_19523,N_19557);
xnor UO_1084 (O_1084,N_19588,N_19514);
and UO_1085 (O_1085,N_19839,N_19888);
or UO_1086 (O_1086,N_19985,N_19994);
and UO_1087 (O_1087,N_19682,N_19623);
nand UO_1088 (O_1088,N_19912,N_19895);
and UO_1089 (O_1089,N_19745,N_19755);
nor UO_1090 (O_1090,N_19631,N_19823);
or UO_1091 (O_1091,N_19744,N_19979);
or UO_1092 (O_1092,N_19613,N_19546);
nand UO_1093 (O_1093,N_19644,N_19898);
or UO_1094 (O_1094,N_19868,N_19900);
and UO_1095 (O_1095,N_19524,N_19993);
or UO_1096 (O_1096,N_19527,N_19554);
or UO_1097 (O_1097,N_19553,N_19994);
nor UO_1098 (O_1098,N_19792,N_19725);
or UO_1099 (O_1099,N_19600,N_19874);
xnor UO_1100 (O_1100,N_19820,N_19505);
and UO_1101 (O_1101,N_19553,N_19724);
or UO_1102 (O_1102,N_19737,N_19585);
or UO_1103 (O_1103,N_19846,N_19997);
or UO_1104 (O_1104,N_19938,N_19773);
nor UO_1105 (O_1105,N_19500,N_19522);
or UO_1106 (O_1106,N_19688,N_19782);
and UO_1107 (O_1107,N_19861,N_19703);
and UO_1108 (O_1108,N_19718,N_19843);
and UO_1109 (O_1109,N_19811,N_19788);
or UO_1110 (O_1110,N_19765,N_19914);
nand UO_1111 (O_1111,N_19870,N_19537);
and UO_1112 (O_1112,N_19609,N_19987);
nor UO_1113 (O_1113,N_19973,N_19581);
xnor UO_1114 (O_1114,N_19567,N_19886);
nand UO_1115 (O_1115,N_19609,N_19666);
nand UO_1116 (O_1116,N_19784,N_19996);
and UO_1117 (O_1117,N_19803,N_19581);
and UO_1118 (O_1118,N_19660,N_19974);
nor UO_1119 (O_1119,N_19779,N_19775);
and UO_1120 (O_1120,N_19526,N_19975);
nand UO_1121 (O_1121,N_19771,N_19660);
nand UO_1122 (O_1122,N_19897,N_19615);
nor UO_1123 (O_1123,N_19875,N_19561);
nor UO_1124 (O_1124,N_19688,N_19781);
nand UO_1125 (O_1125,N_19986,N_19555);
and UO_1126 (O_1126,N_19895,N_19704);
xor UO_1127 (O_1127,N_19785,N_19514);
nand UO_1128 (O_1128,N_19703,N_19842);
nor UO_1129 (O_1129,N_19954,N_19937);
nand UO_1130 (O_1130,N_19788,N_19782);
or UO_1131 (O_1131,N_19788,N_19761);
nor UO_1132 (O_1132,N_19801,N_19806);
or UO_1133 (O_1133,N_19794,N_19683);
nor UO_1134 (O_1134,N_19882,N_19993);
xor UO_1135 (O_1135,N_19631,N_19804);
or UO_1136 (O_1136,N_19719,N_19750);
and UO_1137 (O_1137,N_19728,N_19625);
and UO_1138 (O_1138,N_19728,N_19768);
or UO_1139 (O_1139,N_19964,N_19799);
xnor UO_1140 (O_1140,N_19620,N_19814);
nand UO_1141 (O_1141,N_19762,N_19903);
nand UO_1142 (O_1142,N_19533,N_19706);
nand UO_1143 (O_1143,N_19568,N_19860);
nor UO_1144 (O_1144,N_19911,N_19980);
nand UO_1145 (O_1145,N_19545,N_19628);
xnor UO_1146 (O_1146,N_19845,N_19571);
or UO_1147 (O_1147,N_19615,N_19885);
and UO_1148 (O_1148,N_19750,N_19729);
nand UO_1149 (O_1149,N_19964,N_19916);
xor UO_1150 (O_1150,N_19763,N_19663);
xnor UO_1151 (O_1151,N_19979,N_19828);
nand UO_1152 (O_1152,N_19993,N_19736);
or UO_1153 (O_1153,N_19845,N_19891);
or UO_1154 (O_1154,N_19962,N_19537);
and UO_1155 (O_1155,N_19803,N_19574);
nand UO_1156 (O_1156,N_19910,N_19897);
and UO_1157 (O_1157,N_19683,N_19724);
xor UO_1158 (O_1158,N_19730,N_19916);
or UO_1159 (O_1159,N_19726,N_19575);
or UO_1160 (O_1160,N_19553,N_19665);
nor UO_1161 (O_1161,N_19867,N_19565);
nor UO_1162 (O_1162,N_19809,N_19790);
and UO_1163 (O_1163,N_19632,N_19668);
and UO_1164 (O_1164,N_19702,N_19626);
xnor UO_1165 (O_1165,N_19799,N_19534);
nor UO_1166 (O_1166,N_19843,N_19886);
or UO_1167 (O_1167,N_19973,N_19529);
or UO_1168 (O_1168,N_19896,N_19884);
xor UO_1169 (O_1169,N_19542,N_19753);
or UO_1170 (O_1170,N_19674,N_19934);
or UO_1171 (O_1171,N_19568,N_19522);
nor UO_1172 (O_1172,N_19564,N_19822);
xor UO_1173 (O_1173,N_19663,N_19958);
xor UO_1174 (O_1174,N_19634,N_19656);
or UO_1175 (O_1175,N_19617,N_19794);
or UO_1176 (O_1176,N_19932,N_19723);
or UO_1177 (O_1177,N_19843,N_19865);
xnor UO_1178 (O_1178,N_19683,N_19722);
xor UO_1179 (O_1179,N_19997,N_19967);
or UO_1180 (O_1180,N_19784,N_19776);
and UO_1181 (O_1181,N_19903,N_19751);
or UO_1182 (O_1182,N_19888,N_19504);
xnor UO_1183 (O_1183,N_19510,N_19547);
or UO_1184 (O_1184,N_19603,N_19897);
and UO_1185 (O_1185,N_19511,N_19560);
or UO_1186 (O_1186,N_19824,N_19928);
nand UO_1187 (O_1187,N_19661,N_19747);
nor UO_1188 (O_1188,N_19920,N_19547);
nor UO_1189 (O_1189,N_19857,N_19877);
nand UO_1190 (O_1190,N_19785,N_19929);
nand UO_1191 (O_1191,N_19695,N_19989);
nand UO_1192 (O_1192,N_19908,N_19619);
nand UO_1193 (O_1193,N_19789,N_19530);
or UO_1194 (O_1194,N_19790,N_19757);
nand UO_1195 (O_1195,N_19890,N_19625);
xor UO_1196 (O_1196,N_19876,N_19670);
and UO_1197 (O_1197,N_19504,N_19573);
nand UO_1198 (O_1198,N_19911,N_19769);
xor UO_1199 (O_1199,N_19685,N_19787);
and UO_1200 (O_1200,N_19580,N_19865);
xnor UO_1201 (O_1201,N_19956,N_19555);
or UO_1202 (O_1202,N_19816,N_19942);
nor UO_1203 (O_1203,N_19563,N_19944);
or UO_1204 (O_1204,N_19749,N_19951);
nor UO_1205 (O_1205,N_19923,N_19692);
and UO_1206 (O_1206,N_19615,N_19560);
and UO_1207 (O_1207,N_19541,N_19929);
nand UO_1208 (O_1208,N_19651,N_19617);
nor UO_1209 (O_1209,N_19939,N_19733);
nor UO_1210 (O_1210,N_19989,N_19864);
nor UO_1211 (O_1211,N_19719,N_19748);
xnor UO_1212 (O_1212,N_19755,N_19545);
and UO_1213 (O_1213,N_19860,N_19786);
and UO_1214 (O_1214,N_19702,N_19946);
or UO_1215 (O_1215,N_19855,N_19830);
nand UO_1216 (O_1216,N_19873,N_19581);
xor UO_1217 (O_1217,N_19535,N_19691);
or UO_1218 (O_1218,N_19634,N_19920);
and UO_1219 (O_1219,N_19669,N_19994);
nand UO_1220 (O_1220,N_19974,N_19790);
xor UO_1221 (O_1221,N_19843,N_19617);
nor UO_1222 (O_1222,N_19714,N_19658);
nand UO_1223 (O_1223,N_19981,N_19667);
xnor UO_1224 (O_1224,N_19517,N_19558);
nand UO_1225 (O_1225,N_19526,N_19976);
xnor UO_1226 (O_1226,N_19942,N_19978);
or UO_1227 (O_1227,N_19870,N_19598);
xor UO_1228 (O_1228,N_19589,N_19940);
xnor UO_1229 (O_1229,N_19993,N_19883);
and UO_1230 (O_1230,N_19611,N_19877);
xor UO_1231 (O_1231,N_19591,N_19638);
nand UO_1232 (O_1232,N_19945,N_19684);
and UO_1233 (O_1233,N_19915,N_19922);
xnor UO_1234 (O_1234,N_19626,N_19875);
or UO_1235 (O_1235,N_19952,N_19861);
nand UO_1236 (O_1236,N_19846,N_19686);
and UO_1237 (O_1237,N_19815,N_19905);
xor UO_1238 (O_1238,N_19653,N_19587);
nor UO_1239 (O_1239,N_19617,N_19874);
and UO_1240 (O_1240,N_19966,N_19653);
or UO_1241 (O_1241,N_19546,N_19693);
nand UO_1242 (O_1242,N_19663,N_19628);
and UO_1243 (O_1243,N_19664,N_19529);
nor UO_1244 (O_1244,N_19831,N_19827);
xnor UO_1245 (O_1245,N_19531,N_19743);
and UO_1246 (O_1246,N_19976,N_19884);
or UO_1247 (O_1247,N_19590,N_19609);
nor UO_1248 (O_1248,N_19582,N_19664);
and UO_1249 (O_1249,N_19985,N_19881);
nor UO_1250 (O_1250,N_19668,N_19518);
xor UO_1251 (O_1251,N_19889,N_19580);
and UO_1252 (O_1252,N_19617,N_19668);
nor UO_1253 (O_1253,N_19760,N_19749);
xnor UO_1254 (O_1254,N_19946,N_19814);
and UO_1255 (O_1255,N_19580,N_19970);
nand UO_1256 (O_1256,N_19659,N_19943);
nand UO_1257 (O_1257,N_19812,N_19586);
and UO_1258 (O_1258,N_19533,N_19775);
and UO_1259 (O_1259,N_19792,N_19955);
nor UO_1260 (O_1260,N_19649,N_19972);
nand UO_1261 (O_1261,N_19517,N_19564);
nand UO_1262 (O_1262,N_19919,N_19736);
and UO_1263 (O_1263,N_19757,N_19657);
xnor UO_1264 (O_1264,N_19743,N_19665);
nand UO_1265 (O_1265,N_19932,N_19981);
or UO_1266 (O_1266,N_19958,N_19852);
or UO_1267 (O_1267,N_19787,N_19961);
nand UO_1268 (O_1268,N_19640,N_19711);
nand UO_1269 (O_1269,N_19943,N_19879);
nand UO_1270 (O_1270,N_19964,N_19688);
nor UO_1271 (O_1271,N_19835,N_19589);
nand UO_1272 (O_1272,N_19761,N_19751);
or UO_1273 (O_1273,N_19896,N_19902);
nand UO_1274 (O_1274,N_19982,N_19731);
xor UO_1275 (O_1275,N_19895,N_19573);
and UO_1276 (O_1276,N_19955,N_19878);
or UO_1277 (O_1277,N_19660,N_19542);
and UO_1278 (O_1278,N_19915,N_19776);
and UO_1279 (O_1279,N_19754,N_19715);
and UO_1280 (O_1280,N_19947,N_19981);
xor UO_1281 (O_1281,N_19911,N_19754);
nor UO_1282 (O_1282,N_19776,N_19581);
or UO_1283 (O_1283,N_19873,N_19592);
nor UO_1284 (O_1284,N_19916,N_19712);
nor UO_1285 (O_1285,N_19767,N_19736);
nor UO_1286 (O_1286,N_19734,N_19652);
and UO_1287 (O_1287,N_19670,N_19788);
and UO_1288 (O_1288,N_19826,N_19586);
or UO_1289 (O_1289,N_19620,N_19794);
and UO_1290 (O_1290,N_19940,N_19644);
nand UO_1291 (O_1291,N_19698,N_19751);
nor UO_1292 (O_1292,N_19740,N_19817);
or UO_1293 (O_1293,N_19789,N_19696);
nand UO_1294 (O_1294,N_19556,N_19737);
or UO_1295 (O_1295,N_19728,N_19991);
nor UO_1296 (O_1296,N_19651,N_19501);
xnor UO_1297 (O_1297,N_19787,N_19593);
or UO_1298 (O_1298,N_19999,N_19790);
and UO_1299 (O_1299,N_19871,N_19939);
and UO_1300 (O_1300,N_19803,N_19720);
nand UO_1301 (O_1301,N_19993,N_19791);
nand UO_1302 (O_1302,N_19980,N_19698);
xnor UO_1303 (O_1303,N_19539,N_19605);
nand UO_1304 (O_1304,N_19977,N_19602);
nand UO_1305 (O_1305,N_19788,N_19892);
and UO_1306 (O_1306,N_19709,N_19630);
nor UO_1307 (O_1307,N_19713,N_19751);
and UO_1308 (O_1308,N_19991,N_19821);
and UO_1309 (O_1309,N_19520,N_19853);
nor UO_1310 (O_1310,N_19705,N_19554);
and UO_1311 (O_1311,N_19703,N_19897);
nor UO_1312 (O_1312,N_19538,N_19602);
and UO_1313 (O_1313,N_19981,N_19831);
and UO_1314 (O_1314,N_19573,N_19918);
nand UO_1315 (O_1315,N_19776,N_19545);
nand UO_1316 (O_1316,N_19562,N_19525);
and UO_1317 (O_1317,N_19748,N_19591);
nor UO_1318 (O_1318,N_19510,N_19559);
nor UO_1319 (O_1319,N_19873,N_19633);
and UO_1320 (O_1320,N_19897,N_19633);
xor UO_1321 (O_1321,N_19892,N_19505);
nand UO_1322 (O_1322,N_19572,N_19684);
or UO_1323 (O_1323,N_19621,N_19938);
nor UO_1324 (O_1324,N_19694,N_19749);
or UO_1325 (O_1325,N_19797,N_19668);
or UO_1326 (O_1326,N_19640,N_19906);
xnor UO_1327 (O_1327,N_19719,N_19804);
or UO_1328 (O_1328,N_19520,N_19929);
or UO_1329 (O_1329,N_19649,N_19942);
or UO_1330 (O_1330,N_19678,N_19730);
or UO_1331 (O_1331,N_19924,N_19947);
or UO_1332 (O_1332,N_19596,N_19550);
nand UO_1333 (O_1333,N_19833,N_19860);
and UO_1334 (O_1334,N_19701,N_19730);
and UO_1335 (O_1335,N_19802,N_19959);
or UO_1336 (O_1336,N_19614,N_19695);
and UO_1337 (O_1337,N_19950,N_19633);
nand UO_1338 (O_1338,N_19779,N_19503);
nand UO_1339 (O_1339,N_19994,N_19780);
or UO_1340 (O_1340,N_19786,N_19821);
nor UO_1341 (O_1341,N_19942,N_19850);
nand UO_1342 (O_1342,N_19585,N_19891);
nor UO_1343 (O_1343,N_19688,N_19756);
xor UO_1344 (O_1344,N_19942,N_19726);
nand UO_1345 (O_1345,N_19508,N_19823);
xor UO_1346 (O_1346,N_19969,N_19734);
nor UO_1347 (O_1347,N_19569,N_19929);
nand UO_1348 (O_1348,N_19869,N_19650);
nor UO_1349 (O_1349,N_19555,N_19761);
and UO_1350 (O_1350,N_19524,N_19504);
or UO_1351 (O_1351,N_19573,N_19517);
nand UO_1352 (O_1352,N_19660,N_19891);
or UO_1353 (O_1353,N_19865,N_19784);
nor UO_1354 (O_1354,N_19859,N_19633);
nand UO_1355 (O_1355,N_19702,N_19646);
nand UO_1356 (O_1356,N_19696,N_19589);
xor UO_1357 (O_1357,N_19671,N_19796);
or UO_1358 (O_1358,N_19766,N_19754);
nand UO_1359 (O_1359,N_19828,N_19623);
and UO_1360 (O_1360,N_19570,N_19966);
xor UO_1361 (O_1361,N_19612,N_19851);
nand UO_1362 (O_1362,N_19794,N_19614);
or UO_1363 (O_1363,N_19930,N_19582);
xor UO_1364 (O_1364,N_19506,N_19562);
or UO_1365 (O_1365,N_19955,N_19663);
nand UO_1366 (O_1366,N_19705,N_19863);
and UO_1367 (O_1367,N_19828,N_19843);
and UO_1368 (O_1368,N_19531,N_19553);
or UO_1369 (O_1369,N_19747,N_19534);
and UO_1370 (O_1370,N_19898,N_19839);
xnor UO_1371 (O_1371,N_19692,N_19951);
or UO_1372 (O_1372,N_19786,N_19982);
or UO_1373 (O_1373,N_19974,N_19828);
nor UO_1374 (O_1374,N_19973,N_19503);
or UO_1375 (O_1375,N_19840,N_19626);
xnor UO_1376 (O_1376,N_19683,N_19941);
or UO_1377 (O_1377,N_19967,N_19858);
xnor UO_1378 (O_1378,N_19706,N_19734);
or UO_1379 (O_1379,N_19601,N_19805);
and UO_1380 (O_1380,N_19736,N_19829);
nand UO_1381 (O_1381,N_19684,N_19807);
or UO_1382 (O_1382,N_19960,N_19976);
and UO_1383 (O_1383,N_19884,N_19603);
or UO_1384 (O_1384,N_19705,N_19525);
nor UO_1385 (O_1385,N_19983,N_19796);
nor UO_1386 (O_1386,N_19552,N_19562);
nand UO_1387 (O_1387,N_19645,N_19643);
nand UO_1388 (O_1388,N_19876,N_19919);
and UO_1389 (O_1389,N_19820,N_19822);
or UO_1390 (O_1390,N_19712,N_19974);
nand UO_1391 (O_1391,N_19501,N_19624);
nand UO_1392 (O_1392,N_19825,N_19588);
and UO_1393 (O_1393,N_19906,N_19551);
nor UO_1394 (O_1394,N_19573,N_19674);
or UO_1395 (O_1395,N_19876,N_19711);
or UO_1396 (O_1396,N_19789,N_19676);
xnor UO_1397 (O_1397,N_19849,N_19940);
xor UO_1398 (O_1398,N_19817,N_19651);
nor UO_1399 (O_1399,N_19515,N_19542);
and UO_1400 (O_1400,N_19964,N_19773);
nor UO_1401 (O_1401,N_19866,N_19556);
or UO_1402 (O_1402,N_19953,N_19943);
nor UO_1403 (O_1403,N_19884,N_19905);
or UO_1404 (O_1404,N_19604,N_19514);
xor UO_1405 (O_1405,N_19792,N_19539);
or UO_1406 (O_1406,N_19771,N_19687);
and UO_1407 (O_1407,N_19628,N_19872);
and UO_1408 (O_1408,N_19582,N_19591);
nand UO_1409 (O_1409,N_19539,N_19618);
or UO_1410 (O_1410,N_19819,N_19913);
and UO_1411 (O_1411,N_19756,N_19648);
nand UO_1412 (O_1412,N_19724,N_19670);
nand UO_1413 (O_1413,N_19804,N_19833);
xor UO_1414 (O_1414,N_19773,N_19769);
or UO_1415 (O_1415,N_19938,N_19544);
xnor UO_1416 (O_1416,N_19644,N_19844);
and UO_1417 (O_1417,N_19519,N_19503);
nor UO_1418 (O_1418,N_19811,N_19777);
or UO_1419 (O_1419,N_19510,N_19511);
xnor UO_1420 (O_1420,N_19549,N_19868);
or UO_1421 (O_1421,N_19661,N_19881);
or UO_1422 (O_1422,N_19983,N_19899);
nor UO_1423 (O_1423,N_19912,N_19902);
or UO_1424 (O_1424,N_19764,N_19983);
and UO_1425 (O_1425,N_19873,N_19714);
nor UO_1426 (O_1426,N_19590,N_19720);
nor UO_1427 (O_1427,N_19869,N_19963);
and UO_1428 (O_1428,N_19961,N_19524);
and UO_1429 (O_1429,N_19807,N_19897);
xor UO_1430 (O_1430,N_19681,N_19815);
nor UO_1431 (O_1431,N_19744,N_19895);
xnor UO_1432 (O_1432,N_19956,N_19637);
nor UO_1433 (O_1433,N_19715,N_19757);
nor UO_1434 (O_1434,N_19777,N_19996);
nor UO_1435 (O_1435,N_19649,N_19965);
nand UO_1436 (O_1436,N_19740,N_19506);
nor UO_1437 (O_1437,N_19660,N_19680);
or UO_1438 (O_1438,N_19650,N_19929);
nor UO_1439 (O_1439,N_19691,N_19827);
or UO_1440 (O_1440,N_19842,N_19506);
xnor UO_1441 (O_1441,N_19912,N_19582);
and UO_1442 (O_1442,N_19853,N_19939);
xor UO_1443 (O_1443,N_19786,N_19641);
or UO_1444 (O_1444,N_19722,N_19503);
nand UO_1445 (O_1445,N_19972,N_19528);
or UO_1446 (O_1446,N_19731,N_19609);
and UO_1447 (O_1447,N_19698,N_19670);
nor UO_1448 (O_1448,N_19699,N_19656);
or UO_1449 (O_1449,N_19884,N_19511);
and UO_1450 (O_1450,N_19566,N_19743);
and UO_1451 (O_1451,N_19787,N_19764);
nor UO_1452 (O_1452,N_19578,N_19827);
nand UO_1453 (O_1453,N_19988,N_19640);
and UO_1454 (O_1454,N_19613,N_19883);
nor UO_1455 (O_1455,N_19520,N_19658);
or UO_1456 (O_1456,N_19985,N_19528);
nor UO_1457 (O_1457,N_19605,N_19727);
nor UO_1458 (O_1458,N_19603,N_19540);
nand UO_1459 (O_1459,N_19873,N_19941);
and UO_1460 (O_1460,N_19968,N_19619);
xor UO_1461 (O_1461,N_19819,N_19574);
or UO_1462 (O_1462,N_19723,N_19687);
xor UO_1463 (O_1463,N_19505,N_19612);
nor UO_1464 (O_1464,N_19873,N_19806);
nor UO_1465 (O_1465,N_19583,N_19568);
or UO_1466 (O_1466,N_19884,N_19695);
or UO_1467 (O_1467,N_19753,N_19657);
and UO_1468 (O_1468,N_19724,N_19694);
or UO_1469 (O_1469,N_19570,N_19627);
and UO_1470 (O_1470,N_19929,N_19586);
nor UO_1471 (O_1471,N_19860,N_19671);
nor UO_1472 (O_1472,N_19509,N_19519);
and UO_1473 (O_1473,N_19640,N_19861);
and UO_1474 (O_1474,N_19591,N_19940);
nor UO_1475 (O_1475,N_19740,N_19805);
xor UO_1476 (O_1476,N_19666,N_19528);
or UO_1477 (O_1477,N_19629,N_19632);
nor UO_1478 (O_1478,N_19709,N_19502);
and UO_1479 (O_1479,N_19780,N_19986);
nand UO_1480 (O_1480,N_19933,N_19718);
nand UO_1481 (O_1481,N_19876,N_19683);
nor UO_1482 (O_1482,N_19868,N_19889);
and UO_1483 (O_1483,N_19968,N_19886);
nor UO_1484 (O_1484,N_19945,N_19672);
nor UO_1485 (O_1485,N_19971,N_19974);
nor UO_1486 (O_1486,N_19804,N_19914);
xor UO_1487 (O_1487,N_19527,N_19533);
or UO_1488 (O_1488,N_19705,N_19644);
nand UO_1489 (O_1489,N_19603,N_19922);
xnor UO_1490 (O_1490,N_19956,N_19581);
xor UO_1491 (O_1491,N_19793,N_19844);
or UO_1492 (O_1492,N_19865,N_19721);
or UO_1493 (O_1493,N_19840,N_19792);
and UO_1494 (O_1494,N_19661,N_19562);
nand UO_1495 (O_1495,N_19842,N_19865);
and UO_1496 (O_1496,N_19644,N_19780);
xnor UO_1497 (O_1497,N_19993,N_19701);
nand UO_1498 (O_1498,N_19548,N_19825);
nand UO_1499 (O_1499,N_19754,N_19909);
xor UO_1500 (O_1500,N_19557,N_19744);
and UO_1501 (O_1501,N_19718,N_19639);
and UO_1502 (O_1502,N_19852,N_19822);
and UO_1503 (O_1503,N_19611,N_19592);
nor UO_1504 (O_1504,N_19542,N_19561);
or UO_1505 (O_1505,N_19778,N_19794);
or UO_1506 (O_1506,N_19517,N_19935);
and UO_1507 (O_1507,N_19984,N_19846);
nor UO_1508 (O_1508,N_19795,N_19655);
nor UO_1509 (O_1509,N_19812,N_19831);
and UO_1510 (O_1510,N_19989,N_19907);
nand UO_1511 (O_1511,N_19561,N_19652);
or UO_1512 (O_1512,N_19989,N_19952);
or UO_1513 (O_1513,N_19545,N_19824);
nor UO_1514 (O_1514,N_19803,N_19722);
nor UO_1515 (O_1515,N_19606,N_19725);
or UO_1516 (O_1516,N_19679,N_19949);
xnor UO_1517 (O_1517,N_19747,N_19682);
xnor UO_1518 (O_1518,N_19531,N_19913);
or UO_1519 (O_1519,N_19982,N_19977);
nor UO_1520 (O_1520,N_19838,N_19892);
nand UO_1521 (O_1521,N_19879,N_19986);
or UO_1522 (O_1522,N_19723,N_19653);
and UO_1523 (O_1523,N_19631,N_19691);
nor UO_1524 (O_1524,N_19593,N_19932);
nor UO_1525 (O_1525,N_19572,N_19674);
xor UO_1526 (O_1526,N_19911,N_19895);
and UO_1527 (O_1527,N_19760,N_19647);
or UO_1528 (O_1528,N_19825,N_19838);
and UO_1529 (O_1529,N_19951,N_19754);
nor UO_1530 (O_1530,N_19928,N_19614);
nand UO_1531 (O_1531,N_19537,N_19775);
and UO_1532 (O_1532,N_19801,N_19864);
nand UO_1533 (O_1533,N_19974,N_19739);
nand UO_1534 (O_1534,N_19526,N_19964);
and UO_1535 (O_1535,N_19958,N_19631);
nand UO_1536 (O_1536,N_19658,N_19526);
and UO_1537 (O_1537,N_19607,N_19745);
or UO_1538 (O_1538,N_19911,N_19837);
or UO_1539 (O_1539,N_19870,N_19844);
nor UO_1540 (O_1540,N_19789,N_19527);
nor UO_1541 (O_1541,N_19756,N_19874);
xnor UO_1542 (O_1542,N_19930,N_19597);
or UO_1543 (O_1543,N_19929,N_19672);
xor UO_1544 (O_1544,N_19591,N_19856);
and UO_1545 (O_1545,N_19651,N_19872);
and UO_1546 (O_1546,N_19889,N_19650);
nor UO_1547 (O_1547,N_19643,N_19705);
xnor UO_1548 (O_1548,N_19526,N_19792);
or UO_1549 (O_1549,N_19605,N_19996);
nand UO_1550 (O_1550,N_19635,N_19950);
nor UO_1551 (O_1551,N_19799,N_19974);
and UO_1552 (O_1552,N_19949,N_19957);
xor UO_1553 (O_1553,N_19606,N_19776);
nand UO_1554 (O_1554,N_19576,N_19831);
xor UO_1555 (O_1555,N_19664,N_19889);
or UO_1556 (O_1556,N_19551,N_19713);
and UO_1557 (O_1557,N_19694,N_19740);
and UO_1558 (O_1558,N_19596,N_19635);
nand UO_1559 (O_1559,N_19880,N_19855);
or UO_1560 (O_1560,N_19776,N_19555);
nand UO_1561 (O_1561,N_19575,N_19886);
xor UO_1562 (O_1562,N_19883,N_19833);
nand UO_1563 (O_1563,N_19801,N_19551);
and UO_1564 (O_1564,N_19611,N_19554);
and UO_1565 (O_1565,N_19631,N_19564);
nor UO_1566 (O_1566,N_19642,N_19688);
and UO_1567 (O_1567,N_19687,N_19873);
or UO_1568 (O_1568,N_19873,N_19747);
or UO_1569 (O_1569,N_19987,N_19538);
and UO_1570 (O_1570,N_19543,N_19770);
nor UO_1571 (O_1571,N_19766,N_19827);
or UO_1572 (O_1572,N_19518,N_19868);
nor UO_1573 (O_1573,N_19551,N_19759);
xnor UO_1574 (O_1574,N_19522,N_19949);
nand UO_1575 (O_1575,N_19518,N_19680);
nand UO_1576 (O_1576,N_19614,N_19722);
xor UO_1577 (O_1577,N_19801,N_19866);
xnor UO_1578 (O_1578,N_19582,N_19872);
xor UO_1579 (O_1579,N_19834,N_19553);
or UO_1580 (O_1580,N_19688,N_19766);
nand UO_1581 (O_1581,N_19690,N_19542);
or UO_1582 (O_1582,N_19938,N_19705);
and UO_1583 (O_1583,N_19774,N_19606);
or UO_1584 (O_1584,N_19901,N_19797);
or UO_1585 (O_1585,N_19630,N_19920);
xor UO_1586 (O_1586,N_19906,N_19949);
nor UO_1587 (O_1587,N_19687,N_19519);
nand UO_1588 (O_1588,N_19539,N_19558);
or UO_1589 (O_1589,N_19784,N_19659);
nor UO_1590 (O_1590,N_19690,N_19717);
or UO_1591 (O_1591,N_19888,N_19726);
or UO_1592 (O_1592,N_19945,N_19631);
nor UO_1593 (O_1593,N_19685,N_19544);
or UO_1594 (O_1594,N_19550,N_19879);
nor UO_1595 (O_1595,N_19791,N_19984);
nor UO_1596 (O_1596,N_19527,N_19878);
xor UO_1597 (O_1597,N_19542,N_19935);
and UO_1598 (O_1598,N_19735,N_19826);
xnor UO_1599 (O_1599,N_19889,N_19945);
nand UO_1600 (O_1600,N_19964,N_19524);
xor UO_1601 (O_1601,N_19750,N_19817);
nor UO_1602 (O_1602,N_19975,N_19548);
xnor UO_1603 (O_1603,N_19728,N_19665);
or UO_1604 (O_1604,N_19563,N_19832);
nor UO_1605 (O_1605,N_19731,N_19938);
or UO_1606 (O_1606,N_19862,N_19872);
xnor UO_1607 (O_1607,N_19616,N_19970);
xnor UO_1608 (O_1608,N_19809,N_19593);
and UO_1609 (O_1609,N_19535,N_19533);
or UO_1610 (O_1610,N_19630,N_19561);
nor UO_1611 (O_1611,N_19708,N_19641);
nand UO_1612 (O_1612,N_19738,N_19903);
nand UO_1613 (O_1613,N_19824,N_19744);
or UO_1614 (O_1614,N_19808,N_19690);
nor UO_1615 (O_1615,N_19618,N_19756);
nand UO_1616 (O_1616,N_19861,N_19742);
nand UO_1617 (O_1617,N_19694,N_19922);
or UO_1618 (O_1618,N_19948,N_19965);
nor UO_1619 (O_1619,N_19539,N_19675);
xor UO_1620 (O_1620,N_19570,N_19846);
and UO_1621 (O_1621,N_19555,N_19898);
xor UO_1622 (O_1622,N_19967,N_19894);
or UO_1623 (O_1623,N_19945,N_19701);
and UO_1624 (O_1624,N_19886,N_19959);
nor UO_1625 (O_1625,N_19856,N_19764);
nand UO_1626 (O_1626,N_19812,N_19937);
and UO_1627 (O_1627,N_19862,N_19905);
xor UO_1628 (O_1628,N_19797,N_19592);
and UO_1629 (O_1629,N_19528,N_19742);
xor UO_1630 (O_1630,N_19708,N_19775);
or UO_1631 (O_1631,N_19643,N_19953);
nand UO_1632 (O_1632,N_19795,N_19539);
and UO_1633 (O_1633,N_19659,N_19867);
or UO_1634 (O_1634,N_19525,N_19536);
nor UO_1635 (O_1635,N_19570,N_19801);
xor UO_1636 (O_1636,N_19717,N_19896);
nor UO_1637 (O_1637,N_19961,N_19976);
nand UO_1638 (O_1638,N_19895,N_19555);
nor UO_1639 (O_1639,N_19772,N_19975);
and UO_1640 (O_1640,N_19701,N_19699);
xnor UO_1641 (O_1641,N_19522,N_19549);
xnor UO_1642 (O_1642,N_19556,N_19779);
and UO_1643 (O_1643,N_19982,N_19811);
nor UO_1644 (O_1644,N_19636,N_19801);
nor UO_1645 (O_1645,N_19592,N_19880);
or UO_1646 (O_1646,N_19885,N_19747);
xnor UO_1647 (O_1647,N_19661,N_19706);
nor UO_1648 (O_1648,N_19785,N_19521);
xnor UO_1649 (O_1649,N_19505,N_19638);
nand UO_1650 (O_1650,N_19823,N_19587);
xnor UO_1651 (O_1651,N_19613,N_19662);
or UO_1652 (O_1652,N_19907,N_19639);
nand UO_1653 (O_1653,N_19786,N_19580);
or UO_1654 (O_1654,N_19923,N_19767);
nor UO_1655 (O_1655,N_19516,N_19735);
nor UO_1656 (O_1656,N_19763,N_19875);
nand UO_1657 (O_1657,N_19974,N_19765);
xor UO_1658 (O_1658,N_19824,N_19898);
xnor UO_1659 (O_1659,N_19772,N_19853);
nand UO_1660 (O_1660,N_19853,N_19735);
and UO_1661 (O_1661,N_19526,N_19746);
xnor UO_1662 (O_1662,N_19583,N_19710);
xnor UO_1663 (O_1663,N_19538,N_19723);
and UO_1664 (O_1664,N_19556,N_19650);
nor UO_1665 (O_1665,N_19875,N_19966);
nand UO_1666 (O_1666,N_19966,N_19530);
nand UO_1667 (O_1667,N_19518,N_19538);
nor UO_1668 (O_1668,N_19859,N_19866);
nor UO_1669 (O_1669,N_19868,N_19500);
or UO_1670 (O_1670,N_19874,N_19676);
xor UO_1671 (O_1671,N_19956,N_19559);
and UO_1672 (O_1672,N_19941,N_19619);
and UO_1673 (O_1673,N_19565,N_19513);
nor UO_1674 (O_1674,N_19882,N_19700);
nor UO_1675 (O_1675,N_19794,N_19565);
nor UO_1676 (O_1676,N_19873,N_19628);
xor UO_1677 (O_1677,N_19729,N_19639);
and UO_1678 (O_1678,N_19654,N_19806);
xor UO_1679 (O_1679,N_19593,N_19746);
nor UO_1680 (O_1680,N_19887,N_19597);
and UO_1681 (O_1681,N_19684,N_19535);
and UO_1682 (O_1682,N_19682,N_19804);
nand UO_1683 (O_1683,N_19547,N_19781);
or UO_1684 (O_1684,N_19550,N_19834);
or UO_1685 (O_1685,N_19725,N_19607);
or UO_1686 (O_1686,N_19680,N_19694);
and UO_1687 (O_1687,N_19609,N_19658);
xnor UO_1688 (O_1688,N_19766,N_19864);
and UO_1689 (O_1689,N_19681,N_19618);
xnor UO_1690 (O_1690,N_19983,N_19544);
nand UO_1691 (O_1691,N_19917,N_19589);
nor UO_1692 (O_1692,N_19924,N_19644);
or UO_1693 (O_1693,N_19806,N_19908);
or UO_1694 (O_1694,N_19705,N_19893);
or UO_1695 (O_1695,N_19645,N_19965);
nand UO_1696 (O_1696,N_19786,N_19714);
nor UO_1697 (O_1697,N_19652,N_19644);
and UO_1698 (O_1698,N_19786,N_19885);
and UO_1699 (O_1699,N_19750,N_19876);
or UO_1700 (O_1700,N_19894,N_19710);
nand UO_1701 (O_1701,N_19736,N_19984);
and UO_1702 (O_1702,N_19842,N_19807);
nand UO_1703 (O_1703,N_19534,N_19925);
nand UO_1704 (O_1704,N_19561,N_19841);
nand UO_1705 (O_1705,N_19793,N_19970);
xnor UO_1706 (O_1706,N_19862,N_19647);
nor UO_1707 (O_1707,N_19909,N_19993);
xnor UO_1708 (O_1708,N_19564,N_19737);
and UO_1709 (O_1709,N_19819,N_19680);
or UO_1710 (O_1710,N_19788,N_19978);
nand UO_1711 (O_1711,N_19988,N_19802);
nor UO_1712 (O_1712,N_19867,N_19586);
or UO_1713 (O_1713,N_19679,N_19527);
nor UO_1714 (O_1714,N_19968,N_19536);
and UO_1715 (O_1715,N_19604,N_19761);
or UO_1716 (O_1716,N_19866,N_19938);
nor UO_1717 (O_1717,N_19989,N_19967);
nand UO_1718 (O_1718,N_19839,N_19908);
nand UO_1719 (O_1719,N_19753,N_19807);
nand UO_1720 (O_1720,N_19989,N_19802);
or UO_1721 (O_1721,N_19653,N_19599);
nor UO_1722 (O_1722,N_19501,N_19903);
or UO_1723 (O_1723,N_19855,N_19598);
xor UO_1724 (O_1724,N_19766,N_19939);
or UO_1725 (O_1725,N_19705,N_19868);
nand UO_1726 (O_1726,N_19819,N_19730);
xor UO_1727 (O_1727,N_19768,N_19667);
and UO_1728 (O_1728,N_19646,N_19582);
nand UO_1729 (O_1729,N_19668,N_19600);
xnor UO_1730 (O_1730,N_19815,N_19735);
or UO_1731 (O_1731,N_19613,N_19504);
or UO_1732 (O_1732,N_19664,N_19553);
xor UO_1733 (O_1733,N_19930,N_19845);
and UO_1734 (O_1734,N_19773,N_19795);
nand UO_1735 (O_1735,N_19542,N_19552);
xor UO_1736 (O_1736,N_19830,N_19784);
nor UO_1737 (O_1737,N_19775,N_19851);
nand UO_1738 (O_1738,N_19943,N_19628);
and UO_1739 (O_1739,N_19992,N_19556);
and UO_1740 (O_1740,N_19639,N_19590);
nand UO_1741 (O_1741,N_19549,N_19878);
xnor UO_1742 (O_1742,N_19789,N_19895);
nand UO_1743 (O_1743,N_19801,N_19695);
xnor UO_1744 (O_1744,N_19691,N_19664);
and UO_1745 (O_1745,N_19895,N_19652);
nor UO_1746 (O_1746,N_19797,N_19553);
and UO_1747 (O_1747,N_19635,N_19993);
or UO_1748 (O_1748,N_19868,N_19955);
or UO_1749 (O_1749,N_19892,N_19895);
xnor UO_1750 (O_1750,N_19527,N_19914);
nor UO_1751 (O_1751,N_19924,N_19890);
and UO_1752 (O_1752,N_19733,N_19864);
or UO_1753 (O_1753,N_19874,N_19520);
nor UO_1754 (O_1754,N_19830,N_19808);
nand UO_1755 (O_1755,N_19516,N_19701);
or UO_1756 (O_1756,N_19625,N_19676);
or UO_1757 (O_1757,N_19759,N_19638);
nor UO_1758 (O_1758,N_19911,N_19556);
and UO_1759 (O_1759,N_19630,N_19976);
nand UO_1760 (O_1760,N_19957,N_19634);
xor UO_1761 (O_1761,N_19839,N_19665);
nor UO_1762 (O_1762,N_19734,N_19575);
or UO_1763 (O_1763,N_19503,N_19723);
nand UO_1764 (O_1764,N_19622,N_19819);
xor UO_1765 (O_1765,N_19744,N_19725);
and UO_1766 (O_1766,N_19851,N_19750);
nor UO_1767 (O_1767,N_19761,N_19870);
xnor UO_1768 (O_1768,N_19952,N_19657);
and UO_1769 (O_1769,N_19755,N_19577);
nor UO_1770 (O_1770,N_19934,N_19518);
or UO_1771 (O_1771,N_19628,N_19742);
nor UO_1772 (O_1772,N_19920,N_19515);
nand UO_1773 (O_1773,N_19959,N_19576);
nor UO_1774 (O_1774,N_19955,N_19937);
nor UO_1775 (O_1775,N_19911,N_19922);
nor UO_1776 (O_1776,N_19578,N_19647);
xnor UO_1777 (O_1777,N_19644,N_19615);
xor UO_1778 (O_1778,N_19613,N_19657);
xor UO_1779 (O_1779,N_19708,N_19736);
and UO_1780 (O_1780,N_19934,N_19999);
xor UO_1781 (O_1781,N_19508,N_19995);
or UO_1782 (O_1782,N_19835,N_19578);
nor UO_1783 (O_1783,N_19522,N_19712);
and UO_1784 (O_1784,N_19960,N_19959);
xor UO_1785 (O_1785,N_19866,N_19617);
and UO_1786 (O_1786,N_19521,N_19617);
nor UO_1787 (O_1787,N_19904,N_19710);
nand UO_1788 (O_1788,N_19702,N_19853);
or UO_1789 (O_1789,N_19571,N_19642);
nor UO_1790 (O_1790,N_19727,N_19969);
nand UO_1791 (O_1791,N_19721,N_19654);
and UO_1792 (O_1792,N_19592,N_19824);
nand UO_1793 (O_1793,N_19590,N_19608);
or UO_1794 (O_1794,N_19599,N_19941);
nand UO_1795 (O_1795,N_19776,N_19551);
nand UO_1796 (O_1796,N_19707,N_19613);
nand UO_1797 (O_1797,N_19950,N_19715);
xnor UO_1798 (O_1798,N_19620,N_19653);
xnor UO_1799 (O_1799,N_19660,N_19986);
or UO_1800 (O_1800,N_19619,N_19827);
nor UO_1801 (O_1801,N_19554,N_19911);
xor UO_1802 (O_1802,N_19711,N_19719);
and UO_1803 (O_1803,N_19543,N_19994);
nand UO_1804 (O_1804,N_19988,N_19919);
and UO_1805 (O_1805,N_19570,N_19840);
and UO_1806 (O_1806,N_19691,N_19654);
xnor UO_1807 (O_1807,N_19705,N_19526);
xor UO_1808 (O_1808,N_19515,N_19968);
nand UO_1809 (O_1809,N_19652,N_19679);
nand UO_1810 (O_1810,N_19652,N_19856);
nor UO_1811 (O_1811,N_19931,N_19982);
xnor UO_1812 (O_1812,N_19789,N_19551);
nor UO_1813 (O_1813,N_19716,N_19856);
nand UO_1814 (O_1814,N_19970,N_19757);
nor UO_1815 (O_1815,N_19685,N_19759);
xnor UO_1816 (O_1816,N_19802,N_19671);
xor UO_1817 (O_1817,N_19833,N_19927);
and UO_1818 (O_1818,N_19755,N_19742);
nand UO_1819 (O_1819,N_19961,N_19836);
and UO_1820 (O_1820,N_19614,N_19985);
nor UO_1821 (O_1821,N_19896,N_19683);
and UO_1822 (O_1822,N_19944,N_19862);
or UO_1823 (O_1823,N_19574,N_19938);
and UO_1824 (O_1824,N_19612,N_19689);
or UO_1825 (O_1825,N_19529,N_19954);
nor UO_1826 (O_1826,N_19693,N_19777);
nor UO_1827 (O_1827,N_19960,N_19859);
or UO_1828 (O_1828,N_19591,N_19859);
xor UO_1829 (O_1829,N_19743,N_19905);
nand UO_1830 (O_1830,N_19620,N_19645);
and UO_1831 (O_1831,N_19668,N_19961);
nor UO_1832 (O_1832,N_19931,N_19991);
and UO_1833 (O_1833,N_19971,N_19569);
nor UO_1834 (O_1834,N_19917,N_19621);
nand UO_1835 (O_1835,N_19554,N_19530);
nand UO_1836 (O_1836,N_19608,N_19982);
nand UO_1837 (O_1837,N_19919,N_19914);
xnor UO_1838 (O_1838,N_19718,N_19796);
nand UO_1839 (O_1839,N_19579,N_19528);
and UO_1840 (O_1840,N_19819,N_19510);
xor UO_1841 (O_1841,N_19670,N_19687);
nand UO_1842 (O_1842,N_19503,N_19999);
and UO_1843 (O_1843,N_19660,N_19578);
and UO_1844 (O_1844,N_19634,N_19887);
and UO_1845 (O_1845,N_19603,N_19582);
xor UO_1846 (O_1846,N_19698,N_19997);
nor UO_1847 (O_1847,N_19970,N_19533);
nand UO_1848 (O_1848,N_19948,N_19734);
xnor UO_1849 (O_1849,N_19836,N_19585);
or UO_1850 (O_1850,N_19685,N_19788);
xnor UO_1851 (O_1851,N_19924,N_19556);
and UO_1852 (O_1852,N_19532,N_19942);
nand UO_1853 (O_1853,N_19578,N_19564);
xor UO_1854 (O_1854,N_19976,N_19942);
or UO_1855 (O_1855,N_19791,N_19521);
xor UO_1856 (O_1856,N_19707,N_19603);
and UO_1857 (O_1857,N_19752,N_19805);
nor UO_1858 (O_1858,N_19825,N_19944);
or UO_1859 (O_1859,N_19781,N_19886);
nand UO_1860 (O_1860,N_19945,N_19633);
nor UO_1861 (O_1861,N_19650,N_19535);
nor UO_1862 (O_1862,N_19646,N_19628);
xor UO_1863 (O_1863,N_19788,N_19954);
xor UO_1864 (O_1864,N_19771,N_19733);
or UO_1865 (O_1865,N_19975,N_19706);
xor UO_1866 (O_1866,N_19951,N_19851);
xor UO_1867 (O_1867,N_19972,N_19591);
or UO_1868 (O_1868,N_19698,N_19923);
xor UO_1869 (O_1869,N_19805,N_19666);
xnor UO_1870 (O_1870,N_19631,N_19562);
or UO_1871 (O_1871,N_19535,N_19816);
or UO_1872 (O_1872,N_19897,N_19700);
nand UO_1873 (O_1873,N_19818,N_19758);
and UO_1874 (O_1874,N_19793,N_19861);
nor UO_1875 (O_1875,N_19985,N_19563);
nor UO_1876 (O_1876,N_19806,N_19612);
and UO_1877 (O_1877,N_19912,N_19726);
nand UO_1878 (O_1878,N_19539,N_19680);
or UO_1879 (O_1879,N_19895,N_19693);
nor UO_1880 (O_1880,N_19566,N_19694);
or UO_1881 (O_1881,N_19882,N_19542);
or UO_1882 (O_1882,N_19798,N_19925);
and UO_1883 (O_1883,N_19978,N_19761);
xnor UO_1884 (O_1884,N_19590,N_19506);
xnor UO_1885 (O_1885,N_19880,N_19540);
or UO_1886 (O_1886,N_19587,N_19607);
and UO_1887 (O_1887,N_19676,N_19630);
nor UO_1888 (O_1888,N_19987,N_19560);
and UO_1889 (O_1889,N_19568,N_19816);
and UO_1890 (O_1890,N_19748,N_19809);
nand UO_1891 (O_1891,N_19916,N_19969);
or UO_1892 (O_1892,N_19930,N_19871);
and UO_1893 (O_1893,N_19720,N_19729);
and UO_1894 (O_1894,N_19815,N_19500);
and UO_1895 (O_1895,N_19504,N_19529);
nor UO_1896 (O_1896,N_19980,N_19514);
nor UO_1897 (O_1897,N_19771,N_19858);
nor UO_1898 (O_1898,N_19942,N_19697);
and UO_1899 (O_1899,N_19627,N_19639);
or UO_1900 (O_1900,N_19975,N_19527);
nand UO_1901 (O_1901,N_19891,N_19989);
xnor UO_1902 (O_1902,N_19676,N_19680);
nor UO_1903 (O_1903,N_19866,N_19867);
or UO_1904 (O_1904,N_19925,N_19742);
xor UO_1905 (O_1905,N_19868,N_19720);
nor UO_1906 (O_1906,N_19816,N_19880);
nor UO_1907 (O_1907,N_19721,N_19709);
and UO_1908 (O_1908,N_19650,N_19991);
nor UO_1909 (O_1909,N_19960,N_19877);
and UO_1910 (O_1910,N_19837,N_19711);
or UO_1911 (O_1911,N_19554,N_19932);
or UO_1912 (O_1912,N_19602,N_19839);
xor UO_1913 (O_1913,N_19709,N_19627);
nor UO_1914 (O_1914,N_19877,N_19556);
xor UO_1915 (O_1915,N_19686,N_19627);
or UO_1916 (O_1916,N_19756,N_19966);
or UO_1917 (O_1917,N_19755,N_19642);
or UO_1918 (O_1918,N_19501,N_19787);
and UO_1919 (O_1919,N_19683,N_19663);
nand UO_1920 (O_1920,N_19709,N_19706);
and UO_1921 (O_1921,N_19721,N_19642);
and UO_1922 (O_1922,N_19598,N_19844);
nor UO_1923 (O_1923,N_19911,N_19665);
xor UO_1924 (O_1924,N_19999,N_19544);
nor UO_1925 (O_1925,N_19718,N_19776);
nor UO_1926 (O_1926,N_19722,N_19834);
nor UO_1927 (O_1927,N_19857,N_19598);
and UO_1928 (O_1928,N_19877,N_19860);
and UO_1929 (O_1929,N_19948,N_19888);
or UO_1930 (O_1930,N_19678,N_19726);
and UO_1931 (O_1931,N_19773,N_19525);
xnor UO_1932 (O_1932,N_19537,N_19933);
or UO_1933 (O_1933,N_19757,N_19858);
xor UO_1934 (O_1934,N_19853,N_19503);
or UO_1935 (O_1935,N_19945,N_19662);
xor UO_1936 (O_1936,N_19824,N_19697);
and UO_1937 (O_1937,N_19826,N_19728);
nor UO_1938 (O_1938,N_19680,N_19681);
xnor UO_1939 (O_1939,N_19971,N_19500);
nor UO_1940 (O_1940,N_19982,N_19574);
nor UO_1941 (O_1941,N_19782,N_19906);
nand UO_1942 (O_1942,N_19923,N_19839);
nor UO_1943 (O_1943,N_19768,N_19502);
and UO_1944 (O_1944,N_19543,N_19644);
and UO_1945 (O_1945,N_19743,N_19798);
or UO_1946 (O_1946,N_19833,N_19681);
and UO_1947 (O_1947,N_19871,N_19948);
nand UO_1948 (O_1948,N_19849,N_19661);
and UO_1949 (O_1949,N_19985,N_19649);
or UO_1950 (O_1950,N_19936,N_19839);
xor UO_1951 (O_1951,N_19708,N_19631);
nor UO_1952 (O_1952,N_19893,N_19989);
nand UO_1953 (O_1953,N_19707,N_19845);
nor UO_1954 (O_1954,N_19926,N_19746);
nor UO_1955 (O_1955,N_19687,N_19945);
xnor UO_1956 (O_1956,N_19903,N_19735);
or UO_1957 (O_1957,N_19696,N_19593);
nand UO_1958 (O_1958,N_19730,N_19866);
nor UO_1959 (O_1959,N_19530,N_19504);
and UO_1960 (O_1960,N_19636,N_19966);
nor UO_1961 (O_1961,N_19867,N_19926);
nor UO_1962 (O_1962,N_19620,N_19876);
or UO_1963 (O_1963,N_19718,N_19853);
or UO_1964 (O_1964,N_19730,N_19859);
xnor UO_1965 (O_1965,N_19618,N_19572);
nor UO_1966 (O_1966,N_19517,N_19634);
and UO_1967 (O_1967,N_19680,N_19837);
nand UO_1968 (O_1968,N_19908,N_19537);
nor UO_1969 (O_1969,N_19574,N_19746);
nor UO_1970 (O_1970,N_19853,N_19975);
nor UO_1971 (O_1971,N_19882,N_19741);
nand UO_1972 (O_1972,N_19710,N_19670);
nor UO_1973 (O_1973,N_19952,N_19581);
and UO_1974 (O_1974,N_19773,N_19613);
or UO_1975 (O_1975,N_19788,N_19653);
xor UO_1976 (O_1976,N_19809,N_19732);
nor UO_1977 (O_1977,N_19647,N_19857);
nand UO_1978 (O_1978,N_19673,N_19878);
nor UO_1979 (O_1979,N_19767,N_19882);
nor UO_1980 (O_1980,N_19594,N_19769);
xnor UO_1981 (O_1981,N_19824,N_19747);
nor UO_1982 (O_1982,N_19518,N_19796);
nand UO_1983 (O_1983,N_19975,N_19566);
xor UO_1984 (O_1984,N_19790,N_19882);
nor UO_1985 (O_1985,N_19827,N_19891);
and UO_1986 (O_1986,N_19532,N_19618);
and UO_1987 (O_1987,N_19944,N_19902);
and UO_1988 (O_1988,N_19507,N_19632);
nor UO_1989 (O_1989,N_19782,N_19926);
and UO_1990 (O_1990,N_19534,N_19834);
xor UO_1991 (O_1991,N_19952,N_19508);
and UO_1992 (O_1992,N_19758,N_19861);
nor UO_1993 (O_1993,N_19595,N_19560);
or UO_1994 (O_1994,N_19664,N_19997);
nor UO_1995 (O_1995,N_19760,N_19536);
nand UO_1996 (O_1996,N_19861,N_19701);
nand UO_1997 (O_1997,N_19955,N_19668);
nand UO_1998 (O_1998,N_19628,N_19834);
nand UO_1999 (O_1999,N_19989,N_19623);
xor UO_2000 (O_2000,N_19752,N_19818);
or UO_2001 (O_2001,N_19587,N_19677);
nor UO_2002 (O_2002,N_19847,N_19913);
or UO_2003 (O_2003,N_19748,N_19734);
xnor UO_2004 (O_2004,N_19770,N_19752);
or UO_2005 (O_2005,N_19566,N_19876);
and UO_2006 (O_2006,N_19985,N_19595);
nor UO_2007 (O_2007,N_19872,N_19888);
nand UO_2008 (O_2008,N_19952,N_19638);
and UO_2009 (O_2009,N_19595,N_19599);
nor UO_2010 (O_2010,N_19604,N_19582);
nor UO_2011 (O_2011,N_19678,N_19779);
or UO_2012 (O_2012,N_19530,N_19735);
nor UO_2013 (O_2013,N_19668,N_19552);
or UO_2014 (O_2014,N_19900,N_19601);
nor UO_2015 (O_2015,N_19647,N_19711);
or UO_2016 (O_2016,N_19871,N_19901);
or UO_2017 (O_2017,N_19950,N_19723);
or UO_2018 (O_2018,N_19648,N_19624);
and UO_2019 (O_2019,N_19876,N_19500);
or UO_2020 (O_2020,N_19570,N_19721);
nand UO_2021 (O_2021,N_19566,N_19693);
nor UO_2022 (O_2022,N_19590,N_19816);
nor UO_2023 (O_2023,N_19893,N_19673);
nor UO_2024 (O_2024,N_19778,N_19995);
nand UO_2025 (O_2025,N_19918,N_19945);
or UO_2026 (O_2026,N_19825,N_19509);
and UO_2027 (O_2027,N_19519,N_19536);
nor UO_2028 (O_2028,N_19502,N_19981);
and UO_2029 (O_2029,N_19774,N_19645);
xnor UO_2030 (O_2030,N_19868,N_19893);
nand UO_2031 (O_2031,N_19565,N_19774);
xnor UO_2032 (O_2032,N_19817,N_19548);
nand UO_2033 (O_2033,N_19651,N_19573);
and UO_2034 (O_2034,N_19550,N_19770);
or UO_2035 (O_2035,N_19607,N_19570);
nor UO_2036 (O_2036,N_19508,N_19706);
nand UO_2037 (O_2037,N_19990,N_19870);
or UO_2038 (O_2038,N_19520,N_19834);
and UO_2039 (O_2039,N_19814,N_19575);
and UO_2040 (O_2040,N_19789,N_19784);
nor UO_2041 (O_2041,N_19963,N_19969);
nor UO_2042 (O_2042,N_19547,N_19770);
nor UO_2043 (O_2043,N_19947,N_19821);
nand UO_2044 (O_2044,N_19929,N_19899);
xor UO_2045 (O_2045,N_19807,N_19763);
nand UO_2046 (O_2046,N_19650,N_19938);
nand UO_2047 (O_2047,N_19973,N_19718);
or UO_2048 (O_2048,N_19557,N_19786);
nand UO_2049 (O_2049,N_19775,N_19627);
and UO_2050 (O_2050,N_19836,N_19595);
and UO_2051 (O_2051,N_19626,N_19778);
nand UO_2052 (O_2052,N_19970,N_19605);
and UO_2053 (O_2053,N_19808,N_19700);
and UO_2054 (O_2054,N_19770,N_19844);
nor UO_2055 (O_2055,N_19872,N_19985);
and UO_2056 (O_2056,N_19591,N_19518);
nor UO_2057 (O_2057,N_19600,N_19638);
xnor UO_2058 (O_2058,N_19588,N_19600);
nor UO_2059 (O_2059,N_19505,N_19819);
xor UO_2060 (O_2060,N_19617,N_19536);
nor UO_2061 (O_2061,N_19796,N_19991);
nor UO_2062 (O_2062,N_19815,N_19896);
and UO_2063 (O_2063,N_19930,N_19669);
xnor UO_2064 (O_2064,N_19665,N_19584);
or UO_2065 (O_2065,N_19615,N_19709);
and UO_2066 (O_2066,N_19663,N_19542);
nor UO_2067 (O_2067,N_19560,N_19798);
or UO_2068 (O_2068,N_19622,N_19686);
xnor UO_2069 (O_2069,N_19783,N_19726);
nand UO_2070 (O_2070,N_19878,N_19641);
or UO_2071 (O_2071,N_19901,N_19532);
and UO_2072 (O_2072,N_19957,N_19854);
nand UO_2073 (O_2073,N_19601,N_19985);
nand UO_2074 (O_2074,N_19569,N_19687);
and UO_2075 (O_2075,N_19949,N_19907);
xor UO_2076 (O_2076,N_19990,N_19578);
and UO_2077 (O_2077,N_19533,N_19800);
nand UO_2078 (O_2078,N_19787,N_19786);
nand UO_2079 (O_2079,N_19961,N_19946);
and UO_2080 (O_2080,N_19503,N_19680);
nor UO_2081 (O_2081,N_19901,N_19608);
nor UO_2082 (O_2082,N_19968,N_19986);
xnor UO_2083 (O_2083,N_19584,N_19903);
or UO_2084 (O_2084,N_19834,N_19514);
and UO_2085 (O_2085,N_19607,N_19907);
nand UO_2086 (O_2086,N_19682,N_19738);
xor UO_2087 (O_2087,N_19953,N_19923);
and UO_2088 (O_2088,N_19649,N_19781);
xnor UO_2089 (O_2089,N_19774,N_19603);
xnor UO_2090 (O_2090,N_19620,N_19857);
or UO_2091 (O_2091,N_19743,N_19998);
xor UO_2092 (O_2092,N_19783,N_19962);
nor UO_2093 (O_2093,N_19908,N_19823);
nor UO_2094 (O_2094,N_19540,N_19612);
and UO_2095 (O_2095,N_19940,N_19560);
nand UO_2096 (O_2096,N_19666,N_19577);
xor UO_2097 (O_2097,N_19705,N_19687);
nand UO_2098 (O_2098,N_19543,N_19975);
nor UO_2099 (O_2099,N_19878,N_19890);
nand UO_2100 (O_2100,N_19694,N_19896);
and UO_2101 (O_2101,N_19664,N_19663);
and UO_2102 (O_2102,N_19554,N_19607);
nor UO_2103 (O_2103,N_19715,N_19540);
or UO_2104 (O_2104,N_19802,N_19723);
or UO_2105 (O_2105,N_19741,N_19774);
xor UO_2106 (O_2106,N_19543,N_19929);
nand UO_2107 (O_2107,N_19679,N_19538);
nand UO_2108 (O_2108,N_19723,N_19625);
nor UO_2109 (O_2109,N_19651,N_19960);
xor UO_2110 (O_2110,N_19963,N_19624);
and UO_2111 (O_2111,N_19508,N_19909);
nand UO_2112 (O_2112,N_19665,N_19652);
nor UO_2113 (O_2113,N_19570,N_19974);
xor UO_2114 (O_2114,N_19977,N_19622);
and UO_2115 (O_2115,N_19526,N_19569);
xnor UO_2116 (O_2116,N_19514,N_19799);
nand UO_2117 (O_2117,N_19662,N_19717);
and UO_2118 (O_2118,N_19829,N_19785);
nand UO_2119 (O_2119,N_19951,N_19868);
and UO_2120 (O_2120,N_19915,N_19635);
nor UO_2121 (O_2121,N_19803,N_19952);
xor UO_2122 (O_2122,N_19569,N_19886);
nor UO_2123 (O_2123,N_19941,N_19876);
and UO_2124 (O_2124,N_19633,N_19534);
nand UO_2125 (O_2125,N_19932,N_19695);
and UO_2126 (O_2126,N_19946,N_19514);
xnor UO_2127 (O_2127,N_19711,N_19679);
and UO_2128 (O_2128,N_19628,N_19945);
xor UO_2129 (O_2129,N_19601,N_19910);
and UO_2130 (O_2130,N_19579,N_19909);
nor UO_2131 (O_2131,N_19840,N_19988);
nor UO_2132 (O_2132,N_19831,N_19870);
xnor UO_2133 (O_2133,N_19598,N_19757);
nor UO_2134 (O_2134,N_19866,N_19539);
nor UO_2135 (O_2135,N_19875,N_19702);
nand UO_2136 (O_2136,N_19959,N_19944);
nand UO_2137 (O_2137,N_19995,N_19588);
or UO_2138 (O_2138,N_19529,N_19543);
or UO_2139 (O_2139,N_19579,N_19863);
and UO_2140 (O_2140,N_19542,N_19763);
xor UO_2141 (O_2141,N_19651,N_19735);
xnor UO_2142 (O_2142,N_19972,N_19989);
xnor UO_2143 (O_2143,N_19936,N_19580);
and UO_2144 (O_2144,N_19650,N_19961);
nor UO_2145 (O_2145,N_19796,N_19581);
or UO_2146 (O_2146,N_19789,N_19867);
or UO_2147 (O_2147,N_19993,N_19781);
and UO_2148 (O_2148,N_19747,N_19759);
nor UO_2149 (O_2149,N_19884,N_19689);
and UO_2150 (O_2150,N_19670,N_19667);
xnor UO_2151 (O_2151,N_19820,N_19886);
xnor UO_2152 (O_2152,N_19539,N_19959);
nand UO_2153 (O_2153,N_19645,N_19955);
nand UO_2154 (O_2154,N_19624,N_19645);
or UO_2155 (O_2155,N_19606,N_19763);
and UO_2156 (O_2156,N_19807,N_19518);
nor UO_2157 (O_2157,N_19858,N_19638);
nor UO_2158 (O_2158,N_19822,N_19544);
nand UO_2159 (O_2159,N_19613,N_19558);
and UO_2160 (O_2160,N_19795,N_19514);
or UO_2161 (O_2161,N_19958,N_19525);
nand UO_2162 (O_2162,N_19658,N_19866);
and UO_2163 (O_2163,N_19562,N_19863);
xnor UO_2164 (O_2164,N_19984,N_19752);
nand UO_2165 (O_2165,N_19994,N_19814);
xor UO_2166 (O_2166,N_19750,N_19892);
nand UO_2167 (O_2167,N_19879,N_19544);
nor UO_2168 (O_2168,N_19739,N_19722);
nand UO_2169 (O_2169,N_19989,N_19528);
and UO_2170 (O_2170,N_19761,N_19507);
or UO_2171 (O_2171,N_19643,N_19983);
nand UO_2172 (O_2172,N_19742,N_19933);
nor UO_2173 (O_2173,N_19734,N_19826);
or UO_2174 (O_2174,N_19580,N_19937);
nor UO_2175 (O_2175,N_19566,N_19685);
or UO_2176 (O_2176,N_19812,N_19541);
or UO_2177 (O_2177,N_19740,N_19871);
xnor UO_2178 (O_2178,N_19785,N_19977);
or UO_2179 (O_2179,N_19959,N_19624);
and UO_2180 (O_2180,N_19820,N_19713);
and UO_2181 (O_2181,N_19555,N_19775);
or UO_2182 (O_2182,N_19922,N_19893);
nand UO_2183 (O_2183,N_19570,N_19648);
nand UO_2184 (O_2184,N_19672,N_19581);
nor UO_2185 (O_2185,N_19804,N_19641);
nor UO_2186 (O_2186,N_19658,N_19859);
nand UO_2187 (O_2187,N_19556,N_19543);
xnor UO_2188 (O_2188,N_19530,N_19543);
and UO_2189 (O_2189,N_19701,N_19528);
nand UO_2190 (O_2190,N_19909,N_19700);
xnor UO_2191 (O_2191,N_19882,N_19711);
nand UO_2192 (O_2192,N_19718,N_19657);
and UO_2193 (O_2193,N_19941,N_19844);
or UO_2194 (O_2194,N_19817,N_19582);
and UO_2195 (O_2195,N_19851,N_19664);
or UO_2196 (O_2196,N_19507,N_19631);
nor UO_2197 (O_2197,N_19692,N_19545);
or UO_2198 (O_2198,N_19636,N_19808);
nand UO_2199 (O_2199,N_19650,N_19686);
nor UO_2200 (O_2200,N_19997,N_19687);
nor UO_2201 (O_2201,N_19655,N_19534);
and UO_2202 (O_2202,N_19960,N_19963);
and UO_2203 (O_2203,N_19682,N_19582);
xnor UO_2204 (O_2204,N_19855,N_19533);
and UO_2205 (O_2205,N_19660,N_19866);
or UO_2206 (O_2206,N_19527,N_19605);
nand UO_2207 (O_2207,N_19922,N_19507);
and UO_2208 (O_2208,N_19938,N_19655);
or UO_2209 (O_2209,N_19675,N_19863);
and UO_2210 (O_2210,N_19537,N_19678);
xnor UO_2211 (O_2211,N_19939,N_19779);
nor UO_2212 (O_2212,N_19802,N_19601);
nor UO_2213 (O_2213,N_19741,N_19778);
xnor UO_2214 (O_2214,N_19520,N_19660);
xor UO_2215 (O_2215,N_19527,N_19686);
or UO_2216 (O_2216,N_19776,N_19988);
nor UO_2217 (O_2217,N_19881,N_19593);
and UO_2218 (O_2218,N_19866,N_19808);
and UO_2219 (O_2219,N_19770,N_19525);
or UO_2220 (O_2220,N_19639,N_19612);
and UO_2221 (O_2221,N_19589,N_19726);
xnor UO_2222 (O_2222,N_19564,N_19634);
nor UO_2223 (O_2223,N_19722,N_19833);
and UO_2224 (O_2224,N_19861,N_19857);
and UO_2225 (O_2225,N_19800,N_19572);
or UO_2226 (O_2226,N_19936,N_19699);
or UO_2227 (O_2227,N_19604,N_19861);
xnor UO_2228 (O_2228,N_19851,N_19571);
nand UO_2229 (O_2229,N_19933,N_19791);
and UO_2230 (O_2230,N_19924,N_19674);
or UO_2231 (O_2231,N_19641,N_19961);
nor UO_2232 (O_2232,N_19589,N_19565);
xnor UO_2233 (O_2233,N_19946,N_19770);
nor UO_2234 (O_2234,N_19672,N_19755);
and UO_2235 (O_2235,N_19746,N_19548);
and UO_2236 (O_2236,N_19991,N_19584);
nor UO_2237 (O_2237,N_19672,N_19884);
or UO_2238 (O_2238,N_19598,N_19773);
nand UO_2239 (O_2239,N_19759,N_19640);
or UO_2240 (O_2240,N_19871,N_19621);
nor UO_2241 (O_2241,N_19948,N_19542);
nor UO_2242 (O_2242,N_19718,N_19917);
xor UO_2243 (O_2243,N_19977,N_19775);
and UO_2244 (O_2244,N_19564,N_19989);
nor UO_2245 (O_2245,N_19932,N_19601);
nor UO_2246 (O_2246,N_19603,N_19892);
and UO_2247 (O_2247,N_19635,N_19504);
xor UO_2248 (O_2248,N_19839,N_19703);
or UO_2249 (O_2249,N_19770,N_19567);
nand UO_2250 (O_2250,N_19588,N_19637);
or UO_2251 (O_2251,N_19523,N_19506);
and UO_2252 (O_2252,N_19718,N_19827);
or UO_2253 (O_2253,N_19926,N_19706);
and UO_2254 (O_2254,N_19602,N_19983);
nand UO_2255 (O_2255,N_19826,N_19888);
nand UO_2256 (O_2256,N_19890,N_19897);
nor UO_2257 (O_2257,N_19677,N_19744);
nor UO_2258 (O_2258,N_19890,N_19543);
or UO_2259 (O_2259,N_19904,N_19865);
nand UO_2260 (O_2260,N_19693,N_19607);
xor UO_2261 (O_2261,N_19627,N_19691);
nor UO_2262 (O_2262,N_19901,N_19745);
or UO_2263 (O_2263,N_19689,N_19573);
nor UO_2264 (O_2264,N_19636,N_19707);
and UO_2265 (O_2265,N_19657,N_19956);
and UO_2266 (O_2266,N_19853,N_19839);
or UO_2267 (O_2267,N_19965,N_19571);
or UO_2268 (O_2268,N_19963,N_19751);
xnor UO_2269 (O_2269,N_19824,N_19879);
nor UO_2270 (O_2270,N_19642,N_19648);
and UO_2271 (O_2271,N_19774,N_19619);
xnor UO_2272 (O_2272,N_19829,N_19663);
nor UO_2273 (O_2273,N_19520,N_19727);
and UO_2274 (O_2274,N_19802,N_19710);
and UO_2275 (O_2275,N_19931,N_19654);
or UO_2276 (O_2276,N_19631,N_19873);
nand UO_2277 (O_2277,N_19752,N_19563);
or UO_2278 (O_2278,N_19647,N_19594);
xor UO_2279 (O_2279,N_19924,N_19680);
or UO_2280 (O_2280,N_19645,N_19971);
xnor UO_2281 (O_2281,N_19784,N_19863);
nor UO_2282 (O_2282,N_19915,N_19970);
and UO_2283 (O_2283,N_19875,N_19613);
or UO_2284 (O_2284,N_19978,N_19795);
or UO_2285 (O_2285,N_19631,N_19515);
xor UO_2286 (O_2286,N_19637,N_19933);
nor UO_2287 (O_2287,N_19728,N_19530);
xnor UO_2288 (O_2288,N_19824,N_19669);
xnor UO_2289 (O_2289,N_19943,N_19952);
or UO_2290 (O_2290,N_19516,N_19700);
nand UO_2291 (O_2291,N_19703,N_19890);
and UO_2292 (O_2292,N_19839,N_19806);
or UO_2293 (O_2293,N_19520,N_19903);
nor UO_2294 (O_2294,N_19987,N_19531);
nand UO_2295 (O_2295,N_19917,N_19854);
nor UO_2296 (O_2296,N_19613,N_19925);
nand UO_2297 (O_2297,N_19589,N_19637);
nor UO_2298 (O_2298,N_19964,N_19970);
or UO_2299 (O_2299,N_19696,N_19690);
nor UO_2300 (O_2300,N_19773,N_19828);
xnor UO_2301 (O_2301,N_19985,N_19575);
xnor UO_2302 (O_2302,N_19699,N_19548);
xnor UO_2303 (O_2303,N_19864,N_19798);
nand UO_2304 (O_2304,N_19611,N_19574);
and UO_2305 (O_2305,N_19841,N_19837);
nor UO_2306 (O_2306,N_19967,N_19923);
nand UO_2307 (O_2307,N_19783,N_19596);
nand UO_2308 (O_2308,N_19930,N_19825);
xnor UO_2309 (O_2309,N_19770,N_19706);
and UO_2310 (O_2310,N_19869,N_19953);
or UO_2311 (O_2311,N_19821,N_19554);
or UO_2312 (O_2312,N_19781,N_19973);
xor UO_2313 (O_2313,N_19701,N_19888);
xnor UO_2314 (O_2314,N_19916,N_19829);
xnor UO_2315 (O_2315,N_19740,N_19695);
or UO_2316 (O_2316,N_19509,N_19725);
and UO_2317 (O_2317,N_19767,N_19569);
and UO_2318 (O_2318,N_19720,N_19528);
xnor UO_2319 (O_2319,N_19939,N_19865);
and UO_2320 (O_2320,N_19734,N_19780);
xnor UO_2321 (O_2321,N_19613,N_19740);
nor UO_2322 (O_2322,N_19598,N_19543);
nand UO_2323 (O_2323,N_19506,N_19932);
nor UO_2324 (O_2324,N_19766,N_19882);
or UO_2325 (O_2325,N_19580,N_19732);
or UO_2326 (O_2326,N_19511,N_19934);
nand UO_2327 (O_2327,N_19663,N_19572);
nor UO_2328 (O_2328,N_19946,N_19664);
nand UO_2329 (O_2329,N_19580,N_19884);
nand UO_2330 (O_2330,N_19639,N_19710);
xor UO_2331 (O_2331,N_19790,N_19966);
and UO_2332 (O_2332,N_19879,N_19792);
nand UO_2333 (O_2333,N_19609,N_19807);
xnor UO_2334 (O_2334,N_19531,N_19993);
and UO_2335 (O_2335,N_19930,N_19613);
and UO_2336 (O_2336,N_19601,N_19661);
xnor UO_2337 (O_2337,N_19699,N_19675);
xnor UO_2338 (O_2338,N_19653,N_19894);
and UO_2339 (O_2339,N_19759,N_19847);
nand UO_2340 (O_2340,N_19635,N_19682);
xnor UO_2341 (O_2341,N_19945,N_19882);
xnor UO_2342 (O_2342,N_19621,N_19927);
nand UO_2343 (O_2343,N_19573,N_19843);
and UO_2344 (O_2344,N_19989,N_19881);
xor UO_2345 (O_2345,N_19758,N_19914);
and UO_2346 (O_2346,N_19530,N_19797);
nand UO_2347 (O_2347,N_19681,N_19639);
xnor UO_2348 (O_2348,N_19946,N_19907);
nand UO_2349 (O_2349,N_19994,N_19711);
nand UO_2350 (O_2350,N_19732,N_19615);
xnor UO_2351 (O_2351,N_19954,N_19693);
nor UO_2352 (O_2352,N_19521,N_19606);
nor UO_2353 (O_2353,N_19662,N_19622);
or UO_2354 (O_2354,N_19615,N_19557);
or UO_2355 (O_2355,N_19566,N_19625);
or UO_2356 (O_2356,N_19516,N_19901);
and UO_2357 (O_2357,N_19914,N_19667);
xor UO_2358 (O_2358,N_19978,N_19666);
xor UO_2359 (O_2359,N_19535,N_19521);
xnor UO_2360 (O_2360,N_19707,N_19850);
and UO_2361 (O_2361,N_19597,N_19984);
nor UO_2362 (O_2362,N_19628,N_19501);
or UO_2363 (O_2363,N_19842,N_19959);
nor UO_2364 (O_2364,N_19710,N_19617);
nand UO_2365 (O_2365,N_19890,N_19682);
and UO_2366 (O_2366,N_19971,N_19665);
and UO_2367 (O_2367,N_19965,N_19540);
nor UO_2368 (O_2368,N_19684,N_19927);
and UO_2369 (O_2369,N_19685,N_19870);
nand UO_2370 (O_2370,N_19918,N_19950);
xnor UO_2371 (O_2371,N_19729,N_19724);
nand UO_2372 (O_2372,N_19509,N_19941);
nand UO_2373 (O_2373,N_19956,N_19915);
and UO_2374 (O_2374,N_19922,N_19921);
or UO_2375 (O_2375,N_19828,N_19968);
xor UO_2376 (O_2376,N_19697,N_19962);
nand UO_2377 (O_2377,N_19673,N_19520);
nand UO_2378 (O_2378,N_19638,N_19869);
nor UO_2379 (O_2379,N_19762,N_19750);
nor UO_2380 (O_2380,N_19804,N_19958);
nor UO_2381 (O_2381,N_19663,N_19591);
nor UO_2382 (O_2382,N_19755,N_19771);
nor UO_2383 (O_2383,N_19685,N_19575);
nor UO_2384 (O_2384,N_19828,N_19887);
or UO_2385 (O_2385,N_19954,N_19605);
nand UO_2386 (O_2386,N_19506,N_19623);
nor UO_2387 (O_2387,N_19753,N_19671);
or UO_2388 (O_2388,N_19944,N_19534);
nand UO_2389 (O_2389,N_19958,N_19564);
nand UO_2390 (O_2390,N_19856,N_19524);
and UO_2391 (O_2391,N_19549,N_19873);
or UO_2392 (O_2392,N_19747,N_19896);
xor UO_2393 (O_2393,N_19929,N_19603);
nand UO_2394 (O_2394,N_19908,N_19960);
nand UO_2395 (O_2395,N_19825,N_19974);
or UO_2396 (O_2396,N_19951,N_19565);
nor UO_2397 (O_2397,N_19511,N_19578);
or UO_2398 (O_2398,N_19718,N_19923);
nor UO_2399 (O_2399,N_19565,N_19526);
nand UO_2400 (O_2400,N_19803,N_19505);
xnor UO_2401 (O_2401,N_19755,N_19812);
or UO_2402 (O_2402,N_19572,N_19939);
and UO_2403 (O_2403,N_19735,N_19818);
xnor UO_2404 (O_2404,N_19974,N_19911);
nand UO_2405 (O_2405,N_19773,N_19584);
or UO_2406 (O_2406,N_19637,N_19740);
nand UO_2407 (O_2407,N_19763,N_19572);
and UO_2408 (O_2408,N_19863,N_19972);
nand UO_2409 (O_2409,N_19767,N_19544);
xor UO_2410 (O_2410,N_19741,N_19860);
or UO_2411 (O_2411,N_19829,N_19748);
xnor UO_2412 (O_2412,N_19548,N_19823);
or UO_2413 (O_2413,N_19800,N_19699);
nor UO_2414 (O_2414,N_19825,N_19609);
nor UO_2415 (O_2415,N_19517,N_19678);
xnor UO_2416 (O_2416,N_19685,N_19967);
nor UO_2417 (O_2417,N_19988,N_19948);
and UO_2418 (O_2418,N_19969,N_19539);
and UO_2419 (O_2419,N_19690,N_19781);
xnor UO_2420 (O_2420,N_19511,N_19583);
and UO_2421 (O_2421,N_19572,N_19831);
xnor UO_2422 (O_2422,N_19780,N_19778);
nor UO_2423 (O_2423,N_19786,N_19790);
xnor UO_2424 (O_2424,N_19736,N_19667);
xnor UO_2425 (O_2425,N_19917,N_19978);
nor UO_2426 (O_2426,N_19820,N_19681);
nand UO_2427 (O_2427,N_19611,N_19521);
nor UO_2428 (O_2428,N_19988,N_19714);
and UO_2429 (O_2429,N_19714,N_19796);
xor UO_2430 (O_2430,N_19866,N_19676);
nor UO_2431 (O_2431,N_19991,N_19594);
nor UO_2432 (O_2432,N_19975,N_19667);
or UO_2433 (O_2433,N_19584,N_19977);
nor UO_2434 (O_2434,N_19598,N_19708);
nor UO_2435 (O_2435,N_19564,N_19545);
xnor UO_2436 (O_2436,N_19741,N_19798);
or UO_2437 (O_2437,N_19741,N_19724);
nand UO_2438 (O_2438,N_19674,N_19773);
nor UO_2439 (O_2439,N_19868,N_19563);
nand UO_2440 (O_2440,N_19735,N_19525);
xnor UO_2441 (O_2441,N_19775,N_19661);
and UO_2442 (O_2442,N_19526,N_19851);
and UO_2443 (O_2443,N_19690,N_19635);
xor UO_2444 (O_2444,N_19564,N_19536);
nand UO_2445 (O_2445,N_19996,N_19890);
nand UO_2446 (O_2446,N_19726,N_19784);
xnor UO_2447 (O_2447,N_19592,N_19662);
and UO_2448 (O_2448,N_19983,N_19840);
or UO_2449 (O_2449,N_19725,N_19561);
or UO_2450 (O_2450,N_19681,N_19682);
nand UO_2451 (O_2451,N_19837,N_19974);
xnor UO_2452 (O_2452,N_19624,N_19721);
nor UO_2453 (O_2453,N_19901,N_19755);
nand UO_2454 (O_2454,N_19789,N_19779);
or UO_2455 (O_2455,N_19659,N_19864);
nor UO_2456 (O_2456,N_19680,N_19624);
or UO_2457 (O_2457,N_19627,N_19756);
nand UO_2458 (O_2458,N_19724,N_19900);
xor UO_2459 (O_2459,N_19663,N_19758);
xor UO_2460 (O_2460,N_19625,N_19814);
and UO_2461 (O_2461,N_19936,N_19728);
and UO_2462 (O_2462,N_19552,N_19762);
and UO_2463 (O_2463,N_19975,N_19632);
xnor UO_2464 (O_2464,N_19581,N_19732);
and UO_2465 (O_2465,N_19689,N_19569);
nand UO_2466 (O_2466,N_19743,N_19842);
nand UO_2467 (O_2467,N_19585,N_19526);
xor UO_2468 (O_2468,N_19591,N_19664);
or UO_2469 (O_2469,N_19874,N_19592);
nor UO_2470 (O_2470,N_19624,N_19705);
xor UO_2471 (O_2471,N_19546,N_19718);
or UO_2472 (O_2472,N_19896,N_19615);
and UO_2473 (O_2473,N_19509,N_19996);
nor UO_2474 (O_2474,N_19983,N_19868);
xnor UO_2475 (O_2475,N_19900,N_19711);
xor UO_2476 (O_2476,N_19860,N_19946);
and UO_2477 (O_2477,N_19725,N_19851);
and UO_2478 (O_2478,N_19741,N_19847);
nand UO_2479 (O_2479,N_19560,N_19653);
nor UO_2480 (O_2480,N_19573,N_19855);
nand UO_2481 (O_2481,N_19959,N_19825);
nor UO_2482 (O_2482,N_19572,N_19793);
nand UO_2483 (O_2483,N_19510,N_19734);
nor UO_2484 (O_2484,N_19993,N_19981);
nor UO_2485 (O_2485,N_19914,N_19660);
nor UO_2486 (O_2486,N_19882,N_19540);
xor UO_2487 (O_2487,N_19653,N_19678);
nand UO_2488 (O_2488,N_19661,N_19894);
or UO_2489 (O_2489,N_19693,N_19554);
nand UO_2490 (O_2490,N_19971,N_19814);
nand UO_2491 (O_2491,N_19987,N_19649);
nor UO_2492 (O_2492,N_19647,N_19911);
nand UO_2493 (O_2493,N_19909,N_19688);
and UO_2494 (O_2494,N_19804,N_19702);
nor UO_2495 (O_2495,N_19740,N_19798);
or UO_2496 (O_2496,N_19885,N_19811);
nand UO_2497 (O_2497,N_19687,N_19806);
or UO_2498 (O_2498,N_19785,N_19983);
or UO_2499 (O_2499,N_19919,N_19857);
endmodule