module basic_500_3000_500_30_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_206,In_338);
and U1 (N_1,In_377,In_182);
nor U2 (N_2,In_65,In_410);
or U3 (N_3,In_282,In_96);
and U4 (N_4,In_134,In_184);
or U5 (N_5,In_121,In_496);
nand U6 (N_6,In_268,In_439);
or U7 (N_7,In_205,In_316);
and U8 (N_8,In_10,In_324);
or U9 (N_9,In_331,In_80);
nand U10 (N_10,In_306,In_44);
nand U11 (N_11,In_84,In_265);
and U12 (N_12,In_144,In_11);
or U13 (N_13,In_187,In_7);
or U14 (N_14,In_363,In_153);
and U15 (N_15,In_88,In_118);
or U16 (N_16,In_178,In_6);
nor U17 (N_17,In_87,In_450);
or U18 (N_18,In_440,In_26);
nor U19 (N_19,In_287,In_434);
nand U20 (N_20,In_381,In_412);
nor U21 (N_21,In_365,In_48);
nand U22 (N_22,In_111,In_261);
or U23 (N_23,In_358,In_202);
nand U24 (N_24,In_300,In_173);
nand U25 (N_25,In_57,In_379);
and U26 (N_26,In_176,In_14);
nand U27 (N_27,In_46,In_321);
nor U28 (N_28,In_226,In_390);
nand U29 (N_29,In_426,In_47);
nor U30 (N_30,In_114,In_483);
nand U31 (N_31,In_384,In_0);
xnor U32 (N_32,In_462,In_104);
or U33 (N_33,In_154,In_78);
and U34 (N_34,In_13,In_168);
xnor U35 (N_35,In_214,In_255);
nor U36 (N_36,In_459,In_245);
or U37 (N_37,In_479,In_186);
and U38 (N_38,In_396,In_53);
nand U39 (N_39,In_467,In_119);
nand U40 (N_40,In_42,In_297);
nor U41 (N_41,In_130,In_123);
nor U42 (N_42,In_352,In_110);
nor U43 (N_43,In_313,In_108);
and U44 (N_44,In_120,In_422);
and U45 (N_45,In_376,In_49);
or U46 (N_46,In_256,In_429);
and U47 (N_47,In_498,In_107);
or U48 (N_48,In_50,In_356);
and U49 (N_49,In_436,In_102);
nand U50 (N_50,In_399,In_308);
nand U51 (N_51,In_12,In_418);
nand U52 (N_52,In_335,In_4);
and U53 (N_53,In_407,In_470);
nor U54 (N_54,In_425,In_194);
or U55 (N_55,In_38,In_257);
and U56 (N_56,In_275,In_203);
nor U57 (N_57,In_149,In_269);
nor U58 (N_58,In_368,In_162);
nor U59 (N_59,In_366,In_159);
nor U60 (N_60,In_69,In_473);
nand U61 (N_61,In_132,In_145);
nor U62 (N_62,In_171,In_112);
or U63 (N_63,In_315,In_83);
and U64 (N_64,In_322,In_235);
or U65 (N_65,In_264,In_99);
nand U66 (N_66,In_451,In_273);
nand U67 (N_67,In_125,In_304);
nor U68 (N_68,In_183,In_337);
and U69 (N_69,In_457,In_452);
nand U70 (N_70,In_391,In_63);
xor U71 (N_71,In_86,In_190);
nand U72 (N_72,In_272,In_431);
or U73 (N_73,In_33,In_22);
or U74 (N_74,In_309,In_101);
and U75 (N_75,In_437,In_276);
nand U76 (N_76,In_350,In_317);
nand U77 (N_77,In_198,In_117);
and U78 (N_78,In_274,In_141);
or U79 (N_79,In_223,In_113);
nand U80 (N_80,In_372,In_177);
xnor U81 (N_81,In_165,In_181);
nand U82 (N_82,In_420,In_43);
and U83 (N_83,In_24,In_284);
nand U84 (N_84,In_342,In_404);
and U85 (N_85,In_20,In_218);
nor U86 (N_86,In_385,In_128);
nor U87 (N_87,In_251,In_456);
or U88 (N_88,In_161,In_136);
nand U89 (N_89,In_406,In_137);
and U90 (N_90,In_415,In_39);
or U91 (N_91,In_447,In_90);
nand U92 (N_92,In_71,In_175);
nor U93 (N_93,In_189,In_54);
xor U94 (N_94,In_454,In_30);
nor U95 (N_95,In_330,In_464);
nor U96 (N_96,In_219,In_460);
or U97 (N_97,In_333,In_25);
nor U98 (N_98,In_303,In_77);
or U99 (N_99,In_495,In_277);
nor U100 (N_100,In_241,In_32);
xnor U101 (N_101,In_97,In_405);
and U102 (N_102,N_43,In_427);
nor U103 (N_103,In_15,In_73);
or U104 (N_104,N_70,In_208);
xnor U105 (N_105,In_386,N_94);
nor U106 (N_106,In_209,N_38);
nand U107 (N_107,In_215,N_8);
nor U108 (N_108,In_485,In_89);
or U109 (N_109,In_5,In_448);
and U110 (N_110,In_336,N_21);
nor U111 (N_111,N_55,In_217);
or U112 (N_112,N_44,In_481);
nand U113 (N_113,In_92,In_196);
or U114 (N_114,In_270,In_192);
nand U115 (N_115,N_4,N_62);
or U116 (N_116,In_238,In_61);
and U117 (N_117,N_17,In_400);
nand U118 (N_118,In_311,In_133);
or U119 (N_119,N_29,N_25);
and U120 (N_120,In_152,In_353);
nand U121 (N_121,In_359,N_28);
or U122 (N_122,In_484,In_360);
and U123 (N_123,In_193,In_185);
xnor U124 (N_124,In_9,In_279);
nand U125 (N_125,In_95,In_70);
or U126 (N_126,In_414,N_13);
or U127 (N_127,In_329,N_97);
or U128 (N_128,In_328,In_139);
nor U129 (N_129,In_312,N_87);
or U130 (N_130,In_444,In_357);
nand U131 (N_131,In_224,In_180);
and U132 (N_132,N_6,In_291);
or U133 (N_133,In_258,In_387);
and U134 (N_134,In_234,In_493);
or U135 (N_135,In_252,In_442);
nand U136 (N_136,N_47,In_201);
and U137 (N_137,N_65,N_23);
nand U138 (N_138,In_327,In_487);
xnor U139 (N_139,N_91,N_49);
nand U140 (N_140,N_54,In_413);
and U141 (N_141,N_40,In_494);
and U142 (N_142,In_428,N_63);
and U143 (N_143,In_167,N_51);
nor U144 (N_144,N_20,In_320);
and U145 (N_145,In_438,In_367);
or U146 (N_146,N_2,N_9);
nand U147 (N_147,N_96,In_41);
and U148 (N_148,In_179,In_488);
nand U149 (N_149,In_307,In_271);
nand U150 (N_150,In_93,In_216);
nor U151 (N_151,In_197,In_394);
nor U152 (N_152,In_103,N_37);
nor U153 (N_153,In_403,In_262);
and U154 (N_154,In_109,In_361);
and U155 (N_155,N_36,In_3);
and U156 (N_156,In_74,N_27);
and U157 (N_157,In_294,In_389);
or U158 (N_158,In_55,In_45);
and U159 (N_159,N_15,N_98);
xnor U160 (N_160,In_491,N_30);
or U161 (N_161,In_156,In_370);
nor U162 (N_162,In_98,In_373);
and U163 (N_163,In_59,In_314);
and U164 (N_164,In_126,In_378);
or U165 (N_165,In_380,In_402);
nor U166 (N_166,In_349,In_158);
and U167 (N_167,N_67,In_476);
xor U168 (N_168,In_207,N_58);
nand U169 (N_169,In_302,In_259);
or U170 (N_170,In_75,N_85);
nor U171 (N_171,In_323,In_283);
or U172 (N_172,In_51,In_419);
nor U173 (N_173,In_8,In_472);
nor U174 (N_174,In_85,In_375);
or U175 (N_175,In_35,In_401);
or U176 (N_176,In_423,In_16);
or U177 (N_177,In_115,In_163);
and U178 (N_178,In_72,In_347);
or U179 (N_179,N_48,In_301);
or U180 (N_180,In_204,N_33);
and U181 (N_181,In_441,In_188);
or U182 (N_182,In_263,In_151);
or U183 (N_183,N_79,In_246);
nor U184 (N_184,In_475,In_56);
and U185 (N_185,In_169,In_395);
xnor U186 (N_186,In_281,N_3);
or U187 (N_187,In_67,In_267);
and U188 (N_188,In_369,In_325);
nor U189 (N_189,N_78,In_492);
xor U190 (N_190,In_348,In_408);
nand U191 (N_191,N_82,In_289);
nand U192 (N_192,In_148,N_39);
or U193 (N_193,In_340,In_280);
xnor U194 (N_194,In_463,In_129);
and U195 (N_195,In_305,In_122);
and U196 (N_196,N_64,N_61);
nand U197 (N_197,In_31,N_32);
nand U198 (N_198,In_21,In_453);
and U199 (N_199,N_74,N_0);
xnor U200 (N_200,In_471,N_162);
nand U201 (N_201,In_58,In_81);
and U202 (N_202,N_167,N_72);
and U203 (N_203,N_141,In_362);
or U204 (N_204,N_199,In_298);
nor U205 (N_205,N_175,N_195);
nand U206 (N_206,In_290,N_42);
nand U207 (N_207,N_84,N_182);
xor U208 (N_208,In_296,N_147);
and U209 (N_209,In_499,N_7);
or U210 (N_210,In_354,N_186);
nor U211 (N_211,N_134,N_77);
or U212 (N_212,N_180,N_69);
or U213 (N_213,N_148,N_104);
nand U214 (N_214,In_345,In_489);
or U215 (N_215,In_490,N_129);
nand U216 (N_216,N_150,N_133);
xor U217 (N_217,In_199,N_169);
nor U218 (N_218,N_165,N_115);
xnor U219 (N_219,In_486,In_461);
and U220 (N_220,In_266,In_310);
nor U221 (N_221,In_100,N_109);
or U222 (N_222,N_31,In_346);
nand U223 (N_223,N_89,In_212);
and U224 (N_224,In_430,In_409);
nor U225 (N_225,N_88,N_45);
nor U226 (N_226,N_102,N_111);
nor U227 (N_227,In_288,In_172);
nand U228 (N_228,N_163,N_132);
nand U229 (N_229,In_478,N_80);
and U230 (N_230,In_220,In_200);
nor U231 (N_231,N_114,N_196);
nand U232 (N_232,In_239,In_116);
nand U233 (N_233,In_455,In_482);
xnor U234 (N_234,N_118,N_90);
and U235 (N_235,N_185,In_392);
xor U236 (N_236,In_278,N_24);
xnor U237 (N_237,N_197,N_139);
nor U238 (N_238,N_81,N_190);
nor U239 (N_239,In_374,N_93);
and U240 (N_240,In_435,N_140);
or U241 (N_241,N_105,N_142);
nor U242 (N_242,N_179,In_446);
nand U243 (N_243,N_50,N_173);
nand U244 (N_244,N_146,N_18);
or U245 (N_245,N_131,In_142);
nand U246 (N_246,N_124,In_68);
xnor U247 (N_247,In_326,N_177);
nor U248 (N_248,In_17,N_71);
nand U249 (N_249,In_443,In_106);
or U250 (N_250,In_383,In_371);
and U251 (N_251,N_16,In_213);
and U252 (N_252,N_192,N_128);
nand U253 (N_253,In_147,N_144);
and U254 (N_254,N_123,N_34);
xnor U255 (N_255,N_171,In_91);
nand U256 (N_256,In_28,In_250);
or U257 (N_257,N_157,In_18);
or U258 (N_258,N_95,In_292);
nor U259 (N_259,In_364,N_76);
or U260 (N_260,N_189,N_125);
or U261 (N_261,N_100,In_469);
or U262 (N_262,In_36,In_66);
and U263 (N_263,N_66,In_445);
and U264 (N_264,N_174,In_449);
nand U265 (N_265,N_35,In_286);
nand U266 (N_266,In_332,In_210);
nor U267 (N_267,N_137,In_242);
or U268 (N_268,N_75,N_92);
nand U269 (N_269,In_94,N_41);
nand U270 (N_270,N_164,N_172);
or U271 (N_271,In_293,N_11);
nor U272 (N_272,In_131,In_127);
and U273 (N_273,In_82,In_497);
and U274 (N_274,In_221,In_417);
or U275 (N_275,In_143,In_318);
nor U276 (N_276,N_110,N_181);
or U277 (N_277,N_46,In_237);
or U278 (N_278,In_225,N_143);
or U279 (N_279,In_432,In_249);
nand U280 (N_280,In_164,In_229);
and U281 (N_281,N_112,N_56);
xor U282 (N_282,N_176,In_480);
nand U283 (N_283,N_168,In_319);
nor U284 (N_284,In_34,In_76);
or U285 (N_285,In_334,In_397);
or U286 (N_286,N_127,N_119);
xor U287 (N_287,N_198,In_140);
or U288 (N_288,N_22,N_86);
or U289 (N_289,N_53,N_26);
xnor U290 (N_290,N_191,N_10);
or U291 (N_291,N_73,In_411);
xor U292 (N_292,In_135,N_160);
xnor U293 (N_293,In_230,N_152);
and U294 (N_294,In_382,N_154);
and U295 (N_295,In_468,In_355);
nor U296 (N_296,In_29,N_68);
or U297 (N_297,In_341,N_193);
nand U298 (N_298,In_191,In_146);
nand U299 (N_299,N_194,N_178);
nor U300 (N_300,N_282,In_64);
or U301 (N_301,N_269,N_138);
or U302 (N_302,In_243,N_289);
and U303 (N_303,In_295,N_188);
nand U304 (N_304,N_290,N_271);
nor U305 (N_305,N_113,N_258);
or U306 (N_306,In_393,In_233);
or U307 (N_307,N_206,In_424);
nand U308 (N_308,N_299,N_210);
nand U309 (N_309,N_153,N_52);
xor U310 (N_310,N_101,N_57);
and U311 (N_311,In_60,In_433);
nor U312 (N_312,N_232,In_343);
or U313 (N_313,N_106,N_201);
or U314 (N_314,In_351,N_270);
nor U315 (N_315,N_227,N_107);
or U316 (N_316,In_388,N_103);
or U317 (N_317,In_458,N_155);
nor U318 (N_318,N_219,N_246);
and U319 (N_319,N_247,N_267);
and U320 (N_320,N_291,In_155);
nand U321 (N_321,N_208,In_247);
nand U322 (N_322,N_243,N_216);
nor U323 (N_323,In_157,In_222);
or U324 (N_324,N_242,N_263);
nand U325 (N_325,N_233,N_244);
nor U326 (N_326,In_339,N_248);
nor U327 (N_327,N_108,N_159);
nand U328 (N_328,N_83,In_299);
and U329 (N_329,N_220,N_231);
nand U330 (N_330,N_293,N_122);
and U331 (N_331,In_465,N_251);
nand U332 (N_332,N_126,N_136);
or U333 (N_333,N_240,N_184);
nor U334 (N_334,In_253,In_421);
or U335 (N_335,N_296,In_231);
nor U336 (N_336,N_203,N_215);
xor U337 (N_337,N_295,In_40);
or U338 (N_338,In_254,N_207);
nand U339 (N_339,N_14,N_260);
or U340 (N_340,N_214,N_217);
and U341 (N_341,In_244,In_248);
nor U342 (N_342,N_170,N_273);
nor U343 (N_343,N_60,N_235);
nand U344 (N_344,In_37,In_232);
and U345 (N_345,N_264,N_19);
nand U346 (N_346,In_79,N_211);
and U347 (N_347,In_344,N_151);
or U348 (N_348,N_116,N_283);
or U349 (N_349,N_259,N_280);
or U350 (N_350,N_225,N_249);
xnor U351 (N_351,In_124,In_285);
and U352 (N_352,N_236,N_297);
and U353 (N_353,In_195,In_105);
nor U354 (N_354,N_121,In_150);
nand U355 (N_355,N_202,In_477);
or U356 (N_356,N_223,N_166);
or U357 (N_357,In_466,In_170);
nor U358 (N_358,N_237,N_218);
nor U359 (N_359,N_298,N_245);
or U360 (N_360,In_416,In_236);
or U361 (N_361,N_239,N_222);
nand U362 (N_362,N_204,N_209);
or U363 (N_363,In_19,N_149);
nor U364 (N_364,N_205,In_62);
and U365 (N_365,N_268,N_254);
nor U366 (N_366,In_166,In_52);
xnor U367 (N_367,N_12,N_130);
or U368 (N_368,N_213,N_120);
nor U369 (N_369,N_277,N_284);
nand U370 (N_370,N_288,N_221);
or U371 (N_371,N_145,N_279);
or U372 (N_372,N_156,In_227);
or U373 (N_373,N_135,In_2);
nor U374 (N_374,N_238,In_174);
and U375 (N_375,N_183,N_161);
nor U376 (N_376,N_286,In_1);
or U377 (N_377,N_257,N_276);
or U378 (N_378,N_274,N_275);
and U379 (N_379,N_253,N_228);
nor U380 (N_380,N_187,N_250);
nand U381 (N_381,N_200,In_228);
or U382 (N_382,N_117,N_287);
nand U383 (N_383,N_241,N_252);
and U384 (N_384,N_5,In_27);
nor U385 (N_385,N_294,N_285);
nand U386 (N_386,In_240,N_234);
and U387 (N_387,N_265,N_255);
nand U388 (N_388,N_229,N_99);
nand U389 (N_389,N_256,N_281);
nand U390 (N_390,N_230,In_398);
nor U391 (N_391,N_272,N_158);
nor U392 (N_392,In_160,In_211);
xor U393 (N_393,N_292,In_474);
or U394 (N_394,In_23,N_278);
nand U395 (N_395,N_212,N_261);
or U396 (N_396,N_262,In_260);
or U397 (N_397,In_138,N_59);
nand U398 (N_398,N_1,N_226);
nand U399 (N_399,N_224,N_266);
and U400 (N_400,N_330,N_331);
and U401 (N_401,N_391,N_350);
and U402 (N_402,N_385,N_346);
or U403 (N_403,N_363,N_351);
xor U404 (N_404,N_392,N_327);
nand U405 (N_405,N_301,N_347);
or U406 (N_406,N_316,N_397);
or U407 (N_407,N_336,N_318);
or U408 (N_408,N_380,N_382);
nor U409 (N_409,N_390,N_375);
nor U410 (N_410,N_379,N_357);
or U411 (N_411,N_342,N_307);
nor U412 (N_412,N_388,N_344);
nor U413 (N_413,N_353,N_369);
or U414 (N_414,N_358,N_377);
and U415 (N_415,N_335,N_300);
nand U416 (N_416,N_322,N_368);
nand U417 (N_417,N_343,N_303);
nor U418 (N_418,N_309,N_332);
and U419 (N_419,N_315,N_314);
nor U420 (N_420,N_366,N_365);
or U421 (N_421,N_381,N_361);
nor U422 (N_422,N_319,N_374);
and U423 (N_423,N_389,N_339);
and U424 (N_424,N_313,N_340);
or U425 (N_425,N_304,N_383);
or U426 (N_426,N_338,N_348);
and U427 (N_427,N_396,N_352);
or U428 (N_428,N_371,N_398);
or U429 (N_429,N_394,N_384);
and U430 (N_430,N_372,N_367);
nand U431 (N_431,N_329,N_364);
and U432 (N_432,N_326,N_334);
and U433 (N_433,N_317,N_386);
xor U434 (N_434,N_349,N_305);
or U435 (N_435,N_312,N_328);
xnor U436 (N_436,N_378,N_359);
nor U437 (N_437,N_355,N_376);
nor U438 (N_438,N_323,N_399);
and U439 (N_439,N_360,N_362);
and U440 (N_440,N_320,N_373);
nand U441 (N_441,N_354,N_395);
or U442 (N_442,N_325,N_310);
or U443 (N_443,N_302,N_337);
or U444 (N_444,N_370,N_311);
nor U445 (N_445,N_345,N_324);
and U446 (N_446,N_308,N_321);
or U447 (N_447,N_356,N_341);
nor U448 (N_448,N_333,N_306);
nand U449 (N_449,N_387,N_393);
nand U450 (N_450,N_370,N_307);
nor U451 (N_451,N_317,N_309);
xor U452 (N_452,N_361,N_319);
nand U453 (N_453,N_316,N_377);
nor U454 (N_454,N_306,N_398);
nor U455 (N_455,N_396,N_334);
nor U456 (N_456,N_357,N_358);
and U457 (N_457,N_310,N_301);
and U458 (N_458,N_351,N_394);
or U459 (N_459,N_323,N_356);
or U460 (N_460,N_382,N_322);
xnor U461 (N_461,N_371,N_344);
nor U462 (N_462,N_356,N_375);
nor U463 (N_463,N_380,N_386);
or U464 (N_464,N_340,N_382);
nand U465 (N_465,N_340,N_301);
or U466 (N_466,N_300,N_333);
and U467 (N_467,N_317,N_320);
and U468 (N_468,N_309,N_308);
nor U469 (N_469,N_331,N_321);
nand U470 (N_470,N_350,N_361);
or U471 (N_471,N_362,N_303);
nand U472 (N_472,N_388,N_316);
and U473 (N_473,N_324,N_366);
or U474 (N_474,N_372,N_368);
and U475 (N_475,N_368,N_330);
xnor U476 (N_476,N_382,N_318);
nand U477 (N_477,N_377,N_343);
xnor U478 (N_478,N_328,N_376);
or U479 (N_479,N_353,N_376);
or U480 (N_480,N_348,N_345);
and U481 (N_481,N_344,N_305);
and U482 (N_482,N_364,N_365);
xnor U483 (N_483,N_333,N_366);
and U484 (N_484,N_348,N_325);
nand U485 (N_485,N_351,N_350);
xnor U486 (N_486,N_316,N_380);
and U487 (N_487,N_382,N_367);
nand U488 (N_488,N_354,N_346);
and U489 (N_489,N_319,N_316);
or U490 (N_490,N_305,N_390);
nand U491 (N_491,N_341,N_339);
xnor U492 (N_492,N_314,N_364);
and U493 (N_493,N_361,N_383);
or U494 (N_494,N_330,N_303);
and U495 (N_495,N_399,N_351);
or U496 (N_496,N_332,N_346);
nand U497 (N_497,N_311,N_333);
xnor U498 (N_498,N_318,N_364);
nand U499 (N_499,N_306,N_396);
xor U500 (N_500,N_438,N_444);
xnor U501 (N_501,N_405,N_447);
nand U502 (N_502,N_476,N_489);
and U503 (N_503,N_474,N_425);
or U504 (N_504,N_414,N_436);
nor U505 (N_505,N_432,N_471);
nand U506 (N_506,N_406,N_411);
nor U507 (N_507,N_428,N_434);
nor U508 (N_508,N_452,N_490);
nor U509 (N_509,N_404,N_400);
nand U510 (N_510,N_496,N_492);
nand U511 (N_511,N_479,N_494);
or U512 (N_512,N_424,N_426);
or U513 (N_513,N_421,N_487);
or U514 (N_514,N_430,N_413);
nor U515 (N_515,N_480,N_412);
nor U516 (N_516,N_429,N_491);
or U517 (N_517,N_486,N_483);
nor U518 (N_518,N_427,N_488);
or U519 (N_519,N_437,N_420);
and U520 (N_520,N_475,N_467);
or U521 (N_521,N_466,N_457);
and U522 (N_522,N_461,N_469);
nor U523 (N_523,N_449,N_454);
nor U524 (N_524,N_478,N_495);
or U525 (N_525,N_451,N_497);
nor U526 (N_526,N_456,N_407);
xor U527 (N_527,N_446,N_417);
and U528 (N_528,N_443,N_473);
or U529 (N_529,N_419,N_482);
xor U530 (N_530,N_477,N_439);
nand U531 (N_531,N_498,N_463);
nand U532 (N_532,N_415,N_455);
and U533 (N_533,N_462,N_435);
nand U534 (N_534,N_465,N_458);
or U535 (N_535,N_464,N_440);
nor U536 (N_536,N_410,N_470);
nand U537 (N_537,N_433,N_418);
nand U538 (N_538,N_453,N_403);
nand U539 (N_539,N_459,N_485);
or U540 (N_540,N_450,N_481);
and U541 (N_541,N_445,N_468);
xnor U542 (N_542,N_409,N_442);
nand U543 (N_543,N_499,N_448);
nor U544 (N_544,N_460,N_401);
nor U545 (N_545,N_493,N_484);
xnor U546 (N_546,N_402,N_431);
or U547 (N_547,N_441,N_422);
nor U548 (N_548,N_472,N_416);
xnor U549 (N_549,N_408,N_423);
nor U550 (N_550,N_458,N_496);
and U551 (N_551,N_400,N_491);
nor U552 (N_552,N_484,N_499);
nor U553 (N_553,N_467,N_474);
or U554 (N_554,N_485,N_496);
or U555 (N_555,N_469,N_414);
xnor U556 (N_556,N_426,N_499);
nand U557 (N_557,N_443,N_417);
nor U558 (N_558,N_481,N_439);
or U559 (N_559,N_411,N_457);
or U560 (N_560,N_484,N_415);
and U561 (N_561,N_441,N_438);
nor U562 (N_562,N_483,N_401);
or U563 (N_563,N_463,N_429);
nand U564 (N_564,N_407,N_427);
or U565 (N_565,N_482,N_469);
or U566 (N_566,N_489,N_413);
and U567 (N_567,N_496,N_493);
or U568 (N_568,N_484,N_409);
xnor U569 (N_569,N_438,N_464);
or U570 (N_570,N_416,N_468);
and U571 (N_571,N_434,N_457);
xor U572 (N_572,N_458,N_409);
and U573 (N_573,N_420,N_405);
nor U574 (N_574,N_409,N_493);
nand U575 (N_575,N_443,N_493);
nand U576 (N_576,N_431,N_467);
nor U577 (N_577,N_403,N_444);
and U578 (N_578,N_411,N_473);
or U579 (N_579,N_400,N_477);
nor U580 (N_580,N_437,N_466);
xor U581 (N_581,N_437,N_409);
or U582 (N_582,N_464,N_470);
or U583 (N_583,N_467,N_449);
nor U584 (N_584,N_430,N_418);
and U585 (N_585,N_463,N_488);
or U586 (N_586,N_466,N_423);
or U587 (N_587,N_451,N_426);
or U588 (N_588,N_458,N_470);
nor U589 (N_589,N_474,N_487);
nor U590 (N_590,N_450,N_412);
nand U591 (N_591,N_480,N_402);
and U592 (N_592,N_487,N_429);
xnor U593 (N_593,N_428,N_414);
nand U594 (N_594,N_478,N_426);
xor U595 (N_595,N_450,N_453);
or U596 (N_596,N_474,N_416);
nor U597 (N_597,N_470,N_491);
nor U598 (N_598,N_422,N_485);
and U599 (N_599,N_431,N_424);
and U600 (N_600,N_545,N_587);
and U601 (N_601,N_556,N_516);
nor U602 (N_602,N_533,N_550);
xnor U603 (N_603,N_517,N_562);
or U604 (N_604,N_553,N_567);
or U605 (N_605,N_544,N_530);
or U606 (N_606,N_529,N_570);
xnor U607 (N_607,N_590,N_543);
or U608 (N_608,N_572,N_501);
nand U609 (N_609,N_561,N_571);
or U610 (N_610,N_568,N_591);
and U611 (N_611,N_594,N_549);
nand U612 (N_612,N_514,N_521);
nor U613 (N_613,N_575,N_548);
nor U614 (N_614,N_551,N_523);
and U615 (N_615,N_500,N_505);
nand U616 (N_616,N_558,N_532);
xnor U617 (N_617,N_597,N_522);
nor U618 (N_618,N_566,N_564);
and U619 (N_619,N_569,N_541);
and U620 (N_620,N_579,N_588);
nor U621 (N_621,N_503,N_582);
or U622 (N_622,N_598,N_504);
nand U623 (N_623,N_518,N_547);
nor U624 (N_624,N_512,N_507);
and U625 (N_625,N_509,N_560);
or U626 (N_626,N_515,N_525);
and U627 (N_627,N_513,N_520);
or U628 (N_628,N_535,N_534);
and U629 (N_629,N_559,N_526);
and U630 (N_630,N_593,N_581);
xor U631 (N_631,N_542,N_540);
and U632 (N_632,N_538,N_555);
or U633 (N_633,N_577,N_578);
and U634 (N_634,N_574,N_565);
nand U635 (N_635,N_537,N_592);
nor U636 (N_636,N_552,N_599);
or U637 (N_637,N_528,N_508);
nor U638 (N_638,N_596,N_502);
nor U639 (N_639,N_506,N_573);
nand U640 (N_640,N_586,N_519);
nand U641 (N_641,N_511,N_527);
nand U642 (N_642,N_583,N_531);
and U643 (N_643,N_539,N_589);
nor U644 (N_644,N_585,N_536);
and U645 (N_645,N_524,N_576);
xnor U646 (N_646,N_510,N_546);
and U647 (N_647,N_580,N_563);
nand U648 (N_648,N_595,N_557);
nand U649 (N_649,N_554,N_584);
or U650 (N_650,N_519,N_594);
nor U651 (N_651,N_522,N_554);
and U652 (N_652,N_544,N_521);
or U653 (N_653,N_523,N_526);
or U654 (N_654,N_559,N_548);
nand U655 (N_655,N_587,N_559);
or U656 (N_656,N_521,N_567);
nand U657 (N_657,N_593,N_537);
and U658 (N_658,N_563,N_502);
and U659 (N_659,N_530,N_508);
nand U660 (N_660,N_558,N_587);
or U661 (N_661,N_527,N_565);
or U662 (N_662,N_575,N_537);
xor U663 (N_663,N_537,N_578);
or U664 (N_664,N_528,N_543);
nand U665 (N_665,N_505,N_544);
or U666 (N_666,N_596,N_551);
or U667 (N_667,N_541,N_585);
and U668 (N_668,N_598,N_573);
and U669 (N_669,N_506,N_541);
nand U670 (N_670,N_585,N_563);
and U671 (N_671,N_557,N_571);
or U672 (N_672,N_573,N_500);
and U673 (N_673,N_577,N_506);
nand U674 (N_674,N_561,N_581);
nand U675 (N_675,N_573,N_508);
or U676 (N_676,N_558,N_599);
and U677 (N_677,N_538,N_565);
nand U678 (N_678,N_565,N_505);
xnor U679 (N_679,N_558,N_526);
and U680 (N_680,N_583,N_569);
or U681 (N_681,N_549,N_548);
xor U682 (N_682,N_585,N_566);
nor U683 (N_683,N_510,N_570);
or U684 (N_684,N_507,N_588);
or U685 (N_685,N_529,N_544);
and U686 (N_686,N_561,N_559);
xnor U687 (N_687,N_558,N_513);
nand U688 (N_688,N_566,N_593);
nor U689 (N_689,N_553,N_509);
or U690 (N_690,N_585,N_531);
nor U691 (N_691,N_531,N_517);
nor U692 (N_692,N_507,N_599);
nor U693 (N_693,N_588,N_517);
nand U694 (N_694,N_545,N_532);
nand U695 (N_695,N_518,N_517);
and U696 (N_696,N_568,N_506);
nand U697 (N_697,N_593,N_524);
or U698 (N_698,N_541,N_505);
and U699 (N_699,N_529,N_597);
or U700 (N_700,N_649,N_641);
or U701 (N_701,N_655,N_615);
nand U702 (N_702,N_671,N_636);
and U703 (N_703,N_681,N_622);
nor U704 (N_704,N_674,N_642);
and U705 (N_705,N_666,N_623);
xor U706 (N_706,N_617,N_635);
nor U707 (N_707,N_687,N_698);
nand U708 (N_708,N_624,N_695);
and U709 (N_709,N_611,N_632);
or U710 (N_710,N_601,N_618);
and U711 (N_711,N_663,N_659);
nand U712 (N_712,N_697,N_640);
nand U713 (N_713,N_696,N_684);
or U714 (N_714,N_683,N_680);
nor U715 (N_715,N_682,N_677);
nand U716 (N_716,N_612,N_604);
nor U717 (N_717,N_639,N_690);
nor U718 (N_718,N_646,N_627);
and U719 (N_719,N_619,N_629);
or U720 (N_720,N_699,N_654);
or U721 (N_721,N_633,N_678);
xnor U722 (N_722,N_614,N_667);
nor U723 (N_723,N_691,N_673);
xnor U724 (N_724,N_656,N_648);
nand U725 (N_725,N_665,N_658);
xor U726 (N_726,N_603,N_650);
or U727 (N_727,N_607,N_685);
nand U728 (N_728,N_651,N_672);
or U729 (N_729,N_662,N_676);
nand U730 (N_730,N_688,N_621);
or U731 (N_731,N_609,N_652);
xor U732 (N_732,N_616,N_644);
and U733 (N_733,N_686,N_608);
nor U734 (N_734,N_679,N_653);
or U735 (N_735,N_605,N_613);
or U736 (N_736,N_628,N_606);
or U737 (N_737,N_694,N_630);
or U738 (N_738,N_670,N_626);
nand U739 (N_739,N_600,N_668);
nand U740 (N_740,N_692,N_647);
or U741 (N_741,N_675,N_664);
nand U742 (N_742,N_689,N_669);
and U743 (N_743,N_660,N_643);
nor U744 (N_744,N_693,N_625);
nand U745 (N_745,N_610,N_620);
and U746 (N_746,N_645,N_602);
nor U747 (N_747,N_657,N_634);
nand U748 (N_748,N_631,N_637);
nor U749 (N_749,N_661,N_638);
nand U750 (N_750,N_631,N_644);
or U751 (N_751,N_621,N_626);
nor U752 (N_752,N_666,N_630);
nor U753 (N_753,N_613,N_661);
nor U754 (N_754,N_688,N_616);
and U755 (N_755,N_690,N_643);
or U756 (N_756,N_657,N_682);
nor U757 (N_757,N_680,N_605);
nor U758 (N_758,N_685,N_645);
and U759 (N_759,N_642,N_600);
nand U760 (N_760,N_627,N_600);
nor U761 (N_761,N_614,N_699);
nor U762 (N_762,N_656,N_668);
nand U763 (N_763,N_610,N_684);
or U764 (N_764,N_634,N_669);
or U765 (N_765,N_668,N_643);
nand U766 (N_766,N_617,N_669);
and U767 (N_767,N_629,N_680);
or U768 (N_768,N_619,N_687);
nor U769 (N_769,N_653,N_684);
and U770 (N_770,N_680,N_685);
and U771 (N_771,N_639,N_698);
or U772 (N_772,N_654,N_697);
nand U773 (N_773,N_691,N_643);
and U774 (N_774,N_663,N_623);
nand U775 (N_775,N_679,N_681);
xor U776 (N_776,N_644,N_655);
and U777 (N_777,N_663,N_692);
xor U778 (N_778,N_640,N_620);
and U779 (N_779,N_607,N_614);
or U780 (N_780,N_698,N_611);
or U781 (N_781,N_608,N_615);
nor U782 (N_782,N_650,N_653);
or U783 (N_783,N_612,N_645);
and U784 (N_784,N_669,N_623);
xnor U785 (N_785,N_622,N_687);
nand U786 (N_786,N_609,N_624);
nand U787 (N_787,N_683,N_616);
nand U788 (N_788,N_671,N_681);
nor U789 (N_789,N_640,N_669);
and U790 (N_790,N_611,N_676);
nor U791 (N_791,N_610,N_674);
nor U792 (N_792,N_639,N_655);
nand U793 (N_793,N_629,N_666);
xor U794 (N_794,N_643,N_695);
and U795 (N_795,N_629,N_602);
and U796 (N_796,N_668,N_638);
xor U797 (N_797,N_600,N_651);
or U798 (N_798,N_642,N_673);
or U799 (N_799,N_608,N_609);
nor U800 (N_800,N_749,N_740);
nor U801 (N_801,N_782,N_775);
xor U802 (N_802,N_752,N_767);
nor U803 (N_803,N_738,N_712);
or U804 (N_804,N_714,N_706);
and U805 (N_805,N_783,N_765);
and U806 (N_806,N_725,N_764);
and U807 (N_807,N_736,N_745);
xor U808 (N_808,N_760,N_734);
and U809 (N_809,N_797,N_791);
or U810 (N_810,N_708,N_756);
and U811 (N_811,N_792,N_777);
or U812 (N_812,N_796,N_728);
nor U813 (N_813,N_746,N_747);
nor U814 (N_814,N_784,N_781);
or U815 (N_815,N_750,N_700);
or U816 (N_816,N_757,N_729);
and U817 (N_817,N_785,N_754);
and U818 (N_818,N_771,N_769);
nor U819 (N_819,N_705,N_742);
and U820 (N_820,N_787,N_715);
and U821 (N_821,N_768,N_762);
nor U822 (N_822,N_798,N_743);
or U823 (N_823,N_727,N_763);
nand U824 (N_824,N_794,N_718);
and U825 (N_825,N_730,N_713);
nor U826 (N_826,N_720,N_773);
xor U827 (N_827,N_751,N_793);
and U828 (N_828,N_733,N_724);
xnor U829 (N_829,N_723,N_790);
xor U830 (N_830,N_772,N_799);
or U831 (N_831,N_755,N_789);
nor U832 (N_832,N_721,N_719);
nor U833 (N_833,N_701,N_759);
and U834 (N_834,N_748,N_702);
nor U835 (N_835,N_776,N_741);
nor U836 (N_836,N_795,N_779);
or U837 (N_837,N_780,N_703);
and U838 (N_838,N_709,N_722);
and U839 (N_839,N_726,N_778);
and U840 (N_840,N_739,N_788);
or U841 (N_841,N_744,N_707);
or U842 (N_842,N_735,N_731);
nor U843 (N_843,N_766,N_711);
xnor U844 (N_844,N_732,N_716);
nand U845 (N_845,N_774,N_710);
and U846 (N_846,N_717,N_758);
and U847 (N_847,N_704,N_761);
or U848 (N_848,N_770,N_786);
and U849 (N_849,N_753,N_737);
or U850 (N_850,N_780,N_744);
nand U851 (N_851,N_750,N_762);
or U852 (N_852,N_789,N_704);
and U853 (N_853,N_782,N_721);
nor U854 (N_854,N_796,N_744);
and U855 (N_855,N_763,N_722);
xor U856 (N_856,N_760,N_722);
and U857 (N_857,N_748,N_762);
xnor U858 (N_858,N_742,N_743);
nand U859 (N_859,N_732,N_779);
xnor U860 (N_860,N_758,N_730);
or U861 (N_861,N_753,N_748);
or U862 (N_862,N_767,N_756);
nor U863 (N_863,N_792,N_704);
nor U864 (N_864,N_759,N_788);
and U865 (N_865,N_744,N_799);
nor U866 (N_866,N_770,N_765);
and U867 (N_867,N_753,N_789);
and U868 (N_868,N_793,N_735);
or U869 (N_869,N_758,N_788);
or U870 (N_870,N_782,N_739);
and U871 (N_871,N_703,N_790);
nand U872 (N_872,N_732,N_776);
and U873 (N_873,N_713,N_756);
and U874 (N_874,N_714,N_792);
nor U875 (N_875,N_758,N_706);
nand U876 (N_876,N_752,N_769);
or U877 (N_877,N_792,N_711);
and U878 (N_878,N_795,N_742);
or U879 (N_879,N_776,N_737);
nand U880 (N_880,N_735,N_752);
nand U881 (N_881,N_766,N_771);
nor U882 (N_882,N_779,N_770);
and U883 (N_883,N_774,N_760);
nand U884 (N_884,N_714,N_736);
nor U885 (N_885,N_744,N_728);
and U886 (N_886,N_725,N_799);
and U887 (N_887,N_721,N_767);
nor U888 (N_888,N_707,N_773);
and U889 (N_889,N_761,N_791);
nand U890 (N_890,N_736,N_732);
nor U891 (N_891,N_783,N_727);
nor U892 (N_892,N_766,N_705);
or U893 (N_893,N_784,N_764);
nor U894 (N_894,N_760,N_756);
and U895 (N_895,N_731,N_780);
nor U896 (N_896,N_767,N_711);
nor U897 (N_897,N_742,N_736);
nor U898 (N_898,N_797,N_752);
nand U899 (N_899,N_772,N_769);
and U900 (N_900,N_845,N_895);
xnor U901 (N_901,N_896,N_877);
nor U902 (N_902,N_890,N_851);
and U903 (N_903,N_818,N_844);
nand U904 (N_904,N_857,N_843);
or U905 (N_905,N_865,N_828);
nand U906 (N_906,N_855,N_882);
or U907 (N_907,N_880,N_802);
nor U908 (N_908,N_801,N_864);
or U909 (N_909,N_872,N_878);
nor U910 (N_910,N_846,N_825);
nor U911 (N_911,N_835,N_824);
nand U912 (N_912,N_817,N_815);
or U913 (N_913,N_837,N_812);
and U914 (N_914,N_805,N_819);
or U915 (N_915,N_831,N_868);
or U916 (N_916,N_850,N_849);
or U917 (N_917,N_899,N_842);
nand U918 (N_918,N_883,N_826);
xor U919 (N_919,N_807,N_879);
nand U920 (N_920,N_810,N_803);
and U921 (N_921,N_873,N_884);
and U922 (N_922,N_833,N_813);
and U923 (N_923,N_876,N_829);
nor U924 (N_924,N_869,N_897);
nor U925 (N_925,N_852,N_893);
xnor U926 (N_926,N_839,N_838);
nand U927 (N_927,N_811,N_894);
or U928 (N_928,N_809,N_804);
nand U929 (N_929,N_858,N_863);
or U930 (N_930,N_885,N_822);
and U931 (N_931,N_841,N_871);
nor U932 (N_932,N_832,N_830);
xnor U933 (N_933,N_862,N_816);
or U934 (N_934,N_836,N_867);
nand U935 (N_935,N_840,N_821);
xor U936 (N_936,N_875,N_861);
xnor U937 (N_937,N_892,N_823);
nand U938 (N_938,N_834,N_808);
xor U939 (N_939,N_859,N_856);
nor U940 (N_940,N_886,N_853);
or U941 (N_941,N_874,N_891);
nand U942 (N_942,N_854,N_848);
and U943 (N_943,N_889,N_881);
nor U944 (N_944,N_860,N_814);
or U945 (N_945,N_827,N_800);
xor U946 (N_946,N_887,N_866);
xor U947 (N_947,N_820,N_888);
nand U948 (N_948,N_870,N_847);
nor U949 (N_949,N_806,N_898);
xnor U950 (N_950,N_813,N_892);
and U951 (N_951,N_891,N_882);
xnor U952 (N_952,N_890,N_842);
xnor U953 (N_953,N_867,N_839);
or U954 (N_954,N_802,N_877);
nand U955 (N_955,N_892,N_822);
and U956 (N_956,N_878,N_805);
nand U957 (N_957,N_830,N_825);
and U958 (N_958,N_805,N_843);
or U959 (N_959,N_867,N_821);
nor U960 (N_960,N_890,N_803);
or U961 (N_961,N_864,N_820);
xor U962 (N_962,N_826,N_802);
xnor U963 (N_963,N_833,N_845);
xnor U964 (N_964,N_887,N_858);
nand U965 (N_965,N_883,N_820);
nor U966 (N_966,N_887,N_870);
nand U967 (N_967,N_810,N_873);
and U968 (N_968,N_875,N_816);
nor U969 (N_969,N_859,N_869);
nor U970 (N_970,N_899,N_812);
or U971 (N_971,N_825,N_878);
nand U972 (N_972,N_808,N_821);
nand U973 (N_973,N_802,N_806);
nand U974 (N_974,N_893,N_837);
nand U975 (N_975,N_837,N_874);
xnor U976 (N_976,N_899,N_890);
or U977 (N_977,N_835,N_846);
and U978 (N_978,N_800,N_821);
nand U979 (N_979,N_816,N_865);
xor U980 (N_980,N_852,N_855);
or U981 (N_981,N_878,N_851);
nor U982 (N_982,N_816,N_896);
and U983 (N_983,N_801,N_846);
or U984 (N_984,N_862,N_878);
nand U985 (N_985,N_882,N_811);
or U986 (N_986,N_801,N_869);
or U987 (N_987,N_851,N_885);
xnor U988 (N_988,N_889,N_869);
nor U989 (N_989,N_886,N_831);
xnor U990 (N_990,N_878,N_852);
nand U991 (N_991,N_859,N_871);
nor U992 (N_992,N_893,N_827);
nor U993 (N_993,N_817,N_853);
and U994 (N_994,N_898,N_895);
nor U995 (N_995,N_810,N_893);
and U996 (N_996,N_891,N_842);
nand U997 (N_997,N_848,N_805);
nand U998 (N_998,N_878,N_879);
nor U999 (N_999,N_825,N_856);
nor U1000 (N_1000,N_907,N_971);
nand U1001 (N_1001,N_954,N_969);
nand U1002 (N_1002,N_953,N_920);
or U1003 (N_1003,N_956,N_946);
nand U1004 (N_1004,N_977,N_911);
and U1005 (N_1005,N_993,N_925);
and U1006 (N_1006,N_904,N_912);
and U1007 (N_1007,N_976,N_927);
or U1008 (N_1008,N_959,N_950);
nand U1009 (N_1009,N_937,N_957);
nand U1010 (N_1010,N_929,N_948);
and U1011 (N_1011,N_924,N_960);
nor U1012 (N_1012,N_932,N_915);
nor U1013 (N_1013,N_900,N_952);
nand U1014 (N_1014,N_982,N_903);
nor U1015 (N_1015,N_909,N_930);
nand U1016 (N_1016,N_970,N_905);
or U1017 (N_1017,N_998,N_964);
nor U1018 (N_1018,N_974,N_926);
nor U1019 (N_1019,N_917,N_918);
nand U1020 (N_1020,N_928,N_906);
and U1021 (N_1021,N_963,N_978);
nand U1022 (N_1022,N_989,N_979);
xnor U1023 (N_1023,N_987,N_988);
nor U1024 (N_1024,N_943,N_902);
xor U1025 (N_1025,N_945,N_973);
or U1026 (N_1026,N_922,N_958);
nand U1027 (N_1027,N_992,N_949);
nor U1028 (N_1028,N_955,N_939);
nand U1029 (N_1029,N_935,N_962);
and U1030 (N_1030,N_994,N_916);
nand U1031 (N_1031,N_901,N_990);
or U1032 (N_1032,N_910,N_981);
or U1033 (N_1033,N_986,N_951);
nor U1034 (N_1034,N_947,N_985);
or U1035 (N_1035,N_999,N_934);
nor U1036 (N_1036,N_936,N_967);
and U1037 (N_1037,N_944,N_914);
nor U1038 (N_1038,N_908,N_938);
nand U1039 (N_1039,N_995,N_966);
and U1040 (N_1040,N_941,N_931);
and U1041 (N_1041,N_975,N_997);
xnor U1042 (N_1042,N_983,N_961);
and U1043 (N_1043,N_940,N_913);
nor U1044 (N_1044,N_984,N_942);
or U1045 (N_1045,N_923,N_921);
and U1046 (N_1046,N_965,N_996);
nand U1047 (N_1047,N_972,N_919);
or U1048 (N_1048,N_933,N_991);
or U1049 (N_1049,N_968,N_980);
nand U1050 (N_1050,N_997,N_920);
nor U1051 (N_1051,N_945,N_980);
xor U1052 (N_1052,N_943,N_926);
and U1053 (N_1053,N_953,N_956);
and U1054 (N_1054,N_902,N_993);
or U1055 (N_1055,N_940,N_999);
and U1056 (N_1056,N_932,N_930);
and U1057 (N_1057,N_981,N_982);
and U1058 (N_1058,N_909,N_998);
nand U1059 (N_1059,N_987,N_991);
or U1060 (N_1060,N_913,N_984);
nand U1061 (N_1061,N_953,N_937);
nor U1062 (N_1062,N_961,N_977);
or U1063 (N_1063,N_900,N_958);
or U1064 (N_1064,N_986,N_957);
and U1065 (N_1065,N_933,N_907);
or U1066 (N_1066,N_969,N_904);
nor U1067 (N_1067,N_903,N_940);
nor U1068 (N_1068,N_916,N_964);
and U1069 (N_1069,N_921,N_994);
nor U1070 (N_1070,N_995,N_999);
nand U1071 (N_1071,N_936,N_912);
nor U1072 (N_1072,N_929,N_956);
and U1073 (N_1073,N_918,N_990);
and U1074 (N_1074,N_927,N_951);
nor U1075 (N_1075,N_978,N_920);
nor U1076 (N_1076,N_914,N_948);
or U1077 (N_1077,N_971,N_950);
or U1078 (N_1078,N_965,N_913);
or U1079 (N_1079,N_921,N_943);
nor U1080 (N_1080,N_941,N_993);
and U1081 (N_1081,N_917,N_902);
or U1082 (N_1082,N_957,N_929);
or U1083 (N_1083,N_905,N_978);
nand U1084 (N_1084,N_927,N_943);
nor U1085 (N_1085,N_917,N_995);
and U1086 (N_1086,N_986,N_963);
and U1087 (N_1087,N_913,N_900);
and U1088 (N_1088,N_977,N_983);
nand U1089 (N_1089,N_953,N_924);
and U1090 (N_1090,N_968,N_976);
nor U1091 (N_1091,N_930,N_943);
nor U1092 (N_1092,N_945,N_911);
nor U1093 (N_1093,N_976,N_995);
nand U1094 (N_1094,N_968,N_995);
and U1095 (N_1095,N_947,N_945);
and U1096 (N_1096,N_905,N_997);
nor U1097 (N_1097,N_950,N_964);
nand U1098 (N_1098,N_990,N_932);
and U1099 (N_1099,N_973,N_954);
nor U1100 (N_1100,N_1051,N_1070);
and U1101 (N_1101,N_1072,N_1035);
nand U1102 (N_1102,N_1001,N_1005);
nor U1103 (N_1103,N_1015,N_1002);
nand U1104 (N_1104,N_1099,N_1043);
xnor U1105 (N_1105,N_1026,N_1094);
and U1106 (N_1106,N_1088,N_1027);
nand U1107 (N_1107,N_1092,N_1062);
or U1108 (N_1108,N_1042,N_1041);
and U1109 (N_1109,N_1007,N_1003);
xor U1110 (N_1110,N_1021,N_1038);
nand U1111 (N_1111,N_1048,N_1011);
and U1112 (N_1112,N_1082,N_1028);
xnor U1113 (N_1113,N_1080,N_1052);
and U1114 (N_1114,N_1057,N_1079);
nand U1115 (N_1115,N_1034,N_1000);
nand U1116 (N_1116,N_1061,N_1085);
nand U1117 (N_1117,N_1020,N_1014);
and U1118 (N_1118,N_1076,N_1066);
nand U1119 (N_1119,N_1025,N_1090);
nor U1120 (N_1120,N_1036,N_1059);
nor U1121 (N_1121,N_1084,N_1029);
nand U1122 (N_1122,N_1047,N_1095);
or U1123 (N_1123,N_1096,N_1008);
nor U1124 (N_1124,N_1068,N_1018);
nor U1125 (N_1125,N_1055,N_1097);
or U1126 (N_1126,N_1056,N_1049);
nor U1127 (N_1127,N_1089,N_1016);
and U1128 (N_1128,N_1053,N_1069);
nand U1129 (N_1129,N_1044,N_1045);
and U1130 (N_1130,N_1067,N_1037);
nand U1131 (N_1131,N_1083,N_1054);
xor U1132 (N_1132,N_1031,N_1050);
or U1133 (N_1133,N_1073,N_1032);
nand U1134 (N_1134,N_1023,N_1017);
nor U1135 (N_1135,N_1087,N_1030);
nand U1136 (N_1136,N_1040,N_1091);
and U1137 (N_1137,N_1098,N_1064);
nand U1138 (N_1138,N_1033,N_1013);
xnor U1139 (N_1139,N_1077,N_1046);
nand U1140 (N_1140,N_1022,N_1006);
nand U1141 (N_1141,N_1065,N_1004);
and U1142 (N_1142,N_1081,N_1060);
nor U1143 (N_1143,N_1074,N_1039);
nor U1144 (N_1144,N_1058,N_1078);
nand U1145 (N_1145,N_1086,N_1009);
nand U1146 (N_1146,N_1063,N_1075);
or U1147 (N_1147,N_1019,N_1012);
and U1148 (N_1148,N_1093,N_1071);
nand U1149 (N_1149,N_1024,N_1010);
or U1150 (N_1150,N_1052,N_1065);
or U1151 (N_1151,N_1089,N_1067);
or U1152 (N_1152,N_1053,N_1004);
xor U1153 (N_1153,N_1015,N_1063);
nor U1154 (N_1154,N_1096,N_1001);
and U1155 (N_1155,N_1075,N_1053);
nor U1156 (N_1156,N_1010,N_1071);
and U1157 (N_1157,N_1012,N_1074);
and U1158 (N_1158,N_1019,N_1077);
xor U1159 (N_1159,N_1093,N_1055);
nand U1160 (N_1160,N_1029,N_1066);
and U1161 (N_1161,N_1058,N_1017);
nand U1162 (N_1162,N_1086,N_1061);
and U1163 (N_1163,N_1076,N_1014);
and U1164 (N_1164,N_1069,N_1041);
and U1165 (N_1165,N_1094,N_1080);
xor U1166 (N_1166,N_1050,N_1037);
and U1167 (N_1167,N_1073,N_1071);
or U1168 (N_1168,N_1017,N_1084);
nor U1169 (N_1169,N_1031,N_1081);
or U1170 (N_1170,N_1088,N_1013);
nor U1171 (N_1171,N_1001,N_1012);
nor U1172 (N_1172,N_1015,N_1018);
nor U1173 (N_1173,N_1049,N_1059);
or U1174 (N_1174,N_1099,N_1044);
or U1175 (N_1175,N_1028,N_1025);
nor U1176 (N_1176,N_1055,N_1068);
nand U1177 (N_1177,N_1090,N_1022);
and U1178 (N_1178,N_1067,N_1056);
and U1179 (N_1179,N_1065,N_1094);
nor U1180 (N_1180,N_1021,N_1005);
nand U1181 (N_1181,N_1067,N_1015);
or U1182 (N_1182,N_1067,N_1052);
and U1183 (N_1183,N_1093,N_1066);
xor U1184 (N_1184,N_1029,N_1032);
and U1185 (N_1185,N_1019,N_1070);
or U1186 (N_1186,N_1073,N_1022);
nor U1187 (N_1187,N_1064,N_1006);
nor U1188 (N_1188,N_1098,N_1028);
xnor U1189 (N_1189,N_1067,N_1016);
or U1190 (N_1190,N_1084,N_1085);
or U1191 (N_1191,N_1022,N_1071);
nand U1192 (N_1192,N_1087,N_1097);
and U1193 (N_1193,N_1001,N_1062);
or U1194 (N_1194,N_1037,N_1035);
nor U1195 (N_1195,N_1079,N_1033);
nor U1196 (N_1196,N_1083,N_1020);
and U1197 (N_1197,N_1092,N_1060);
nand U1198 (N_1198,N_1081,N_1091);
nand U1199 (N_1199,N_1025,N_1088);
and U1200 (N_1200,N_1153,N_1197);
xor U1201 (N_1201,N_1152,N_1130);
and U1202 (N_1202,N_1134,N_1127);
or U1203 (N_1203,N_1131,N_1188);
or U1204 (N_1204,N_1124,N_1119);
xor U1205 (N_1205,N_1113,N_1145);
xnor U1206 (N_1206,N_1191,N_1129);
and U1207 (N_1207,N_1176,N_1112);
nor U1208 (N_1208,N_1158,N_1163);
nand U1209 (N_1209,N_1147,N_1143);
nor U1210 (N_1210,N_1198,N_1116);
nand U1211 (N_1211,N_1120,N_1137);
nand U1212 (N_1212,N_1182,N_1135);
nand U1213 (N_1213,N_1150,N_1104);
nor U1214 (N_1214,N_1110,N_1155);
or U1215 (N_1215,N_1169,N_1146);
or U1216 (N_1216,N_1105,N_1107);
and U1217 (N_1217,N_1175,N_1173);
and U1218 (N_1218,N_1194,N_1149);
nand U1219 (N_1219,N_1195,N_1156);
nor U1220 (N_1220,N_1144,N_1189);
or U1221 (N_1221,N_1177,N_1114);
xnor U1222 (N_1222,N_1159,N_1133);
and U1223 (N_1223,N_1164,N_1170);
or U1224 (N_1224,N_1103,N_1115);
or U1225 (N_1225,N_1192,N_1122);
or U1226 (N_1226,N_1117,N_1108);
or U1227 (N_1227,N_1126,N_1100);
or U1228 (N_1228,N_1154,N_1157);
nand U1229 (N_1229,N_1180,N_1162);
nand U1230 (N_1230,N_1179,N_1125);
or U1231 (N_1231,N_1165,N_1166);
and U1232 (N_1232,N_1139,N_1102);
and U1233 (N_1233,N_1184,N_1196);
or U1234 (N_1234,N_1181,N_1140);
nand U1235 (N_1235,N_1199,N_1141);
nand U1236 (N_1236,N_1148,N_1178);
and U1237 (N_1237,N_1128,N_1151);
or U1238 (N_1238,N_1167,N_1121);
nor U1239 (N_1239,N_1138,N_1193);
or U1240 (N_1240,N_1136,N_1186);
and U1241 (N_1241,N_1160,N_1174);
or U1242 (N_1242,N_1161,N_1168);
or U1243 (N_1243,N_1132,N_1106);
or U1244 (N_1244,N_1109,N_1187);
or U1245 (N_1245,N_1118,N_1190);
or U1246 (N_1246,N_1123,N_1171);
and U1247 (N_1247,N_1185,N_1142);
nand U1248 (N_1248,N_1111,N_1101);
and U1249 (N_1249,N_1183,N_1172);
nand U1250 (N_1250,N_1196,N_1178);
and U1251 (N_1251,N_1142,N_1151);
nand U1252 (N_1252,N_1116,N_1138);
nand U1253 (N_1253,N_1175,N_1152);
nand U1254 (N_1254,N_1141,N_1155);
nor U1255 (N_1255,N_1146,N_1148);
and U1256 (N_1256,N_1191,N_1146);
xor U1257 (N_1257,N_1180,N_1186);
or U1258 (N_1258,N_1169,N_1174);
and U1259 (N_1259,N_1142,N_1141);
and U1260 (N_1260,N_1118,N_1110);
nor U1261 (N_1261,N_1187,N_1151);
nor U1262 (N_1262,N_1109,N_1148);
or U1263 (N_1263,N_1159,N_1135);
and U1264 (N_1264,N_1109,N_1136);
or U1265 (N_1265,N_1174,N_1102);
nor U1266 (N_1266,N_1176,N_1157);
and U1267 (N_1267,N_1103,N_1186);
nor U1268 (N_1268,N_1129,N_1110);
nand U1269 (N_1269,N_1168,N_1129);
nand U1270 (N_1270,N_1107,N_1122);
nor U1271 (N_1271,N_1155,N_1179);
or U1272 (N_1272,N_1136,N_1175);
nand U1273 (N_1273,N_1187,N_1179);
and U1274 (N_1274,N_1149,N_1161);
nand U1275 (N_1275,N_1172,N_1142);
nand U1276 (N_1276,N_1186,N_1140);
xor U1277 (N_1277,N_1169,N_1102);
nand U1278 (N_1278,N_1168,N_1130);
and U1279 (N_1279,N_1161,N_1180);
or U1280 (N_1280,N_1149,N_1120);
nor U1281 (N_1281,N_1183,N_1105);
nand U1282 (N_1282,N_1117,N_1199);
and U1283 (N_1283,N_1186,N_1143);
nand U1284 (N_1284,N_1187,N_1123);
and U1285 (N_1285,N_1138,N_1165);
nor U1286 (N_1286,N_1159,N_1139);
nand U1287 (N_1287,N_1173,N_1168);
nor U1288 (N_1288,N_1164,N_1175);
and U1289 (N_1289,N_1122,N_1118);
nor U1290 (N_1290,N_1114,N_1198);
nor U1291 (N_1291,N_1127,N_1137);
nand U1292 (N_1292,N_1199,N_1107);
or U1293 (N_1293,N_1144,N_1129);
nand U1294 (N_1294,N_1190,N_1149);
nand U1295 (N_1295,N_1113,N_1137);
and U1296 (N_1296,N_1101,N_1195);
and U1297 (N_1297,N_1192,N_1196);
nor U1298 (N_1298,N_1197,N_1109);
or U1299 (N_1299,N_1160,N_1183);
nand U1300 (N_1300,N_1248,N_1258);
nor U1301 (N_1301,N_1260,N_1211);
and U1302 (N_1302,N_1271,N_1202);
nand U1303 (N_1303,N_1231,N_1250);
nor U1304 (N_1304,N_1272,N_1278);
and U1305 (N_1305,N_1216,N_1294);
or U1306 (N_1306,N_1263,N_1277);
nand U1307 (N_1307,N_1295,N_1241);
or U1308 (N_1308,N_1243,N_1230);
nor U1309 (N_1309,N_1268,N_1283);
nand U1310 (N_1310,N_1238,N_1235);
nand U1311 (N_1311,N_1289,N_1214);
nand U1312 (N_1312,N_1215,N_1297);
and U1313 (N_1313,N_1265,N_1286);
or U1314 (N_1314,N_1227,N_1267);
xor U1315 (N_1315,N_1254,N_1229);
and U1316 (N_1316,N_1249,N_1274);
or U1317 (N_1317,N_1221,N_1270);
xnor U1318 (N_1318,N_1222,N_1220);
and U1319 (N_1319,N_1223,N_1240);
nor U1320 (N_1320,N_1237,N_1273);
nand U1321 (N_1321,N_1233,N_1252);
xor U1322 (N_1322,N_1208,N_1280);
nand U1323 (N_1323,N_1219,N_1262);
or U1324 (N_1324,N_1224,N_1225);
and U1325 (N_1325,N_1200,N_1204);
or U1326 (N_1326,N_1244,N_1247);
or U1327 (N_1327,N_1293,N_1291);
xor U1328 (N_1328,N_1251,N_1264);
or U1329 (N_1329,N_1209,N_1239);
nand U1330 (N_1330,N_1218,N_1207);
nor U1331 (N_1331,N_1269,N_1228);
nor U1332 (N_1332,N_1255,N_1256);
nor U1333 (N_1333,N_1210,N_1201);
nor U1334 (N_1334,N_1246,N_1282);
nor U1335 (N_1335,N_1290,N_1203);
and U1336 (N_1336,N_1234,N_1279);
nand U1337 (N_1337,N_1298,N_1212);
or U1338 (N_1338,N_1281,N_1266);
and U1339 (N_1339,N_1261,N_1276);
and U1340 (N_1340,N_1284,N_1206);
and U1341 (N_1341,N_1232,N_1205);
nor U1342 (N_1342,N_1245,N_1299);
nor U1343 (N_1343,N_1288,N_1296);
nor U1344 (N_1344,N_1292,N_1253);
nor U1345 (N_1345,N_1236,N_1259);
and U1346 (N_1346,N_1275,N_1285);
nor U1347 (N_1347,N_1226,N_1217);
nand U1348 (N_1348,N_1213,N_1287);
or U1349 (N_1349,N_1242,N_1257);
nor U1350 (N_1350,N_1216,N_1246);
and U1351 (N_1351,N_1267,N_1244);
or U1352 (N_1352,N_1231,N_1221);
nor U1353 (N_1353,N_1255,N_1276);
or U1354 (N_1354,N_1299,N_1274);
xnor U1355 (N_1355,N_1237,N_1248);
and U1356 (N_1356,N_1262,N_1258);
and U1357 (N_1357,N_1253,N_1282);
nand U1358 (N_1358,N_1222,N_1268);
nand U1359 (N_1359,N_1284,N_1209);
nand U1360 (N_1360,N_1238,N_1265);
nand U1361 (N_1361,N_1284,N_1226);
and U1362 (N_1362,N_1283,N_1260);
and U1363 (N_1363,N_1250,N_1247);
and U1364 (N_1364,N_1223,N_1280);
or U1365 (N_1365,N_1254,N_1246);
nor U1366 (N_1366,N_1206,N_1247);
nand U1367 (N_1367,N_1296,N_1291);
nor U1368 (N_1368,N_1269,N_1291);
nand U1369 (N_1369,N_1254,N_1287);
and U1370 (N_1370,N_1204,N_1263);
or U1371 (N_1371,N_1285,N_1234);
xnor U1372 (N_1372,N_1263,N_1268);
or U1373 (N_1373,N_1297,N_1246);
or U1374 (N_1374,N_1206,N_1235);
and U1375 (N_1375,N_1213,N_1226);
or U1376 (N_1376,N_1247,N_1259);
or U1377 (N_1377,N_1258,N_1228);
xnor U1378 (N_1378,N_1255,N_1218);
nand U1379 (N_1379,N_1270,N_1247);
or U1380 (N_1380,N_1293,N_1240);
nand U1381 (N_1381,N_1279,N_1258);
nand U1382 (N_1382,N_1270,N_1239);
nand U1383 (N_1383,N_1231,N_1263);
nor U1384 (N_1384,N_1256,N_1264);
nor U1385 (N_1385,N_1257,N_1221);
and U1386 (N_1386,N_1206,N_1262);
and U1387 (N_1387,N_1227,N_1274);
and U1388 (N_1388,N_1202,N_1229);
or U1389 (N_1389,N_1218,N_1295);
and U1390 (N_1390,N_1288,N_1287);
nor U1391 (N_1391,N_1257,N_1209);
or U1392 (N_1392,N_1265,N_1272);
or U1393 (N_1393,N_1229,N_1204);
and U1394 (N_1394,N_1256,N_1298);
or U1395 (N_1395,N_1274,N_1271);
nor U1396 (N_1396,N_1285,N_1291);
nor U1397 (N_1397,N_1206,N_1278);
xnor U1398 (N_1398,N_1244,N_1219);
nor U1399 (N_1399,N_1210,N_1271);
nor U1400 (N_1400,N_1368,N_1345);
nor U1401 (N_1401,N_1381,N_1308);
nand U1402 (N_1402,N_1356,N_1319);
and U1403 (N_1403,N_1397,N_1349);
or U1404 (N_1404,N_1393,N_1377);
and U1405 (N_1405,N_1370,N_1364);
xnor U1406 (N_1406,N_1379,N_1355);
or U1407 (N_1407,N_1365,N_1310);
and U1408 (N_1408,N_1362,N_1351);
nor U1409 (N_1409,N_1309,N_1382);
nand U1410 (N_1410,N_1367,N_1300);
and U1411 (N_1411,N_1388,N_1336);
nor U1412 (N_1412,N_1389,N_1337);
nor U1413 (N_1413,N_1338,N_1305);
nor U1414 (N_1414,N_1306,N_1354);
and U1415 (N_1415,N_1311,N_1361);
and U1416 (N_1416,N_1374,N_1347);
and U1417 (N_1417,N_1399,N_1391);
xnor U1418 (N_1418,N_1334,N_1357);
nor U1419 (N_1419,N_1380,N_1318);
nand U1420 (N_1420,N_1316,N_1341);
nand U1421 (N_1421,N_1392,N_1396);
or U1422 (N_1422,N_1307,N_1394);
nand U1423 (N_1423,N_1387,N_1328);
or U1424 (N_1424,N_1378,N_1371);
nor U1425 (N_1425,N_1320,N_1329);
nand U1426 (N_1426,N_1342,N_1304);
nor U1427 (N_1427,N_1395,N_1369);
and U1428 (N_1428,N_1330,N_1385);
or U1429 (N_1429,N_1358,N_1322);
nand U1430 (N_1430,N_1398,N_1343);
and U1431 (N_1431,N_1373,N_1327);
and U1432 (N_1432,N_1323,N_1359);
nand U1433 (N_1433,N_1333,N_1372);
xor U1434 (N_1434,N_1335,N_1303);
nor U1435 (N_1435,N_1352,N_1360);
nor U1436 (N_1436,N_1344,N_1331);
nor U1437 (N_1437,N_1386,N_1302);
nor U1438 (N_1438,N_1346,N_1339);
nand U1439 (N_1439,N_1348,N_1332);
and U1440 (N_1440,N_1313,N_1376);
and U1441 (N_1441,N_1324,N_1326);
xor U1442 (N_1442,N_1312,N_1317);
nor U1443 (N_1443,N_1325,N_1353);
xnor U1444 (N_1444,N_1314,N_1375);
and U1445 (N_1445,N_1390,N_1383);
and U1446 (N_1446,N_1301,N_1340);
nand U1447 (N_1447,N_1363,N_1384);
and U1448 (N_1448,N_1366,N_1321);
nand U1449 (N_1449,N_1350,N_1315);
nor U1450 (N_1450,N_1351,N_1328);
and U1451 (N_1451,N_1389,N_1362);
and U1452 (N_1452,N_1316,N_1346);
xor U1453 (N_1453,N_1335,N_1352);
nand U1454 (N_1454,N_1321,N_1388);
nor U1455 (N_1455,N_1345,N_1329);
nand U1456 (N_1456,N_1343,N_1323);
nand U1457 (N_1457,N_1342,N_1307);
or U1458 (N_1458,N_1308,N_1302);
and U1459 (N_1459,N_1329,N_1336);
or U1460 (N_1460,N_1348,N_1328);
or U1461 (N_1461,N_1364,N_1337);
and U1462 (N_1462,N_1377,N_1300);
nand U1463 (N_1463,N_1360,N_1395);
nor U1464 (N_1464,N_1315,N_1325);
xor U1465 (N_1465,N_1344,N_1307);
nor U1466 (N_1466,N_1335,N_1379);
xnor U1467 (N_1467,N_1334,N_1332);
nand U1468 (N_1468,N_1379,N_1350);
or U1469 (N_1469,N_1320,N_1359);
xnor U1470 (N_1470,N_1324,N_1358);
or U1471 (N_1471,N_1309,N_1314);
and U1472 (N_1472,N_1382,N_1351);
or U1473 (N_1473,N_1393,N_1313);
and U1474 (N_1474,N_1386,N_1329);
nor U1475 (N_1475,N_1361,N_1392);
nor U1476 (N_1476,N_1363,N_1374);
nor U1477 (N_1477,N_1377,N_1391);
xnor U1478 (N_1478,N_1393,N_1341);
nor U1479 (N_1479,N_1361,N_1359);
nand U1480 (N_1480,N_1350,N_1383);
and U1481 (N_1481,N_1372,N_1364);
nand U1482 (N_1482,N_1327,N_1356);
nand U1483 (N_1483,N_1322,N_1344);
or U1484 (N_1484,N_1378,N_1332);
and U1485 (N_1485,N_1376,N_1321);
and U1486 (N_1486,N_1352,N_1320);
or U1487 (N_1487,N_1387,N_1317);
and U1488 (N_1488,N_1387,N_1336);
nand U1489 (N_1489,N_1338,N_1309);
xor U1490 (N_1490,N_1356,N_1387);
xnor U1491 (N_1491,N_1391,N_1316);
nand U1492 (N_1492,N_1383,N_1349);
or U1493 (N_1493,N_1307,N_1326);
or U1494 (N_1494,N_1362,N_1320);
nand U1495 (N_1495,N_1351,N_1334);
nor U1496 (N_1496,N_1346,N_1394);
nor U1497 (N_1497,N_1381,N_1361);
nor U1498 (N_1498,N_1364,N_1321);
or U1499 (N_1499,N_1343,N_1317);
nand U1500 (N_1500,N_1402,N_1465);
nor U1501 (N_1501,N_1438,N_1401);
nor U1502 (N_1502,N_1457,N_1454);
and U1503 (N_1503,N_1450,N_1452);
and U1504 (N_1504,N_1418,N_1419);
nand U1505 (N_1505,N_1445,N_1473);
xor U1506 (N_1506,N_1494,N_1469);
nand U1507 (N_1507,N_1478,N_1437);
nor U1508 (N_1508,N_1484,N_1427);
and U1509 (N_1509,N_1479,N_1458);
or U1510 (N_1510,N_1434,N_1409);
nand U1511 (N_1511,N_1470,N_1485);
and U1512 (N_1512,N_1475,N_1449);
or U1513 (N_1513,N_1423,N_1425);
or U1514 (N_1514,N_1481,N_1428);
nor U1515 (N_1515,N_1430,N_1424);
and U1516 (N_1516,N_1443,N_1406);
nor U1517 (N_1517,N_1412,N_1422);
and U1518 (N_1518,N_1456,N_1461);
and U1519 (N_1519,N_1415,N_1477);
xnor U1520 (N_1520,N_1468,N_1466);
and U1521 (N_1521,N_1487,N_1493);
nor U1522 (N_1522,N_1492,N_1490);
and U1523 (N_1523,N_1472,N_1462);
and U1524 (N_1524,N_1496,N_1421);
or U1525 (N_1525,N_1439,N_1433);
nor U1526 (N_1526,N_1414,N_1480);
and U1527 (N_1527,N_1460,N_1467);
nand U1528 (N_1528,N_1459,N_1488);
nor U1529 (N_1529,N_1455,N_1448);
and U1530 (N_1530,N_1498,N_1476);
and U1531 (N_1531,N_1429,N_1436);
nor U1532 (N_1532,N_1432,N_1497);
nor U1533 (N_1533,N_1441,N_1453);
xnor U1534 (N_1534,N_1411,N_1495);
nand U1535 (N_1535,N_1451,N_1440);
or U1536 (N_1536,N_1408,N_1463);
and U1537 (N_1537,N_1499,N_1400);
nand U1538 (N_1538,N_1447,N_1404);
xor U1539 (N_1539,N_1446,N_1489);
and U1540 (N_1540,N_1486,N_1417);
or U1541 (N_1541,N_1471,N_1407);
or U1542 (N_1542,N_1405,N_1474);
nor U1543 (N_1543,N_1482,N_1416);
nand U1544 (N_1544,N_1444,N_1431);
nor U1545 (N_1545,N_1426,N_1483);
and U1546 (N_1546,N_1491,N_1420);
nor U1547 (N_1547,N_1464,N_1413);
nor U1548 (N_1548,N_1442,N_1435);
nor U1549 (N_1549,N_1410,N_1403);
or U1550 (N_1550,N_1474,N_1458);
nand U1551 (N_1551,N_1443,N_1408);
nand U1552 (N_1552,N_1484,N_1466);
and U1553 (N_1553,N_1438,N_1419);
nand U1554 (N_1554,N_1496,N_1468);
or U1555 (N_1555,N_1450,N_1490);
nand U1556 (N_1556,N_1418,N_1401);
nor U1557 (N_1557,N_1414,N_1460);
xor U1558 (N_1558,N_1486,N_1422);
and U1559 (N_1559,N_1481,N_1455);
nand U1560 (N_1560,N_1412,N_1403);
nand U1561 (N_1561,N_1466,N_1486);
nand U1562 (N_1562,N_1487,N_1419);
nor U1563 (N_1563,N_1420,N_1400);
or U1564 (N_1564,N_1496,N_1445);
or U1565 (N_1565,N_1448,N_1441);
nor U1566 (N_1566,N_1489,N_1437);
nor U1567 (N_1567,N_1488,N_1499);
and U1568 (N_1568,N_1457,N_1405);
and U1569 (N_1569,N_1443,N_1459);
nor U1570 (N_1570,N_1408,N_1495);
nand U1571 (N_1571,N_1444,N_1483);
or U1572 (N_1572,N_1405,N_1423);
nor U1573 (N_1573,N_1454,N_1442);
nand U1574 (N_1574,N_1492,N_1458);
or U1575 (N_1575,N_1427,N_1402);
nor U1576 (N_1576,N_1446,N_1495);
and U1577 (N_1577,N_1437,N_1485);
nor U1578 (N_1578,N_1401,N_1465);
xnor U1579 (N_1579,N_1476,N_1407);
xor U1580 (N_1580,N_1446,N_1406);
nor U1581 (N_1581,N_1481,N_1435);
and U1582 (N_1582,N_1479,N_1442);
and U1583 (N_1583,N_1476,N_1483);
nand U1584 (N_1584,N_1468,N_1409);
nor U1585 (N_1585,N_1412,N_1410);
and U1586 (N_1586,N_1420,N_1434);
nor U1587 (N_1587,N_1432,N_1492);
nor U1588 (N_1588,N_1480,N_1465);
and U1589 (N_1589,N_1417,N_1460);
nand U1590 (N_1590,N_1477,N_1442);
nand U1591 (N_1591,N_1411,N_1438);
nor U1592 (N_1592,N_1494,N_1498);
nand U1593 (N_1593,N_1425,N_1475);
nor U1594 (N_1594,N_1475,N_1470);
or U1595 (N_1595,N_1460,N_1456);
nor U1596 (N_1596,N_1419,N_1425);
or U1597 (N_1597,N_1454,N_1467);
and U1598 (N_1598,N_1409,N_1496);
nand U1599 (N_1599,N_1439,N_1418);
nor U1600 (N_1600,N_1533,N_1558);
nand U1601 (N_1601,N_1524,N_1511);
or U1602 (N_1602,N_1554,N_1535);
or U1603 (N_1603,N_1517,N_1542);
nand U1604 (N_1604,N_1530,N_1564);
xnor U1605 (N_1605,N_1546,N_1581);
nor U1606 (N_1606,N_1504,N_1589);
nor U1607 (N_1607,N_1591,N_1528);
or U1608 (N_1608,N_1599,N_1527);
nand U1609 (N_1609,N_1566,N_1534);
nand U1610 (N_1610,N_1519,N_1590);
and U1611 (N_1611,N_1565,N_1521);
or U1612 (N_1612,N_1568,N_1550);
or U1613 (N_1613,N_1583,N_1540);
and U1614 (N_1614,N_1513,N_1512);
or U1615 (N_1615,N_1573,N_1575);
nor U1616 (N_1616,N_1580,N_1506);
nand U1617 (N_1617,N_1520,N_1525);
nor U1618 (N_1618,N_1538,N_1532);
or U1619 (N_1619,N_1507,N_1588);
or U1620 (N_1620,N_1503,N_1544);
xnor U1621 (N_1621,N_1505,N_1571);
nor U1622 (N_1622,N_1537,N_1570);
nor U1623 (N_1623,N_1502,N_1598);
nor U1624 (N_1624,N_1529,N_1593);
or U1625 (N_1625,N_1563,N_1594);
or U1626 (N_1626,N_1569,N_1548);
or U1627 (N_1627,N_1584,N_1510);
and U1628 (N_1628,N_1578,N_1592);
or U1629 (N_1629,N_1543,N_1560);
nor U1630 (N_1630,N_1547,N_1531);
or U1631 (N_1631,N_1576,N_1509);
xnor U1632 (N_1632,N_1508,N_1555);
and U1633 (N_1633,N_1586,N_1579);
or U1634 (N_1634,N_1541,N_1522);
xor U1635 (N_1635,N_1526,N_1557);
xor U1636 (N_1636,N_1597,N_1574);
nand U1637 (N_1637,N_1587,N_1582);
xor U1638 (N_1638,N_1552,N_1562);
or U1639 (N_1639,N_1518,N_1536);
or U1640 (N_1640,N_1553,N_1523);
nand U1641 (N_1641,N_1515,N_1516);
or U1642 (N_1642,N_1514,N_1539);
or U1643 (N_1643,N_1545,N_1585);
or U1644 (N_1644,N_1556,N_1595);
nand U1645 (N_1645,N_1500,N_1549);
nand U1646 (N_1646,N_1596,N_1551);
and U1647 (N_1647,N_1561,N_1567);
or U1648 (N_1648,N_1501,N_1559);
nor U1649 (N_1649,N_1577,N_1572);
nand U1650 (N_1650,N_1517,N_1586);
or U1651 (N_1651,N_1588,N_1565);
or U1652 (N_1652,N_1583,N_1562);
and U1653 (N_1653,N_1536,N_1573);
nand U1654 (N_1654,N_1532,N_1515);
xnor U1655 (N_1655,N_1587,N_1528);
nor U1656 (N_1656,N_1500,N_1577);
nand U1657 (N_1657,N_1525,N_1503);
and U1658 (N_1658,N_1523,N_1557);
and U1659 (N_1659,N_1508,N_1599);
or U1660 (N_1660,N_1528,N_1515);
or U1661 (N_1661,N_1552,N_1570);
or U1662 (N_1662,N_1562,N_1542);
nor U1663 (N_1663,N_1545,N_1538);
nand U1664 (N_1664,N_1516,N_1576);
and U1665 (N_1665,N_1555,N_1548);
or U1666 (N_1666,N_1528,N_1584);
or U1667 (N_1667,N_1574,N_1569);
nor U1668 (N_1668,N_1592,N_1528);
or U1669 (N_1669,N_1552,N_1540);
nand U1670 (N_1670,N_1508,N_1590);
or U1671 (N_1671,N_1507,N_1530);
or U1672 (N_1672,N_1535,N_1589);
or U1673 (N_1673,N_1536,N_1563);
nand U1674 (N_1674,N_1593,N_1568);
nor U1675 (N_1675,N_1589,N_1585);
nand U1676 (N_1676,N_1574,N_1553);
nand U1677 (N_1677,N_1542,N_1509);
nand U1678 (N_1678,N_1501,N_1512);
xor U1679 (N_1679,N_1548,N_1510);
and U1680 (N_1680,N_1501,N_1507);
nand U1681 (N_1681,N_1559,N_1591);
xnor U1682 (N_1682,N_1514,N_1530);
nor U1683 (N_1683,N_1556,N_1596);
nand U1684 (N_1684,N_1575,N_1591);
or U1685 (N_1685,N_1539,N_1552);
and U1686 (N_1686,N_1557,N_1554);
xnor U1687 (N_1687,N_1527,N_1583);
and U1688 (N_1688,N_1598,N_1561);
xor U1689 (N_1689,N_1531,N_1593);
nor U1690 (N_1690,N_1538,N_1560);
nand U1691 (N_1691,N_1531,N_1526);
nand U1692 (N_1692,N_1536,N_1531);
and U1693 (N_1693,N_1570,N_1502);
or U1694 (N_1694,N_1516,N_1526);
or U1695 (N_1695,N_1545,N_1569);
or U1696 (N_1696,N_1510,N_1597);
or U1697 (N_1697,N_1514,N_1587);
and U1698 (N_1698,N_1518,N_1579);
nor U1699 (N_1699,N_1540,N_1594);
xnor U1700 (N_1700,N_1684,N_1691);
nor U1701 (N_1701,N_1613,N_1652);
nor U1702 (N_1702,N_1675,N_1623);
or U1703 (N_1703,N_1664,N_1648);
and U1704 (N_1704,N_1660,N_1692);
nand U1705 (N_1705,N_1699,N_1602);
nand U1706 (N_1706,N_1661,N_1680);
nand U1707 (N_1707,N_1682,N_1672);
xnor U1708 (N_1708,N_1609,N_1637);
xor U1709 (N_1709,N_1697,N_1612);
and U1710 (N_1710,N_1658,N_1616);
and U1711 (N_1711,N_1641,N_1649);
and U1712 (N_1712,N_1610,N_1636);
nor U1713 (N_1713,N_1656,N_1694);
nor U1714 (N_1714,N_1624,N_1678);
or U1715 (N_1715,N_1628,N_1689);
nand U1716 (N_1716,N_1647,N_1614);
or U1717 (N_1717,N_1620,N_1631);
nand U1718 (N_1718,N_1653,N_1622);
and U1719 (N_1719,N_1695,N_1617);
nor U1720 (N_1720,N_1643,N_1674);
or U1721 (N_1721,N_1632,N_1625);
or U1722 (N_1722,N_1644,N_1685);
or U1723 (N_1723,N_1650,N_1662);
or U1724 (N_1724,N_1642,N_1626);
nor U1725 (N_1725,N_1671,N_1657);
nor U1726 (N_1726,N_1698,N_1600);
nand U1727 (N_1727,N_1619,N_1606);
or U1728 (N_1728,N_1608,N_1640);
or U1729 (N_1729,N_1654,N_1630);
nor U1730 (N_1730,N_1683,N_1611);
and U1731 (N_1731,N_1665,N_1601);
nor U1732 (N_1732,N_1655,N_1645);
nor U1733 (N_1733,N_1696,N_1635);
and U1734 (N_1734,N_1669,N_1651);
nor U1735 (N_1735,N_1634,N_1687);
and U1736 (N_1736,N_1639,N_1646);
nand U1737 (N_1737,N_1676,N_1605);
or U1738 (N_1738,N_1668,N_1686);
nand U1739 (N_1739,N_1615,N_1667);
and U1740 (N_1740,N_1638,N_1607);
nand U1741 (N_1741,N_1633,N_1688);
and U1742 (N_1742,N_1690,N_1629);
xor U1743 (N_1743,N_1666,N_1618);
nor U1744 (N_1744,N_1663,N_1673);
or U1745 (N_1745,N_1681,N_1659);
or U1746 (N_1746,N_1693,N_1603);
and U1747 (N_1747,N_1621,N_1677);
xor U1748 (N_1748,N_1670,N_1604);
nand U1749 (N_1749,N_1679,N_1627);
and U1750 (N_1750,N_1636,N_1639);
xor U1751 (N_1751,N_1681,N_1622);
or U1752 (N_1752,N_1636,N_1663);
nand U1753 (N_1753,N_1698,N_1614);
nor U1754 (N_1754,N_1692,N_1623);
nand U1755 (N_1755,N_1646,N_1688);
or U1756 (N_1756,N_1668,N_1631);
nor U1757 (N_1757,N_1684,N_1666);
nor U1758 (N_1758,N_1649,N_1676);
xor U1759 (N_1759,N_1687,N_1667);
nand U1760 (N_1760,N_1687,N_1675);
or U1761 (N_1761,N_1687,N_1673);
nor U1762 (N_1762,N_1640,N_1650);
xnor U1763 (N_1763,N_1641,N_1664);
or U1764 (N_1764,N_1641,N_1608);
and U1765 (N_1765,N_1637,N_1658);
or U1766 (N_1766,N_1600,N_1623);
nor U1767 (N_1767,N_1666,N_1693);
and U1768 (N_1768,N_1614,N_1684);
or U1769 (N_1769,N_1651,N_1646);
nand U1770 (N_1770,N_1619,N_1669);
nand U1771 (N_1771,N_1671,N_1665);
nand U1772 (N_1772,N_1660,N_1687);
and U1773 (N_1773,N_1626,N_1601);
nand U1774 (N_1774,N_1695,N_1658);
nand U1775 (N_1775,N_1607,N_1692);
and U1776 (N_1776,N_1621,N_1657);
and U1777 (N_1777,N_1682,N_1638);
and U1778 (N_1778,N_1688,N_1630);
nand U1779 (N_1779,N_1648,N_1691);
and U1780 (N_1780,N_1671,N_1684);
or U1781 (N_1781,N_1694,N_1692);
or U1782 (N_1782,N_1637,N_1675);
and U1783 (N_1783,N_1697,N_1601);
xor U1784 (N_1784,N_1696,N_1627);
or U1785 (N_1785,N_1684,N_1697);
nand U1786 (N_1786,N_1623,N_1689);
nor U1787 (N_1787,N_1693,N_1602);
xnor U1788 (N_1788,N_1615,N_1668);
nand U1789 (N_1789,N_1648,N_1614);
nand U1790 (N_1790,N_1609,N_1679);
or U1791 (N_1791,N_1648,N_1656);
and U1792 (N_1792,N_1682,N_1697);
xnor U1793 (N_1793,N_1660,N_1614);
nor U1794 (N_1794,N_1607,N_1646);
and U1795 (N_1795,N_1688,N_1658);
or U1796 (N_1796,N_1692,N_1614);
nand U1797 (N_1797,N_1635,N_1647);
nand U1798 (N_1798,N_1664,N_1643);
or U1799 (N_1799,N_1678,N_1689);
nand U1800 (N_1800,N_1790,N_1701);
nand U1801 (N_1801,N_1733,N_1795);
and U1802 (N_1802,N_1777,N_1751);
nand U1803 (N_1803,N_1798,N_1793);
and U1804 (N_1804,N_1796,N_1719);
xnor U1805 (N_1805,N_1782,N_1784);
nor U1806 (N_1806,N_1762,N_1773);
or U1807 (N_1807,N_1730,N_1759);
or U1808 (N_1808,N_1703,N_1723);
or U1809 (N_1809,N_1738,N_1713);
and U1810 (N_1810,N_1729,N_1712);
xor U1811 (N_1811,N_1724,N_1768);
nor U1812 (N_1812,N_1743,N_1722);
and U1813 (N_1813,N_1706,N_1714);
or U1814 (N_1814,N_1732,N_1772);
nor U1815 (N_1815,N_1755,N_1774);
nor U1816 (N_1816,N_1744,N_1700);
and U1817 (N_1817,N_1702,N_1710);
xor U1818 (N_1818,N_1717,N_1767);
and U1819 (N_1819,N_1731,N_1704);
nor U1820 (N_1820,N_1766,N_1791);
and U1821 (N_1821,N_1742,N_1776);
nand U1822 (N_1822,N_1705,N_1780);
nand U1823 (N_1823,N_1725,N_1747);
nand U1824 (N_1824,N_1760,N_1736);
or U1825 (N_1825,N_1771,N_1765);
nor U1826 (N_1826,N_1779,N_1745);
nor U1827 (N_1827,N_1770,N_1789);
or U1828 (N_1828,N_1769,N_1721);
or U1829 (N_1829,N_1781,N_1709);
nor U1830 (N_1830,N_1788,N_1707);
nor U1831 (N_1831,N_1734,N_1740);
nand U1832 (N_1832,N_1764,N_1757);
nor U1833 (N_1833,N_1786,N_1756);
and U1834 (N_1834,N_1754,N_1720);
nor U1835 (N_1835,N_1708,N_1727);
nand U1836 (N_1836,N_1728,N_1792);
nor U1837 (N_1837,N_1799,N_1746);
and U1838 (N_1838,N_1763,N_1750);
or U1839 (N_1839,N_1752,N_1715);
nand U1840 (N_1840,N_1783,N_1785);
or U1841 (N_1841,N_1718,N_1726);
and U1842 (N_1842,N_1797,N_1758);
or U1843 (N_1843,N_1741,N_1761);
nand U1844 (N_1844,N_1778,N_1748);
nand U1845 (N_1845,N_1737,N_1787);
nand U1846 (N_1846,N_1749,N_1739);
and U1847 (N_1847,N_1735,N_1794);
nor U1848 (N_1848,N_1716,N_1711);
nor U1849 (N_1849,N_1775,N_1753);
nor U1850 (N_1850,N_1781,N_1728);
xnor U1851 (N_1851,N_1719,N_1780);
nand U1852 (N_1852,N_1739,N_1770);
nand U1853 (N_1853,N_1707,N_1747);
nor U1854 (N_1854,N_1738,N_1733);
xor U1855 (N_1855,N_1785,N_1715);
and U1856 (N_1856,N_1714,N_1799);
nor U1857 (N_1857,N_1704,N_1791);
or U1858 (N_1858,N_1779,N_1717);
xor U1859 (N_1859,N_1787,N_1727);
and U1860 (N_1860,N_1701,N_1719);
and U1861 (N_1861,N_1793,N_1788);
nor U1862 (N_1862,N_1758,N_1727);
and U1863 (N_1863,N_1782,N_1773);
xnor U1864 (N_1864,N_1764,N_1751);
xor U1865 (N_1865,N_1708,N_1763);
and U1866 (N_1866,N_1761,N_1754);
xnor U1867 (N_1867,N_1752,N_1771);
and U1868 (N_1868,N_1703,N_1736);
or U1869 (N_1869,N_1715,N_1726);
nand U1870 (N_1870,N_1768,N_1719);
nand U1871 (N_1871,N_1760,N_1713);
xnor U1872 (N_1872,N_1750,N_1778);
and U1873 (N_1873,N_1709,N_1796);
xnor U1874 (N_1874,N_1757,N_1758);
nor U1875 (N_1875,N_1779,N_1768);
nand U1876 (N_1876,N_1755,N_1776);
nor U1877 (N_1877,N_1793,N_1750);
xor U1878 (N_1878,N_1794,N_1731);
and U1879 (N_1879,N_1702,N_1780);
nand U1880 (N_1880,N_1760,N_1749);
and U1881 (N_1881,N_1748,N_1796);
or U1882 (N_1882,N_1784,N_1702);
xor U1883 (N_1883,N_1749,N_1702);
nand U1884 (N_1884,N_1727,N_1746);
and U1885 (N_1885,N_1756,N_1726);
nand U1886 (N_1886,N_1763,N_1779);
or U1887 (N_1887,N_1721,N_1783);
xnor U1888 (N_1888,N_1745,N_1799);
and U1889 (N_1889,N_1712,N_1711);
nor U1890 (N_1890,N_1797,N_1763);
xnor U1891 (N_1891,N_1701,N_1752);
nand U1892 (N_1892,N_1747,N_1733);
or U1893 (N_1893,N_1771,N_1795);
nor U1894 (N_1894,N_1745,N_1758);
xor U1895 (N_1895,N_1757,N_1714);
nor U1896 (N_1896,N_1724,N_1701);
nor U1897 (N_1897,N_1760,N_1763);
nand U1898 (N_1898,N_1772,N_1739);
and U1899 (N_1899,N_1701,N_1780);
and U1900 (N_1900,N_1801,N_1836);
nand U1901 (N_1901,N_1889,N_1871);
or U1902 (N_1902,N_1845,N_1806);
nor U1903 (N_1903,N_1852,N_1892);
or U1904 (N_1904,N_1878,N_1816);
nand U1905 (N_1905,N_1858,N_1808);
nand U1906 (N_1906,N_1813,N_1809);
xnor U1907 (N_1907,N_1865,N_1869);
nor U1908 (N_1908,N_1807,N_1846);
or U1909 (N_1909,N_1803,N_1837);
xor U1910 (N_1910,N_1853,N_1859);
nor U1911 (N_1911,N_1823,N_1882);
and U1912 (N_1912,N_1811,N_1812);
nor U1913 (N_1913,N_1824,N_1840);
and U1914 (N_1914,N_1819,N_1839);
nand U1915 (N_1915,N_1874,N_1861);
xor U1916 (N_1916,N_1815,N_1832);
nand U1917 (N_1917,N_1873,N_1887);
or U1918 (N_1918,N_1821,N_1827);
or U1919 (N_1919,N_1817,N_1800);
or U1920 (N_1920,N_1885,N_1842);
and U1921 (N_1921,N_1895,N_1851);
nor U1922 (N_1922,N_1850,N_1838);
or U1923 (N_1923,N_1890,N_1894);
nor U1924 (N_1924,N_1857,N_1814);
and U1925 (N_1925,N_1841,N_1891);
or U1926 (N_1926,N_1883,N_1867);
nand U1927 (N_1927,N_1864,N_1802);
nand U1928 (N_1928,N_1893,N_1835);
or U1929 (N_1929,N_1884,N_1829);
nand U1930 (N_1930,N_1805,N_1897);
nor U1931 (N_1931,N_1828,N_1855);
or U1932 (N_1932,N_1881,N_1880);
nor U1933 (N_1933,N_1818,N_1877);
nand U1934 (N_1934,N_1804,N_1886);
or U1935 (N_1935,N_1875,N_1810);
xnor U1936 (N_1936,N_1854,N_1896);
nand U1937 (N_1937,N_1822,N_1848);
xnor U1938 (N_1938,N_1868,N_1888);
and U1939 (N_1939,N_1830,N_1866);
or U1940 (N_1940,N_1870,N_1843);
nand U1941 (N_1941,N_1856,N_1872);
or U1942 (N_1942,N_1820,N_1847);
or U1943 (N_1943,N_1849,N_1834);
or U1944 (N_1944,N_1899,N_1844);
nand U1945 (N_1945,N_1860,N_1863);
or U1946 (N_1946,N_1833,N_1876);
xor U1947 (N_1947,N_1825,N_1826);
and U1948 (N_1948,N_1831,N_1862);
and U1949 (N_1949,N_1879,N_1898);
or U1950 (N_1950,N_1841,N_1872);
and U1951 (N_1951,N_1892,N_1883);
or U1952 (N_1952,N_1873,N_1849);
nor U1953 (N_1953,N_1882,N_1839);
or U1954 (N_1954,N_1804,N_1892);
or U1955 (N_1955,N_1856,N_1865);
nand U1956 (N_1956,N_1848,N_1838);
nand U1957 (N_1957,N_1872,N_1820);
or U1958 (N_1958,N_1873,N_1855);
nand U1959 (N_1959,N_1805,N_1817);
xor U1960 (N_1960,N_1885,N_1879);
nand U1961 (N_1961,N_1876,N_1853);
nand U1962 (N_1962,N_1889,N_1846);
or U1963 (N_1963,N_1860,N_1805);
nand U1964 (N_1964,N_1854,N_1809);
nor U1965 (N_1965,N_1896,N_1899);
nor U1966 (N_1966,N_1895,N_1884);
and U1967 (N_1967,N_1800,N_1822);
and U1968 (N_1968,N_1879,N_1874);
nor U1969 (N_1969,N_1891,N_1823);
or U1970 (N_1970,N_1874,N_1859);
and U1971 (N_1971,N_1895,N_1829);
nand U1972 (N_1972,N_1849,N_1875);
and U1973 (N_1973,N_1866,N_1882);
and U1974 (N_1974,N_1875,N_1812);
nor U1975 (N_1975,N_1882,N_1855);
and U1976 (N_1976,N_1876,N_1830);
nor U1977 (N_1977,N_1810,N_1825);
nand U1978 (N_1978,N_1879,N_1820);
and U1979 (N_1979,N_1886,N_1868);
nand U1980 (N_1980,N_1804,N_1808);
or U1981 (N_1981,N_1862,N_1852);
and U1982 (N_1982,N_1846,N_1883);
nor U1983 (N_1983,N_1838,N_1858);
nor U1984 (N_1984,N_1807,N_1875);
nor U1985 (N_1985,N_1854,N_1856);
nor U1986 (N_1986,N_1805,N_1886);
or U1987 (N_1987,N_1880,N_1887);
and U1988 (N_1988,N_1808,N_1800);
nand U1989 (N_1989,N_1893,N_1827);
nor U1990 (N_1990,N_1843,N_1824);
or U1991 (N_1991,N_1872,N_1808);
xor U1992 (N_1992,N_1867,N_1850);
nand U1993 (N_1993,N_1814,N_1877);
and U1994 (N_1994,N_1847,N_1872);
or U1995 (N_1995,N_1848,N_1871);
and U1996 (N_1996,N_1821,N_1888);
nand U1997 (N_1997,N_1870,N_1876);
or U1998 (N_1998,N_1854,N_1870);
and U1999 (N_1999,N_1832,N_1826);
nor U2000 (N_2000,N_1994,N_1946);
and U2001 (N_2001,N_1930,N_1902);
nor U2002 (N_2002,N_1915,N_1922);
nor U2003 (N_2003,N_1925,N_1985);
or U2004 (N_2004,N_1980,N_1940);
xor U2005 (N_2005,N_1935,N_1957);
xnor U2006 (N_2006,N_1908,N_1991);
and U2007 (N_2007,N_1976,N_1974);
and U2008 (N_2008,N_1956,N_1927);
nand U2009 (N_2009,N_1916,N_1997);
and U2010 (N_2010,N_1942,N_1993);
nand U2011 (N_2011,N_1962,N_1917);
nor U2012 (N_2012,N_1909,N_1937);
nor U2013 (N_2013,N_1914,N_1960);
or U2014 (N_2014,N_1911,N_1972);
and U2015 (N_2015,N_1968,N_1981);
and U2016 (N_2016,N_1951,N_1919);
nor U2017 (N_2017,N_1920,N_1961);
xnor U2018 (N_2018,N_1963,N_1933);
nand U2019 (N_2019,N_1967,N_1912);
xor U2020 (N_2020,N_1947,N_1907);
and U2021 (N_2021,N_1928,N_1936);
and U2022 (N_2022,N_1979,N_1969);
nor U2023 (N_2023,N_1959,N_1924);
nand U2024 (N_2024,N_1926,N_1954);
xnor U2025 (N_2025,N_1970,N_1905);
xnor U2026 (N_2026,N_1929,N_1965);
nand U2027 (N_2027,N_1943,N_1987);
and U2028 (N_2028,N_1934,N_1918);
xnor U2029 (N_2029,N_1990,N_1932);
and U2030 (N_2030,N_1999,N_1906);
or U2031 (N_2031,N_1939,N_1913);
xnor U2032 (N_2032,N_1982,N_1955);
nand U2033 (N_2033,N_1975,N_1949);
or U2034 (N_2034,N_1971,N_1923);
xnor U2035 (N_2035,N_1921,N_1977);
nand U2036 (N_2036,N_1983,N_1941);
xnor U2037 (N_2037,N_1904,N_1978);
and U2038 (N_2038,N_1992,N_1995);
xnor U2039 (N_2039,N_1901,N_1986);
nand U2040 (N_2040,N_1958,N_1988);
nand U2041 (N_2041,N_1931,N_1952);
xor U2042 (N_2042,N_1945,N_1966);
nand U2043 (N_2043,N_1910,N_1989);
nand U2044 (N_2044,N_1964,N_1950);
and U2045 (N_2045,N_1900,N_1948);
or U2046 (N_2046,N_1998,N_1973);
nand U2047 (N_2047,N_1938,N_1944);
or U2048 (N_2048,N_1996,N_1984);
nand U2049 (N_2049,N_1903,N_1953);
nor U2050 (N_2050,N_1913,N_1906);
or U2051 (N_2051,N_1982,N_1989);
or U2052 (N_2052,N_1995,N_1974);
xor U2053 (N_2053,N_1902,N_1909);
nand U2054 (N_2054,N_1932,N_1955);
nand U2055 (N_2055,N_1913,N_1929);
or U2056 (N_2056,N_1919,N_1993);
nor U2057 (N_2057,N_1939,N_1945);
nor U2058 (N_2058,N_1947,N_1977);
or U2059 (N_2059,N_1924,N_1989);
xnor U2060 (N_2060,N_1925,N_1929);
nand U2061 (N_2061,N_1967,N_1950);
nor U2062 (N_2062,N_1936,N_1959);
and U2063 (N_2063,N_1936,N_1945);
or U2064 (N_2064,N_1926,N_1903);
and U2065 (N_2065,N_1976,N_1956);
and U2066 (N_2066,N_1984,N_1997);
or U2067 (N_2067,N_1968,N_1950);
and U2068 (N_2068,N_1918,N_1979);
and U2069 (N_2069,N_1900,N_1979);
or U2070 (N_2070,N_1987,N_1956);
nand U2071 (N_2071,N_1928,N_1905);
and U2072 (N_2072,N_1975,N_1907);
nand U2073 (N_2073,N_1963,N_1988);
and U2074 (N_2074,N_1986,N_1963);
or U2075 (N_2075,N_1916,N_1928);
nand U2076 (N_2076,N_1987,N_1920);
and U2077 (N_2077,N_1992,N_1945);
xor U2078 (N_2078,N_1974,N_1939);
xor U2079 (N_2079,N_1995,N_1924);
nor U2080 (N_2080,N_1943,N_1924);
or U2081 (N_2081,N_1913,N_1924);
nand U2082 (N_2082,N_1900,N_1984);
nor U2083 (N_2083,N_1929,N_1996);
and U2084 (N_2084,N_1938,N_1901);
or U2085 (N_2085,N_1913,N_1933);
nor U2086 (N_2086,N_1932,N_1961);
and U2087 (N_2087,N_1954,N_1977);
nand U2088 (N_2088,N_1928,N_1947);
nand U2089 (N_2089,N_1935,N_1965);
nand U2090 (N_2090,N_1953,N_1999);
nand U2091 (N_2091,N_1977,N_1915);
nor U2092 (N_2092,N_1975,N_1927);
and U2093 (N_2093,N_1933,N_1952);
nor U2094 (N_2094,N_1906,N_1970);
xnor U2095 (N_2095,N_1989,N_1993);
nor U2096 (N_2096,N_1915,N_1945);
nand U2097 (N_2097,N_1967,N_1992);
nor U2098 (N_2098,N_1994,N_1982);
or U2099 (N_2099,N_1956,N_1982);
nor U2100 (N_2100,N_2069,N_2082);
nand U2101 (N_2101,N_2059,N_2013);
and U2102 (N_2102,N_2077,N_2066);
nand U2103 (N_2103,N_2098,N_2081);
and U2104 (N_2104,N_2095,N_2027);
nand U2105 (N_2105,N_2000,N_2005);
xor U2106 (N_2106,N_2061,N_2044);
nor U2107 (N_2107,N_2017,N_2006);
xnor U2108 (N_2108,N_2091,N_2033);
nor U2109 (N_2109,N_2079,N_2052);
xnor U2110 (N_2110,N_2010,N_2080);
and U2111 (N_2111,N_2040,N_2036);
or U2112 (N_2112,N_2025,N_2031);
or U2113 (N_2113,N_2020,N_2050);
nand U2114 (N_2114,N_2014,N_2076);
and U2115 (N_2115,N_2011,N_2093);
or U2116 (N_2116,N_2028,N_2053);
or U2117 (N_2117,N_2002,N_2021);
nand U2118 (N_2118,N_2024,N_2007);
nand U2119 (N_2119,N_2001,N_2023);
nand U2120 (N_2120,N_2087,N_2008);
or U2121 (N_2121,N_2029,N_2072);
or U2122 (N_2122,N_2019,N_2042);
and U2123 (N_2123,N_2039,N_2030);
xor U2124 (N_2124,N_2012,N_2041);
or U2125 (N_2125,N_2089,N_2068);
xor U2126 (N_2126,N_2038,N_2067);
nand U2127 (N_2127,N_2074,N_2083);
xnor U2128 (N_2128,N_2064,N_2070);
nand U2129 (N_2129,N_2056,N_2003);
nand U2130 (N_2130,N_2009,N_2078);
and U2131 (N_2131,N_2022,N_2060);
or U2132 (N_2132,N_2035,N_2084);
nand U2133 (N_2133,N_2071,N_2048);
xnor U2134 (N_2134,N_2099,N_2047);
or U2135 (N_2135,N_2088,N_2073);
nand U2136 (N_2136,N_2049,N_2075);
nor U2137 (N_2137,N_2016,N_2004);
nor U2138 (N_2138,N_2051,N_2046);
nor U2139 (N_2139,N_2054,N_2043);
or U2140 (N_2140,N_2045,N_2085);
and U2141 (N_2141,N_2062,N_2032);
and U2142 (N_2142,N_2086,N_2057);
and U2143 (N_2143,N_2034,N_2065);
nor U2144 (N_2144,N_2063,N_2094);
and U2145 (N_2145,N_2055,N_2058);
or U2146 (N_2146,N_2096,N_2092);
or U2147 (N_2147,N_2026,N_2018);
nor U2148 (N_2148,N_2090,N_2015);
nor U2149 (N_2149,N_2097,N_2037);
and U2150 (N_2150,N_2045,N_2080);
nor U2151 (N_2151,N_2074,N_2093);
and U2152 (N_2152,N_2050,N_2013);
nand U2153 (N_2153,N_2024,N_2062);
nand U2154 (N_2154,N_2063,N_2019);
or U2155 (N_2155,N_2038,N_2092);
nand U2156 (N_2156,N_2042,N_2071);
nor U2157 (N_2157,N_2086,N_2005);
or U2158 (N_2158,N_2085,N_2006);
nor U2159 (N_2159,N_2005,N_2096);
and U2160 (N_2160,N_2062,N_2066);
nor U2161 (N_2161,N_2090,N_2083);
xor U2162 (N_2162,N_2078,N_2064);
nand U2163 (N_2163,N_2012,N_2028);
nor U2164 (N_2164,N_2073,N_2002);
or U2165 (N_2165,N_2064,N_2008);
nand U2166 (N_2166,N_2001,N_2094);
or U2167 (N_2167,N_2070,N_2067);
nor U2168 (N_2168,N_2099,N_2024);
xor U2169 (N_2169,N_2033,N_2098);
or U2170 (N_2170,N_2071,N_2070);
nor U2171 (N_2171,N_2042,N_2000);
nand U2172 (N_2172,N_2001,N_2044);
xor U2173 (N_2173,N_2077,N_2035);
nor U2174 (N_2174,N_2039,N_2018);
nand U2175 (N_2175,N_2006,N_2067);
or U2176 (N_2176,N_2040,N_2039);
xor U2177 (N_2177,N_2036,N_2017);
nor U2178 (N_2178,N_2034,N_2045);
nor U2179 (N_2179,N_2039,N_2035);
or U2180 (N_2180,N_2061,N_2090);
and U2181 (N_2181,N_2061,N_2074);
nand U2182 (N_2182,N_2010,N_2077);
nand U2183 (N_2183,N_2029,N_2067);
or U2184 (N_2184,N_2085,N_2099);
nor U2185 (N_2185,N_2045,N_2078);
and U2186 (N_2186,N_2066,N_2000);
nand U2187 (N_2187,N_2062,N_2018);
nor U2188 (N_2188,N_2008,N_2005);
and U2189 (N_2189,N_2041,N_2076);
nand U2190 (N_2190,N_2084,N_2018);
nor U2191 (N_2191,N_2013,N_2016);
xor U2192 (N_2192,N_2005,N_2087);
nand U2193 (N_2193,N_2043,N_2022);
nand U2194 (N_2194,N_2033,N_2079);
and U2195 (N_2195,N_2005,N_2002);
and U2196 (N_2196,N_2058,N_2037);
nand U2197 (N_2197,N_2068,N_2084);
or U2198 (N_2198,N_2009,N_2074);
and U2199 (N_2199,N_2042,N_2033);
xnor U2200 (N_2200,N_2190,N_2137);
xor U2201 (N_2201,N_2149,N_2135);
nand U2202 (N_2202,N_2133,N_2154);
nor U2203 (N_2203,N_2103,N_2102);
nor U2204 (N_2204,N_2116,N_2157);
and U2205 (N_2205,N_2125,N_2171);
nor U2206 (N_2206,N_2175,N_2170);
xor U2207 (N_2207,N_2161,N_2134);
nand U2208 (N_2208,N_2199,N_2146);
and U2209 (N_2209,N_2115,N_2136);
and U2210 (N_2210,N_2144,N_2127);
nor U2211 (N_2211,N_2112,N_2183);
and U2212 (N_2212,N_2111,N_2173);
xor U2213 (N_2213,N_2126,N_2123);
or U2214 (N_2214,N_2142,N_2174);
and U2215 (N_2215,N_2158,N_2152);
and U2216 (N_2216,N_2108,N_2121);
and U2217 (N_2217,N_2156,N_2182);
and U2218 (N_2218,N_2113,N_2155);
or U2219 (N_2219,N_2181,N_2179);
or U2220 (N_2220,N_2151,N_2110);
or U2221 (N_2221,N_2166,N_2148);
or U2222 (N_2222,N_2167,N_2191);
nor U2223 (N_2223,N_2143,N_2195);
nand U2224 (N_2224,N_2162,N_2109);
nand U2225 (N_2225,N_2131,N_2159);
nand U2226 (N_2226,N_2197,N_2153);
or U2227 (N_2227,N_2145,N_2184);
nor U2228 (N_2228,N_2105,N_2187);
nand U2229 (N_2229,N_2128,N_2130);
nor U2230 (N_2230,N_2177,N_2100);
and U2231 (N_2231,N_2192,N_2196);
nand U2232 (N_2232,N_2114,N_2180);
and U2233 (N_2233,N_2178,N_2140);
and U2234 (N_2234,N_2169,N_2106);
or U2235 (N_2235,N_2117,N_2176);
nand U2236 (N_2236,N_2107,N_2139);
xor U2237 (N_2237,N_2164,N_2104);
or U2238 (N_2238,N_2118,N_2120);
and U2239 (N_2239,N_2160,N_2172);
or U2240 (N_2240,N_2129,N_2138);
nor U2241 (N_2241,N_2132,N_2119);
or U2242 (N_2242,N_2186,N_2188);
or U2243 (N_2243,N_2101,N_2165);
nor U2244 (N_2244,N_2185,N_2141);
nor U2245 (N_2245,N_2168,N_2193);
xor U2246 (N_2246,N_2198,N_2147);
nand U2247 (N_2247,N_2189,N_2194);
and U2248 (N_2248,N_2122,N_2163);
and U2249 (N_2249,N_2150,N_2124);
nand U2250 (N_2250,N_2120,N_2160);
and U2251 (N_2251,N_2151,N_2148);
nor U2252 (N_2252,N_2168,N_2112);
nand U2253 (N_2253,N_2106,N_2150);
and U2254 (N_2254,N_2196,N_2114);
nor U2255 (N_2255,N_2103,N_2192);
nand U2256 (N_2256,N_2106,N_2187);
nand U2257 (N_2257,N_2141,N_2113);
or U2258 (N_2258,N_2171,N_2181);
xnor U2259 (N_2259,N_2166,N_2156);
or U2260 (N_2260,N_2143,N_2175);
xnor U2261 (N_2261,N_2139,N_2191);
or U2262 (N_2262,N_2131,N_2198);
and U2263 (N_2263,N_2100,N_2167);
xnor U2264 (N_2264,N_2176,N_2113);
nand U2265 (N_2265,N_2153,N_2132);
nand U2266 (N_2266,N_2167,N_2129);
or U2267 (N_2267,N_2180,N_2195);
nor U2268 (N_2268,N_2108,N_2164);
and U2269 (N_2269,N_2133,N_2198);
nor U2270 (N_2270,N_2155,N_2144);
nand U2271 (N_2271,N_2169,N_2192);
nand U2272 (N_2272,N_2147,N_2191);
or U2273 (N_2273,N_2146,N_2158);
and U2274 (N_2274,N_2151,N_2156);
nand U2275 (N_2275,N_2139,N_2103);
xor U2276 (N_2276,N_2106,N_2112);
nor U2277 (N_2277,N_2151,N_2100);
nor U2278 (N_2278,N_2128,N_2123);
nand U2279 (N_2279,N_2100,N_2125);
and U2280 (N_2280,N_2125,N_2102);
nor U2281 (N_2281,N_2180,N_2120);
nor U2282 (N_2282,N_2178,N_2106);
nand U2283 (N_2283,N_2190,N_2121);
or U2284 (N_2284,N_2116,N_2132);
nand U2285 (N_2285,N_2144,N_2125);
or U2286 (N_2286,N_2129,N_2115);
nor U2287 (N_2287,N_2123,N_2158);
nand U2288 (N_2288,N_2184,N_2169);
xor U2289 (N_2289,N_2104,N_2123);
nand U2290 (N_2290,N_2162,N_2148);
nand U2291 (N_2291,N_2138,N_2182);
nand U2292 (N_2292,N_2115,N_2132);
xor U2293 (N_2293,N_2152,N_2182);
nor U2294 (N_2294,N_2183,N_2182);
nor U2295 (N_2295,N_2125,N_2163);
nor U2296 (N_2296,N_2168,N_2116);
nor U2297 (N_2297,N_2104,N_2148);
nand U2298 (N_2298,N_2159,N_2171);
nand U2299 (N_2299,N_2123,N_2157);
nor U2300 (N_2300,N_2210,N_2260);
and U2301 (N_2301,N_2270,N_2229);
and U2302 (N_2302,N_2263,N_2253);
nor U2303 (N_2303,N_2289,N_2287);
and U2304 (N_2304,N_2291,N_2209);
and U2305 (N_2305,N_2279,N_2231);
nand U2306 (N_2306,N_2294,N_2217);
or U2307 (N_2307,N_2225,N_2295);
or U2308 (N_2308,N_2245,N_2273);
nor U2309 (N_2309,N_2283,N_2268);
nand U2310 (N_2310,N_2241,N_2286);
nor U2311 (N_2311,N_2278,N_2257);
nor U2312 (N_2312,N_2211,N_2298);
or U2313 (N_2313,N_2256,N_2297);
and U2314 (N_2314,N_2236,N_2276);
or U2315 (N_2315,N_2285,N_2200);
and U2316 (N_2316,N_2226,N_2234);
nand U2317 (N_2317,N_2237,N_2214);
nor U2318 (N_2318,N_2259,N_2204);
nor U2319 (N_2319,N_2233,N_2222);
nor U2320 (N_2320,N_2271,N_2269);
and U2321 (N_2321,N_2261,N_2235);
nor U2322 (N_2322,N_2280,N_2219);
nand U2323 (N_2323,N_2293,N_2272);
or U2324 (N_2324,N_2213,N_2274);
xnor U2325 (N_2325,N_2249,N_2258);
nor U2326 (N_2326,N_2218,N_2242);
nand U2327 (N_2327,N_2250,N_2230);
nor U2328 (N_2328,N_2299,N_2201);
xor U2329 (N_2329,N_2223,N_2252);
nand U2330 (N_2330,N_2238,N_2292);
and U2331 (N_2331,N_2207,N_2224);
or U2332 (N_2332,N_2221,N_2243);
nor U2333 (N_2333,N_2288,N_2264);
or U2334 (N_2334,N_2254,N_2262);
and U2335 (N_2335,N_2275,N_2284);
and U2336 (N_2336,N_2296,N_2228);
or U2337 (N_2337,N_2208,N_2220);
or U2338 (N_2338,N_2277,N_2203);
xnor U2339 (N_2339,N_2215,N_2246);
or U2340 (N_2340,N_2247,N_2251);
xor U2341 (N_2341,N_2232,N_2212);
nand U2342 (N_2342,N_2282,N_2202);
or U2343 (N_2343,N_2265,N_2206);
nor U2344 (N_2344,N_2244,N_2205);
nand U2345 (N_2345,N_2267,N_2281);
or U2346 (N_2346,N_2216,N_2255);
nor U2347 (N_2347,N_2248,N_2227);
and U2348 (N_2348,N_2290,N_2240);
or U2349 (N_2349,N_2239,N_2266);
nor U2350 (N_2350,N_2244,N_2291);
nor U2351 (N_2351,N_2289,N_2207);
xor U2352 (N_2352,N_2228,N_2287);
and U2353 (N_2353,N_2200,N_2216);
xor U2354 (N_2354,N_2282,N_2289);
or U2355 (N_2355,N_2278,N_2233);
or U2356 (N_2356,N_2265,N_2254);
and U2357 (N_2357,N_2278,N_2270);
or U2358 (N_2358,N_2226,N_2247);
or U2359 (N_2359,N_2253,N_2268);
nand U2360 (N_2360,N_2217,N_2256);
nor U2361 (N_2361,N_2234,N_2208);
nand U2362 (N_2362,N_2253,N_2203);
or U2363 (N_2363,N_2255,N_2289);
and U2364 (N_2364,N_2202,N_2250);
and U2365 (N_2365,N_2233,N_2210);
nor U2366 (N_2366,N_2245,N_2281);
xnor U2367 (N_2367,N_2277,N_2299);
or U2368 (N_2368,N_2218,N_2238);
xor U2369 (N_2369,N_2261,N_2283);
xor U2370 (N_2370,N_2233,N_2243);
nand U2371 (N_2371,N_2267,N_2205);
or U2372 (N_2372,N_2265,N_2249);
nor U2373 (N_2373,N_2263,N_2298);
nand U2374 (N_2374,N_2260,N_2207);
nor U2375 (N_2375,N_2229,N_2267);
nor U2376 (N_2376,N_2274,N_2252);
nor U2377 (N_2377,N_2263,N_2233);
or U2378 (N_2378,N_2215,N_2235);
nor U2379 (N_2379,N_2247,N_2266);
or U2380 (N_2380,N_2204,N_2233);
and U2381 (N_2381,N_2204,N_2240);
nand U2382 (N_2382,N_2205,N_2201);
nand U2383 (N_2383,N_2248,N_2268);
nor U2384 (N_2384,N_2204,N_2268);
nand U2385 (N_2385,N_2220,N_2295);
nand U2386 (N_2386,N_2242,N_2210);
nand U2387 (N_2387,N_2223,N_2273);
and U2388 (N_2388,N_2272,N_2245);
or U2389 (N_2389,N_2298,N_2248);
or U2390 (N_2390,N_2252,N_2206);
and U2391 (N_2391,N_2260,N_2281);
and U2392 (N_2392,N_2211,N_2281);
or U2393 (N_2393,N_2273,N_2214);
nor U2394 (N_2394,N_2258,N_2246);
nor U2395 (N_2395,N_2254,N_2231);
nor U2396 (N_2396,N_2209,N_2266);
or U2397 (N_2397,N_2209,N_2271);
nor U2398 (N_2398,N_2209,N_2249);
nor U2399 (N_2399,N_2225,N_2260);
nor U2400 (N_2400,N_2364,N_2330);
nor U2401 (N_2401,N_2313,N_2310);
xor U2402 (N_2402,N_2362,N_2356);
nor U2403 (N_2403,N_2319,N_2300);
nand U2404 (N_2404,N_2386,N_2388);
and U2405 (N_2405,N_2392,N_2399);
or U2406 (N_2406,N_2389,N_2385);
or U2407 (N_2407,N_2322,N_2374);
and U2408 (N_2408,N_2328,N_2382);
or U2409 (N_2409,N_2326,N_2303);
nor U2410 (N_2410,N_2355,N_2344);
and U2411 (N_2411,N_2312,N_2354);
or U2412 (N_2412,N_2357,N_2349);
nor U2413 (N_2413,N_2302,N_2376);
and U2414 (N_2414,N_2398,N_2338);
nand U2415 (N_2415,N_2383,N_2372);
nor U2416 (N_2416,N_2314,N_2375);
or U2417 (N_2417,N_2305,N_2324);
or U2418 (N_2418,N_2301,N_2323);
xor U2419 (N_2419,N_2352,N_2333);
nand U2420 (N_2420,N_2351,N_2315);
nor U2421 (N_2421,N_2304,N_2335);
nand U2422 (N_2422,N_2379,N_2308);
nand U2423 (N_2423,N_2337,N_2348);
and U2424 (N_2424,N_2371,N_2329);
and U2425 (N_2425,N_2395,N_2359);
or U2426 (N_2426,N_2306,N_2360);
and U2427 (N_2427,N_2361,N_2378);
and U2428 (N_2428,N_2368,N_2341);
or U2429 (N_2429,N_2396,N_2307);
nor U2430 (N_2430,N_2342,N_2334);
and U2431 (N_2431,N_2321,N_2390);
nand U2432 (N_2432,N_2370,N_2377);
nor U2433 (N_2433,N_2332,N_2346);
xnor U2434 (N_2434,N_2331,N_2369);
nor U2435 (N_2435,N_2340,N_2327);
or U2436 (N_2436,N_2343,N_2320);
and U2437 (N_2437,N_2373,N_2393);
xnor U2438 (N_2438,N_2397,N_2316);
nor U2439 (N_2439,N_2366,N_2318);
and U2440 (N_2440,N_2347,N_2358);
nand U2441 (N_2441,N_2339,N_2391);
nor U2442 (N_2442,N_2384,N_2309);
and U2443 (N_2443,N_2387,N_2365);
and U2444 (N_2444,N_2367,N_2350);
nand U2445 (N_2445,N_2381,N_2317);
xnor U2446 (N_2446,N_2311,N_2353);
xnor U2447 (N_2447,N_2336,N_2363);
nor U2448 (N_2448,N_2380,N_2325);
and U2449 (N_2449,N_2345,N_2394);
nand U2450 (N_2450,N_2331,N_2326);
nand U2451 (N_2451,N_2301,N_2331);
or U2452 (N_2452,N_2323,N_2316);
or U2453 (N_2453,N_2305,N_2350);
xnor U2454 (N_2454,N_2308,N_2306);
or U2455 (N_2455,N_2391,N_2395);
or U2456 (N_2456,N_2303,N_2346);
or U2457 (N_2457,N_2362,N_2344);
nand U2458 (N_2458,N_2374,N_2348);
nor U2459 (N_2459,N_2357,N_2345);
nand U2460 (N_2460,N_2335,N_2316);
and U2461 (N_2461,N_2369,N_2384);
nand U2462 (N_2462,N_2300,N_2350);
nand U2463 (N_2463,N_2303,N_2320);
nor U2464 (N_2464,N_2375,N_2352);
nand U2465 (N_2465,N_2378,N_2353);
nor U2466 (N_2466,N_2321,N_2359);
or U2467 (N_2467,N_2362,N_2376);
and U2468 (N_2468,N_2371,N_2368);
or U2469 (N_2469,N_2380,N_2372);
and U2470 (N_2470,N_2328,N_2394);
nor U2471 (N_2471,N_2388,N_2349);
nand U2472 (N_2472,N_2351,N_2369);
nor U2473 (N_2473,N_2373,N_2341);
nand U2474 (N_2474,N_2336,N_2346);
nor U2475 (N_2475,N_2365,N_2382);
nand U2476 (N_2476,N_2373,N_2330);
nand U2477 (N_2477,N_2307,N_2329);
or U2478 (N_2478,N_2343,N_2362);
or U2479 (N_2479,N_2387,N_2356);
and U2480 (N_2480,N_2384,N_2356);
nor U2481 (N_2481,N_2308,N_2344);
nor U2482 (N_2482,N_2355,N_2312);
and U2483 (N_2483,N_2393,N_2304);
and U2484 (N_2484,N_2327,N_2312);
nor U2485 (N_2485,N_2333,N_2313);
nand U2486 (N_2486,N_2367,N_2394);
nand U2487 (N_2487,N_2381,N_2334);
and U2488 (N_2488,N_2354,N_2360);
nor U2489 (N_2489,N_2307,N_2388);
nand U2490 (N_2490,N_2304,N_2385);
or U2491 (N_2491,N_2345,N_2343);
nand U2492 (N_2492,N_2372,N_2316);
and U2493 (N_2493,N_2369,N_2366);
xnor U2494 (N_2494,N_2397,N_2355);
xor U2495 (N_2495,N_2327,N_2362);
xnor U2496 (N_2496,N_2302,N_2371);
and U2497 (N_2497,N_2371,N_2393);
or U2498 (N_2498,N_2308,N_2386);
and U2499 (N_2499,N_2390,N_2323);
and U2500 (N_2500,N_2444,N_2493);
nand U2501 (N_2501,N_2407,N_2470);
nor U2502 (N_2502,N_2458,N_2468);
and U2503 (N_2503,N_2434,N_2474);
or U2504 (N_2504,N_2404,N_2400);
nor U2505 (N_2505,N_2473,N_2451);
nand U2506 (N_2506,N_2440,N_2438);
nand U2507 (N_2507,N_2463,N_2462);
and U2508 (N_2508,N_2431,N_2401);
or U2509 (N_2509,N_2478,N_2464);
xnor U2510 (N_2510,N_2467,N_2413);
nand U2511 (N_2511,N_2418,N_2454);
and U2512 (N_2512,N_2439,N_2410);
and U2513 (N_2513,N_2479,N_2452);
or U2514 (N_2514,N_2483,N_2442);
nor U2515 (N_2515,N_2417,N_2480);
or U2516 (N_2516,N_2406,N_2494);
and U2517 (N_2517,N_2497,N_2414);
nor U2518 (N_2518,N_2420,N_2455);
nand U2519 (N_2519,N_2476,N_2456);
nor U2520 (N_2520,N_2485,N_2446);
nor U2521 (N_2521,N_2492,N_2486);
nor U2522 (N_2522,N_2472,N_2402);
or U2523 (N_2523,N_2498,N_2419);
and U2524 (N_2524,N_2482,N_2430);
nor U2525 (N_2525,N_2465,N_2426);
nand U2526 (N_2526,N_2457,N_2499);
or U2527 (N_2527,N_2435,N_2437);
nand U2528 (N_2528,N_2460,N_2412);
nor U2529 (N_2529,N_2490,N_2469);
xnor U2530 (N_2530,N_2447,N_2484);
nor U2531 (N_2531,N_2495,N_2405);
and U2532 (N_2532,N_2441,N_2403);
nand U2533 (N_2533,N_2448,N_2461);
or U2534 (N_2534,N_2422,N_2475);
nand U2535 (N_2535,N_2487,N_2489);
and U2536 (N_2536,N_2423,N_2488);
xnor U2537 (N_2537,N_2429,N_2477);
xor U2538 (N_2538,N_2409,N_2449);
and U2539 (N_2539,N_2471,N_2481);
and U2540 (N_2540,N_2416,N_2428);
and U2541 (N_2541,N_2424,N_2408);
nor U2542 (N_2542,N_2496,N_2411);
and U2543 (N_2543,N_2453,N_2491);
xor U2544 (N_2544,N_2427,N_2433);
nand U2545 (N_2545,N_2415,N_2443);
nand U2546 (N_2546,N_2450,N_2425);
nor U2547 (N_2547,N_2432,N_2421);
xnor U2548 (N_2548,N_2445,N_2459);
xor U2549 (N_2549,N_2436,N_2466);
nand U2550 (N_2550,N_2413,N_2424);
nor U2551 (N_2551,N_2467,N_2430);
nor U2552 (N_2552,N_2415,N_2437);
or U2553 (N_2553,N_2450,N_2439);
or U2554 (N_2554,N_2422,N_2444);
nand U2555 (N_2555,N_2479,N_2494);
nor U2556 (N_2556,N_2437,N_2496);
or U2557 (N_2557,N_2413,N_2428);
or U2558 (N_2558,N_2468,N_2454);
and U2559 (N_2559,N_2416,N_2447);
and U2560 (N_2560,N_2424,N_2490);
nand U2561 (N_2561,N_2464,N_2481);
nor U2562 (N_2562,N_2483,N_2424);
and U2563 (N_2563,N_2420,N_2444);
and U2564 (N_2564,N_2442,N_2490);
nor U2565 (N_2565,N_2423,N_2477);
or U2566 (N_2566,N_2475,N_2479);
or U2567 (N_2567,N_2485,N_2455);
nor U2568 (N_2568,N_2408,N_2454);
nand U2569 (N_2569,N_2469,N_2403);
nand U2570 (N_2570,N_2480,N_2495);
or U2571 (N_2571,N_2417,N_2495);
nor U2572 (N_2572,N_2401,N_2492);
or U2573 (N_2573,N_2432,N_2473);
and U2574 (N_2574,N_2454,N_2435);
xnor U2575 (N_2575,N_2490,N_2493);
and U2576 (N_2576,N_2436,N_2432);
nor U2577 (N_2577,N_2408,N_2453);
nand U2578 (N_2578,N_2486,N_2497);
nor U2579 (N_2579,N_2498,N_2457);
and U2580 (N_2580,N_2459,N_2470);
nand U2581 (N_2581,N_2463,N_2431);
and U2582 (N_2582,N_2465,N_2406);
nor U2583 (N_2583,N_2447,N_2450);
nor U2584 (N_2584,N_2429,N_2450);
or U2585 (N_2585,N_2463,N_2404);
xor U2586 (N_2586,N_2402,N_2477);
and U2587 (N_2587,N_2412,N_2490);
or U2588 (N_2588,N_2402,N_2483);
or U2589 (N_2589,N_2451,N_2452);
nor U2590 (N_2590,N_2451,N_2401);
nand U2591 (N_2591,N_2471,N_2483);
and U2592 (N_2592,N_2432,N_2495);
and U2593 (N_2593,N_2449,N_2490);
nand U2594 (N_2594,N_2458,N_2431);
and U2595 (N_2595,N_2404,N_2432);
nand U2596 (N_2596,N_2496,N_2472);
nor U2597 (N_2597,N_2400,N_2483);
or U2598 (N_2598,N_2426,N_2461);
or U2599 (N_2599,N_2409,N_2403);
or U2600 (N_2600,N_2521,N_2554);
nand U2601 (N_2601,N_2520,N_2563);
nor U2602 (N_2602,N_2553,N_2541);
or U2603 (N_2603,N_2531,N_2509);
nand U2604 (N_2604,N_2548,N_2556);
nor U2605 (N_2605,N_2587,N_2591);
nor U2606 (N_2606,N_2524,N_2588);
and U2607 (N_2607,N_2551,N_2528);
and U2608 (N_2608,N_2533,N_2530);
nor U2609 (N_2609,N_2576,N_2523);
or U2610 (N_2610,N_2595,N_2580);
nand U2611 (N_2611,N_2557,N_2542);
nor U2612 (N_2612,N_2590,N_2532);
nand U2613 (N_2613,N_2577,N_2514);
nor U2614 (N_2614,N_2596,N_2510);
or U2615 (N_2615,N_2589,N_2584);
nor U2616 (N_2616,N_2566,N_2593);
or U2617 (N_2617,N_2581,N_2516);
nor U2618 (N_2618,N_2540,N_2561);
nor U2619 (N_2619,N_2578,N_2569);
and U2620 (N_2620,N_2547,N_2594);
nor U2621 (N_2621,N_2518,N_2529);
and U2622 (N_2622,N_2573,N_2568);
nor U2623 (N_2623,N_2574,N_2534);
or U2624 (N_2624,N_2599,N_2558);
or U2625 (N_2625,N_2539,N_2597);
nor U2626 (N_2626,N_2567,N_2544);
and U2627 (N_2627,N_2560,N_2503);
nand U2628 (N_2628,N_2545,N_2526);
and U2629 (N_2629,N_2527,N_2517);
nand U2630 (N_2630,N_2506,N_2582);
and U2631 (N_2631,N_2592,N_2512);
and U2632 (N_2632,N_2583,N_2570);
nand U2633 (N_2633,N_2511,N_2502);
and U2634 (N_2634,N_2549,N_2519);
nand U2635 (N_2635,N_2598,N_2513);
nor U2636 (N_2636,N_2537,N_2535);
or U2637 (N_2637,N_2571,N_2565);
nand U2638 (N_2638,N_2505,N_2515);
nor U2639 (N_2639,N_2525,N_2536);
or U2640 (N_2640,N_2572,N_2586);
nand U2641 (N_2641,N_2500,N_2564);
xor U2642 (N_2642,N_2579,N_2501);
xnor U2643 (N_2643,N_2507,N_2538);
nand U2644 (N_2644,N_2562,N_2550);
and U2645 (N_2645,N_2555,N_2559);
nand U2646 (N_2646,N_2585,N_2575);
or U2647 (N_2647,N_2504,N_2543);
or U2648 (N_2648,N_2546,N_2508);
nor U2649 (N_2649,N_2522,N_2552);
nand U2650 (N_2650,N_2546,N_2529);
or U2651 (N_2651,N_2538,N_2530);
and U2652 (N_2652,N_2567,N_2528);
and U2653 (N_2653,N_2573,N_2562);
and U2654 (N_2654,N_2593,N_2509);
nand U2655 (N_2655,N_2532,N_2504);
nor U2656 (N_2656,N_2536,N_2562);
and U2657 (N_2657,N_2567,N_2502);
and U2658 (N_2658,N_2500,N_2544);
or U2659 (N_2659,N_2553,N_2589);
xor U2660 (N_2660,N_2580,N_2553);
and U2661 (N_2661,N_2583,N_2564);
and U2662 (N_2662,N_2545,N_2511);
xnor U2663 (N_2663,N_2545,N_2508);
nand U2664 (N_2664,N_2514,N_2575);
nor U2665 (N_2665,N_2525,N_2507);
xor U2666 (N_2666,N_2555,N_2546);
nor U2667 (N_2667,N_2516,N_2578);
nand U2668 (N_2668,N_2520,N_2571);
nand U2669 (N_2669,N_2513,N_2544);
nand U2670 (N_2670,N_2529,N_2505);
and U2671 (N_2671,N_2563,N_2515);
nor U2672 (N_2672,N_2585,N_2554);
and U2673 (N_2673,N_2561,N_2553);
nor U2674 (N_2674,N_2521,N_2510);
nor U2675 (N_2675,N_2500,N_2587);
xnor U2676 (N_2676,N_2582,N_2507);
xor U2677 (N_2677,N_2521,N_2570);
nor U2678 (N_2678,N_2567,N_2508);
nor U2679 (N_2679,N_2557,N_2507);
or U2680 (N_2680,N_2539,N_2565);
nand U2681 (N_2681,N_2575,N_2508);
nand U2682 (N_2682,N_2523,N_2502);
nand U2683 (N_2683,N_2513,N_2548);
nor U2684 (N_2684,N_2581,N_2571);
nand U2685 (N_2685,N_2512,N_2513);
xor U2686 (N_2686,N_2500,N_2536);
xor U2687 (N_2687,N_2599,N_2547);
and U2688 (N_2688,N_2539,N_2574);
nor U2689 (N_2689,N_2557,N_2503);
and U2690 (N_2690,N_2573,N_2581);
or U2691 (N_2691,N_2508,N_2500);
xnor U2692 (N_2692,N_2516,N_2528);
or U2693 (N_2693,N_2522,N_2544);
nand U2694 (N_2694,N_2592,N_2532);
nand U2695 (N_2695,N_2583,N_2512);
and U2696 (N_2696,N_2570,N_2563);
and U2697 (N_2697,N_2550,N_2574);
nand U2698 (N_2698,N_2576,N_2571);
nor U2699 (N_2699,N_2509,N_2597);
xor U2700 (N_2700,N_2688,N_2604);
nand U2701 (N_2701,N_2665,N_2620);
nor U2702 (N_2702,N_2606,N_2649);
or U2703 (N_2703,N_2648,N_2615);
or U2704 (N_2704,N_2651,N_2694);
nor U2705 (N_2705,N_2643,N_2631);
and U2706 (N_2706,N_2674,N_2669);
and U2707 (N_2707,N_2600,N_2605);
or U2708 (N_2708,N_2610,N_2660);
and U2709 (N_2709,N_2612,N_2607);
nand U2710 (N_2710,N_2618,N_2636);
and U2711 (N_2711,N_2638,N_2642);
and U2712 (N_2712,N_2623,N_2690);
nor U2713 (N_2713,N_2678,N_2691);
or U2714 (N_2714,N_2661,N_2680);
and U2715 (N_2715,N_2628,N_2699);
and U2716 (N_2716,N_2656,N_2632);
or U2717 (N_2717,N_2622,N_2676);
nand U2718 (N_2718,N_2626,N_2639);
nand U2719 (N_2719,N_2663,N_2617);
nand U2720 (N_2720,N_2664,N_2602);
nand U2721 (N_2721,N_2670,N_2689);
and U2722 (N_2722,N_2673,N_2629);
xnor U2723 (N_2723,N_2662,N_2653);
nand U2724 (N_2724,N_2698,N_2697);
xor U2725 (N_2725,N_2646,N_2667);
or U2726 (N_2726,N_2640,N_2672);
or U2727 (N_2727,N_2645,N_2654);
nor U2728 (N_2728,N_2637,N_2635);
xnor U2729 (N_2729,N_2686,N_2652);
xnor U2730 (N_2730,N_2601,N_2695);
or U2731 (N_2731,N_2677,N_2693);
and U2732 (N_2732,N_2633,N_2641);
and U2733 (N_2733,N_2644,N_2658);
and U2734 (N_2734,N_2692,N_2621);
and U2735 (N_2735,N_2616,N_2668);
nand U2736 (N_2736,N_2647,N_2681);
xnor U2737 (N_2737,N_2655,N_2630);
and U2738 (N_2738,N_2666,N_2679);
or U2739 (N_2739,N_2619,N_2609);
nand U2740 (N_2740,N_2671,N_2650);
nor U2741 (N_2741,N_2603,N_2657);
or U2742 (N_2742,N_2611,N_2624);
nor U2743 (N_2743,N_2634,N_2627);
and U2744 (N_2744,N_2687,N_2685);
or U2745 (N_2745,N_2614,N_2683);
or U2746 (N_2746,N_2675,N_2608);
xnor U2747 (N_2747,N_2613,N_2684);
nor U2748 (N_2748,N_2659,N_2696);
nand U2749 (N_2749,N_2625,N_2682);
nand U2750 (N_2750,N_2647,N_2646);
and U2751 (N_2751,N_2689,N_2673);
nor U2752 (N_2752,N_2656,N_2600);
nand U2753 (N_2753,N_2662,N_2650);
nand U2754 (N_2754,N_2612,N_2674);
nor U2755 (N_2755,N_2697,N_2624);
xor U2756 (N_2756,N_2619,N_2662);
nand U2757 (N_2757,N_2636,N_2668);
nor U2758 (N_2758,N_2634,N_2673);
nand U2759 (N_2759,N_2614,N_2654);
and U2760 (N_2760,N_2663,N_2696);
or U2761 (N_2761,N_2648,N_2684);
nand U2762 (N_2762,N_2658,N_2641);
nand U2763 (N_2763,N_2633,N_2690);
and U2764 (N_2764,N_2617,N_2681);
nor U2765 (N_2765,N_2643,N_2682);
nor U2766 (N_2766,N_2610,N_2607);
nor U2767 (N_2767,N_2695,N_2620);
and U2768 (N_2768,N_2620,N_2601);
or U2769 (N_2769,N_2606,N_2697);
nor U2770 (N_2770,N_2685,N_2611);
or U2771 (N_2771,N_2607,N_2693);
and U2772 (N_2772,N_2692,N_2684);
and U2773 (N_2773,N_2661,N_2646);
or U2774 (N_2774,N_2634,N_2611);
nand U2775 (N_2775,N_2655,N_2615);
and U2776 (N_2776,N_2648,N_2677);
nand U2777 (N_2777,N_2640,N_2648);
or U2778 (N_2778,N_2671,N_2651);
nand U2779 (N_2779,N_2613,N_2632);
or U2780 (N_2780,N_2640,N_2628);
xnor U2781 (N_2781,N_2663,N_2671);
and U2782 (N_2782,N_2676,N_2671);
or U2783 (N_2783,N_2685,N_2604);
nand U2784 (N_2784,N_2689,N_2692);
and U2785 (N_2785,N_2661,N_2660);
and U2786 (N_2786,N_2665,N_2644);
nand U2787 (N_2787,N_2669,N_2684);
and U2788 (N_2788,N_2664,N_2634);
nor U2789 (N_2789,N_2616,N_2672);
nor U2790 (N_2790,N_2650,N_2667);
nand U2791 (N_2791,N_2672,N_2663);
and U2792 (N_2792,N_2616,N_2636);
or U2793 (N_2793,N_2634,N_2662);
nor U2794 (N_2794,N_2625,N_2670);
and U2795 (N_2795,N_2636,N_2640);
nand U2796 (N_2796,N_2690,N_2630);
nor U2797 (N_2797,N_2674,N_2601);
nor U2798 (N_2798,N_2673,N_2619);
or U2799 (N_2799,N_2666,N_2612);
nand U2800 (N_2800,N_2776,N_2751);
and U2801 (N_2801,N_2724,N_2710);
or U2802 (N_2802,N_2770,N_2764);
nor U2803 (N_2803,N_2763,N_2754);
and U2804 (N_2804,N_2740,N_2775);
nand U2805 (N_2805,N_2708,N_2767);
and U2806 (N_2806,N_2747,N_2753);
and U2807 (N_2807,N_2795,N_2705);
nand U2808 (N_2808,N_2723,N_2784);
or U2809 (N_2809,N_2756,N_2755);
nand U2810 (N_2810,N_2752,N_2716);
or U2811 (N_2811,N_2771,N_2766);
nand U2812 (N_2812,N_2799,N_2703);
xnor U2813 (N_2813,N_2717,N_2727);
nor U2814 (N_2814,N_2790,N_2701);
nand U2815 (N_2815,N_2736,N_2748);
nor U2816 (N_2816,N_2725,N_2792);
nand U2817 (N_2817,N_2788,N_2741);
nand U2818 (N_2818,N_2706,N_2712);
or U2819 (N_2819,N_2729,N_2787);
nand U2820 (N_2820,N_2772,N_2789);
nand U2821 (N_2821,N_2750,N_2738);
or U2822 (N_2822,N_2715,N_2700);
nor U2823 (N_2823,N_2720,N_2782);
or U2824 (N_2824,N_2728,N_2735);
nor U2825 (N_2825,N_2704,N_2732);
nor U2826 (N_2826,N_2757,N_2737);
nor U2827 (N_2827,N_2733,N_2734);
and U2828 (N_2828,N_2768,N_2722);
xor U2829 (N_2829,N_2713,N_2797);
nor U2830 (N_2830,N_2709,N_2746);
nand U2831 (N_2831,N_2783,N_2726);
nand U2832 (N_2832,N_2780,N_2798);
xnor U2833 (N_2833,N_2786,N_2739);
nand U2834 (N_2834,N_2745,N_2759);
xor U2835 (N_2835,N_2796,N_2742);
xnor U2836 (N_2836,N_2707,N_2779);
or U2837 (N_2837,N_2794,N_2730);
nor U2838 (N_2838,N_2711,N_2791);
and U2839 (N_2839,N_2765,N_2718);
xor U2840 (N_2840,N_2761,N_2744);
nor U2841 (N_2841,N_2719,N_2778);
or U2842 (N_2842,N_2758,N_2731);
or U2843 (N_2843,N_2760,N_2721);
or U2844 (N_2844,N_2785,N_2773);
nor U2845 (N_2845,N_2702,N_2777);
nor U2846 (N_2846,N_2762,N_2714);
nand U2847 (N_2847,N_2793,N_2781);
nor U2848 (N_2848,N_2749,N_2743);
xnor U2849 (N_2849,N_2769,N_2774);
nor U2850 (N_2850,N_2705,N_2744);
nand U2851 (N_2851,N_2770,N_2789);
nor U2852 (N_2852,N_2739,N_2720);
and U2853 (N_2853,N_2753,N_2786);
nor U2854 (N_2854,N_2722,N_2741);
xnor U2855 (N_2855,N_2732,N_2731);
nor U2856 (N_2856,N_2744,N_2732);
nand U2857 (N_2857,N_2767,N_2741);
nor U2858 (N_2858,N_2715,N_2723);
nand U2859 (N_2859,N_2735,N_2773);
or U2860 (N_2860,N_2770,N_2776);
or U2861 (N_2861,N_2791,N_2737);
and U2862 (N_2862,N_2791,N_2793);
or U2863 (N_2863,N_2712,N_2719);
and U2864 (N_2864,N_2732,N_2782);
and U2865 (N_2865,N_2792,N_2714);
nand U2866 (N_2866,N_2711,N_2709);
or U2867 (N_2867,N_2700,N_2794);
xnor U2868 (N_2868,N_2718,N_2743);
and U2869 (N_2869,N_2760,N_2789);
nor U2870 (N_2870,N_2788,N_2773);
and U2871 (N_2871,N_2730,N_2763);
and U2872 (N_2872,N_2755,N_2742);
and U2873 (N_2873,N_2739,N_2793);
nand U2874 (N_2874,N_2719,N_2769);
or U2875 (N_2875,N_2714,N_2753);
nor U2876 (N_2876,N_2747,N_2763);
nand U2877 (N_2877,N_2739,N_2754);
and U2878 (N_2878,N_2780,N_2760);
or U2879 (N_2879,N_2713,N_2711);
or U2880 (N_2880,N_2714,N_2716);
or U2881 (N_2881,N_2724,N_2768);
or U2882 (N_2882,N_2728,N_2741);
nand U2883 (N_2883,N_2763,N_2701);
or U2884 (N_2884,N_2790,N_2726);
and U2885 (N_2885,N_2795,N_2736);
or U2886 (N_2886,N_2723,N_2782);
and U2887 (N_2887,N_2777,N_2738);
and U2888 (N_2888,N_2732,N_2711);
and U2889 (N_2889,N_2702,N_2793);
nand U2890 (N_2890,N_2730,N_2753);
or U2891 (N_2891,N_2795,N_2714);
or U2892 (N_2892,N_2792,N_2742);
nand U2893 (N_2893,N_2701,N_2735);
and U2894 (N_2894,N_2719,N_2797);
or U2895 (N_2895,N_2733,N_2747);
nor U2896 (N_2896,N_2784,N_2756);
or U2897 (N_2897,N_2751,N_2732);
and U2898 (N_2898,N_2710,N_2736);
or U2899 (N_2899,N_2703,N_2735);
nand U2900 (N_2900,N_2893,N_2825);
nor U2901 (N_2901,N_2819,N_2889);
and U2902 (N_2902,N_2809,N_2865);
and U2903 (N_2903,N_2859,N_2858);
xor U2904 (N_2904,N_2830,N_2860);
nor U2905 (N_2905,N_2872,N_2895);
or U2906 (N_2906,N_2879,N_2815);
and U2907 (N_2907,N_2814,N_2840);
or U2908 (N_2908,N_2861,N_2854);
nand U2909 (N_2909,N_2803,N_2816);
and U2910 (N_2910,N_2882,N_2826);
xor U2911 (N_2911,N_2802,N_2828);
nor U2912 (N_2912,N_2834,N_2876);
and U2913 (N_2913,N_2898,N_2870);
nand U2914 (N_2914,N_2884,N_2863);
and U2915 (N_2915,N_2899,N_2806);
nor U2916 (N_2916,N_2837,N_2812);
nor U2917 (N_2917,N_2843,N_2867);
or U2918 (N_2918,N_2810,N_2857);
and U2919 (N_2919,N_2888,N_2887);
nand U2920 (N_2920,N_2801,N_2846);
and U2921 (N_2921,N_2877,N_2841);
nand U2922 (N_2922,N_2896,N_2866);
xor U2923 (N_2923,N_2847,N_2852);
or U2924 (N_2924,N_2845,N_2856);
nand U2925 (N_2925,N_2850,N_2868);
nor U2926 (N_2926,N_2823,N_2851);
nor U2927 (N_2927,N_2832,N_2805);
nor U2928 (N_2928,N_2892,N_2897);
or U2929 (N_2929,N_2848,N_2849);
nand U2930 (N_2930,N_2875,N_2883);
and U2931 (N_2931,N_2821,N_2873);
and U2932 (N_2932,N_2894,N_2890);
nand U2933 (N_2933,N_2833,N_2835);
and U2934 (N_2934,N_2813,N_2804);
nand U2935 (N_2935,N_2817,N_2878);
nand U2936 (N_2936,N_2886,N_2829);
and U2937 (N_2937,N_2807,N_2831);
nand U2938 (N_2938,N_2808,N_2874);
nand U2939 (N_2939,N_2836,N_2800);
or U2940 (N_2940,N_2842,N_2822);
nor U2941 (N_2941,N_2881,N_2824);
nor U2942 (N_2942,N_2871,N_2869);
nor U2943 (N_2943,N_2885,N_2839);
and U2944 (N_2944,N_2862,N_2880);
nand U2945 (N_2945,N_2818,N_2855);
nor U2946 (N_2946,N_2811,N_2827);
nand U2947 (N_2947,N_2838,N_2891);
nand U2948 (N_2948,N_2844,N_2853);
nand U2949 (N_2949,N_2864,N_2820);
or U2950 (N_2950,N_2883,N_2856);
nor U2951 (N_2951,N_2865,N_2860);
nand U2952 (N_2952,N_2888,N_2884);
or U2953 (N_2953,N_2843,N_2800);
nor U2954 (N_2954,N_2870,N_2880);
and U2955 (N_2955,N_2823,N_2866);
nor U2956 (N_2956,N_2824,N_2832);
nor U2957 (N_2957,N_2886,N_2869);
or U2958 (N_2958,N_2899,N_2844);
and U2959 (N_2959,N_2808,N_2891);
nand U2960 (N_2960,N_2888,N_2839);
and U2961 (N_2961,N_2803,N_2827);
and U2962 (N_2962,N_2843,N_2834);
or U2963 (N_2963,N_2808,N_2803);
or U2964 (N_2964,N_2800,N_2835);
or U2965 (N_2965,N_2878,N_2849);
and U2966 (N_2966,N_2859,N_2841);
and U2967 (N_2967,N_2807,N_2855);
or U2968 (N_2968,N_2880,N_2839);
nor U2969 (N_2969,N_2861,N_2864);
xor U2970 (N_2970,N_2833,N_2844);
and U2971 (N_2971,N_2820,N_2844);
nor U2972 (N_2972,N_2830,N_2845);
nor U2973 (N_2973,N_2882,N_2868);
and U2974 (N_2974,N_2841,N_2852);
or U2975 (N_2975,N_2899,N_2853);
xnor U2976 (N_2976,N_2862,N_2867);
or U2977 (N_2977,N_2864,N_2819);
and U2978 (N_2978,N_2873,N_2831);
xnor U2979 (N_2979,N_2821,N_2816);
or U2980 (N_2980,N_2894,N_2840);
nor U2981 (N_2981,N_2825,N_2804);
nor U2982 (N_2982,N_2817,N_2865);
xnor U2983 (N_2983,N_2830,N_2854);
nand U2984 (N_2984,N_2835,N_2830);
or U2985 (N_2985,N_2833,N_2884);
xor U2986 (N_2986,N_2870,N_2871);
xnor U2987 (N_2987,N_2805,N_2879);
nand U2988 (N_2988,N_2810,N_2843);
xnor U2989 (N_2989,N_2852,N_2818);
or U2990 (N_2990,N_2878,N_2899);
and U2991 (N_2991,N_2877,N_2886);
nor U2992 (N_2992,N_2861,N_2890);
nor U2993 (N_2993,N_2814,N_2855);
or U2994 (N_2994,N_2890,N_2853);
nand U2995 (N_2995,N_2804,N_2851);
and U2996 (N_2996,N_2885,N_2820);
or U2997 (N_2997,N_2863,N_2873);
xnor U2998 (N_2998,N_2859,N_2862);
nor U2999 (N_2999,N_2846,N_2872);
xnor UO_0 (O_0,N_2999,N_2966);
or UO_1 (O_1,N_2901,N_2997);
nor UO_2 (O_2,N_2926,N_2962);
and UO_3 (O_3,N_2985,N_2956);
nand UO_4 (O_4,N_2964,N_2935);
nor UO_5 (O_5,N_2909,N_2971);
nand UO_6 (O_6,N_2900,N_2978);
nand UO_7 (O_7,N_2994,N_2911);
or UO_8 (O_8,N_2995,N_2979);
and UO_9 (O_9,N_2970,N_2948);
nor UO_10 (O_10,N_2986,N_2975);
nor UO_11 (O_11,N_2980,N_2912);
xor UO_12 (O_12,N_2936,N_2907);
xor UO_13 (O_13,N_2944,N_2902);
or UO_14 (O_14,N_2928,N_2998);
nand UO_15 (O_15,N_2996,N_2968);
nand UO_16 (O_16,N_2977,N_2941);
nor UO_17 (O_17,N_2989,N_2992);
and UO_18 (O_18,N_2987,N_2984);
nand UO_19 (O_19,N_2967,N_2945);
nand UO_20 (O_20,N_2933,N_2934);
xnor UO_21 (O_21,N_2908,N_2983);
and UO_22 (O_22,N_2939,N_2957);
and UO_23 (O_23,N_2981,N_2915);
or UO_24 (O_24,N_2931,N_2958);
nand UO_25 (O_25,N_2924,N_2917);
and UO_26 (O_26,N_2969,N_2918);
or UO_27 (O_27,N_2930,N_2914);
or UO_28 (O_28,N_2993,N_2929);
or UO_29 (O_29,N_2988,N_2932);
xnor UO_30 (O_30,N_2953,N_2910);
and UO_31 (O_31,N_2972,N_2974);
xor UO_32 (O_32,N_2904,N_2946);
nor UO_33 (O_33,N_2991,N_2965);
and UO_34 (O_34,N_2959,N_2973);
and UO_35 (O_35,N_2937,N_2919);
xor UO_36 (O_36,N_2951,N_2922);
or UO_37 (O_37,N_2921,N_2954);
nand UO_38 (O_38,N_2942,N_2916);
or UO_39 (O_39,N_2949,N_2920);
nor UO_40 (O_40,N_2955,N_2976);
nor UO_41 (O_41,N_2990,N_2903);
or UO_42 (O_42,N_2905,N_2950);
and UO_43 (O_43,N_2952,N_2960);
nand UO_44 (O_44,N_2943,N_2927);
and UO_45 (O_45,N_2906,N_2982);
nor UO_46 (O_46,N_2947,N_2925);
xnor UO_47 (O_47,N_2913,N_2923);
nand UO_48 (O_48,N_2938,N_2940);
and UO_49 (O_49,N_2961,N_2963);
or UO_50 (O_50,N_2911,N_2909);
nand UO_51 (O_51,N_2962,N_2932);
or UO_52 (O_52,N_2953,N_2991);
nor UO_53 (O_53,N_2938,N_2944);
xnor UO_54 (O_54,N_2927,N_2998);
xor UO_55 (O_55,N_2949,N_2900);
and UO_56 (O_56,N_2997,N_2912);
nor UO_57 (O_57,N_2998,N_2934);
nand UO_58 (O_58,N_2942,N_2979);
nor UO_59 (O_59,N_2902,N_2962);
nor UO_60 (O_60,N_2931,N_2905);
nand UO_61 (O_61,N_2965,N_2977);
or UO_62 (O_62,N_2968,N_2911);
xnor UO_63 (O_63,N_2912,N_2991);
or UO_64 (O_64,N_2929,N_2989);
and UO_65 (O_65,N_2945,N_2934);
xor UO_66 (O_66,N_2968,N_2930);
nand UO_67 (O_67,N_2905,N_2924);
nand UO_68 (O_68,N_2900,N_2916);
xor UO_69 (O_69,N_2934,N_2962);
xor UO_70 (O_70,N_2981,N_2989);
and UO_71 (O_71,N_2988,N_2913);
xor UO_72 (O_72,N_2937,N_2942);
nand UO_73 (O_73,N_2967,N_2949);
nand UO_74 (O_74,N_2976,N_2960);
nor UO_75 (O_75,N_2906,N_2913);
and UO_76 (O_76,N_2906,N_2943);
xnor UO_77 (O_77,N_2933,N_2956);
or UO_78 (O_78,N_2904,N_2954);
or UO_79 (O_79,N_2946,N_2924);
xor UO_80 (O_80,N_2945,N_2909);
and UO_81 (O_81,N_2932,N_2925);
or UO_82 (O_82,N_2901,N_2907);
nand UO_83 (O_83,N_2902,N_2967);
or UO_84 (O_84,N_2971,N_2958);
nand UO_85 (O_85,N_2938,N_2943);
and UO_86 (O_86,N_2947,N_2996);
or UO_87 (O_87,N_2987,N_2946);
xor UO_88 (O_88,N_2964,N_2997);
or UO_89 (O_89,N_2906,N_2963);
nor UO_90 (O_90,N_2903,N_2963);
nand UO_91 (O_91,N_2972,N_2947);
nand UO_92 (O_92,N_2935,N_2930);
xnor UO_93 (O_93,N_2957,N_2975);
or UO_94 (O_94,N_2936,N_2992);
nand UO_95 (O_95,N_2972,N_2940);
nor UO_96 (O_96,N_2964,N_2922);
nand UO_97 (O_97,N_2911,N_2967);
or UO_98 (O_98,N_2917,N_2935);
and UO_99 (O_99,N_2963,N_2968);
nor UO_100 (O_100,N_2981,N_2961);
or UO_101 (O_101,N_2985,N_2908);
nor UO_102 (O_102,N_2924,N_2940);
nor UO_103 (O_103,N_2926,N_2905);
or UO_104 (O_104,N_2994,N_2948);
nand UO_105 (O_105,N_2940,N_2956);
nand UO_106 (O_106,N_2924,N_2902);
and UO_107 (O_107,N_2998,N_2982);
nor UO_108 (O_108,N_2970,N_2934);
or UO_109 (O_109,N_2939,N_2996);
or UO_110 (O_110,N_2955,N_2915);
nor UO_111 (O_111,N_2933,N_2920);
nor UO_112 (O_112,N_2925,N_2938);
or UO_113 (O_113,N_2982,N_2977);
nand UO_114 (O_114,N_2961,N_2900);
nand UO_115 (O_115,N_2915,N_2923);
nand UO_116 (O_116,N_2953,N_2913);
or UO_117 (O_117,N_2975,N_2989);
nand UO_118 (O_118,N_2992,N_2910);
xor UO_119 (O_119,N_2965,N_2939);
and UO_120 (O_120,N_2974,N_2921);
nand UO_121 (O_121,N_2970,N_2960);
nor UO_122 (O_122,N_2959,N_2908);
nand UO_123 (O_123,N_2923,N_2984);
nor UO_124 (O_124,N_2989,N_2908);
nor UO_125 (O_125,N_2962,N_2938);
nand UO_126 (O_126,N_2967,N_2981);
and UO_127 (O_127,N_2942,N_2952);
nand UO_128 (O_128,N_2972,N_2954);
and UO_129 (O_129,N_2912,N_2959);
and UO_130 (O_130,N_2956,N_2984);
nor UO_131 (O_131,N_2955,N_2993);
nand UO_132 (O_132,N_2931,N_2975);
and UO_133 (O_133,N_2996,N_2922);
nor UO_134 (O_134,N_2962,N_2942);
nand UO_135 (O_135,N_2907,N_2974);
nor UO_136 (O_136,N_2903,N_2920);
or UO_137 (O_137,N_2996,N_2982);
nand UO_138 (O_138,N_2984,N_2950);
and UO_139 (O_139,N_2901,N_2964);
and UO_140 (O_140,N_2979,N_2994);
nand UO_141 (O_141,N_2906,N_2981);
nand UO_142 (O_142,N_2952,N_2948);
or UO_143 (O_143,N_2994,N_2952);
nand UO_144 (O_144,N_2918,N_2924);
nand UO_145 (O_145,N_2993,N_2939);
nand UO_146 (O_146,N_2968,N_2922);
nor UO_147 (O_147,N_2935,N_2927);
and UO_148 (O_148,N_2912,N_2924);
nand UO_149 (O_149,N_2976,N_2987);
nand UO_150 (O_150,N_2973,N_2914);
nor UO_151 (O_151,N_2975,N_2944);
and UO_152 (O_152,N_2977,N_2909);
nand UO_153 (O_153,N_2963,N_2973);
and UO_154 (O_154,N_2996,N_2985);
or UO_155 (O_155,N_2997,N_2914);
nor UO_156 (O_156,N_2939,N_2924);
nor UO_157 (O_157,N_2939,N_2972);
xnor UO_158 (O_158,N_2944,N_2961);
nor UO_159 (O_159,N_2952,N_2980);
or UO_160 (O_160,N_2912,N_2937);
nand UO_161 (O_161,N_2910,N_2942);
nor UO_162 (O_162,N_2907,N_2957);
nor UO_163 (O_163,N_2931,N_2981);
or UO_164 (O_164,N_2983,N_2918);
nor UO_165 (O_165,N_2978,N_2945);
nand UO_166 (O_166,N_2967,N_2966);
nor UO_167 (O_167,N_2948,N_2901);
nand UO_168 (O_168,N_2974,N_2989);
nand UO_169 (O_169,N_2952,N_2966);
nand UO_170 (O_170,N_2926,N_2986);
or UO_171 (O_171,N_2999,N_2977);
and UO_172 (O_172,N_2913,N_2950);
or UO_173 (O_173,N_2984,N_2925);
xor UO_174 (O_174,N_2973,N_2945);
nand UO_175 (O_175,N_2909,N_2918);
nor UO_176 (O_176,N_2928,N_2905);
xor UO_177 (O_177,N_2982,N_2965);
or UO_178 (O_178,N_2982,N_2957);
and UO_179 (O_179,N_2984,N_2976);
and UO_180 (O_180,N_2946,N_2993);
nor UO_181 (O_181,N_2985,N_2951);
xor UO_182 (O_182,N_2956,N_2941);
or UO_183 (O_183,N_2935,N_2916);
nor UO_184 (O_184,N_2970,N_2980);
and UO_185 (O_185,N_2928,N_2991);
nor UO_186 (O_186,N_2973,N_2965);
or UO_187 (O_187,N_2950,N_2996);
nand UO_188 (O_188,N_2976,N_2995);
nand UO_189 (O_189,N_2998,N_2977);
nor UO_190 (O_190,N_2951,N_2983);
or UO_191 (O_191,N_2989,N_2907);
nor UO_192 (O_192,N_2986,N_2984);
and UO_193 (O_193,N_2972,N_2943);
or UO_194 (O_194,N_2971,N_2906);
or UO_195 (O_195,N_2913,N_2990);
and UO_196 (O_196,N_2978,N_2910);
nor UO_197 (O_197,N_2949,N_2907);
nor UO_198 (O_198,N_2900,N_2960);
or UO_199 (O_199,N_2972,N_2992);
or UO_200 (O_200,N_2930,N_2995);
or UO_201 (O_201,N_2937,N_2940);
or UO_202 (O_202,N_2964,N_2932);
nor UO_203 (O_203,N_2988,N_2906);
nor UO_204 (O_204,N_2957,N_2962);
or UO_205 (O_205,N_2911,N_2938);
or UO_206 (O_206,N_2904,N_2912);
or UO_207 (O_207,N_2913,N_2939);
and UO_208 (O_208,N_2921,N_2933);
and UO_209 (O_209,N_2925,N_2985);
nor UO_210 (O_210,N_2980,N_2963);
and UO_211 (O_211,N_2932,N_2917);
or UO_212 (O_212,N_2924,N_2954);
and UO_213 (O_213,N_2975,N_2949);
or UO_214 (O_214,N_2998,N_2960);
or UO_215 (O_215,N_2913,N_2928);
xnor UO_216 (O_216,N_2975,N_2951);
xor UO_217 (O_217,N_2933,N_2932);
or UO_218 (O_218,N_2916,N_2933);
xnor UO_219 (O_219,N_2905,N_2951);
or UO_220 (O_220,N_2911,N_2925);
nor UO_221 (O_221,N_2928,N_2967);
nand UO_222 (O_222,N_2968,N_2939);
and UO_223 (O_223,N_2991,N_2931);
or UO_224 (O_224,N_2953,N_2946);
nor UO_225 (O_225,N_2950,N_2983);
nand UO_226 (O_226,N_2942,N_2982);
and UO_227 (O_227,N_2930,N_2916);
nor UO_228 (O_228,N_2980,N_2951);
nor UO_229 (O_229,N_2983,N_2955);
and UO_230 (O_230,N_2992,N_2909);
nor UO_231 (O_231,N_2932,N_2902);
nor UO_232 (O_232,N_2906,N_2954);
or UO_233 (O_233,N_2970,N_2958);
xor UO_234 (O_234,N_2979,N_2980);
nor UO_235 (O_235,N_2950,N_2975);
nor UO_236 (O_236,N_2927,N_2965);
and UO_237 (O_237,N_2900,N_2982);
or UO_238 (O_238,N_2962,N_2958);
nand UO_239 (O_239,N_2940,N_2982);
nand UO_240 (O_240,N_2902,N_2951);
and UO_241 (O_241,N_2942,N_2922);
and UO_242 (O_242,N_2936,N_2904);
nor UO_243 (O_243,N_2983,N_2978);
or UO_244 (O_244,N_2926,N_2915);
xor UO_245 (O_245,N_2966,N_2945);
nor UO_246 (O_246,N_2915,N_2956);
or UO_247 (O_247,N_2944,N_2970);
nor UO_248 (O_248,N_2934,N_2954);
or UO_249 (O_249,N_2926,N_2928);
xnor UO_250 (O_250,N_2947,N_2951);
nand UO_251 (O_251,N_2900,N_2974);
nand UO_252 (O_252,N_2941,N_2938);
nand UO_253 (O_253,N_2964,N_2927);
and UO_254 (O_254,N_2996,N_2907);
and UO_255 (O_255,N_2927,N_2937);
nor UO_256 (O_256,N_2977,N_2973);
nand UO_257 (O_257,N_2914,N_2947);
and UO_258 (O_258,N_2970,N_2952);
and UO_259 (O_259,N_2970,N_2907);
nand UO_260 (O_260,N_2937,N_2989);
or UO_261 (O_261,N_2943,N_2920);
and UO_262 (O_262,N_2908,N_2902);
or UO_263 (O_263,N_2937,N_2953);
nor UO_264 (O_264,N_2963,N_2945);
nand UO_265 (O_265,N_2967,N_2940);
nand UO_266 (O_266,N_2923,N_2998);
and UO_267 (O_267,N_2940,N_2998);
or UO_268 (O_268,N_2939,N_2974);
xor UO_269 (O_269,N_2994,N_2933);
or UO_270 (O_270,N_2907,N_2959);
nand UO_271 (O_271,N_2948,N_2979);
nor UO_272 (O_272,N_2973,N_2942);
nand UO_273 (O_273,N_2904,N_2910);
or UO_274 (O_274,N_2991,N_2910);
xor UO_275 (O_275,N_2944,N_2980);
nor UO_276 (O_276,N_2970,N_2923);
xnor UO_277 (O_277,N_2961,N_2988);
xor UO_278 (O_278,N_2959,N_2991);
nand UO_279 (O_279,N_2967,N_2927);
or UO_280 (O_280,N_2906,N_2931);
or UO_281 (O_281,N_2912,N_2988);
nor UO_282 (O_282,N_2900,N_2937);
nor UO_283 (O_283,N_2960,N_2939);
nor UO_284 (O_284,N_2999,N_2947);
nand UO_285 (O_285,N_2962,N_2982);
xnor UO_286 (O_286,N_2973,N_2946);
and UO_287 (O_287,N_2920,N_2912);
and UO_288 (O_288,N_2993,N_2934);
or UO_289 (O_289,N_2945,N_2952);
nor UO_290 (O_290,N_2942,N_2919);
nand UO_291 (O_291,N_2971,N_2905);
and UO_292 (O_292,N_2966,N_2985);
nor UO_293 (O_293,N_2982,N_2999);
and UO_294 (O_294,N_2986,N_2993);
or UO_295 (O_295,N_2918,N_2962);
and UO_296 (O_296,N_2965,N_2942);
and UO_297 (O_297,N_2935,N_2979);
xor UO_298 (O_298,N_2918,N_2953);
nand UO_299 (O_299,N_2934,N_2943);
and UO_300 (O_300,N_2901,N_2995);
and UO_301 (O_301,N_2994,N_2913);
or UO_302 (O_302,N_2922,N_2972);
and UO_303 (O_303,N_2972,N_2971);
or UO_304 (O_304,N_2906,N_2949);
and UO_305 (O_305,N_2970,N_2973);
nor UO_306 (O_306,N_2960,N_2947);
nor UO_307 (O_307,N_2902,N_2950);
nor UO_308 (O_308,N_2910,N_2924);
and UO_309 (O_309,N_2929,N_2988);
nor UO_310 (O_310,N_2900,N_2922);
nand UO_311 (O_311,N_2951,N_2978);
or UO_312 (O_312,N_2959,N_2914);
nor UO_313 (O_313,N_2903,N_2941);
nor UO_314 (O_314,N_2988,N_2909);
xnor UO_315 (O_315,N_2908,N_2945);
or UO_316 (O_316,N_2966,N_2911);
or UO_317 (O_317,N_2953,N_2997);
or UO_318 (O_318,N_2924,N_2992);
and UO_319 (O_319,N_2966,N_2988);
nor UO_320 (O_320,N_2921,N_2989);
nor UO_321 (O_321,N_2956,N_2998);
and UO_322 (O_322,N_2907,N_2933);
or UO_323 (O_323,N_2927,N_2928);
nand UO_324 (O_324,N_2960,N_2943);
nor UO_325 (O_325,N_2964,N_2944);
or UO_326 (O_326,N_2968,N_2919);
nor UO_327 (O_327,N_2977,N_2950);
nor UO_328 (O_328,N_2962,N_2911);
and UO_329 (O_329,N_2919,N_2971);
or UO_330 (O_330,N_2940,N_2941);
and UO_331 (O_331,N_2920,N_2929);
nor UO_332 (O_332,N_2980,N_2977);
nand UO_333 (O_333,N_2917,N_2967);
xor UO_334 (O_334,N_2984,N_2921);
nand UO_335 (O_335,N_2901,N_2918);
or UO_336 (O_336,N_2947,N_2950);
or UO_337 (O_337,N_2948,N_2923);
and UO_338 (O_338,N_2994,N_2981);
or UO_339 (O_339,N_2966,N_2914);
or UO_340 (O_340,N_2974,N_2931);
xnor UO_341 (O_341,N_2977,N_2925);
nand UO_342 (O_342,N_2977,N_2906);
and UO_343 (O_343,N_2981,N_2903);
and UO_344 (O_344,N_2912,N_2944);
nand UO_345 (O_345,N_2987,N_2990);
or UO_346 (O_346,N_2943,N_2907);
and UO_347 (O_347,N_2915,N_2964);
nand UO_348 (O_348,N_2999,N_2984);
or UO_349 (O_349,N_2931,N_2902);
nor UO_350 (O_350,N_2925,N_2940);
nor UO_351 (O_351,N_2959,N_2981);
or UO_352 (O_352,N_2958,N_2928);
or UO_353 (O_353,N_2932,N_2919);
nand UO_354 (O_354,N_2990,N_2940);
nand UO_355 (O_355,N_2932,N_2999);
and UO_356 (O_356,N_2943,N_2963);
nand UO_357 (O_357,N_2974,N_2901);
and UO_358 (O_358,N_2958,N_2975);
xor UO_359 (O_359,N_2982,N_2947);
xnor UO_360 (O_360,N_2998,N_2904);
or UO_361 (O_361,N_2994,N_2909);
nor UO_362 (O_362,N_2937,N_2984);
nor UO_363 (O_363,N_2947,N_2957);
nand UO_364 (O_364,N_2905,N_2987);
nand UO_365 (O_365,N_2922,N_2988);
and UO_366 (O_366,N_2961,N_2962);
and UO_367 (O_367,N_2938,N_2977);
or UO_368 (O_368,N_2907,N_2965);
or UO_369 (O_369,N_2900,N_2918);
nand UO_370 (O_370,N_2910,N_2996);
nand UO_371 (O_371,N_2970,N_2938);
nand UO_372 (O_372,N_2976,N_2931);
or UO_373 (O_373,N_2950,N_2981);
nor UO_374 (O_374,N_2942,N_2932);
or UO_375 (O_375,N_2921,N_2988);
and UO_376 (O_376,N_2941,N_2909);
or UO_377 (O_377,N_2963,N_2900);
or UO_378 (O_378,N_2915,N_2957);
nor UO_379 (O_379,N_2922,N_2905);
nor UO_380 (O_380,N_2921,N_2918);
and UO_381 (O_381,N_2985,N_2946);
or UO_382 (O_382,N_2973,N_2985);
nor UO_383 (O_383,N_2936,N_2956);
nor UO_384 (O_384,N_2982,N_2919);
nand UO_385 (O_385,N_2951,N_2981);
nor UO_386 (O_386,N_2906,N_2975);
nor UO_387 (O_387,N_2992,N_2913);
nor UO_388 (O_388,N_2987,N_2907);
or UO_389 (O_389,N_2937,N_2904);
or UO_390 (O_390,N_2965,N_2930);
nor UO_391 (O_391,N_2997,N_2933);
or UO_392 (O_392,N_2942,N_2998);
or UO_393 (O_393,N_2992,N_2955);
or UO_394 (O_394,N_2927,N_2980);
nor UO_395 (O_395,N_2903,N_2947);
and UO_396 (O_396,N_2968,N_2993);
and UO_397 (O_397,N_2919,N_2965);
and UO_398 (O_398,N_2938,N_2974);
nor UO_399 (O_399,N_2937,N_2997);
and UO_400 (O_400,N_2927,N_2984);
and UO_401 (O_401,N_2932,N_2910);
or UO_402 (O_402,N_2918,N_2940);
xnor UO_403 (O_403,N_2993,N_2973);
or UO_404 (O_404,N_2931,N_2997);
nor UO_405 (O_405,N_2968,N_2929);
nor UO_406 (O_406,N_2904,N_2934);
nor UO_407 (O_407,N_2954,N_2952);
nand UO_408 (O_408,N_2951,N_2963);
and UO_409 (O_409,N_2915,N_2945);
nand UO_410 (O_410,N_2942,N_2939);
xor UO_411 (O_411,N_2942,N_2931);
and UO_412 (O_412,N_2923,N_2973);
and UO_413 (O_413,N_2924,N_2997);
nor UO_414 (O_414,N_2914,N_2984);
and UO_415 (O_415,N_2995,N_2919);
nand UO_416 (O_416,N_2948,N_2919);
or UO_417 (O_417,N_2982,N_2972);
or UO_418 (O_418,N_2916,N_2924);
and UO_419 (O_419,N_2915,N_2910);
and UO_420 (O_420,N_2968,N_2941);
and UO_421 (O_421,N_2932,N_2981);
nand UO_422 (O_422,N_2913,N_2917);
nor UO_423 (O_423,N_2963,N_2913);
and UO_424 (O_424,N_2999,N_2964);
or UO_425 (O_425,N_2990,N_2953);
nor UO_426 (O_426,N_2926,N_2976);
nand UO_427 (O_427,N_2972,N_2997);
nand UO_428 (O_428,N_2924,N_2903);
and UO_429 (O_429,N_2955,N_2968);
or UO_430 (O_430,N_2947,N_2934);
nand UO_431 (O_431,N_2998,N_2983);
or UO_432 (O_432,N_2928,N_2929);
or UO_433 (O_433,N_2928,N_2900);
nor UO_434 (O_434,N_2928,N_2977);
nand UO_435 (O_435,N_2940,N_2910);
xor UO_436 (O_436,N_2912,N_2943);
or UO_437 (O_437,N_2921,N_2987);
nand UO_438 (O_438,N_2945,N_2948);
nor UO_439 (O_439,N_2925,N_2906);
nand UO_440 (O_440,N_2934,N_2935);
nor UO_441 (O_441,N_2906,N_2987);
or UO_442 (O_442,N_2929,N_2916);
nor UO_443 (O_443,N_2981,N_2923);
or UO_444 (O_444,N_2908,N_2978);
or UO_445 (O_445,N_2999,N_2965);
nand UO_446 (O_446,N_2902,N_2968);
nor UO_447 (O_447,N_2960,N_2921);
and UO_448 (O_448,N_2954,N_2935);
nor UO_449 (O_449,N_2906,N_2997);
nand UO_450 (O_450,N_2966,N_2971);
nor UO_451 (O_451,N_2949,N_2941);
nand UO_452 (O_452,N_2904,N_2975);
nand UO_453 (O_453,N_2919,N_2911);
or UO_454 (O_454,N_2900,N_2956);
nand UO_455 (O_455,N_2966,N_2959);
nor UO_456 (O_456,N_2975,N_2929);
xnor UO_457 (O_457,N_2909,N_2900);
and UO_458 (O_458,N_2968,N_2900);
or UO_459 (O_459,N_2945,N_2972);
or UO_460 (O_460,N_2976,N_2973);
nand UO_461 (O_461,N_2920,N_2919);
nand UO_462 (O_462,N_2979,N_2996);
nand UO_463 (O_463,N_2925,N_2996);
nor UO_464 (O_464,N_2984,N_2916);
xor UO_465 (O_465,N_2939,N_2931);
nor UO_466 (O_466,N_2921,N_2931);
nand UO_467 (O_467,N_2986,N_2974);
nor UO_468 (O_468,N_2945,N_2977);
nand UO_469 (O_469,N_2928,N_2916);
nand UO_470 (O_470,N_2944,N_2992);
nand UO_471 (O_471,N_2904,N_2992);
nand UO_472 (O_472,N_2922,N_2950);
nor UO_473 (O_473,N_2928,N_2956);
and UO_474 (O_474,N_2930,N_2961);
and UO_475 (O_475,N_2944,N_2990);
or UO_476 (O_476,N_2933,N_2993);
and UO_477 (O_477,N_2951,N_2945);
xor UO_478 (O_478,N_2998,N_2966);
or UO_479 (O_479,N_2991,N_2938);
xor UO_480 (O_480,N_2945,N_2914);
nor UO_481 (O_481,N_2915,N_2968);
or UO_482 (O_482,N_2941,N_2994);
nand UO_483 (O_483,N_2982,N_2960);
nand UO_484 (O_484,N_2948,N_2927);
nor UO_485 (O_485,N_2923,N_2953);
nand UO_486 (O_486,N_2900,N_2988);
nor UO_487 (O_487,N_2951,N_2911);
nor UO_488 (O_488,N_2908,N_2974);
and UO_489 (O_489,N_2940,N_2936);
and UO_490 (O_490,N_2975,N_2997);
or UO_491 (O_491,N_2944,N_2969);
or UO_492 (O_492,N_2954,N_2920);
nand UO_493 (O_493,N_2996,N_2954);
xnor UO_494 (O_494,N_2911,N_2956);
nor UO_495 (O_495,N_2981,N_2983);
nor UO_496 (O_496,N_2930,N_2974);
nor UO_497 (O_497,N_2986,N_2931);
nand UO_498 (O_498,N_2945,N_2901);
nor UO_499 (O_499,N_2980,N_2936);
endmodule