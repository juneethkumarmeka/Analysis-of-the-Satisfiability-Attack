module basic_2500_25000_3000_100_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
and U0 (N_0,In_580,In_1424);
nand U1 (N_1,In_1231,In_1940);
nor U2 (N_2,In_1551,In_1625);
or U3 (N_3,In_248,In_457);
or U4 (N_4,In_200,In_286);
nand U5 (N_5,In_682,In_1018);
and U6 (N_6,In_741,In_98);
and U7 (N_7,In_61,In_65);
or U8 (N_8,In_331,In_19);
nand U9 (N_9,In_1339,In_298);
or U10 (N_10,In_823,In_781);
nor U11 (N_11,In_1246,In_1948);
and U12 (N_12,In_58,In_564);
xnor U13 (N_13,In_41,In_118);
nor U14 (N_14,In_1730,In_579);
nor U15 (N_15,In_1875,In_1089);
and U16 (N_16,In_538,In_0);
nand U17 (N_17,In_738,In_1974);
and U18 (N_18,In_2498,In_1902);
and U19 (N_19,In_1545,In_503);
nor U20 (N_20,In_2289,In_384);
nand U21 (N_21,In_2244,In_2127);
nor U22 (N_22,In_971,In_2496);
and U23 (N_23,In_991,In_84);
or U24 (N_24,In_951,In_1238);
and U25 (N_25,In_2386,In_1316);
or U26 (N_26,In_1618,In_1623);
and U27 (N_27,In_1282,In_835);
or U28 (N_28,In_2248,In_2427);
nor U29 (N_29,In_2382,In_1372);
and U30 (N_30,In_428,In_1607);
xnor U31 (N_31,In_1472,In_2217);
or U32 (N_32,In_2345,In_1756);
nor U33 (N_33,In_1589,In_2195);
nand U34 (N_34,In_2161,In_1490);
nor U35 (N_35,In_476,In_1999);
and U36 (N_36,In_2369,In_2006);
and U37 (N_37,In_802,In_1679);
or U38 (N_38,In_2179,In_2495);
or U39 (N_39,In_917,In_1991);
nand U40 (N_40,In_1990,In_397);
or U41 (N_41,In_48,In_825);
nand U42 (N_42,In_661,In_861);
nor U43 (N_43,In_2075,In_1924);
nor U44 (N_44,In_488,In_1746);
nor U45 (N_45,In_841,In_1301);
nand U46 (N_46,In_973,In_2461);
nand U47 (N_47,In_2485,In_344);
and U48 (N_48,In_96,In_1349);
and U49 (N_49,In_153,In_1907);
and U50 (N_50,In_1156,In_309);
xnor U51 (N_51,In_2199,In_2231);
nand U52 (N_52,In_2104,In_24);
nor U53 (N_53,In_1776,In_2259);
nor U54 (N_54,In_2260,In_2170);
nor U55 (N_55,In_7,In_458);
nand U56 (N_56,In_1021,In_856);
nor U57 (N_57,In_750,In_2061);
or U58 (N_58,In_1159,In_1785);
or U59 (N_59,In_585,In_2058);
or U60 (N_60,In_1494,In_2304);
nor U61 (N_61,In_1193,In_1540);
and U62 (N_62,In_1788,In_95);
or U63 (N_63,In_2144,In_591);
or U64 (N_64,In_43,In_27);
or U65 (N_65,In_2204,In_1058);
and U66 (N_66,In_1187,In_1103);
xor U67 (N_67,In_2100,In_1641);
and U68 (N_68,In_928,In_2401);
nand U69 (N_69,In_1614,In_1538);
nor U70 (N_70,In_132,In_401);
or U71 (N_71,In_968,In_1227);
and U72 (N_72,In_370,In_1181);
and U73 (N_73,In_848,In_2022);
or U74 (N_74,In_1520,In_1169);
or U75 (N_75,In_2439,In_649);
nand U76 (N_76,In_2245,In_2354);
xor U77 (N_77,In_1405,In_2014);
xor U78 (N_78,In_1844,In_2065);
nand U79 (N_79,In_1460,In_2145);
and U80 (N_80,In_867,In_716);
nand U81 (N_81,In_2008,In_654);
and U82 (N_82,In_2380,In_2157);
nor U83 (N_83,In_226,In_1505);
and U84 (N_84,In_616,In_385);
nand U85 (N_85,In_2407,In_1119);
nand U86 (N_86,In_313,In_2239);
and U87 (N_87,In_358,In_1558);
or U88 (N_88,In_1039,In_921);
nor U89 (N_89,In_2379,In_1210);
nand U90 (N_90,In_1543,In_77);
or U91 (N_91,In_1951,In_1737);
nor U92 (N_92,In_337,In_1218);
nor U93 (N_93,In_705,In_28);
and U94 (N_94,In_587,In_668);
and U95 (N_95,In_2436,In_1661);
or U96 (N_96,In_2007,In_2385);
nor U97 (N_97,In_1222,In_1113);
nor U98 (N_98,In_1828,In_1565);
and U99 (N_99,In_1692,In_149);
and U100 (N_100,In_1886,In_1431);
or U101 (N_101,In_253,In_1098);
nor U102 (N_102,In_1985,In_2060);
nand U103 (N_103,In_1393,In_2394);
and U104 (N_104,In_296,In_757);
nand U105 (N_105,In_441,In_1344);
or U106 (N_106,In_1161,In_1324);
or U107 (N_107,In_552,In_2049);
nand U108 (N_108,In_1586,In_708);
nand U109 (N_109,In_605,In_1237);
and U110 (N_110,In_1590,In_1584);
nand U111 (N_111,In_355,In_1603);
or U112 (N_112,In_1763,In_1779);
nor U113 (N_113,In_1022,In_1175);
and U114 (N_114,In_2112,In_285);
nor U115 (N_115,In_1033,In_448);
nand U116 (N_116,In_123,In_536);
and U117 (N_117,In_411,In_2435);
nand U118 (N_118,In_1622,In_287);
xnor U119 (N_119,In_1030,In_931);
nand U120 (N_120,In_1445,In_1698);
nor U121 (N_121,In_188,In_1228);
and U122 (N_122,In_364,In_1583);
and U123 (N_123,In_1394,In_2428);
and U124 (N_124,In_162,In_2201);
nor U125 (N_125,In_104,In_1579);
nand U126 (N_126,In_1760,In_134);
and U127 (N_127,In_1125,In_2335);
xnor U128 (N_128,In_889,In_395);
nand U129 (N_129,In_1307,In_810);
nor U130 (N_130,In_2465,In_2238);
and U131 (N_131,In_1845,In_1473);
nand U132 (N_132,In_1167,In_115);
or U133 (N_133,In_246,In_466);
or U134 (N_134,In_2307,In_81);
nand U135 (N_135,In_452,In_790);
and U136 (N_136,In_1765,In_643);
nand U137 (N_137,In_2291,In_229);
nand U138 (N_138,In_1462,In_1678);
or U139 (N_139,In_2082,In_1670);
nand U140 (N_140,In_2448,In_2137);
or U141 (N_141,In_187,In_450);
nor U142 (N_142,In_2039,In_1997);
nand U143 (N_143,In_1983,In_2357);
nand U144 (N_144,In_111,In_1609);
nand U145 (N_145,In_596,In_1850);
or U146 (N_146,In_1702,In_256);
and U147 (N_147,In_2109,In_1501);
and U148 (N_148,In_1384,In_1176);
and U149 (N_149,In_2175,In_851);
nand U150 (N_150,In_2298,In_473);
or U151 (N_151,In_812,In_2301);
nor U152 (N_152,In_879,In_2055);
or U153 (N_153,In_2486,In_1006);
or U154 (N_154,In_237,In_912);
and U155 (N_155,In_853,In_71);
or U156 (N_156,In_1489,In_2117);
and U157 (N_157,In_1696,In_1793);
nor U158 (N_158,In_718,In_1455);
or U159 (N_159,In_2440,In_33);
or U160 (N_160,In_1743,In_927);
nor U161 (N_161,In_1832,In_547);
nand U162 (N_162,In_2377,In_1596);
or U163 (N_163,In_255,In_2225);
or U164 (N_164,In_947,In_732);
nor U165 (N_165,In_194,In_1686);
and U166 (N_166,In_1736,In_534);
nand U167 (N_167,In_1152,In_1560);
and U168 (N_168,In_2292,In_1637);
and U169 (N_169,In_1754,In_1352);
nand U170 (N_170,In_1153,In_988);
nor U171 (N_171,In_1725,In_813);
xnor U172 (N_172,In_1977,In_1268);
nor U173 (N_173,In_1166,In_1525);
or U174 (N_174,In_1087,In_622);
and U175 (N_175,In_1710,In_799);
and U176 (N_176,In_593,In_292);
or U177 (N_177,In_295,In_1220);
nor U178 (N_178,In_1370,In_495);
and U179 (N_179,In_1003,In_2091);
and U180 (N_180,In_873,In_2000);
or U181 (N_181,In_811,In_1254);
or U182 (N_182,In_82,In_902);
xor U183 (N_183,In_2420,In_443);
or U184 (N_184,In_883,In_939);
xor U185 (N_185,In_352,In_1711);
nand U186 (N_186,In_1441,In_1972);
xnor U187 (N_187,In_224,In_1256);
and U188 (N_188,In_975,In_502);
and U189 (N_189,In_1477,In_576);
nand U190 (N_190,In_1331,In_474);
and U191 (N_191,In_2419,In_254);
nor U192 (N_192,In_94,In_239);
or U193 (N_193,In_1910,In_1595);
or U194 (N_194,In_878,In_1036);
nand U195 (N_195,In_1482,In_2094);
xor U196 (N_196,In_858,In_2499);
nand U197 (N_197,In_2315,In_2153);
xnor U198 (N_198,In_1364,In_1880);
nor U199 (N_199,In_276,In_1293);
and U200 (N_200,In_1134,In_1248);
xnor U201 (N_201,In_2410,In_1873);
or U202 (N_202,In_624,In_1470);
and U203 (N_203,In_2024,In_1052);
and U204 (N_204,In_335,In_2140);
nand U205 (N_205,In_2336,In_1688);
xor U206 (N_206,In_2371,In_1687);
or U207 (N_207,In_1149,In_343);
nand U208 (N_208,In_266,In_14);
or U209 (N_209,In_1044,In_877);
nand U210 (N_210,In_53,In_294);
or U211 (N_211,In_2167,In_744);
and U212 (N_212,In_1762,In_173);
nand U213 (N_213,In_1734,In_1797);
and U214 (N_214,In_1911,In_1196);
and U215 (N_215,In_293,In_2430);
nor U216 (N_216,In_809,In_1487);
nor U217 (N_217,In_2185,In_1009);
nand U218 (N_218,In_409,In_332);
or U219 (N_219,In_6,In_120);
nand U220 (N_220,In_1106,In_1396);
nand U221 (N_221,In_854,In_1613);
and U222 (N_222,In_1913,In_2158);
or U223 (N_223,In_2093,In_1615);
nand U224 (N_224,In_602,In_481);
nor U225 (N_225,In_201,In_1608);
xnor U226 (N_226,In_2230,In_197);
nand U227 (N_227,In_866,In_2413);
and U228 (N_228,In_1047,In_2176);
and U229 (N_229,In_2032,In_914);
nor U230 (N_230,In_993,In_566);
and U231 (N_231,In_489,In_1904);
and U232 (N_232,In_946,In_1480);
nand U233 (N_233,In_1000,In_376);
and U234 (N_234,In_388,In_1707);
xnor U235 (N_235,In_1390,In_1981);
or U236 (N_236,In_1385,In_2090);
or U237 (N_237,In_2222,In_2476);
and U238 (N_238,In_1013,In_1336);
nor U239 (N_239,In_637,In_2051);
or U240 (N_240,In_1067,In_264);
xor U241 (N_241,In_766,In_156);
xor U242 (N_242,In_2142,In_1280);
or U243 (N_243,In_594,In_2202);
xor U244 (N_244,In_1712,In_1038);
and U245 (N_245,In_392,In_2274);
nand U246 (N_246,In_2253,In_311);
and U247 (N_247,In_1059,In_1406);
and U248 (N_248,In_1323,In_2279);
and U249 (N_249,In_653,In_898);
nand U250 (N_250,In_350,In_203);
and U251 (N_251,In_2156,In_628);
nor U252 (N_252,In_754,In_2460);
or U253 (N_253,In_970,In_673);
nand U254 (N_254,In_2453,In_671);
or U255 (N_255,In_1750,In_2290);
and U256 (N_256,In_2205,In_421);
nor U257 (N_257,In_496,In_1150);
nor U258 (N_258,In_597,N_10);
xor U259 (N_259,In_839,In_2360);
nor U260 (N_260,In_1082,N_115);
and U261 (N_261,In_1899,In_122);
nand U262 (N_262,N_23,In_1708);
and U263 (N_263,N_114,In_2009);
nor U264 (N_264,In_789,In_692);
nand U265 (N_265,In_2387,N_138);
and U266 (N_266,In_273,In_956);
nor U267 (N_267,In_1439,N_57);
or U268 (N_268,N_1,In_1831);
nor U269 (N_269,In_208,N_139);
xnor U270 (N_270,In_570,In_507);
and U271 (N_271,In_1314,In_357);
or U272 (N_272,In_189,In_948);
or U273 (N_273,In_23,N_120);
xor U274 (N_274,In_1140,N_7);
and U275 (N_275,N_34,In_107);
or U276 (N_276,In_913,In_2002);
or U277 (N_277,In_306,In_1954);
or U278 (N_278,In_1935,In_2418);
nand U279 (N_279,In_1715,In_1141);
nor U280 (N_280,In_918,In_190);
nor U281 (N_281,N_148,In_1056);
or U282 (N_282,In_2267,In_483);
nor U283 (N_283,In_1459,In_1582);
nor U284 (N_284,In_911,In_967);
nand U285 (N_285,In_1345,In_1533);
or U286 (N_286,In_1656,In_2297);
or U287 (N_287,In_903,In_2442);
nor U288 (N_288,In_1027,In_261);
or U289 (N_289,In_1341,In_1635);
and U290 (N_290,In_1279,In_920);
nor U291 (N_291,In_2406,In_1570);
nand U292 (N_292,In_1124,In_847);
nand U293 (N_293,In_26,In_961);
nor U294 (N_294,In_2316,In_1160);
nand U295 (N_295,In_1937,In_2042);
and U296 (N_296,In_1350,In_2263);
nand U297 (N_297,In_1436,In_1217);
and U298 (N_298,In_1475,In_1251);
or U299 (N_299,In_2188,In_2057);
nor U300 (N_300,In_1457,In_1856);
and U301 (N_301,In_130,In_815);
and U302 (N_302,In_1214,N_112);
and U303 (N_303,In_1509,In_862);
and U304 (N_304,In_2240,In_479);
nor U305 (N_305,In_1205,In_513);
xnor U306 (N_306,In_2062,In_2318);
xnor U307 (N_307,In_1898,In_859);
xnor U308 (N_308,In_685,In_734);
nand U309 (N_309,In_2079,In_195);
nor U310 (N_310,In_985,In_758);
or U311 (N_311,In_2071,In_636);
nor U312 (N_312,In_307,In_1008);
or U313 (N_313,In_2050,In_437);
nor U314 (N_314,N_171,In_833);
nand U315 (N_315,N_64,In_179);
nand U316 (N_316,N_54,In_1534);
nor U317 (N_317,In_2101,N_158);
xor U318 (N_318,In_1334,In_1592);
nor U319 (N_319,In_2027,In_1877);
or U320 (N_320,In_1162,In_1742);
nand U321 (N_321,N_63,In_663);
xnor U322 (N_322,In_586,In_2005);
or U323 (N_323,In_680,In_1236);
nand U324 (N_324,In_1518,In_1893);
or U325 (N_325,In_157,In_1781);
and U326 (N_326,In_535,In_1049);
xor U327 (N_327,In_509,In_1452);
or U328 (N_328,In_537,In_2069);
xor U329 (N_329,In_124,In_804);
nor U330 (N_330,In_1878,In_405);
nand U331 (N_331,In_962,In_740);
or U332 (N_332,In_1870,In_1857);
nor U333 (N_333,In_1195,In_35);
xor U334 (N_334,In_1662,In_2192);
xnor U335 (N_335,In_1598,In_1631);
xor U336 (N_336,In_291,In_2469);
nand U337 (N_337,In_2034,In_1933);
nor U338 (N_338,In_339,In_2452);
nor U339 (N_339,In_792,N_22);
or U340 (N_340,In_589,In_780);
or U341 (N_341,In_976,In_1519);
or U342 (N_342,In_731,In_213);
nor U343 (N_343,N_164,In_822);
or U344 (N_344,In_1397,In_2472);
nor U345 (N_345,In_2012,In_2228);
or U346 (N_346,In_613,In_152);
xor U347 (N_347,In_752,In_1239);
and U348 (N_348,N_122,In_234);
nor U349 (N_349,In_1611,In_445);
or U350 (N_350,In_2356,In_1325);
nor U351 (N_351,In_413,In_66);
or U352 (N_352,In_1034,In_391);
nand U353 (N_353,In_1814,In_2344);
nor U354 (N_354,N_107,N_73);
and U355 (N_355,In_1665,In_268);
nor U356 (N_356,In_145,In_1638);
nor U357 (N_357,In_1772,In_222);
nor U358 (N_358,In_1121,In_583);
xor U359 (N_359,In_1953,In_2132);
or U360 (N_360,N_147,N_8);
nand U361 (N_361,In_371,In_315);
nor U362 (N_362,In_1650,In_1966);
nand U363 (N_363,In_349,In_1945);
nor U364 (N_364,In_1155,In_1199);
nand U365 (N_365,In_241,In_2294);
or U366 (N_366,In_341,In_714);
nand U367 (N_367,In_706,In_1759);
nand U368 (N_368,N_30,In_10);
and U369 (N_369,In_2484,In_1848);
or U370 (N_370,In_876,In_1961);
or U371 (N_371,N_103,In_1079);
nand U372 (N_372,In_733,In_1269);
and U373 (N_373,In_2374,In_2128);
nand U374 (N_374,In_522,In_1724);
and U375 (N_375,In_178,In_2334);
nor U376 (N_376,In_1054,In_270);
or U377 (N_377,In_803,In_8);
or U378 (N_378,In_746,In_161);
or U379 (N_379,In_1758,In_461);
nor U380 (N_380,In_475,In_1895);
nand U381 (N_381,In_484,N_155);
nand U382 (N_382,In_2246,In_1517);
and U383 (N_383,In_888,In_2445);
xor U384 (N_384,N_60,N_104);
nor U385 (N_385,In_2402,In_1621);
and U386 (N_386,In_272,In_2467);
nand U387 (N_387,In_762,In_1354);
xor U388 (N_388,In_1819,In_1949);
and U389 (N_389,In_1495,In_303);
and U390 (N_390,In_737,In_2323);
xnor U391 (N_391,In_342,In_1398);
nand U392 (N_392,In_723,In_1243);
nor U393 (N_393,N_146,In_160);
nor U394 (N_394,In_891,In_1726);
or U395 (N_395,In_818,In_957);
nor U396 (N_396,N_191,In_1430);
and U397 (N_397,In_1073,In_1387);
xnor U398 (N_398,In_543,In_742);
nor U399 (N_399,In_216,In_1469);
and U400 (N_400,In_1854,In_1629);
or U401 (N_401,In_1440,In_717);
and U402 (N_402,In_1453,In_2256);
nand U403 (N_403,N_127,N_32);
and U404 (N_404,In_2431,In_722);
nand U405 (N_405,In_2362,In_715);
and U406 (N_406,In_1813,In_105);
nand U407 (N_407,In_1820,In_516);
xnor U408 (N_408,In_683,In_1492);
nor U409 (N_409,In_2198,In_545);
nor U410 (N_410,N_224,In_1926);
xor U411 (N_411,In_2031,In_1908);
nand U412 (N_412,In_2415,In_2481);
and U413 (N_413,In_699,In_1465);
nor U414 (N_414,In_926,In_184);
or U415 (N_415,In_1729,N_80);
or U416 (N_416,In_989,In_2092);
and U417 (N_417,In_568,In_1105);
or U418 (N_418,In_1174,In_166);
nor U419 (N_419,In_1980,In_625);
or U420 (N_420,In_147,In_319);
nand U421 (N_421,N_44,In_1065);
nand U422 (N_422,In_638,In_978);
and U423 (N_423,In_1332,In_2479);
xnor U424 (N_424,N_38,In_765);
nor U425 (N_425,In_1839,In_1179);
or U426 (N_426,In_1225,In_1836);
xnor U427 (N_427,In_2025,In_1806);
or U428 (N_428,In_1941,In_381);
nand U429 (N_429,In_2028,In_1956);
or U430 (N_430,In_1164,In_174);
or U431 (N_431,N_237,In_1567);
nand U432 (N_432,In_1017,In_1932);
nand U433 (N_433,In_1978,In_1510);
or U434 (N_434,In_333,In_2073);
and U435 (N_435,In_2309,In_56);
and U436 (N_436,In_2126,N_163);
or U437 (N_437,In_1516,In_2019);
nor U438 (N_438,In_1840,In_1508);
nor U439 (N_439,In_396,In_986);
and U440 (N_440,In_1348,In_1437);
and U441 (N_441,In_389,In_592);
or U442 (N_442,In_1011,In_1226);
nor U443 (N_443,N_100,In_1186);
nand U444 (N_444,In_2338,In_100);
and U445 (N_445,In_1433,In_69);
or U446 (N_446,In_80,N_233);
nor U447 (N_447,In_2133,In_460);
or U448 (N_448,In_595,In_1401);
nand U449 (N_449,In_2416,In_497);
nand U450 (N_450,In_1992,In_2);
and U451 (N_451,In_182,In_399);
and U452 (N_452,In_710,In_642);
nor U453 (N_453,In_2317,In_372);
or U454 (N_454,In_531,N_31);
nor U455 (N_455,N_137,In_1604);
and U456 (N_456,In_1443,In_1203);
nand U457 (N_457,In_2348,N_216);
and U458 (N_458,In_2138,N_12);
nand U459 (N_459,In_2373,In_1561);
nor U460 (N_460,In_567,In_665);
nand U461 (N_461,N_25,In_219);
nor U462 (N_462,In_487,In_1064);
nand U463 (N_463,In_359,N_96);
nor U464 (N_464,N_149,In_1694);
nand U465 (N_465,In_632,In_2363);
or U466 (N_466,In_2313,In_794);
nand U467 (N_467,In_1311,In_1241);
nand U468 (N_468,In_1346,In_459);
and U469 (N_469,In_1102,In_2310);
xor U470 (N_470,In_1136,In_1532);
or U471 (N_471,In_1588,In_932);
or U472 (N_472,In_90,In_2166);
and U473 (N_473,In_674,In_560);
or U474 (N_474,In_1157,In_265);
nand U475 (N_475,In_1807,In_1964);
or U476 (N_476,N_231,In_453);
nor U477 (N_477,In_1467,In_1309);
nand U478 (N_478,In_944,N_174);
xnor U479 (N_479,In_2067,In_1865);
and U480 (N_480,In_1996,In_2261);
and U481 (N_481,In_361,In_631);
and U482 (N_482,In_617,In_2319);
and U483 (N_483,In_852,In_1984);
nor U484 (N_484,In_288,In_1019);
nand U485 (N_485,In_751,In_1326);
nand U486 (N_486,In_916,N_116);
nor U487 (N_487,In_2221,In_1817);
or U488 (N_488,N_21,N_33);
and U489 (N_489,In_1802,In_832);
nand U490 (N_490,In_1675,In_212);
or U491 (N_491,In_377,In_2129);
xor U492 (N_492,In_1804,N_186);
nand U493 (N_493,In_1014,In_2236);
and U494 (N_494,N_156,In_1053);
nand U495 (N_495,In_155,In_351);
nand U496 (N_496,In_1496,In_704);
or U497 (N_497,In_582,In_806);
or U498 (N_498,In_930,In_561);
nor U499 (N_499,In_1207,In_2054);
or U500 (N_500,In_1329,N_355);
and U501 (N_501,N_212,In_1969);
nand U502 (N_502,In_2337,In_1288);
and U503 (N_503,In_2141,In_753);
and U504 (N_504,In_2123,In_1846);
and U505 (N_505,In_2257,In_1605);
or U506 (N_506,In_941,In_1795);
nor U507 (N_507,In_1805,In_2155);
or U508 (N_508,In_1177,N_235);
and U509 (N_509,In_1782,N_254);
nand U510 (N_510,In_1550,In_669);
and U511 (N_511,N_20,In_656);
nand U512 (N_512,In_1328,In_934);
nor U513 (N_513,In_1417,In_689);
nor U514 (N_514,N_272,N_89);
or U515 (N_515,In_1537,In_429);
and U516 (N_516,N_129,In_398);
nand U517 (N_517,In_1620,In_1273);
nand U518 (N_518,In_1915,N_273);
nand U519 (N_519,In_2471,In_1420);
or U520 (N_520,N_496,In_1194);
xnor U521 (N_521,N_318,N_194);
nor U522 (N_522,In_1330,In_652);
and U523 (N_523,In_698,N_181);
and U524 (N_524,In_1697,In_2178);
nor U525 (N_525,In_2455,In_1610);
nor U526 (N_526,In_1407,In_553);
xor U527 (N_527,In_1291,In_1094);
nand U528 (N_528,N_202,In_204);
xor U529 (N_529,In_937,In_1816);
or U530 (N_530,N_183,In_635);
nand U531 (N_531,N_342,In_2449);
nand U532 (N_532,In_2020,In_778);
nand U533 (N_533,N_67,In_1653);
xnor U534 (N_534,In_735,In_910);
or U535 (N_535,In_2023,In_782);
nand U536 (N_536,In_958,In_112);
nand U537 (N_537,In_805,N_327);
xor U538 (N_538,In_2306,In_284);
nor U539 (N_539,In_992,N_404);
and U540 (N_540,In_963,N_372);
nor U541 (N_541,In_1552,In_837);
nor U542 (N_542,In_1823,In_4);
nor U543 (N_543,In_842,In_64);
or U544 (N_544,In_2001,In_1357);
and U545 (N_545,N_281,In_1619);
nor U546 (N_546,In_630,In_1863);
nor U547 (N_547,N_471,N_482);
nand U548 (N_548,In_380,In_2483);
and U549 (N_549,In_1626,N_215);
or U550 (N_550,N_354,In_1403);
or U551 (N_551,In_695,In_982);
nand U552 (N_552,In_2432,In_907);
or U553 (N_553,In_1914,In_1666);
or U554 (N_554,In_55,In_2326);
nand U555 (N_555,N_132,In_260);
nor U556 (N_556,In_1204,In_2349);
nand U557 (N_557,N_15,In_1110);
or U558 (N_558,N_374,In_419);
and U559 (N_559,In_60,In_365);
nand U560 (N_560,N_265,In_1716);
or U561 (N_561,In_1982,N_141);
nor U562 (N_562,In_21,In_2229);
and U563 (N_563,N_467,In_231);
or U564 (N_564,In_1645,N_108);
or U565 (N_565,N_317,In_882);
and U566 (N_566,In_1135,In_2096);
and U567 (N_567,In_2045,In_2311);
nand U568 (N_568,In_687,In_1444);
and U569 (N_569,N_14,In_1809);
nor U570 (N_570,In_2412,In_1025);
nand U571 (N_571,In_1450,In_2266);
nand U572 (N_572,N_401,In_1960);
or U573 (N_573,In_972,In_2392);
and U574 (N_574,N_257,N_406);
nor U575 (N_575,In_79,In_1731);
nor U576 (N_576,In_1827,N_213);
nor U577 (N_577,In_2235,N_192);
and U578 (N_578,In_2036,N_227);
nor U579 (N_579,In_1513,In_954);
and U580 (N_580,In_1422,In_1695);
nor U581 (N_581,In_1970,In_896);
nand U582 (N_582,In_514,In_1659);
nand U583 (N_583,In_1100,In_1245);
and U584 (N_584,In_830,N_362);
or U585 (N_585,In_238,In_1667);
or U586 (N_586,In_1182,In_375);
nand U587 (N_587,In_834,In_1642);
nor U588 (N_588,In_1868,In_2254);
nand U589 (N_589,In_1930,In_1060);
and U590 (N_590,In_1147,In_1032);
xor U591 (N_591,In_91,In_322);
and U592 (N_592,N_479,N_296);
or U593 (N_593,In_2115,In_1818);
or U594 (N_594,In_2441,In_2283);
nor U595 (N_595,In_244,In_38);
nand U596 (N_596,In_2491,In_2237);
and U597 (N_597,In_301,N_306);
nor U598 (N_598,In_78,N_415);
or U599 (N_599,N_266,In_1080);
nor U600 (N_600,In_1029,In_578);
xnor U601 (N_601,In_1847,In_1287);
and U602 (N_602,N_370,In_89);
xor U603 (N_603,In_1931,In_2321);
xor U604 (N_604,N_199,N_200);
nand U605 (N_605,In_528,In_76);
or U606 (N_606,In_282,N_83);
nand U607 (N_607,In_1471,In_346);
nand U608 (N_608,In_1685,In_230);
nor U609 (N_609,In_1306,N_161);
nand U610 (N_610,In_1950,N_140);
and U611 (N_611,In_2210,In_434);
and U612 (N_612,In_517,In_1178);
and U613 (N_613,In_1936,N_459);
or U614 (N_614,In_964,In_324);
and U615 (N_615,In_2194,In_1713);
nor U616 (N_616,In_641,N_309);
xnor U617 (N_617,In_1419,N_388);
nand U618 (N_618,In_1976,In_1024);
and U619 (N_619,In_759,In_170);
and U620 (N_620,In_2056,In_666);
xnor U621 (N_621,In_1593,In_1906);
xnor U622 (N_622,In_1201,In_997);
nor U623 (N_623,N_135,In_1284);
and U624 (N_624,In_467,N_383);
or U625 (N_625,N_70,In_1770);
or U626 (N_626,N_144,In_205);
or U627 (N_627,In_1689,N_275);
nand U628 (N_628,In_1378,N_326);
or U629 (N_629,In_44,N_377);
or U630 (N_630,In_506,In_320);
and U631 (N_631,In_1066,In_1297);
nor U632 (N_632,N_430,In_196);
or U633 (N_633,In_2068,In_1252);
nand U634 (N_634,In_31,In_1800);
xnor U635 (N_635,N_62,N_313);
nor U636 (N_636,In_713,In_1229);
nand U637 (N_637,In_1247,In_729);
nor U638 (N_638,In_225,N_214);
or U639 (N_639,In_369,In_1521);
nor U640 (N_640,In_2186,In_829);
nor U641 (N_641,N_105,In_1646);
nand U642 (N_642,In_1481,In_672);
nor U643 (N_643,In_2102,In_1223);
and U644 (N_644,In_562,In_1085);
or U645 (N_645,In_183,In_621);
and U646 (N_646,In_119,In_485);
nand U647 (N_647,In_432,N_259);
or U648 (N_648,In_1312,N_86);
and U649 (N_649,In_240,In_1627);
nor U650 (N_650,N_491,In_2376);
xor U651 (N_651,N_95,In_16);
nand U652 (N_652,In_185,In_2272);
xnor U653 (N_653,In_378,In_70);
and U654 (N_654,In_1581,In_1253);
nand U655 (N_655,N_268,In_305);
nand U656 (N_656,In_1771,In_646);
and U657 (N_657,In_1173,In_2242);
nand U658 (N_658,N_375,In_739);
and U659 (N_659,In_1946,In_1794);
or U660 (N_660,N_416,N_448);
nor U661 (N_661,In_2275,In_1617);
nand U662 (N_662,In_1512,N_428);
or U663 (N_663,N_270,In_68);
nand U664 (N_664,In_1356,N_263);
or U665 (N_665,In_1084,In_2293);
or U666 (N_666,In_39,In_1568);
nand U667 (N_667,In_1628,N_97);
xor U668 (N_668,In_508,N_405);
nand U669 (N_669,N_50,N_466);
or U670 (N_670,In_1365,In_1057);
nand U671 (N_671,In_1074,In_435);
or U672 (N_672,In_849,In_1528);
and U673 (N_673,In_1108,In_186);
nand U674 (N_674,In_2043,In_233);
nor U675 (N_675,In_1359,In_1644);
and U676 (N_676,In_797,N_42);
nor U677 (N_677,N_450,N_285);
and U678 (N_678,In_1995,In_1342);
and U679 (N_679,In_1647,In_348);
nor U680 (N_680,N_204,In_1305);
or U681 (N_681,In_2081,In_2097);
nand U682 (N_682,In_2383,In_855);
nand U683 (N_683,In_950,In_942);
and U684 (N_684,In_2414,In_463);
nand U685 (N_685,N_456,In_3);
nand U686 (N_686,In_639,N_299);
nor U687 (N_687,In_180,In_2164);
nand U688 (N_688,In_312,In_110);
nor U689 (N_689,In_1606,In_422);
or U690 (N_690,In_336,In_258);
nor U691 (N_691,In_252,In_1078);
or U692 (N_692,In_2473,In_2220);
xnor U693 (N_693,In_681,In_1144);
or U694 (N_694,N_367,In_2087);
nand U695 (N_695,In_1677,In_1703);
or U696 (N_696,In_607,In_277);
or U697 (N_697,In_721,In_1993);
nor U698 (N_698,In_1088,N_488);
nor U699 (N_699,In_1979,N_180);
nor U700 (N_700,In_1298,In_2152);
nand U701 (N_701,In_1574,In_2351);
nor U702 (N_702,In_2403,In_1884);
nand U703 (N_703,N_451,N_59);
and U704 (N_704,In_1504,In_1751);
nor U705 (N_705,In_1004,In_1529);
and U706 (N_706,In_1881,In_1752);
nand U707 (N_707,In_1843,In_191);
xor U708 (N_708,In_1916,In_109);
xor U709 (N_709,In_959,N_99);
nand U710 (N_710,In_1885,In_657);
nor U711 (N_711,In_555,In_577);
and U712 (N_712,In_1154,In_99);
xnor U713 (N_713,In_965,N_350);
and U714 (N_714,In_1923,In_278);
nand U715 (N_715,In_325,In_1723);
xnor U716 (N_716,In_1261,N_111);
nand U717 (N_717,In_2411,In_1585);
or U718 (N_718,In_1304,In_2322);
or U719 (N_719,N_175,In_990);
or U720 (N_720,In_2111,N_480);
or U721 (N_721,In_2187,In_321);
xnor U722 (N_722,N_439,In_2346);
nor U723 (N_723,N_201,In_1859);
and U724 (N_724,In_1310,In_259);
or U725 (N_725,In_2191,In_1043);
or U726 (N_726,In_727,In_1429);
nand U727 (N_727,N_475,In_1943);
nand U728 (N_728,In_2295,N_423);
xor U729 (N_729,In_798,In_556);
nor U730 (N_730,In_915,N_101);
and U731 (N_731,N_391,In_1037);
or U732 (N_732,In_29,In_374);
or U733 (N_733,In_1163,N_356);
xnor U734 (N_734,In_345,In_1200);
or U735 (N_735,In_1571,In_1815);
nor U736 (N_736,In_2287,In_2116);
and U737 (N_737,N_499,In_1171);
nor U738 (N_738,N_392,In_2433);
nand U739 (N_739,In_2262,In_774);
nor U740 (N_740,In_1657,N_128);
nand U741 (N_741,In_360,In_843);
and U742 (N_742,In_2330,In_2277);
nor U743 (N_743,In_2180,In_1673);
and U744 (N_744,N_81,In_1929);
nand U745 (N_745,In_13,In_2331);
and U746 (N_746,In_1668,In_999);
xor U747 (N_747,In_1001,N_193);
nand U748 (N_748,In_144,In_511);
nor U749 (N_749,N_126,In_909);
nor U750 (N_750,In_1891,N_218);
and U751 (N_751,In_1727,N_420);
or U752 (N_752,In_1303,N_411);
nor U753 (N_753,In_1858,In_519);
nor U754 (N_754,In_827,In_575);
or U755 (N_755,In_688,In_2183);
or U756 (N_756,N_655,In_899);
nand U757 (N_757,In_2300,In_1896);
nor U758 (N_758,N_583,N_642);
nand U759 (N_759,In_116,N_550);
nand U760 (N_760,In_2233,In_2099);
or U761 (N_761,In_667,N_694);
and U762 (N_762,In_146,N_48);
and U763 (N_763,In_2284,N_500);
and U764 (N_764,In_2196,In_1418);
or U765 (N_765,N_610,In_12);
nand U766 (N_766,In_1825,N_165);
or U767 (N_767,In_894,In_1072);
or U768 (N_768,N_315,In_1192);
nand U769 (N_769,In_1198,In_1573);
nor U770 (N_770,In_2251,In_2247);
and U771 (N_771,In_387,In_2125);
xnor U772 (N_772,N_674,In_236);
nand U773 (N_773,In_2118,N_300);
nor U774 (N_774,N_330,In_1023);
or U775 (N_775,N_303,In_2120);
nor U776 (N_776,In_366,N_697);
or U777 (N_777,In_2444,In_1612);
nor U778 (N_778,N_705,In_1454);
and U779 (N_779,In_1562,In_18);
nor U780 (N_780,In_210,In_317);
nor U781 (N_781,In_2364,N_223);
and U782 (N_782,N_289,N_436);
or U783 (N_783,In_386,N_486);
xnor U784 (N_784,In_2312,In_1852);
and U785 (N_785,N_74,N_119);
nand U786 (N_786,N_187,In_648);
nand U787 (N_787,N_82,In_2426);
and U788 (N_788,In_1002,N_221);
nand U789 (N_789,In_1527,In_1391);
or U790 (N_790,In_1068,N_39);
nor U791 (N_791,In_2135,In_838);
xnor U792 (N_792,N_358,In_677);
nor U793 (N_793,N_574,N_91);
and U794 (N_794,In_2437,N_725);
nor U795 (N_795,N_539,In_1476);
nor U796 (N_796,In_820,In_2395);
nor U797 (N_797,N_305,In_221);
or U798 (N_798,N_483,In_1837);
or U799 (N_799,N_631,In_1569);
nand U800 (N_800,In_469,In_1704);
and U801 (N_801,In_2488,N_143);
nand U802 (N_802,In_232,In_1426);
and U803 (N_803,In_1764,N_559);
nor U804 (N_804,N_446,In_52);
and U805 (N_805,In_1374,N_153);
or U806 (N_806,In_1112,In_46);
nand U807 (N_807,In_1276,In_1031);
or U808 (N_808,In_1446,In_1499);
and U809 (N_809,In_1554,In_243);
and U810 (N_810,In_1841,In_420);
or U811 (N_811,N_637,In_1905);
nand U812 (N_812,N_40,In_2397);
xor U813 (N_813,In_1427,In_73);
and U814 (N_814,N_136,In_42);
or U815 (N_815,In_974,N_682);
or U816 (N_816,In_106,In_1706);
nor U817 (N_817,N_614,N_46);
or U818 (N_818,In_1971,In_1086);
nor U819 (N_819,In_2107,In_1413);
or U820 (N_820,In_1632,In_2454);
or U821 (N_821,N_676,In_1539);
or U822 (N_822,N_177,In_2468);
or U823 (N_823,In_618,In_181);
xnor U824 (N_824,N_670,N_568);
and U825 (N_825,In_1524,In_269);
xor U826 (N_826,In_640,N_596);
nand U827 (N_827,In_1721,N_76);
and U828 (N_828,In_1563,In_1867);
nor U829 (N_829,N_578,N_336);
and U830 (N_830,N_540,N_733);
nor U831 (N_831,In_2273,N_185);
nor U832 (N_832,In_845,In_1866);
nand U833 (N_833,N_570,In_1281);
and U834 (N_834,N_561,In_1381);
nor U835 (N_835,In_1206,In_863);
and U836 (N_836,In_1757,In_1285);
xor U837 (N_837,N_162,N_666);
nand U838 (N_838,In_1338,In_1738);
nand U839 (N_839,In_444,In_1506);
or U840 (N_840,In_2169,N_345);
nor U841 (N_841,N_206,In_2457);
nor U842 (N_842,In_2378,In_787);
nor U843 (N_843,In_2494,In_1691);
and U844 (N_844,In_1684,In_1787);
nand U845 (N_845,In_390,In_623);
or U846 (N_846,N_279,In_1753);
nand U847 (N_847,In_426,N_553);
and U848 (N_848,N_609,N_498);
nor U849 (N_849,N_4,In_15);
nor U850 (N_850,In_1012,In_518);
nor U851 (N_851,In_2299,In_400);
and U852 (N_852,N_222,N_53);
and U853 (N_853,In_711,N_320);
and U854 (N_854,In_634,N_719);
nor U855 (N_855,In_2214,N_79);
or U856 (N_856,N_3,N_522);
nor U857 (N_857,In_684,In_165);
xor U858 (N_858,In_2106,In_2059);
and U859 (N_859,In_1414,In_2086);
and U860 (N_860,In_647,In_1783);
or U861 (N_861,In_442,In_1128);
xnor U862 (N_862,N_603,N_0);
xor U863 (N_863,In_979,N_399);
and U864 (N_864,N_649,In_1546);
and U865 (N_865,In_455,N_662);
or U866 (N_866,N_386,N_556);
xnor U867 (N_867,In_242,In_1761);
and U868 (N_868,In_417,In_664);
or U869 (N_869,N_530,In_67);
or U870 (N_870,In_775,In_299);
nor U871 (N_871,In_697,In_2255);
xor U872 (N_872,In_169,In_512);
nor U873 (N_873,N_369,In_50);
nor U874 (N_874,N_660,N_602);
nand U875 (N_875,In_2066,In_726);
nor U876 (N_876,In_969,N_441);
or U877 (N_877,In_1786,In_1158);
nor U878 (N_878,In_1922,In_2148);
xor U879 (N_879,N_371,N_131);
nor U880 (N_880,In_1046,In_1600);
xnor U881 (N_881,N_88,In_1485);
xnor U882 (N_882,In_326,N_509);
nand U883 (N_883,In_1920,In_763);
nand U884 (N_884,In_1232,In_85);
or U885 (N_885,N_248,In_2162);
nor U886 (N_886,In_2048,In_49);
nand U887 (N_887,N_468,N_142);
nand U888 (N_888,In_1005,In_828);
or U889 (N_889,In_193,In_83);
nor U890 (N_890,In_1139,N_503);
nor U891 (N_891,In_1718,N_749);
and U892 (N_892,In_108,In_2475);
xnor U893 (N_893,In_464,In_1769);
nor U894 (N_894,N_597,In_2425);
or U895 (N_895,In_2070,In_207);
nor U896 (N_896,N_663,In_702);
nor U897 (N_897,In_2174,In_1890);
nand U898 (N_898,In_764,N_85);
nor U899 (N_899,In_645,N_292);
and U900 (N_900,N_363,N_238);
nand U901 (N_901,In_981,N_61);
nor U902 (N_902,In_1479,In_22);
and U903 (N_903,In_1957,In_151);
xnor U904 (N_904,In_554,N_295);
or U905 (N_905,N_658,In_2434);
nand U906 (N_906,N_742,N_690);
or U907 (N_907,In_619,N_661);
xnor U908 (N_908,In_1077,N_517);
nand U909 (N_909,In_504,N_669);
nand U910 (N_910,In_2168,N_692);
or U911 (N_911,N_708,In_2451);
nor U912 (N_912,In_1601,In_694);
or U913 (N_913,N_493,In_1402);
and U914 (N_914,In_235,In_440);
nor U915 (N_915,N_548,N_424);
or U916 (N_916,N_24,In_300);
nor U917 (N_917,In_884,In_2359);
nand U918 (N_918,In_874,In_51);
nor U919 (N_919,N_152,In_2458);
xnor U920 (N_920,In_527,In_2302);
and U921 (N_921,In_767,N_668);
xor U922 (N_922,In_1576,In_707);
or U923 (N_923,In_279,In_1835);
xor U924 (N_924,N_412,N_335);
nor U925 (N_925,N_656,N_581);
or U926 (N_926,In_1466,In_1015);
or U927 (N_927,In_1934,In_1821);
or U928 (N_928,In_2409,N_189);
nand U929 (N_929,In_1145,In_1714);
or U930 (N_930,N_710,In_316);
xnor U931 (N_931,In_2268,In_218);
xnor U932 (N_932,N_173,In_1432);
or U933 (N_933,N_182,N_72);
nand U934 (N_934,In_1190,In_885);
or U935 (N_935,N_334,In_1514);
xor U936 (N_936,N_179,In_1717);
or U937 (N_937,In_1129,N_277);
or U938 (N_938,In_1327,In_2037);
nand U939 (N_939,In_2035,In_1408);
nand U940 (N_940,N_713,In_2160);
nand U941 (N_941,In_17,In_470);
nand U942 (N_942,In_327,N_640);
nand U943 (N_943,In_1587,In_2480);
or U944 (N_944,N_536,In_164);
and U945 (N_945,In_1368,In_2456);
and U946 (N_946,N_364,In_1486);
nand U947 (N_947,N_124,In_814);
or U948 (N_948,In_2203,N_621);
nor U949 (N_949,In_1451,In_895);
nor U950 (N_950,In_1360,In_1249);
and U951 (N_951,N_47,In_1655);
or U952 (N_952,In_908,In_1386);
or U953 (N_953,In_1321,In_2438);
xor U954 (N_954,In_1107,In_1292);
nand U955 (N_955,In_2400,In_2250);
or U956 (N_956,In_1484,N_87);
nor U957 (N_957,In_1221,In_20);
nand U958 (N_958,In_1189,In_573);
xor U959 (N_959,N_495,In_1322);
or U960 (N_960,In_2241,In_678);
and U961 (N_961,N_529,N_121);
nor U962 (N_962,N_440,In_900);
and U963 (N_963,N_366,N_688);
nor U964 (N_964,In_2218,In_427);
nand U965 (N_965,In_403,In_2417);
xnor U966 (N_966,In_1502,In_1130);
and U967 (N_967,In_544,In_1296);
and U968 (N_968,In_328,In_2150);
nand U969 (N_969,In_725,In_1438);
and U970 (N_970,In_676,In_2463);
or U971 (N_971,In_826,N_437);
and U972 (N_972,In_2095,N_351);
nor U973 (N_973,In_9,N_560);
xor U974 (N_974,N_249,In_1063);
nand U975 (N_975,In_1071,In_1442);
nand U976 (N_976,In_1137,In_1040);
or U977 (N_977,In_2216,N_477);
nand U978 (N_978,In_1741,In_129);
nand U979 (N_979,N_558,In_1375);
or U980 (N_980,In_2173,In_557);
and U981 (N_981,In_1968,N_312);
and U982 (N_982,In_1892,In_633);
and U983 (N_983,In_1523,In_1051);
and U984 (N_984,In_206,In_2388);
nand U985 (N_985,N_154,In_1912);
or U986 (N_986,In_784,In_1808);
or U987 (N_987,In_603,In_1633);
nand U988 (N_988,In_1719,In_1942);
or U989 (N_989,In_881,N_619);
nand U990 (N_990,In_353,In_1114);
nand U991 (N_991,In_1493,N_504);
and U992 (N_992,In_1313,N_528);
nor U993 (N_993,N_217,N_341);
xnor U994 (N_994,In_1897,In_1680);
nor U995 (N_995,In_608,In_1449);
or U996 (N_996,N_741,In_40);
and U997 (N_997,N_269,In_1020);
nand U998 (N_998,In_1215,In_408);
or U999 (N_999,N_634,In_1975);
or U1000 (N_1000,N_29,In_2353);
nor U1001 (N_1001,N_242,N_897);
or U1002 (N_1002,In_808,N_851);
nor U1003 (N_1003,In_2320,In_1883);
or U1004 (N_1004,N_321,In_501);
nor U1005 (N_1005,N_999,In_1639);
or U1006 (N_1006,In_368,N_739);
nor U1007 (N_1007,N_639,In_1266);
nor U1008 (N_1008,N_992,In_1651);
or U1009 (N_1009,N_620,In_86);
and U1010 (N_1010,In_1283,In_480);
or U1011 (N_1011,In_228,N_452);
or U1012 (N_1012,In_1803,N_651);
nand U1013 (N_1013,In_2276,N_779);
nand U1014 (N_1014,N_847,In_565);
and U1015 (N_1015,N_447,In_868);
and U1016 (N_1016,In_192,N_795);
or U1017 (N_1017,In_297,In_745);
nand U1018 (N_1018,N_970,In_776);
nor U1019 (N_1019,In_75,N_902);
nand U1020 (N_1020,N_308,N_931);
xor U1021 (N_1021,In_996,In_1766);
and U1022 (N_1022,In_1343,N_197);
nand U1023 (N_1023,In_2013,N_382);
xor U1024 (N_1024,In_2085,In_2328);
nor U1025 (N_1025,In_2038,In_1909);
or U1026 (N_1026,In_1952,N_723);
nand U1027 (N_1027,N_271,In_227);
or U1028 (N_1028,In_655,In_177);
and U1029 (N_1029,In_1767,N_839);
and U1030 (N_1030,In_1464,N_298);
and U1031 (N_1031,In_449,N_52);
xor U1032 (N_1032,In_923,In_675);
and U1033 (N_1033,In_2366,In_1042);
nand U1034 (N_1034,N_938,In_1270);
or U1035 (N_1035,N_647,In_1488);
nor U1036 (N_1036,N_911,In_363);
nor U1037 (N_1037,In_1522,N_332);
or U1038 (N_1038,In_1599,In_394);
xor U1039 (N_1039,In_362,N_572);
and U1040 (N_1040,In_2029,In_1109);
and U1041 (N_1041,In_691,In_2470);
or U1042 (N_1042,In_304,N_435);
or U1043 (N_1043,N_982,In_2159);
xnor U1044 (N_1044,In_821,In_2390);
or U1045 (N_1045,In_1448,N_178);
and U1046 (N_1046,In_572,In_2462);
nand U1047 (N_1047,In_701,In_433);
nor U1048 (N_1048,N_790,N_627);
or U1049 (N_1049,In_2286,In_2224);
or U1050 (N_1050,In_1547,N_808);
and U1051 (N_1051,In_2193,In_1654);
nand U1052 (N_1052,In_121,In_1888);
nor U1053 (N_1053,In_615,N_978);
and U1054 (N_1054,N_962,In_542);
and U1055 (N_1055,N_203,In_1216);
xnor U1056 (N_1056,N_645,N_680);
or U1057 (N_1057,In_1274,In_1197);
nor U1058 (N_1058,N_49,N_826);
nor U1059 (N_1059,In_34,In_1111);
or U1060 (N_1060,N_715,In_1693);
xnor U1061 (N_1061,N_125,In_550);
nand U1062 (N_1062,In_1302,N_283);
and U1063 (N_1063,In_2052,In_1998);
nor U1064 (N_1064,N_585,In_1855);
and U1065 (N_1065,N_325,In_2103);
nor U1066 (N_1066,N_755,N_511);
and U1067 (N_1067,In_2030,N_66);
nor U1068 (N_1068,N_626,N_909);
nor U1069 (N_1069,In_819,In_283);
xor U1070 (N_1070,N_35,In_1491);
and U1071 (N_1071,In_171,N_699);
nand U1072 (N_1072,In_2281,In_1498);
nand U1073 (N_1073,In_949,In_1842);
and U1074 (N_1074,In_1090,In_143);
nand U1075 (N_1075,In_36,In_2282);
nand U1076 (N_1076,In_2384,N_785);
or U1077 (N_1077,In_1986,N_226);
and U1078 (N_1078,N_109,In_2122);
and U1079 (N_1079,N_307,N_869);
and U1080 (N_1080,In_995,N_787);
and U1081 (N_1081,N_340,N_290);
nor U1082 (N_1082,N_252,N_616);
xor U1083 (N_1083,N_258,In_2130);
nor U1084 (N_1084,In_1242,In_943);
and U1085 (N_1085,N_291,N_789);
and U1086 (N_1086,In_2446,In_1643);
nand U1087 (N_1087,N_624,In_2340);
nand U1088 (N_1088,In_126,N_494);
or U1089 (N_1089,In_318,N_729);
and U1090 (N_1090,N_980,N_533);
and U1091 (N_1091,In_1796,N_219);
and U1092 (N_1092,In_1286,N_594);
nand U1093 (N_1093,N_37,N_13);
and U1094 (N_1094,In_525,N_469);
and U1095 (N_1095,In_530,In_2110);
and U1096 (N_1096,In_549,In_1700);
or U1097 (N_1097,In_1127,In_2271);
or U1098 (N_1098,In_771,In_2389);
xor U1099 (N_1099,In_2305,In_2477);
and U1100 (N_1100,In_1871,N_801);
nand U1101 (N_1101,N_497,In_1860);
nand U1102 (N_1102,In_1219,N_267);
and U1103 (N_1103,In_2026,In_1849);
or U1104 (N_1104,In_1862,In_505);
nand U1105 (N_1105,In_1389,In_1315);
nor U1106 (N_1106,In_1955,In_2098);
nor U1107 (N_1107,N_714,In_486);
and U1108 (N_1108,In_439,N_943);
and U1109 (N_1109,In_2226,N_623);
or U1110 (N_1110,N_562,N_679);
nor U1111 (N_1111,N_403,In_1705);
nor U1112 (N_1112,In_1097,In_836);
nand U1113 (N_1113,In_446,N_958);
and U1114 (N_1114,In_945,In_2147);
nor U1115 (N_1115,N_98,In_1959);
xnor U1116 (N_1116,In_1235,N_535);
xnor U1117 (N_1117,In_142,In_245);
nand U1118 (N_1118,In_2207,N_780);
nand U1119 (N_1119,N_433,N_989);
or U1120 (N_1120,In_1774,N_895);
or U1121 (N_1121,In_559,In_679);
or U1122 (N_1122,N_716,N_934);
nor U1123 (N_1123,In_2350,N_246);
nor U1124 (N_1124,N_520,N_976);
nor U1125 (N_1125,In_2053,N_671);
nor U1126 (N_1126,In_1876,In_1096);
and U1127 (N_1127,N_593,In_330);
nand U1128 (N_1128,In_1822,N_898);
and U1129 (N_1129,In_720,In_2131);
nand U1130 (N_1130,In_709,In_1262);
nor U1131 (N_1131,In_977,In_1463);
and U1132 (N_1132,In_2136,In_407);
or U1133 (N_1133,In_2232,N_990);
xnor U1134 (N_1134,N_629,In_563);
xor U1135 (N_1135,In_1833,N_445);
and U1136 (N_1136,N_860,In_870);
or U1137 (N_1137,N_17,N_906);
or U1138 (N_1138,In_1652,In_45);
nand U1139 (N_1139,N_393,In_1095);
nor U1140 (N_1140,In_2223,In_1965);
nand U1141 (N_1141,In_471,In_984);
and U1142 (N_1142,In_924,N_170);
xnor U1143 (N_1143,N_914,In_1347);
and U1144 (N_1144,In_783,In_2165);
and U1145 (N_1145,In_2003,N_863);
and U1146 (N_1146,N_395,N_378);
or U1147 (N_1147,N_961,N_357);
and U1148 (N_1148,N_134,In_2399);
nor U1149 (N_1149,In_1212,In_1900);
and U1150 (N_1150,In_736,In_1671);
and U1151 (N_1151,N_188,N_912);
or U1152 (N_1152,In_47,In_2429);
or U1153 (N_1153,N_580,N_685);
nor U1154 (N_1154,N_130,In_590);
and U1155 (N_1155,N_346,N_775);
nand U1156 (N_1156,N_280,In_1333);
nand U1157 (N_1157,N_577,In_1530);
or U1158 (N_1158,N_782,N_868);
and U1159 (N_1159,N_555,In_1755);
nor U1160 (N_1160,In_1829,In_1483);
xnor U1161 (N_1161,N_549,In_393);
or U1162 (N_1162,N_525,In_1864);
xnor U1163 (N_1163,In_620,N_956);
or U1164 (N_1164,N_969,In_2370);
xor U1165 (N_1165,N_967,In_1143);
and U1166 (N_1166,N_294,In_1461);
and U1167 (N_1167,N_380,N_352);
and U1168 (N_1168,N_939,N_361);
nand U1169 (N_1169,N_390,In_2119);
or U1170 (N_1170,In_1555,In_2391);
or U1171 (N_1171,In_2332,N_880);
nand U1172 (N_1172,In_1591,N_829);
nand U1173 (N_1173,N_945,In_447);
nand U1174 (N_1174,In_329,In_93);
and U1175 (N_1175,In_438,In_1099);
or U1176 (N_1176,N_882,N_879);
nand U1177 (N_1177,In_770,In_532);
and U1178 (N_1178,In_612,N_544);
or U1179 (N_1179,In_2355,N_665);
nor U1180 (N_1180,N_648,In_693);
and U1181 (N_1181,In_163,N_490);
nor U1182 (N_1182,In_1010,In_1115);
nor U1183 (N_1183,N_748,In_2206);
and U1184 (N_1184,In_262,In_367);
and U1185 (N_1185,N_542,In_2421);
or U1186 (N_1186,N_51,N_852);
nor U1187 (N_1187,In_1901,In_875);
nand U1188 (N_1188,N_871,In_795);
and U1189 (N_1189,In_2341,In_600);
nor U1190 (N_1190,In_1104,In_2487);
and U1191 (N_1191,In_338,In_1791);
nand U1192 (N_1192,N_359,In_1674);
and U1193 (N_1193,N_858,In_1168);
nand U1194 (N_1194,N_590,N_804);
nor U1195 (N_1195,N_750,N_732);
nand U1196 (N_1196,In_1191,In_1497);
and U1197 (N_1197,In_1272,N_903);
or U1198 (N_1198,In_2114,N_709);
nand U1199 (N_1199,N_870,In_2404);
nor U1200 (N_1200,In_610,N_41);
and U1201 (N_1201,In_1869,N_510);
and U1202 (N_1202,In_686,In_289);
and U1203 (N_1203,In_1967,N_472);
or U1204 (N_1204,In_1874,N_381);
xnor U1205 (N_1205,In_1026,In_1264);
nand U1206 (N_1206,N_343,In_1882);
xor U1207 (N_1207,In_1541,N_862);
nand U1208 (N_1208,N_145,N_937);
nor U1209 (N_1209,N_84,N_696);
or U1210 (N_1210,N_461,In_1180);
or U1211 (N_1211,N_877,N_575);
nand U1212 (N_1212,In_1240,In_2288);
or U1213 (N_1213,In_2365,In_2208);
nand U1214 (N_1214,In_1597,In_529);
or U1215 (N_1215,In_2044,In_1660);
xnor U1216 (N_1216,In_1542,N_796);
or U1217 (N_1217,In_478,In_1081);
nand U1218 (N_1218,In_141,N_949);
nand U1219 (N_1219,In_749,In_2269);
nand U1220 (N_1220,In_1811,N_726);
and U1221 (N_1221,In_2352,In_548);
nor U1222 (N_1222,In_1557,N_508);
nand U1223 (N_1223,In_987,N_516);
or U1224 (N_1224,In_994,N_657);
or U1225 (N_1225,In_1224,N_855);
xor U1226 (N_1226,N_474,N_947);
and U1227 (N_1227,N_239,N_442);
and U1228 (N_1228,In_168,In_2381);
and U1229 (N_1229,N_579,In_2047);
xnor U1230 (N_1230,In_425,In_1244);
nand U1231 (N_1231,N_427,In_1784);
and U1232 (N_1232,In_1376,In_500);
nand U1233 (N_1233,N_773,N_598);
xor U1234 (N_1234,In_609,N_557);
or U1235 (N_1235,N_915,In_850);
nor U1236 (N_1236,N_722,N_878);
nand U1237 (N_1237,N_481,In_373);
or U1238 (N_1238,In_807,In_1958);
nor U1239 (N_1239,In_1927,In_1123);
and U1240 (N_1240,N_409,N_738);
nor U1241 (N_1241,N_638,In_541);
or U1242 (N_1242,In_1379,N_830);
nand U1243 (N_1243,In_2209,In_2280);
and U1244 (N_1244,In_2084,In_2325);
nor U1245 (N_1245,N_834,N_964);
nor U1246 (N_1246,N_458,N_56);
nor U1247 (N_1247,In_1151,In_30);
or U1248 (N_1248,In_1938,N_379);
or U1249 (N_1249,In_113,N_942);
nor U1250 (N_1250,N_337,In_703);
nor U1251 (N_1251,In_1745,In_769);
nand U1252 (N_1252,N_819,In_2249);
nor U1253 (N_1253,In_551,In_728);
or U1254 (N_1254,N_1152,N_418);
nor U1255 (N_1255,In_2375,In_524);
nor U1256 (N_1256,N_1162,N_1038);
and U1257 (N_1257,N_1180,N_711);
or U1258 (N_1258,In_887,In_1055);
and U1259 (N_1259,In_1564,In_1265);
and U1260 (N_1260,In_599,N_1044);
nand U1261 (N_1261,N_963,N_274);
nand U1262 (N_1262,In_904,N_1246);
nor U1263 (N_1263,N_1236,N_1135);
nor U1264 (N_1264,N_316,In_482);
and U1265 (N_1265,N_650,In_220);
and U1266 (N_1266,N_1120,N_524);
nand U1267 (N_1267,N_975,N_118);
nor U1268 (N_1268,In_1255,In_1853);
and U1269 (N_1269,In_2333,N_925);
nor U1270 (N_1270,N_1178,In_383);
nand U1271 (N_1271,N_230,N_979);
and U1272 (N_1272,In_379,N_476);
or U1273 (N_1273,In_334,N_684);
and U1274 (N_1274,N_211,N_1209);
and U1275 (N_1275,N_434,In_1861);
nand U1276 (N_1276,In_1838,In_1183);
or U1277 (N_1277,In_102,N_768);
xnor U1278 (N_1278,In_2393,In_1616);
xor U1279 (N_1279,In_436,N_1203);
xnor U1280 (N_1280,N_1244,In_1709);
and U1281 (N_1281,N_1102,N_1176);
xor U1282 (N_1282,N_1141,In_2040);
and U1283 (N_1283,In_1367,N_948);
or U1284 (N_1284,N_928,N_410);
or U1285 (N_1285,In_1701,N_241);
or U1286 (N_1286,N_261,In_412);
or U1287 (N_1287,N_534,N_526);
nand U1288 (N_1288,N_986,N_747);
or U1289 (N_1289,In_1395,N_740);
nand U1290 (N_1290,N_176,In_302);
nand U1291 (N_1291,In_271,In_1425);
xor U1292 (N_1292,In_2076,N_1006);
nor U1293 (N_1293,N_565,N_1169);
nand U1294 (N_1294,N_720,N_457);
or U1295 (N_1295,In_2234,N_735);
or U1296 (N_1296,In_59,N_900);
or U1297 (N_1297,N_1031,In_454);
nand U1298 (N_1298,In_404,In_2033);
or U1299 (N_1299,In_249,N_554);
nand U1300 (N_1300,In_651,N_611);
nand U1301 (N_1301,N_617,N_991);
nand U1302 (N_1302,In_1559,N_90);
nor U1303 (N_1303,N_922,N_1230);
nor U1304 (N_1304,N_933,N_1098);
nor U1305 (N_1305,N_1082,N_1182);
or U1306 (N_1306,N_478,In_1233);
and U1307 (N_1307,N_489,N_195);
nor U1308 (N_1308,In_148,N_1144);
or U1309 (N_1309,In_2464,N_1020);
nor U1310 (N_1310,In_2154,In_998);
nor U1311 (N_1311,N_26,In_905);
and U1312 (N_1312,N_110,N_253);
and U1313 (N_1313,N_1047,N_1061);
nor U1314 (N_1314,In_601,In_1250);
xor U1315 (N_1315,In_2408,N_225);
nor U1316 (N_1316,In_2072,N_784);
nor U1317 (N_1317,N_1243,N_944);
and U1318 (N_1318,In_2146,N_576);
xnor U1319 (N_1319,N_1042,In_354);
and U1320 (N_1320,In_2064,In_1035);
and U1321 (N_1321,N_408,N_817);
or U1322 (N_1322,N_950,N_890);
and U1323 (N_1323,In_451,N_205);
xnor U1324 (N_1324,N_444,In_569);
and U1325 (N_1325,N_288,In_760);
xor U1326 (N_1326,In_2270,N_5);
xnor U1327 (N_1327,N_1043,In_340);
nand U1328 (N_1328,N_1123,In_2004);
nor U1329 (N_1329,In_263,N_77);
nand U1330 (N_1330,In_133,N_1118);
nor U1331 (N_1331,In_1549,N_633);
nor U1332 (N_1332,N_1248,N_523);
nor U1333 (N_1333,In_922,N_1233);
nand U1334 (N_1334,N_1214,In_1148);
and U1335 (N_1335,In_54,N_923);
or U1336 (N_1336,N_764,In_172);
xor U1337 (N_1337,In_890,N_396);
nor U1338 (N_1338,N_443,N_1156);
nand U1339 (N_1339,In_983,N_1148);
and U1340 (N_1340,In_574,In_1320);
nand U1341 (N_1341,N_348,N_1129);
nor U1342 (N_1342,N_635,N_985);
nand U1343 (N_1343,N_762,In_2041);
nand U1344 (N_1344,In_611,N_734);
and U1345 (N_1345,In_2074,N_605);
xnor U1346 (N_1346,N_1110,In_2015);
or U1347 (N_1347,In_1382,N_1015);
nor U1348 (N_1348,N_1133,N_1062);
and U1349 (N_1349,N_673,N_894);
nand U1350 (N_1350,In_87,N_1093);
nor U1351 (N_1351,N_492,In_1416);
nor U1352 (N_1352,In_2046,N_763);
nand U1353 (N_1353,N_1245,N_236);
nor U1354 (N_1354,In_1447,In_2063);
and U1355 (N_1355,N_196,N_1012);
and U1356 (N_1356,In_2339,In_57);
nand U1357 (N_1357,N_1134,N_803);
nand U1358 (N_1358,In_1335,N_1139);
nand U1359 (N_1359,N_974,In_1624);
nor U1360 (N_1360,In_2424,N_850);
or U1361 (N_1361,In_1801,In_2213);
nor U1362 (N_1362,N_1228,N_2);
xor U1363 (N_1363,N_636,N_150);
and U1364 (N_1364,N_329,N_133);
nand U1365 (N_1365,In_1317,N_806);
and U1366 (N_1366,N_1018,In_1415);
and U1367 (N_1367,N_761,In_614);
nor U1368 (N_1368,N_587,In_1824);
xor U1369 (N_1369,N_1019,N_717);
and U1370 (N_1370,In_604,In_1578);
nand U1371 (N_1371,In_1070,In_659);
and U1372 (N_1372,In_490,N_1237);
or U1373 (N_1373,N_872,N_916);
and U1374 (N_1374,In_1580,In_1663);
or U1375 (N_1375,In_1556,N_1009);
and U1376 (N_1376,In_280,In_743);
or U1377 (N_1377,N_1140,N_9);
and U1378 (N_1378,N_19,N_756);
xor U1379 (N_1379,N_812,N_11);
nor U1380 (N_1380,N_28,N_856);
nand U1381 (N_1381,N_301,N_552);
nand U1382 (N_1382,N_724,N_1112);
nor U1383 (N_1383,In_1319,In_800);
or U1384 (N_1384,N_1083,N_93);
nand U1385 (N_1385,N_844,In_290);
and U1386 (N_1386,N_930,In_1409);
or U1387 (N_1387,In_1744,N_551);
and U1388 (N_1388,In_2265,N_1194);
nand U1389 (N_1389,In_2121,In_2459);
nand U1390 (N_1390,In_1478,In_415);
and U1391 (N_1391,N_1094,In_1775);
and U1392 (N_1392,N_455,In_2113);
nor U1393 (N_1393,In_2303,In_1503);
and U1394 (N_1394,N_888,In_893);
nand U1395 (N_1395,N_169,In_131);
and U1396 (N_1396,N_347,In_1630);
or U1397 (N_1397,In_1101,In_154);
and U1398 (N_1398,N_1146,N_573);
nor U1399 (N_1399,N_1053,In_1507);
nand U1400 (N_1400,N_1185,N_977);
nor U1401 (N_1401,In_491,In_1048);
nor U1402 (N_1402,In_2478,In_1351);
nor U1403 (N_1403,In_1681,N_1153);
or U1404 (N_1404,In_606,In_670);
nand U1405 (N_1405,N_1100,In_2211);
xnor U1406 (N_1406,N_1174,In_938);
nor U1407 (N_1407,N_1201,N_731);
and U1408 (N_1408,In_2308,In_952);
or U1409 (N_1409,In_1749,In_761);
and U1410 (N_1410,In_629,In_1566);
or U1411 (N_1411,In_1511,N_1034);
nor U1412 (N_1412,N_286,N_1132);
or U1413 (N_1413,In_1369,N_571);
nand U1414 (N_1414,N_867,N_588);
nand U1415 (N_1415,N_918,N_569);
xnor U1416 (N_1416,In_558,N_825);
and U1417 (N_1417,N_453,N_1109);
nor U1418 (N_1418,N_774,In_2497);
nor U1419 (N_1419,N_546,In_2264);
nor U1420 (N_1420,In_1973,N_777);
and U1421 (N_1421,In_1400,In_980);
or U1422 (N_1422,In_1536,N_1101);
nor U1423 (N_1423,N_338,N_997);
nor U1424 (N_1424,N_625,N_512);
nor U1425 (N_1425,N_564,In_2016);
nor U1426 (N_1426,In_74,N_1071);
nor U1427 (N_1427,N_1215,N_896);
xnor U1428 (N_1428,In_724,In_933);
nand U1429 (N_1429,In_1720,N_389);
nor U1430 (N_1430,In_772,N_693);
or U1431 (N_1431,N_1191,N_686);
nor U1432 (N_1432,In_247,In_158);
nor U1433 (N_1433,N_893,In_267);
nor U1434 (N_1434,N_816,N_955);
nand U1435 (N_1435,In_136,N_1216);
nand U1436 (N_1436,In_700,In_1300);
nor U1437 (N_1437,N_1088,In_310);
nor U1438 (N_1438,N_65,N_106);
nand U1439 (N_1439,In_1515,In_2405);
nand U1440 (N_1440,In_1602,N_953);
xnor U1441 (N_1441,N_102,In_1735);
xor U1442 (N_1442,N_1160,N_1087);
nand U1443 (N_1443,In_2358,N_531);
and U1444 (N_1444,In_2077,N_243);
nor U1445 (N_1445,In_1777,N_1151);
nor U1446 (N_1446,N_840,N_841);
nor U1447 (N_1447,In_1290,In_1358);
and U1448 (N_1448,N_304,In_801);
and U1449 (N_1449,In_1392,N_584);
or U1450 (N_1450,In_465,In_314);
xor U1451 (N_1451,N_891,N_1202);
and U1452 (N_1452,N_1161,In_730);
or U1453 (N_1453,N_772,In_1676);
nand U1454 (N_1454,N_36,In_796);
nand U1455 (N_1455,N_1104,N_887);
and U1456 (N_1456,N_384,In_546);
xor U1457 (N_1457,In_2215,N_1124);
xnor U1458 (N_1458,N_1143,In_176);
nand U1459 (N_1459,In_223,N_972);
or U1460 (N_1460,N_1108,N_917);
or U1461 (N_1461,N_1219,N_545);
and U1462 (N_1462,N_776,N_1131);
nor U1463 (N_1463,N_707,N_667);
or U1464 (N_1464,In_1799,N_1234);
or U1465 (N_1465,N_957,N_1217);
and U1466 (N_1466,N_814,N_160);
or U1467 (N_1467,In_1423,In_323);
or U1468 (N_1468,N_328,N_43);
and U1469 (N_1469,N_425,In_11);
or U1470 (N_1470,In_2278,In_523);
nand U1471 (N_1471,In_125,N_1002);
and U1472 (N_1472,N_1218,In_786);
or U1473 (N_1473,In_2347,In_2139);
nand U1474 (N_1474,In_1594,N_1045);
or U1475 (N_1475,In_135,N_1165);
or U1476 (N_1476,N_876,In_1748);
or U1477 (N_1477,N_1138,N_960);
nand U1478 (N_1478,N_1058,N_1079);
nand U1479 (N_1479,In_817,N_473);
and U1480 (N_1480,N_794,In_1411);
nand U1481 (N_1481,N_1051,N_1207);
or U1482 (N_1482,N_324,N_276);
and U1483 (N_1483,In_250,N_1028);
nor U1484 (N_1484,N_618,N_1184);
nor U1485 (N_1485,In_1373,In_275);
nand U1486 (N_1486,In_5,In_540);
or U1487 (N_1487,In_1988,In_1792);
nor U1488 (N_1488,N_521,In_2343);
and U1489 (N_1489,N_1142,N_157);
nor U1490 (N_1490,N_797,N_940);
and U1491 (N_1491,In_1383,N_1072);
and U1492 (N_1492,N_1008,N_865);
xnor U1493 (N_1493,N_706,N_432);
xor U1494 (N_1494,In_1165,N_278);
nor U1495 (N_1495,In_1404,N_1130);
or U1496 (N_1496,In_1208,N_843);
nor U1497 (N_1497,N_421,In_308);
or U1498 (N_1498,In_382,In_2010);
and U1499 (N_1499,In_2212,N_815);
or U1500 (N_1500,N_310,N_1323);
and U1501 (N_1501,In_1826,N_394);
nor U1502 (N_1502,N_92,N_537);
xnor U1503 (N_1503,N_566,In_1211);
and U1504 (N_1504,N_835,N_1242);
and U1505 (N_1505,N_1402,N_1367);
nand U1506 (N_1506,N_1326,In_1275);
and U1507 (N_1507,N_1173,In_865);
nand U1508 (N_1508,N_1375,N_1415);
or U1509 (N_1509,N_1336,N_1264);
and U1510 (N_1510,N_698,N_1493);
nor U1511 (N_1511,N_1434,N_966);
or U1512 (N_1512,N_1273,In_872);
or U1513 (N_1513,N_1171,In_960);
nor U1514 (N_1514,In_1353,N_207);
nor U1515 (N_1515,N_1190,N_1260);
and U1516 (N_1516,In_499,In_1648);
xor U1517 (N_1517,In_2171,N_1249);
nand U1518 (N_1518,In_1075,N_1479);
and U1519 (N_1519,N_1231,N_45);
or U1520 (N_1520,N_1250,N_1366);
or U1521 (N_1521,N_1181,In_748);
or U1522 (N_1522,N_1314,In_2149);
nor U1523 (N_1523,N_1103,N_1289);
or U1524 (N_1524,N_1384,N_1001);
and U1525 (N_1525,N_886,In_1263);
nand U1526 (N_1526,N_463,In_840);
or U1527 (N_1527,N_1052,N_622);
or U1528 (N_1528,In_857,In_2474);
nand U1529 (N_1529,N_1345,N_1294);
xnor U1530 (N_1530,N_746,N_262);
and U1531 (N_1531,N_1369,N_832);
nor U1532 (N_1532,N_1351,In_1294);
and U1533 (N_1533,In_468,N_27);
nand U1534 (N_1534,N_1374,In_114);
and U1535 (N_1535,N_1362,In_598);
nand U1536 (N_1536,In_650,N_971);
and U1537 (N_1537,N_1077,N_998);
nor U1538 (N_1538,N_1491,In_211);
and U1539 (N_1539,In_747,N_323);
nand U1540 (N_1540,N_752,In_1267);
nand U1541 (N_1541,In_1258,N_532);
nor U1542 (N_1542,N_1145,N_995);
nand U1543 (N_1543,N_449,N_1484);
nand U1544 (N_1544,N_1349,N_792);
and U1545 (N_1545,N_1443,N_541);
xor U1546 (N_1546,N_1128,N_1368);
nand U1547 (N_1547,N_331,In_1812);
nand U1548 (N_1548,N_1205,N_854);
nor U1549 (N_1549,In_2296,N_718);
nand U1550 (N_1550,In_1531,In_1146);
or U1551 (N_1551,N_1497,N_1428);
nand U1552 (N_1552,In_584,In_756);
nand U1553 (N_1553,N_1258,N_613);
nand U1554 (N_1554,N_1433,In_1428);
xor U1555 (N_1555,N_1227,N_1423);
nand U1556 (N_1556,N_1247,N_628);
and U1557 (N_1557,N_198,N_592);
nor U1558 (N_1558,N_1167,N_1412);
nor U1559 (N_1559,In_140,In_955);
or U1560 (N_1560,N_824,N_1357);
and U1561 (N_1561,N_172,N_385);
nand U1562 (N_1562,N_1409,N_282);
or U1563 (N_1563,In_418,N_260);
nand U1564 (N_1564,In_2088,In_526);
or U1565 (N_1565,In_2466,N_1495);
nor U1566 (N_1566,N_913,In_423);
nand U1567 (N_1567,N_1419,N_744);
or U1568 (N_1568,In_2011,In_779);
nor U1569 (N_1569,N_941,N_1445);
and U1570 (N_1570,N_586,N_1026);
nand U1571 (N_1571,In_1458,In_128);
and U1572 (N_1572,In_1669,N_1000);
xor U1573 (N_1573,N_1268,N_1159);
nor U1574 (N_1574,N_1195,N_1401);
or U1575 (N_1575,N_820,N_689);
or U1576 (N_1576,In_159,N_702);
and U1577 (N_1577,N_1192,In_2151);
or U1578 (N_1578,N_921,N_759);
nor U1579 (N_1579,In_2177,N_1256);
and U1580 (N_1580,N_78,N_1457);
nand U1581 (N_1581,In_2258,N_1424);
or U1582 (N_1582,N_712,N_1039);
nor U1583 (N_1583,N_1193,N_1251);
or U1584 (N_1584,N_1085,In_1658);
and U1585 (N_1585,In_217,N_1395);
or U1586 (N_1586,In_864,N_1347);
or U1587 (N_1587,N_885,In_1944);
or U1588 (N_1588,N_55,N_1252);
nand U1589 (N_1589,N_360,In_498);
and U1590 (N_1590,N_1150,N_1400);
nand U1591 (N_1591,N_884,N_1430);
nor U1592 (N_1592,In_1091,In_410);
nor U1593 (N_1593,N_1494,N_256);
and U1594 (N_1594,N_646,N_1489);
and U1595 (N_1595,N_1035,N_1288);
and U1596 (N_1596,N_1290,N_919);
or U1597 (N_1597,In_1919,N_1298);
xnor U1598 (N_1598,N_936,In_1184);
or U1599 (N_1599,In_2134,N_1292);
or U1600 (N_1600,In_1947,N_1106);
xnor U1601 (N_1601,N_1383,N_612);
nand U1602 (N_1602,In_88,N_1024);
or U1603 (N_1603,N_1377,N_1453);
or U1604 (N_1604,N_1320,In_719);
nand U1605 (N_1605,In_493,N_1059);
xor U1606 (N_1606,In_1747,N_1277);
nand U1607 (N_1607,In_824,N_1446);
xnor U1608 (N_1608,N_778,In_627);
nor U1609 (N_1609,N_823,N_632);
nand U1610 (N_1610,N_71,N_1163);
nor U1611 (N_1611,In_793,In_1989);
or U1612 (N_1612,In_935,In_1733);
and U1613 (N_1613,N_881,In_494);
nor U1614 (N_1614,N_1387,N_1056);
and U1615 (N_1615,N_615,N_1390);
nand U1616 (N_1616,N_1389,N_1472);
or U1617 (N_1617,N_1348,In_1007);
xor U1618 (N_1618,N_501,In_2143);
and U1619 (N_1619,N_419,In_1834);
and U1620 (N_1620,N_245,In_966);
or U1621 (N_1621,N_251,N_454);
or U1622 (N_1622,In_1388,In_456);
nor U1623 (N_1623,N_659,N_1498);
or U1624 (N_1624,In_1131,N_166);
nor U1625 (N_1625,In_2182,In_1016);
or U1626 (N_1626,N_168,N_1429);
or U1627 (N_1627,N_1335,N_1490);
or U1628 (N_1628,N_1027,N_1386);
or U1629 (N_1629,N_866,In_1230);
or U1630 (N_1630,N_837,N_1346);
nand U1631 (N_1631,In_1468,N_1302);
or U1632 (N_1632,N_1470,N_757);
nor U1633 (N_1633,N_1313,N_1378);
and U1634 (N_1634,In_2314,In_1234);
and U1635 (N_1635,In_1778,In_1649);
nor U1636 (N_1636,N_1370,N_255);
nor U1637 (N_1637,N_1281,In_773);
xnor U1638 (N_1638,In_281,N_1426);
nor U1639 (N_1639,N_786,N_1235);
nor U1640 (N_1640,N_751,In_138);
and U1641 (N_1641,In_251,In_940);
and U1642 (N_1642,N_1054,N_464);
or U1643 (N_1643,In_2021,N_1328);
and U1644 (N_1644,N_1421,In_117);
nor U1645 (N_1645,N_1333,N_833);
nor U1646 (N_1646,In_1963,N_1291);
nor U1647 (N_1647,N_874,N_1186);
nand U1648 (N_1648,N_1473,In_1879);
or U1649 (N_1649,In_520,In_953);
xor U1650 (N_1650,In_2083,N_653);
nand U1651 (N_1651,N_1399,In_72);
nor U1652 (N_1652,In_2089,N_1040);
or U1653 (N_1653,In_1142,In_1041);
or U1654 (N_1654,N_1063,N_1282);
nand U1655 (N_1655,In_2490,In_897);
nand U1656 (N_1656,N_438,N_1253);
and U1657 (N_1657,N_1004,In_2489);
or U1658 (N_1658,In_860,N_487);
nand U1659 (N_1659,In_215,In_1062);
xnor U1660 (N_1660,In_1260,In_1126);
or U1661 (N_1661,N_1444,N_1361);
nor U1662 (N_1662,N_771,In_892);
or U1663 (N_1663,N_743,N_1461);
nand U1664 (N_1664,N_1422,N_1211);
or U1665 (N_1665,N_1011,N_1439);
nand U1666 (N_1666,In_1299,N_1474);
or U1667 (N_1667,In_1790,In_777);
xnor U1668 (N_1668,N_1404,N_1239);
or U1669 (N_1669,N_1496,In_347);
xor U1670 (N_1670,N_704,N_1299);
nand U1671 (N_1671,N_1017,N_1226);
nand U1672 (N_1672,N_1065,In_1308);
nand U1673 (N_1673,N_987,N_822);
and U1674 (N_1674,In_2372,N_1316);
or U1675 (N_1675,N_1483,N_1050);
or U1676 (N_1676,In_1202,N_1324);
nand U1677 (N_1677,N_58,N_783);
nor U1678 (N_1678,N_1221,In_515);
or U1679 (N_1679,N_675,N_1080);
xnor U1680 (N_1680,N_664,In_1363);
xnor U1681 (N_1681,In_1699,N_1212);
and U1682 (N_1682,In_2219,In_1050);
nand U1683 (N_1683,N_1398,N_721);
or U1684 (N_1684,N_836,N_1304);
and U1685 (N_1685,N_1278,In_1371);
nor U1686 (N_1686,N_1391,In_150);
and U1687 (N_1687,N_387,N_1274);
nand U1688 (N_1688,In_1337,N_905);
nand U1689 (N_1689,In_32,N_344);
and U1690 (N_1690,N_1057,In_97);
nor U1691 (N_1691,N_1475,N_319);
or U1692 (N_1692,In_127,N_864);
nor U1693 (N_1693,N_1459,N_1344);
or U1694 (N_1694,N_861,N_1147);
nor U1695 (N_1695,N_952,In_2423);
and U1696 (N_1696,N_1223,N_515);
or U1697 (N_1697,N_981,N_1437);
xnor U1698 (N_1698,N_920,In_1209);
nand U1699 (N_1699,In_1768,N_994);
or U1700 (N_1700,N_1224,N_400);
nand U1701 (N_1701,N_1280,N_1319);
nand U1702 (N_1702,N_1175,N_1388);
and U1703 (N_1703,N_1265,N_210);
nand U1704 (N_1704,N_229,N_805);
or U1705 (N_1705,In_712,N_996);
nand U1706 (N_1706,N_293,In_2200);
xnor U1707 (N_1707,N_1255,In_472);
and U1708 (N_1708,N_1308,In_919);
and U1709 (N_1709,N_859,N_506);
nand U1710 (N_1710,N_1301,N_284);
and U1711 (N_1711,In_880,N_601);
xor U1712 (N_1712,N_220,N_1275);
nor U1713 (N_1713,N_1452,In_1798);
and U1714 (N_1714,N_767,N_353);
and U1715 (N_1715,In_2080,In_2367);
and U1716 (N_1716,N_314,N_754);
or U1717 (N_1717,In_101,N_1416);
xor U1718 (N_1718,N_431,In_1664);
or U1719 (N_1719,N_184,N_1410);
or U1720 (N_1720,N_968,In_477);
and U1721 (N_1721,In_1138,N_765);
nand U1722 (N_1722,In_1921,N_701);
nand U1723 (N_1723,N_1168,In_1278);
and U1724 (N_1724,N_413,N_1436);
nor U1725 (N_1725,N_1097,In_1925);
nor U1726 (N_1726,N_1064,N_1067);
nor U1727 (N_1727,N_1435,In_886);
nand U1728 (N_1728,N_1449,N_932);
nor U1729 (N_1729,N_1382,N_1078);
or U1730 (N_1730,N_538,In_1894);
or U1731 (N_1731,N_376,N_687);
or U1732 (N_1732,In_2243,N_1392);
or U1733 (N_1733,N_802,In_1028);
nand U1734 (N_1734,N_695,N_1411);
and U1735 (N_1735,N_1441,In_1366);
nor U1736 (N_1736,N_770,In_2190);
nor U1737 (N_1737,N_1089,In_92);
nor U1738 (N_1738,In_2329,N_1121);
or U1739 (N_1739,N_547,N_368);
or U1740 (N_1740,In_274,N_677);
and U1741 (N_1741,N_857,N_1488);
xor U1742 (N_1742,N_1477,N_1451);
nand U1743 (N_1743,In_1410,In_626);
or U1744 (N_1744,N_1354,In_1117);
and U1745 (N_1745,N_1467,N_398);
nor U1746 (N_1746,N_1066,In_1133);
nor U1747 (N_1747,N_1438,In_871);
and U1748 (N_1748,N_402,In_402);
nor U1749 (N_1749,In_844,N_1166);
and U1750 (N_1750,N_1626,N_1570);
or U1751 (N_1751,N_828,N_1721);
nor U1752 (N_1752,In_1120,N_630);
and U1753 (N_1753,N_1705,In_1340);
and U1754 (N_1754,N_1530,N_1709);
and U1755 (N_1755,In_1362,In_430);
and U1756 (N_1756,N_1512,In_936);
or U1757 (N_1757,N_1114,In_1773);
or U1758 (N_1758,In_2443,N_875);
nor U1759 (N_1759,In_1500,N_1270);
or U1760 (N_1760,In_539,N_1200);
nand U1761 (N_1761,N_567,In_62);
nand U1762 (N_1762,N_1728,N_505);
nor U1763 (N_1763,N_904,N_1342);
or U1764 (N_1764,N_946,N_1048);
nand U1765 (N_1765,N_1726,N_1718);
and U1766 (N_1766,N_563,N_1632);
or U1767 (N_1767,In_209,N_1325);
and U1768 (N_1768,N_1648,N_973);
or U1769 (N_1769,N_1565,N_827);
nor U1770 (N_1770,In_1683,N_1700);
and U1771 (N_1771,N_1117,N_1515);
or U1772 (N_1772,N_1105,N_1521);
nor U1773 (N_1773,N_1229,N_1704);
nand U1774 (N_1774,N_1458,N_1533);
nand U1775 (N_1775,N_1727,In_755);
nand U1776 (N_1776,N_1287,N_1465);
or U1777 (N_1777,N_94,In_2017);
nor U1778 (N_1778,N_1394,N_1672);
nor U1779 (N_1779,N_1698,N_339);
nor U1780 (N_1780,N_678,N_1296);
xor U1781 (N_1781,N_1579,N_1293);
and U1782 (N_1782,N_209,N_1725);
or U1783 (N_1783,In_1672,N_1719);
nand U1784 (N_1784,N_1126,N_1023);
and U1785 (N_1785,N_652,In_1722);
nand U1786 (N_1786,N_113,In_869);
and U1787 (N_1787,N_1691,In_1185);
or U1788 (N_1788,In_1380,N_1076);
nor U1789 (N_1789,N_1330,N_244);
nor U1790 (N_1790,N_1310,N_1210);
nor U1791 (N_1791,N_1359,In_1553);
or U1792 (N_1792,N_1582,In_2482);
or U1793 (N_1793,N_1538,N_1608);
nand U1794 (N_1794,N_1482,In_791);
and U1795 (N_1795,In_1132,N_1610);
nand U1796 (N_1796,N_1571,N_1694);
nand U1797 (N_1797,N_1055,N_1664);
nand U1798 (N_1798,N_927,N_1604);
nor U1799 (N_1799,N_1550,N_1030);
or U1800 (N_1800,N_1518,In_1421);
nand U1801 (N_1801,N_1074,N_1086);
or U1802 (N_1802,In_1069,N_1137);
nand U1803 (N_1803,N_728,In_1577);
nor U1804 (N_1804,N_1541,N_1283);
nor U1805 (N_1805,N_1600,N_1561);
and U1806 (N_1806,In_139,N_365);
nor U1807 (N_1807,In_1789,N_167);
nor U1808 (N_1808,N_1730,N_1371);
nand U1809 (N_1809,In_846,N_683);
or U1810 (N_1810,N_414,In_1);
xor U1811 (N_1811,N_1337,In_1810);
nand U1812 (N_1812,N_926,N_644);
nor U1813 (N_1813,In_175,In_1903);
or U1814 (N_1814,N_1513,In_1739);
nand U1815 (N_1815,N_1641,N_951);
nand U1816 (N_1816,N_1681,N_1507);
and U1817 (N_1817,N_1674,N_1511);
nand U1818 (N_1818,N_1689,N_1624);
xnor U1819 (N_1819,In_2324,N_1732);
or U1820 (N_1820,N_1334,N_1376);
and U1821 (N_1821,In_1994,In_1399);
or U1822 (N_1822,N_1450,N_811);
nand U1823 (N_1823,N_1746,N_1408);
or U1824 (N_1824,N_1396,N_1545);
nand U1825 (N_1825,In_1188,N_1655);
nand U1826 (N_1826,N_1712,In_658);
nor U1827 (N_1827,N_1206,N_429);
and U1828 (N_1828,N_935,N_1266);
nor U1829 (N_1829,N_1590,N_1542);
nor U1830 (N_1830,N_1514,In_1535);
or U1831 (N_1831,N_462,N_470);
nor U1832 (N_1832,N_1637,In_416);
and U1833 (N_1833,N_959,In_1434);
nand U1834 (N_1834,N_1623,N_1639);
nand U1835 (N_1835,N_1297,In_37);
xor U1836 (N_1836,N_1125,N_1568);
and U1837 (N_1837,In_1213,N_1081);
or U1838 (N_1838,N_1733,N_1673);
and U1839 (N_1839,N_1612,N_845);
xor U1840 (N_1840,N_1321,In_356);
and U1841 (N_1841,N_1688,N_1650);
or U1842 (N_1842,N_1536,N_800);
nand U1843 (N_1843,N_1627,In_1271);
xor U1844 (N_1844,In_103,In_831);
or U1845 (N_1845,In_1889,N_1358);
or U1846 (N_1846,N_1676,In_2172);
or U1847 (N_1847,N_1197,N_1431);
nor U1848 (N_1848,N_1406,N_1284);
and U1849 (N_1849,N_159,N_1107);
or U1850 (N_1850,N_1021,In_1093);
and U1851 (N_1851,N_527,N_1642);
xor U1852 (N_1852,N_1238,N_1257);
or U1853 (N_1853,N_1022,N_1596);
nand U1854 (N_1854,N_1448,In_2285);
nand U1855 (N_1855,In_1887,In_492);
or U1856 (N_1856,N_1666,N_1353);
nor U1857 (N_1857,N_984,N_1432);
xor U1858 (N_1858,N_1605,In_1076);
or U1859 (N_1859,N_1699,N_1569);
and U1860 (N_1860,N_1481,N_766);
and U1861 (N_1861,N_1096,N_1090);
nor U1862 (N_1862,N_1647,N_1649);
nor U1863 (N_1863,N_1462,N_518);
or U1864 (N_1864,N_889,N_1456);
or U1865 (N_1865,N_1615,In_2422);
nand U1866 (N_1866,N_1463,N_1095);
nand U1867 (N_1867,N_190,N_607);
or U1868 (N_1868,N_1690,N_1341);
and U1869 (N_1869,N_1322,In_137);
nand U1870 (N_1870,In_2252,N_1745);
nand U1871 (N_1871,N_1480,N_1269);
xnor U1872 (N_1872,N_1352,N_1136);
and U1873 (N_1873,In_571,N_1524);
nor U1874 (N_1874,N_1609,N_1747);
and U1875 (N_1875,N_818,N_910);
or U1876 (N_1876,N_1403,In_2124);
and U1877 (N_1877,N_1622,N_1583);
nand U1878 (N_1878,N_1303,N_1241);
or U1879 (N_1879,N_760,N_849);
or U1880 (N_1880,N_1340,In_1544);
nor U1881 (N_1881,N_1695,In_2450);
or U1882 (N_1882,N_1662,N_1585);
or U1883 (N_1883,N_1505,N_1598);
nand U1884 (N_1884,N_1540,N_1625);
nor U1885 (N_1885,N_681,N_1199);
and U1886 (N_1886,N_1678,In_1277);
or U1887 (N_1887,In_1361,N_1737);
nand U1888 (N_1888,N_1735,In_1575);
nor U1889 (N_1889,N_1263,N_1535);
xor U1890 (N_1890,N_333,N_1711);
and U1891 (N_1891,N_519,N_1307);
nor U1892 (N_1892,N_1621,N_1501);
and U1893 (N_1893,N_117,N_1716);
or U1894 (N_1894,In_1640,N_1271);
and U1895 (N_1895,N_1385,N_1309);
and U1896 (N_1896,In_1682,In_2398);
nor U1897 (N_1897,N_1597,N_1560);
nor U1898 (N_1898,In_1289,In_414);
or U1899 (N_1899,N_1591,N_417);
nor U1900 (N_1900,N_1528,N_1566);
xor U1901 (N_1901,N_1157,N_1425);
xor U1902 (N_1902,N_1552,In_581);
and U1903 (N_1903,N_1355,N_1555);
or U1904 (N_1904,In_406,N_703);
nand U1905 (N_1905,N_1232,N_1099);
or U1906 (N_1906,N_1669,N_1653);
and U1907 (N_1907,N_589,N_1559);
and U1908 (N_1908,N_821,N_1736);
nand U1909 (N_1909,In_1572,In_257);
nand U1910 (N_1910,N_1187,In_662);
nand U1911 (N_1911,In_1083,N_1279);
nor U1912 (N_1912,N_1070,N_1628);
or U1913 (N_1913,N_654,N_1049);
nand U1914 (N_1914,N_1317,N_1196);
and U1915 (N_1915,In_63,N_1119);
nand U1916 (N_1916,N_322,In_431);
nand U1917 (N_1917,N_1485,N_1742);
or U1918 (N_1918,N_1363,N_1413);
xnor U1919 (N_1919,N_643,N_853);
and U1920 (N_1920,In_1092,In_2227);
nand U1921 (N_1921,In_2105,N_1442);
or U1922 (N_1922,N_1602,N_1734);
nand U1923 (N_1923,N_16,N_1259);
and U1924 (N_1924,In_1780,In_2108);
nand U1925 (N_1925,N_1155,N_1654);
or U1926 (N_1926,N_1068,In_925);
and U1927 (N_1927,In_202,N_1658);
nor U1928 (N_1928,In_1412,N_1286);
xor U1929 (N_1929,N_1516,N_1478);
and U1930 (N_1930,N_1611,N_1492);
or U1931 (N_1931,N_465,N_1525);
and U1932 (N_1932,N_793,In_198);
and U1933 (N_1933,N_1033,N_1687);
nor U1934 (N_1934,In_2342,N_1717);
nor U1935 (N_1935,In_167,N_807);
nand U1936 (N_1936,N_1715,N_1075);
nand U1937 (N_1937,N_1724,N_1170);
or U1938 (N_1938,N_1373,N_1414);
or U1939 (N_1939,N_1466,N_1714);
or U1940 (N_1940,N_1262,N_1683);
nor U1941 (N_1941,N_1339,N_1276);
and U1942 (N_1942,N_848,N_1537);
nand U1943 (N_1943,N_1127,N_1577);
or U1944 (N_1944,N_1738,In_1851);
nor U1945 (N_1945,In_2078,N_247);
or U1946 (N_1946,N_460,N_1356);
or U1947 (N_1947,N_1381,N_1427);
nor U1948 (N_1948,N_595,N_1731);
nand U1949 (N_1949,N_1558,N_1003);
nor U1950 (N_1950,N_1188,N_831);
and U1951 (N_1951,In_1045,N_1667);
nand U1952 (N_1952,N_6,N_1060);
or U1953 (N_1953,In_644,N_1041);
xnor U1954 (N_1954,In_2493,N_1254);
or U1955 (N_1955,In_1917,In_1257);
nor U1956 (N_1956,N_1420,N_1520);
xor U1957 (N_1957,N_1305,In_1172);
nand U1958 (N_1958,N_1703,N_1680);
and U1959 (N_1959,N_1557,N_1179);
or U1960 (N_1960,N_1455,N_1748);
xnor U1961 (N_1961,N_1172,N_1014);
nor U1962 (N_1962,N_1722,N_1713);
nor U1963 (N_1963,N_983,In_1939);
and U1964 (N_1964,In_1872,N_397);
nand U1965 (N_1965,N_75,N_1372);
xnor U1966 (N_1966,N_993,N_485);
or U1967 (N_1967,N_1701,In_1377);
or U1968 (N_1968,N_929,In_2189);
nor U1969 (N_1969,N_1630,N_954);
nand U1970 (N_1970,N_1594,N_1222);
or U1971 (N_1971,In_1061,N_582);
nor U1972 (N_1972,In_1918,In_2018);
and U1973 (N_1973,N_1634,N_1572);
or U1974 (N_1974,N_1551,N_1029);
and U1975 (N_1975,N_745,N_1671);
nor U1976 (N_1976,N_1640,N_1743);
and U1977 (N_1977,N_1531,N_1696);
or U1978 (N_1978,N_1587,N_1013);
nand U1979 (N_1979,N_591,N_1405);
nor U1980 (N_1980,N_641,N_1380);
nand U1981 (N_1981,N_1225,N_1510);
xnor U1982 (N_1982,N_1468,N_791);
xnor U1983 (N_1983,In_1116,In_1962);
nand U1984 (N_1984,N_1025,In_1728);
xnor U1985 (N_1985,N_1331,N_1614);
or U1986 (N_1986,N_769,N_600);
or U1987 (N_1987,N_1710,N_907);
xnor U1988 (N_1988,In_690,N_924);
nand U1989 (N_1989,N_1682,N_1661);
or U1990 (N_1990,In_1548,N_1149);
nor U1991 (N_1991,N_1272,N_1261);
and U1992 (N_1992,N_1584,N_1684);
nor U1993 (N_1993,In_533,N_1633);
nor U1994 (N_1994,N_1295,N_1729);
xor U1995 (N_1995,In_1636,N_892);
nor U1996 (N_1996,In_1259,In_660);
or U1997 (N_1997,N_1506,N_1300);
and U1998 (N_1998,N_1589,N_234);
and U1999 (N_1999,N_228,N_846);
or U2000 (N_2000,N_1417,N_1668);
and U2001 (N_2001,N_507,N_1613);
or U2002 (N_2002,N_1997,N_1856);
nor U2003 (N_2003,N_1754,N_1998);
and U2004 (N_2004,N_1768,N_1502);
and U2005 (N_2005,N_1036,N_1757);
nor U2006 (N_2006,N_1900,N_1586);
nand U2007 (N_2007,N_1883,N_1947);
or U2008 (N_2008,N_1851,N_1783);
nand U2009 (N_2009,N_1046,N_788);
nor U2010 (N_2010,N_1969,N_1645);
nor U2011 (N_2011,N_1845,N_1799);
nor U2012 (N_2012,N_1539,N_1876);
or U2013 (N_2013,N_1885,N_700);
nand U2014 (N_2014,N_1213,N_1616);
or U2015 (N_2015,N_1122,N_1988);
and U2016 (N_2016,N_1464,N_1720);
or U2017 (N_2017,N_69,N_1220);
nand U2018 (N_2018,N_1974,N_1805);
and U2019 (N_2019,N_781,N_1834);
nand U2020 (N_2020,N_1460,N_1999);
and U2021 (N_2021,N_1758,N_1762);
nand U2022 (N_2022,N_1957,N_1978);
and U2023 (N_2023,N_1877,N_1926);
nand U2024 (N_2024,N_1901,N_1808);
nor U2025 (N_2025,N_1764,N_1504);
nand U2026 (N_2026,N_1774,In_199);
and U2027 (N_2027,N_1824,N_1332);
nor U2028 (N_2028,In_1830,N_1573);
nand U2029 (N_2029,N_1005,N_1795);
nand U2030 (N_2030,N_1809,N_1526);
or U2031 (N_2031,N_1894,In_1170);
nand U2032 (N_2032,N_1581,N_1941);
nand U2033 (N_2033,In_2447,N_1983);
nand U2034 (N_2034,N_1971,N_1606);
or U2035 (N_2035,N_1707,N_1943);
nor U2036 (N_2036,N_1702,N_1767);
or U2037 (N_2037,N_1846,N_1267);
xnor U2038 (N_2038,In_1456,N_1850);
or U2039 (N_2039,N_1828,N_1111);
xnor U2040 (N_2040,N_1787,In_2197);
and U2041 (N_2041,N_1867,N_1849);
nor U2042 (N_2042,N_1855,N_1951);
nor U2043 (N_2043,In_785,N_1818);
nand U2044 (N_2044,In_1526,N_1939);
xnor U2045 (N_2045,N_1091,N_1554);
nand U2046 (N_2046,N_1930,N_1844);
xor U2047 (N_2047,N_1904,N_1189);
or U2048 (N_2048,N_1899,N_1775);
or U2049 (N_2049,In_1634,In_2368);
xor U2050 (N_2050,N_18,N_1619);
nand U2051 (N_2051,N_1546,N_1553);
xnor U2052 (N_2052,In_2361,N_1183);
nand U2053 (N_2053,N_1852,N_753);
and U2054 (N_2054,N_1972,N_901);
or U2055 (N_2055,N_1990,N_883);
nor U2056 (N_2056,N_1929,In_510);
nor U2057 (N_2057,In_25,In_2181);
nor U2058 (N_2058,N_1154,N_1925);
and U2059 (N_2059,In_1118,N_899);
nor U2060 (N_2060,N_1875,N_1948);
and U2061 (N_2061,N_1306,N_1800);
and U2062 (N_2062,N_1796,N_1995);
nor U2063 (N_2063,N_1994,N_1486);
and U2064 (N_2064,N_1812,N_1870);
nand U2065 (N_2065,N_1895,N_1908);
nand U2066 (N_2066,N_1873,N_1932);
and U2067 (N_2067,N_1547,In_2396);
xor U2068 (N_2068,N_1891,N_1847);
nor U2069 (N_2069,N_604,N_1567);
or U2070 (N_2070,N_232,N_988);
or U2071 (N_2071,N_1918,N_1781);
or U2072 (N_2072,N_1970,N_407);
nand U2073 (N_2073,N_151,N_1741);
nand U2074 (N_2074,N_1863,N_311);
or U2075 (N_2075,N_1869,N_1996);
nand U2076 (N_2076,N_1786,N_1917);
nand U2077 (N_2077,N_798,N_1984);
xnor U2078 (N_2078,N_1804,N_1788);
or U2079 (N_2079,N_1910,N_1838);
or U2080 (N_2080,N_1752,N_1753);
or U2081 (N_2081,N_1440,N_1866);
and U2082 (N_2082,N_1791,N_1685);
or U2083 (N_2083,N_1360,N_1364);
nand U2084 (N_2084,In_2163,N_250);
nand U2085 (N_2085,N_1549,N_1989);
or U2086 (N_2086,N_208,N_1878);
nand U2087 (N_2087,In_768,N_1723);
or U2088 (N_2088,N_349,N_1407);
nor U2089 (N_2089,N_1840,N_1797);
nor U2090 (N_2090,N_1037,N_287);
nand U2091 (N_2091,N_1755,N_1927);
or U2092 (N_2092,N_1898,N_1208);
or U2093 (N_2093,N_1793,N_1909);
and U2094 (N_2094,N_1907,N_1770);
or U2095 (N_2095,N_1789,N_1740);
and U2096 (N_2096,N_1861,N_1914);
nand U2097 (N_2097,N_1836,N_1903);
xor U2098 (N_2098,N_1902,In_424);
nand U2099 (N_2099,N_1823,N_1476);
and U2100 (N_2100,N_1896,N_1693);
or U2101 (N_2101,N_1778,N_1811);
nor U2102 (N_2102,In_1474,N_513);
or U2103 (N_2103,N_1841,N_1500);
nand U2104 (N_2104,N_737,N_799);
nand U2105 (N_2105,N_1853,N_1643);
or U2106 (N_2106,N_1563,N_240);
nand U2107 (N_2107,N_1928,N_1198);
xnor U2108 (N_2108,N_1821,N_302);
and U2109 (N_2109,N_1487,N_1964);
and U2110 (N_2110,N_1950,N_1697);
and U2111 (N_2111,N_1780,N_1769);
nand U2112 (N_2112,N_1952,N_1979);
or U2113 (N_2113,N_1393,N_1350);
nand U2114 (N_2114,N_1635,N_1675);
and U2115 (N_2115,In_1122,N_1519);
xnor U2116 (N_2116,N_1859,N_1946);
nor U2117 (N_2117,In_214,N_1759);
nor U2118 (N_2118,N_1766,N_1985);
and U2119 (N_2119,N_1240,N_1285);
nand U2120 (N_2120,N_1825,N_1776);
nand U2121 (N_2121,N_1819,N_1889);
and U2122 (N_2122,N_1343,N_1813);
and U2123 (N_2123,N_1660,In_2184);
or U2124 (N_2124,N_1032,N_1593);
nand U2125 (N_2125,N_1858,N_1798);
or U2126 (N_2126,N_1912,N_1069);
nor U2127 (N_2127,N_1670,N_1888);
nand U2128 (N_2128,N_1792,N_1544);
and U2129 (N_2129,In_1318,N_1397);
xor U2130 (N_2130,N_1857,N_908);
or U2131 (N_2131,N_1976,N_608);
nor U2132 (N_2132,N_1588,N_1692);
nand U2133 (N_2133,N_1508,N_1084);
or U2134 (N_2134,N_68,N_1679);
nor U2135 (N_2135,In_2327,N_1865);
or U2136 (N_2136,N_1454,N_1469);
and U2137 (N_2137,N_1807,N_1966);
nand U2138 (N_2138,In_1690,N_1827);
nand U2139 (N_2139,N_1773,N_1802);
xor U2140 (N_2140,N_1794,N_1574);
and U2141 (N_2141,N_1522,N_1158);
nor U2142 (N_2142,N_1938,N_1936);
nor U2143 (N_2143,N_1871,In_901);
nor U2144 (N_2144,N_1312,N_1955);
and U2145 (N_2145,N_1517,N_1777);
and U2146 (N_2146,N_1592,N_1646);
xor U2147 (N_2147,N_1967,N_1527);
nor U2148 (N_2148,N_1578,N_1993);
and U2149 (N_2149,N_1881,N_1897);
nor U2150 (N_2150,N_1204,N_1879);
and U2151 (N_2151,N_1911,In_929);
or U2152 (N_2152,N_1651,N_1815);
nand U2153 (N_2153,N_1945,N_727);
or U2154 (N_2154,N_1784,N_1916);
nor U2155 (N_2155,N_1905,N_1923);
nor U2156 (N_2156,N_1618,In_1295);
and U2157 (N_2157,N_1933,N_1644);
xor U2158 (N_2158,N_1744,N_1657);
and U2159 (N_2159,N_1953,N_1595);
or U2160 (N_2160,N_1931,N_1772);
xor U2161 (N_2161,N_1315,N_1636);
and U2162 (N_2162,N_1806,N_1365);
or U2163 (N_2163,N_1503,N_1509);
nand U2164 (N_2164,N_1379,N_1782);
or U2165 (N_2165,N_1822,N_1543);
and U2166 (N_2166,N_1924,N_1874);
and U2167 (N_2167,N_1779,N_1765);
and U2168 (N_2168,N_1499,N_1471);
xor U2169 (N_2169,N_1832,N_1954);
nand U2170 (N_2170,N_873,N_1607);
or U2171 (N_2171,N_1810,N_1880);
nor U2172 (N_2172,N_1663,N_1826);
xor U2173 (N_2173,In_588,N_1790);
nor U2174 (N_2174,N_1962,In_906);
nor U2175 (N_2175,N_543,N_123);
nand U2176 (N_2176,N_1601,N_1906);
and U2177 (N_2177,N_1116,N_422);
or U2178 (N_2178,N_1652,N_1771);
nor U2179 (N_2179,In_462,N_1739);
or U2180 (N_2180,In_788,N_1638);
nand U2181 (N_2181,N_1991,N_1418);
and U2182 (N_2182,N_1816,N_606);
nor U2183 (N_2183,N_1835,N_1886);
and U2184 (N_2184,N_1751,N_1007);
nand U2185 (N_2185,N_1992,In_696);
nand U2186 (N_2186,N_1763,N_1884);
nand U2187 (N_2187,N_1575,N_1843);
nand U2188 (N_2188,N_1915,N_1934);
nand U2189 (N_2189,N_1921,N_1750);
nor U2190 (N_2190,N_809,N_1338);
nand U2191 (N_2191,N_758,N_1982);
nand U2192 (N_2192,N_1890,N_1961);
or U2193 (N_2193,In_816,N_838);
nor U2194 (N_2194,N_1801,In_1928);
nor U2195 (N_2195,N_1833,N_1603);
nand U2196 (N_2196,In_1740,N_1708);
and U2197 (N_2197,N_1920,N_1944);
xnor U2198 (N_2198,N_1706,N_297);
and U2199 (N_2199,N_502,In_1987);
xnor U2200 (N_2200,N_672,N_1576);
or U2201 (N_2201,N_813,N_1958);
nand U2202 (N_2202,N_1529,N_1803);
nand U2203 (N_2203,N_1665,N_1556);
nand U2204 (N_2204,N_1913,N_1523);
xnor U2205 (N_2205,N_1820,N_1629);
nor U2206 (N_2206,N_691,N_1756);
or U2207 (N_2207,N_1617,N_1548);
or U2208 (N_2208,N_1564,N_1760);
nor U2209 (N_2209,In_2492,N_1937);
nand U2210 (N_2210,N_1973,N_1935);
xor U2211 (N_2211,N_1968,N_1318);
xnor U2212 (N_2212,N_1831,N_1686);
or U2213 (N_2213,N_1963,N_1919);
xor U2214 (N_2214,N_1872,N_1631);
nand U2215 (N_2215,N_1860,N_1862);
or U2216 (N_2216,N_965,N_1854);
nand U2217 (N_2217,N_1659,N_1922);
and U2218 (N_2218,N_1940,N_1327);
nor U2219 (N_2219,N_1977,In_1355);
or U2220 (N_2220,N_1839,N_1177);
nand U2221 (N_2221,In_1732,N_1677);
nor U2222 (N_2222,N_1893,N_1956);
nor U2223 (N_2223,N_842,N_1842);
or U2224 (N_2224,N_1562,N_1532);
and U2225 (N_2225,N_1620,N_1599);
nor U2226 (N_2226,N_1959,N_1092);
or U2227 (N_2227,N_1164,N_426);
nor U2228 (N_2228,N_1311,N_1868);
nand U2229 (N_2229,N_1656,N_373);
nor U2230 (N_2230,N_1986,N_1987);
nand U2231 (N_2231,In_521,N_1837);
or U2232 (N_2232,N_1848,N_1965);
and U2233 (N_2233,N_1749,N_1830);
nor U2234 (N_2234,N_1942,N_1785);
nand U2235 (N_2235,N_1975,N_264);
or U2236 (N_2236,N_1534,N_484);
and U2237 (N_2237,N_1010,N_730);
nor U2238 (N_2238,N_1115,N_810);
nor U2239 (N_2239,N_1887,N_1329);
or U2240 (N_2240,N_1447,N_599);
and U2241 (N_2241,N_1113,N_1864);
nor U2242 (N_2242,N_1980,N_736);
and U2243 (N_2243,In_1435,N_1829);
or U2244 (N_2244,N_1949,N_1817);
nand U2245 (N_2245,N_1761,N_1016);
nand U2246 (N_2246,N_1981,N_1892);
and U2247 (N_2247,N_514,N_1814);
nor U2248 (N_2248,N_1580,N_1073);
nor U2249 (N_2249,N_1882,N_1960);
xor U2250 (N_2250,N_2179,N_2074);
nand U2251 (N_2251,N_2029,N_2107);
nor U2252 (N_2252,N_2161,N_2227);
xor U2253 (N_2253,N_2061,N_2109);
nor U2254 (N_2254,N_2019,N_2209);
or U2255 (N_2255,N_2197,N_2015);
nand U2256 (N_2256,N_2073,N_2186);
xor U2257 (N_2257,N_2068,N_2177);
and U2258 (N_2258,N_2143,N_2136);
nor U2259 (N_2259,N_2009,N_2016);
or U2260 (N_2260,N_2071,N_2167);
nand U2261 (N_2261,N_2024,N_2121);
and U2262 (N_2262,N_2156,N_2183);
nand U2263 (N_2263,N_2021,N_2214);
and U2264 (N_2264,N_2118,N_2044);
or U2265 (N_2265,N_2105,N_2081);
nand U2266 (N_2266,N_2211,N_2224);
nor U2267 (N_2267,N_2028,N_2228);
and U2268 (N_2268,N_2083,N_2114);
nor U2269 (N_2269,N_2180,N_2087);
or U2270 (N_2270,N_2023,N_2100);
nor U2271 (N_2271,N_2160,N_2047);
nand U2272 (N_2272,N_2150,N_2003);
nand U2273 (N_2273,N_2201,N_2056);
xor U2274 (N_2274,N_2146,N_2172);
and U2275 (N_2275,N_2220,N_2088);
and U2276 (N_2276,N_2244,N_2005);
nand U2277 (N_2277,N_2122,N_2090);
nand U2278 (N_2278,N_2207,N_2239);
nor U2279 (N_2279,N_2093,N_2216);
and U2280 (N_2280,N_2240,N_2153);
or U2281 (N_2281,N_2165,N_2010);
or U2282 (N_2282,N_2147,N_2219);
and U2283 (N_2283,N_2135,N_2204);
nor U2284 (N_2284,N_2098,N_2069);
and U2285 (N_2285,N_2189,N_2158);
and U2286 (N_2286,N_2119,N_2092);
or U2287 (N_2287,N_2238,N_2134);
nor U2288 (N_2288,N_2064,N_2110);
and U2289 (N_2289,N_2234,N_2140);
nor U2290 (N_2290,N_2006,N_2163);
and U2291 (N_2291,N_2085,N_2062);
or U2292 (N_2292,N_2182,N_2013);
xor U2293 (N_2293,N_2039,N_2001);
and U2294 (N_2294,N_2196,N_2187);
and U2295 (N_2295,N_2067,N_2106);
and U2296 (N_2296,N_2034,N_2116);
xor U2297 (N_2297,N_2066,N_2011);
nand U2298 (N_2298,N_2195,N_2155);
nor U2299 (N_2299,N_2082,N_2203);
nand U2300 (N_2300,N_2157,N_2049);
and U2301 (N_2301,N_2117,N_2230);
nand U2302 (N_2302,N_2149,N_2101);
nand U2303 (N_2303,N_2038,N_2032);
or U2304 (N_2304,N_2128,N_2170);
or U2305 (N_2305,N_2113,N_2070);
or U2306 (N_2306,N_2036,N_2089);
and U2307 (N_2307,N_2248,N_2226);
nor U2308 (N_2308,N_2137,N_2190);
and U2309 (N_2309,N_2014,N_2022);
xnor U2310 (N_2310,N_2169,N_2027);
nand U2311 (N_2311,N_2102,N_2017);
nand U2312 (N_2312,N_2030,N_2237);
or U2313 (N_2313,N_2052,N_2046);
or U2314 (N_2314,N_2151,N_2096);
xor U2315 (N_2315,N_2188,N_2130);
nand U2316 (N_2316,N_2141,N_2075);
and U2317 (N_2317,N_2041,N_2176);
and U2318 (N_2318,N_2205,N_2144);
nand U2319 (N_2319,N_2051,N_2040);
xnor U2320 (N_2320,N_2080,N_2037);
or U2321 (N_2321,N_2111,N_2063);
or U2322 (N_2322,N_2054,N_2020);
nand U2323 (N_2323,N_2164,N_2221);
and U2324 (N_2324,N_2095,N_2104);
nand U2325 (N_2325,N_2000,N_2139);
nor U2326 (N_2326,N_2133,N_2200);
nor U2327 (N_2327,N_2231,N_2241);
or U2328 (N_2328,N_2159,N_2191);
and U2329 (N_2329,N_2076,N_2175);
and U2330 (N_2330,N_2152,N_2242);
nand U2331 (N_2331,N_2232,N_2249);
nand U2332 (N_2332,N_2112,N_2060);
or U2333 (N_2333,N_2126,N_2091);
and U2334 (N_2334,N_2086,N_2045);
xnor U2335 (N_2335,N_2131,N_2192);
or U2336 (N_2336,N_2129,N_2185);
and U2337 (N_2337,N_2184,N_2178);
nand U2338 (N_2338,N_2043,N_2138);
and U2339 (N_2339,N_2078,N_2168);
and U2340 (N_2340,N_2053,N_2245);
and U2341 (N_2341,N_2198,N_2099);
nand U2342 (N_2342,N_2025,N_2142);
and U2343 (N_2343,N_2035,N_2145);
or U2344 (N_2344,N_2193,N_2057);
xor U2345 (N_2345,N_2103,N_2199);
nor U2346 (N_2346,N_2072,N_2213);
xor U2347 (N_2347,N_2018,N_2115);
nor U2348 (N_2348,N_2065,N_2222);
nand U2349 (N_2349,N_2059,N_2246);
and U2350 (N_2350,N_2123,N_2055);
nand U2351 (N_2351,N_2174,N_2132);
nor U2352 (N_2352,N_2166,N_2004);
nand U2353 (N_2353,N_2026,N_2148);
nor U2354 (N_2354,N_2127,N_2181);
nand U2355 (N_2355,N_2007,N_2084);
or U2356 (N_2356,N_2050,N_2079);
or U2357 (N_2357,N_2173,N_2002);
nand U2358 (N_2358,N_2108,N_2218);
or U2359 (N_2359,N_2058,N_2217);
and U2360 (N_2360,N_2154,N_2077);
nand U2361 (N_2361,N_2031,N_2210);
or U2362 (N_2362,N_2233,N_2223);
xnor U2363 (N_2363,N_2012,N_2008);
and U2364 (N_2364,N_2243,N_2208);
and U2365 (N_2365,N_2162,N_2048);
xor U2366 (N_2366,N_2212,N_2120);
and U2367 (N_2367,N_2235,N_2033);
and U2368 (N_2368,N_2215,N_2097);
and U2369 (N_2369,N_2094,N_2125);
and U2370 (N_2370,N_2042,N_2236);
nor U2371 (N_2371,N_2124,N_2247);
nor U2372 (N_2372,N_2194,N_2171);
nand U2373 (N_2373,N_2225,N_2202);
nand U2374 (N_2374,N_2229,N_2206);
nor U2375 (N_2375,N_2040,N_2128);
or U2376 (N_2376,N_2145,N_2201);
xor U2377 (N_2377,N_2087,N_2214);
nor U2378 (N_2378,N_2143,N_2241);
nor U2379 (N_2379,N_2037,N_2059);
nor U2380 (N_2380,N_2031,N_2061);
or U2381 (N_2381,N_2103,N_2030);
xor U2382 (N_2382,N_2166,N_2027);
nand U2383 (N_2383,N_2102,N_2223);
or U2384 (N_2384,N_2119,N_2167);
nor U2385 (N_2385,N_2166,N_2209);
and U2386 (N_2386,N_2143,N_2150);
nor U2387 (N_2387,N_2003,N_2171);
nor U2388 (N_2388,N_2118,N_2229);
nand U2389 (N_2389,N_2085,N_2223);
xor U2390 (N_2390,N_2145,N_2042);
nand U2391 (N_2391,N_2115,N_2210);
nor U2392 (N_2392,N_2083,N_2089);
and U2393 (N_2393,N_2055,N_2011);
nand U2394 (N_2394,N_2175,N_2014);
nor U2395 (N_2395,N_2201,N_2069);
and U2396 (N_2396,N_2031,N_2127);
or U2397 (N_2397,N_2048,N_2167);
or U2398 (N_2398,N_2159,N_2128);
or U2399 (N_2399,N_2000,N_2072);
and U2400 (N_2400,N_2172,N_2095);
nor U2401 (N_2401,N_2053,N_2137);
nor U2402 (N_2402,N_2090,N_2114);
or U2403 (N_2403,N_2060,N_2247);
nand U2404 (N_2404,N_2082,N_2174);
nand U2405 (N_2405,N_2099,N_2200);
xnor U2406 (N_2406,N_2140,N_2177);
and U2407 (N_2407,N_2132,N_2162);
xor U2408 (N_2408,N_2037,N_2223);
nor U2409 (N_2409,N_2083,N_2235);
nand U2410 (N_2410,N_2103,N_2015);
nor U2411 (N_2411,N_2222,N_2074);
nor U2412 (N_2412,N_2059,N_2175);
and U2413 (N_2413,N_2026,N_2106);
or U2414 (N_2414,N_2127,N_2008);
or U2415 (N_2415,N_2214,N_2228);
nand U2416 (N_2416,N_2208,N_2044);
nand U2417 (N_2417,N_2227,N_2185);
and U2418 (N_2418,N_2181,N_2214);
nand U2419 (N_2419,N_2242,N_2234);
or U2420 (N_2420,N_2172,N_2140);
nor U2421 (N_2421,N_2170,N_2209);
xnor U2422 (N_2422,N_2177,N_2207);
xnor U2423 (N_2423,N_2014,N_2045);
or U2424 (N_2424,N_2092,N_2167);
nand U2425 (N_2425,N_2203,N_2008);
nand U2426 (N_2426,N_2215,N_2007);
or U2427 (N_2427,N_2024,N_2082);
or U2428 (N_2428,N_2183,N_2212);
nor U2429 (N_2429,N_2105,N_2178);
nand U2430 (N_2430,N_2091,N_2048);
nand U2431 (N_2431,N_2205,N_2219);
or U2432 (N_2432,N_2062,N_2120);
or U2433 (N_2433,N_2088,N_2155);
nor U2434 (N_2434,N_2220,N_2120);
nor U2435 (N_2435,N_2014,N_2217);
nand U2436 (N_2436,N_2229,N_2084);
nor U2437 (N_2437,N_2060,N_2081);
and U2438 (N_2438,N_2024,N_2045);
nor U2439 (N_2439,N_2125,N_2087);
xor U2440 (N_2440,N_2183,N_2025);
and U2441 (N_2441,N_2074,N_2024);
or U2442 (N_2442,N_2166,N_2144);
and U2443 (N_2443,N_2098,N_2113);
nor U2444 (N_2444,N_2121,N_2010);
and U2445 (N_2445,N_2032,N_2093);
or U2446 (N_2446,N_2204,N_2237);
and U2447 (N_2447,N_2103,N_2075);
nand U2448 (N_2448,N_2191,N_2156);
nand U2449 (N_2449,N_2150,N_2228);
nand U2450 (N_2450,N_2114,N_2202);
nand U2451 (N_2451,N_2117,N_2000);
nor U2452 (N_2452,N_2166,N_2121);
nor U2453 (N_2453,N_2151,N_2089);
nand U2454 (N_2454,N_2050,N_2160);
and U2455 (N_2455,N_2042,N_2043);
or U2456 (N_2456,N_2073,N_2156);
and U2457 (N_2457,N_2048,N_2208);
nor U2458 (N_2458,N_2242,N_2062);
or U2459 (N_2459,N_2077,N_2020);
nor U2460 (N_2460,N_2020,N_2165);
or U2461 (N_2461,N_2050,N_2172);
or U2462 (N_2462,N_2137,N_2149);
and U2463 (N_2463,N_2141,N_2179);
nor U2464 (N_2464,N_2114,N_2157);
nand U2465 (N_2465,N_2053,N_2110);
and U2466 (N_2466,N_2064,N_2059);
or U2467 (N_2467,N_2213,N_2113);
xnor U2468 (N_2468,N_2048,N_2076);
or U2469 (N_2469,N_2186,N_2058);
nand U2470 (N_2470,N_2083,N_2084);
or U2471 (N_2471,N_2073,N_2070);
nand U2472 (N_2472,N_2044,N_2085);
nand U2473 (N_2473,N_2133,N_2213);
nor U2474 (N_2474,N_2088,N_2233);
nand U2475 (N_2475,N_2126,N_2068);
or U2476 (N_2476,N_2166,N_2179);
and U2477 (N_2477,N_2218,N_2001);
and U2478 (N_2478,N_2124,N_2198);
and U2479 (N_2479,N_2138,N_2062);
xnor U2480 (N_2480,N_2248,N_2246);
or U2481 (N_2481,N_2141,N_2140);
nor U2482 (N_2482,N_2151,N_2024);
or U2483 (N_2483,N_2081,N_2087);
and U2484 (N_2484,N_2015,N_2037);
and U2485 (N_2485,N_2049,N_2034);
nand U2486 (N_2486,N_2091,N_2196);
or U2487 (N_2487,N_2223,N_2011);
or U2488 (N_2488,N_2171,N_2137);
or U2489 (N_2489,N_2121,N_2049);
and U2490 (N_2490,N_2181,N_2104);
nand U2491 (N_2491,N_2137,N_2033);
and U2492 (N_2492,N_2038,N_2245);
and U2493 (N_2493,N_2214,N_2011);
or U2494 (N_2494,N_2201,N_2130);
nor U2495 (N_2495,N_2171,N_2157);
or U2496 (N_2496,N_2116,N_2085);
nor U2497 (N_2497,N_2190,N_2104);
or U2498 (N_2498,N_2067,N_2071);
nand U2499 (N_2499,N_2124,N_2069);
and U2500 (N_2500,N_2284,N_2325);
and U2501 (N_2501,N_2471,N_2440);
nor U2502 (N_2502,N_2361,N_2420);
or U2503 (N_2503,N_2289,N_2391);
nor U2504 (N_2504,N_2334,N_2276);
and U2505 (N_2505,N_2435,N_2388);
and U2506 (N_2506,N_2465,N_2343);
or U2507 (N_2507,N_2485,N_2404);
nor U2508 (N_2508,N_2381,N_2346);
nor U2509 (N_2509,N_2429,N_2487);
and U2510 (N_2510,N_2492,N_2446);
nor U2511 (N_2511,N_2432,N_2396);
nand U2512 (N_2512,N_2384,N_2287);
or U2513 (N_2513,N_2433,N_2356);
nor U2514 (N_2514,N_2459,N_2374);
and U2515 (N_2515,N_2299,N_2430);
nor U2516 (N_2516,N_2498,N_2401);
nand U2517 (N_2517,N_2417,N_2392);
or U2518 (N_2518,N_2320,N_2257);
nand U2519 (N_2519,N_2281,N_2264);
nor U2520 (N_2520,N_2300,N_2321);
nand U2521 (N_2521,N_2315,N_2260);
nand U2522 (N_2522,N_2378,N_2395);
nand U2523 (N_2523,N_2274,N_2479);
or U2524 (N_2524,N_2478,N_2473);
nand U2525 (N_2525,N_2372,N_2453);
or U2526 (N_2526,N_2326,N_2493);
nor U2527 (N_2527,N_2332,N_2458);
xor U2528 (N_2528,N_2288,N_2428);
nand U2529 (N_2529,N_2328,N_2421);
and U2530 (N_2530,N_2385,N_2292);
nor U2531 (N_2531,N_2387,N_2296);
xnor U2532 (N_2532,N_2301,N_2383);
and U2533 (N_2533,N_2280,N_2489);
nor U2534 (N_2534,N_2450,N_2494);
xnor U2535 (N_2535,N_2317,N_2483);
or U2536 (N_2536,N_2357,N_2336);
and U2537 (N_2537,N_2393,N_2291);
and U2538 (N_2538,N_2386,N_2457);
and U2539 (N_2539,N_2297,N_2303);
nor U2540 (N_2540,N_2347,N_2394);
nor U2541 (N_2541,N_2345,N_2362);
nor U2542 (N_2542,N_2273,N_2363);
and U2543 (N_2543,N_2255,N_2348);
nand U2544 (N_2544,N_2431,N_2376);
xor U2545 (N_2545,N_2298,N_2414);
nand U2546 (N_2546,N_2360,N_2278);
and U2547 (N_2547,N_2262,N_2309);
and U2548 (N_2548,N_2382,N_2466);
nor U2549 (N_2549,N_2438,N_2412);
nor U2550 (N_2550,N_2495,N_2441);
and U2551 (N_2551,N_2250,N_2472);
nor U2552 (N_2552,N_2474,N_2481);
nand U2553 (N_2553,N_2369,N_2377);
or U2554 (N_2554,N_2469,N_2364);
or U2555 (N_2555,N_2444,N_2439);
and U2556 (N_2556,N_2259,N_2454);
nand U2557 (N_2557,N_2285,N_2352);
or U2558 (N_2558,N_2290,N_2355);
or U2559 (N_2559,N_2305,N_2482);
and U2560 (N_2560,N_2442,N_2366);
or U2561 (N_2561,N_2310,N_2252);
xnor U2562 (N_2562,N_2316,N_2497);
and U2563 (N_2563,N_2415,N_2426);
nand U2564 (N_2564,N_2451,N_2476);
nor U2565 (N_2565,N_2283,N_2452);
xnor U2566 (N_2566,N_2409,N_2413);
nand U2567 (N_2567,N_2354,N_2330);
or U2568 (N_2568,N_2389,N_2256);
or U2569 (N_2569,N_2323,N_2486);
nor U2570 (N_2570,N_2445,N_2265);
or U2571 (N_2571,N_2258,N_2272);
and U2572 (N_2572,N_2405,N_2277);
or U2573 (N_2573,N_2335,N_2302);
and U2574 (N_2574,N_2436,N_2324);
and U2575 (N_2575,N_2367,N_2403);
nand U2576 (N_2576,N_2496,N_2267);
nand U2577 (N_2577,N_2398,N_2279);
or U2578 (N_2578,N_2397,N_2339);
nor U2579 (N_2579,N_2340,N_2411);
and U2580 (N_2580,N_2418,N_2477);
nor U2581 (N_2581,N_2268,N_2447);
nor U2582 (N_2582,N_2353,N_2344);
and U2583 (N_2583,N_2307,N_2434);
and U2584 (N_2584,N_2308,N_2448);
and U2585 (N_2585,N_2464,N_2311);
and U2586 (N_2586,N_2375,N_2449);
and U2587 (N_2587,N_2271,N_2419);
nor U2588 (N_2588,N_2251,N_2312);
and U2589 (N_2589,N_2400,N_2463);
nor U2590 (N_2590,N_2304,N_2484);
nor U2591 (N_2591,N_2314,N_2365);
nand U2592 (N_2592,N_2318,N_2253);
and U2593 (N_2593,N_2480,N_2390);
nor U2594 (N_2594,N_2406,N_2468);
xor U2595 (N_2595,N_2293,N_2488);
nor U2596 (N_2596,N_2349,N_2270);
nand U2597 (N_2597,N_2410,N_2266);
xnor U2598 (N_2598,N_2461,N_2467);
nor U2599 (N_2599,N_2313,N_2416);
or U2600 (N_2600,N_2424,N_2373);
or U2601 (N_2601,N_2423,N_2342);
nand U2602 (N_2602,N_2456,N_2380);
and U2603 (N_2603,N_2425,N_2261);
nand U2604 (N_2604,N_2269,N_2370);
or U2605 (N_2605,N_2358,N_2333);
or U2606 (N_2606,N_2350,N_2338);
and U2607 (N_2607,N_2408,N_2371);
nor U2608 (N_2608,N_2402,N_2407);
and U2609 (N_2609,N_2306,N_2399);
or U2610 (N_2610,N_2275,N_2368);
nand U2611 (N_2611,N_2329,N_2254);
or U2612 (N_2612,N_2490,N_2475);
xnor U2613 (N_2613,N_2379,N_2455);
nand U2614 (N_2614,N_2331,N_2422);
xor U2615 (N_2615,N_2286,N_2294);
nand U2616 (N_2616,N_2341,N_2282);
nand U2617 (N_2617,N_2319,N_2295);
or U2618 (N_2618,N_2499,N_2437);
and U2619 (N_2619,N_2427,N_2351);
or U2620 (N_2620,N_2359,N_2322);
and U2621 (N_2621,N_2460,N_2462);
and U2622 (N_2622,N_2443,N_2263);
or U2623 (N_2623,N_2470,N_2327);
nor U2624 (N_2624,N_2337,N_2491);
and U2625 (N_2625,N_2472,N_2306);
nor U2626 (N_2626,N_2255,N_2471);
or U2627 (N_2627,N_2460,N_2385);
nand U2628 (N_2628,N_2280,N_2351);
nor U2629 (N_2629,N_2445,N_2335);
and U2630 (N_2630,N_2371,N_2312);
nand U2631 (N_2631,N_2415,N_2368);
xnor U2632 (N_2632,N_2468,N_2382);
xnor U2633 (N_2633,N_2448,N_2311);
or U2634 (N_2634,N_2496,N_2404);
and U2635 (N_2635,N_2429,N_2256);
and U2636 (N_2636,N_2324,N_2318);
or U2637 (N_2637,N_2486,N_2459);
and U2638 (N_2638,N_2360,N_2382);
or U2639 (N_2639,N_2429,N_2455);
xnor U2640 (N_2640,N_2260,N_2263);
nand U2641 (N_2641,N_2453,N_2251);
nand U2642 (N_2642,N_2254,N_2454);
nor U2643 (N_2643,N_2451,N_2427);
and U2644 (N_2644,N_2335,N_2347);
or U2645 (N_2645,N_2408,N_2363);
nand U2646 (N_2646,N_2355,N_2294);
xnor U2647 (N_2647,N_2395,N_2269);
or U2648 (N_2648,N_2267,N_2435);
nand U2649 (N_2649,N_2338,N_2375);
or U2650 (N_2650,N_2360,N_2261);
nor U2651 (N_2651,N_2324,N_2462);
nor U2652 (N_2652,N_2492,N_2470);
nand U2653 (N_2653,N_2267,N_2293);
or U2654 (N_2654,N_2353,N_2347);
nor U2655 (N_2655,N_2402,N_2322);
nand U2656 (N_2656,N_2268,N_2458);
nand U2657 (N_2657,N_2455,N_2418);
xor U2658 (N_2658,N_2387,N_2394);
or U2659 (N_2659,N_2339,N_2309);
nand U2660 (N_2660,N_2346,N_2367);
or U2661 (N_2661,N_2365,N_2398);
or U2662 (N_2662,N_2489,N_2403);
xnor U2663 (N_2663,N_2305,N_2456);
nand U2664 (N_2664,N_2331,N_2426);
nand U2665 (N_2665,N_2419,N_2445);
or U2666 (N_2666,N_2496,N_2259);
nor U2667 (N_2667,N_2333,N_2293);
or U2668 (N_2668,N_2297,N_2285);
nand U2669 (N_2669,N_2476,N_2456);
and U2670 (N_2670,N_2337,N_2417);
and U2671 (N_2671,N_2313,N_2415);
nor U2672 (N_2672,N_2464,N_2421);
nor U2673 (N_2673,N_2430,N_2490);
nand U2674 (N_2674,N_2351,N_2278);
and U2675 (N_2675,N_2362,N_2413);
nor U2676 (N_2676,N_2448,N_2299);
xnor U2677 (N_2677,N_2325,N_2411);
or U2678 (N_2678,N_2299,N_2260);
and U2679 (N_2679,N_2258,N_2349);
and U2680 (N_2680,N_2449,N_2317);
nand U2681 (N_2681,N_2427,N_2449);
or U2682 (N_2682,N_2364,N_2351);
and U2683 (N_2683,N_2321,N_2473);
or U2684 (N_2684,N_2440,N_2431);
and U2685 (N_2685,N_2282,N_2262);
or U2686 (N_2686,N_2263,N_2336);
or U2687 (N_2687,N_2255,N_2379);
or U2688 (N_2688,N_2485,N_2336);
and U2689 (N_2689,N_2415,N_2316);
nand U2690 (N_2690,N_2399,N_2490);
and U2691 (N_2691,N_2264,N_2274);
or U2692 (N_2692,N_2485,N_2446);
nor U2693 (N_2693,N_2399,N_2345);
or U2694 (N_2694,N_2400,N_2371);
and U2695 (N_2695,N_2411,N_2289);
and U2696 (N_2696,N_2372,N_2332);
nand U2697 (N_2697,N_2406,N_2378);
nand U2698 (N_2698,N_2421,N_2315);
or U2699 (N_2699,N_2471,N_2337);
nor U2700 (N_2700,N_2302,N_2498);
nor U2701 (N_2701,N_2459,N_2381);
or U2702 (N_2702,N_2481,N_2269);
and U2703 (N_2703,N_2340,N_2252);
and U2704 (N_2704,N_2499,N_2416);
nor U2705 (N_2705,N_2471,N_2412);
or U2706 (N_2706,N_2332,N_2370);
nand U2707 (N_2707,N_2302,N_2485);
and U2708 (N_2708,N_2345,N_2426);
nor U2709 (N_2709,N_2430,N_2330);
and U2710 (N_2710,N_2258,N_2392);
nor U2711 (N_2711,N_2415,N_2439);
xor U2712 (N_2712,N_2406,N_2467);
xor U2713 (N_2713,N_2326,N_2396);
nor U2714 (N_2714,N_2287,N_2483);
nor U2715 (N_2715,N_2458,N_2387);
nand U2716 (N_2716,N_2441,N_2372);
xnor U2717 (N_2717,N_2382,N_2368);
xor U2718 (N_2718,N_2328,N_2263);
nand U2719 (N_2719,N_2491,N_2406);
nor U2720 (N_2720,N_2300,N_2330);
or U2721 (N_2721,N_2441,N_2488);
or U2722 (N_2722,N_2463,N_2341);
nor U2723 (N_2723,N_2460,N_2394);
or U2724 (N_2724,N_2466,N_2287);
and U2725 (N_2725,N_2399,N_2317);
nor U2726 (N_2726,N_2284,N_2452);
or U2727 (N_2727,N_2490,N_2497);
and U2728 (N_2728,N_2346,N_2401);
and U2729 (N_2729,N_2253,N_2259);
and U2730 (N_2730,N_2478,N_2364);
xnor U2731 (N_2731,N_2435,N_2309);
nor U2732 (N_2732,N_2291,N_2256);
or U2733 (N_2733,N_2445,N_2472);
and U2734 (N_2734,N_2323,N_2459);
or U2735 (N_2735,N_2269,N_2393);
xor U2736 (N_2736,N_2279,N_2322);
and U2737 (N_2737,N_2365,N_2449);
nand U2738 (N_2738,N_2402,N_2499);
or U2739 (N_2739,N_2435,N_2360);
nor U2740 (N_2740,N_2488,N_2391);
xnor U2741 (N_2741,N_2258,N_2326);
and U2742 (N_2742,N_2396,N_2417);
nand U2743 (N_2743,N_2344,N_2485);
xnor U2744 (N_2744,N_2372,N_2274);
nand U2745 (N_2745,N_2378,N_2262);
and U2746 (N_2746,N_2427,N_2384);
nor U2747 (N_2747,N_2300,N_2475);
or U2748 (N_2748,N_2392,N_2472);
or U2749 (N_2749,N_2473,N_2370);
and U2750 (N_2750,N_2516,N_2677);
nand U2751 (N_2751,N_2679,N_2571);
nand U2752 (N_2752,N_2712,N_2504);
nand U2753 (N_2753,N_2724,N_2729);
nor U2754 (N_2754,N_2664,N_2593);
and U2755 (N_2755,N_2613,N_2601);
nand U2756 (N_2756,N_2596,N_2718);
nand U2757 (N_2757,N_2536,N_2542);
or U2758 (N_2758,N_2628,N_2534);
nand U2759 (N_2759,N_2731,N_2708);
nor U2760 (N_2760,N_2735,N_2649);
or U2761 (N_2761,N_2556,N_2739);
and U2762 (N_2762,N_2698,N_2555);
xnor U2763 (N_2763,N_2558,N_2627);
nand U2764 (N_2764,N_2560,N_2624);
nor U2765 (N_2765,N_2648,N_2513);
xnor U2766 (N_2766,N_2654,N_2551);
and U2767 (N_2767,N_2573,N_2579);
and U2768 (N_2768,N_2709,N_2638);
or U2769 (N_2769,N_2687,N_2655);
nand U2770 (N_2770,N_2642,N_2727);
xnor U2771 (N_2771,N_2612,N_2572);
nor U2772 (N_2772,N_2584,N_2583);
or U2773 (N_2773,N_2692,N_2671);
nand U2774 (N_2774,N_2725,N_2641);
xor U2775 (N_2775,N_2640,N_2635);
nor U2776 (N_2776,N_2650,N_2524);
nor U2777 (N_2777,N_2645,N_2566);
or U2778 (N_2778,N_2744,N_2651);
nor U2779 (N_2779,N_2505,N_2631);
nand U2780 (N_2780,N_2552,N_2569);
and U2781 (N_2781,N_2738,N_2644);
nor U2782 (N_2782,N_2723,N_2512);
nand U2783 (N_2783,N_2716,N_2599);
nor U2784 (N_2784,N_2678,N_2511);
nand U2785 (N_2785,N_2539,N_2674);
or U2786 (N_2786,N_2538,N_2515);
nand U2787 (N_2787,N_2694,N_2529);
and U2788 (N_2788,N_2587,N_2608);
xor U2789 (N_2789,N_2656,N_2549);
nor U2790 (N_2790,N_2637,N_2730);
and U2791 (N_2791,N_2726,N_2706);
and U2792 (N_2792,N_2563,N_2682);
nand U2793 (N_2793,N_2688,N_2592);
nand U2794 (N_2794,N_2745,N_2672);
xor U2795 (N_2795,N_2620,N_2550);
nand U2796 (N_2796,N_2728,N_2585);
and U2797 (N_2797,N_2531,N_2606);
nand U2798 (N_2798,N_2575,N_2622);
nand U2799 (N_2799,N_2600,N_2561);
nand U2800 (N_2800,N_2553,N_2567);
nor U2801 (N_2801,N_2615,N_2673);
and U2802 (N_2802,N_2713,N_2721);
or U2803 (N_2803,N_2625,N_2665);
or U2804 (N_2804,N_2697,N_2522);
and U2805 (N_2805,N_2506,N_2736);
or U2806 (N_2806,N_2733,N_2541);
and U2807 (N_2807,N_2710,N_2748);
or U2808 (N_2808,N_2702,N_2604);
nand U2809 (N_2809,N_2746,N_2545);
nor U2810 (N_2810,N_2720,N_2670);
and U2811 (N_2811,N_2707,N_2557);
nor U2812 (N_2812,N_2686,N_2737);
xnor U2813 (N_2813,N_2619,N_2684);
and U2814 (N_2814,N_2714,N_2594);
nor U2815 (N_2815,N_2500,N_2740);
nand U2816 (N_2816,N_2582,N_2581);
and U2817 (N_2817,N_2732,N_2660);
nand U2818 (N_2818,N_2667,N_2704);
xnor U2819 (N_2819,N_2653,N_2646);
and U2820 (N_2820,N_2652,N_2680);
nand U2821 (N_2821,N_2501,N_2546);
nor U2822 (N_2822,N_2683,N_2611);
nor U2823 (N_2823,N_2547,N_2701);
nand U2824 (N_2824,N_2564,N_2617);
and U2825 (N_2825,N_2526,N_2562);
and U2826 (N_2826,N_2554,N_2548);
nand U2827 (N_2827,N_2630,N_2633);
or U2828 (N_2828,N_2609,N_2603);
or U2829 (N_2829,N_2540,N_2577);
nor U2830 (N_2830,N_2634,N_2528);
and U2831 (N_2831,N_2743,N_2568);
nand U2832 (N_2832,N_2711,N_2703);
nand U2833 (N_2833,N_2605,N_2508);
or U2834 (N_2834,N_2636,N_2741);
nand U2835 (N_2835,N_2537,N_2700);
nor U2836 (N_2836,N_2742,N_2695);
and U2837 (N_2837,N_2580,N_2610);
and U2838 (N_2838,N_2507,N_2717);
and U2839 (N_2839,N_2639,N_2535);
nor U2840 (N_2840,N_2696,N_2715);
and U2841 (N_2841,N_2629,N_2693);
nand U2842 (N_2842,N_2676,N_2734);
xnor U2843 (N_2843,N_2647,N_2520);
nand U2844 (N_2844,N_2509,N_2632);
nand U2845 (N_2845,N_2527,N_2576);
or U2846 (N_2846,N_2589,N_2597);
nor U2847 (N_2847,N_2574,N_2586);
or U2848 (N_2848,N_2578,N_2518);
or U2849 (N_2849,N_2685,N_2747);
nand U2850 (N_2850,N_2689,N_2588);
nand U2851 (N_2851,N_2532,N_2559);
nor U2852 (N_2852,N_2517,N_2657);
or U2853 (N_2853,N_2749,N_2669);
or U2854 (N_2854,N_2626,N_2661);
xnor U2855 (N_2855,N_2591,N_2618);
nand U2856 (N_2856,N_2668,N_2521);
nand U2857 (N_2857,N_2722,N_2514);
nor U2858 (N_2858,N_2602,N_2699);
nand U2859 (N_2859,N_2659,N_2503);
and U2860 (N_2860,N_2544,N_2543);
or U2861 (N_2861,N_2502,N_2570);
nor U2862 (N_2862,N_2681,N_2662);
or U2863 (N_2863,N_2565,N_2621);
and U2864 (N_2864,N_2616,N_2590);
or U2865 (N_2865,N_2623,N_2663);
and U2866 (N_2866,N_2598,N_2666);
or U2867 (N_2867,N_2614,N_2525);
or U2868 (N_2868,N_2523,N_2690);
xor U2869 (N_2869,N_2691,N_2643);
and U2870 (N_2870,N_2705,N_2530);
nand U2871 (N_2871,N_2533,N_2607);
and U2872 (N_2872,N_2719,N_2595);
and U2873 (N_2873,N_2658,N_2675);
and U2874 (N_2874,N_2519,N_2510);
xnor U2875 (N_2875,N_2663,N_2721);
and U2876 (N_2876,N_2668,N_2670);
nand U2877 (N_2877,N_2668,N_2618);
nor U2878 (N_2878,N_2718,N_2612);
or U2879 (N_2879,N_2557,N_2585);
or U2880 (N_2880,N_2711,N_2667);
nand U2881 (N_2881,N_2589,N_2586);
nand U2882 (N_2882,N_2683,N_2713);
nor U2883 (N_2883,N_2662,N_2650);
or U2884 (N_2884,N_2546,N_2649);
and U2885 (N_2885,N_2664,N_2657);
nand U2886 (N_2886,N_2657,N_2687);
or U2887 (N_2887,N_2606,N_2615);
nor U2888 (N_2888,N_2619,N_2535);
or U2889 (N_2889,N_2706,N_2744);
or U2890 (N_2890,N_2720,N_2669);
nor U2891 (N_2891,N_2591,N_2562);
and U2892 (N_2892,N_2606,N_2539);
or U2893 (N_2893,N_2521,N_2584);
nand U2894 (N_2894,N_2676,N_2662);
or U2895 (N_2895,N_2672,N_2643);
nor U2896 (N_2896,N_2628,N_2642);
or U2897 (N_2897,N_2669,N_2678);
xor U2898 (N_2898,N_2699,N_2668);
and U2899 (N_2899,N_2562,N_2731);
nand U2900 (N_2900,N_2604,N_2637);
or U2901 (N_2901,N_2532,N_2534);
nand U2902 (N_2902,N_2695,N_2585);
or U2903 (N_2903,N_2680,N_2584);
and U2904 (N_2904,N_2621,N_2683);
nand U2905 (N_2905,N_2683,N_2615);
and U2906 (N_2906,N_2749,N_2510);
or U2907 (N_2907,N_2624,N_2738);
or U2908 (N_2908,N_2527,N_2520);
nor U2909 (N_2909,N_2594,N_2524);
nor U2910 (N_2910,N_2683,N_2692);
nor U2911 (N_2911,N_2705,N_2743);
nor U2912 (N_2912,N_2618,N_2718);
nand U2913 (N_2913,N_2626,N_2641);
xnor U2914 (N_2914,N_2523,N_2656);
nand U2915 (N_2915,N_2566,N_2642);
nand U2916 (N_2916,N_2684,N_2687);
or U2917 (N_2917,N_2640,N_2559);
nor U2918 (N_2918,N_2739,N_2730);
and U2919 (N_2919,N_2733,N_2582);
and U2920 (N_2920,N_2747,N_2514);
or U2921 (N_2921,N_2714,N_2628);
nor U2922 (N_2922,N_2501,N_2644);
and U2923 (N_2923,N_2590,N_2726);
xnor U2924 (N_2924,N_2659,N_2551);
nand U2925 (N_2925,N_2588,N_2505);
nor U2926 (N_2926,N_2514,N_2594);
or U2927 (N_2927,N_2588,N_2710);
nand U2928 (N_2928,N_2738,N_2574);
nor U2929 (N_2929,N_2594,N_2504);
and U2930 (N_2930,N_2515,N_2688);
nand U2931 (N_2931,N_2532,N_2680);
and U2932 (N_2932,N_2662,N_2636);
xnor U2933 (N_2933,N_2666,N_2639);
and U2934 (N_2934,N_2609,N_2526);
nor U2935 (N_2935,N_2550,N_2622);
and U2936 (N_2936,N_2686,N_2539);
or U2937 (N_2937,N_2522,N_2725);
and U2938 (N_2938,N_2548,N_2744);
or U2939 (N_2939,N_2527,N_2566);
or U2940 (N_2940,N_2501,N_2654);
or U2941 (N_2941,N_2673,N_2737);
or U2942 (N_2942,N_2708,N_2506);
nand U2943 (N_2943,N_2548,N_2569);
nand U2944 (N_2944,N_2513,N_2709);
nor U2945 (N_2945,N_2531,N_2675);
and U2946 (N_2946,N_2712,N_2684);
xor U2947 (N_2947,N_2584,N_2546);
xnor U2948 (N_2948,N_2604,N_2656);
nand U2949 (N_2949,N_2640,N_2749);
nand U2950 (N_2950,N_2523,N_2555);
or U2951 (N_2951,N_2508,N_2613);
nor U2952 (N_2952,N_2651,N_2610);
or U2953 (N_2953,N_2546,N_2515);
and U2954 (N_2954,N_2574,N_2741);
or U2955 (N_2955,N_2659,N_2655);
nand U2956 (N_2956,N_2740,N_2647);
nand U2957 (N_2957,N_2586,N_2542);
nand U2958 (N_2958,N_2584,N_2514);
or U2959 (N_2959,N_2661,N_2594);
or U2960 (N_2960,N_2562,N_2531);
xnor U2961 (N_2961,N_2582,N_2638);
xnor U2962 (N_2962,N_2636,N_2743);
and U2963 (N_2963,N_2683,N_2654);
or U2964 (N_2964,N_2645,N_2734);
xnor U2965 (N_2965,N_2602,N_2748);
or U2966 (N_2966,N_2511,N_2589);
and U2967 (N_2967,N_2581,N_2685);
xnor U2968 (N_2968,N_2578,N_2607);
nor U2969 (N_2969,N_2709,N_2582);
and U2970 (N_2970,N_2569,N_2639);
xor U2971 (N_2971,N_2645,N_2665);
and U2972 (N_2972,N_2632,N_2550);
nand U2973 (N_2973,N_2569,N_2501);
and U2974 (N_2974,N_2563,N_2657);
nand U2975 (N_2975,N_2505,N_2648);
or U2976 (N_2976,N_2520,N_2597);
nor U2977 (N_2977,N_2708,N_2562);
xor U2978 (N_2978,N_2702,N_2652);
or U2979 (N_2979,N_2706,N_2598);
and U2980 (N_2980,N_2517,N_2586);
and U2981 (N_2981,N_2686,N_2664);
xnor U2982 (N_2982,N_2517,N_2681);
nor U2983 (N_2983,N_2745,N_2719);
or U2984 (N_2984,N_2619,N_2694);
nor U2985 (N_2985,N_2597,N_2649);
nand U2986 (N_2986,N_2660,N_2697);
nor U2987 (N_2987,N_2560,N_2631);
and U2988 (N_2988,N_2723,N_2747);
and U2989 (N_2989,N_2563,N_2527);
and U2990 (N_2990,N_2728,N_2620);
and U2991 (N_2991,N_2564,N_2616);
nand U2992 (N_2992,N_2523,N_2625);
nand U2993 (N_2993,N_2575,N_2663);
and U2994 (N_2994,N_2505,N_2605);
or U2995 (N_2995,N_2659,N_2746);
nor U2996 (N_2996,N_2716,N_2607);
nor U2997 (N_2997,N_2721,N_2594);
nor U2998 (N_2998,N_2648,N_2580);
or U2999 (N_2999,N_2570,N_2714);
or U3000 (N_3000,N_2907,N_2842);
and U3001 (N_3001,N_2799,N_2761);
and U3002 (N_3002,N_2817,N_2812);
nand U3003 (N_3003,N_2762,N_2835);
and U3004 (N_3004,N_2836,N_2877);
or U3005 (N_3005,N_2838,N_2750);
or U3006 (N_3006,N_2795,N_2926);
or U3007 (N_3007,N_2798,N_2934);
and U3008 (N_3008,N_2765,N_2963);
nand U3009 (N_3009,N_2902,N_2950);
and U3010 (N_3010,N_2942,N_2814);
nor U3011 (N_3011,N_2751,N_2851);
and U3012 (N_3012,N_2821,N_2763);
nand U3013 (N_3013,N_2833,N_2793);
nand U3014 (N_3014,N_2978,N_2925);
nand U3015 (N_3015,N_2891,N_2752);
nor U3016 (N_3016,N_2916,N_2875);
and U3017 (N_3017,N_2971,N_2989);
nor U3018 (N_3018,N_2809,N_2786);
nor U3019 (N_3019,N_2981,N_2767);
and U3020 (N_3020,N_2810,N_2895);
or U3021 (N_3021,N_2945,N_2860);
nor U3022 (N_3022,N_2951,N_2889);
or U3023 (N_3023,N_2936,N_2943);
nor U3024 (N_3024,N_2852,N_2892);
and U3025 (N_3025,N_2998,N_2960);
and U3026 (N_3026,N_2755,N_2830);
nor U3027 (N_3027,N_2959,N_2898);
nor U3028 (N_3028,N_2976,N_2893);
nand U3029 (N_3029,N_2756,N_2988);
nor U3030 (N_3030,N_2953,N_2828);
nor U3031 (N_3031,N_2856,N_2944);
nor U3032 (N_3032,N_2802,N_2791);
nand U3033 (N_3033,N_2825,N_2894);
nand U3034 (N_3034,N_2864,N_2826);
nand U3035 (N_3035,N_2858,N_2947);
nor U3036 (N_3036,N_2969,N_2939);
nor U3037 (N_3037,N_2783,N_2957);
or U3038 (N_3038,N_2941,N_2999);
or U3039 (N_3039,N_2949,N_2993);
xnor U3040 (N_3040,N_2946,N_2857);
nor U3041 (N_3041,N_2768,N_2918);
and U3042 (N_3042,N_2774,N_2766);
nor U3043 (N_3043,N_2840,N_2787);
or U3044 (N_3044,N_2868,N_2871);
and U3045 (N_3045,N_2986,N_2772);
nand U3046 (N_3046,N_2757,N_2880);
or U3047 (N_3047,N_2804,N_2940);
or U3048 (N_3048,N_2967,N_2775);
or U3049 (N_3049,N_2824,N_2844);
nor U3050 (N_3050,N_2987,N_2778);
xnor U3051 (N_3051,N_2754,N_2921);
and U3052 (N_3052,N_2792,N_2972);
nor U3053 (N_3053,N_2924,N_2827);
or U3054 (N_3054,N_2917,N_2848);
or U3055 (N_3055,N_2965,N_2784);
nor U3056 (N_3056,N_2872,N_2901);
nor U3057 (N_3057,N_2769,N_2862);
or U3058 (N_3058,N_2923,N_2829);
or U3059 (N_3059,N_2759,N_2956);
xor U3060 (N_3060,N_2878,N_2760);
or U3061 (N_3061,N_2776,N_2900);
and U3062 (N_3062,N_2758,N_2906);
nor U3063 (N_3063,N_2847,N_2797);
or U3064 (N_3064,N_2905,N_2948);
and U3065 (N_3065,N_2850,N_2980);
nor U3066 (N_3066,N_2876,N_2927);
or U3067 (N_3067,N_2996,N_2865);
and U3068 (N_3068,N_2977,N_2818);
or U3069 (N_3069,N_2785,N_2883);
nor U3070 (N_3070,N_2834,N_2803);
nor U3071 (N_3071,N_2968,N_2973);
and U3072 (N_3072,N_2777,N_2909);
and U3073 (N_3073,N_2870,N_2845);
nand U3074 (N_3074,N_2979,N_2753);
nor U3075 (N_3075,N_2952,N_2807);
nor U3076 (N_3076,N_2962,N_2914);
and U3077 (N_3077,N_2819,N_2932);
xnor U3078 (N_3078,N_2970,N_2904);
or U3079 (N_3079,N_2808,N_2888);
and U3080 (N_3080,N_2882,N_2899);
xor U3081 (N_3081,N_2854,N_2781);
or U3082 (N_3082,N_2975,N_2855);
or U3083 (N_3083,N_2874,N_2822);
nand U3084 (N_3084,N_2782,N_2832);
or U3085 (N_3085,N_2958,N_2839);
and U3086 (N_3086,N_2897,N_2796);
and U3087 (N_3087,N_2867,N_2984);
and U3088 (N_3088,N_2866,N_2890);
and U3089 (N_3089,N_2790,N_2933);
nor U3090 (N_3090,N_2990,N_2800);
nand U3091 (N_3091,N_2928,N_2823);
nor U3092 (N_3092,N_2873,N_2794);
and U3093 (N_3093,N_2982,N_2779);
or U3094 (N_3094,N_2966,N_2911);
nor U3095 (N_3095,N_2954,N_2997);
nand U3096 (N_3096,N_2831,N_2903);
nor U3097 (N_3097,N_2843,N_2811);
or U3098 (N_3098,N_2859,N_2884);
nand U3099 (N_3099,N_2770,N_2974);
and U3100 (N_3100,N_2773,N_2881);
nand U3101 (N_3101,N_2985,N_2994);
nand U3102 (N_3102,N_2983,N_2764);
and U3103 (N_3103,N_2915,N_2910);
or U3104 (N_3104,N_2771,N_2920);
or U3105 (N_3105,N_2919,N_2861);
nor U3106 (N_3106,N_2913,N_2937);
nor U3107 (N_3107,N_2841,N_2991);
or U3108 (N_3108,N_2801,N_2853);
nor U3109 (N_3109,N_2805,N_2849);
or U3110 (N_3110,N_2931,N_2846);
xnor U3111 (N_3111,N_2863,N_2869);
and U3112 (N_3112,N_2813,N_2815);
nand U3113 (N_3113,N_2938,N_2930);
or U3114 (N_3114,N_2820,N_2885);
and U3115 (N_3115,N_2789,N_2896);
and U3116 (N_3116,N_2788,N_2961);
or U3117 (N_3117,N_2886,N_2879);
nor U3118 (N_3118,N_2887,N_2935);
and U3119 (N_3119,N_2955,N_2995);
and U3120 (N_3120,N_2908,N_2816);
or U3121 (N_3121,N_2806,N_2964);
nor U3122 (N_3122,N_2992,N_2780);
nand U3123 (N_3123,N_2922,N_2837);
nand U3124 (N_3124,N_2929,N_2912);
and U3125 (N_3125,N_2865,N_2772);
and U3126 (N_3126,N_2870,N_2880);
xnor U3127 (N_3127,N_2787,N_2944);
nand U3128 (N_3128,N_2844,N_2837);
xnor U3129 (N_3129,N_2943,N_2975);
or U3130 (N_3130,N_2950,N_2896);
nand U3131 (N_3131,N_2847,N_2877);
or U3132 (N_3132,N_2844,N_2971);
or U3133 (N_3133,N_2866,N_2849);
nor U3134 (N_3134,N_2757,N_2828);
or U3135 (N_3135,N_2764,N_2889);
xor U3136 (N_3136,N_2844,N_2772);
nand U3137 (N_3137,N_2752,N_2957);
or U3138 (N_3138,N_2976,N_2793);
or U3139 (N_3139,N_2883,N_2984);
and U3140 (N_3140,N_2961,N_2818);
and U3141 (N_3141,N_2848,N_2936);
xor U3142 (N_3142,N_2915,N_2873);
nor U3143 (N_3143,N_2962,N_2904);
xor U3144 (N_3144,N_2924,N_2777);
nor U3145 (N_3145,N_2857,N_2925);
nor U3146 (N_3146,N_2889,N_2760);
xnor U3147 (N_3147,N_2825,N_2908);
nor U3148 (N_3148,N_2986,N_2782);
nand U3149 (N_3149,N_2864,N_2980);
or U3150 (N_3150,N_2800,N_2782);
and U3151 (N_3151,N_2930,N_2888);
nand U3152 (N_3152,N_2784,N_2783);
or U3153 (N_3153,N_2892,N_2809);
and U3154 (N_3154,N_2821,N_2919);
xor U3155 (N_3155,N_2809,N_2941);
and U3156 (N_3156,N_2885,N_2913);
nand U3157 (N_3157,N_2946,N_2952);
xnor U3158 (N_3158,N_2875,N_2753);
nand U3159 (N_3159,N_2844,N_2775);
and U3160 (N_3160,N_2780,N_2947);
nand U3161 (N_3161,N_2829,N_2781);
or U3162 (N_3162,N_2974,N_2778);
or U3163 (N_3163,N_2950,N_2925);
nand U3164 (N_3164,N_2830,N_2963);
xnor U3165 (N_3165,N_2944,N_2891);
and U3166 (N_3166,N_2969,N_2800);
or U3167 (N_3167,N_2975,N_2877);
xor U3168 (N_3168,N_2955,N_2779);
or U3169 (N_3169,N_2955,N_2980);
nor U3170 (N_3170,N_2752,N_2851);
or U3171 (N_3171,N_2959,N_2951);
or U3172 (N_3172,N_2781,N_2985);
nor U3173 (N_3173,N_2826,N_2821);
nor U3174 (N_3174,N_2855,N_2854);
nand U3175 (N_3175,N_2758,N_2766);
nor U3176 (N_3176,N_2812,N_2949);
nor U3177 (N_3177,N_2973,N_2841);
or U3178 (N_3178,N_2799,N_2927);
or U3179 (N_3179,N_2782,N_2992);
or U3180 (N_3180,N_2858,N_2953);
nor U3181 (N_3181,N_2983,N_2989);
nand U3182 (N_3182,N_2990,N_2919);
nand U3183 (N_3183,N_2816,N_2864);
or U3184 (N_3184,N_2771,N_2848);
and U3185 (N_3185,N_2896,N_2790);
and U3186 (N_3186,N_2959,N_2762);
and U3187 (N_3187,N_2803,N_2817);
and U3188 (N_3188,N_2809,N_2838);
xnor U3189 (N_3189,N_2768,N_2975);
nor U3190 (N_3190,N_2909,N_2852);
and U3191 (N_3191,N_2805,N_2884);
nand U3192 (N_3192,N_2999,N_2981);
and U3193 (N_3193,N_2980,N_2802);
nand U3194 (N_3194,N_2954,N_2774);
nor U3195 (N_3195,N_2921,N_2906);
nand U3196 (N_3196,N_2914,N_2906);
nor U3197 (N_3197,N_2878,N_2999);
or U3198 (N_3198,N_2882,N_2830);
and U3199 (N_3199,N_2987,N_2864);
or U3200 (N_3200,N_2793,N_2790);
or U3201 (N_3201,N_2855,N_2993);
nor U3202 (N_3202,N_2806,N_2822);
or U3203 (N_3203,N_2966,N_2804);
or U3204 (N_3204,N_2857,N_2801);
or U3205 (N_3205,N_2751,N_2752);
or U3206 (N_3206,N_2996,N_2754);
nor U3207 (N_3207,N_2826,N_2882);
nor U3208 (N_3208,N_2918,N_2861);
nor U3209 (N_3209,N_2950,N_2777);
nand U3210 (N_3210,N_2785,N_2866);
or U3211 (N_3211,N_2797,N_2822);
and U3212 (N_3212,N_2947,N_2812);
nand U3213 (N_3213,N_2821,N_2881);
nor U3214 (N_3214,N_2751,N_2806);
nand U3215 (N_3215,N_2995,N_2765);
and U3216 (N_3216,N_2787,N_2763);
nand U3217 (N_3217,N_2986,N_2834);
and U3218 (N_3218,N_2919,N_2755);
xnor U3219 (N_3219,N_2871,N_2834);
or U3220 (N_3220,N_2920,N_2950);
nor U3221 (N_3221,N_2856,N_2966);
nor U3222 (N_3222,N_2782,N_2847);
nor U3223 (N_3223,N_2781,N_2807);
nor U3224 (N_3224,N_2870,N_2884);
nand U3225 (N_3225,N_2921,N_2969);
xor U3226 (N_3226,N_2952,N_2902);
nor U3227 (N_3227,N_2779,N_2788);
nor U3228 (N_3228,N_2904,N_2873);
nor U3229 (N_3229,N_2930,N_2908);
nor U3230 (N_3230,N_2795,N_2996);
nand U3231 (N_3231,N_2797,N_2917);
xor U3232 (N_3232,N_2776,N_2935);
nand U3233 (N_3233,N_2784,N_2892);
nor U3234 (N_3234,N_2813,N_2885);
nor U3235 (N_3235,N_2804,N_2820);
and U3236 (N_3236,N_2786,N_2820);
and U3237 (N_3237,N_2787,N_2845);
xnor U3238 (N_3238,N_2957,N_2775);
nand U3239 (N_3239,N_2763,N_2996);
or U3240 (N_3240,N_2765,N_2932);
or U3241 (N_3241,N_2772,N_2794);
and U3242 (N_3242,N_2771,N_2804);
xnor U3243 (N_3243,N_2758,N_2759);
and U3244 (N_3244,N_2939,N_2793);
nor U3245 (N_3245,N_2829,N_2824);
or U3246 (N_3246,N_2857,N_2915);
and U3247 (N_3247,N_2905,N_2965);
nor U3248 (N_3248,N_2828,N_2880);
nand U3249 (N_3249,N_2851,N_2855);
nand U3250 (N_3250,N_3196,N_3082);
nor U3251 (N_3251,N_3128,N_3167);
and U3252 (N_3252,N_3040,N_3103);
xor U3253 (N_3253,N_3051,N_3073);
nor U3254 (N_3254,N_3116,N_3079);
or U3255 (N_3255,N_3009,N_3044);
nand U3256 (N_3256,N_3070,N_3094);
nor U3257 (N_3257,N_3003,N_3118);
nand U3258 (N_3258,N_3187,N_3151);
and U3259 (N_3259,N_3112,N_3234);
nor U3260 (N_3260,N_3205,N_3138);
and U3261 (N_3261,N_3123,N_3063);
nor U3262 (N_3262,N_3159,N_3023);
and U3263 (N_3263,N_3002,N_3247);
or U3264 (N_3264,N_3188,N_3028);
or U3265 (N_3265,N_3110,N_3072);
or U3266 (N_3266,N_3207,N_3027);
or U3267 (N_3267,N_3194,N_3013);
or U3268 (N_3268,N_3184,N_3032);
xor U3269 (N_3269,N_3107,N_3133);
or U3270 (N_3270,N_3046,N_3201);
and U3271 (N_3271,N_3136,N_3043);
and U3272 (N_3272,N_3031,N_3066);
xnor U3273 (N_3273,N_3149,N_3111);
nor U3274 (N_3274,N_3239,N_3039);
and U3275 (N_3275,N_3007,N_3172);
or U3276 (N_3276,N_3024,N_3176);
or U3277 (N_3277,N_3047,N_3122);
or U3278 (N_3278,N_3181,N_3085);
nand U3279 (N_3279,N_3091,N_3143);
nor U3280 (N_3280,N_3134,N_3035);
nand U3281 (N_3281,N_3147,N_3223);
xnor U3282 (N_3282,N_3217,N_3087);
and U3283 (N_3283,N_3202,N_3193);
or U3284 (N_3284,N_3076,N_3016);
nand U3285 (N_3285,N_3120,N_3050);
nor U3286 (N_3286,N_3019,N_3090);
nor U3287 (N_3287,N_3242,N_3204);
nor U3288 (N_3288,N_3077,N_3121);
xnor U3289 (N_3289,N_3001,N_3211);
xnor U3290 (N_3290,N_3071,N_3177);
nand U3291 (N_3291,N_3059,N_3097);
xnor U3292 (N_3292,N_3052,N_3240);
and U3293 (N_3293,N_3164,N_3086);
or U3294 (N_3294,N_3198,N_3233);
and U3295 (N_3295,N_3174,N_3175);
nor U3296 (N_3296,N_3119,N_3064);
nor U3297 (N_3297,N_3171,N_3238);
or U3298 (N_3298,N_3225,N_3126);
nand U3299 (N_3299,N_3130,N_3236);
and U3300 (N_3300,N_3034,N_3022);
xnor U3301 (N_3301,N_3135,N_3065);
or U3302 (N_3302,N_3095,N_3124);
nor U3303 (N_3303,N_3101,N_3197);
nand U3304 (N_3304,N_3131,N_3179);
or U3305 (N_3305,N_3089,N_3155);
nand U3306 (N_3306,N_3221,N_3140);
or U3307 (N_3307,N_3006,N_3154);
xnor U3308 (N_3308,N_3041,N_3098);
nand U3309 (N_3309,N_3132,N_3144);
or U3310 (N_3310,N_3212,N_3092);
nand U3311 (N_3311,N_3075,N_3061);
and U3312 (N_3312,N_3102,N_3104);
or U3313 (N_3313,N_3057,N_3195);
xnor U3314 (N_3314,N_3020,N_3005);
and U3315 (N_3315,N_3190,N_3241);
nor U3316 (N_3316,N_3108,N_3117);
nand U3317 (N_3317,N_3105,N_3088);
and U3318 (N_3318,N_3146,N_3083);
and U3319 (N_3319,N_3017,N_3045);
and U3320 (N_3320,N_3100,N_3080);
and U3321 (N_3321,N_3030,N_3200);
nand U3322 (N_3322,N_3231,N_3000);
nand U3323 (N_3323,N_3150,N_3008);
nand U3324 (N_3324,N_3173,N_3226);
nand U3325 (N_3325,N_3142,N_3222);
nor U3326 (N_3326,N_3067,N_3074);
xnor U3327 (N_3327,N_3156,N_3049);
and U3328 (N_3328,N_3014,N_3230);
and U3329 (N_3329,N_3199,N_3168);
or U3330 (N_3330,N_3021,N_3180);
nor U3331 (N_3331,N_3216,N_3191);
and U3332 (N_3332,N_3113,N_3068);
nor U3333 (N_3333,N_3186,N_3206);
and U3334 (N_3334,N_3153,N_3178);
or U3335 (N_3335,N_3227,N_3185);
nand U3336 (N_3336,N_3157,N_3096);
nor U3337 (N_3337,N_3249,N_3048);
and U3338 (N_3338,N_3192,N_3213);
nand U3339 (N_3339,N_3158,N_3145);
and U3340 (N_3340,N_3078,N_3125);
or U3341 (N_3341,N_3203,N_3210);
or U3342 (N_3342,N_3010,N_3127);
and U3343 (N_3343,N_3243,N_3169);
or U3344 (N_3344,N_3115,N_3232);
nand U3345 (N_3345,N_3218,N_3037);
nor U3346 (N_3346,N_3038,N_3081);
nand U3347 (N_3347,N_3161,N_3129);
nor U3348 (N_3348,N_3170,N_3183);
and U3349 (N_3349,N_3114,N_3141);
and U3350 (N_3350,N_3053,N_3036);
or U3351 (N_3351,N_3189,N_3162);
nand U3352 (N_3352,N_3084,N_3015);
nand U3353 (N_3353,N_3228,N_3099);
and U3354 (N_3354,N_3033,N_3182);
and U3355 (N_3355,N_3209,N_3069);
nand U3356 (N_3356,N_3152,N_3166);
and U3357 (N_3357,N_3093,N_3244);
or U3358 (N_3358,N_3163,N_3248);
nor U3359 (N_3359,N_3026,N_3025);
nor U3360 (N_3360,N_3056,N_3060);
nor U3361 (N_3361,N_3139,N_3246);
and U3362 (N_3362,N_3148,N_3237);
or U3363 (N_3363,N_3029,N_3109);
or U3364 (N_3364,N_3245,N_3229);
nand U3365 (N_3365,N_3160,N_3054);
or U3366 (N_3366,N_3011,N_3062);
nor U3367 (N_3367,N_3165,N_3220);
nand U3368 (N_3368,N_3012,N_3224);
or U3369 (N_3369,N_3055,N_3058);
or U3370 (N_3370,N_3214,N_3004);
or U3371 (N_3371,N_3042,N_3235);
xnor U3372 (N_3372,N_3018,N_3137);
nor U3373 (N_3373,N_3106,N_3219);
or U3374 (N_3374,N_3208,N_3215);
and U3375 (N_3375,N_3172,N_3113);
or U3376 (N_3376,N_3240,N_3021);
nor U3377 (N_3377,N_3017,N_3152);
and U3378 (N_3378,N_3091,N_3183);
nand U3379 (N_3379,N_3189,N_3053);
nor U3380 (N_3380,N_3083,N_3053);
nand U3381 (N_3381,N_3170,N_3038);
or U3382 (N_3382,N_3061,N_3051);
nand U3383 (N_3383,N_3089,N_3022);
and U3384 (N_3384,N_3148,N_3100);
and U3385 (N_3385,N_3249,N_3147);
nand U3386 (N_3386,N_3017,N_3166);
nand U3387 (N_3387,N_3052,N_3209);
or U3388 (N_3388,N_3135,N_3002);
nand U3389 (N_3389,N_3064,N_3161);
nand U3390 (N_3390,N_3155,N_3043);
or U3391 (N_3391,N_3171,N_3210);
or U3392 (N_3392,N_3146,N_3150);
and U3393 (N_3393,N_3017,N_3099);
nor U3394 (N_3394,N_3082,N_3134);
or U3395 (N_3395,N_3120,N_3069);
xor U3396 (N_3396,N_3190,N_3166);
nand U3397 (N_3397,N_3029,N_3097);
xnor U3398 (N_3398,N_3075,N_3156);
and U3399 (N_3399,N_3234,N_3074);
and U3400 (N_3400,N_3083,N_3038);
and U3401 (N_3401,N_3213,N_3052);
or U3402 (N_3402,N_3223,N_3114);
nor U3403 (N_3403,N_3094,N_3129);
and U3404 (N_3404,N_3156,N_3158);
nand U3405 (N_3405,N_3106,N_3246);
xor U3406 (N_3406,N_3083,N_3047);
and U3407 (N_3407,N_3228,N_3165);
or U3408 (N_3408,N_3096,N_3091);
and U3409 (N_3409,N_3194,N_3165);
and U3410 (N_3410,N_3043,N_3148);
or U3411 (N_3411,N_3050,N_3021);
or U3412 (N_3412,N_3106,N_3068);
nand U3413 (N_3413,N_3037,N_3131);
nand U3414 (N_3414,N_3147,N_3207);
nand U3415 (N_3415,N_3173,N_3054);
or U3416 (N_3416,N_3114,N_3181);
or U3417 (N_3417,N_3227,N_3099);
nor U3418 (N_3418,N_3154,N_3239);
or U3419 (N_3419,N_3093,N_3018);
nand U3420 (N_3420,N_3169,N_3233);
nor U3421 (N_3421,N_3213,N_3218);
nand U3422 (N_3422,N_3020,N_3004);
and U3423 (N_3423,N_3089,N_3110);
or U3424 (N_3424,N_3048,N_3222);
nand U3425 (N_3425,N_3238,N_3166);
or U3426 (N_3426,N_3141,N_3061);
nand U3427 (N_3427,N_3060,N_3064);
nor U3428 (N_3428,N_3161,N_3006);
and U3429 (N_3429,N_3151,N_3056);
nor U3430 (N_3430,N_3107,N_3222);
or U3431 (N_3431,N_3218,N_3120);
nand U3432 (N_3432,N_3209,N_3248);
or U3433 (N_3433,N_3190,N_3033);
nand U3434 (N_3434,N_3161,N_3134);
and U3435 (N_3435,N_3119,N_3175);
xnor U3436 (N_3436,N_3015,N_3138);
and U3437 (N_3437,N_3173,N_3113);
and U3438 (N_3438,N_3235,N_3241);
and U3439 (N_3439,N_3067,N_3190);
nand U3440 (N_3440,N_3106,N_3086);
nor U3441 (N_3441,N_3071,N_3060);
nand U3442 (N_3442,N_3123,N_3150);
nand U3443 (N_3443,N_3214,N_3003);
or U3444 (N_3444,N_3194,N_3163);
nor U3445 (N_3445,N_3154,N_3238);
nor U3446 (N_3446,N_3228,N_3169);
or U3447 (N_3447,N_3008,N_3045);
and U3448 (N_3448,N_3198,N_3224);
and U3449 (N_3449,N_3117,N_3012);
nor U3450 (N_3450,N_3100,N_3059);
xnor U3451 (N_3451,N_3243,N_3134);
or U3452 (N_3452,N_3100,N_3136);
and U3453 (N_3453,N_3135,N_3101);
nor U3454 (N_3454,N_3161,N_3130);
or U3455 (N_3455,N_3200,N_3024);
nor U3456 (N_3456,N_3029,N_3103);
xor U3457 (N_3457,N_3075,N_3094);
nand U3458 (N_3458,N_3195,N_3233);
nor U3459 (N_3459,N_3220,N_3111);
and U3460 (N_3460,N_3001,N_3186);
xor U3461 (N_3461,N_3066,N_3131);
nand U3462 (N_3462,N_3014,N_3202);
and U3463 (N_3463,N_3113,N_3074);
nor U3464 (N_3464,N_3007,N_3058);
xnor U3465 (N_3465,N_3038,N_3166);
nor U3466 (N_3466,N_3186,N_3204);
xnor U3467 (N_3467,N_3113,N_3243);
or U3468 (N_3468,N_3174,N_3151);
or U3469 (N_3469,N_3190,N_3015);
nand U3470 (N_3470,N_3142,N_3140);
and U3471 (N_3471,N_3027,N_3010);
xnor U3472 (N_3472,N_3125,N_3074);
and U3473 (N_3473,N_3169,N_3056);
nor U3474 (N_3474,N_3172,N_3028);
xnor U3475 (N_3475,N_3026,N_3190);
nand U3476 (N_3476,N_3195,N_3019);
and U3477 (N_3477,N_3148,N_3202);
nand U3478 (N_3478,N_3122,N_3080);
or U3479 (N_3479,N_3160,N_3220);
nand U3480 (N_3480,N_3166,N_3016);
and U3481 (N_3481,N_3014,N_3168);
and U3482 (N_3482,N_3168,N_3056);
xnor U3483 (N_3483,N_3142,N_3113);
nand U3484 (N_3484,N_3000,N_3137);
nor U3485 (N_3485,N_3171,N_3152);
nor U3486 (N_3486,N_3027,N_3093);
nor U3487 (N_3487,N_3105,N_3054);
and U3488 (N_3488,N_3199,N_3138);
and U3489 (N_3489,N_3145,N_3011);
xor U3490 (N_3490,N_3019,N_3184);
xnor U3491 (N_3491,N_3125,N_3178);
or U3492 (N_3492,N_3118,N_3210);
nand U3493 (N_3493,N_3248,N_3162);
and U3494 (N_3494,N_3163,N_3063);
nand U3495 (N_3495,N_3108,N_3238);
or U3496 (N_3496,N_3072,N_3100);
nand U3497 (N_3497,N_3075,N_3155);
or U3498 (N_3498,N_3065,N_3076);
nor U3499 (N_3499,N_3073,N_3069);
nand U3500 (N_3500,N_3282,N_3406);
or U3501 (N_3501,N_3359,N_3486);
nand U3502 (N_3502,N_3450,N_3410);
or U3503 (N_3503,N_3252,N_3395);
and U3504 (N_3504,N_3447,N_3440);
xor U3505 (N_3505,N_3496,N_3421);
and U3506 (N_3506,N_3307,N_3444);
xor U3507 (N_3507,N_3376,N_3328);
xor U3508 (N_3508,N_3475,N_3477);
or U3509 (N_3509,N_3377,N_3433);
nor U3510 (N_3510,N_3474,N_3429);
nor U3511 (N_3511,N_3363,N_3420);
and U3512 (N_3512,N_3455,N_3375);
nand U3513 (N_3513,N_3344,N_3296);
or U3514 (N_3514,N_3281,N_3451);
or U3515 (N_3515,N_3471,N_3497);
xnor U3516 (N_3516,N_3371,N_3273);
or U3517 (N_3517,N_3330,N_3286);
and U3518 (N_3518,N_3367,N_3487);
xor U3519 (N_3519,N_3460,N_3457);
and U3520 (N_3520,N_3260,N_3306);
and U3521 (N_3521,N_3384,N_3289);
or U3522 (N_3522,N_3357,N_3480);
or U3523 (N_3523,N_3326,N_3324);
or U3524 (N_3524,N_3295,N_3255);
or U3525 (N_3525,N_3332,N_3453);
and U3526 (N_3526,N_3396,N_3464);
xor U3527 (N_3527,N_3272,N_3360);
and U3528 (N_3528,N_3492,N_3391);
and U3529 (N_3529,N_3370,N_3342);
nand U3530 (N_3530,N_3257,N_3473);
nand U3531 (N_3531,N_3358,N_3254);
nand U3532 (N_3532,N_3308,N_3408);
nand U3533 (N_3533,N_3339,N_3442);
or U3534 (N_3534,N_3274,N_3347);
or U3535 (N_3535,N_3491,N_3291);
nor U3536 (N_3536,N_3399,N_3428);
or U3537 (N_3537,N_3418,N_3351);
nor U3538 (N_3538,N_3362,N_3387);
and U3539 (N_3539,N_3490,N_3298);
nand U3540 (N_3540,N_3317,N_3338);
and U3541 (N_3541,N_3299,N_3319);
and U3542 (N_3542,N_3304,N_3393);
and U3543 (N_3543,N_3456,N_3264);
or U3544 (N_3544,N_3305,N_3270);
nand U3545 (N_3545,N_3413,N_3314);
or U3546 (N_3546,N_3427,N_3432);
nand U3547 (N_3547,N_3335,N_3383);
nand U3548 (N_3548,N_3280,N_3364);
nor U3549 (N_3549,N_3345,N_3300);
and U3550 (N_3550,N_3278,N_3417);
and U3551 (N_3551,N_3355,N_3388);
or U3552 (N_3552,N_3368,N_3262);
nor U3553 (N_3553,N_3318,N_3253);
and U3554 (N_3554,N_3416,N_3284);
or U3555 (N_3555,N_3365,N_3354);
and U3556 (N_3556,N_3398,N_3379);
nor U3557 (N_3557,N_3467,N_3385);
and U3558 (N_3558,N_3381,N_3414);
nor U3559 (N_3559,N_3378,N_3343);
xnor U3560 (N_3560,N_3250,N_3315);
xor U3561 (N_3561,N_3405,N_3403);
nor U3562 (N_3562,N_3266,N_3293);
and U3563 (N_3563,N_3484,N_3415);
nand U3564 (N_3564,N_3348,N_3337);
nand U3565 (N_3565,N_3320,N_3312);
or U3566 (N_3566,N_3470,N_3472);
nand U3567 (N_3567,N_3369,N_3481);
nor U3568 (N_3568,N_3466,N_3443);
xor U3569 (N_3569,N_3448,N_3404);
nand U3570 (N_3570,N_3439,N_3271);
xnor U3571 (N_3571,N_3275,N_3498);
or U3572 (N_3572,N_3259,N_3340);
and U3573 (N_3573,N_3325,N_3435);
and U3574 (N_3574,N_3465,N_3302);
or U3575 (N_3575,N_3283,N_3454);
nor U3576 (N_3576,N_3438,N_3494);
and U3577 (N_3577,N_3287,N_3469);
nor U3578 (N_3578,N_3279,N_3452);
or U3579 (N_3579,N_3483,N_3353);
or U3580 (N_3580,N_3411,N_3301);
or U3581 (N_3581,N_3321,N_3482);
xor U3582 (N_3582,N_3309,N_3402);
and U3583 (N_3583,N_3495,N_3366);
and U3584 (N_3584,N_3419,N_3445);
and U3585 (N_3585,N_3441,N_3478);
and U3586 (N_3586,N_3251,N_3311);
and U3587 (N_3587,N_3316,N_3380);
xor U3588 (N_3588,N_3336,N_3374);
or U3589 (N_3589,N_3462,N_3261);
nand U3590 (N_3590,N_3485,N_3263);
nand U3591 (N_3591,N_3493,N_3422);
and U3592 (N_3592,N_3392,N_3488);
nor U3593 (N_3593,N_3436,N_3268);
and U3594 (N_3594,N_3256,N_3499);
or U3595 (N_3595,N_3382,N_3310);
nor U3596 (N_3596,N_3400,N_3258);
and U3597 (N_3597,N_3269,N_3285);
nor U3598 (N_3598,N_3333,N_3350);
and U3599 (N_3599,N_3276,N_3458);
nor U3600 (N_3600,N_3334,N_3361);
and U3601 (N_3601,N_3329,N_3409);
xor U3602 (N_3602,N_3277,N_3322);
nand U3603 (N_3603,N_3390,N_3401);
nor U3604 (N_3604,N_3424,N_3294);
or U3605 (N_3605,N_3412,N_3394);
or U3606 (N_3606,N_3431,N_3423);
or U3607 (N_3607,N_3463,N_3459);
nand U3608 (N_3608,N_3476,N_3303);
nor U3609 (N_3609,N_3346,N_3372);
xnor U3610 (N_3610,N_3468,N_3449);
nand U3611 (N_3611,N_3267,N_3425);
or U3612 (N_3612,N_3434,N_3430);
nor U3613 (N_3613,N_3352,N_3437);
nor U3614 (N_3614,N_3331,N_3489);
nand U3615 (N_3615,N_3292,N_3479);
nand U3616 (N_3616,N_3341,N_3389);
and U3617 (N_3617,N_3356,N_3386);
and U3618 (N_3618,N_3446,N_3327);
and U3619 (N_3619,N_3373,N_3288);
and U3620 (N_3620,N_3290,N_3461);
or U3621 (N_3621,N_3323,N_3313);
or U3622 (N_3622,N_3349,N_3407);
or U3623 (N_3623,N_3265,N_3426);
and U3624 (N_3624,N_3397,N_3297);
nor U3625 (N_3625,N_3373,N_3265);
and U3626 (N_3626,N_3274,N_3442);
and U3627 (N_3627,N_3250,N_3396);
or U3628 (N_3628,N_3416,N_3275);
nand U3629 (N_3629,N_3465,N_3350);
or U3630 (N_3630,N_3308,N_3403);
nor U3631 (N_3631,N_3368,N_3365);
nor U3632 (N_3632,N_3488,N_3436);
nor U3633 (N_3633,N_3389,N_3266);
or U3634 (N_3634,N_3497,N_3339);
or U3635 (N_3635,N_3482,N_3265);
nand U3636 (N_3636,N_3300,N_3324);
nand U3637 (N_3637,N_3440,N_3341);
nor U3638 (N_3638,N_3294,N_3498);
nand U3639 (N_3639,N_3393,N_3295);
nand U3640 (N_3640,N_3320,N_3362);
nand U3641 (N_3641,N_3267,N_3389);
or U3642 (N_3642,N_3352,N_3441);
nor U3643 (N_3643,N_3346,N_3265);
and U3644 (N_3644,N_3270,N_3291);
and U3645 (N_3645,N_3316,N_3399);
or U3646 (N_3646,N_3486,N_3441);
nand U3647 (N_3647,N_3425,N_3466);
or U3648 (N_3648,N_3419,N_3416);
xor U3649 (N_3649,N_3270,N_3256);
or U3650 (N_3650,N_3350,N_3413);
nor U3651 (N_3651,N_3430,N_3310);
nor U3652 (N_3652,N_3471,N_3296);
or U3653 (N_3653,N_3267,N_3310);
nor U3654 (N_3654,N_3441,N_3434);
or U3655 (N_3655,N_3479,N_3439);
and U3656 (N_3656,N_3401,N_3334);
or U3657 (N_3657,N_3484,N_3433);
or U3658 (N_3658,N_3432,N_3395);
or U3659 (N_3659,N_3429,N_3293);
or U3660 (N_3660,N_3482,N_3286);
and U3661 (N_3661,N_3499,N_3488);
or U3662 (N_3662,N_3316,N_3308);
nor U3663 (N_3663,N_3322,N_3391);
nand U3664 (N_3664,N_3346,N_3411);
nor U3665 (N_3665,N_3409,N_3420);
nor U3666 (N_3666,N_3250,N_3324);
nand U3667 (N_3667,N_3391,N_3355);
nor U3668 (N_3668,N_3396,N_3335);
nor U3669 (N_3669,N_3479,N_3445);
nor U3670 (N_3670,N_3284,N_3378);
or U3671 (N_3671,N_3290,N_3251);
or U3672 (N_3672,N_3462,N_3352);
nand U3673 (N_3673,N_3393,N_3283);
or U3674 (N_3674,N_3446,N_3274);
nor U3675 (N_3675,N_3315,N_3311);
and U3676 (N_3676,N_3460,N_3250);
nand U3677 (N_3677,N_3498,N_3386);
or U3678 (N_3678,N_3385,N_3402);
nor U3679 (N_3679,N_3423,N_3331);
nand U3680 (N_3680,N_3454,N_3461);
or U3681 (N_3681,N_3353,N_3438);
or U3682 (N_3682,N_3370,N_3254);
nand U3683 (N_3683,N_3322,N_3308);
xnor U3684 (N_3684,N_3318,N_3339);
nand U3685 (N_3685,N_3466,N_3474);
and U3686 (N_3686,N_3250,N_3498);
and U3687 (N_3687,N_3289,N_3342);
or U3688 (N_3688,N_3375,N_3436);
or U3689 (N_3689,N_3394,N_3283);
and U3690 (N_3690,N_3446,N_3456);
xor U3691 (N_3691,N_3439,N_3451);
or U3692 (N_3692,N_3337,N_3373);
nand U3693 (N_3693,N_3471,N_3410);
nor U3694 (N_3694,N_3369,N_3396);
nor U3695 (N_3695,N_3299,N_3463);
or U3696 (N_3696,N_3372,N_3386);
and U3697 (N_3697,N_3330,N_3408);
nand U3698 (N_3698,N_3430,N_3375);
and U3699 (N_3699,N_3406,N_3258);
or U3700 (N_3700,N_3436,N_3461);
nand U3701 (N_3701,N_3270,N_3325);
nor U3702 (N_3702,N_3467,N_3328);
nand U3703 (N_3703,N_3256,N_3498);
nor U3704 (N_3704,N_3272,N_3442);
nand U3705 (N_3705,N_3461,N_3434);
and U3706 (N_3706,N_3448,N_3258);
or U3707 (N_3707,N_3296,N_3348);
and U3708 (N_3708,N_3453,N_3365);
or U3709 (N_3709,N_3267,N_3446);
nor U3710 (N_3710,N_3348,N_3432);
and U3711 (N_3711,N_3409,N_3419);
nand U3712 (N_3712,N_3351,N_3471);
or U3713 (N_3713,N_3322,N_3281);
or U3714 (N_3714,N_3422,N_3463);
nand U3715 (N_3715,N_3401,N_3406);
or U3716 (N_3716,N_3398,N_3441);
nor U3717 (N_3717,N_3421,N_3475);
nand U3718 (N_3718,N_3407,N_3304);
or U3719 (N_3719,N_3476,N_3425);
and U3720 (N_3720,N_3309,N_3373);
nand U3721 (N_3721,N_3358,N_3480);
nand U3722 (N_3722,N_3428,N_3353);
and U3723 (N_3723,N_3385,N_3373);
and U3724 (N_3724,N_3296,N_3334);
xnor U3725 (N_3725,N_3297,N_3385);
and U3726 (N_3726,N_3484,N_3428);
xor U3727 (N_3727,N_3383,N_3474);
nor U3728 (N_3728,N_3421,N_3372);
and U3729 (N_3729,N_3457,N_3273);
nor U3730 (N_3730,N_3273,N_3414);
xnor U3731 (N_3731,N_3402,N_3488);
nand U3732 (N_3732,N_3329,N_3288);
xor U3733 (N_3733,N_3323,N_3285);
or U3734 (N_3734,N_3490,N_3372);
or U3735 (N_3735,N_3490,N_3485);
or U3736 (N_3736,N_3315,N_3296);
nor U3737 (N_3737,N_3430,N_3338);
nor U3738 (N_3738,N_3403,N_3322);
and U3739 (N_3739,N_3353,N_3392);
nor U3740 (N_3740,N_3408,N_3283);
or U3741 (N_3741,N_3268,N_3441);
and U3742 (N_3742,N_3462,N_3444);
or U3743 (N_3743,N_3442,N_3285);
nand U3744 (N_3744,N_3267,N_3296);
nand U3745 (N_3745,N_3277,N_3305);
and U3746 (N_3746,N_3299,N_3284);
nor U3747 (N_3747,N_3460,N_3334);
or U3748 (N_3748,N_3328,N_3348);
and U3749 (N_3749,N_3443,N_3337);
nor U3750 (N_3750,N_3526,N_3748);
and U3751 (N_3751,N_3565,N_3722);
and U3752 (N_3752,N_3564,N_3556);
nand U3753 (N_3753,N_3504,N_3613);
or U3754 (N_3754,N_3629,N_3721);
nand U3755 (N_3755,N_3543,N_3637);
nor U3756 (N_3756,N_3732,N_3743);
or U3757 (N_3757,N_3635,N_3723);
nand U3758 (N_3758,N_3636,N_3671);
nand U3759 (N_3759,N_3575,N_3674);
or U3760 (N_3760,N_3606,N_3547);
nand U3761 (N_3761,N_3655,N_3570);
or U3762 (N_3762,N_3622,N_3514);
and U3763 (N_3763,N_3625,N_3580);
nand U3764 (N_3764,N_3612,N_3610);
nor U3765 (N_3765,N_3587,N_3739);
nor U3766 (N_3766,N_3714,N_3686);
nor U3767 (N_3767,N_3687,N_3599);
nor U3768 (N_3768,N_3713,N_3663);
nor U3769 (N_3769,N_3561,N_3503);
or U3770 (N_3770,N_3501,N_3520);
xor U3771 (N_3771,N_3654,N_3708);
and U3772 (N_3772,N_3670,N_3640);
nor U3773 (N_3773,N_3676,N_3525);
or U3774 (N_3774,N_3720,N_3736);
xnor U3775 (N_3775,N_3604,N_3729);
and U3776 (N_3776,N_3649,N_3740);
nand U3777 (N_3777,N_3683,N_3523);
nand U3778 (N_3778,N_3596,N_3505);
nand U3779 (N_3779,N_3704,N_3672);
nor U3780 (N_3780,N_3725,N_3518);
or U3781 (N_3781,N_3567,N_3553);
nor U3782 (N_3782,N_3638,N_3726);
nand U3783 (N_3783,N_3691,N_3656);
nand U3784 (N_3784,N_3516,N_3517);
nor U3785 (N_3785,N_3552,N_3696);
nor U3786 (N_3786,N_3593,N_3569);
nand U3787 (N_3787,N_3572,N_3560);
or U3788 (N_3788,N_3662,N_3749);
or U3789 (N_3789,N_3633,N_3549);
nor U3790 (N_3790,N_3632,N_3614);
nor U3791 (N_3791,N_3621,N_3643);
or U3792 (N_3792,N_3602,N_3694);
nor U3793 (N_3793,N_3534,N_3512);
xnor U3794 (N_3794,N_3611,N_3646);
or U3795 (N_3795,N_3650,N_3581);
or U3796 (N_3796,N_3521,N_3700);
or U3797 (N_3797,N_3678,N_3727);
nor U3798 (N_3798,N_3506,N_3571);
nand U3799 (N_3799,N_3542,N_3529);
and U3800 (N_3800,N_3680,N_3698);
or U3801 (N_3801,N_3738,N_3710);
nand U3802 (N_3802,N_3617,N_3665);
nor U3803 (N_3803,N_3668,N_3681);
nor U3804 (N_3804,N_3550,N_3509);
or U3805 (N_3805,N_3563,N_3623);
or U3806 (N_3806,N_3579,N_3568);
xnor U3807 (N_3807,N_3536,N_3711);
nor U3808 (N_3808,N_3511,N_3741);
nand U3809 (N_3809,N_3519,N_3634);
nand U3810 (N_3810,N_3719,N_3688);
nor U3811 (N_3811,N_3648,N_3557);
nor U3812 (N_3812,N_3685,N_3695);
nor U3813 (N_3813,N_3666,N_3583);
or U3814 (N_3814,N_3538,N_3507);
nor U3815 (N_3815,N_3664,N_3528);
or U3816 (N_3816,N_3692,N_3619);
nand U3817 (N_3817,N_3645,N_3652);
or U3818 (N_3818,N_3631,N_3618);
nand U3819 (N_3819,N_3690,N_3537);
nor U3820 (N_3820,N_3582,N_3734);
and U3821 (N_3821,N_3624,N_3546);
and U3822 (N_3822,N_3535,N_3597);
nand U3823 (N_3823,N_3598,N_3594);
xor U3824 (N_3824,N_3545,N_3591);
nand U3825 (N_3825,N_3705,N_3508);
nand U3826 (N_3826,N_3669,N_3628);
nand U3827 (N_3827,N_3554,N_3745);
xor U3828 (N_3828,N_3715,N_3703);
nand U3829 (N_3829,N_3717,N_3607);
or U3830 (N_3830,N_3532,N_3589);
or U3831 (N_3831,N_3707,N_3500);
nor U3832 (N_3832,N_3527,N_3724);
nor U3833 (N_3833,N_3588,N_3513);
or U3834 (N_3834,N_3658,N_3573);
nand U3835 (N_3835,N_3679,N_3544);
or U3836 (N_3836,N_3586,N_3706);
nand U3837 (N_3837,N_3559,N_3601);
and U3838 (N_3838,N_3524,N_3716);
xor U3839 (N_3839,N_3620,N_3510);
and U3840 (N_3840,N_3592,N_3697);
xor U3841 (N_3841,N_3639,N_3728);
nand U3842 (N_3842,N_3630,N_3747);
nor U3843 (N_3843,N_3677,N_3585);
and U3844 (N_3844,N_3533,N_3584);
and U3845 (N_3845,N_3699,N_3627);
nand U3846 (N_3846,N_3737,N_3718);
nand U3847 (N_3847,N_3644,N_3608);
and U3848 (N_3848,N_3651,N_3641);
nor U3849 (N_3849,N_3548,N_3661);
xnor U3850 (N_3850,N_3642,N_3733);
xnor U3851 (N_3851,N_3702,N_3660);
or U3852 (N_3852,N_3590,N_3647);
nor U3853 (N_3853,N_3730,N_3735);
and U3854 (N_3854,N_3530,N_3653);
and U3855 (N_3855,N_3657,N_3682);
nor U3856 (N_3856,N_3566,N_3689);
nor U3857 (N_3857,N_3540,N_3551);
nand U3858 (N_3858,N_3574,N_3609);
or U3859 (N_3859,N_3709,N_3531);
and U3860 (N_3860,N_3515,N_3712);
nand U3861 (N_3861,N_3576,N_3701);
or U3862 (N_3862,N_3562,N_3667);
or U3863 (N_3863,N_3742,N_3684);
and U3864 (N_3864,N_3522,N_3616);
nor U3865 (N_3865,N_3595,N_3746);
nor U3866 (N_3866,N_3577,N_3673);
nor U3867 (N_3867,N_3675,N_3731);
and U3868 (N_3868,N_3539,N_3600);
nand U3869 (N_3869,N_3578,N_3744);
nand U3870 (N_3870,N_3558,N_3615);
nand U3871 (N_3871,N_3605,N_3502);
nor U3872 (N_3872,N_3541,N_3693);
nor U3873 (N_3873,N_3659,N_3555);
xor U3874 (N_3874,N_3626,N_3603);
nor U3875 (N_3875,N_3741,N_3527);
nand U3876 (N_3876,N_3511,N_3654);
nor U3877 (N_3877,N_3628,N_3606);
nor U3878 (N_3878,N_3708,N_3685);
and U3879 (N_3879,N_3602,N_3541);
xnor U3880 (N_3880,N_3606,N_3666);
xor U3881 (N_3881,N_3726,N_3653);
nor U3882 (N_3882,N_3579,N_3677);
and U3883 (N_3883,N_3716,N_3665);
nor U3884 (N_3884,N_3678,N_3728);
nor U3885 (N_3885,N_3742,N_3565);
or U3886 (N_3886,N_3730,N_3521);
or U3887 (N_3887,N_3610,N_3542);
or U3888 (N_3888,N_3619,N_3572);
or U3889 (N_3889,N_3701,N_3682);
xnor U3890 (N_3890,N_3694,N_3651);
or U3891 (N_3891,N_3681,N_3606);
nand U3892 (N_3892,N_3508,N_3643);
nand U3893 (N_3893,N_3569,N_3536);
or U3894 (N_3894,N_3577,N_3625);
nand U3895 (N_3895,N_3723,N_3715);
or U3896 (N_3896,N_3627,N_3574);
or U3897 (N_3897,N_3563,N_3666);
or U3898 (N_3898,N_3699,N_3705);
and U3899 (N_3899,N_3747,N_3586);
or U3900 (N_3900,N_3693,N_3711);
or U3901 (N_3901,N_3686,N_3530);
nand U3902 (N_3902,N_3636,N_3595);
and U3903 (N_3903,N_3554,N_3555);
and U3904 (N_3904,N_3516,N_3624);
nor U3905 (N_3905,N_3746,N_3544);
and U3906 (N_3906,N_3664,N_3706);
and U3907 (N_3907,N_3696,N_3613);
xnor U3908 (N_3908,N_3744,N_3669);
or U3909 (N_3909,N_3536,N_3742);
or U3910 (N_3910,N_3593,N_3638);
and U3911 (N_3911,N_3628,N_3588);
or U3912 (N_3912,N_3503,N_3611);
nor U3913 (N_3913,N_3745,N_3542);
and U3914 (N_3914,N_3516,N_3676);
xnor U3915 (N_3915,N_3719,N_3660);
nor U3916 (N_3916,N_3613,N_3559);
nor U3917 (N_3917,N_3679,N_3525);
nor U3918 (N_3918,N_3663,N_3526);
or U3919 (N_3919,N_3532,N_3669);
and U3920 (N_3920,N_3684,N_3552);
xnor U3921 (N_3921,N_3734,N_3663);
nand U3922 (N_3922,N_3514,N_3643);
xnor U3923 (N_3923,N_3622,N_3702);
and U3924 (N_3924,N_3720,N_3625);
nand U3925 (N_3925,N_3573,N_3671);
nand U3926 (N_3926,N_3742,N_3747);
nor U3927 (N_3927,N_3621,N_3571);
nor U3928 (N_3928,N_3520,N_3671);
nand U3929 (N_3929,N_3558,N_3549);
nand U3930 (N_3930,N_3621,N_3636);
nand U3931 (N_3931,N_3550,N_3586);
and U3932 (N_3932,N_3613,N_3690);
xor U3933 (N_3933,N_3506,N_3640);
nand U3934 (N_3934,N_3634,N_3521);
and U3935 (N_3935,N_3685,N_3709);
or U3936 (N_3936,N_3682,N_3547);
nand U3937 (N_3937,N_3586,N_3605);
and U3938 (N_3938,N_3650,N_3686);
or U3939 (N_3939,N_3558,N_3617);
and U3940 (N_3940,N_3625,N_3705);
and U3941 (N_3941,N_3584,N_3597);
and U3942 (N_3942,N_3671,N_3740);
xnor U3943 (N_3943,N_3595,N_3516);
nor U3944 (N_3944,N_3555,N_3562);
nand U3945 (N_3945,N_3610,N_3574);
or U3946 (N_3946,N_3625,N_3559);
xnor U3947 (N_3947,N_3619,N_3649);
nand U3948 (N_3948,N_3523,N_3610);
and U3949 (N_3949,N_3552,N_3503);
nand U3950 (N_3950,N_3554,N_3546);
nand U3951 (N_3951,N_3630,N_3745);
nor U3952 (N_3952,N_3502,N_3505);
nand U3953 (N_3953,N_3519,N_3746);
and U3954 (N_3954,N_3575,N_3620);
or U3955 (N_3955,N_3743,N_3703);
and U3956 (N_3956,N_3681,N_3589);
nor U3957 (N_3957,N_3539,N_3687);
or U3958 (N_3958,N_3549,N_3574);
or U3959 (N_3959,N_3608,N_3564);
nand U3960 (N_3960,N_3641,N_3543);
nor U3961 (N_3961,N_3728,N_3614);
nand U3962 (N_3962,N_3570,N_3649);
nor U3963 (N_3963,N_3610,N_3516);
nand U3964 (N_3964,N_3676,N_3724);
nand U3965 (N_3965,N_3550,N_3531);
xnor U3966 (N_3966,N_3701,N_3631);
xnor U3967 (N_3967,N_3743,N_3500);
xor U3968 (N_3968,N_3627,N_3679);
or U3969 (N_3969,N_3739,N_3559);
or U3970 (N_3970,N_3506,N_3655);
and U3971 (N_3971,N_3576,N_3544);
nand U3972 (N_3972,N_3539,N_3683);
nor U3973 (N_3973,N_3683,N_3541);
nand U3974 (N_3974,N_3512,N_3700);
nor U3975 (N_3975,N_3735,N_3507);
nand U3976 (N_3976,N_3723,N_3642);
nand U3977 (N_3977,N_3638,N_3557);
nor U3978 (N_3978,N_3518,N_3606);
and U3979 (N_3979,N_3745,N_3703);
xor U3980 (N_3980,N_3613,N_3557);
nor U3981 (N_3981,N_3657,N_3624);
or U3982 (N_3982,N_3585,N_3630);
or U3983 (N_3983,N_3503,N_3647);
and U3984 (N_3984,N_3671,N_3576);
nand U3985 (N_3985,N_3731,N_3557);
nor U3986 (N_3986,N_3733,N_3573);
nor U3987 (N_3987,N_3627,N_3706);
or U3988 (N_3988,N_3576,N_3696);
nand U3989 (N_3989,N_3592,N_3580);
nor U3990 (N_3990,N_3706,N_3640);
nand U3991 (N_3991,N_3550,N_3699);
and U3992 (N_3992,N_3584,N_3519);
or U3993 (N_3993,N_3523,N_3696);
nand U3994 (N_3994,N_3663,N_3637);
nor U3995 (N_3995,N_3587,N_3554);
nand U3996 (N_3996,N_3747,N_3500);
nor U3997 (N_3997,N_3602,N_3593);
and U3998 (N_3998,N_3705,N_3581);
xnor U3999 (N_3999,N_3642,N_3562);
or U4000 (N_4000,N_3872,N_3878);
or U4001 (N_4001,N_3943,N_3805);
or U4002 (N_4002,N_3856,N_3893);
or U4003 (N_4003,N_3808,N_3799);
or U4004 (N_4004,N_3840,N_3790);
nand U4005 (N_4005,N_3863,N_3947);
or U4006 (N_4006,N_3951,N_3935);
xor U4007 (N_4007,N_3940,N_3980);
nand U4008 (N_4008,N_3802,N_3798);
nor U4009 (N_4009,N_3841,N_3931);
xor U4010 (N_4010,N_3792,N_3838);
nor U4011 (N_4011,N_3864,N_3993);
nand U4012 (N_4012,N_3787,N_3986);
xnor U4013 (N_4013,N_3826,N_3967);
nand U4014 (N_4014,N_3906,N_3887);
or U4015 (N_4015,N_3877,N_3773);
and U4016 (N_4016,N_3825,N_3903);
and U4017 (N_4017,N_3891,N_3890);
nand U4018 (N_4018,N_3859,N_3937);
xor U4019 (N_4019,N_3844,N_3982);
nor U4020 (N_4020,N_3954,N_3833);
and U4021 (N_4021,N_3981,N_3973);
nor U4022 (N_4022,N_3902,N_3865);
xnor U4023 (N_4023,N_3920,N_3882);
and U4024 (N_4024,N_3901,N_3997);
nor U4025 (N_4025,N_3999,N_3950);
nor U4026 (N_4026,N_3911,N_3928);
and U4027 (N_4027,N_3813,N_3765);
nor U4028 (N_4028,N_3834,N_3794);
and U4029 (N_4029,N_3975,N_3827);
nor U4030 (N_4030,N_3884,N_3946);
or U4031 (N_4031,N_3914,N_3912);
nor U4032 (N_4032,N_3924,N_3953);
xnor U4033 (N_4033,N_3754,N_3839);
and U4034 (N_4034,N_3803,N_3855);
or U4035 (N_4035,N_3910,N_3780);
nand U4036 (N_4036,N_3849,N_3806);
nand U4037 (N_4037,N_3857,N_3752);
xor U4038 (N_4038,N_3976,N_3934);
nand U4039 (N_4039,N_3768,N_3845);
and U4040 (N_4040,N_3847,N_3883);
nand U4041 (N_4041,N_3867,N_3918);
nor U4042 (N_4042,N_3835,N_3843);
nor U4043 (N_4043,N_3944,N_3995);
xor U4044 (N_4044,N_3945,N_3783);
or U4045 (N_4045,N_3930,N_3786);
nand U4046 (N_4046,N_3971,N_3756);
nand U4047 (N_4047,N_3926,N_3992);
or U4048 (N_4048,N_3774,N_3972);
nor U4049 (N_4049,N_3956,N_3896);
nor U4050 (N_4050,N_3764,N_3824);
or U4051 (N_4051,N_3990,N_3957);
and U4052 (N_4052,N_3758,N_3929);
nand U4053 (N_4053,N_3797,N_3988);
and U4054 (N_4054,N_3819,N_3942);
or U4055 (N_4055,N_3842,N_3895);
or U4056 (N_4056,N_3941,N_3804);
or U4057 (N_4057,N_3948,N_3927);
and U4058 (N_4058,N_3828,N_3860);
and U4059 (N_4059,N_3770,N_3791);
and U4060 (N_4060,N_3757,N_3868);
or U4061 (N_4061,N_3955,N_3753);
nor U4062 (N_4062,N_3899,N_3919);
nand U4063 (N_4063,N_3760,N_3885);
nor U4064 (N_4064,N_3831,N_3852);
or U4065 (N_4065,N_3905,N_3952);
nor U4066 (N_4066,N_3904,N_3888);
or U4067 (N_4067,N_3858,N_3932);
xor U4068 (N_4068,N_3894,N_3866);
and U4069 (N_4069,N_3820,N_3966);
and U4070 (N_4070,N_3854,N_3875);
or U4071 (N_4071,N_3936,N_3889);
xnor U4072 (N_4072,N_3968,N_3830);
nand U4073 (N_4073,N_3969,N_3994);
or U4074 (N_4074,N_3874,N_3816);
nand U4075 (N_4075,N_3811,N_3836);
or U4076 (N_4076,N_3818,N_3892);
or U4077 (N_4077,N_3881,N_3822);
nand U4078 (N_4078,N_3989,N_3909);
and U4079 (N_4079,N_3978,N_3761);
and U4080 (N_4080,N_3755,N_3751);
or U4081 (N_4081,N_3987,N_3962);
or U4082 (N_4082,N_3938,N_3795);
or U4083 (N_4083,N_3823,N_3861);
or U4084 (N_4084,N_3829,N_3977);
nor U4085 (N_4085,N_3789,N_3897);
nand U4086 (N_4086,N_3913,N_3873);
nand U4087 (N_4087,N_3851,N_3772);
nor U4088 (N_4088,N_3915,N_3961);
nor U4089 (N_4089,N_3782,N_3776);
nand U4090 (N_4090,N_3763,N_3846);
nor U4091 (N_4091,N_3779,N_3777);
and U4092 (N_4092,N_3917,N_3898);
or U4093 (N_4093,N_3809,N_3817);
and U4094 (N_4094,N_3921,N_3964);
and U4095 (N_4095,N_3862,N_3869);
nor U4096 (N_4096,N_3750,N_3985);
nand U4097 (N_4097,N_3771,N_3810);
or U4098 (N_4098,N_3949,N_3886);
and U4099 (N_4099,N_3815,N_3916);
nand U4100 (N_4100,N_3970,N_3963);
or U4101 (N_4101,N_3974,N_3832);
nor U4102 (N_4102,N_3960,N_3759);
nor U4103 (N_4103,N_3979,N_3933);
nor U4104 (N_4104,N_3991,N_3923);
or U4105 (N_4105,N_3853,N_3796);
nand U4106 (N_4106,N_3925,N_3922);
or U4107 (N_4107,N_3784,N_3837);
nor U4108 (N_4108,N_3907,N_3939);
or U4109 (N_4109,N_3801,N_3800);
or U4110 (N_4110,N_3876,N_3778);
xor U4111 (N_4111,N_3984,N_3958);
nor U4112 (N_4112,N_3781,N_3793);
or U4113 (N_4113,N_3879,N_3965);
and U4114 (N_4114,N_3767,N_3983);
nor U4115 (N_4115,N_3766,N_3996);
and U4116 (N_4116,N_3870,N_3769);
nor U4117 (N_4117,N_3807,N_3788);
and U4118 (N_4118,N_3775,N_3908);
and U4119 (N_4119,N_3871,N_3812);
or U4120 (N_4120,N_3762,N_3814);
nand U4121 (N_4121,N_3821,N_3785);
or U4122 (N_4122,N_3959,N_3998);
nand U4123 (N_4123,N_3850,N_3880);
or U4124 (N_4124,N_3848,N_3900);
nand U4125 (N_4125,N_3797,N_3854);
and U4126 (N_4126,N_3867,N_3758);
and U4127 (N_4127,N_3761,N_3788);
xor U4128 (N_4128,N_3810,N_3968);
and U4129 (N_4129,N_3975,N_3756);
or U4130 (N_4130,N_3835,N_3955);
nor U4131 (N_4131,N_3854,N_3788);
or U4132 (N_4132,N_3834,N_3994);
nor U4133 (N_4133,N_3865,N_3798);
and U4134 (N_4134,N_3970,N_3973);
and U4135 (N_4135,N_3974,N_3896);
and U4136 (N_4136,N_3997,N_3753);
nand U4137 (N_4137,N_3844,N_3961);
xnor U4138 (N_4138,N_3923,N_3970);
or U4139 (N_4139,N_3894,N_3845);
or U4140 (N_4140,N_3926,N_3938);
nor U4141 (N_4141,N_3843,N_3819);
or U4142 (N_4142,N_3841,N_3797);
nand U4143 (N_4143,N_3938,N_3762);
nand U4144 (N_4144,N_3905,N_3896);
xor U4145 (N_4145,N_3908,N_3816);
or U4146 (N_4146,N_3988,N_3990);
nand U4147 (N_4147,N_3881,N_3928);
xor U4148 (N_4148,N_3978,N_3988);
nor U4149 (N_4149,N_3884,N_3860);
and U4150 (N_4150,N_3835,N_3761);
and U4151 (N_4151,N_3901,N_3920);
nor U4152 (N_4152,N_3842,N_3799);
nor U4153 (N_4153,N_3898,N_3972);
and U4154 (N_4154,N_3953,N_3857);
nand U4155 (N_4155,N_3816,N_3854);
nand U4156 (N_4156,N_3771,N_3977);
nor U4157 (N_4157,N_3869,N_3951);
and U4158 (N_4158,N_3762,N_3980);
xor U4159 (N_4159,N_3933,N_3846);
and U4160 (N_4160,N_3888,N_3929);
nor U4161 (N_4161,N_3752,N_3924);
and U4162 (N_4162,N_3801,N_3970);
xnor U4163 (N_4163,N_3922,N_3834);
and U4164 (N_4164,N_3811,N_3826);
and U4165 (N_4165,N_3939,N_3801);
and U4166 (N_4166,N_3869,N_3860);
nor U4167 (N_4167,N_3799,N_3821);
and U4168 (N_4168,N_3787,N_3925);
xnor U4169 (N_4169,N_3826,N_3773);
and U4170 (N_4170,N_3968,N_3890);
xnor U4171 (N_4171,N_3873,N_3882);
nand U4172 (N_4172,N_3896,N_3939);
or U4173 (N_4173,N_3987,N_3776);
and U4174 (N_4174,N_3915,N_3951);
nor U4175 (N_4175,N_3788,N_3992);
or U4176 (N_4176,N_3785,N_3765);
or U4177 (N_4177,N_3766,N_3895);
nand U4178 (N_4178,N_3888,N_3882);
or U4179 (N_4179,N_3753,N_3798);
and U4180 (N_4180,N_3751,N_3901);
or U4181 (N_4181,N_3995,N_3835);
nand U4182 (N_4182,N_3793,N_3942);
or U4183 (N_4183,N_3990,N_3947);
nor U4184 (N_4184,N_3768,N_3963);
nor U4185 (N_4185,N_3785,N_3816);
nor U4186 (N_4186,N_3991,N_3987);
nor U4187 (N_4187,N_3813,N_3957);
nand U4188 (N_4188,N_3882,N_3918);
nor U4189 (N_4189,N_3918,N_3883);
nand U4190 (N_4190,N_3842,N_3984);
xnor U4191 (N_4191,N_3915,N_3752);
nor U4192 (N_4192,N_3886,N_3874);
and U4193 (N_4193,N_3796,N_3888);
nor U4194 (N_4194,N_3891,N_3819);
nor U4195 (N_4195,N_3938,N_3880);
or U4196 (N_4196,N_3787,N_3902);
xor U4197 (N_4197,N_3755,N_3969);
or U4198 (N_4198,N_3758,N_3936);
nand U4199 (N_4199,N_3773,N_3786);
or U4200 (N_4200,N_3766,N_3828);
nor U4201 (N_4201,N_3930,N_3988);
nor U4202 (N_4202,N_3770,N_3915);
xor U4203 (N_4203,N_3816,N_3803);
or U4204 (N_4204,N_3782,N_3887);
or U4205 (N_4205,N_3802,N_3750);
nor U4206 (N_4206,N_3793,N_3910);
or U4207 (N_4207,N_3833,N_3835);
and U4208 (N_4208,N_3874,N_3977);
xnor U4209 (N_4209,N_3800,N_3978);
and U4210 (N_4210,N_3974,N_3856);
or U4211 (N_4211,N_3919,N_3787);
nor U4212 (N_4212,N_3885,N_3955);
nor U4213 (N_4213,N_3953,N_3866);
nand U4214 (N_4214,N_3912,N_3805);
and U4215 (N_4215,N_3854,N_3970);
or U4216 (N_4216,N_3776,N_3837);
and U4217 (N_4217,N_3945,N_3831);
nand U4218 (N_4218,N_3817,N_3825);
and U4219 (N_4219,N_3952,N_3960);
nand U4220 (N_4220,N_3862,N_3994);
nor U4221 (N_4221,N_3752,N_3751);
and U4222 (N_4222,N_3875,N_3785);
or U4223 (N_4223,N_3754,N_3797);
xnor U4224 (N_4224,N_3781,N_3962);
and U4225 (N_4225,N_3893,N_3778);
nor U4226 (N_4226,N_3798,N_3787);
nor U4227 (N_4227,N_3782,N_3758);
nor U4228 (N_4228,N_3923,N_3932);
and U4229 (N_4229,N_3842,N_3827);
and U4230 (N_4230,N_3903,N_3790);
nor U4231 (N_4231,N_3940,N_3853);
nor U4232 (N_4232,N_3755,N_3797);
nor U4233 (N_4233,N_3756,N_3833);
nand U4234 (N_4234,N_3903,N_3883);
and U4235 (N_4235,N_3775,N_3946);
nor U4236 (N_4236,N_3896,N_3838);
xnor U4237 (N_4237,N_3867,N_3860);
nand U4238 (N_4238,N_3914,N_3757);
or U4239 (N_4239,N_3986,N_3852);
and U4240 (N_4240,N_3758,N_3786);
or U4241 (N_4241,N_3763,N_3999);
nor U4242 (N_4242,N_3763,N_3833);
nor U4243 (N_4243,N_3925,N_3803);
and U4244 (N_4244,N_3990,N_3763);
nand U4245 (N_4245,N_3824,N_3752);
or U4246 (N_4246,N_3878,N_3998);
nor U4247 (N_4247,N_3819,N_3758);
nor U4248 (N_4248,N_3841,N_3883);
nor U4249 (N_4249,N_3950,N_3855);
nor U4250 (N_4250,N_4117,N_4027);
or U4251 (N_4251,N_4131,N_4119);
nor U4252 (N_4252,N_4014,N_4082);
and U4253 (N_4253,N_4056,N_4174);
or U4254 (N_4254,N_4102,N_4028);
nor U4255 (N_4255,N_4228,N_4158);
xnor U4256 (N_4256,N_4184,N_4035);
and U4257 (N_4257,N_4021,N_4142);
nand U4258 (N_4258,N_4114,N_4006);
or U4259 (N_4259,N_4019,N_4076);
or U4260 (N_4260,N_4176,N_4079);
nand U4261 (N_4261,N_4078,N_4236);
and U4262 (N_4262,N_4081,N_4206);
nor U4263 (N_4263,N_4179,N_4189);
and U4264 (N_4264,N_4048,N_4151);
nor U4265 (N_4265,N_4045,N_4138);
and U4266 (N_4266,N_4002,N_4003);
nor U4267 (N_4267,N_4197,N_4192);
nand U4268 (N_4268,N_4169,N_4153);
nand U4269 (N_4269,N_4000,N_4004);
xor U4270 (N_4270,N_4108,N_4230);
xor U4271 (N_4271,N_4055,N_4245);
nor U4272 (N_4272,N_4183,N_4188);
and U4273 (N_4273,N_4135,N_4218);
and U4274 (N_4274,N_4011,N_4080);
nor U4275 (N_4275,N_4094,N_4084);
or U4276 (N_4276,N_4034,N_4193);
nand U4277 (N_4277,N_4167,N_4017);
or U4278 (N_4278,N_4064,N_4009);
nor U4279 (N_4279,N_4145,N_4171);
nor U4280 (N_4280,N_4132,N_4224);
and U4281 (N_4281,N_4246,N_4057);
or U4282 (N_4282,N_4225,N_4186);
or U4283 (N_4283,N_4140,N_4178);
or U4284 (N_4284,N_4089,N_4065);
or U4285 (N_4285,N_4198,N_4097);
or U4286 (N_4286,N_4166,N_4243);
nor U4287 (N_4287,N_4182,N_4205);
or U4288 (N_4288,N_4038,N_4195);
and U4289 (N_4289,N_4058,N_4149);
nand U4290 (N_4290,N_4073,N_4180);
and U4291 (N_4291,N_4051,N_4147);
and U4292 (N_4292,N_4042,N_4077);
nor U4293 (N_4293,N_4146,N_4024);
and U4294 (N_4294,N_4120,N_4063);
or U4295 (N_4295,N_4227,N_4143);
or U4296 (N_4296,N_4249,N_4122);
and U4297 (N_4297,N_4223,N_4157);
or U4298 (N_4298,N_4110,N_4068);
xor U4299 (N_4299,N_4026,N_4125);
or U4300 (N_4300,N_4099,N_4204);
and U4301 (N_4301,N_4163,N_4177);
or U4302 (N_4302,N_4067,N_4098);
xor U4303 (N_4303,N_4118,N_4032);
or U4304 (N_4304,N_4010,N_4015);
nand U4305 (N_4305,N_4170,N_4112);
nand U4306 (N_4306,N_4164,N_4020);
or U4307 (N_4307,N_4095,N_4106);
or U4308 (N_4308,N_4066,N_4093);
or U4309 (N_4309,N_4185,N_4181);
or U4310 (N_4310,N_4041,N_4115);
nand U4311 (N_4311,N_4231,N_4159);
nor U4312 (N_4312,N_4005,N_4072);
and U4313 (N_4313,N_4237,N_4070);
nor U4314 (N_4314,N_4203,N_4054);
nand U4315 (N_4315,N_4071,N_4124);
or U4316 (N_4316,N_4133,N_4136);
nand U4317 (N_4317,N_4012,N_4216);
and U4318 (N_4318,N_4208,N_4105);
and U4319 (N_4319,N_4202,N_4085);
nor U4320 (N_4320,N_4060,N_4104);
or U4321 (N_4321,N_4239,N_4199);
and U4322 (N_4322,N_4008,N_4226);
nor U4323 (N_4323,N_4049,N_4156);
nor U4324 (N_4324,N_4052,N_4129);
xor U4325 (N_4325,N_4152,N_4241);
or U4326 (N_4326,N_4137,N_4123);
and U4327 (N_4327,N_4150,N_4144);
and U4328 (N_4328,N_4059,N_4130);
nor U4329 (N_4329,N_4212,N_4083);
or U4330 (N_4330,N_4211,N_4061);
or U4331 (N_4331,N_4096,N_4221);
and U4332 (N_4332,N_4215,N_4107);
nand U4333 (N_4333,N_4175,N_4030);
or U4334 (N_4334,N_4191,N_4037);
xor U4335 (N_4335,N_4207,N_4187);
or U4336 (N_4336,N_4190,N_4141);
nor U4337 (N_4337,N_4214,N_4062);
nand U4338 (N_4338,N_4162,N_4222);
nand U4339 (N_4339,N_4160,N_4007);
xnor U4340 (N_4340,N_4116,N_4016);
xnor U4341 (N_4341,N_4023,N_4217);
xnor U4342 (N_4342,N_4113,N_4047);
and U4343 (N_4343,N_4154,N_4039);
xor U4344 (N_4344,N_4242,N_4139);
nand U4345 (N_4345,N_4234,N_4069);
nor U4346 (N_4346,N_4018,N_4235);
nor U4347 (N_4347,N_4075,N_4155);
and U4348 (N_4348,N_4092,N_4161);
and U4349 (N_4349,N_4134,N_4050);
and U4350 (N_4350,N_4238,N_4173);
nor U4351 (N_4351,N_4046,N_4091);
xnor U4352 (N_4352,N_4240,N_4232);
or U4353 (N_4353,N_4033,N_4088);
and U4354 (N_4354,N_4087,N_4165);
and U4355 (N_4355,N_4148,N_4111);
nand U4356 (N_4356,N_4127,N_4194);
nand U4357 (N_4357,N_4220,N_4036);
nand U4358 (N_4358,N_4025,N_4040);
and U4359 (N_4359,N_4200,N_4090);
or U4360 (N_4360,N_4086,N_4168);
or U4361 (N_4361,N_4128,N_4126);
or U4362 (N_4362,N_4209,N_4013);
nor U4363 (N_4363,N_4213,N_4043);
nor U4364 (N_4364,N_4201,N_4247);
and U4365 (N_4365,N_4229,N_4031);
or U4366 (N_4366,N_4001,N_4053);
nor U4367 (N_4367,N_4233,N_4100);
nor U4368 (N_4368,N_4074,N_4044);
nor U4369 (N_4369,N_4103,N_4244);
or U4370 (N_4370,N_4121,N_4248);
and U4371 (N_4371,N_4101,N_4210);
or U4372 (N_4372,N_4022,N_4109);
and U4373 (N_4373,N_4029,N_4219);
and U4374 (N_4374,N_4172,N_4196);
or U4375 (N_4375,N_4117,N_4003);
and U4376 (N_4376,N_4152,N_4134);
nand U4377 (N_4377,N_4202,N_4225);
nand U4378 (N_4378,N_4137,N_4144);
and U4379 (N_4379,N_4224,N_4099);
and U4380 (N_4380,N_4149,N_4151);
and U4381 (N_4381,N_4236,N_4111);
or U4382 (N_4382,N_4047,N_4230);
or U4383 (N_4383,N_4071,N_4117);
nor U4384 (N_4384,N_4237,N_4152);
xor U4385 (N_4385,N_4010,N_4020);
nand U4386 (N_4386,N_4167,N_4025);
or U4387 (N_4387,N_4061,N_4066);
xnor U4388 (N_4388,N_4117,N_4113);
and U4389 (N_4389,N_4039,N_4076);
and U4390 (N_4390,N_4062,N_4157);
and U4391 (N_4391,N_4224,N_4036);
nand U4392 (N_4392,N_4058,N_4086);
and U4393 (N_4393,N_4046,N_4126);
or U4394 (N_4394,N_4186,N_4118);
nand U4395 (N_4395,N_4243,N_4083);
and U4396 (N_4396,N_4201,N_4182);
and U4397 (N_4397,N_4077,N_4143);
nand U4398 (N_4398,N_4172,N_4179);
and U4399 (N_4399,N_4074,N_4028);
or U4400 (N_4400,N_4241,N_4072);
nand U4401 (N_4401,N_4215,N_4236);
nand U4402 (N_4402,N_4115,N_4227);
xnor U4403 (N_4403,N_4044,N_4212);
and U4404 (N_4404,N_4054,N_4060);
nand U4405 (N_4405,N_4237,N_4174);
nor U4406 (N_4406,N_4069,N_4106);
nor U4407 (N_4407,N_4013,N_4023);
and U4408 (N_4408,N_4050,N_4090);
and U4409 (N_4409,N_4048,N_4132);
nand U4410 (N_4410,N_4021,N_4151);
or U4411 (N_4411,N_4198,N_4164);
and U4412 (N_4412,N_4020,N_4182);
and U4413 (N_4413,N_4196,N_4033);
and U4414 (N_4414,N_4044,N_4157);
nor U4415 (N_4415,N_4089,N_4211);
or U4416 (N_4416,N_4191,N_4163);
or U4417 (N_4417,N_4079,N_4033);
nor U4418 (N_4418,N_4110,N_4001);
nand U4419 (N_4419,N_4243,N_4155);
and U4420 (N_4420,N_4128,N_4087);
nor U4421 (N_4421,N_4237,N_4004);
and U4422 (N_4422,N_4142,N_4215);
or U4423 (N_4423,N_4015,N_4211);
nor U4424 (N_4424,N_4192,N_4176);
nand U4425 (N_4425,N_4232,N_4007);
nand U4426 (N_4426,N_4241,N_4134);
or U4427 (N_4427,N_4085,N_4223);
or U4428 (N_4428,N_4012,N_4037);
nand U4429 (N_4429,N_4177,N_4130);
or U4430 (N_4430,N_4093,N_4182);
nand U4431 (N_4431,N_4123,N_4071);
or U4432 (N_4432,N_4162,N_4106);
nor U4433 (N_4433,N_4061,N_4121);
nand U4434 (N_4434,N_4180,N_4100);
or U4435 (N_4435,N_4124,N_4006);
and U4436 (N_4436,N_4037,N_4022);
nor U4437 (N_4437,N_4110,N_4048);
and U4438 (N_4438,N_4016,N_4159);
and U4439 (N_4439,N_4166,N_4171);
or U4440 (N_4440,N_4050,N_4213);
and U4441 (N_4441,N_4088,N_4133);
nor U4442 (N_4442,N_4081,N_4129);
and U4443 (N_4443,N_4035,N_4102);
nand U4444 (N_4444,N_4249,N_4153);
and U4445 (N_4445,N_4221,N_4235);
or U4446 (N_4446,N_4054,N_4055);
nor U4447 (N_4447,N_4200,N_4244);
and U4448 (N_4448,N_4098,N_4041);
or U4449 (N_4449,N_4208,N_4152);
and U4450 (N_4450,N_4053,N_4079);
nor U4451 (N_4451,N_4081,N_4115);
nor U4452 (N_4452,N_4224,N_4064);
nor U4453 (N_4453,N_4095,N_4091);
nand U4454 (N_4454,N_4204,N_4078);
nand U4455 (N_4455,N_4225,N_4174);
or U4456 (N_4456,N_4054,N_4129);
nand U4457 (N_4457,N_4245,N_4086);
nor U4458 (N_4458,N_4157,N_4103);
or U4459 (N_4459,N_4139,N_4151);
nor U4460 (N_4460,N_4184,N_4213);
and U4461 (N_4461,N_4101,N_4100);
or U4462 (N_4462,N_4095,N_4002);
or U4463 (N_4463,N_4141,N_4233);
xor U4464 (N_4464,N_4238,N_4112);
xnor U4465 (N_4465,N_4035,N_4134);
xnor U4466 (N_4466,N_4227,N_4199);
xnor U4467 (N_4467,N_4190,N_4037);
nand U4468 (N_4468,N_4008,N_4126);
and U4469 (N_4469,N_4228,N_4128);
nand U4470 (N_4470,N_4234,N_4160);
nor U4471 (N_4471,N_4084,N_4010);
nor U4472 (N_4472,N_4028,N_4101);
or U4473 (N_4473,N_4027,N_4199);
nor U4474 (N_4474,N_4004,N_4045);
and U4475 (N_4475,N_4168,N_4116);
and U4476 (N_4476,N_4158,N_4196);
xnor U4477 (N_4477,N_4174,N_4051);
nor U4478 (N_4478,N_4011,N_4118);
nand U4479 (N_4479,N_4221,N_4129);
and U4480 (N_4480,N_4248,N_4144);
or U4481 (N_4481,N_4031,N_4011);
or U4482 (N_4482,N_4185,N_4029);
and U4483 (N_4483,N_4019,N_4103);
nor U4484 (N_4484,N_4001,N_4097);
or U4485 (N_4485,N_4176,N_4172);
or U4486 (N_4486,N_4152,N_4094);
xor U4487 (N_4487,N_4207,N_4176);
or U4488 (N_4488,N_4101,N_4116);
xor U4489 (N_4489,N_4144,N_4102);
xnor U4490 (N_4490,N_4247,N_4000);
nor U4491 (N_4491,N_4051,N_4187);
nor U4492 (N_4492,N_4107,N_4147);
nand U4493 (N_4493,N_4077,N_4228);
xnor U4494 (N_4494,N_4024,N_4121);
and U4495 (N_4495,N_4179,N_4003);
and U4496 (N_4496,N_4049,N_4062);
and U4497 (N_4497,N_4171,N_4089);
nand U4498 (N_4498,N_4175,N_4228);
nand U4499 (N_4499,N_4246,N_4172);
and U4500 (N_4500,N_4399,N_4499);
xor U4501 (N_4501,N_4268,N_4324);
nor U4502 (N_4502,N_4252,N_4352);
nor U4503 (N_4503,N_4262,N_4431);
or U4504 (N_4504,N_4486,N_4373);
or U4505 (N_4505,N_4314,N_4384);
or U4506 (N_4506,N_4250,N_4468);
nand U4507 (N_4507,N_4488,N_4365);
xnor U4508 (N_4508,N_4329,N_4278);
nand U4509 (N_4509,N_4267,N_4328);
and U4510 (N_4510,N_4393,N_4427);
xnor U4511 (N_4511,N_4439,N_4382);
or U4512 (N_4512,N_4291,N_4321);
or U4513 (N_4513,N_4317,N_4490);
and U4514 (N_4514,N_4419,N_4425);
and U4515 (N_4515,N_4454,N_4369);
and U4516 (N_4516,N_4270,N_4397);
or U4517 (N_4517,N_4361,N_4390);
or U4518 (N_4518,N_4303,N_4379);
and U4519 (N_4519,N_4304,N_4280);
or U4520 (N_4520,N_4380,N_4484);
nand U4521 (N_4521,N_4335,N_4357);
or U4522 (N_4522,N_4482,N_4414);
nand U4523 (N_4523,N_4338,N_4334);
or U4524 (N_4524,N_4487,N_4356);
and U4525 (N_4525,N_4446,N_4496);
or U4526 (N_4526,N_4322,N_4353);
xor U4527 (N_4527,N_4387,N_4416);
and U4528 (N_4528,N_4288,N_4445);
nor U4529 (N_4529,N_4421,N_4358);
or U4530 (N_4530,N_4481,N_4308);
or U4531 (N_4531,N_4346,N_4343);
or U4532 (N_4532,N_4271,N_4437);
and U4533 (N_4533,N_4377,N_4438);
nand U4534 (N_4534,N_4277,N_4279);
nand U4535 (N_4535,N_4348,N_4312);
or U4536 (N_4536,N_4261,N_4441);
or U4537 (N_4537,N_4259,N_4459);
nor U4538 (N_4538,N_4444,N_4404);
or U4539 (N_4539,N_4287,N_4294);
nor U4540 (N_4540,N_4360,N_4396);
or U4541 (N_4541,N_4363,N_4429);
nand U4542 (N_4542,N_4462,N_4333);
xor U4543 (N_4543,N_4350,N_4285);
or U4544 (N_4544,N_4465,N_4415);
nor U4545 (N_4545,N_4264,N_4275);
or U4546 (N_4546,N_4448,N_4455);
xnor U4547 (N_4547,N_4469,N_4319);
or U4548 (N_4548,N_4283,N_4458);
and U4549 (N_4549,N_4491,N_4394);
and U4550 (N_4550,N_4495,N_4493);
and U4551 (N_4551,N_4383,N_4436);
nand U4552 (N_4552,N_4432,N_4286);
nor U4553 (N_4553,N_4476,N_4412);
or U4554 (N_4554,N_4260,N_4310);
and U4555 (N_4555,N_4435,N_4418);
nor U4556 (N_4556,N_4355,N_4354);
or U4557 (N_4557,N_4479,N_4344);
xnor U4558 (N_4558,N_4424,N_4385);
or U4559 (N_4559,N_4320,N_4254);
and U4560 (N_4560,N_4461,N_4265);
or U4561 (N_4561,N_4290,N_4256);
nor U4562 (N_4562,N_4306,N_4295);
or U4563 (N_4563,N_4400,N_4451);
or U4564 (N_4564,N_4410,N_4388);
nor U4565 (N_4565,N_4340,N_4473);
and U4566 (N_4566,N_4330,N_4318);
or U4567 (N_4567,N_4342,N_4475);
nor U4568 (N_4568,N_4366,N_4457);
and U4569 (N_4569,N_4339,N_4362);
nor U4570 (N_4570,N_4297,N_4422);
nand U4571 (N_4571,N_4299,N_4443);
and U4572 (N_4572,N_4258,N_4257);
nand U4573 (N_4573,N_4313,N_4347);
or U4574 (N_4574,N_4472,N_4309);
nand U4575 (N_4575,N_4426,N_4368);
and U4576 (N_4576,N_4289,N_4401);
or U4577 (N_4577,N_4316,N_4349);
and U4578 (N_4578,N_4452,N_4332);
or U4579 (N_4579,N_4282,N_4315);
nand U4580 (N_4580,N_4351,N_4375);
and U4581 (N_4581,N_4371,N_4440);
and U4582 (N_4582,N_4428,N_4374);
or U4583 (N_4583,N_4274,N_4325);
and U4584 (N_4584,N_4447,N_4483);
and U4585 (N_4585,N_4359,N_4434);
and U4586 (N_4586,N_4301,N_4417);
and U4587 (N_4587,N_4272,N_4389);
or U4588 (N_4588,N_4407,N_4485);
nand U4589 (N_4589,N_4292,N_4391);
or U4590 (N_4590,N_4463,N_4253);
nand U4591 (N_4591,N_4456,N_4423);
and U4592 (N_4592,N_4266,N_4326);
xor U4593 (N_4593,N_4386,N_4413);
nor U4594 (N_4594,N_4494,N_4269);
nand U4595 (N_4595,N_4395,N_4449);
xor U4596 (N_4596,N_4281,N_4466);
xnor U4597 (N_4597,N_4311,N_4403);
nor U4598 (N_4598,N_4398,N_4376);
and U4599 (N_4599,N_4497,N_4470);
nor U4600 (N_4600,N_4341,N_4450);
and U4601 (N_4601,N_4323,N_4336);
xor U4602 (N_4602,N_4255,N_4442);
nand U4603 (N_4603,N_4331,N_4433);
nand U4604 (N_4604,N_4302,N_4345);
nor U4605 (N_4605,N_4409,N_4477);
or U4606 (N_4606,N_4337,N_4467);
nor U4607 (N_4607,N_4464,N_4305);
nand U4608 (N_4608,N_4471,N_4284);
and U4609 (N_4609,N_4293,N_4367);
or U4610 (N_4610,N_4381,N_4478);
nor U4611 (N_4611,N_4298,N_4402);
nor U4612 (N_4612,N_4378,N_4296);
nand U4613 (N_4613,N_4251,N_4411);
or U4614 (N_4614,N_4480,N_4372);
or U4615 (N_4615,N_4392,N_4364);
nor U4616 (N_4616,N_4300,N_4408);
nand U4617 (N_4617,N_4498,N_4263);
nor U4618 (N_4618,N_4327,N_4276);
nand U4619 (N_4619,N_4406,N_4453);
xnor U4620 (N_4620,N_4307,N_4430);
nor U4621 (N_4621,N_4489,N_4492);
nor U4622 (N_4622,N_4370,N_4420);
nor U4623 (N_4623,N_4474,N_4405);
nor U4624 (N_4624,N_4273,N_4460);
or U4625 (N_4625,N_4359,N_4255);
nand U4626 (N_4626,N_4273,N_4325);
nor U4627 (N_4627,N_4415,N_4275);
nor U4628 (N_4628,N_4331,N_4258);
and U4629 (N_4629,N_4473,N_4343);
or U4630 (N_4630,N_4254,N_4309);
and U4631 (N_4631,N_4355,N_4261);
nor U4632 (N_4632,N_4333,N_4477);
and U4633 (N_4633,N_4265,N_4260);
or U4634 (N_4634,N_4451,N_4429);
nor U4635 (N_4635,N_4414,N_4418);
nand U4636 (N_4636,N_4354,N_4311);
and U4637 (N_4637,N_4309,N_4370);
xor U4638 (N_4638,N_4482,N_4302);
or U4639 (N_4639,N_4467,N_4317);
nor U4640 (N_4640,N_4373,N_4261);
nand U4641 (N_4641,N_4311,N_4343);
nand U4642 (N_4642,N_4486,N_4267);
or U4643 (N_4643,N_4447,N_4484);
or U4644 (N_4644,N_4378,N_4317);
and U4645 (N_4645,N_4314,N_4493);
nand U4646 (N_4646,N_4447,N_4303);
or U4647 (N_4647,N_4326,N_4487);
or U4648 (N_4648,N_4442,N_4365);
nor U4649 (N_4649,N_4335,N_4422);
or U4650 (N_4650,N_4354,N_4463);
or U4651 (N_4651,N_4486,N_4391);
xor U4652 (N_4652,N_4463,N_4362);
nand U4653 (N_4653,N_4347,N_4420);
and U4654 (N_4654,N_4373,N_4414);
or U4655 (N_4655,N_4479,N_4478);
nor U4656 (N_4656,N_4404,N_4467);
nand U4657 (N_4657,N_4416,N_4352);
nor U4658 (N_4658,N_4399,N_4270);
and U4659 (N_4659,N_4349,N_4318);
or U4660 (N_4660,N_4434,N_4441);
nor U4661 (N_4661,N_4439,N_4385);
nor U4662 (N_4662,N_4373,N_4251);
or U4663 (N_4663,N_4495,N_4264);
and U4664 (N_4664,N_4366,N_4251);
or U4665 (N_4665,N_4257,N_4495);
and U4666 (N_4666,N_4280,N_4496);
and U4667 (N_4667,N_4325,N_4348);
or U4668 (N_4668,N_4403,N_4350);
or U4669 (N_4669,N_4384,N_4305);
and U4670 (N_4670,N_4261,N_4315);
and U4671 (N_4671,N_4302,N_4400);
nor U4672 (N_4672,N_4438,N_4284);
nor U4673 (N_4673,N_4315,N_4376);
xnor U4674 (N_4674,N_4388,N_4457);
or U4675 (N_4675,N_4401,N_4462);
nor U4676 (N_4676,N_4449,N_4295);
or U4677 (N_4677,N_4398,N_4294);
and U4678 (N_4678,N_4308,N_4283);
nand U4679 (N_4679,N_4267,N_4481);
and U4680 (N_4680,N_4265,N_4351);
nand U4681 (N_4681,N_4483,N_4346);
and U4682 (N_4682,N_4323,N_4426);
or U4683 (N_4683,N_4382,N_4468);
or U4684 (N_4684,N_4304,N_4407);
nor U4685 (N_4685,N_4474,N_4359);
or U4686 (N_4686,N_4367,N_4452);
and U4687 (N_4687,N_4332,N_4454);
xor U4688 (N_4688,N_4377,N_4323);
or U4689 (N_4689,N_4280,N_4456);
and U4690 (N_4690,N_4378,N_4347);
and U4691 (N_4691,N_4420,N_4379);
or U4692 (N_4692,N_4312,N_4325);
and U4693 (N_4693,N_4495,N_4487);
nand U4694 (N_4694,N_4281,N_4367);
xnor U4695 (N_4695,N_4489,N_4363);
or U4696 (N_4696,N_4368,N_4283);
and U4697 (N_4697,N_4344,N_4452);
or U4698 (N_4698,N_4342,N_4372);
and U4699 (N_4699,N_4312,N_4408);
or U4700 (N_4700,N_4432,N_4464);
xnor U4701 (N_4701,N_4416,N_4478);
nor U4702 (N_4702,N_4296,N_4484);
and U4703 (N_4703,N_4463,N_4379);
and U4704 (N_4704,N_4399,N_4360);
and U4705 (N_4705,N_4344,N_4328);
and U4706 (N_4706,N_4282,N_4494);
and U4707 (N_4707,N_4269,N_4374);
nand U4708 (N_4708,N_4343,N_4312);
nor U4709 (N_4709,N_4302,N_4268);
nor U4710 (N_4710,N_4286,N_4352);
or U4711 (N_4711,N_4365,N_4276);
xnor U4712 (N_4712,N_4483,N_4429);
nor U4713 (N_4713,N_4388,N_4262);
nand U4714 (N_4714,N_4420,N_4438);
nor U4715 (N_4715,N_4288,N_4443);
or U4716 (N_4716,N_4444,N_4336);
nor U4717 (N_4717,N_4498,N_4415);
nand U4718 (N_4718,N_4307,N_4368);
nand U4719 (N_4719,N_4389,N_4422);
and U4720 (N_4720,N_4466,N_4426);
or U4721 (N_4721,N_4296,N_4489);
or U4722 (N_4722,N_4424,N_4260);
or U4723 (N_4723,N_4444,N_4362);
nand U4724 (N_4724,N_4413,N_4320);
or U4725 (N_4725,N_4495,N_4308);
and U4726 (N_4726,N_4312,N_4446);
nor U4727 (N_4727,N_4336,N_4443);
and U4728 (N_4728,N_4265,N_4270);
or U4729 (N_4729,N_4266,N_4340);
or U4730 (N_4730,N_4379,N_4272);
xor U4731 (N_4731,N_4399,N_4328);
nand U4732 (N_4732,N_4349,N_4476);
or U4733 (N_4733,N_4264,N_4343);
nand U4734 (N_4734,N_4290,N_4360);
and U4735 (N_4735,N_4405,N_4351);
nor U4736 (N_4736,N_4327,N_4461);
and U4737 (N_4737,N_4441,N_4467);
or U4738 (N_4738,N_4426,N_4252);
and U4739 (N_4739,N_4427,N_4377);
and U4740 (N_4740,N_4294,N_4386);
nor U4741 (N_4741,N_4332,N_4268);
xnor U4742 (N_4742,N_4414,N_4275);
nand U4743 (N_4743,N_4277,N_4250);
nor U4744 (N_4744,N_4331,N_4447);
nand U4745 (N_4745,N_4297,N_4432);
and U4746 (N_4746,N_4395,N_4345);
nor U4747 (N_4747,N_4481,N_4463);
nor U4748 (N_4748,N_4255,N_4286);
xor U4749 (N_4749,N_4335,N_4251);
and U4750 (N_4750,N_4707,N_4529);
nor U4751 (N_4751,N_4598,N_4585);
nor U4752 (N_4752,N_4721,N_4611);
or U4753 (N_4753,N_4570,N_4663);
and U4754 (N_4754,N_4723,N_4531);
nand U4755 (N_4755,N_4580,N_4504);
nor U4756 (N_4756,N_4674,N_4587);
nand U4757 (N_4757,N_4632,N_4558);
nand U4758 (N_4758,N_4676,N_4704);
and U4759 (N_4759,N_4745,N_4718);
and U4760 (N_4760,N_4739,N_4625);
and U4761 (N_4761,N_4686,N_4618);
xnor U4762 (N_4762,N_4574,N_4560);
and U4763 (N_4763,N_4639,N_4727);
and U4764 (N_4764,N_4719,N_4628);
nand U4765 (N_4765,N_4641,N_4657);
nand U4766 (N_4766,N_4502,N_4582);
and U4767 (N_4767,N_4536,N_4682);
xor U4768 (N_4768,N_4732,N_4593);
nor U4769 (N_4769,N_4517,N_4678);
nor U4770 (N_4770,N_4552,N_4594);
nor U4771 (N_4771,N_4722,N_4622);
or U4772 (N_4772,N_4522,N_4629);
nor U4773 (N_4773,N_4556,N_4533);
or U4774 (N_4774,N_4561,N_4519);
nor U4775 (N_4775,N_4726,N_4636);
nand U4776 (N_4776,N_4528,N_4656);
nor U4777 (N_4777,N_4684,N_4566);
and U4778 (N_4778,N_4717,N_4691);
nor U4779 (N_4779,N_4644,N_4661);
nand U4780 (N_4780,N_4701,N_4665);
nor U4781 (N_4781,N_4526,N_4518);
nor U4782 (N_4782,N_4507,N_4700);
and U4783 (N_4783,N_4550,N_4591);
nand U4784 (N_4784,N_4520,N_4709);
nand U4785 (N_4785,N_4606,N_4554);
nor U4786 (N_4786,N_4597,N_4545);
xnor U4787 (N_4787,N_4649,N_4596);
or U4788 (N_4788,N_4735,N_4694);
or U4789 (N_4789,N_4509,N_4546);
or U4790 (N_4790,N_4549,N_4690);
and U4791 (N_4791,N_4681,N_4605);
and U4792 (N_4792,N_4720,N_4600);
nand U4793 (N_4793,N_4680,N_4563);
xor U4794 (N_4794,N_4608,N_4713);
nand U4795 (N_4795,N_4512,N_4671);
nand U4796 (N_4796,N_4621,N_4541);
or U4797 (N_4797,N_4592,N_4508);
nor U4798 (N_4798,N_4642,N_4643);
nor U4799 (N_4799,N_4573,N_4568);
or U4800 (N_4800,N_4724,N_4711);
and U4801 (N_4801,N_4620,N_4510);
nor U4802 (N_4802,N_4640,N_4693);
or U4803 (N_4803,N_4633,N_4532);
nand U4804 (N_4804,N_4503,N_4583);
nand U4805 (N_4805,N_4679,N_4734);
nand U4806 (N_4806,N_4740,N_4715);
or U4807 (N_4807,N_4523,N_4653);
nand U4808 (N_4808,N_4699,N_4505);
and U4809 (N_4809,N_4527,N_4516);
and U4810 (N_4810,N_4637,N_4544);
and U4811 (N_4811,N_4685,N_4728);
nand U4812 (N_4812,N_4652,N_4572);
nor U4813 (N_4813,N_4645,N_4589);
or U4814 (N_4814,N_4630,N_4500);
nor U4815 (N_4815,N_4648,N_4683);
nor U4816 (N_4816,N_4737,N_4654);
nand U4817 (N_4817,N_4571,N_4710);
or U4818 (N_4818,N_4537,N_4581);
or U4819 (N_4819,N_4506,N_4603);
and U4820 (N_4820,N_4631,N_4595);
nor U4821 (N_4821,N_4524,N_4667);
xnor U4822 (N_4822,N_4655,N_4702);
or U4823 (N_4823,N_4543,N_4624);
or U4824 (N_4824,N_4731,N_4747);
and U4825 (N_4825,N_4538,N_4736);
and U4826 (N_4826,N_4688,N_4738);
and U4827 (N_4827,N_4542,N_4578);
or U4828 (N_4828,N_4647,N_4539);
and U4829 (N_4829,N_4623,N_4730);
or U4830 (N_4830,N_4540,N_4689);
nand U4831 (N_4831,N_4599,N_4646);
nand U4832 (N_4832,N_4610,N_4616);
nor U4833 (N_4833,N_4562,N_4659);
nor U4834 (N_4834,N_4501,N_4627);
or U4835 (N_4835,N_4565,N_4743);
and U4836 (N_4836,N_4551,N_4634);
or U4837 (N_4837,N_4607,N_4521);
nor U4838 (N_4838,N_4725,N_4687);
nor U4839 (N_4839,N_4609,N_4564);
nand U4840 (N_4840,N_4706,N_4741);
xnor U4841 (N_4841,N_4660,N_4513);
nor U4842 (N_4842,N_4677,N_4601);
nand U4843 (N_4843,N_4666,N_4530);
or U4844 (N_4844,N_4658,N_4712);
nand U4845 (N_4845,N_4588,N_4692);
xor U4846 (N_4846,N_4547,N_4744);
and U4847 (N_4847,N_4515,N_4626);
and U4848 (N_4848,N_4708,N_4698);
and U4849 (N_4849,N_4619,N_4703);
nor U4850 (N_4850,N_4559,N_4534);
nor U4851 (N_4851,N_4638,N_4567);
xnor U4852 (N_4852,N_4670,N_4672);
nor U4853 (N_4853,N_4548,N_4749);
nor U4854 (N_4854,N_4695,N_4602);
or U4855 (N_4855,N_4664,N_4576);
and U4856 (N_4856,N_4635,N_4586);
nand U4857 (N_4857,N_4733,N_4662);
or U4858 (N_4858,N_4579,N_4729);
nand U4859 (N_4859,N_4590,N_4746);
and U4860 (N_4860,N_4748,N_4650);
xor U4861 (N_4861,N_4511,N_4705);
and U4862 (N_4862,N_4604,N_4553);
and U4863 (N_4863,N_4535,N_4696);
or U4864 (N_4864,N_4613,N_4669);
and U4865 (N_4865,N_4714,N_4577);
nand U4866 (N_4866,N_4557,N_4716);
nand U4867 (N_4867,N_4612,N_4668);
nand U4868 (N_4868,N_4614,N_4569);
or U4869 (N_4869,N_4525,N_4514);
nor U4870 (N_4870,N_4651,N_4673);
nor U4871 (N_4871,N_4742,N_4615);
or U4872 (N_4872,N_4575,N_4555);
nor U4873 (N_4873,N_4675,N_4617);
nor U4874 (N_4874,N_4584,N_4697);
nand U4875 (N_4875,N_4576,N_4699);
xnor U4876 (N_4876,N_4514,N_4706);
and U4877 (N_4877,N_4616,N_4528);
nor U4878 (N_4878,N_4555,N_4727);
nor U4879 (N_4879,N_4534,N_4545);
or U4880 (N_4880,N_4589,N_4658);
nand U4881 (N_4881,N_4711,N_4735);
or U4882 (N_4882,N_4567,N_4502);
nor U4883 (N_4883,N_4726,N_4715);
or U4884 (N_4884,N_4509,N_4611);
and U4885 (N_4885,N_4742,N_4542);
nand U4886 (N_4886,N_4526,N_4646);
and U4887 (N_4887,N_4535,N_4500);
nor U4888 (N_4888,N_4685,N_4618);
xor U4889 (N_4889,N_4703,N_4549);
nor U4890 (N_4890,N_4574,N_4573);
nor U4891 (N_4891,N_4536,N_4500);
xnor U4892 (N_4892,N_4737,N_4692);
nand U4893 (N_4893,N_4727,N_4695);
nor U4894 (N_4894,N_4527,N_4663);
or U4895 (N_4895,N_4535,N_4550);
nand U4896 (N_4896,N_4551,N_4663);
and U4897 (N_4897,N_4601,N_4629);
and U4898 (N_4898,N_4721,N_4561);
or U4899 (N_4899,N_4730,N_4588);
nor U4900 (N_4900,N_4741,N_4632);
nor U4901 (N_4901,N_4718,N_4627);
or U4902 (N_4902,N_4610,N_4641);
xnor U4903 (N_4903,N_4500,N_4588);
nor U4904 (N_4904,N_4569,N_4518);
nand U4905 (N_4905,N_4539,N_4631);
and U4906 (N_4906,N_4699,N_4566);
and U4907 (N_4907,N_4596,N_4553);
nor U4908 (N_4908,N_4550,N_4720);
or U4909 (N_4909,N_4580,N_4679);
nor U4910 (N_4910,N_4732,N_4690);
xnor U4911 (N_4911,N_4734,N_4656);
and U4912 (N_4912,N_4598,N_4700);
xnor U4913 (N_4913,N_4746,N_4619);
or U4914 (N_4914,N_4512,N_4641);
or U4915 (N_4915,N_4514,N_4618);
nor U4916 (N_4916,N_4666,N_4667);
and U4917 (N_4917,N_4704,N_4544);
or U4918 (N_4918,N_4710,N_4723);
and U4919 (N_4919,N_4635,N_4695);
and U4920 (N_4920,N_4707,N_4537);
nor U4921 (N_4921,N_4587,N_4545);
nor U4922 (N_4922,N_4549,N_4569);
or U4923 (N_4923,N_4630,N_4613);
and U4924 (N_4924,N_4708,N_4618);
xor U4925 (N_4925,N_4707,N_4594);
or U4926 (N_4926,N_4574,N_4654);
or U4927 (N_4927,N_4694,N_4592);
and U4928 (N_4928,N_4598,N_4540);
nand U4929 (N_4929,N_4715,N_4680);
and U4930 (N_4930,N_4501,N_4747);
nor U4931 (N_4931,N_4723,N_4737);
xnor U4932 (N_4932,N_4647,N_4653);
and U4933 (N_4933,N_4706,N_4565);
nor U4934 (N_4934,N_4666,N_4626);
nor U4935 (N_4935,N_4509,N_4503);
or U4936 (N_4936,N_4682,N_4685);
nand U4937 (N_4937,N_4605,N_4613);
or U4938 (N_4938,N_4749,N_4547);
or U4939 (N_4939,N_4593,N_4723);
nor U4940 (N_4940,N_4630,N_4533);
or U4941 (N_4941,N_4622,N_4565);
and U4942 (N_4942,N_4636,N_4535);
nand U4943 (N_4943,N_4579,N_4683);
nor U4944 (N_4944,N_4666,N_4523);
or U4945 (N_4945,N_4681,N_4660);
nor U4946 (N_4946,N_4558,N_4670);
or U4947 (N_4947,N_4522,N_4679);
or U4948 (N_4948,N_4594,N_4628);
nor U4949 (N_4949,N_4573,N_4602);
xnor U4950 (N_4950,N_4711,N_4512);
nand U4951 (N_4951,N_4607,N_4675);
or U4952 (N_4952,N_4558,N_4507);
nand U4953 (N_4953,N_4737,N_4531);
xnor U4954 (N_4954,N_4601,N_4581);
nand U4955 (N_4955,N_4719,N_4709);
and U4956 (N_4956,N_4724,N_4540);
xnor U4957 (N_4957,N_4747,N_4626);
and U4958 (N_4958,N_4703,N_4732);
and U4959 (N_4959,N_4522,N_4690);
nand U4960 (N_4960,N_4623,N_4557);
or U4961 (N_4961,N_4701,N_4517);
nand U4962 (N_4962,N_4604,N_4717);
nand U4963 (N_4963,N_4681,N_4569);
nand U4964 (N_4964,N_4513,N_4591);
nand U4965 (N_4965,N_4673,N_4585);
or U4966 (N_4966,N_4501,N_4517);
or U4967 (N_4967,N_4675,N_4572);
or U4968 (N_4968,N_4554,N_4648);
and U4969 (N_4969,N_4646,N_4514);
and U4970 (N_4970,N_4691,N_4592);
nand U4971 (N_4971,N_4603,N_4690);
nor U4972 (N_4972,N_4708,N_4673);
and U4973 (N_4973,N_4630,N_4708);
nor U4974 (N_4974,N_4639,N_4666);
and U4975 (N_4975,N_4625,N_4733);
nor U4976 (N_4976,N_4530,N_4590);
and U4977 (N_4977,N_4500,N_4703);
and U4978 (N_4978,N_4627,N_4533);
and U4979 (N_4979,N_4500,N_4746);
xnor U4980 (N_4980,N_4520,N_4596);
or U4981 (N_4981,N_4505,N_4723);
xnor U4982 (N_4982,N_4505,N_4524);
or U4983 (N_4983,N_4601,N_4583);
nor U4984 (N_4984,N_4620,N_4718);
xnor U4985 (N_4985,N_4668,N_4596);
or U4986 (N_4986,N_4596,N_4692);
nor U4987 (N_4987,N_4541,N_4746);
nor U4988 (N_4988,N_4729,N_4707);
and U4989 (N_4989,N_4542,N_4719);
or U4990 (N_4990,N_4556,N_4616);
or U4991 (N_4991,N_4666,N_4728);
or U4992 (N_4992,N_4669,N_4648);
nor U4993 (N_4993,N_4615,N_4530);
nand U4994 (N_4994,N_4672,N_4704);
xnor U4995 (N_4995,N_4733,N_4554);
nand U4996 (N_4996,N_4568,N_4620);
nand U4997 (N_4997,N_4746,N_4630);
nor U4998 (N_4998,N_4548,N_4743);
and U4999 (N_4999,N_4640,N_4690);
or U5000 (N_5000,N_4995,N_4991);
nand U5001 (N_5001,N_4824,N_4889);
nor U5002 (N_5002,N_4882,N_4777);
and U5003 (N_5003,N_4838,N_4771);
and U5004 (N_5004,N_4922,N_4778);
and U5005 (N_5005,N_4796,N_4880);
nand U5006 (N_5006,N_4957,N_4927);
nand U5007 (N_5007,N_4809,N_4794);
or U5008 (N_5008,N_4986,N_4805);
xor U5009 (N_5009,N_4930,N_4960);
and U5010 (N_5010,N_4770,N_4863);
nand U5011 (N_5011,N_4842,N_4821);
and U5012 (N_5012,N_4786,N_4984);
nand U5013 (N_5013,N_4994,N_4812);
nand U5014 (N_5014,N_4755,N_4964);
nand U5015 (N_5015,N_4885,N_4774);
or U5016 (N_5016,N_4907,N_4945);
and U5017 (N_5017,N_4846,N_4855);
xor U5018 (N_5018,N_4856,N_4938);
xnor U5019 (N_5019,N_4905,N_4868);
or U5020 (N_5020,N_4993,N_4811);
xor U5021 (N_5021,N_4802,N_4963);
and U5022 (N_5022,N_4823,N_4955);
nor U5023 (N_5023,N_4997,N_4941);
or U5024 (N_5024,N_4841,N_4954);
and U5025 (N_5025,N_4881,N_4756);
nor U5026 (N_5026,N_4886,N_4869);
nand U5027 (N_5027,N_4990,N_4827);
and U5028 (N_5028,N_4894,N_4864);
and U5029 (N_5029,N_4888,N_4897);
nand U5030 (N_5030,N_4830,N_4813);
or U5031 (N_5031,N_4903,N_4866);
xnor U5032 (N_5032,N_4834,N_4998);
nand U5033 (N_5033,N_4877,N_4949);
nor U5034 (N_5034,N_4883,N_4873);
nor U5035 (N_5035,N_4839,N_4792);
nor U5036 (N_5036,N_4942,N_4752);
nand U5037 (N_5037,N_4845,N_4865);
xor U5038 (N_5038,N_4988,N_4766);
and U5039 (N_5039,N_4789,N_4790);
or U5040 (N_5040,N_4832,N_4853);
nand U5041 (N_5041,N_4909,N_4931);
nand U5042 (N_5042,N_4914,N_4912);
and U5043 (N_5043,N_4773,N_4843);
nor U5044 (N_5044,N_4765,N_4944);
nor U5045 (N_5045,N_4937,N_4852);
nand U5046 (N_5046,N_4982,N_4936);
xor U5047 (N_5047,N_4753,N_4916);
nand U5048 (N_5048,N_4776,N_4918);
and U5049 (N_5049,N_4782,N_4861);
nand U5050 (N_5050,N_4919,N_4879);
nor U5051 (N_5051,N_4913,N_4962);
nor U5052 (N_5052,N_4763,N_4822);
or U5053 (N_5053,N_4965,N_4850);
or U5054 (N_5054,N_4884,N_4859);
nor U5055 (N_5055,N_4992,N_4785);
xnor U5056 (N_5056,N_4972,N_4761);
nand U5057 (N_5057,N_4840,N_4780);
and U5058 (N_5058,N_4906,N_4910);
and U5059 (N_5059,N_4779,N_4967);
nor U5060 (N_5060,N_4947,N_4784);
and U5061 (N_5061,N_4872,N_4951);
or U5062 (N_5062,N_4799,N_4975);
or U5063 (N_5063,N_4767,N_4871);
nand U5064 (N_5064,N_4925,N_4801);
and U5065 (N_5065,N_4898,N_4961);
xnor U5066 (N_5066,N_4870,N_4769);
nand U5067 (N_5067,N_4791,N_4929);
and U5068 (N_5068,N_4849,N_4973);
nor U5069 (N_5069,N_4754,N_4950);
nand U5070 (N_5070,N_4847,N_4795);
and U5071 (N_5071,N_4900,N_4875);
nor U5072 (N_5072,N_4893,N_4924);
nor U5073 (N_5073,N_4904,N_4862);
nand U5074 (N_5074,N_4958,N_4974);
nor U5075 (N_5075,N_4835,N_4921);
or U5076 (N_5076,N_4768,N_4851);
nor U5077 (N_5077,N_4971,N_4977);
nor U5078 (N_5078,N_4876,N_4858);
and U5079 (N_5079,N_4939,N_4783);
or U5080 (N_5080,N_4760,N_4978);
or U5081 (N_5081,N_4902,N_4987);
xnor U5082 (N_5082,N_4887,N_4814);
and U5083 (N_5083,N_4908,N_4933);
nand U5084 (N_5084,N_4917,N_4979);
xor U5085 (N_5085,N_4969,N_4999);
nand U5086 (N_5086,N_4788,N_4829);
nor U5087 (N_5087,N_4837,N_4816);
or U5088 (N_5088,N_4890,N_4985);
and U5089 (N_5089,N_4940,N_4848);
nor U5090 (N_5090,N_4874,N_4983);
xor U5091 (N_5091,N_4935,N_4759);
nand U5092 (N_5092,N_4828,N_4926);
xor U5093 (N_5093,N_4833,N_4920);
nand U5094 (N_5094,N_4826,N_4797);
nor U5095 (N_5095,N_4803,N_4923);
nor U5096 (N_5096,N_4952,N_4758);
nor U5097 (N_5097,N_4932,N_4867);
and U5098 (N_5098,N_4787,N_4892);
xor U5099 (N_5099,N_4793,N_4953);
and U5100 (N_5100,N_4895,N_4934);
and U5101 (N_5101,N_4825,N_4775);
nand U5102 (N_5102,N_4831,N_4891);
and U5103 (N_5103,N_4857,N_4948);
nand U5104 (N_5104,N_4996,N_4807);
and U5105 (N_5105,N_4901,N_4970);
or U5106 (N_5106,N_4878,N_4817);
nand U5107 (N_5107,N_4946,N_4810);
nor U5108 (N_5108,N_4844,N_4751);
and U5109 (N_5109,N_4854,N_4764);
and U5110 (N_5110,N_4968,N_4899);
nand U5111 (N_5111,N_4989,N_4750);
and U5112 (N_5112,N_4928,N_4896);
nor U5113 (N_5113,N_4836,N_4808);
nor U5114 (N_5114,N_4911,N_4762);
and U5115 (N_5115,N_4800,N_4966);
nand U5116 (N_5116,N_4772,N_4981);
nor U5117 (N_5117,N_4860,N_4806);
or U5118 (N_5118,N_4820,N_4915);
nand U5119 (N_5119,N_4815,N_4959);
or U5120 (N_5120,N_4781,N_4757);
or U5121 (N_5121,N_4976,N_4943);
or U5122 (N_5122,N_4980,N_4956);
or U5123 (N_5123,N_4819,N_4804);
nand U5124 (N_5124,N_4798,N_4818);
nand U5125 (N_5125,N_4984,N_4949);
and U5126 (N_5126,N_4923,N_4842);
nand U5127 (N_5127,N_4784,N_4765);
nor U5128 (N_5128,N_4891,N_4788);
nor U5129 (N_5129,N_4918,N_4750);
nor U5130 (N_5130,N_4954,N_4870);
nand U5131 (N_5131,N_4887,N_4753);
and U5132 (N_5132,N_4784,N_4887);
or U5133 (N_5133,N_4862,N_4900);
or U5134 (N_5134,N_4911,N_4909);
nor U5135 (N_5135,N_4773,N_4872);
or U5136 (N_5136,N_4780,N_4910);
nor U5137 (N_5137,N_4921,N_4984);
and U5138 (N_5138,N_4829,N_4985);
or U5139 (N_5139,N_4842,N_4775);
or U5140 (N_5140,N_4847,N_4831);
or U5141 (N_5141,N_4801,N_4781);
nor U5142 (N_5142,N_4883,N_4967);
or U5143 (N_5143,N_4855,N_4775);
nand U5144 (N_5144,N_4767,N_4890);
or U5145 (N_5145,N_4765,N_4834);
nor U5146 (N_5146,N_4780,N_4909);
nor U5147 (N_5147,N_4801,N_4993);
nor U5148 (N_5148,N_4986,N_4985);
nor U5149 (N_5149,N_4995,N_4888);
nor U5150 (N_5150,N_4983,N_4789);
and U5151 (N_5151,N_4802,N_4978);
and U5152 (N_5152,N_4932,N_4759);
or U5153 (N_5153,N_4984,N_4787);
nand U5154 (N_5154,N_4979,N_4861);
nand U5155 (N_5155,N_4932,N_4972);
and U5156 (N_5156,N_4875,N_4755);
nor U5157 (N_5157,N_4826,N_4805);
and U5158 (N_5158,N_4952,N_4909);
or U5159 (N_5159,N_4914,N_4976);
xor U5160 (N_5160,N_4962,N_4904);
nand U5161 (N_5161,N_4992,N_4867);
and U5162 (N_5162,N_4861,N_4912);
nand U5163 (N_5163,N_4925,N_4879);
nand U5164 (N_5164,N_4796,N_4920);
nand U5165 (N_5165,N_4851,N_4836);
nor U5166 (N_5166,N_4813,N_4865);
or U5167 (N_5167,N_4828,N_4865);
or U5168 (N_5168,N_4913,N_4792);
or U5169 (N_5169,N_4896,N_4789);
nor U5170 (N_5170,N_4957,N_4829);
or U5171 (N_5171,N_4762,N_4837);
nand U5172 (N_5172,N_4880,N_4974);
and U5173 (N_5173,N_4793,N_4782);
nand U5174 (N_5174,N_4993,N_4855);
nand U5175 (N_5175,N_4900,N_4922);
and U5176 (N_5176,N_4780,N_4834);
nor U5177 (N_5177,N_4948,N_4898);
xnor U5178 (N_5178,N_4770,N_4885);
nand U5179 (N_5179,N_4811,N_4788);
or U5180 (N_5180,N_4887,N_4828);
and U5181 (N_5181,N_4969,N_4759);
and U5182 (N_5182,N_4928,N_4825);
or U5183 (N_5183,N_4928,N_4841);
nand U5184 (N_5184,N_4923,N_4962);
xor U5185 (N_5185,N_4835,N_4916);
or U5186 (N_5186,N_4791,N_4973);
nor U5187 (N_5187,N_4877,N_4904);
and U5188 (N_5188,N_4848,N_4957);
or U5189 (N_5189,N_4827,N_4924);
nor U5190 (N_5190,N_4849,N_4865);
and U5191 (N_5191,N_4881,N_4755);
and U5192 (N_5192,N_4993,N_4934);
xnor U5193 (N_5193,N_4985,N_4895);
nand U5194 (N_5194,N_4998,N_4873);
and U5195 (N_5195,N_4923,N_4993);
or U5196 (N_5196,N_4799,N_4925);
nor U5197 (N_5197,N_4823,N_4788);
nor U5198 (N_5198,N_4901,N_4914);
and U5199 (N_5199,N_4929,N_4956);
or U5200 (N_5200,N_4923,N_4858);
or U5201 (N_5201,N_4753,N_4934);
or U5202 (N_5202,N_4944,N_4810);
or U5203 (N_5203,N_4860,N_4787);
nand U5204 (N_5204,N_4974,N_4806);
or U5205 (N_5205,N_4918,N_4879);
nand U5206 (N_5206,N_4801,N_4949);
nor U5207 (N_5207,N_4991,N_4957);
or U5208 (N_5208,N_4781,N_4818);
nor U5209 (N_5209,N_4888,N_4931);
nor U5210 (N_5210,N_4863,N_4751);
nand U5211 (N_5211,N_4846,N_4770);
and U5212 (N_5212,N_4836,N_4801);
nand U5213 (N_5213,N_4924,N_4948);
xor U5214 (N_5214,N_4811,N_4766);
nand U5215 (N_5215,N_4805,N_4865);
nor U5216 (N_5216,N_4850,N_4854);
or U5217 (N_5217,N_4814,N_4807);
nor U5218 (N_5218,N_4972,N_4941);
nor U5219 (N_5219,N_4895,N_4954);
and U5220 (N_5220,N_4916,N_4844);
or U5221 (N_5221,N_4919,N_4951);
nor U5222 (N_5222,N_4833,N_4899);
and U5223 (N_5223,N_4815,N_4981);
nand U5224 (N_5224,N_4808,N_4754);
nor U5225 (N_5225,N_4817,N_4911);
xor U5226 (N_5226,N_4923,N_4901);
nand U5227 (N_5227,N_4990,N_4938);
xnor U5228 (N_5228,N_4982,N_4866);
nor U5229 (N_5229,N_4797,N_4852);
and U5230 (N_5230,N_4778,N_4757);
or U5231 (N_5231,N_4994,N_4889);
nand U5232 (N_5232,N_4818,N_4869);
nor U5233 (N_5233,N_4961,N_4960);
nor U5234 (N_5234,N_4805,N_4761);
and U5235 (N_5235,N_4862,N_4760);
xnor U5236 (N_5236,N_4901,N_4830);
nor U5237 (N_5237,N_4810,N_4979);
and U5238 (N_5238,N_4816,N_4948);
nor U5239 (N_5239,N_4773,N_4936);
or U5240 (N_5240,N_4846,N_4985);
or U5241 (N_5241,N_4805,N_4755);
and U5242 (N_5242,N_4842,N_4879);
or U5243 (N_5243,N_4854,N_4986);
nor U5244 (N_5244,N_4922,N_4893);
and U5245 (N_5245,N_4879,N_4754);
nor U5246 (N_5246,N_4936,N_4780);
and U5247 (N_5247,N_4825,N_4751);
nand U5248 (N_5248,N_4954,N_4848);
nor U5249 (N_5249,N_4758,N_4751);
nor U5250 (N_5250,N_5031,N_5146);
or U5251 (N_5251,N_5021,N_5237);
or U5252 (N_5252,N_5168,N_5193);
and U5253 (N_5253,N_5184,N_5171);
or U5254 (N_5254,N_5159,N_5017);
and U5255 (N_5255,N_5071,N_5186);
nor U5256 (N_5256,N_5144,N_5213);
and U5257 (N_5257,N_5209,N_5054);
nand U5258 (N_5258,N_5156,N_5037);
and U5259 (N_5259,N_5056,N_5117);
or U5260 (N_5260,N_5133,N_5124);
nand U5261 (N_5261,N_5103,N_5226);
and U5262 (N_5262,N_5162,N_5099);
nor U5263 (N_5263,N_5132,N_5008);
or U5264 (N_5264,N_5069,N_5070);
nor U5265 (N_5265,N_5010,N_5085);
nor U5266 (N_5266,N_5195,N_5104);
nor U5267 (N_5267,N_5157,N_5084);
and U5268 (N_5268,N_5126,N_5147);
nor U5269 (N_5269,N_5196,N_5148);
xnor U5270 (N_5270,N_5022,N_5136);
or U5271 (N_5271,N_5172,N_5077);
nand U5272 (N_5272,N_5248,N_5067);
nor U5273 (N_5273,N_5178,N_5044);
and U5274 (N_5274,N_5115,N_5138);
nand U5275 (N_5275,N_5075,N_5055);
or U5276 (N_5276,N_5145,N_5102);
nand U5277 (N_5277,N_5151,N_5236);
nor U5278 (N_5278,N_5016,N_5107);
nor U5279 (N_5279,N_5210,N_5176);
nand U5280 (N_5280,N_5000,N_5129);
nor U5281 (N_5281,N_5123,N_5039);
or U5282 (N_5282,N_5189,N_5116);
and U5283 (N_5283,N_5029,N_5153);
xnor U5284 (N_5284,N_5066,N_5224);
nor U5285 (N_5285,N_5142,N_5072);
nand U5286 (N_5286,N_5087,N_5205);
xnor U5287 (N_5287,N_5166,N_5112);
nand U5288 (N_5288,N_5105,N_5165);
nor U5289 (N_5289,N_5191,N_5231);
nor U5290 (N_5290,N_5011,N_5245);
nor U5291 (N_5291,N_5026,N_5064);
nor U5292 (N_5292,N_5217,N_5177);
and U5293 (N_5293,N_5113,N_5180);
nand U5294 (N_5294,N_5238,N_5023);
nor U5295 (N_5295,N_5201,N_5110);
and U5296 (N_5296,N_5033,N_5076);
or U5297 (N_5297,N_5208,N_5154);
xnor U5298 (N_5298,N_5218,N_5198);
nor U5299 (N_5299,N_5019,N_5025);
nor U5300 (N_5300,N_5013,N_5060);
nor U5301 (N_5301,N_5216,N_5139);
nor U5302 (N_5302,N_5083,N_5163);
nand U5303 (N_5303,N_5135,N_5249);
nand U5304 (N_5304,N_5074,N_5122);
nand U5305 (N_5305,N_5212,N_5015);
xnor U5306 (N_5306,N_5080,N_5003);
nor U5307 (N_5307,N_5004,N_5247);
nor U5308 (N_5308,N_5188,N_5053);
nand U5309 (N_5309,N_5170,N_5152);
and U5310 (N_5310,N_5227,N_5040);
and U5311 (N_5311,N_5230,N_5190);
xnor U5312 (N_5312,N_5091,N_5079);
and U5313 (N_5313,N_5052,N_5078);
or U5314 (N_5314,N_5062,N_5141);
and U5315 (N_5315,N_5118,N_5240);
nor U5316 (N_5316,N_5158,N_5223);
and U5317 (N_5317,N_5203,N_5035);
or U5318 (N_5318,N_5014,N_5174);
xor U5319 (N_5319,N_5081,N_5073);
and U5320 (N_5320,N_5187,N_5120);
xnor U5321 (N_5321,N_5086,N_5179);
or U5322 (N_5322,N_5088,N_5125);
nor U5323 (N_5323,N_5106,N_5030);
nor U5324 (N_5324,N_5009,N_5090);
and U5325 (N_5325,N_5194,N_5127);
and U5326 (N_5326,N_5137,N_5095);
nor U5327 (N_5327,N_5233,N_5235);
nand U5328 (N_5328,N_5169,N_5092);
nor U5329 (N_5329,N_5097,N_5128);
xnor U5330 (N_5330,N_5134,N_5045);
and U5331 (N_5331,N_5059,N_5038);
nand U5332 (N_5332,N_5057,N_5131);
or U5333 (N_5333,N_5228,N_5093);
nand U5334 (N_5334,N_5049,N_5161);
or U5335 (N_5335,N_5024,N_5200);
and U5336 (N_5336,N_5063,N_5155);
or U5337 (N_5337,N_5047,N_5058);
nor U5338 (N_5338,N_5130,N_5041);
nor U5339 (N_5339,N_5220,N_5051);
or U5340 (N_5340,N_5150,N_5160);
and U5341 (N_5341,N_5175,N_5219);
nor U5342 (N_5342,N_5046,N_5101);
nand U5343 (N_5343,N_5012,N_5202);
nand U5344 (N_5344,N_5143,N_5002);
xnor U5345 (N_5345,N_5239,N_5246);
or U5346 (N_5346,N_5032,N_5244);
and U5347 (N_5347,N_5183,N_5225);
or U5348 (N_5348,N_5204,N_5034);
and U5349 (N_5349,N_5048,N_5007);
nand U5350 (N_5350,N_5121,N_5036);
xor U5351 (N_5351,N_5082,N_5020);
nand U5352 (N_5352,N_5001,N_5111);
xor U5353 (N_5353,N_5028,N_5065);
or U5354 (N_5354,N_5042,N_5094);
xor U5355 (N_5355,N_5068,N_5109);
and U5356 (N_5356,N_5241,N_5243);
or U5357 (N_5357,N_5119,N_5096);
and U5358 (N_5358,N_5098,N_5050);
and U5359 (N_5359,N_5061,N_5234);
xor U5360 (N_5360,N_5114,N_5181);
or U5361 (N_5361,N_5182,N_5018);
or U5362 (N_5362,N_5100,N_5199);
xor U5363 (N_5363,N_5167,N_5089);
nor U5364 (N_5364,N_5206,N_5221);
nor U5365 (N_5365,N_5222,N_5149);
and U5366 (N_5366,N_5173,N_5108);
nor U5367 (N_5367,N_5211,N_5214);
nand U5368 (N_5368,N_5197,N_5006);
or U5369 (N_5369,N_5215,N_5043);
nand U5370 (N_5370,N_5164,N_5229);
nand U5371 (N_5371,N_5185,N_5232);
and U5372 (N_5372,N_5005,N_5027);
or U5373 (N_5373,N_5207,N_5242);
or U5374 (N_5374,N_5140,N_5192);
nand U5375 (N_5375,N_5216,N_5132);
and U5376 (N_5376,N_5234,N_5132);
xnor U5377 (N_5377,N_5064,N_5022);
xnor U5378 (N_5378,N_5099,N_5174);
xor U5379 (N_5379,N_5022,N_5026);
nand U5380 (N_5380,N_5058,N_5045);
and U5381 (N_5381,N_5209,N_5117);
and U5382 (N_5382,N_5232,N_5223);
nand U5383 (N_5383,N_5008,N_5089);
nor U5384 (N_5384,N_5216,N_5078);
nor U5385 (N_5385,N_5102,N_5128);
nand U5386 (N_5386,N_5047,N_5231);
nor U5387 (N_5387,N_5208,N_5197);
nand U5388 (N_5388,N_5247,N_5134);
nand U5389 (N_5389,N_5200,N_5102);
nor U5390 (N_5390,N_5061,N_5131);
xnor U5391 (N_5391,N_5079,N_5089);
nand U5392 (N_5392,N_5116,N_5143);
xor U5393 (N_5393,N_5104,N_5084);
and U5394 (N_5394,N_5140,N_5126);
or U5395 (N_5395,N_5137,N_5103);
nand U5396 (N_5396,N_5075,N_5235);
nand U5397 (N_5397,N_5179,N_5033);
nor U5398 (N_5398,N_5162,N_5156);
and U5399 (N_5399,N_5021,N_5034);
or U5400 (N_5400,N_5095,N_5071);
xor U5401 (N_5401,N_5135,N_5081);
and U5402 (N_5402,N_5145,N_5081);
nor U5403 (N_5403,N_5025,N_5191);
nand U5404 (N_5404,N_5135,N_5086);
or U5405 (N_5405,N_5194,N_5161);
or U5406 (N_5406,N_5232,N_5168);
or U5407 (N_5407,N_5205,N_5164);
nor U5408 (N_5408,N_5245,N_5094);
nor U5409 (N_5409,N_5001,N_5242);
or U5410 (N_5410,N_5150,N_5032);
or U5411 (N_5411,N_5054,N_5088);
nor U5412 (N_5412,N_5201,N_5240);
or U5413 (N_5413,N_5243,N_5092);
and U5414 (N_5414,N_5030,N_5068);
nor U5415 (N_5415,N_5218,N_5119);
and U5416 (N_5416,N_5040,N_5064);
nor U5417 (N_5417,N_5035,N_5146);
nand U5418 (N_5418,N_5227,N_5001);
or U5419 (N_5419,N_5080,N_5050);
or U5420 (N_5420,N_5039,N_5070);
and U5421 (N_5421,N_5032,N_5151);
nand U5422 (N_5422,N_5075,N_5001);
nand U5423 (N_5423,N_5141,N_5205);
xor U5424 (N_5424,N_5188,N_5076);
or U5425 (N_5425,N_5087,N_5108);
or U5426 (N_5426,N_5235,N_5063);
or U5427 (N_5427,N_5225,N_5201);
or U5428 (N_5428,N_5124,N_5246);
and U5429 (N_5429,N_5064,N_5112);
or U5430 (N_5430,N_5225,N_5159);
and U5431 (N_5431,N_5228,N_5160);
and U5432 (N_5432,N_5058,N_5056);
xnor U5433 (N_5433,N_5058,N_5012);
nand U5434 (N_5434,N_5040,N_5167);
or U5435 (N_5435,N_5186,N_5214);
and U5436 (N_5436,N_5043,N_5038);
nand U5437 (N_5437,N_5231,N_5156);
nand U5438 (N_5438,N_5172,N_5029);
nand U5439 (N_5439,N_5047,N_5121);
nor U5440 (N_5440,N_5118,N_5140);
nor U5441 (N_5441,N_5120,N_5209);
nand U5442 (N_5442,N_5231,N_5175);
nand U5443 (N_5443,N_5137,N_5074);
or U5444 (N_5444,N_5026,N_5153);
nand U5445 (N_5445,N_5007,N_5094);
nor U5446 (N_5446,N_5174,N_5126);
or U5447 (N_5447,N_5175,N_5078);
xnor U5448 (N_5448,N_5070,N_5175);
nor U5449 (N_5449,N_5082,N_5036);
or U5450 (N_5450,N_5218,N_5095);
nand U5451 (N_5451,N_5066,N_5105);
nand U5452 (N_5452,N_5062,N_5206);
xor U5453 (N_5453,N_5142,N_5109);
nor U5454 (N_5454,N_5028,N_5236);
or U5455 (N_5455,N_5137,N_5234);
or U5456 (N_5456,N_5245,N_5205);
and U5457 (N_5457,N_5218,N_5030);
and U5458 (N_5458,N_5242,N_5075);
or U5459 (N_5459,N_5146,N_5051);
nand U5460 (N_5460,N_5114,N_5017);
nor U5461 (N_5461,N_5029,N_5090);
nor U5462 (N_5462,N_5176,N_5249);
and U5463 (N_5463,N_5236,N_5233);
or U5464 (N_5464,N_5170,N_5120);
nand U5465 (N_5465,N_5036,N_5041);
nor U5466 (N_5466,N_5155,N_5031);
and U5467 (N_5467,N_5214,N_5029);
or U5468 (N_5468,N_5165,N_5055);
nand U5469 (N_5469,N_5081,N_5143);
nand U5470 (N_5470,N_5031,N_5247);
and U5471 (N_5471,N_5241,N_5188);
or U5472 (N_5472,N_5064,N_5136);
nand U5473 (N_5473,N_5222,N_5007);
or U5474 (N_5474,N_5201,N_5106);
and U5475 (N_5475,N_5084,N_5143);
and U5476 (N_5476,N_5003,N_5049);
and U5477 (N_5477,N_5117,N_5182);
nand U5478 (N_5478,N_5248,N_5074);
and U5479 (N_5479,N_5190,N_5173);
and U5480 (N_5480,N_5032,N_5187);
and U5481 (N_5481,N_5101,N_5174);
nand U5482 (N_5482,N_5210,N_5067);
nand U5483 (N_5483,N_5216,N_5242);
and U5484 (N_5484,N_5214,N_5007);
nor U5485 (N_5485,N_5199,N_5207);
nor U5486 (N_5486,N_5224,N_5215);
nand U5487 (N_5487,N_5054,N_5014);
nand U5488 (N_5488,N_5117,N_5113);
nor U5489 (N_5489,N_5142,N_5141);
and U5490 (N_5490,N_5111,N_5143);
or U5491 (N_5491,N_5123,N_5121);
xor U5492 (N_5492,N_5180,N_5175);
nand U5493 (N_5493,N_5049,N_5153);
and U5494 (N_5494,N_5210,N_5102);
nor U5495 (N_5495,N_5005,N_5015);
and U5496 (N_5496,N_5173,N_5195);
nor U5497 (N_5497,N_5049,N_5203);
nor U5498 (N_5498,N_5245,N_5012);
nor U5499 (N_5499,N_5126,N_5032);
or U5500 (N_5500,N_5445,N_5353);
nand U5501 (N_5501,N_5256,N_5391);
xor U5502 (N_5502,N_5356,N_5434);
nand U5503 (N_5503,N_5496,N_5355);
and U5504 (N_5504,N_5296,N_5429);
nand U5505 (N_5505,N_5457,N_5494);
and U5506 (N_5506,N_5367,N_5447);
nand U5507 (N_5507,N_5286,N_5425);
nand U5508 (N_5508,N_5412,N_5416);
nor U5509 (N_5509,N_5350,N_5274);
and U5510 (N_5510,N_5382,N_5323);
and U5511 (N_5511,N_5394,N_5433);
nor U5512 (N_5512,N_5285,N_5459);
xnor U5513 (N_5513,N_5450,N_5368);
and U5514 (N_5514,N_5280,N_5366);
xor U5515 (N_5515,N_5465,N_5493);
nor U5516 (N_5516,N_5390,N_5287);
nand U5517 (N_5517,N_5283,N_5384);
and U5518 (N_5518,N_5275,N_5332);
nand U5519 (N_5519,N_5329,N_5359);
nand U5520 (N_5520,N_5486,N_5320);
nor U5521 (N_5521,N_5262,N_5308);
nor U5522 (N_5522,N_5363,N_5357);
xor U5523 (N_5523,N_5378,N_5253);
nor U5524 (N_5524,N_5351,N_5341);
nand U5525 (N_5525,N_5468,N_5288);
xnor U5526 (N_5526,N_5347,N_5463);
and U5527 (N_5527,N_5354,N_5432);
or U5528 (N_5528,N_5272,N_5497);
nand U5529 (N_5529,N_5265,N_5331);
nor U5530 (N_5530,N_5271,N_5279);
nand U5531 (N_5531,N_5325,N_5362);
nand U5532 (N_5532,N_5303,N_5410);
nor U5533 (N_5533,N_5428,N_5430);
or U5534 (N_5534,N_5315,N_5392);
nor U5535 (N_5535,N_5344,N_5312);
nand U5536 (N_5536,N_5259,N_5282);
nand U5537 (N_5537,N_5388,N_5414);
and U5538 (N_5538,N_5476,N_5498);
or U5539 (N_5539,N_5495,N_5490);
and U5540 (N_5540,N_5301,N_5266);
and U5541 (N_5541,N_5387,N_5349);
and U5542 (N_5542,N_5261,N_5376);
and U5543 (N_5543,N_5369,N_5278);
or U5544 (N_5544,N_5260,N_5379);
nand U5545 (N_5545,N_5313,N_5302);
and U5546 (N_5546,N_5322,N_5334);
or U5547 (N_5547,N_5451,N_5327);
nor U5548 (N_5548,N_5257,N_5473);
and U5549 (N_5549,N_5402,N_5294);
nand U5550 (N_5550,N_5305,N_5297);
or U5551 (N_5551,N_5273,N_5328);
or U5552 (N_5552,N_5460,N_5400);
or U5553 (N_5553,N_5374,N_5335);
or U5554 (N_5554,N_5461,N_5291);
nand U5555 (N_5555,N_5491,N_5267);
nand U5556 (N_5556,N_5338,N_5485);
nor U5557 (N_5557,N_5479,N_5466);
nand U5558 (N_5558,N_5483,N_5270);
nand U5559 (N_5559,N_5406,N_5469);
nor U5560 (N_5560,N_5499,N_5333);
nor U5561 (N_5561,N_5393,N_5438);
nand U5562 (N_5562,N_5324,N_5300);
or U5563 (N_5563,N_5467,N_5321);
nand U5564 (N_5564,N_5263,N_5371);
xnor U5565 (N_5565,N_5352,N_5306);
or U5566 (N_5566,N_5255,N_5318);
nor U5567 (N_5567,N_5440,N_5441);
and U5568 (N_5568,N_5252,N_5385);
nor U5569 (N_5569,N_5277,N_5250);
or U5570 (N_5570,N_5389,N_5492);
nand U5571 (N_5571,N_5437,N_5417);
nor U5572 (N_5572,N_5456,N_5290);
xnor U5573 (N_5573,N_5442,N_5413);
and U5574 (N_5574,N_5386,N_5330);
nor U5575 (N_5575,N_5474,N_5422);
nor U5576 (N_5576,N_5427,N_5372);
or U5577 (N_5577,N_5471,N_5405);
nand U5578 (N_5578,N_5449,N_5408);
xnor U5579 (N_5579,N_5345,N_5311);
and U5580 (N_5580,N_5293,N_5480);
or U5581 (N_5581,N_5304,N_5264);
nand U5582 (N_5582,N_5299,N_5348);
and U5583 (N_5583,N_5383,N_5276);
xor U5584 (N_5584,N_5292,N_5342);
and U5585 (N_5585,N_5401,N_5375);
nand U5586 (N_5586,N_5439,N_5398);
nor U5587 (N_5587,N_5289,N_5418);
nor U5588 (N_5588,N_5488,N_5319);
xnor U5589 (N_5589,N_5444,N_5337);
nand U5590 (N_5590,N_5431,N_5436);
nand U5591 (N_5591,N_5472,N_5481);
and U5592 (N_5592,N_5396,N_5446);
or U5593 (N_5593,N_5251,N_5360);
nand U5594 (N_5594,N_5316,N_5424);
nand U5595 (N_5595,N_5370,N_5364);
or U5596 (N_5596,N_5454,N_5307);
and U5597 (N_5597,N_5380,N_5397);
nand U5598 (N_5598,N_5281,N_5309);
and U5599 (N_5599,N_5452,N_5420);
nor U5600 (N_5600,N_5298,N_5407);
xor U5601 (N_5601,N_5475,N_5373);
nand U5602 (N_5602,N_5268,N_5326);
or U5603 (N_5603,N_5395,N_5448);
nor U5604 (N_5604,N_5269,N_5423);
nor U5605 (N_5605,N_5295,N_5478);
and U5606 (N_5606,N_5415,N_5317);
nor U5607 (N_5607,N_5421,N_5487);
nor U5608 (N_5608,N_5455,N_5419);
and U5609 (N_5609,N_5409,N_5404);
and U5610 (N_5610,N_5314,N_5426);
and U5611 (N_5611,N_5343,N_5361);
nand U5612 (N_5612,N_5258,N_5484);
or U5613 (N_5613,N_5435,N_5284);
nand U5614 (N_5614,N_5381,N_5358);
nor U5615 (N_5615,N_5399,N_5458);
and U5616 (N_5616,N_5377,N_5340);
or U5617 (N_5617,N_5462,N_5470);
nor U5618 (N_5618,N_5365,N_5443);
and U5619 (N_5619,N_5346,N_5336);
nand U5620 (N_5620,N_5482,N_5254);
nor U5621 (N_5621,N_5403,N_5411);
nand U5622 (N_5622,N_5453,N_5464);
or U5623 (N_5623,N_5489,N_5477);
xor U5624 (N_5624,N_5310,N_5339);
and U5625 (N_5625,N_5422,N_5429);
xnor U5626 (N_5626,N_5412,N_5260);
nor U5627 (N_5627,N_5398,N_5368);
and U5628 (N_5628,N_5275,N_5462);
nor U5629 (N_5629,N_5294,N_5396);
xor U5630 (N_5630,N_5397,N_5288);
nor U5631 (N_5631,N_5494,N_5454);
nor U5632 (N_5632,N_5432,N_5273);
nor U5633 (N_5633,N_5397,N_5495);
or U5634 (N_5634,N_5328,N_5287);
nor U5635 (N_5635,N_5485,N_5285);
nand U5636 (N_5636,N_5385,N_5388);
nor U5637 (N_5637,N_5262,N_5418);
and U5638 (N_5638,N_5429,N_5271);
nor U5639 (N_5639,N_5463,N_5489);
xnor U5640 (N_5640,N_5452,N_5262);
and U5641 (N_5641,N_5251,N_5300);
nand U5642 (N_5642,N_5450,N_5400);
nor U5643 (N_5643,N_5316,N_5395);
or U5644 (N_5644,N_5451,N_5410);
and U5645 (N_5645,N_5355,N_5434);
nand U5646 (N_5646,N_5353,N_5390);
nor U5647 (N_5647,N_5294,N_5310);
nor U5648 (N_5648,N_5280,N_5423);
or U5649 (N_5649,N_5465,N_5468);
nor U5650 (N_5650,N_5464,N_5338);
or U5651 (N_5651,N_5363,N_5253);
nor U5652 (N_5652,N_5429,N_5311);
nand U5653 (N_5653,N_5436,N_5285);
nand U5654 (N_5654,N_5370,N_5356);
nand U5655 (N_5655,N_5316,N_5257);
and U5656 (N_5656,N_5346,N_5357);
and U5657 (N_5657,N_5278,N_5385);
or U5658 (N_5658,N_5293,N_5342);
or U5659 (N_5659,N_5338,N_5345);
nand U5660 (N_5660,N_5351,N_5458);
and U5661 (N_5661,N_5420,N_5437);
nand U5662 (N_5662,N_5270,N_5463);
and U5663 (N_5663,N_5406,N_5250);
nor U5664 (N_5664,N_5383,N_5433);
or U5665 (N_5665,N_5309,N_5360);
or U5666 (N_5666,N_5256,N_5444);
nand U5667 (N_5667,N_5474,N_5456);
and U5668 (N_5668,N_5279,N_5497);
or U5669 (N_5669,N_5486,N_5487);
nor U5670 (N_5670,N_5480,N_5425);
or U5671 (N_5671,N_5315,N_5433);
nor U5672 (N_5672,N_5472,N_5444);
and U5673 (N_5673,N_5312,N_5298);
or U5674 (N_5674,N_5349,N_5495);
nand U5675 (N_5675,N_5286,N_5268);
xor U5676 (N_5676,N_5370,N_5458);
nand U5677 (N_5677,N_5354,N_5425);
nor U5678 (N_5678,N_5370,N_5325);
and U5679 (N_5679,N_5280,N_5373);
nor U5680 (N_5680,N_5341,N_5316);
and U5681 (N_5681,N_5497,N_5414);
nor U5682 (N_5682,N_5386,N_5479);
nor U5683 (N_5683,N_5339,N_5403);
and U5684 (N_5684,N_5365,N_5487);
nand U5685 (N_5685,N_5471,N_5356);
and U5686 (N_5686,N_5445,N_5469);
xor U5687 (N_5687,N_5404,N_5320);
or U5688 (N_5688,N_5491,N_5359);
or U5689 (N_5689,N_5394,N_5498);
or U5690 (N_5690,N_5378,N_5348);
nor U5691 (N_5691,N_5470,N_5444);
nor U5692 (N_5692,N_5368,N_5383);
nand U5693 (N_5693,N_5450,N_5481);
and U5694 (N_5694,N_5442,N_5414);
or U5695 (N_5695,N_5464,N_5277);
xor U5696 (N_5696,N_5356,N_5448);
and U5697 (N_5697,N_5261,N_5375);
nor U5698 (N_5698,N_5308,N_5437);
nor U5699 (N_5699,N_5467,N_5390);
xor U5700 (N_5700,N_5250,N_5444);
nor U5701 (N_5701,N_5276,N_5250);
and U5702 (N_5702,N_5387,N_5473);
xor U5703 (N_5703,N_5471,N_5434);
nand U5704 (N_5704,N_5492,N_5400);
and U5705 (N_5705,N_5341,N_5386);
nand U5706 (N_5706,N_5334,N_5417);
or U5707 (N_5707,N_5405,N_5495);
and U5708 (N_5708,N_5349,N_5414);
nor U5709 (N_5709,N_5360,N_5252);
or U5710 (N_5710,N_5497,N_5367);
nand U5711 (N_5711,N_5288,N_5403);
and U5712 (N_5712,N_5307,N_5436);
and U5713 (N_5713,N_5296,N_5435);
and U5714 (N_5714,N_5344,N_5471);
or U5715 (N_5715,N_5338,N_5280);
and U5716 (N_5716,N_5367,N_5498);
nor U5717 (N_5717,N_5367,N_5377);
nand U5718 (N_5718,N_5334,N_5471);
nor U5719 (N_5719,N_5418,N_5357);
nor U5720 (N_5720,N_5375,N_5371);
nand U5721 (N_5721,N_5284,N_5359);
and U5722 (N_5722,N_5288,N_5435);
or U5723 (N_5723,N_5469,N_5380);
nand U5724 (N_5724,N_5486,N_5378);
nand U5725 (N_5725,N_5491,N_5470);
and U5726 (N_5726,N_5377,N_5391);
and U5727 (N_5727,N_5251,N_5449);
nand U5728 (N_5728,N_5304,N_5462);
nor U5729 (N_5729,N_5481,N_5344);
nor U5730 (N_5730,N_5332,N_5391);
nand U5731 (N_5731,N_5312,N_5297);
nand U5732 (N_5732,N_5350,N_5436);
or U5733 (N_5733,N_5415,N_5310);
xor U5734 (N_5734,N_5383,N_5490);
or U5735 (N_5735,N_5262,N_5386);
nor U5736 (N_5736,N_5466,N_5455);
and U5737 (N_5737,N_5259,N_5408);
nand U5738 (N_5738,N_5421,N_5443);
nor U5739 (N_5739,N_5442,N_5479);
nand U5740 (N_5740,N_5295,N_5496);
nand U5741 (N_5741,N_5495,N_5484);
or U5742 (N_5742,N_5405,N_5293);
and U5743 (N_5743,N_5453,N_5351);
and U5744 (N_5744,N_5298,N_5485);
or U5745 (N_5745,N_5451,N_5313);
nand U5746 (N_5746,N_5377,N_5301);
nor U5747 (N_5747,N_5309,N_5273);
nand U5748 (N_5748,N_5458,N_5485);
nor U5749 (N_5749,N_5283,N_5423);
or U5750 (N_5750,N_5545,N_5663);
or U5751 (N_5751,N_5664,N_5748);
and U5752 (N_5752,N_5525,N_5673);
and U5753 (N_5753,N_5518,N_5665);
xnor U5754 (N_5754,N_5612,N_5619);
nor U5755 (N_5755,N_5745,N_5668);
and U5756 (N_5756,N_5586,N_5740);
or U5757 (N_5757,N_5706,N_5692);
nor U5758 (N_5758,N_5542,N_5615);
or U5759 (N_5759,N_5544,N_5656);
nand U5760 (N_5760,N_5547,N_5608);
or U5761 (N_5761,N_5594,N_5725);
nor U5762 (N_5762,N_5620,N_5727);
or U5763 (N_5763,N_5502,N_5593);
nand U5764 (N_5764,N_5702,N_5667);
and U5765 (N_5765,N_5681,N_5738);
xor U5766 (N_5766,N_5685,N_5712);
or U5767 (N_5767,N_5647,N_5552);
nand U5768 (N_5768,N_5556,N_5659);
nand U5769 (N_5769,N_5573,N_5511);
and U5770 (N_5770,N_5504,N_5603);
or U5771 (N_5771,N_5650,N_5683);
and U5772 (N_5772,N_5626,N_5676);
or U5773 (N_5773,N_5624,N_5666);
or U5774 (N_5774,N_5597,N_5590);
nand U5775 (N_5775,N_5661,N_5598);
nor U5776 (N_5776,N_5694,N_5737);
nor U5777 (N_5777,N_5609,N_5730);
or U5778 (N_5778,N_5601,N_5582);
or U5779 (N_5779,N_5526,N_5679);
xor U5780 (N_5780,N_5726,N_5648);
nand U5781 (N_5781,N_5691,N_5690);
or U5782 (N_5782,N_5560,N_5553);
nor U5783 (N_5783,N_5527,N_5651);
or U5784 (N_5784,N_5655,N_5600);
and U5785 (N_5785,N_5623,N_5522);
or U5786 (N_5786,N_5696,N_5529);
or U5787 (N_5787,N_5572,N_5705);
nand U5788 (N_5788,N_5640,N_5537);
nor U5789 (N_5789,N_5717,N_5596);
nor U5790 (N_5790,N_5704,N_5652);
nor U5791 (N_5791,N_5606,N_5604);
and U5792 (N_5792,N_5563,N_5741);
xor U5793 (N_5793,N_5549,N_5639);
xor U5794 (N_5794,N_5575,N_5589);
and U5795 (N_5795,N_5568,N_5703);
nor U5796 (N_5796,N_5687,N_5524);
and U5797 (N_5797,N_5627,N_5714);
xnor U5798 (N_5798,N_5610,N_5660);
nand U5799 (N_5799,N_5557,N_5721);
or U5800 (N_5800,N_5645,N_5658);
and U5801 (N_5801,N_5543,N_5503);
and U5802 (N_5802,N_5551,N_5535);
xnor U5803 (N_5803,N_5585,N_5709);
nand U5804 (N_5804,N_5622,N_5718);
nand U5805 (N_5805,N_5588,N_5538);
or U5806 (N_5806,N_5574,N_5613);
and U5807 (N_5807,N_5630,N_5695);
nand U5808 (N_5808,N_5719,N_5617);
and U5809 (N_5809,N_5599,N_5723);
or U5810 (N_5810,N_5662,N_5735);
nor U5811 (N_5811,N_5644,N_5716);
xnor U5812 (N_5812,N_5583,N_5744);
nor U5813 (N_5813,N_5672,N_5711);
and U5814 (N_5814,N_5528,N_5578);
and U5815 (N_5815,N_5633,N_5724);
nand U5816 (N_5816,N_5515,N_5634);
nand U5817 (N_5817,N_5629,N_5713);
and U5818 (N_5818,N_5671,N_5602);
nand U5819 (N_5819,N_5507,N_5517);
xor U5820 (N_5820,N_5616,N_5592);
and U5821 (N_5821,N_5567,N_5684);
nor U5822 (N_5822,N_5708,N_5570);
and U5823 (N_5823,N_5631,N_5710);
or U5824 (N_5824,N_5732,N_5577);
nand U5825 (N_5825,N_5584,N_5506);
or U5826 (N_5826,N_5611,N_5564);
nor U5827 (N_5827,N_5579,N_5731);
nand U5828 (N_5828,N_5698,N_5642);
nand U5829 (N_5829,N_5500,N_5733);
or U5830 (N_5830,N_5566,N_5657);
nor U5831 (N_5831,N_5635,N_5505);
and U5832 (N_5832,N_5519,N_5734);
nand U5833 (N_5833,N_5674,N_5530);
nand U5834 (N_5834,N_5536,N_5675);
xnor U5835 (N_5835,N_5746,N_5539);
and U5836 (N_5836,N_5653,N_5677);
or U5837 (N_5837,N_5632,N_5621);
nor U5838 (N_5838,N_5540,N_5722);
nand U5839 (N_5839,N_5701,N_5670);
nor U5840 (N_5840,N_5641,N_5680);
nor U5841 (N_5841,N_5739,N_5513);
nand U5842 (N_5842,N_5646,N_5747);
or U5843 (N_5843,N_5689,N_5686);
nor U5844 (N_5844,N_5546,N_5554);
nand U5845 (N_5845,N_5532,N_5576);
nand U5846 (N_5846,N_5729,N_5520);
and U5847 (N_5847,N_5533,N_5669);
xnor U5848 (N_5848,N_5595,N_5605);
nand U5849 (N_5849,N_5742,N_5749);
or U5850 (N_5850,N_5587,N_5521);
and U5851 (N_5851,N_5580,N_5514);
and U5852 (N_5852,N_5501,N_5565);
nand U5853 (N_5853,N_5720,N_5509);
and U5854 (N_5854,N_5736,N_5649);
nor U5855 (N_5855,N_5561,N_5558);
nor U5856 (N_5856,N_5699,N_5510);
and U5857 (N_5857,N_5548,N_5555);
or U5858 (N_5858,N_5591,N_5707);
or U5859 (N_5859,N_5614,N_5654);
nor U5860 (N_5860,N_5728,N_5571);
and U5861 (N_5861,N_5607,N_5637);
and U5862 (N_5862,N_5559,N_5678);
and U5863 (N_5863,N_5743,N_5636);
nor U5864 (N_5864,N_5697,N_5638);
or U5865 (N_5865,N_5531,N_5569);
nand U5866 (N_5866,N_5700,N_5523);
nor U5867 (N_5867,N_5508,N_5581);
nor U5868 (N_5868,N_5682,N_5618);
xor U5869 (N_5869,N_5688,N_5562);
nor U5870 (N_5870,N_5512,N_5625);
xnor U5871 (N_5871,N_5541,N_5693);
nor U5872 (N_5872,N_5534,N_5628);
nand U5873 (N_5873,N_5643,N_5550);
nand U5874 (N_5874,N_5715,N_5516);
and U5875 (N_5875,N_5660,N_5613);
nand U5876 (N_5876,N_5561,N_5579);
or U5877 (N_5877,N_5637,N_5554);
nand U5878 (N_5878,N_5531,N_5623);
or U5879 (N_5879,N_5632,N_5532);
nand U5880 (N_5880,N_5713,N_5529);
nand U5881 (N_5881,N_5600,N_5675);
nand U5882 (N_5882,N_5707,N_5540);
and U5883 (N_5883,N_5746,N_5500);
or U5884 (N_5884,N_5605,N_5666);
nor U5885 (N_5885,N_5590,N_5603);
or U5886 (N_5886,N_5588,N_5700);
nand U5887 (N_5887,N_5511,N_5655);
and U5888 (N_5888,N_5681,N_5579);
nand U5889 (N_5889,N_5720,N_5619);
xor U5890 (N_5890,N_5729,N_5715);
nand U5891 (N_5891,N_5608,N_5699);
or U5892 (N_5892,N_5502,N_5672);
xnor U5893 (N_5893,N_5712,N_5686);
and U5894 (N_5894,N_5541,N_5617);
nand U5895 (N_5895,N_5687,N_5622);
and U5896 (N_5896,N_5630,N_5623);
or U5897 (N_5897,N_5524,N_5537);
nand U5898 (N_5898,N_5627,N_5547);
or U5899 (N_5899,N_5571,N_5542);
nand U5900 (N_5900,N_5717,N_5618);
and U5901 (N_5901,N_5614,N_5588);
nand U5902 (N_5902,N_5595,N_5638);
nor U5903 (N_5903,N_5597,N_5546);
or U5904 (N_5904,N_5722,N_5584);
or U5905 (N_5905,N_5601,N_5503);
nand U5906 (N_5906,N_5664,N_5532);
nor U5907 (N_5907,N_5685,N_5573);
nand U5908 (N_5908,N_5668,N_5722);
or U5909 (N_5909,N_5510,N_5504);
nor U5910 (N_5910,N_5633,N_5670);
xnor U5911 (N_5911,N_5632,N_5528);
and U5912 (N_5912,N_5548,N_5626);
nor U5913 (N_5913,N_5651,N_5579);
and U5914 (N_5914,N_5520,N_5536);
nor U5915 (N_5915,N_5696,N_5547);
or U5916 (N_5916,N_5657,N_5675);
nor U5917 (N_5917,N_5575,N_5619);
and U5918 (N_5918,N_5577,N_5678);
and U5919 (N_5919,N_5739,N_5743);
nor U5920 (N_5920,N_5690,N_5671);
nor U5921 (N_5921,N_5743,N_5622);
xor U5922 (N_5922,N_5673,N_5661);
nand U5923 (N_5923,N_5717,N_5580);
nand U5924 (N_5924,N_5517,N_5627);
and U5925 (N_5925,N_5513,N_5608);
or U5926 (N_5926,N_5658,N_5725);
nand U5927 (N_5927,N_5671,N_5538);
or U5928 (N_5928,N_5732,N_5542);
or U5929 (N_5929,N_5717,N_5506);
nand U5930 (N_5930,N_5705,N_5738);
nand U5931 (N_5931,N_5656,N_5607);
nand U5932 (N_5932,N_5627,N_5678);
nand U5933 (N_5933,N_5508,N_5543);
nand U5934 (N_5934,N_5616,N_5530);
nor U5935 (N_5935,N_5527,N_5525);
nand U5936 (N_5936,N_5693,N_5675);
or U5937 (N_5937,N_5601,N_5573);
nand U5938 (N_5938,N_5656,N_5708);
nand U5939 (N_5939,N_5618,N_5539);
nand U5940 (N_5940,N_5741,N_5517);
or U5941 (N_5941,N_5651,N_5567);
nor U5942 (N_5942,N_5649,N_5746);
nand U5943 (N_5943,N_5695,N_5593);
and U5944 (N_5944,N_5731,N_5540);
nor U5945 (N_5945,N_5557,N_5708);
nor U5946 (N_5946,N_5665,N_5591);
xor U5947 (N_5947,N_5553,N_5577);
or U5948 (N_5948,N_5541,N_5627);
and U5949 (N_5949,N_5664,N_5583);
and U5950 (N_5950,N_5682,N_5559);
or U5951 (N_5951,N_5707,N_5558);
and U5952 (N_5952,N_5724,N_5681);
xnor U5953 (N_5953,N_5726,N_5678);
and U5954 (N_5954,N_5746,N_5608);
and U5955 (N_5955,N_5730,N_5566);
nor U5956 (N_5956,N_5646,N_5681);
nand U5957 (N_5957,N_5560,N_5686);
or U5958 (N_5958,N_5693,N_5733);
nand U5959 (N_5959,N_5694,N_5666);
and U5960 (N_5960,N_5554,N_5548);
and U5961 (N_5961,N_5526,N_5570);
nor U5962 (N_5962,N_5623,N_5559);
and U5963 (N_5963,N_5602,N_5500);
nand U5964 (N_5964,N_5656,N_5565);
nand U5965 (N_5965,N_5629,N_5742);
nor U5966 (N_5966,N_5630,N_5564);
and U5967 (N_5967,N_5634,N_5741);
nor U5968 (N_5968,N_5525,N_5560);
xnor U5969 (N_5969,N_5526,N_5540);
nor U5970 (N_5970,N_5632,N_5736);
nor U5971 (N_5971,N_5667,N_5726);
nor U5972 (N_5972,N_5642,N_5594);
nand U5973 (N_5973,N_5586,N_5508);
and U5974 (N_5974,N_5721,N_5578);
and U5975 (N_5975,N_5687,N_5740);
nand U5976 (N_5976,N_5565,N_5732);
or U5977 (N_5977,N_5523,N_5547);
nand U5978 (N_5978,N_5731,N_5670);
nor U5979 (N_5979,N_5555,N_5602);
and U5980 (N_5980,N_5610,N_5516);
nand U5981 (N_5981,N_5547,N_5545);
xor U5982 (N_5982,N_5526,N_5527);
nand U5983 (N_5983,N_5691,N_5585);
or U5984 (N_5984,N_5593,N_5637);
or U5985 (N_5985,N_5516,N_5521);
and U5986 (N_5986,N_5559,N_5747);
nand U5987 (N_5987,N_5592,N_5574);
nor U5988 (N_5988,N_5581,N_5579);
xnor U5989 (N_5989,N_5666,N_5576);
and U5990 (N_5990,N_5540,N_5699);
nand U5991 (N_5991,N_5514,N_5664);
and U5992 (N_5992,N_5501,N_5597);
nand U5993 (N_5993,N_5647,N_5559);
nand U5994 (N_5994,N_5631,N_5520);
and U5995 (N_5995,N_5742,N_5560);
xnor U5996 (N_5996,N_5649,N_5506);
nand U5997 (N_5997,N_5515,N_5565);
or U5998 (N_5998,N_5727,N_5713);
or U5999 (N_5999,N_5570,N_5689);
nor U6000 (N_6000,N_5918,N_5862);
nand U6001 (N_6001,N_5794,N_5785);
or U6002 (N_6002,N_5905,N_5786);
nor U6003 (N_6003,N_5756,N_5939);
xnor U6004 (N_6004,N_5961,N_5945);
xor U6005 (N_6005,N_5814,N_5885);
nand U6006 (N_6006,N_5847,N_5942);
or U6007 (N_6007,N_5883,N_5988);
nand U6008 (N_6008,N_5818,N_5992);
or U6009 (N_6009,N_5788,N_5768);
or U6010 (N_6010,N_5861,N_5923);
nor U6011 (N_6011,N_5895,N_5835);
nand U6012 (N_6012,N_5770,N_5948);
or U6013 (N_6013,N_5826,N_5931);
xnor U6014 (N_6014,N_5886,N_5804);
nand U6015 (N_6015,N_5935,N_5878);
or U6016 (N_6016,N_5784,N_5852);
or U6017 (N_6017,N_5925,N_5975);
and U6018 (N_6018,N_5901,N_5860);
or U6019 (N_6019,N_5941,N_5867);
and U6020 (N_6020,N_5970,N_5985);
and U6021 (N_6021,N_5780,N_5774);
or U6022 (N_6022,N_5787,N_5930);
nand U6023 (N_6023,N_5772,N_5778);
nor U6024 (N_6024,N_5877,N_5789);
xor U6025 (N_6025,N_5907,N_5954);
nor U6026 (N_6026,N_5953,N_5764);
nor U6027 (N_6027,N_5868,N_5910);
or U6028 (N_6028,N_5996,N_5915);
nor U6029 (N_6029,N_5997,N_5932);
nand U6030 (N_6030,N_5851,N_5916);
or U6031 (N_6031,N_5872,N_5995);
and U6032 (N_6032,N_5924,N_5849);
nand U6033 (N_6033,N_5951,N_5783);
nand U6034 (N_6034,N_5928,N_5803);
nand U6035 (N_6035,N_5882,N_5856);
nor U6036 (N_6036,N_5834,N_5864);
and U6037 (N_6037,N_5810,N_5753);
nor U6038 (N_6038,N_5972,N_5936);
nand U6039 (N_6039,N_5974,N_5843);
nand U6040 (N_6040,N_5919,N_5822);
and U6041 (N_6041,N_5800,N_5828);
nor U6042 (N_6042,N_5891,N_5889);
and U6043 (N_6043,N_5806,N_5871);
or U6044 (N_6044,N_5848,N_5993);
and U6045 (N_6045,N_5781,N_5902);
nand U6046 (N_6046,N_5755,N_5884);
or U6047 (N_6047,N_5824,N_5807);
nor U6048 (N_6048,N_5790,N_5754);
nand U6049 (N_6049,N_5782,N_5898);
or U6050 (N_6050,N_5816,N_5908);
xor U6051 (N_6051,N_5855,N_5842);
or U6052 (N_6052,N_5829,N_5765);
xor U6053 (N_6053,N_5815,N_5840);
nand U6054 (N_6054,N_5808,N_5964);
nor U6055 (N_6055,N_5944,N_5926);
nor U6056 (N_6056,N_5998,N_5811);
nor U6057 (N_6057,N_5809,N_5832);
and U6058 (N_6058,N_5821,N_5999);
and U6059 (N_6059,N_5759,N_5962);
nor U6060 (N_6060,N_5819,N_5771);
nand U6061 (N_6061,N_5767,N_5792);
or U6062 (N_6062,N_5853,N_5960);
xor U6063 (N_6063,N_5823,N_5817);
nand U6064 (N_6064,N_5946,N_5986);
nor U6065 (N_6065,N_5760,N_5874);
nor U6066 (N_6066,N_5865,N_5949);
or U6067 (N_6067,N_5831,N_5869);
and U6068 (N_6068,N_5906,N_5887);
nand U6069 (N_6069,N_5921,N_5904);
nand U6070 (N_6070,N_5825,N_5897);
and U6071 (N_6071,N_5799,N_5859);
or U6072 (N_6072,N_5796,N_5967);
nor U6073 (N_6073,N_5894,N_5977);
nand U6074 (N_6074,N_5980,N_5779);
or U6075 (N_6075,N_5845,N_5857);
and U6076 (N_6076,N_5888,N_5952);
or U6077 (N_6077,N_5890,N_5973);
or U6078 (N_6078,N_5879,N_5955);
xor U6079 (N_6079,N_5933,N_5795);
or U6080 (N_6080,N_5776,N_5989);
nor U6081 (N_6081,N_5758,N_5751);
or U6082 (N_6082,N_5880,N_5802);
and U6083 (N_6083,N_5797,N_5854);
xnor U6084 (N_6084,N_5801,N_5820);
nor U6085 (N_6085,N_5947,N_5841);
nor U6086 (N_6086,N_5994,N_5899);
xnor U6087 (N_6087,N_5892,N_5846);
and U6088 (N_6088,N_5775,N_5893);
nor U6089 (N_6089,N_5982,N_5863);
and U6090 (N_6090,N_5833,N_5757);
nand U6091 (N_6091,N_5913,N_5762);
or U6092 (N_6092,N_5876,N_5940);
nor U6093 (N_6093,N_5763,N_5870);
xnor U6094 (N_6094,N_5793,N_5896);
and U6095 (N_6095,N_5903,N_5912);
nor U6096 (N_6096,N_5881,N_5837);
xnor U6097 (N_6097,N_5812,N_5965);
xor U6098 (N_6098,N_5805,N_5858);
or U6099 (N_6099,N_5791,N_5766);
nand U6100 (N_6100,N_5979,N_5917);
nand U6101 (N_6101,N_5978,N_5927);
and U6102 (N_6102,N_5963,N_5950);
nand U6103 (N_6103,N_5866,N_5971);
or U6104 (N_6104,N_5911,N_5830);
nand U6105 (N_6105,N_5922,N_5990);
nor U6106 (N_6106,N_5934,N_5914);
nor U6107 (N_6107,N_5957,N_5813);
and U6108 (N_6108,N_5966,N_5909);
or U6109 (N_6109,N_5968,N_5850);
nor U6110 (N_6110,N_5838,N_5983);
or U6111 (N_6111,N_5929,N_5777);
nor U6112 (N_6112,N_5836,N_5873);
and U6113 (N_6113,N_5943,N_5798);
nand U6114 (N_6114,N_5844,N_5750);
and U6115 (N_6115,N_5991,N_5752);
nand U6116 (N_6116,N_5937,N_5875);
xnor U6117 (N_6117,N_5900,N_5956);
or U6118 (N_6118,N_5769,N_5920);
or U6119 (N_6119,N_5938,N_5969);
nand U6120 (N_6120,N_5761,N_5976);
nand U6121 (N_6121,N_5959,N_5981);
or U6122 (N_6122,N_5827,N_5958);
and U6123 (N_6123,N_5987,N_5984);
nand U6124 (N_6124,N_5773,N_5839);
nor U6125 (N_6125,N_5877,N_5970);
or U6126 (N_6126,N_5950,N_5784);
or U6127 (N_6127,N_5850,N_5922);
nand U6128 (N_6128,N_5876,N_5992);
and U6129 (N_6129,N_5819,N_5807);
nor U6130 (N_6130,N_5899,N_5999);
and U6131 (N_6131,N_5893,N_5819);
or U6132 (N_6132,N_5754,N_5983);
nor U6133 (N_6133,N_5873,N_5842);
and U6134 (N_6134,N_5835,N_5773);
nand U6135 (N_6135,N_5898,N_5975);
or U6136 (N_6136,N_5828,N_5871);
nor U6137 (N_6137,N_5853,N_5967);
xnor U6138 (N_6138,N_5907,N_5808);
and U6139 (N_6139,N_5762,N_5824);
or U6140 (N_6140,N_5861,N_5794);
nand U6141 (N_6141,N_5808,N_5835);
nor U6142 (N_6142,N_5831,N_5936);
and U6143 (N_6143,N_5857,N_5987);
nor U6144 (N_6144,N_5882,N_5956);
nand U6145 (N_6145,N_5950,N_5937);
nand U6146 (N_6146,N_5930,N_5770);
nand U6147 (N_6147,N_5867,N_5779);
or U6148 (N_6148,N_5799,N_5821);
nand U6149 (N_6149,N_5950,N_5871);
nor U6150 (N_6150,N_5829,N_5893);
and U6151 (N_6151,N_5822,N_5977);
nand U6152 (N_6152,N_5963,N_5848);
or U6153 (N_6153,N_5885,N_5772);
or U6154 (N_6154,N_5928,N_5850);
nor U6155 (N_6155,N_5938,N_5868);
nand U6156 (N_6156,N_5822,N_5763);
nand U6157 (N_6157,N_5861,N_5971);
xnor U6158 (N_6158,N_5979,N_5835);
xor U6159 (N_6159,N_5841,N_5956);
and U6160 (N_6160,N_5984,N_5878);
xor U6161 (N_6161,N_5968,N_5764);
or U6162 (N_6162,N_5786,N_5983);
and U6163 (N_6163,N_5894,N_5786);
and U6164 (N_6164,N_5982,N_5771);
and U6165 (N_6165,N_5866,N_5876);
nand U6166 (N_6166,N_5798,N_5931);
or U6167 (N_6167,N_5779,N_5952);
nand U6168 (N_6168,N_5816,N_5919);
nand U6169 (N_6169,N_5905,N_5757);
xnor U6170 (N_6170,N_5806,N_5888);
nand U6171 (N_6171,N_5857,N_5898);
or U6172 (N_6172,N_5954,N_5784);
nand U6173 (N_6173,N_5974,N_5827);
and U6174 (N_6174,N_5960,N_5889);
nand U6175 (N_6175,N_5819,N_5798);
or U6176 (N_6176,N_5901,N_5855);
or U6177 (N_6177,N_5872,N_5802);
and U6178 (N_6178,N_5961,N_5939);
or U6179 (N_6179,N_5913,N_5866);
nor U6180 (N_6180,N_5766,N_5943);
or U6181 (N_6181,N_5774,N_5790);
and U6182 (N_6182,N_5960,N_5855);
nand U6183 (N_6183,N_5859,N_5768);
and U6184 (N_6184,N_5895,N_5924);
or U6185 (N_6185,N_5805,N_5904);
nand U6186 (N_6186,N_5941,N_5791);
nand U6187 (N_6187,N_5919,N_5856);
or U6188 (N_6188,N_5815,N_5884);
nand U6189 (N_6189,N_5863,N_5751);
xor U6190 (N_6190,N_5818,N_5766);
nand U6191 (N_6191,N_5883,N_5808);
and U6192 (N_6192,N_5980,N_5978);
xnor U6193 (N_6193,N_5754,N_5910);
nand U6194 (N_6194,N_5795,N_5759);
nor U6195 (N_6195,N_5874,N_5785);
nor U6196 (N_6196,N_5795,N_5784);
and U6197 (N_6197,N_5812,N_5862);
nand U6198 (N_6198,N_5828,N_5923);
and U6199 (N_6199,N_5972,N_5797);
or U6200 (N_6200,N_5908,N_5780);
nor U6201 (N_6201,N_5989,N_5951);
nand U6202 (N_6202,N_5810,N_5976);
xor U6203 (N_6203,N_5870,N_5899);
nand U6204 (N_6204,N_5774,N_5945);
and U6205 (N_6205,N_5963,N_5821);
nor U6206 (N_6206,N_5767,N_5865);
nor U6207 (N_6207,N_5984,N_5940);
or U6208 (N_6208,N_5996,N_5821);
nand U6209 (N_6209,N_5999,N_5879);
and U6210 (N_6210,N_5929,N_5916);
and U6211 (N_6211,N_5986,N_5987);
nand U6212 (N_6212,N_5947,N_5820);
nand U6213 (N_6213,N_5808,N_5973);
xor U6214 (N_6214,N_5840,N_5931);
xnor U6215 (N_6215,N_5768,N_5779);
nor U6216 (N_6216,N_5888,N_5938);
or U6217 (N_6217,N_5879,N_5993);
or U6218 (N_6218,N_5870,N_5856);
and U6219 (N_6219,N_5778,N_5897);
or U6220 (N_6220,N_5926,N_5853);
and U6221 (N_6221,N_5764,N_5836);
or U6222 (N_6222,N_5932,N_5951);
and U6223 (N_6223,N_5881,N_5976);
and U6224 (N_6224,N_5952,N_5803);
or U6225 (N_6225,N_5773,N_5998);
nand U6226 (N_6226,N_5873,N_5800);
nor U6227 (N_6227,N_5918,N_5856);
or U6228 (N_6228,N_5766,N_5768);
or U6229 (N_6229,N_5922,N_5966);
or U6230 (N_6230,N_5751,N_5871);
nand U6231 (N_6231,N_5974,N_5770);
and U6232 (N_6232,N_5775,N_5840);
or U6233 (N_6233,N_5889,N_5930);
nand U6234 (N_6234,N_5889,N_5798);
nand U6235 (N_6235,N_5786,N_5958);
nand U6236 (N_6236,N_5961,N_5973);
or U6237 (N_6237,N_5785,N_5902);
nand U6238 (N_6238,N_5906,N_5969);
and U6239 (N_6239,N_5827,N_5930);
and U6240 (N_6240,N_5788,N_5974);
nand U6241 (N_6241,N_5991,N_5864);
or U6242 (N_6242,N_5917,N_5763);
xor U6243 (N_6243,N_5892,N_5822);
and U6244 (N_6244,N_5822,N_5854);
xor U6245 (N_6245,N_5959,N_5797);
nor U6246 (N_6246,N_5947,N_5907);
and U6247 (N_6247,N_5890,N_5760);
nand U6248 (N_6248,N_5819,N_5815);
and U6249 (N_6249,N_5916,N_5923);
nor U6250 (N_6250,N_6238,N_6022);
nor U6251 (N_6251,N_6227,N_6013);
and U6252 (N_6252,N_6019,N_6021);
and U6253 (N_6253,N_6216,N_6158);
nor U6254 (N_6254,N_6240,N_6125);
and U6255 (N_6255,N_6218,N_6073);
nor U6256 (N_6256,N_6220,N_6152);
and U6257 (N_6257,N_6169,N_6214);
nor U6258 (N_6258,N_6011,N_6069);
nor U6259 (N_6259,N_6053,N_6048);
nand U6260 (N_6260,N_6050,N_6204);
nand U6261 (N_6261,N_6217,N_6180);
or U6262 (N_6262,N_6185,N_6042);
nand U6263 (N_6263,N_6175,N_6205);
nor U6264 (N_6264,N_6004,N_6157);
or U6265 (N_6265,N_6224,N_6056);
nor U6266 (N_6266,N_6115,N_6028);
nand U6267 (N_6267,N_6101,N_6191);
nor U6268 (N_6268,N_6201,N_6149);
or U6269 (N_6269,N_6159,N_6140);
xor U6270 (N_6270,N_6243,N_6009);
and U6271 (N_6271,N_6138,N_6177);
and U6272 (N_6272,N_6110,N_6148);
and U6273 (N_6273,N_6129,N_6064);
xnor U6274 (N_6274,N_6198,N_6131);
and U6275 (N_6275,N_6135,N_6167);
nand U6276 (N_6276,N_6113,N_6223);
nand U6277 (N_6277,N_6104,N_6040);
nor U6278 (N_6278,N_6139,N_6160);
xor U6279 (N_6279,N_6176,N_6183);
or U6280 (N_6280,N_6207,N_6033);
and U6281 (N_6281,N_6059,N_6174);
and U6282 (N_6282,N_6111,N_6061);
or U6283 (N_6283,N_6074,N_6194);
and U6284 (N_6284,N_6234,N_6147);
and U6285 (N_6285,N_6193,N_6086);
or U6286 (N_6286,N_6051,N_6249);
nand U6287 (N_6287,N_6245,N_6213);
nand U6288 (N_6288,N_6209,N_6170);
and U6289 (N_6289,N_6195,N_6229);
nor U6290 (N_6290,N_6097,N_6079);
xnor U6291 (N_6291,N_6067,N_6047);
or U6292 (N_6292,N_6242,N_6016);
nand U6293 (N_6293,N_6102,N_6235);
nor U6294 (N_6294,N_6124,N_6150);
xor U6295 (N_6295,N_6117,N_6137);
and U6296 (N_6296,N_6200,N_6247);
nand U6297 (N_6297,N_6151,N_6038);
nand U6298 (N_6298,N_6092,N_6196);
or U6299 (N_6299,N_6060,N_6001);
and U6300 (N_6300,N_6121,N_6027);
nor U6301 (N_6301,N_6057,N_6142);
and U6302 (N_6302,N_6231,N_6202);
xor U6303 (N_6303,N_6046,N_6233);
nand U6304 (N_6304,N_6232,N_6164);
nand U6305 (N_6305,N_6029,N_6222);
xor U6306 (N_6306,N_6144,N_6211);
or U6307 (N_6307,N_6132,N_6237);
nor U6308 (N_6308,N_6017,N_6020);
and U6309 (N_6309,N_6078,N_6199);
or U6310 (N_6310,N_6099,N_6108);
or U6311 (N_6311,N_6153,N_6025);
nand U6312 (N_6312,N_6126,N_6036);
nand U6313 (N_6313,N_6094,N_6246);
xor U6314 (N_6314,N_6228,N_6130);
and U6315 (N_6315,N_6041,N_6003);
nand U6316 (N_6316,N_6244,N_6080);
and U6317 (N_6317,N_6122,N_6024);
nand U6318 (N_6318,N_6105,N_6189);
or U6319 (N_6319,N_6037,N_6184);
or U6320 (N_6320,N_6045,N_6081);
xnor U6321 (N_6321,N_6039,N_6058);
or U6322 (N_6322,N_6206,N_6109);
or U6323 (N_6323,N_6123,N_6187);
or U6324 (N_6324,N_6043,N_6212);
nand U6325 (N_6325,N_6171,N_6188);
nand U6326 (N_6326,N_6221,N_6141);
or U6327 (N_6327,N_6182,N_6178);
or U6328 (N_6328,N_6186,N_6192);
nand U6329 (N_6329,N_6119,N_6236);
xnor U6330 (N_6330,N_6156,N_6225);
nor U6331 (N_6331,N_6166,N_6095);
and U6332 (N_6332,N_6068,N_6098);
nor U6333 (N_6333,N_6049,N_6173);
or U6334 (N_6334,N_6035,N_6062);
or U6335 (N_6335,N_6026,N_6100);
or U6336 (N_6336,N_6179,N_6018);
and U6337 (N_6337,N_6063,N_6226);
and U6338 (N_6338,N_6168,N_6072);
nor U6339 (N_6339,N_6219,N_6143);
nor U6340 (N_6340,N_6076,N_6008);
or U6341 (N_6341,N_6203,N_6083);
nor U6342 (N_6342,N_6210,N_6114);
nand U6343 (N_6343,N_6002,N_6208);
xnor U6344 (N_6344,N_6055,N_6145);
nor U6345 (N_6345,N_6103,N_6087);
nand U6346 (N_6346,N_6084,N_6248);
or U6347 (N_6347,N_6155,N_6165);
nor U6348 (N_6348,N_6000,N_6136);
nor U6349 (N_6349,N_6012,N_6128);
nor U6350 (N_6350,N_6093,N_6118);
nor U6351 (N_6351,N_6023,N_6044);
nand U6352 (N_6352,N_6162,N_6120);
nor U6353 (N_6353,N_6082,N_6107);
nor U6354 (N_6354,N_6241,N_6070);
and U6355 (N_6355,N_6146,N_6065);
or U6356 (N_6356,N_6181,N_6230);
xor U6357 (N_6357,N_6075,N_6014);
nand U6358 (N_6358,N_6088,N_6015);
xor U6359 (N_6359,N_6032,N_6163);
xnor U6360 (N_6360,N_6090,N_6089);
and U6361 (N_6361,N_6116,N_6096);
nor U6362 (N_6362,N_6085,N_6172);
or U6363 (N_6363,N_6239,N_6066);
or U6364 (N_6364,N_6106,N_6197);
nor U6365 (N_6365,N_6030,N_6007);
or U6366 (N_6366,N_6006,N_6054);
or U6367 (N_6367,N_6190,N_6052);
or U6368 (N_6368,N_6071,N_6127);
nand U6369 (N_6369,N_6077,N_6031);
and U6370 (N_6370,N_6161,N_6134);
and U6371 (N_6371,N_6112,N_6215);
nor U6372 (N_6372,N_6133,N_6034);
nor U6373 (N_6373,N_6005,N_6010);
nor U6374 (N_6374,N_6154,N_6091);
xnor U6375 (N_6375,N_6190,N_6170);
or U6376 (N_6376,N_6241,N_6020);
and U6377 (N_6377,N_6166,N_6229);
nand U6378 (N_6378,N_6150,N_6068);
and U6379 (N_6379,N_6024,N_6151);
and U6380 (N_6380,N_6019,N_6222);
nand U6381 (N_6381,N_6201,N_6102);
nor U6382 (N_6382,N_6212,N_6169);
and U6383 (N_6383,N_6135,N_6139);
xnor U6384 (N_6384,N_6204,N_6094);
xor U6385 (N_6385,N_6193,N_6191);
nand U6386 (N_6386,N_6197,N_6118);
nor U6387 (N_6387,N_6108,N_6026);
or U6388 (N_6388,N_6101,N_6152);
and U6389 (N_6389,N_6244,N_6022);
nand U6390 (N_6390,N_6117,N_6213);
nand U6391 (N_6391,N_6036,N_6047);
nor U6392 (N_6392,N_6036,N_6025);
nor U6393 (N_6393,N_6025,N_6079);
nand U6394 (N_6394,N_6096,N_6066);
nand U6395 (N_6395,N_6206,N_6092);
nor U6396 (N_6396,N_6238,N_6204);
and U6397 (N_6397,N_6243,N_6084);
or U6398 (N_6398,N_6185,N_6169);
nand U6399 (N_6399,N_6038,N_6115);
nor U6400 (N_6400,N_6129,N_6121);
nand U6401 (N_6401,N_6248,N_6031);
nor U6402 (N_6402,N_6116,N_6052);
or U6403 (N_6403,N_6098,N_6108);
nand U6404 (N_6404,N_6038,N_6122);
nand U6405 (N_6405,N_6086,N_6115);
nor U6406 (N_6406,N_6137,N_6065);
nand U6407 (N_6407,N_6195,N_6113);
nand U6408 (N_6408,N_6123,N_6141);
and U6409 (N_6409,N_6063,N_6084);
or U6410 (N_6410,N_6244,N_6153);
or U6411 (N_6411,N_6210,N_6003);
or U6412 (N_6412,N_6066,N_6016);
and U6413 (N_6413,N_6020,N_6032);
nor U6414 (N_6414,N_6041,N_6160);
and U6415 (N_6415,N_6125,N_6008);
xnor U6416 (N_6416,N_6150,N_6248);
nor U6417 (N_6417,N_6146,N_6046);
or U6418 (N_6418,N_6036,N_6221);
and U6419 (N_6419,N_6057,N_6088);
nand U6420 (N_6420,N_6132,N_6097);
and U6421 (N_6421,N_6005,N_6224);
and U6422 (N_6422,N_6021,N_6035);
nor U6423 (N_6423,N_6083,N_6174);
and U6424 (N_6424,N_6224,N_6084);
and U6425 (N_6425,N_6210,N_6246);
or U6426 (N_6426,N_6191,N_6128);
xnor U6427 (N_6427,N_6072,N_6231);
nand U6428 (N_6428,N_6207,N_6098);
or U6429 (N_6429,N_6134,N_6150);
or U6430 (N_6430,N_6101,N_6083);
nor U6431 (N_6431,N_6236,N_6102);
nand U6432 (N_6432,N_6191,N_6162);
or U6433 (N_6433,N_6165,N_6005);
nor U6434 (N_6434,N_6120,N_6013);
or U6435 (N_6435,N_6225,N_6239);
nand U6436 (N_6436,N_6231,N_6046);
nand U6437 (N_6437,N_6124,N_6154);
and U6438 (N_6438,N_6143,N_6196);
nand U6439 (N_6439,N_6094,N_6126);
xor U6440 (N_6440,N_6207,N_6235);
and U6441 (N_6441,N_6021,N_6204);
nand U6442 (N_6442,N_6114,N_6198);
and U6443 (N_6443,N_6144,N_6240);
nand U6444 (N_6444,N_6125,N_6186);
nor U6445 (N_6445,N_6191,N_6039);
nand U6446 (N_6446,N_6218,N_6215);
nand U6447 (N_6447,N_6066,N_6107);
or U6448 (N_6448,N_6214,N_6124);
nor U6449 (N_6449,N_6158,N_6174);
and U6450 (N_6450,N_6224,N_6037);
and U6451 (N_6451,N_6179,N_6045);
or U6452 (N_6452,N_6004,N_6191);
nor U6453 (N_6453,N_6141,N_6101);
or U6454 (N_6454,N_6117,N_6050);
xnor U6455 (N_6455,N_6052,N_6177);
nand U6456 (N_6456,N_6134,N_6142);
nor U6457 (N_6457,N_6039,N_6017);
nor U6458 (N_6458,N_6142,N_6110);
nand U6459 (N_6459,N_6183,N_6089);
xor U6460 (N_6460,N_6085,N_6048);
or U6461 (N_6461,N_6228,N_6058);
or U6462 (N_6462,N_6149,N_6082);
or U6463 (N_6463,N_6238,N_6090);
and U6464 (N_6464,N_6214,N_6237);
xor U6465 (N_6465,N_6176,N_6022);
nand U6466 (N_6466,N_6219,N_6070);
xnor U6467 (N_6467,N_6168,N_6057);
nand U6468 (N_6468,N_6038,N_6014);
nor U6469 (N_6469,N_6007,N_6238);
or U6470 (N_6470,N_6120,N_6035);
and U6471 (N_6471,N_6091,N_6152);
and U6472 (N_6472,N_6051,N_6179);
nand U6473 (N_6473,N_6247,N_6126);
or U6474 (N_6474,N_6094,N_6239);
and U6475 (N_6475,N_6162,N_6123);
and U6476 (N_6476,N_6196,N_6164);
or U6477 (N_6477,N_6033,N_6123);
nand U6478 (N_6478,N_6230,N_6051);
and U6479 (N_6479,N_6168,N_6015);
nand U6480 (N_6480,N_6186,N_6058);
xnor U6481 (N_6481,N_6112,N_6220);
or U6482 (N_6482,N_6182,N_6120);
xnor U6483 (N_6483,N_6068,N_6041);
nor U6484 (N_6484,N_6123,N_6226);
and U6485 (N_6485,N_6107,N_6245);
nand U6486 (N_6486,N_6106,N_6203);
or U6487 (N_6487,N_6015,N_6046);
nor U6488 (N_6488,N_6106,N_6032);
nor U6489 (N_6489,N_6021,N_6193);
nand U6490 (N_6490,N_6104,N_6032);
nand U6491 (N_6491,N_6019,N_6009);
nor U6492 (N_6492,N_6067,N_6019);
nand U6493 (N_6493,N_6187,N_6163);
xor U6494 (N_6494,N_6020,N_6090);
nor U6495 (N_6495,N_6223,N_6173);
nor U6496 (N_6496,N_6230,N_6157);
nor U6497 (N_6497,N_6098,N_6051);
nand U6498 (N_6498,N_6213,N_6176);
or U6499 (N_6499,N_6060,N_6110);
or U6500 (N_6500,N_6493,N_6402);
or U6501 (N_6501,N_6406,N_6453);
or U6502 (N_6502,N_6262,N_6319);
nor U6503 (N_6503,N_6255,N_6480);
or U6504 (N_6504,N_6369,N_6428);
or U6505 (N_6505,N_6296,N_6275);
nand U6506 (N_6506,N_6434,N_6418);
nand U6507 (N_6507,N_6318,N_6464);
nor U6508 (N_6508,N_6450,N_6397);
and U6509 (N_6509,N_6462,N_6423);
nand U6510 (N_6510,N_6472,N_6494);
or U6511 (N_6511,N_6475,N_6299);
nand U6512 (N_6512,N_6270,N_6272);
and U6513 (N_6513,N_6457,N_6368);
nand U6514 (N_6514,N_6370,N_6485);
nand U6515 (N_6515,N_6348,N_6286);
xnor U6516 (N_6516,N_6306,N_6358);
nand U6517 (N_6517,N_6456,N_6386);
and U6518 (N_6518,N_6400,N_6335);
nor U6519 (N_6519,N_6304,N_6316);
or U6520 (N_6520,N_6308,N_6284);
xnor U6521 (N_6521,N_6341,N_6343);
xnor U6522 (N_6522,N_6467,N_6412);
and U6523 (N_6523,N_6401,N_6411);
nand U6524 (N_6524,N_6263,N_6486);
xor U6525 (N_6525,N_6357,N_6309);
and U6526 (N_6526,N_6466,N_6391);
nand U6527 (N_6527,N_6461,N_6322);
nand U6528 (N_6528,N_6291,N_6327);
nor U6529 (N_6529,N_6484,N_6459);
nor U6530 (N_6530,N_6435,N_6429);
or U6531 (N_6531,N_6394,N_6372);
or U6532 (N_6532,N_6392,N_6454);
nand U6533 (N_6533,N_6385,N_6478);
or U6534 (N_6534,N_6452,N_6324);
nor U6535 (N_6535,N_6366,N_6265);
or U6536 (N_6536,N_6387,N_6251);
nor U6537 (N_6537,N_6356,N_6274);
or U6538 (N_6538,N_6490,N_6367);
nor U6539 (N_6539,N_6378,N_6253);
or U6540 (N_6540,N_6381,N_6463);
or U6541 (N_6541,N_6331,N_6476);
nand U6542 (N_6542,N_6442,N_6474);
nand U6543 (N_6543,N_6311,N_6469);
nand U6544 (N_6544,N_6393,N_6373);
and U6545 (N_6545,N_6376,N_6471);
nor U6546 (N_6546,N_6436,N_6482);
and U6547 (N_6547,N_6266,N_6346);
nor U6548 (N_6548,N_6354,N_6427);
nand U6549 (N_6549,N_6420,N_6439);
nor U6550 (N_6550,N_6398,N_6300);
or U6551 (N_6551,N_6399,N_6279);
and U6552 (N_6552,N_6430,N_6336);
nor U6553 (N_6553,N_6325,N_6499);
or U6554 (N_6554,N_6449,N_6421);
nor U6555 (N_6555,N_6285,N_6252);
or U6556 (N_6556,N_6277,N_6440);
nand U6557 (N_6557,N_6473,N_6498);
xor U6558 (N_6558,N_6448,N_6298);
and U6559 (N_6559,N_6334,N_6329);
nand U6560 (N_6560,N_6477,N_6388);
nor U6561 (N_6561,N_6465,N_6353);
nand U6562 (N_6562,N_6384,N_6424);
nor U6563 (N_6563,N_6332,N_6441);
nor U6564 (N_6564,N_6405,N_6446);
and U6565 (N_6565,N_6416,N_6347);
xnor U6566 (N_6566,N_6414,N_6264);
nor U6567 (N_6567,N_6433,N_6413);
nor U6568 (N_6568,N_6451,N_6349);
and U6569 (N_6569,N_6288,N_6377);
nand U6570 (N_6570,N_6407,N_6403);
nor U6571 (N_6571,N_6330,N_6293);
and U6572 (N_6572,N_6488,N_6437);
or U6573 (N_6573,N_6497,N_6305);
or U6574 (N_6574,N_6491,N_6294);
or U6575 (N_6575,N_6315,N_6282);
nand U6576 (N_6576,N_6408,N_6438);
or U6577 (N_6577,N_6390,N_6383);
nor U6578 (N_6578,N_6364,N_6261);
nand U6579 (N_6579,N_6458,N_6404);
and U6580 (N_6580,N_6443,N_6268);
and U6581 (N_6581,N_6321,N_6415);
nand U6582 (N_6582,N_6361,N_6360);
or U6583 (N_6583,N_6307,N_6278);
or U6584 (N_6584,N_6302,N_6310);
or U6585 (N_6585,N_6374,N_6328);
and U6586 (N_6586,N_6283,N_6496);
and U6587 (N_6587,N_6320,N_6483);
and U6588 (N_6588,N_6396,N_6344);
nor U6589 (N_6589,N_6269,N_6260);
nor U6590 (N_6590,N_6342,N_6410);
or U6591 (N_6591,N_6455,N_6492);
xnor U6592 (N_6592,N_6409,N_6312);
nor U6593 (N_6593,N_6301,N_6431);
xnor U6594 (N_6594,N_6313,N_6379);
and U6595 (N_6595,N_6445,N_6259);
nand U6596 (N_6596,N_6382,N_6337);
and U6597 (N_6597,N_6287,N_6326);
and U6598 (N_6598,N_6460,N_6338);
nand U6599 (N_6599,N_6340,N_6432);
nor U6600 (N_6600,N_6363,N_6487);
or U6601 (N_6601,N_6375,N_6419);
nor U6602 (N_6602,N_6447,N_6495);
or U6603 (N_6603,N_6250,N_6303);
or U6604 (N_6604,N_6290,N_6289);
or U6605 (N_6605,N_6479,N_6350);
nor U6606 (N_6606,N_6254,N_6426);
nor U6607 (N_6607,N_6425,N_6323);
and U6608 (N_6608,N_6417,N_6395);
and U6609 (N_6609,N_6481,N_6292);
nor U6610 (N_6610,N_6258,N_6333);
xor U6611 (N_6611,N_6422,N_6365);
xnor U6612 (N_6612,N_6380,N_6271);
nand U6613 (N_6613,N_6351,N_6280);
nor U6614 (N_6614,N_6276,N_6345);
nor U6615 (N_6615,N_6297,N_6470);
nor U6616 (N_6616,N_6489,N_6317);
and U6617 (N_6617,N_6339,N_6389);
and U6618 (N_6618,N_6359,N_6295);
or U6619 (N_6619,N_6444,N_6371);
nor U6620 (N_6620,N_6314,N_6281);
nor U6621 (N_6621,N_6256,N_6362);
or U6622 (N_6622,N_6257,N_6355);
nor U6623 (N_6623,N_6267,N_6273);
nand U6624 (N_6624,N_6352,N_6468);
or U6625 (N_6625,N_6325,N_6276);
or U6626 (N_6626,N_6386,N_6315);
xnor U6627 (N_6627,N_6493,N_6273);
and U6628 (N_6628,N_6459,N_6497);
nor U6629 (N_6629,N_6477,N_6480);
nand U6630 (N_6630,N_6383,N_6465);
nand U6631 (N_6631,N_6303,N_6493);
and U6632 (N_6632,N_6328,N_6361);
nor U6633 (N_6633,N_6380,N_6277);
nand U6634 (N_6634,N_6272,N_6275);
nor U6635 (N_6635,N_6447,N_6445);
xnor U6636 (N_6636,N_6337,N_6390);
or U6637 (N_6637,N_6336,N_6370);
nor U6638 (N_6638,N_6391,N_6363);
nand U6639 (N_6639,N_6251,N_6483);
xor U6640 (N_6640,N_6378,N_6271);
or U6641 (N_6641,N_6494,N_6462);
xnor U6642 (N_6642,N_6434,N_6452);
and U6643 (N_6643,N_6457,N_6320);
or U6644 (N_6644,N_6282,N_6476);
nor U6645 (N_6645,N_6392,N_6452);
and U6646 (N_6646,N_6456,N_6341);
xor U6647 (N_6647,N_6486,N_6374);
xor U6648 (N_6648,N_6324,N_6345);
nand U6649 (N_6649,N_6374,N_6294);
nor U6650 (N_6650,N_6439,N_6370);
nand U6651 (N_6651,N_6321,N_6369);
xnor U6652 (N_6652,N_6429,N_6371);
nor U6653 (N_6653,N_6464,N_6376);
nand U6654 (N_6654,N_6302,N_6399);
nor U6655 (N_6655,N_6258,N_6269);
nand U6656 (N_6656,N_6251,N_6366);
nor U6657 (N_6657,N_6291,N_6495);
nor U6658 (N_6658,N_6290,N_6344);
nor U6659 (N_6659,N_6370,N_6495);
nand U6660 (N_6660,N_6469,N_6251);
and U6661 (N_6661,N_6301,N_6497);
nor U6662 (N_6662,N_6454,N_6280);
xnor U6663 (N_6663,N_6443,N_6475);
or U6664 (N_6664,N_6393,N_6462);
and U6665 (N_6665,N_6468,N_6457);
xnor U6666 (N_6666,N_6371,N_6268);
nor U6667 (N_6667,N_6427,N_6258);
xnor U6668 (N_6668,N_6274,N_6344);
xnor U6669 (N_6669,N_6339,N_6401);
or U6670 (N_6670,N_6414,N_6293);
nor U6671 (N_6671,N_6253,N_6469);
and U6672 (N_6672,N_6374,N_6325);
nand U6673 (N_6673,N_6270,N_6498);
nand U6674 (N_6674,N_6325,N_6364);
nand U6675 (N_6675,N_6266,N_6396);
or U6676 (N_6676,N_6337,N_6375);
and U6677 (N_6677,N_6484,N_6263);
nor U6678 (N_6678,N_6316,N_6401);
nor U6679 (N_6679,N_6484,N_6302);
or U6680 (N_6680,N_6490,N_6335);
nand U6681 (N_6681,N_6377,N_6423);
or U6682 (N_6682,N_6344,N_6439);
nand U6683 (N_6683,N_6371,N_6297);
nand U6684 (N_6684,N_6303,N_6346);
xnor U6685 (N_6685,N_6391,N_6427);
or U6686 (N_6686,N_6253,N_6293);
nor U6687 (N_6687,N_6293,N_6299);
xnor U6688 (N_6688,N_6383,N_6400);
nand U6689 (N_6689,N_6307,N_6434);
nor U6690 (N_6690,N_6329,N_6445);
xnor U6691 (N_6691,N_6282,N_6268);
nor U6692 (N_6692,N_6488,N_6436);
xnor U6693 (N_6693,N_6461,N_6264);
or U6694 (N_6694,N_6493,N_6391);
nand U6695 (N_6695,N_6389,N_6288);
or U6696 (N_6696,N_6385,N_6386);
nand U6697 (N_6697,N_6358,N_6394);
nor U6698 (N_6698,N_6435,N_6488);
nand U6699 (N_6699,N_6473,N_6385);
and U6700 (N_6700,N_6417,N_6273);
and U6701 (N_6701,N_6405,N_6408);
or U6702 (N_6702,N_6360,N_6400);
xnor U6703 (N_6703,N_6313,N_6302);
nand U6704 (N_6704,N_6448,N_6394);
and U6705 (N_6705,N_6342,N_6451);
nand U6706 (N_6706,N_6370,N_6407);
nand U6707 (N_6707,N_6433,N_6479);
and U6708 (N_6708,N_6479,N_6450);
nor U6709 (N_6709,N_6444,N_6397);
or U6710 (N_6710,N_6274,N_6489);
nand U6711 (N_6711,N_6251,N_6451);
nand U6712 (N_6712,N_6342,N_6415);
or U6713 (N_6713,N_6470,N_6440);
or U6714 (N_6714,N_6389,N_6391);
and U6715 (N_6715,N_6382,N_6425);
or U6716 (N_6716,N_6350,N_6471);
nor U6717 (N_6717,N_6251,N_6382);
and U6718 (N_6718,N_6293,N_6365);
xnor U6719 (N_6719,N_6338,N_6305);
or U6720 (N_6720,N_6464,N_6461);
nor U6721 (N_6721,N_6372,N_6262);
nand U6722 (N_6722,N_6315,N_6307);
and U6723 (N_6723,N_6417,N_6348);
and U6724 (N_6724,N_6373,N_6478);
and U6725 (N_6725,N_6308,N_6369);
nor U6726 (N_6726,N_6475,N_6493);
nand U6727 (N_6727,N_6310,N_6345);
and U6728 (N_6728,N_6260,N_6266);
or U6729 (N_6729,N_6352,N_6420);
and U6730 (N_6730,N_6452,N_6278);
or U6731 (N_6731,N_6433,N_6289);
or U6732 (N_6732,N_6492,N_6475);
nor U6733 (N_6733,N_6489,N_6306);
nor U6734 (N_6734,N_6382,N_6343);
or U6735 (N_6735,N_6487,N_6310);
nor U6736 (N_6736,N_6449,N_6391);
and U6737 (N_6737,N_6452,N_6378);
nor U6738 (N_6738,N_6403,N_6323);
or U6739 (N_6739,N_6350,N_6468);
and U6740 (N_6740,N_6395,N_6268);
xnor U6741 (N_6741,N_6423,N_6484);
or U6742 (N_6742,N_6477,N_6305);
and U6743 (N_6743,N_6461,N_6479);
xnor U6744 (N_6744,N_6386,N_6252);
nand U6745 (N_6745,N_6419,N_6372);
or U6746 (N_6746,N_6375,N_6310);
nor U6747 (N_6747,N_6258,N_6349);
and U6748 (N_6748,N_6309,N_6440);
nor U6749 (N_6749,N_6487,N_6482);
or U6750 (N_6750,N_6618,N_6512);
or U6751 (N_6751,N_6517,N_6720);
xor U6752 (N_6752,N_6559,N_6581);
and U6753 (N_6753,N_6513,N_6729);
and U6754 (N_6754,N_6554,N_6711);
xnor U6755 (N_6755,N_6586,N_6507);
and U6756 (N_6756,N_6599,N_6632);
nor U6757 (N_6757,N_6552,N_6604);
or U6758 (N_6758,N_6545,N_6539);
nor U6759 (N_6759,N_6540,N_6743);
or U6760 (N_6760,N_6621,N_6637);
xor U6761 (N_6761,N_6629,N_6667);
nand U6762 (N_6762,N_6701,N_6610);
or U6763 (N_6763,N_6707,N_6580);
nand U6764 (N_6764,N_6665,N_6589);
or U6765 (N_6765,N_6690,N_6746);
or U6766 (N_6766,N_6567,N_6547);
and U6767 (N_6767,N_6504,N_6679);
nand U6768 (N_6768,N_6601,N_6689);
or U6769 (N_6769,N_6616,N_6646);
or U6770 (N_6770,N_6509,N_6605);
or U6771 (N_6771,N_6566,N_6570);
or U6772 (N_6772,N_6553,N_6696);
or U6773 (N_6773,N_6597,N_6732);
nor U6774 (N_6774,N_6682,N_6515);
nor U6775 (N_6775,N_6523,N_6565);
and U6776 (N_6776,N_6591,N_6587);
or U6777 (N_6777,N_6676,N_6653);
and U6778 (N_6778,N_6607,N_6651);
or U6779 (N_6779,N_6652,N_6639);
and U6780 (N_6780,N_6733,N_6630);
and U6781 (N_6781,N_6669,N_6683);
nand U6782 (N_6782,N_6698,N_6568);
nand U6783 (N_6783,N_6658,N_6631);
nand U6784 (N_6784,N_6674,N_6500);
or U6785 (N_6785,N_6520,N_6694);
and U6786 (N_6786,N_6514,N_6526);
nand U6787 (N_6787,N_6572,N_6542);
and U6788 (N_6788,N_6502,N_6728);
nor U6789 (N_6789,N_6702,N_6649);
nand U6790 (N_6790,N_6555,N_6541);
and U6791 (N_6791,N_6535,N_6548);
and U6792 (N_6792,N_6569,N_6534);
or U6793 (N_6793,N_6685,N_6739);
nor U6794 (N_6794,N_6584,N_6664);
nor U6795 (N_6795,N_6706,N_6742);
nor U6796 (N_6796,N_6609,N_6564);
nand U6797 (N_6797,N_6722,N_6666);
or U6798 (N_6798,N_6672,N_6704);
nand U6799 (N_6799,N_6735,N_6716);
nand U6800 (N_6800,N_6747,N_6655);
nor U6801 (N_6801,N_6576,N_6647);
or U6802 (N_6802,N_6582,N_6590);
or U6803 (N_6803,N_6510,N_6525);
nand U6804 (N_6804,N_6638,N_6612);
or U6805 (N_6805,N_6724,N_6537);
nand U6806 (N_6806,N_6622,N_6501);
or U6807 (N_6807,N_6546,N_6533);
nor U6808 (N_6808,N_6745,N_6709);
and U6809 (N_6809,N_6660,N_6579);
xor U6810 (N_6810,N_6519,N_6668);
nor U6811 (N_6811,N_6573,N_6532);
and U6812 (N_6812,N_6516,N_6538);
nor U6813 (N_6813,N_6644,N_6677);
or U6814 (N_6814,N_6562,N_6611);
nand U6815 (N_6815,N_6592,N_6680);
nor U6816 (N_6816,N_6661,N_6606);
and U6817 (N_6817,N_6657,N_6717);
or U6818 (N_6818,N_6634,N_6615);
and U6819 (N_6819,N_6692,N_6583);
nand U6820 (N_6820,N_6748,N_6527);
or U6821 (N_6821,N_6730,N_6563);
nand U6822 (N_6822,N_6503,N_6714);
and U6823 (N_6823,N_6725,N_6673);
and U6824 (N_6824,N_6619,N_6528);
nand U6825 (N_6825,N_6662,N_6684);
or U6826 (N_6826,N_6640,N_6712);
or U6827 (N_6827,N_6594,N_6617);
nor U6828 (N_6828,N_6595,N_6686);
nor U6829 (N_6829,N_6643,N_6633);
nand U6830 (N_6830,N_6627,N_6588);
or U6831 (N_6831,N_6671,N_6530);
nand U6832 (N_6832,N_6598,N_6575);
nor U6833 (N_6833,N_6659,N_6736);
nor U6834 (N_6834,N_6726,N_6697);
and U6835 (N_6835,N_6719,N_6635);
nand U6836 (N_6836,N_6613,N_6718);
and U6837 (N_6837,N_6585,N_6600);
and U6838 (N_6838,N_6744,N_6681);
nor U6839 (N_6839,N_6734,N_6508);
nand U6840 (N_6840,N_6678,N_6505);
or U6841 (N_6841,N_6624,N_6731);
nor U6842 (N_6842,N_6543,N_6703);
or U6843 (N_6843,N_6556,N_6710);
and U6844 (N_6844,N_6614,N_6740);
xnor U6845 (N_6845,N_6636,N_6648);
nor U6846 (N_6846,N_6511,N_6656);
xnor U6847 (N_6847,N_6691,N_6695);
and U6848 (N_6848,N_6721,N_6620);
and U6849 (N_6849,N_6593,N_6518);
or U6850 (N_6850,N_6623,N_6551);
xor U6851 (N_6851,N_6670,N_6557);
and U6852 (N_6852,N_6529,N_6650);
or U6853 (N_6853,N_6550,N_6749);
or U6854 (N_6854,N_6524,N_6642);
nand U6855 (N_6855,N_6506,N_6603);
nor U6856 (N_6856,N_6705,N_6693);
nand U6857 (N_6857,N_6708,N_6663);
xnor U6858 (N_6858,N_6561,N_6715);
or U6859 (N_6859,N_6578,N_6713);
nand U6860 (N_6860,N_6688,N_6645);
nor U6861 (N_6861,N_6521,N_6536);
and U6862 (N_6862,N_6723,N_6727);
and U6863 (N_6863,N_6571,N_6549);
nor U6864 (N_6864,N_6602,N_6641);
xor U6865 (N_6865,N_6628,N_6737);
nand U6866 (N_6866,N_6522,N_6544);
nand U6867 (N_6867,N_6531,N_6560);
or U6868 (N_6868,N_6738,N_6596);
or U6869 (N_6869,N_6699,N_6654);
or U6870 (N_6870,N_6741,N_6608);
and U6871 (N_6871,N_6625,N_6577);
and U6872 (N_6872,N_6626,N_6700);
nor U6873 (N_6873,N_6558,N_6675);
nand U6874 (N_6874,N_6687,N_6574);
or U6875 (N_6875,N_6595,N_6692);
or U6876 (N_6876,N_6617,N_6532);
nand U6877 (N_6877,N_6724,N_6584);
xor U6878 (N_6878,N_6661,N_6639);
and U6879 (N_6879,N_6564,N_6739);
nor U6880 (N_6880,N_6736,N_6511);
or U6881 (N_6881,N_6739,N_6614);
or U6882 (N_6882,N_6677,N_6522);
or U6883 (N_6883,N_6619,N_6628);
and U6884 (N_6884,N_6623,N_6728);
and U6885 (N_6885,N_6689,N_6523);
xnor U6886 (N_6886,N_6654,N_6650);
nand U6887 (N_6887,N_6725,N_6667);
and U6888 (N_6888,N_6603,N_6616);
nand U6889 (N_6889,N_6679,N_6610);
or U6890 (N_6890,N_6565,N_6653);
and U6891 (N_6891,N_6621,N_6558);
nor U6892 (N_6892,N_6708,N_6734);
nor U6893 (N_6893,N_6614,N_6662);
nand U6894 (N_6894,N_6642,N_6712);
nand U6895 (N_6895,N_6660,N_6717);
or U6896 (N_6896,N_6533,N_6508);
nor U6897 (N_6897,N_6685,N_6560);
nand U6898 (N_6898,N_6655,N_6624);
xnor U6899 (N_6899,N_6683,N_6587);
or U6900 (N_6900,N_6615,N_6663);
nor U6901 (N_6901,N_6688,N_6572);
and U6902 (N_6902,N_6745,N_6695);
nand U6903 (N_6903,N_6603,N_6744);
nand U6904 (N_6904,N_6694,N_6603);
nor U6905 (N_6905,N_6727,N_6742);
and U6906 (N_6906,N_6743,N_6577);
or U6907 (N_6907,N_6640,N_6630);
or U6908 (N_6908,N_6539,N_6657);
nand U6909 (N_6909,N_6674,N_6520);
nor U6910 (N_6910,N_6641,N_6524);
nor U6911 (N_6911,N_6727,N_6719);
nand U6912 (N_6912,N_6591,N_6718);
and U6913 (N_6913,N_6678,N_6567);
or U6914 (N_6914,N_6733,N_6557);
and U6915 (N_6915,N_6697,N_6636);
nand U6916 (N_6916,N_6591,N_6693);
and U6917 (N_6917,N_6737,N_6681);
and U6918 (N_6918,N_6732,N_6672);
nor U6919 (N_6919,N_6666,N_6623);
nor U6920 (N_6920,N_6613,N_6581);
nand U6921 (N_6921,N_6656,N_6513);
and U6922 (N_6922,N_6613,N_6640);
and U6923 (N_6923,N_6655,N_6717);
and U6924 (N_6924,N_6574,N_6675);
nand U6925 (N_6925,N_6543,N_6505);
nor U6926 (N_6926,N_6680,N_6609);
and U6927 (N_6927,N_6631,N_6536);
and U6928 (N_6928,N_6624,N_6682);
nor U6929 (N_6929,N_6559,N_6579);
and U6930 (N_6930,N_6516,N_6537);
nor U6931 (N_6931,N_6702,N_6628);
and U6932 (N_6932,N_6556,N_6684);
nand U6933 (N_6933,N_6619,N_6555);
and U6934 (N_6934,N_6541,N_6689);
nor U6935 (N_6935,N_6512,N_6541);
or U6936 (N_6936,N_6676,N_6543);
or U6937 (N_6937,N_6601,N_6518);
and U6938 (N_6938,N_6732,N_6501);
nor U6939 (N_6939,N_6643,N_6696);
and U6940 (N_6940,N_6704,N_6590);
nor U6941 (N_6941,N_6666,N_6542);
or U6942 (N_6942,N_6501,N_6519);
nand U6943 (N_6943,N_6740,N_6647);
and U6944 (N_6944,N_6668,N_6538);
nand U6945 (N_6945,N_6681,N_6721);
and U6946 (N_6946,N_6652,N_6720);
nor U6947 (N_6947,N_6624,N_6538);
or U6948 (N_6948,N_6701,N_6525);
nor U6949 (N_6949,N_6572,N_6507);
or U6950 (N_6950,N_6565,N_6728);
nand U6951 (N_6951,N_6731,N_6536);
and U6952 (N_6952,N_6743,N_6563);
nor U6953 (N_6953,N_6677,N_6527);
nor U6954 (N_6954,N_6577,N_6504);
nor U6955 (N_6955,N_6518,N_6710);
or U6956 (N_6956,N_6613,N_6661);
and U6957 (N_6957,N_6546,N_6739);
and U6958 (N_6958,N_6550,N_6647);
nand U6959 (N_6959,N_6664,N_6634);
nand U6960 (N_6960,N_6587,N_6512);
or U6961 (N_6961,N_6641,N_6715);
or U6962 (N_6962,N_6593,N_6743);
or U6963 (N_6963,N_6543,N_6723);
and U6964 (N_6964,N_6730,N_6543);
or U6965 (N_6965,N_6538,N_6524);
xnor U6966 (N_6966,N_6594,N_6626);
and U6967 (N_6967,N_6600,N_6597);
nand U6968 (N_6968,N_6678,N_6616);
or U6969 (N_6969,N_6577,N_6731);
nand U6970 (N_6970,N_6744,N_6618);
and U6971 (N_6971,N_6522,N_6501);
nor U6972 (N_6972,N_6647,N_6655);
nor U6973 (N_6973,N_6515,N_6574);
xor U6974 (N_6974,N_6554,N_6529);
xnor U6975 (N_6975,N_6714,N_6517);
xnor U6976 (N_6976,N_6731,N_6703);
or U6977 (N_6977,N_6560,N_6504);
nor U6978 (N_6978,N_6573,N_6566);
and U6979 (N_6979,N_6583,N_6539);
or U6980 (N_6980,N_6684,N_6668);
or U6981 (N_6981,N_6684,N_6694);
nor U6982 (N_6982,N_6670,N_6650);
nor U6983 (N_6983,N_6560,N_6505);
nor U6984 (N_6984,N_6636,N_6622);
or U6985 (N_6985,N_6549,N_6701);
and U6986 (N_6986,N_6591,N_6585);
nor U6987 (N_6987,N_6654,N_6618);
nand U6988 (N_6988,N_6648,N_6740);
or U6989 (N_6989,N_6561,N_6550);
and U6990 (N_6990,N_6655,N_6599);
nor U6991 (N_6991,N_6515,N_6743);
xor U6992 (N_6992,N_6644,N_6720);
and U6993 (N_6993,N_6604,N_6730);
nand U6994 (N_6994,N_6543,N_6741);
nor U6995 (N_6995,N_6517,N_6591);
nand U6996 (N_6996,N_6560,N_6515);
and U6997 (N_6997,N_6600,N_6549);
nor U6998 (N_6998,N_6704,N_6713);
nor U6999 (N_6999,N_6583,N_6582);
and U7000 (N_7000,N_6826,N_6921);
or U7001 (N_7001,N_6815,N_6855);
nand U7002 (N_7002,N_6878,N_6973);
nor U7003 (N_7003,N_6892,N_6792);
nand U7004 (N_7004,N_6947,N_6999);
nand U7005 (N_7005,N_6965,N_6964);
and U7006 (N_7006,N_6821,N_6846);
or U7007 (N_7007,N_6771,N_6995);
and U7008 (N_7008,N_6988,N_6848);
nand U7009 (N_7009,N_6939,N_6928);
nor U7010 (N_7010,N_6997,N_6959);
or U7011 (N_7011,N_6931,N_6836);
or U7012 (N_7012,N_6924,N_6969);
nand U7013 (N_7013,N_6993,N_6797);
or U7014 (N_7014,N_6856,N_6946);
nand U7015 (N_7015,N_6904,N_6934);
and U7016 (N_7016,N_6906,N_6952);
nand U7017 (N_7017,N_6767,N_6943);
and U7018 (N_7018,N_6851,N_6838);
nor U7019 (N_7019,N_6844,N_6978);
nand U7020 (N_7020,N_6834,N_6756);
or U7021 (N_7021,N_6835,N_6967);
and U7022 (N_7022,N_6827,N_6781);
and U7023 (N_7023,N_6902,N_6982);
and U7024 (N_7024,N_6789,N_6912);
and U7025 (N_7025,N_6857,N_6918);
or U7026 (N_7026,N_6891,N_6905);
nand U7027 (N_7027,N_6832,N_6841);
nor U7028 (N_7028,N_6872,N_6954);
nor U7029 (N_7029,N_6887,N_6992);
or U7030 (N_7030,N_6955,N_6784);
and U7031 (N_7031,N_6927,N_6884);
or U7032 (N_7032,N_6817,N_6914);
nor U7033 (N_7033,N_6929,N_6812);
or U7034 (N_7034,N_6800,N_6974);
or U7035 (N_7035,N_6975,N_6831);
nor U7036 (N_7036,N_6896,N_6989);
nand U7037 (N_7037,N_6942,N_6897);
or U7038 (N_7038,N_6865,N_6907);
nand U7039 (N_7039,N_6802,N_6795);
and U7040 (N_7040,N_6869,N_6875);
nor U7041 (N_7041,N_6805,N_6966);
nand U7042 (N_7042,N_6825,N_6909);
or U7043 (N_7043,N_6908,N_6977);
nand U7044 (N_7044,N_6833,N_6940);
or U7045 (N_7045,N_6783,N_6796);
and U7046 (N_7046,N_6814,N_6752);
nand U7047 (N_7047,N_6819,N_6863);
or U7048 (N_7048,N_6866,N_6903);
nand U7049 (N_7049,N_6945,N_6935);
xor U7050 (N_7050,N_6813,N_6956);
or U7051 (N_7051,N_6948,N_6976);
or U7052 (N_7052,N_6822,N_6885);
and U7053 (N_7053,N_6925,N_6782);
and U7054 (N_7054,N_6913,N_6766);
nor U7055 (N_7055,N_6890,N_6911);
nand U7056 (N_7056,N_6778,N_6861);
nand U7057 (N_7057,N_6842,N_6985);
nand U7058 (N_7058,N_6930,N_6829);
nand U7059 (N_7059,N_6895,N_6768);
or U7060 (N_7060,N_6936,N_6791);
nand U7061 (N_7061,N_6777,N_6873);
xnor U7062 (N_7062,N_6980,N_6810);
and U7063 (N_7063,N_6770,N_6759);
and U7064 (N_7064,N_6764,N_6763);
or U7065 (N_7065,N_6774,N_6760);
nor U7066 (N_7066,N_6773,N_6881);
and U7067 (N_7067,N_6779,N_6972);
or U7068 (N_7068,N_6868,N_6755);
or U7069 (N_7069,N_6910,N_6837);
and U7070 (N_7070,N_6990,N_6958);
nor U7071 (N_7071,N_6996,N_6788);
and U7072 (N_7072,N_6807,N_6970);
or U7073 (N_7073,N_6816,N_6953);
or U7074 (N_7074,N_6867,N_6849);
and U7075 (N_7075,N_6984,N_6850);
or U7076 (N_7076,N_6981,N_6762);
and U7077 (N_7077,N_6960,N_6961);
xor U7078 (N_7078,N_6858,N_6859);
or U7079 (N_7079,N_6776,N_6804);
nand U7080 (N_7080,N_6994,N_6983);
nand U7081 (N_7081,N_6801,N_6758);
nand U7082 (N_7082,N_6853,N_6951);
xor U7083 (N_7083,N_6820,N_6811);
xor U7084 (N_7084,N_6775,N_6894);
nor U7085 (N_7085,N_6920,N_6847);
xnor U7086 (N_7086,N_6932,N_6786);
nand U7087 (N_7087,N_6840,N_6798);
and U7088 (N_7088,N_6852,N_6823);
or U7089 (N_7089,N_6901,N_6769);
nor U7090 (N_7090,N_6991,N_6941);
xor U7091 (N_7091,N_6922,N_6916);
and U7092 (N_7092,N_6998,N_6862);
and U7093 (N_7093,N_6799,N_6893);
nand U7094 (N_7094,N_6919,N_6888);
nand U7095 (N_7095,N_6963,N_6818);
or U7096 (N_7096,N_6877,N_6898);
nand U7097 (N_7097,N_6882,N_6923);
and U7098 (N_7098,N_6750,N_6864);
nor U7099 (N_7099,N_6854,N_6900);
nor U7100 (N_7100,N_6794,N_6933);
and U7101 (N_7101,N_6879,N_6968);
nor U7102 (N_7102,N_6780,N_6874);
nor U7103 (N_7103,N_6839,N_6772);
and U7104 (N_7104,N_6889,N_6944);
nand U7105 (N_7105,N_6830,N_6785);
and U7106 (N_7106,N_6790,N_6886);
and U7107 (N_7107,N_6753,N_6880);
nor U7108 (N_7108,N_6824,N_6937);
and U7109 (N_7109,N_6828,N_6979);
or U7110 (N_7110,N_6803,N_6987);
xnor U7111 (N_7111,N_6917,N_6860);
or U7112 (N_7112,N_6787,N_6949);
nor U7113 (N_7113,N_6761,N_6957);
xor U7114 (N_7114,N_6870,N_6883);
or U7115 (N_7115,N_6754,N_6845);
and U7116 (N_7116,N_6899,N_6938);
and U7117 (N_7117,N_6871,N_6962);
nand U7118 (N_7118,N_6751,N_6809);
and U7119 (N_7119,N_6876,N_6793);
nand U7120 (N_7120,N_6986,N_6765);
nand U7121 (N_7121,N_6926,N_6843);
and U7122 (N_7122,N_6808,N_6915);
nor U7123 (N_7123,N_6971,N_6950);
xnor U7124 (N_7124,N_6757,N_6806);
xnor U7125 (N_7125,N_6780,N_6915);
xnor U7126 (N_7126,N_6967,N_6904);
nand U7127 (N_7127,N_6999,N_6777);
nand U7128 (N_7128,N_6765,N_6898);
or U7129 (N_7129,N_6757,N_6827);
or U7130 (N_7130,N_6810,N_6927);
and U7131 (N_7131,N_6848,N_6760);
nand U7132 (N_7132,N_6792,N_6948);
xor U7133 (N_7133,N_6901,N_6793);
or U7134 (N_7134,N_6768,N_6805);
or U7135 (N_7135,N_6864,N_6872);
nor U7136 (N_7136,N_6772,N_6840);
nand U7137 (N_7137,N_6779,N_6801);
nand U7138 (N_7138,N_6956,N_6881);
and U7139 (N_7139,N_6908,N_6882);
nor U7140 (N_7140,N_6912,N_6870);
nor U7141 (N_7141,N_6772,N_6792);
nor U7142 (N_7142,N_6957,N_6815);
and U7143 (N_7143,N_6870,N_6925);
nor U7144 (N_7144,N_6755,N_6922);
and U7145 (N_7145,N_6833,N_6904);
nand U7146 (N_7146,N_6842,N_6836);
nand U7147 (N_7147,N_6941,N_6808);
or U7148 (N_7148,N_6964,N_6881);
xor U7149 (N_7149,N_6892,N_6876);
nand U7150 (N_7150,N_6925,N_6912);
nor U7151 (N_7151,N_6999,N_6867);
xnor U7152 (N_7152,N_6812,N_6818);
nor U7153 (N_7153,N_6836,N_6979);
nor U7154 (N_7154,N_6942,N_6964);
nor U7155 (N_7155,N_6841,N_6768);
nand U7156 (N_7156,N_6883,N_6914);
and U7157 (N_7157,N_6827,N_6960);
and U7158 (N_7158,N_6871,N_6946);
or U7159 (N_7159,N_6824,N_6950);
xnor U7160 (N_7160,N_6957,N_6856);
nand U7161 (N_7161,N_6859,N_6824);
nor U7162 (N_7162,N_6861,N_6886);
and U7163 (N_7163,N_6992,N_6834);
nand U7164 (N_7164,N_6895,N_6848);
nand U7165 (N_7165,N_6804,N_6961);
xor U7166 (N_7166,N_6847,N_6807);
nor U7167 (N_7167,N_6845,N_6979);
nor U7168 (N_7168,N_6906,N_6919);
xnor U7169 (N_7169,N_6759,N_6934);
nor U7170 (N_7170,N_6766,N_6866);
nor U7171 (N_7171,N_6839,N_6766);
nor U7172 (N_7172,N_6912,N_6894);
or U7173 (N_7173,N_6891,N_6979);
nand U7174 (N_7174,N_6998,N_6976);
and U7175 (N_7175,N_6954,N_6859);
and U7176 (N_7176,N_6949,N_6975);
or U7177 (N_7177,N_6806,N_6755);
and U7178 (N_7178,N_6887,N_6763);
or U7179 (N_7179,N_6915,N_6999);
or U7180 (N_7180,N_6970,N_6759);
or U7181 (N_7181,N_6952,N_6842);
nand U7182 (N_7182,N_6757,N_6860);
xor U7183 (N_7183,N_6997,N_6961);
xor U7184 (N_7184,N_6922,N_6765);
nand U7185 (N_7185,N_6838,N_6895);
nor U7186 (N_7186,N_6798,N_6893);
and U7187 (N_7187,N_6996,N_6836);
xor U7188 (N_7188,N_6880,N_6810);
or U7189 (N_7189,N_6953,N_6915);
or U7190 (N_7190,N_6861,N_6902);
or U7191 (N_7191,N_6827,N_6969);
or U7192 (N_7192,N_6776,N_6891);
and U7193 (N_7193,N_6829,N_6796);
nor U7194 (N_7194,N_6891,N_6947);
and U7195 (N_7195,N_6864,N_6768);
nand U7196 (N_7196,N_6819,N_6938);
nand U7197 (N_7197,N_6972,N_6950);
or U7198 (N_7198,N_6947,N_6778);
and U7199 (N_7199,N_6808,N_6885);
xor U7200 (N_7200,N_6928,N_6844);
nand U7201 (N_7201,N_6763,N_6966);
nor U7202 (N_7202,N_6764,N_6875);
xor U7203 (N_7203,N_6759,N_6884);
nand U7204 (N_7204,N_6879,N_6897);
or U7205 (N_7205,N_6794,N_6800);
or U7206 (N_7206,N_6753,N_6845);
and U7207 (N_7207,N_6752,N_6866);
nor U7208 (N_7208,N_6847,N_6840);
xor U7209 (N_7209,N_6784,N_6964);
nand U7210 (N_7210,N_6964,N_6751);
or U7211 (N_7211,N_6813,N_6865);
or U7212 (N_7212,N_6812,N_6750);
xnor U7213 (N_7213,N_6751,N_6784);
nand U7214 (N_7214,N_6810,N_6940);
and U7215 (N_7215,N_6826,N_6831);
and U7216 (N_7216,N_6870,N_6798);
and U7217 (N_7217,N_6753,N_6971);
nand U7218 (N_7218,N_6882,N_6779);
nor U7219 (N_7219,N_6996,N_6887);
or U7220 (N_7220,N_6762,N_6801);
nor U7221 (N_7221,N_6937,N_6883);
xnor U7222 (N_7222,N_6990,N_6899);
xor U7223 (N_7223,N_6986,N_6839);
nand U7224 (N_7224,N_6857,N_6760);
or U7225 (N_7225,N_6833,N_6819);
nor U7226 (N_7226,N_6753,N_6893);
or U7227 (N_7227,N_6842,N_6803);
nand U7228 (N_7228,N_6883,N_6809);
or U7229 (N_7229,N_6791,N_6810);
nor U7230 (N_7230,N_6786,N_6841);
or U7231 (N_7231,N_6788,N_6867);
nor U7232 (N_7232,N_6972,N_6831);
or U7233 (N_7233,N_6865,N_6926);
nor U7234 (N_7234,N_6876,N_6851);
or U7235 (N_7235,N_6812,N_6767);
nor U7236 (N_7236,N_6856,N_6827);
nand U7237 (N_7237,N_6908,N_6796);
nor U7238 (N_7238,N_6919,N_6946);
or U7239 (N_7239,N_6929,N_6961);
and U7240 (N_7240,N_6961,N_6949);
and U7241 (N_7241,N_6941,N_6956);
nor U7242 (N_7242,N_6802,N_6878);
or U7243 (N_7243,N_6989,N_6881);
nand U7244 (N_7244,N_6852,N_6787);
nor U7245 (N_7245,N_6885,N_6930);
or U7246 (N_7246,N_6878,N_6824);
or U7247 (N_7247,N_6829,N_6818);
nor U7248 (N_7248,N_6780,N_6909);
nand U7249 (N_7249,N_6837,N_6883);
and U7250 (N_7250,N_7194,N_7152);
nor U7251 (N_7251,N_7093,N_7209);
nor U7252 (N_7252,N_7095,N_7235);
nor U7253 (N_7253,N_7021,N_7188);
and U7254 (N_7254,N_7006,N_7217);
nand U7255 (N_7255,N_7125,N_7054);
and U7256 (N_7256,N_7077,N_7058);
or U7257 (N_7257,N_7110,N_7202);
and U7258 (N_7258,N_7249,N_7090);
nand U7259 (N_7259,N_7035,N_7016);
and U7260 (N_7260,N_7086,N_7190);
or U7261 (N_7261,N_7225,N_7172);
and U7262 (N_7262,N_7153,N_7040);
xnor U7263 (N_7263,N_7206,N_7178);
or U7264 (N_7264,N_7003,N_7230);
and U7265 (N_7265,N_7109,N_7124);
nand U7266 (N_7266,N_7134,N_7213);
and U7267 (N_7267,N_7002,N_7037);
and U7268 (N_7268,N_7214,N_7234);
or U7269 (N_7269,N_7221,N_7210);
nand U7270 (N_7270,N_7026,N_7047);
or U7271 (N_7271,N_7068,N_7032);
or U7272 (N_7272,N_7157,N_7119);
nor U7273 (N_7273,N_7145,N_7014);
and U7274 (N_7274,N_7105,N_7085);
nand U7275 (N_7275,N_7089,N_7091);
or U7276 (N_7276,N_7144,N_7177);
or U7277 (N_7277,N_7075,N_7101);
nor U7278 (N_7278,N_7150,N_7163);
or U7279 (N_7279,N_7175,N_7098);
or U7280 (N_7280,N_7142,N_7132);
and U7281 (N_7281,N_7232,N_7061);
nand U7282 (N_7282,N_7166,N_7120);
and U7283 (N_7283,N_7147,N_7201);
nor U7284 (N_7284,N_7080,N_7216);
or U7285 (N_7285,N_7176,N_7103);
or U7286 (N_7286,N_7180,N_7231);
or U7287 (N_7287,N_7036,N_7123);
and U7288 (N_7288,N_7169,N_7004);
nand U7289 (N_7289,N_7156,N_7115);
and U7290 (N_7290,N_7233,N_7242);
or U7291 (N_7291,N_7070,N_7087);
and U7292 (N_7292,N_7174,N_7126);
nand U7293 (N_7293,N_7154,N_7107);
nor U7294 (N_7294,N_7240,N_7059);
nand U7295 (N_7295,N_7139,N_7034);
and U7296 (N_7296,N_7155,N_7094);
xor U7297 (N_7297,N_7027,N_7069);
nor U7298 (N_7298,N_7076,N_7010);
or U7299 (N_7299,N_7192,N_7072);
nand U7300 (N_7300,N_7013,N_7168);
nand U7301 (N_7301,N_7025,N_7161);
xnor U7302 (N_7302,N_7195,N_7066);
xor U7303 (N_7303,N_7019,N_7171);
nor U7304 (N_7304,N_7020,N_7011);
or U7305 (N_7305,N_7030,N_7204);
and U7306 (N_7306,N_7099,N_7131);
and U7307 (N_7307,N_7050,N_7022);
nor U7308 (N_7308,N_7081,N_7096);
and U7309 (N_7309,N_7084,N_7159);
nand U7310 (N_7310,N_7043,N_7015);
and U7311 (N_7311,N_7128,N_7029);
nand U7312 (N_7312,N_7111,N_7223);
and U7313 (N_7313,N_7246,N_7009);
or U7314 (N_7314,N_7062,N_7113);
or U7315 (N_7315,N_7205,N_7116);
nand U7316 (N_7316,N_7173,N_7042);
or U7317 (N_7317,N_7181,N_7044);
or U7318 (N_7318,N_7057,N_7189);
and U7319 (N_7319,N_7247,N_7212);
nand U7320 (N_7320,N_7237,N_7148);
and U7321 (N_7321,N_7164,N_7102);
or U7322 (N_7322,N_7211,N_7135);
nor U7323 (N_7323,N_7244,N_7196);
nand U7324 (N_7324,N_7063,N_7220);
nand U7325 (N_7325,N_7039,N_7067);
nor U7326 (N_7326,N_7187,N_7088);
nor U7327 (N_7327,N_7141,N_7114);
and U7328 (N_7328,N_7207,N_7053);
nand U7329 (N_7329,N_7127,N_7208);
xor U7330 (N_7330,N_7143,N_7200);
and U7331 (N_7331,N_7136,N_7198);
nand U7332 (N_7332,N_7106,N_7118);
or U7333 (N_7333,N_7218,N_7241);
and U7334 (N_7334,N_7001,N_7033);
and U7335 (N_7335,N_7100,N_7012);
and U7336 (N_7336,N_7104,N_7023);
nand U7337 (N_7337,N_7183,N_7005);
and U7338 (N_7338,N_7065,N_7162);
nand U7339 (N_7339,N_7193,N_7024);
and U7340 (N_7340,N_7078,N_7028);
nor U7341 (N_7341,N_7222,N_7165);
xnor U7342 (N_7342,N_7236,N_7170);
xnor U7343 (N_7343,N_7122,N_7179);
and U7344 (N_7344,N_7046,N_7137);
nor U7345 (N_7345,N_7041,N_7248);
or U7346 (N_7346,N_7184,N_7229);
and U7347 (N_7347,N_7160,N_7018);
or U7348 (N_7348,N_7064,N_7227);
nand U7349 (N_7349,N_7243,N_7060);
nand U7350 (N_7350,N_7224,N_7239);
nand U7351 (N_7351,N_7238,N_7138);
nor U7352 (N_7352,N_7197,N_7112);
nand U7353 (N_7353,N_7133,N_7051);
nor U7354 (N_7354,N_7049,N_7052);
nor U7355 (N_7355,N_7117,N_7056);
xnor U7356 (N_7356,N_7199,N_7121);
nor U7357 (N_7357,N_7130,N_7219);
nand U7358 (N_7358,N_7203,N_7045);
nor U7359 (N_7359,N_7228,N_7071);
or U7360 (N_7360,N_7007,N_7031);
nor U7361 (N_7361,N_7092,N_7017);
nor U7362 (N_7362,N_7083,N_7008);
nor U7363 (N_7363,N_7082,N_7186);
and U7364 (N_7364,N_7000,N_7185);
nand U7365 (N_7365,N_7140,N_7108);
and U7366 (N_7366,N_7245,N_7151);
nand U7367 (N_7367,N_7167,N_7074);
xnor U7368 (N_7368,N_7226,N_7048);
nor U7369 (N_7369,N_7038,N_7073);
or U7370 (N_7370,N_7158,N_7055);
and U7371 (N_7371,N_7191,N_7097);
xnor U7372 (N_7372,N_7182,N_7149);
nand U7373 (N_7373,N_7215,N_7129);
nand U7374 (N_7374,N_7079,N_7146);
nor U7375 (N_7375,N_7030,N_7225);
nand U7376 (N_7376,N_7149,N_7133);
nand U7377 (N_7377,N_7089,N_7160);
nor U7378 (N_7378,N_7150,N_7047);
or U7379 (N_7379,N_7057,N_7022);
and U7380 (N_7380,N_7136,N_7055);
nand U7381 (N_7381,N_7158,N_7137);
nand U7382 (N_7382,N_7144,N_7141);
xor U7383 (N_7383,N_7024,N_7124);
or U7384 (N_7384,N_7249,N_7035);
or U7385 (N_7385,N_7082,N_7124);
or U7386 (N_7386,N_7155,N_7093);
nor U7387 (N_7387,N_7130,N_7041);
nand U7388 (N_7388,N_7070,N_7246);
nand U7389 (N_7389,N_7085,N_7123);
and U7390 (N_7390,N_7226,N_7093);
and U7391 (N_7391,N_7195,N_7181);
nand U7392 (N_7392,N_7170,N_7140);
nand U7393 (N_7393,N_7234,N_7142);
nor U7394 (N_7394,N_7089,N_7138);
or U7395 (N_7395,N_7031,N_7184);
nor U7396 (N_7396,N_7150,N_7074);
nand U7397 (N_7397,N_7008,N_7198);
nand U7398 (N_7398,N_7075,N_7038);
and U7399 (N_7399,N_7056,N_7165);
nand U7400 (N_7400,N_7089,N_7203);
and U7401 (N_7401,N_7012,N_7052);
or U7402 (N_7402,N_7065,N_7078);
or U7403 (N_7403,N_7153,N_7193);
and U7404 (N_7404,N_7031,N_7157);
xor U7405 (N_7405,N_7012,N_7074);
and U7406 (N_7406,N_7187,N_7201);
and U7407 (N_7407,N_7062,N_7048);
xnor U7408 (N_7408,N_7134,N_7029);
nand U7409 (N_7409,N_7167,N_7171);
and U7410 (N_7410,N_7177,N_7066);
nand U7411 (N_7411,N_7036,N_7194);
or U7412 (N_7412,N_7090,N_7202);
nand U7413 (N_7413,N_7214,N_7156);
nor U7414 (N_7414,N_7215,N_7007);
nand U7415 (N_7415,N_7006,N_7236);
and U7416 (N_7416,N_7048,N_7010);
nand U7417 (N_7417,N_7008,N_7088);
nor U7418 (N_7418,N_7122,N_7075);
nor U7419 (N_7419,N_7204,N_7081);
nand U7420 (N_7420,N_7105,N_7057);
xor U7421 (N_7421,N_7038,N_7165);
and U7422 (N_7422,N_7038,N_7140);
and U7423 (N_7423,N_7162,N_7082);
and U7424 (N_7424,N_7032,N_7176);
or U7425 (N_7425,N_7020,N_7115);
xnor U7426 (N_7426,N_7122,N_7015);
nor U7427 (N_7427,N_7144,N_7159);
and U7428 (N_7428,N_7016,N_7041);
nand U7429 (N_7429,N_7030,N_7012);
nor U7430 (N_7430,N_7201,N_7222);
and U7431 (N_7431,N_7202,N_7061);
nor U7432 (N_7432,N_7039,N_7164);
nor U7433 (N_7433,N_7008,N_7070);
nand U7434 (N_7434,N_7110,N_7017);
nand U7435 (N_7435,N_7198,N_7201);
nor U7436 (N_7436,N_7224,N_7170);
nor U7437 (N_7437,N_7060,N_7122);
or U7438 (N_7438,N_7154,N_7062);
nor U7439 (N_7439,N_7190,N_7197);
nor U7440 (N_7440,N_7110,N_7249);
nand U7441 (N_7441,N_7239,N_7036);
or U7442 (N_7442,N_7038,N_7021);
nor U7443 (N_7443,N_7221,N_7017);
or U7444 (N_7444,N_7210,N_7242);
nand U7445 (N_7445,N_7221,N_7106);
nor U7446 (N_7446,N_7192,N_7169);
nand U7447 (N_7447,N_7181,N_7108);
nand U7448 (N_7448,N_7055,N_7191);
nor U7449 (N_7449,N_7142,N_7194);
or U7450 (N_7450,N_7174,N_7224);
nand U7451 (N_7451,N_7223,N_7027);
nor U7452 (N_7452,N_7198,N_7042);
or U7453 (N_7453,N_7156,N_7129);
and U7454 (N_7454,N_7140,N_7200);
nor U7455 (N_7455,N_7186,N_7188);
or U7456 (N_7456,N_7037,N_7134);
nand U7457 (N_7457,N_7169,N_7076);
and U7458 (N_7458,N_7184,N_7124);
nand U7459 (N_7459,N_7148,N_7041);
nor U7460 (N_7460,N_7061,N_7167);
nor U7461 (N_7461,N_7153,N_7056);
nand U7462 (N_7462,N_7238,N_7239);
nand U7463 (N_7463,N_7087,N_7084);
nand U7464 (N_7464,N_7077,N_7137);
xor U7465 (N_7465,N_7031,N_7205);
or U7466 (N_7466,N_7025,N_7227);
nand U7467 (N_7467,N_7093,N_7048);
nor U7468 (N_7468,N_7202,N_7063);
nand U7469 (N_7469,N_7018,N_7158);
nor U7470 (N_7470,N_7103,N_7175);
nand U7471 (N_7471,N_7177,N_7160);
or U7472 (N_7472,N_7221,N_7014);
nand U7473 (N_7473,N_7236,N_7068);
or U7474 (N_7474,N_7101,N_7146);
nor U7475 (N_7475,N_7144,N_7216);
or U7476 (N_7476,N_7060,N_7005);
xor U7477 (N_7477,N_7223,N_7188);
xnor U7478 (N_7478,N_7155,N_7193);
and U7479 (N_7479,N_7118,N_7195);
and U7480 (N_7480,N_7031,N_7169);
or U7481 (N_7481,N_7192,N_7139);
nor U7482 (N_7482,N_7013,N_7041);
nand U7483 (N_7483,N_7013,N_7137);
nor U7484 (N_7484,N_7166,N_7058);
nand U7485 (N_7485,N_7004,N_7184);
nor U7486 (N_7486,N_7181,N_7192);
nand U7487 (N_7487,N_7014,N_7061);
nor U7488 (N_7488,N_7040,N_7177);
and U7489 (N_7489,N_7191,N_7098);
nand U7490 (N_7490,N_7004,N_7187);
nor U7491 (N_7491,N_7112,N_7052);
nor U7492 (N_7492,N_7032,N_7018);
nor U7493 (N_7493,N_7075,N_7032);
or U7494 (N_7494,N_7081,N_7135);
nand U7495 (N_7495,N_7096,N_7181);
nand U7496 (N_7496,N_7110,N_7085);
nor U7497 (N_7497,N_7034,N_7209);
or U7498 (N_7498,N_7030,N_7071);
nand U7499 (N_7499,N_7247,N_7095);
nor U7500 (N_7500,N_7264,N_7312);
nand U7501 (N_7501,N_7339,N_7322);
nand U7502 (N_7502,N_7392,N_7408);
and U7503 (N_7503,N_7304,N_7474);
or U7504 (N_7504,N_7395,N_7337);
nor U7505 (N_7505,N_7252,N_7356);
nor U7506 (N_7506,N_7327,N_7288);
nand U7507 (N_7507,N_7325,N_7467);
or U7508 (N_7508,N_7274,N_7295);
and U7509 (N_7509,N_7420,N_7409);
xor U7510 (N_7510,N_7482,N_7316);
and U7511 (N_7511,N_7499,N_7340);
nor U7512 (N_7512,N_7478,N_7367);
and U7513 (N_7513,N_7493,N_7463);
nor U7514 (N_7514,N_7353,N_7390);
or U7515 (N_7515,N_7426,N_7419);
or U7516 (N_7516,N_7459,N_7328);
nand U7517 (N_7517,N_7451,N_7351);
or U7518 (N_7518,N_7399,N_7434);
and U7519 (N_7519,N_7344,N_7260);
nor U7520 (N_7520,N_7365,N_7330);
nor U7521 (N_7521,N_7277,N_7314);
and U7522 (N_7522,N_7379,N_7446);
or U7523 (N_7523,N_7321,N_7303);
and U7524 (N_7524,N_7291,N_7455);
nand U7525 (N_7525,N_7435,N_7282);
and U7526 (N_7526,N_7380,N_7452);
nor U7527 (N_7527,N_7266,N_7471);
or U7528 (N_7528,N_7403,N_7355);
nand U7529 (N_7529,N_7432,N_7374);
or U7530 (N_7530,N_7453,N_7410);
and U7531 (N_7531,N_7338,N_7342);
nand U7532 (N_7532,N_7425,N_7414);
and U7533 (N_7533,N_7270,N_7491);
nand U7534 (N_7534,N_7498,N_7402);
nor U7535 (N_7535,N_7472,N_7269);
nand U7536 (N_7536,N_7258,N_7318);
or U7537 (N_7537,N_7464,N_7494);
or U7538 (N_7538,N_7400,N_7406);
and U7539 (N_7539,N_7440,N_7438);
nand U7540 (N_7540,N_7369,N_7299);
or U7541 (N_7541,N_7412,N_7313);
xnor U7542 (N_7542,N_7481,N_7263);
or U7543 (N_7543,N_7335,N_7450);
or U7544 (N_7544,N_7462,N_7473);
nor U7545 (N_7545,N_7305,N_7372);
and U7546 (N_7546,N_7255,N_7376);
and U7547 (N_7547,N_7490,N_7417);
nor U7548 (N_7548,N_7306,N_7273);
and U7549 (N_7549,N_7259,N_7430);
nor U7550 (N_7550,N_7495,N_7407);
or U7551 (N_7551,N_7416,N_7293);
nor U7552 (N_7552,N_7307,N_7466);
nand U7553 (N_7553,N_7480,N_7289);
or U7554 (N_7554,N_7354,N_7284);
and U7555 (N_7555,N_7411,N_7324);
nor U7556 (N_7556,N_7447,N_7253);
nand U7557 (N_7557,N_7294,N_7265);
or U7558 (N_7558,N_7309,N_7429);
nand U7559 (N_7559,N_7456,N_7320);
and U7560 (N_7560,N_7468,N_7326);
xor U7561 (N_7561,N_7345,N_7271);
or U7562 (N_7562,N_7397,N_7415);
nor U7563 (N_7563,N_7413,N_7443);
xnor U7564 (N_7564,N_7377,N_7332);
or U7565 (N_7565,N_7348,N_7254);
nor U7566 (N_7566,N_7476,N_7445);
or U7567 (N_7567,N_7475,N_7334);
and U7568 (N_7568,N_7387,N_7457);
or U7569 (N_7569,N_7371,N_7444);
nor U7570 (N_7570,N_7378,N_7331);
or U7571 (N_7571,N_7404,N_7461);
nor U7572 (N_7572,N_7276,N_7267);
nand U7573 (N_7573,N_7319,N_7391);
or U7574 (N_7574,N_7479,N_7427);
xor U7575 (N_7575,N_7477,N_7347);
and U7576 (N_7576,N_7424,N_7496);
and U7577 (N_7577,N_7442,N_7405);
nand U7578 (N_7578,N_7317,N_7300);
nor U7579 (N_7579,N_7280,N_7439);
and U7580 (N_7580,N_7261,N_7394);
xnor U7581 (N_7581,N_7336,N_7302);
or U7582 (N_7582,N_7448,N_7352);
nand U7583 (N_7583,N_7349,N_7292);
xnor U7584 (N_7584,N_7279,N_7283);
nor U7585 (N_7585,N_7418,N_7308);
and U7586 (N_7586,N_7396,N_7441);
nand U7587 (N_7587,N_7398,N_7290);
and U7588 (N_7588,N_7373,N_7384);
nor U7589 (N_7589,N_7484,N_7454);
nor U7590 (N_7590,N_7423,N_7485);
and U7591 (N_7591,N_7486,N_7470);
nor U7592 (N_7592,N_7436,N_7382);
or U7593 (N_7593,N_7311,N_7431);
nor U7594 (N_7594,N_7361,N_7257);
xnor U7595 (N_7595,N_7362,N_7323);
and U7596 (N_7596,N_7278,N_7393);
nand U7597 (N_7597,N_7341,N_7256);
and U7598 (N_7598,N_7250,N_7268);
xnor U7599 (N_7599,N_7437,N_7497);
nor U7600 (N_7600,N_7389,N_7489);
or U7601 (N_7601,N_7286,N_7488);
and U7602 (N_7602,N_7433,N_7383);
nand U7603 (N_7603,N_7375,N_7492);
xnor U7604 (N_7604,N_7329,N_7366);
or U7605 (N_7605,N_7458,N_7298);
nor U7606 (N_7606,N_7460,N_7333);
and U7607 (N_7607,N_7469,N_7449);
nor U7608 (N_7608,N_7357,N_7386);
or U7609 (N_7609,N_7297,N_7285);
nand U7610 (N_7610,N_7310,N_7381);
xor U7611 (N_7611,N_7421,N_7422);
nor U7612 (N_7612,N_7281,N_7296);
xnor U7613 (N_7613,N_7363,N_7487);
or U7614 (N_7614,N_7272,N_7388);
xor U7615 (N_7615,N_7343,N_7360);
or U7616 (N_7616,N_7465,N_7364);
or U7617 (N_7617,N_7483,N_7262);
nor U7618 (N_7618,N_7428,N_7385);
nor U7619 (N_7619,N_7287,N_7275);
nand U7620 (N_7620,N_7301,N_7370);
and U7621 (N_7621,N_7401,N_7251);
and U7622 (N_7622,N_7359,N_7350);
nor U7623 (N_7623,N_7346,N_7368);
xnor U7624 (N_7624,N_7315,N_7358);
or U7625 (N_7625,N_7356,N_7496);
nor U7626 (N_7626,N_7489,N_7265);
nor U7627 (N_7627,N_7377,N_7266);
nor U7628 (N_7628,N_7493,N_7484);
and U7629 (N_7629,N_7289,N_7262);
and U7630 (N_7630,N_7363,N_7456);
or U7631 (N_7631,N_7449,N_7250);
nand U7632 (N_7632,N_7459,N_7472);
or U7633 (N_7633,N_7469,N_7306);
nand U7634 (N_7634,N_7369,N_7388);
and U7635 (N_7635,N_7425,N_7284);
nor U7636 (N_7636,N_7497,N_7280);
and U7637 (N_7637,N_7484,N_7359);
and U7638 (N_7638,N_7468,N_7287);
xnor U7639 (N_7639,N_7256,N_7459);
or U7640 (N_7640,N_7464,N_7252);
nand U7641 (N_7641,N_7434,N_7323);
nand U7642 (N_7642,N_7335,N_7262);
nor U7643 (N_7643,N_7269,N_7382);
nor U7644 (N_7644,N_7411,N_7401);
nor U7645 (N_7645,N_7482,N_7278);
nor U7646 (N_7646,N_7450,N_7314);
and U7647 (N_7647,N_7253,N_7398);
nor U7648 (N_7648,N_7468,N_7465);
xnor U7649 (N_7649,N_7269,N_7475);
nor U7650 (N_7650,N_7359,N_7499);
and U7651 (N_7651,N_7405,N_7433);
and U7652 (N_7652,N_7256,N_7458);
or U7653 (N_7653,N_7288,N_7490);
and U7654 (N_7654,N_7419,N_7433);
nand U7655 (N_7655,N_7366,N_7486);
or U7656 (N_7656,N_7469,N_7321);
nand U7657 (N_7657,N_7384,N_7369);
and U7658 (N_7658,N_7332,N_7330);
and U7659 (N_7659,N_7313,N_7393);
nand U7660 (N_7660,N_7434,N_7360);
and U7661 (N_7661,N_7377,N_7264);
and U7662 (N_7662,N_7383,N_7461);
nor U7663 (N_7663,N_7279,N_7388);
xnor U7664 (N_7664,N_7481,N_7402);
and U7665 (N_7665,N_7375,N_7387);
or U7666 (N_7666,N_7280,N_7481);
or U7667 (N_7667,N_7433,N_7481);
nor U7668 (N_7668,N_7337,N_7371);
nor U7669 (N_7669,N_7416,N_7478);
nand U7670 (N_7670,N_7355,N_7379);
nor U7671 (N_7671,N_7360,N_7288);
nor U7672 (N_7672,N_7447,N_7285);
nand U7673 (N_7673,N_7447,N_7495);
nand U7674 (N_7674,N_7336,N_7410);
nand U7675 (N_7675,N_7324,N_7480);
or U7676 (N_7676,N_7366,N_7260);
or U7677 (N_7677,N_7344,N_7379);
and U7678 (N_7678,N_7425,N_7370);
or U7679 (N_7679,N_7359,N_7377);
and U7680 (N_7680,N_7304,N_7434);
nor U7681 (N_7681,N_7499,N_7429);
and U7682 (N_7682,N_7341,N_7314);
or U7683 (N_7683,N_7385,N_7261);
or U7684 (N_7684,N_7466,N_7301);
and U7685 (N_7685,N_7348,N_7415);
or U7686 (N_7686,N_7339,N_7279);
and U7687 (N_7687,N_7317,N_7388);
nor U7688 (N_7688,N_7250,N_7475);
nand U7689 (N_7689,N_7375,N_7294);
and U7690 (N_7690,N_7255,N_7374);
nor U7691 (N_7691,N_7353,N_7444);
nand U7692 (N_7692,N_7371,N_7493);
nand U7693 (N_7693,N_7399,N_7431);
nand U7694 (N_7694,N_7410,N_7421);
and U7695 (N_7695,N_7499,N_7462);
and U7696 (N_7696,N_7488,N_7313);
nor U7697 (N_7697,N_7328,N_7312);
nand U7698 (N_7698,N_7296,N_7496);
and U7699 (N_7699,N_7379,N_7478);
and U7700 (N_7700,N_7260,N_7404);
nand U7701 (N_7701,N_7498,N_7384);
and U7702 (N_7702,N_7379,N_7466);
nor U7703 (N_7703,N_7330,N_7391);
nand U7704 (N_7704,N_7286,N_7492);
or U7705 (N_7705,N_7451,N_7324);
and U7706 (N_7706,N_7387,N_7263);
and U7707 (N_7707,N_7256,N_7331);
nand U7708 (N_7708,N_7458,N_7337);
nor U7709 (N_7709,N_7427,N_7281);
or U7710 (N_7710,N_7326,N_7345);
nor U7711 (N_7711,N_7397,N_7451);
or U7712 (N_7712,N_7290,N_7484);
nor U7713 (N_7713,N_7318,N_7418);
or U7714 (N_7714,N_7417,N_7333);
nand U7715 (N_7715,N_7329,N_7325);
nor U7716 (N_7716,N_7413,N_7482);
nor U7717 (N_7717,N_7264,N_7378);
nor U7718 (N_7718,N_7484,N_7388);
and U7719 (N_7719,N_7475,N_7414);
or U7720 (N_7720,N_7277,N_7258);
or U7721 (N_7721,N_7416,N_7336);
nand U7722 (N_7722,N_7301,N_7363);
or U7723 (N_7723,N_7476,N_7375);
nor U7724 (N_7724,N_7252,N_7408);
xor U7725 (N_7725,N_7499,N_7294);
nor U7726 (N_7726,N_7285,N_7282);
or U7727 (N_7727,N_7495,N_7318);
nor U7728 (N_7728,N_7326,N_7431);
and U7729 (N_7729,N_7277,N_7469);
and U7730 (N_7730,N_7403,N_7289);
nor U7731 (N_7731,N_7257,N_7335);
nand U7732 (N_7732,N_7453,N_7497);
or U7733 (N_7733,N_7311,N_7318);
nor U7734 (N_7734,N_7478,N_7372);
and U7735 (N_7735,N_7299,N_7457);
and U7736 (N_7736,N_7255,N_7451);
and U7737 (N_7737,N_7453,N_7331);
nor U7738 (N_7738,N_7326,N_7410);
and U7739 (N_7739,N_7320,N_7446);
or U7740 (N_7740,N_7316,N_7330);
or U7741 (N_7741,N_7381,N_7430);
or U7742 (N_7742,N_7457,N_7490);
nor U7743 (N_7743,N_7255,N_7314);
nand U7744 (N_7744,N_7427,N_7409);
nor U7745 (N_7745,N_7429,N_7350);
or U7746 (N_7746,N_7469,N_7447);
nor U7747 (N_7747,N_7276,N_7319);
nand U7748 (N_7748,N_7254,N_7363);
nor U7749 (N_7749,N_7497,N_7458);
xor U7750 (N_7750,N_7594,N_7688);
or U7751 (N_7751,N_7698,N_7505);
and U7752 (N_7752,N_7684,N_7508);
or U7753 (N_7753,N_7607,N_7747);
nor U7754 (N_7754,N_7545,N_7740);
nor U7755 (N_7755,N_7660,N_7673);
and U7756 (N_7756,N_7531,N_7520);
xor U7757 (N_7757,N_7669,N_7577);
or U7758 (N_7758,N_7693,N_7552);
nand U7759 (N_7759,N_7540,N_7565);
nand U7760 (N_7760,N_7676,N_7674);
or U7761 (N_7761,N_7600,N_7610);
nor U7762 (N_7762,N_7644,N_7548);
nand U7763 (N_7763,N_7665,N_7662);
nand U7764 (N_7764,N_7609,N_7556);
nor U7765 (N_7765,N_7561,N_7538);
or U7766 (N_7766,N_7687,N_7584);
nor U7767 (N_7767,N_7575,N_7746);
nand U7768 (N_7768,N_7624,N_7566);
and U7769 (N_7769,N_7646,N_7569);
and U7770 (N_7770,N_7586,N_7555);
or U7771 (N_7771,N_7721,N_7722);
nand U7772 (N_7772,N_7703,N_7554);
or U7773 (N_7773,N_7679,N_7745);
and U7774 (N_7774,N_7710,N_7590);
nand U7775 (N_7775,N_7602,N_7510);
and U7776 (N_7776,N_7603,N_7578);
nand U7777 (N_7777,N_7534,N_7516);
and U7778 (N_7778,N_7638,N_7513);
nor U7779 (N_7779,N_7705,N_7654);
and U7780 (N_7780,N_7535,N_7635);
or U7781 (N_7781,N_7546,N_7637);
and U7782 (N_7782,N_7592,N_7567);
xnor U7783 (N_7783,N_7648,N_7649);
or U7784 (N_7784,N_7570,N_7620);
and U7785 (N_7785,N_7668,N_7736);
nor U7786 (N_7786,N_7670,N_7606);
and U7787 (N_7787,N_7541,N_7542);
and U7788 (N_7788,N_7621,N_7580);
or U7789 (N_7789,N_7625,N_7595);
or U7790 (N_7790,N_7686,N_7514);
nor U7791 (N_7791,N_7737,N_7656);
nor U7792 (N_7792,N_7587,N_7573);
nand U7793 (N_7793,N_7604,N_7616);
and U7794 (N_7794,N_7618,N_7739);
nor U7795 (N_7795,N_7658,N_7591);
and U7796 (N_7796,N_7553,N_7713);
xnor U7797 (N_7797,N_7536,N_7731);
nor U7798 (N_7798,N_7559,N_7568);
nor U7799 (N_7799,N_7666,N_7675);
and U7800 (N_7800,N_7558,N_7551);
nor U7801 (N_7801,N_7633,N_7515);
or U7802 (N_7802,N_7533,N_7527);
or U7803 (N_7803,N_7589,N_7564);
and U7804 (N_7804,N_7506,N_7547);
nand U7805 (N_7805,N_7702,N_7652);
nand U7806 (N_7806,N_7598,N_7504);
nand U7807 (N_7807,N_7704,N_7639);
nor U7808 (N_7808,N_7733,N_7730);
or U7809 (N_7809,N_7507,N_7729);
nor U7810 (N_7810,N_7735,N_7683);
and U7811 (N_7811,N_7611,N_7585);
xnor U7812 (N_7812,N_7700,N_7734);
nand U7813 (N_7813,N_7711,N_7509);
nand U7814 (N_7814,N_7550,N_7629);
or U7815 (N_7815,N_7664,N_7701);
nand U7816 (N_7816,N_7615,N_7579);
and U7817 (N_7817,N_7605,N_7628);
and U7818 (N_7818,N_7715,N_7574);
nand U7819 (N_7819,N_7719,N_7503);
or U7820 (N_7820,N_7582,N_7697);
and U7821 (N_7821,N_7692,N_7712);
nor U7822 (N_7822,N_7716,N_7691);
nand U7823 (N_7823,N_7522,N_7651);
nor U7824 (N_7824,N_7653,N_7742);
and U7825 (N_7825,N_7709,N_7521);
nor U7826 (N_7826,N_7523,N_7690);
or U7827 (N_7827,N_7749,N_7725);
and U7828 (N_7828,N_7529,N_7677);
nor U7829 (N_7829,N_7655,N_7727);
nand U7830 (N_7830,N_7659,N_7557);
nor U7831 (N_7831,N_7650,N_7512);
or U7832 (N_7832,N_7622,N_7572);
nand U7833 (N_7833,N_7597,N_7549);
and U7834 (N_7834,N_7593,N_7748);
nor U7835 (N_7835,N_7608,N_7714);
nand U7836 (N_7836,N_7563,N_7699);
or U7837 (N_7837,N_7641,N_7617);
nor U7838 (N_7838,N_7718,N_7744);
or U7839 (N_7839,N_7627,N_7681);
or U7840 (N_7840,N_7539,N_7502);
nand U7841 (N_7841,N_7500,N_7511);
xnor U7842 (N_7842,N_7525,N_7623);
nor U7843 (N_7843,N_7501,N_7720);
and U7844 (N_7844,N_7560,N_7612);
or U7845 (N_7845,N_7738,N_7678);
nor U7846 (N_7846,N_7667,N_7632);
and U7847 (N_7847,N_7657,N_7518);
nand U7848 (N_7848,N_7614,N_7583);
or U7849 (N_7849,N_7647,N_7680);
xnor U7850 (N_7850,N_7626,N_7613);
and U7851 (N_7851,N_7519,N_7689);
nor U7852 (N_7852,N_7708,N_7741);
or U7853 (N_7853,N_7696,N_7707);
nand U7854 (N_7854,N_7532,N_7724);
or U7855 (N_7855,N_7588,N_7601);
nor U7856 (N_7856,N_7596,N_7671);
or U7857 (N_7857,N_7723,N_7661);
and U7858 (N_7858,N_7642,N_7576);
xnor U7859 (N_7859,N_7717,N_7694);
nor U7860 (N_7860,N_7728,N_7524);
nand U7861 (N_7861,N_7543,N_7528);
and U7862 (N_7862,N_7695,N_7643);
and U7863 (N_7863,N_7636,N_7571);
or U7864 (N_7864,N_7544,N_7663);
nor U7865 (N_7865,N_7526,N_7640);
xnor U7866 (N_7866,N_7682,N_7537);
nor U7867 (N_7867,N_7530,N_7685);
nor U7868 (N_7868,N_7619,N_7630);
and U7869 (N_7869,N_7631,N_7634);
nor U7870 (N_7870,N_7517,N_7562);
nor U7871 (N_7871,N_7732,N_7706);
or U7872 (N_7872,N_7599,N_7726);
nand U7873 (N_7873,N_7672,N_7645);
and U7874 (N_7874,N_7581,N_7743);
and U7875 (N_7875,N_7703,N_7571);
nand U7876 (N_7876,N_7635,N_7746);
nand U7877 (N_7877,N_7527,N_7580);
or U7878 (N_7878,N_7631,N_7743);
nor U7879 (N_7879,N_7517,N_7559);
nand U7880 (N_7880,N_7555,N_7502);
and U7881 (N_7881,N_7503,N_7502);
nand U7882 (N_7882,N_7522,N_7682);
nor U7883 (N_7883,N_7505,N_7740);
or U7884 (N_7884,N_7539,N_7718);
and U7885 (N_7885,N_7680,N_7529);
and U7886 (N_7886,N_7718,N_7660);
and U7887 (N_7887,N_7625,N_7693);
nand U7888 (N_7888,N_7745,N_7541);
xnor U7889 (N_7889,N_7667,N_7510);
nor U7890 (N_7890,N_7734,N_7641);
nor U7891 (N_7891,N_7536,N_7601);
or U7892 (N_7892,N_7643,N_7744);
nand U7893 (N_7893,N_7529,N_7738);
xnor U7894 (N_7894,N_7547,N_7630);
nand U7895 (N_7895,N_7659,N_7624);
nand U7896 (N_7896,N_7551,N_7576);
or U7897 (N_7897,N_7646,N_7630);
or U7898 (N_7898,N_7582,N_7704);
xor U7899 (N_7899,N_7586,N_7630);
nand U7900 (N_7900,N_7655,N_7536);
and U7901 (N_7901,N_7638,N_7654);
xnor U7902 (N_7902,N_7681,N_7576);
or U7903 (N_7903,N_7663,N_7619);
nand U7904 (N_7904,N_7604,N_7565);
nand U7905 (N_7905,N_7634,N_7718);
xor U7906 (N_7906,N_7513,N_7690);
nand U7907 (N_7907,N_7682,N_7589);
and U7908 (N_7908,N_7638,N_7554);
nor U7909 (N_7909,N_7741,N_7717);
or U7910 (N_7910,N_7510,N_7511);
xor U7911 (N_7911,N_7551,N_7628);
and U7912 (N_7912,N_7637,N_7506);
and U7913 (N_7913,N_7742,N_7689);
or U7914 (N_7914,N_7554,N_7697);
xnor U7915 (N_7915,N_7640,N_7565);
nor U7916 (N_7916,N_7719,N_7712);
and U7917 (N_7917,N_7706,N_7601);
or U7918 (N_7918,N_7654,N_7660);
or U7919 (N_7919,N_7553,N_7631);
nand U7920 (N_7920,N_7697,N_7719);
and U7921 (N_7921,N_7682,N_7642);
nor U7922 (N_7922,N_7599,N_7735);
or U7923 (N_7923,N_7574,N_7526);
nand U7924 (N_7924,N_7749,N_7631);
or U7925 (N_7925,N_7631,N_7664);
and U7926 (N_7926,N_7635,N_7638);
nand U7927 (N_7927,N_7555,N_7677);
or U7928 (N_7928,N_7564,N_7509);
nor U7929 (N_7929,N_7504,N_7624);
and U7930 (N_7930,N_7690,N_7737);
or U7931 (N_7931,N_7646,N_7521);
and U7932 (N_7932,N_7576,N_7684);
nor U7933 (N_7933,N_7659,N_7636);
and U7934 (N_7934,N_7685,N_7679);
nor U7935 (N_7935,N_7625,N_7706);
nor U7936 (N_7936,N_7549,N_7640);
nand U7937 (N_7937,N_7684,N_7553);
xnor U7938 (N_7938,N_7691,N_7624);
nand U7939 (N_7939,N_7610,N_7593);
nand U7940 (N_7940,N_7554,N_7522);
nand U7941 (N_7941,N_7500,N_7723);
xor U7942 (N_7942,N_7587,N_7670);
nor U7943 (N_7943,N_7665,N_7645);
nand U7944 (N_7944,N_7574,N_7575);
and U7945 (N_7945,N_7736,N_7550);
nor U7946 (N_7946,N_7588,N_7542);
and U7947 (N_7947,N_7699,N_7723);
or U7948 (N_7948,N_7632,N_7518);
nand U7949 (N_7949,N_7542,N_7646);
or U7950 (N_7950,N_7581,N_7613);
nor U7951 (N_7951,N_7677,N_7563);
nand U7952 (N_7952,N_7705,N_7573);
or U7953 (N_7953,N_7727,N_7503);
nor U7954 (N_7954,N_7564,N_7710);
nor U7955 (N_7955,N_7582,N_7500);
and U7956 (N_7956,N_7548,N_7748);
nor U7957 (N_7957,N_7559,N_7564);
and U7958 (N_7958,N_7662,N_7548);
nor U7959 (N_7959,N_7694,N_7719);
or U7960 (N_7960,N_7704,N_7513);
nor U7961 (N_7961,N_7592,N_7570);
nor U7962 (N_7962,N_7557,N_7609);
or U7963 (N_7963,N_7718,N_7689);
or U7964 (N_7964,N_7643,N_7544);
nor U7965 (N_7965,N_7620,N_7538);
nand U7966 (N_7966,N_7590,N_7735);
nor U7967 (N_7967,N_7609,N_7589);
or U7968 (N_7968,N_7581,N_7722);
or U7969 (N_7969,N_7623,N_7597);
or U7970 (N_7970,N_7723,N_7536);
nand U7971 (N_7971,N_7658,N_7615);
nor U7972 (N_7972,N_7603,N_7535);
nor U7973 (N_7973,N_7531,N_7530);
nor U7974 (N_7974,N_7637,N_7623);
nor U7975 (N_7975,N_7740,N_7624);
nor U7976 (N_7976,N_7636,N_7641);
nor U7977 (N_7977,N_7739,N_7531);
and U7978 (N_7978,N_7510,N_7580);
nand U7979 (N_7979,N_7644,N_7710);
nor U7980 (N_7980,N_7609,N_7532);
nor U7981 (N_7981,N_7667,N_7596);
xnor U7982 (N_7982,N_7570,N_7530);
or U7983 (N_7983,N_7591,N_7515);
nand U7984 (N_7984,N_7659,N_7514);
xor U7985 (N_7985,N_7674,N_7508);
nand U7986 (N_7986,N_7552,N_7507);
and U7987 (N_7987,N_7592,N_7673);
nand U7988 (N_7988,N_7673,N_7560);
nand U7989 (N_7989,N_7701,N_7679);
or U7990 (N_7990,N_7574,N_7670);
nor U7991 (N_7991,N_7735,N_7658);
nor U7992 (N_7992,N_7573,N_7681);
and U7993 (N_7993,N_7612,N_7501);
and U7994 (N_7994,N_7635,N_7610);
xnor U7995 (N_7995,N_7715,N_7639);
nor U7996 (N_7996,N_7598,N_7603);
nand U7997 (N_7997,N_7749,N_7624);
xor U7998 (N_7998,N_7675,N_7503);
and U7999 (N_7999,N_7667,N_7725);
and U8000 (N_8000,N_7846,N_7930);
nand U8001 (N_8001,N_7990,N_7993);
nand U8002 (N_8002,N_7776,N_7849);
or U8003 (N_8003,N_7772,N_7841);
nor U8004 (N_8004,N_7911,N_7751);
or U8005 (N_8005,N_7853,N_7754);
or U8006 (N_8006,N_7997,N_7908);
or U8007 (N_8007,N_7855,N_7770);
nand U8008 (N_8008,N_7904,N_7813);
and U8009 (N_8009,N_7869,N_7866);
nor U8010 (N_8010,N_7795,N_7757);
and U8011 (N_8011,N_7948,N_7859);
nand U8012 (N_8012,N_7825,N_7839);
nor U8013 (N_8013,N_7890,N_7919);
xnor U8014 (N_8014,N_7774,N_7845);
xor U8015 (N_8015,N_7935,N_7955);
nor U8016 (N_8016,N_7932,N_7898);
and U8017 (N_8017,N_7791,N_7817);
nor U8018 (N_8018,N_7802,N_7984);
and U8019 (N_8019,N_7937,N_7941);
and U8020 (N_8020,N_7758,N_7934);
or U8021 (N_8021,N_7992,N_7820);
and U8022 (N_8022,N_7793,N_7856);
nand U8023 (N_8023,N_7848,N_7933);
nand U8024 (N_8024,N_7969,N_7819);
or U8025 (N_8025,N_7868,N_7837);
nand U8026 (N_8026,N_7957,N_7756);
or U8027 (N_8027,N_7906,N_7854);
or U8028 (N_8028,N_7925,N_7794);
or U8029 (N_8029,N_7750,N_7939);
xnor U8030 (N_8030,N_7796,N_7987);
xnor U8031 (N_8031,N_7885,N_7901);
xor U8032 (N_8032,N_7840,N_7959);
and U8033 (N_8033,N_7809,N_7886);
nor U8034 (N_8034,N_7927,N_7781);
or U8035 (N_8035,N_7807,N_7755);
nor U8036 (N_8036,N_7910,N_7780);
or U8037 (N_8037,N_7893,N_7828);
nor U8038 (N_8038,N_7940,N_7827);
nand U8039 (N_8039,N_7778,N_7752);
and U8040 (N_8040,N_7982,N_7980);
or U8041 (N_8041,N_7870,N_7924);
nor U8042 (N_8042,N_7892,N_7769);
or U8043 (N_8043,N_7804,N_7888);
xnor U8044 (N_8044,N_7943,N_7865);
nor U8045 (N_8045,N_7788,N_7958);
nor U8046 (N_8046,N_7917,N_7949);
nand U8047 (N_8047,N_7862,N_7902);
nand U8048 (N_8048,N_7831,N_7792);
or U8049 (N_8049,N_7830,N_7883);
nor U8050 (N_8050,N_7852,N_7929);
or U8051 (N_8051,N_7844,N_7847);
and U8052 (N_8052,N_7767,N_7873);
nor U8053 (N_8053,N_7981,N_7962);
or U8054 (N_8054,N_7834,N_7971);
or U8055 (N_8055,N_7833,N_7832);
or U8056 (N_8056,N_7814,N_7961);
nor U8057 (N_8057,N_7995,N_7826);
or U8058 (N_8058,N_7864,N_7976);
nor U8059 (N_8059,N_7900,N_7956);
and U8060 (N_8060,N_7871,N_7775);
nor U8061 (N_8061,N_7763,N_7936);
nor U8062 (N_8062,N_7996,N_7963);
nand U8063 (N_8063,N_7920,N_7979);
and U8064 (N_8064,N_7838,N_7875);
or U8065 (N_8065,N_7913,N_7761);
nand U8066 (N_8066,N_7880,N_7782);
and U8067 (N_8067,N_7994,N_7765);
or U8068 (N_8068,N_7822,N_7882);
xnor U8069 (N_8069,N_7811,N_7973);
nand U8070 (N_8070,N_7968,N_7881);
nor U8071 (N_8071,N_7786,N_7824);
and U8072 (N_8072,N_7815,N_7787);
or U8073 (N_8073,N_7887,N_7966);
nand U8074 (N_8074,N_7779,N_7896);
nand U8075 (N_8075,N_7857,N_7800);
or U8076 (N_8076,N_7914,N_7867);
nor U8077 (N_8077,N_7829,N_7816);
and U8078 (N_8078,N_7912,N_7773);
nand U8079 (N_8079,N_7860,N_7874);
nor U8080 (N_8080,N_7998,N_7823);
nand U8081 (N_8081,N_7954,N_7762);
nor U8082 (N_8082,N_7897,N_7999);
nor U8083 (N_8083,N_7797,N_7808);
nand U8084 (N_8084,N_7926,N_7953);
nand U8085 (N_8085,N_7812,N_7783);
and U8086 (N_8086,N_7952,N_7806);
and U8087 (N_8087,N_7766,N_7799);
and U8088 (N_8088,N_7991,N_7798);
nand U8089 (N_8089,N_7891,N_7965);
nand U8090 (N_8090,N_7876,N_7843);
nor U8091 (N_8091,N_7821,N_7905);
nor U8092 (N_8092,N_7916,N_7803);
nor U8093 (N_8093,N_7805,N_7789);
and U8094 (N_8094,N_7771,N_7921);
nand U8095 (N_8095,N_7877,N_7790);
or U8096 (N_8096,N_7967,N_7836);
and U8097 (N_8097,N_7760,N_7974);
xnor U8098 (N_8098,N_7960,N_7938);
nor U8099 (N_8099,N_7764,N_7909);
nor U8100 (N_8100,N_7989,N_7858);
and U8101 (N_8101,N_7946,N_7851);
nor U8102 (N_8102,N_7879,N_7988);
or U8103 (N_8103,N_7759,N_7923);
or U8104 (N_8104,N_7872,N_7889);
and U8105 (N_8105,N_7915,N_7977);
or U8106 (N_8106,N_7978,N_7907);
or U8107 (N_8107,N_7947,N_7928);
nor U8108 (N_8108,N_7903,N_7861);
or U8109 (N_8109,N_7951,N_7918);
or U8110 (N_8110,N_7970,N_7884);
nor U8111 (N_8111,N_7768,N_7942);
nor U8112 (N_8112,N_7842,N_7753);
nor U8113 (N_8113,N_7835,N_7777);
nand U8114 (N_8114,N_7922,N_7878);
or U8115 (N_8115,N_7785,N_7945);
and U8116 (N_8116,N_7801,N_7895);
nand U8117 (N_8117,N_7985,N_7986);
nand U8118 (N_8118,N_7950,N_7894);
nor U8119 (N_8119,N_7784,N_7899);
and U8120 (N_8120,N_7810,N_7972);
xor U8121 (N_8121,N_7850,N_7944);
and U8122 (N_8122,N_7975,N_7983);
nor U8123 (N_8123,N_7931,N_7964);
or U8124 (N_8124,N_7818,N_7863);
nand U8125 (N_8125,N_7942,N_7839);
and U8126 (N_8126,N_7824,N_7967);
and U8127 (N_8127,N_7968,N_7817);
xnor U8128 (N_8128,N_7897,N_7979);
nand U8129 (N_8129,N_7866,N_7780);
nand U8130 (N_8130,N_7981,N_7865);
nand U8131 (N_8131,N_7838,N_7777);
nor U8132 (N_8132,N_7949,N_7943);
nor U8133 (N_8133,N_7777,N_7903);
nor U8134 (N_8134,N_7953,N_7975);
nand U8135 (N_8135,N_7998,N_7990);
and U8136 (N_8136,N_7972,N_7953);
nor U8137 (N_8137,N_7821,N_7966);
or U8138 (N_8138,N_7871,N_7856);
xnor U8139 (N_8139,N_7911,N_7859);
nor U8140 (N_8140,N_7887,N_7929);
nor U8141 (N_8141,N_7917,N_7836);
or U8142 (N_8142,N_7958,N_7999);
and U8143 (N_8143,N_7856,N_7772);
xor U8144 (N_8144,N_7784,N_7845);
or U8145 (N_8145,N_7773,N_7851);
and U8146 (N_8146,N_7977,N_7945);
nor U8147 (N_8147,N_7775,N_7768);
xnor U8148 (N_8148,N_7830,N_7907);
nor U8149 (N_8149,N_7845,N_7773);
xnor U8150 (N_8150,N_7977,N_7901);
and U8151 (N_8151,N_7907,N_7920);
nand U8152 (N_8152,N_7763,N_7867);
and U8153 (N_8153,N_7993,N_7883);
and U8154 (N_8154,N_7953,N_7911);
nor U8155 (N_8155,N_7998,N_7866);
nor U8156 (N_8156,N_7987,N_7835);
xnor U8157 (N_8157,N_7972,N_7815);
and U8158 (N_8158,N_7967,N_7842);
nand U8159 (N_8159,N_7986,N_7965);
and U8160 (N_8160,N_7919,N_7900);
xnor U8161 (N_8161,N_7925,N_7931);
nor U8162 (N_8162,N_7865,N_7835);
nor U8163 (N_8163,N_7923,N_7812);
and U8164 (N_8164,N_7835,N_7901);
nand U8165 (N_8165,N_7973,N_7816);
nand U8166 (N_8166,N_7766,N_7964);
or U8167 (N_8167,N_7956,N_7875);
nor U8168 (N_8168,N_7765,N_7881);
xnor U8169 (N_8169,N_7896,N_7846);
or U8170 (N_8170,N_7889,N_7995);
or U8171 (N_8171,N_7958,N_7854);
xor U8172 (N_8172,N_7905,N_7767);
or U8173 (N_8173,N_7976,N_7967);
nand U8174 (N_8174,N_7888,N_7797);
nor U8175 (N_8175,N_7855,N_7881);
or U8176 (N_8176,N_7843,N_7809);
or U8177 (N_8177,N_7842,N_7767);
xnor U8178 (N_8178,N_7961,N_7860);
nor U8179 (N_8179,N_7753,N_7909);
nand U8180 (N_8180,N_7974,N_7947);
xor U8181 (N_8181,N_7962,N_7893);
and U8182 (N_8182,N_7913,N_7940);
and U8183 (N_8183,N_7758,N_7899);
xor U8184 (N_8184,N_7928,N_7891);
nor U8185 (N_8185,N_7760,N_7937);
xnor U8186 (N_8186,N_7946,N_7756);
or U8187 (N_8187,N_7965,N_7868);
nor U8188 (N_8188,N_7758,N_7869);
and U8189 (N_8189,N_7888,N_7830);
nand U8190 (N_8190,N_7811,N_7993);
or U8191 (N_8191,N_7986,N_7831);
or U8192 (N_8192,N_7869,N_7780);
nand U8193 (N_8193,N_7804,N_7849);
nor U8194 (N_8194,N_7850,N_7762);
or U8195 (N_8195,N_7901,N_7762);
nand U8196 (N_8196,N_7947,N_7793);
and U8197 (N_8197,N_7913,N_7783);
nand U8198 (N_8198,N_7823,N_7844);
nor U8199 (N_8199,N_7792,N_7795);
and U8200 (N_8200,N_7801,N_7826);
xnor U8201 (N_8201,N_7764,N_7873);
nor U8202 (N_8202,N_7836,N_7901);
nand U8203 (N_8203,N_7883,N_7898);
nor U8204 (N_8204,N_7866,N_7897);
or U8205 (N_8205,N_7964,N_7753);
nor U8206 (N_8206,N_7848,N_7971);
or U8207 (N_8207,N_7965,N_7916);
and U8208 (N_8208,N_7998,N_7876);
and U8209 (N_8209,N_7982,N_7941);
nor U8210 (N_8210,N_7835,N_7827);
nor U8211 (N_8211,N_7799,N_7753);
or U8212 (N_8212,N_7947,N_7875);
nor U8213 (N_8213,N_7830,N_7903);
and U8214 (N_8214,N_7897,N_7889);
and U8215 (N_8215,N_7869,N_7794);
nand U8216 (N_8216,N_7829,N_7919);
nand U8217 (N_8217,N_7843,N_7901);
nand U8218 (N_8218,N_7939,N_7992);
nand U8219 (N_8219,N_7768,N_7896);
nand U8220 (N_8220,N_7753,N_7943);
nor U8221 (N_8221,N_7964,N_7922);
xor U8222 (N_8222,N_7949,N_7912);
and U8223 (N_8223,N_7798,N_7985);
nand U8224 (N_8224,N_7962,N_7836);
nor U8225 (N_8225,N_7990,N_7850);
nand U8226 (N_8226,N_7819,N_7847);
nand U8227 (N_8227,N_7761,N_7861);
or U8228 (N_8228,N_7918,N_7790);
or U8229 (N_8229,N_7912,N_7940);
and U8230 (N_8230,N_7829,N_7926);
nand U8231 (N_8231,N_7897,N_7765);
nor U8232 (N_8232,N_7900,N_7996);
or U8233 (N_8233,N_7848,N_7751);
nor U8234 (N_8234,N_7844,N_7991);
xnor U8235 (N_8235,N_7793,N_7955);
nand U8236 (N_8236,N_7778,N_7761);
or U8237 (N_8237,N_7973,N_7828);
xor U8238 (N_8238,N_7889,N_7867);
or U8239 (N_8239,N_7956,N_7771);
and U8240 (N_8240,N_7786,N_7780);
nand U8241 (N_8241,N_7865,N_7903);
and U8242 (N_8242,N_7932,N_7767);
or U8243 (N_8243,N_7918,N_7892);
and U8244 (N_8244,N_7869,N_7941);
nor U8245 (N_8245,N_7988,N_7952);
xor U8246 (N_8246,N_7800,N_7851);
and U8247 (N_8247,N_7988,N_7813);
or U8248 (N_8248,N_7883,N_7891);
nor U8249 (N_8249,N_7864,N_7986);
nor U8250 (N_8250,N_8106,N_8159);
and U8251 (N_8251,N_8061,N_8152);
and U8252 (N_8252,N_8191,N_8000);
and U8253 (N_8253,N_8079,N_8050);
nand U8254 (N_8254,N_8036,N_8066);
and U8255 (N_8255,N_8199,N_8005);
nand U8256 (N_8256,N_8096,N_8082);
nor U8257 (N_8257,N_8025,N_8116);
nor U8258 (N_8258,N_8167,N_8124);
xnor U8259 (N_8259,N_8042,N_8112);
nand U8260 (N_8260,N_8032,N_8026);
and U8261 (N_8261,N_8238,N_8186);
and U8262 (N_8262,N_8184,N_8245);
xnor U8263 (N_8263,N_8097,N_8049);
nor U8264 (N_8264,N_8142,N_8192);
and U8265 (N_8265,N_8002,N_8239);
nor U8266 (N_8266,N_8157,N_8154);
nor U8267 (N_8267,N_8168,N_8110);
or U8268 (N_8268,N_8017,N_8072);
or U8269 (N_8269,N_8104,N_8003);
and U8270 (N_8270,N_8070,N_8100);
or U8271 (N_8271,N_8113,N_8114);
nand U8272 (N_8272,N_8021,N_8170);
nand U8273 (N_8273,N_8211,N_8014);
and U8274 (N_8274,N_8055,N_8132);
xnor U8275 (N_8275,N_8065,N_8009);
nor U8276 (N_8276,N_8094,N_8229);
or U8277 (N_8277,N_8040,N_8206);
or U8278 (N_8278,N_8024,N_8108);
nand U8279 (N_8279,N_8087,N_8053);
or U8280 (N_8280,N_8085,N_8174);
or U8281 (N_8281,N_8135,N_8225);
nor U8282 (N_8282,N_8016,N_8139);
and U8283 (N_8283,N_8189,N_8218);
and U8284 (N_8284,N_8173,N_8056);
nand U8285 (N_8285,N_8144,N_8099);
xor U8286 (N_8286,N_8249,N_8151);
nand U8287 (N_8287,N_8160,N_8177);
nand U8288 (N_8288,N_8080,N_8234);
nand U8289 (N_8289,N_8196,N_8149);
nor U8290 (N_8290,N_8084,N_8204);
nand U8291 (N_8291,N_8020,N_8242);
nor U8292 (N_8292,N_8076,N_8063);
and U8293 (N_8293,N_8019,N_8122);
and U8294 (N_8294,N_8134,N_8248);
nor U8295 (N_8295,N_8128,N_8010);
nor U8296 (N_8296,N_8045,N_8227);
or U8297 (N_8297,N_8190,N_8233);
and U8298 (N_8298,N_8075,N_8074);
or U8299 (N_8299,N_8059,N_8086);
and U8300 (N_8300,N_8240,N_8247);
nand U8301 (N_8301,N_8064,N_8081);
or U8302 (N_8302,N_8230,N_8164);
xnor U8303 (N_8303,N_8047,N_8237);
nand U8304 (N_8304,N_8095,N_8031);
nand U8305 (N_8305,N_8223,N_8208);
or U8306 (N_8306,N_8029,N_8001);
nand U8307 (N_8307,N_8103,N_8155);
xor U8308 (N_8308,N_8101,N_8068);
xor U8309 (N_8309,N_8058,N_8198);
nor U8310 (N_8310,N_8111,N_8035);
and U8311 (N_8311,N_8102,N_8119);
xnor U8312 (N_8312,N_8083,N_8156);
and U8313 (N_8313,N_8052,N_8127);
and U8314 (N_8314,N_8243,N_8188);
or U8315 (N_8315,N_8141,N_8018);
xor U8316 (N_8316,N_8090,N_8200);
nand U8317 (N_8317,N_8057,N_8030);
and U8318 (N_8318,N_8203,N_8219);
or U8319 (N_8319,N_8163,N_8140);
nor U8320 (N_8320,N_8091,N_8013);
nor U8321 (N_8321,N_8232,N_8185);
and U8322 (N_8322,N_8143,N_8041);
or U8323 (N_8323,N_8246,N_8228);
and U8324 (N_8324,N_8201,N_8109);
xor U8325 (N_8325,N_8202,N_8088);
and U8326 (N_8326,N_8118,N_8078);
and U8327 (N_8327,N_8209,N_8214);
nand U8328 (N_8328,N_8165,N_8092);
or U8329 (N_8329,N_8044,N_8027);
nand U8330 (N_8330,N_8015,N_8069);
and U8331 (N_8331,N_8137,N_8023);
xnor U8332 (N_8332,N_8236,N_8187);
nand U8333 (N_8333,N_8171,N_8241);
or U8334 (N_8334,N_8235,N_8126);
xnor U8335 (N_8335,N_8034,N_8008);
or U8336 (N_8336,N_8117,N_8205);
xnor U8337 (N_8337,N_8007,N_8130);
or U8338 (N_8338,N_8123,N_8129);
xor U8339 (N_8339,N_8048,N_8136);
or U8340 (N_8340,N_8226,N_8105);
nand U8341 (N_8341,N_8178,N_8153);
xnor U8342 (N_8342,N_8212,N_8176);
and U8343 (N_8343,N_8093,N_8133);
nand U8344 (N_8344,N_8125,N_8158);
xnor U8345 (N_8345,N_8175,N_8166);
and U8346 (N_8346,N_8194,N_8181);
nor U8347 (N_8347,N_8231,N_8077);
and U8348 (N_8348,N_8221,N_8067);
nor U8349 (N_8349,N_8146,N_8162);
or U8350 (N_8350,N_8089,N_8147);
nor U8351 (N_8351,N_8180,N_8131);
nor U8352 (N_8352,N_8033,N_8216);
xnor U8353 (N_8353,N_8207,N_8098);
and U8354 (N_8354,N_8222,N_8004);
nand U8355 (N_8355,N_8107,N_8182);
or U8356 (N_8356,N_8043,N_8138);
or U8357 (N_8357,N_8195,N_8054);
nand U8358 (N_8358,N_8224,N_8179);
xnor U8359 (N_8359,N_8051,N_8150);
nor U8360 (N_8360,N_8148,N_8213);
nor U8361 (N_8361,N_8006,N_8038);
nand U8362 (N_8362,N_8172,N_8039);
and U8363 (N_8363,N_8183,N_8193);
or U8364 (N_8364,N_8046,N_8220);
nand U8365 (N_8365,N_8217,N_8197);
and U8366 (N_8366,N_8071,N_8037);
nor U8367 (N_8367,N_8121,N_8161);
and U8368 (N_8368,N_8115,N_8060);
and U8369 (N_8369,N_8210,N_8011);
nor U8370 (N_8370,N_8145,N_8073);
or U8371 (N_8371,N_8215,N_8028);
nor U8372 (N_8372,N_8022,N_8062);
or U8373 (N_8373,N_8120,N_8244);
and U8374 (N_8374,N_8012,N_8169);
nor U8375 (N_8375,N_8008,N_8106);
and U8376 (N_8376,N_8024,N_8084);
or U8377 (N_8377,N_8117,N_8005);
nand U8378 (N_8378,N_8223,N_8224);
nor U8379 (N_8379,N_8036,N_8096);
nor U8380 (N_8380,N_8247,N_8168);
nand U8381 (N_8381,N_8064,N_8058);
and U8382 (N_8382,N_8131,N_8184);
xor U8383 (N_8383,N_8157,N_8036);
nand U8384 (N_8384,N_8232,N_8207);
or U8385 (N_8385,N_8004,N_8157);
nand U8386 (N_8386,N_8153,N_8056);
nand U8387 (N_8387,N_8078,N_8081);
and U8388 (N_8388,N_8137,N_8187);
nand U8389 (N_8389,N_8046,N_8048);
nor U8390 (N_8390,N_8195,N_8239);
nand U8391 (N_8391,N_8070,N_8014);
nand U8392 (N_8392,N_8022,N_8090);
and U8393 (N_8393,N_8069,N_8064);
and U8394 (N_8394,N_8132,N_8096);
nor U8395 (N_8395,N_8143,N_8052);
nor U8396 (N_8396,N_8097,N_8009);
nor U8397 (N_8397,N_8121,N_8005);
or U8398 (N_8398,N_8152,N_8159);
and U8399 (N_8399,N_8172,N_8249);
nor U8400 (N_8400,N_8071,N_8244);
nor U8401 (N_8401,N_8122,N_8182);
and U8402 (N_8402,N_8091,N_8050);
and U8403 (N_8403,N_8068,N_8192);
and U8404 (N_8404,N_8205,N_8089);
xnor U8405 (N_8405,N_8125,N_8008);
nand U8406 (N_8406,N_8071,N_8156);
or U8407 (N_8407,N_8185,N_8001);
or U8408 (N_8408,N_8101,N_8020);
xor U8409 (N_8409,N_8041,N_8038);
or U8410 (N_8410,N_8000,N_8177);
or U8411 (N_8411,N_8034,N_8196);
and U8412 (N_8412,N_8161,N_8082);
nor U8413 (N_8413,N_8215,N_8162);
nand U8414 (N_8414,N_8130,N_8123);
nor U8415 (N_8415,N_8202,N_8010);
or U8416 (N_8416,N_8030,N_8042);
nor U8417 (N_8417,N_8100,N_8064);
or U8418 (N_8418,N_8103,N_8029);
xnor U8419 (N_8419,N_8034,N_8221);
and U8420 (N_8420,N_8192,N_8219);
or U8421 (N_8421,N_8202,N_8008);
or U8422 (N_8422,N_8157,N_8099);
and U8423 (N_8423,N_8196,N_8219);
nand U8424 (N_8424,N_8111,N_8051);
or U8425 (N_8425,N_8034,N_8200);
or U8426 (N_8426,N_8069,N_8144);
and U8427 (N_8427,N_8177,N_8071);
nand U8428 (N_8428,N_8200,N_8037);
nor U8429 (N_8429,N_8216,N_8041);
nor U8430 (N_8430,N_8217,N_8181);
and U8431 (N_8431,N_8137,N_8210);
nor U8432 (N_8432,N_8237,N_8029);
nand U8433 (N_8433,N_8060,N_8211);
or U8434 (N_8434,N_8177,N_8241);
xnor U8435 (N_8435,N_8227,N_8051);
nand U8436 (N_8436,N_8071,N_8095);
or U8437 (N_8437,N_8125,N_8169);
xnor U8438 (N_8438,N_8163,N_8080);
nor U8439 (N_8439,N_8120,N_8042);
and U8440 (N_8440,N_8073,N_8171);
or U8441 (N_8441,N_8048,N_8118);
nor U8442 (N_8442,N_8004,N_8242);
xor U8443 (N_8443,N_8069,N_8155);
nor U8444 (N_8444,N_8115,N_8218);
xnor U8445 (N_8445,N_8245,N_8061);
and U8446 (N_8446,N_8074,N_8130);
and U8447 (N_8447,N_8113,N_8109);
nor U8448 (N_8448,N_8176,N_8227);
nand U8449 (N_8449,N_8002,N_8195);
xnor U8450 (N_8450,N_8063,N_8112);
xnor U8451 (N_8451,N_8217,N_8025);
or U8452 (N_8452,N_8125,N_8136);
and U8453 (N_8453,N_8159,N_8161);
nand U8454 (N_8454,N_8166,N_8071);
or U8455 (N_8455,N_8156,N_8200);
nor U8456 (N_8456,N_8241,N_8228);
nor U8457 (N_8457,N_8175,N_8011);
or U8458 (N_8458,N_8210,N_8031);
and U8459 (N_8459,N_8201,N_8069);
nand U8460 (N_8460,N_8160,N_8037);
nor U8461 (N_8461,N_8150,N_8085);
nor U8462 (N_8462,N_8036,N_8114);
and U8463 (N_8463,N_8104,N_8186);
and U8464 (N_8464,N_8207,N_8094);
nand U8465 (N_8465,N_8024,N_8055);
or U8466 (N_8466,N_8045,N_8039);
xor U8467 (N_8467,N_8069,N_8098);
nand U8468 (N_8468,N_8168,N_8116);
nor U8469 (N_8469,N_8247,N_8010);
xnor U8470 (N_8470,N_8053,N_8043);
nand U8471 (N_8471,N_8104,N_8216);
nand U8472 (N_8472,N_8169,N_8160);
or U8473 (N_8473,N_8057,N_8042);
nand U8474 (N_8474,N_8246,N_8111);
and U8475 (N_8475,N_8017,N_8223);
nand U8476 (N_8476,N_8077,N_8196);
or U8477 (N_8477,N_8109,N_8120);
nor U8478 (N_8478,N_8037,N_8233);
nand U8479 (N_8479,N_8200,N_8116);
and U8480 (N_8480,N_8167,N_8166);
and U8481 (N_8481,N_8170,N_8061);
nor U8482 (N_8482,N_8010,N_8017);
nand U8483 (N_8483,N_8119,N_8132);
and U8484 (N_8484,N_8171,N_8195);
nand U8485 (N_8485,N_8176,N_8083);
xnor U8486 (N_8486,N_8167,N_8204);
xnor U8487 (N_8487,N_8066,N_8215);
nand U8488 (N_8488,N_8233,N_8212);
nor U8489 (N_8489,N_8209,N_8137);
nor U8490 (N_8490,N_8039,N_8070);
nor U8491 (N_8491,N_8044,N_8203);
nor U8492 (N_8492,N_8004,N_8083);
or U8493 (N_8493,N_8102,N_8104);
nand U8494 (N_8494,N_8064,N_8068);
xor U8495 (N_8495,N_8130,N_8042);
and U8496 (N_8496,N_8159,N_8183);
or U8497 (N_8497,N_8142,N_8201);
nor U8498 (N_8498,N_8022,N_8002);
and U8499 (N_8499,N_8243,N_8203);
or U8500 (N_8500,N_8409,N_8460);
nand U8501 (N_8501,N_8384,N_8440);
or U8502 (N_8502,N_8345,N_8378);
nand U8503 (N_8503,N_8447,N_8433);
nand U8504 (N_8504,N_8297,N_8252);
nand U8505 (N_8505,N_8369,N_8438);
and U8506 (N_8506,N_8296,N_8272);
nand U8507 (N_8507,N_8284,N_8387);
nand U8508 (N_8508,N_8388,N_8307);
or U8509 (N_8509,N_8318,N_8482);
xor U8510 (N_8510,N_8453,N_8494);
or U8511 (N_8511,N_8335,N_8465);
nor U8512 (N_8512,N_8302,N_8487);
and U8513 (N_8513,N_8483,N_8491);
nand U8514 (N_8514,N_8313,N_8385);
and U8515 (N_8515,N_8344,N_8396);
or U8516 (N_8516,N_8416,N_8414);
and U8517 (N_8517,N_8295,N_8292);
nand U8518 (N_8518,N_8357,N_8455);
xor U8519 (N_8519,N_8469,N_8490);
and U8520 (N_8520,N_8265,N_8368);
nand U8521 (N_8521,N_8356,N_8410);
or U8522 (N_8522,N_8278,N_8445);
or U8523 (N_8523,N_8383,N_8379);
and U8524 (N_8524,N_8471,N_8449);
xor U8525 (N_8525,N_8289,N_8404);
or U8526 (N_8526,N_8261,N_8314);
nor U8527 (N_8527,N_8452,N_8285);
or U8528 (N_8528,N_8370,N_8463);
or U8529 (N_8529,N_8264,N_8342);
nor U8530 (N_8530,N_8464,N_8254);
or U8531 (N_8531,N_8436,N_8303);
nor U8532 (N_8532,N_8391,N_8477);
and U8533 (N_8533,N_8390,N_8327);
nor U8534 (N_8534,N_8446,N_8435);
nor U8535 (N_8535,N_8301,N_8402);
nand U8536 (N_8536,N_8484,N_8458);
nor U8537 (N_8537,N_8499,N_8389);
or U8538 (N_8538,N_8263,N_8280);
nor U8539 (N_8539,N_8317,N_8485);
and U8540 (N_8540,N_8415,N_8334);
nor U8541 (N_8541,N_8277,N_8258);
nand U8542 (N_8542,N_8444,N_8359);
nor U8543 (N_8543,N_8260,N_8308);
and U8544 (N_8544,N_8478,N_8405);
xnor U8545 (N_8545,N_8443,N_8325);
and U8546 (N_8546,N_8266,N_8286);
nand U8547 (N_8547,N_8288,N_8293);
and U8548 (N_8548,N_8290,N_8256);
or U8549 (N_8549,N_8337,N_8320);
or U8550 (N_8550,N_8456,N_8412);
and U8551 (N_8551,N_8399,N_8495);
or U8552 (N_8552,N_8372,N_8321);
and U8553 (N_8553,N_8418,N_8343);
nand U8554 (N_8554,N_8498,N_8281);
or U8555 (N_8555,N_8459,N_8376);
nor U8556 (N_8556,N_8255,N_8466);
and U8557 (N_8557,N_8393,N_8341);
and U8558 (N_8558,N_8291,N_8322);
or U8559 (N_8559,N_8274,N_8431);
nand U8560 (N_8560,N_8309,N_8421);
or U8561 (N_8561,N_8294,N_8442);
nor U8562 (N_8562,N_8437,N_8319);
and U8563 (N_8563,N_8411,N_8331);
or U8564 (N_8564,N_8400,N_8493);
and U8565 (N_8565,N_8353,N_8394);
nor U8566 (N_8566,N_8408,N_8324);
nor U8567 (N_8567,N_8271,N_8417);
or U8568 (N_8568,N_8364,N_8282);
nand U8569 (N_8569,N_8304,N_8473);
xor U8570 (N_8570,N_8413,N_8333);
or U8571 (N_8571,N_8323,N_8434);
xnor U8572 (N_8572,N_8428,N_8315);
nand U8573 (N_8573,N_8312,N_8496);
or U8574 (N_8574,N_8339,N_8480);
xor U8575 (N_8575,N_8423,N_8276);
nand U8576 (N_8576,N_8475,N_8283);
and U8577 (N_8577,N_8358,N_8497);
xor U8578 (N_8578,N_8360,N_8373);
nand U8579 (N_8579,N_8430,N_8250);
or U8580 (N_8580,N_8305,N_8316);
and U8581 (N_8581,N_8425,N_8457);
or U8582 (N_8582,N_8349,N_8299);
and U8583 (N_8583,N_8448,N_8382);
or U8584 (N_8584,N_8406,N_8287);
nand U8585 (N_8585,N_8377,N_8251);
or U8586 (N_8586,N_8467,N_8361);
nand U8587 (N_8587,N_8298,N_8439);
nor U8588 (N_8588,N_8386,N_8340);
nor U8589 (N_8589,N_8450,N_8338);
xor U8590 (N_8590,N_8311,N_8374);
nand U8591 (N_8591,N_8259,N_8269);
or U8592 (N_8592,N_8367,N_8474);
xnor U8593 (N_8593,N_8429,N_8489);
and U8594 (N_8594,N_8420,N_8257);
nor U8595 (N_8595,N_8461,N_8306);
nor U8596 (N_8596,N_8352,N_8486);
and U8597 (N_8597,N_8300,N_8363);
or U8598 (N_8598,N_8268,N_8347);
nor U8599 (N_8599,N_8365,N_8351);
or U8600 (N_8600,N_8488,N_8419);
and U8601 (N_8601,N_8479,N_8381);
and U8602 (N_8602,N_8326,N_8468);
and U8603 (N_8603,N_8262,N_8427);
or U8604 (N_8604,N_8441,N_8273);
nor U8605 (N_8605,N_8350,N_8375);
xor U8606 (N_8606,N_8422,N_8462);
and U8607 (N_8607,N_8279,N_8366);
nand U8608 (N_8608,N_8392,N_8476);
nor U8609 (N_8609,N_8398,N_8401);
nor U8610 (N_8610,N_8270,N_8424);
or U8611 (N_8611,N_8332,N_8310);
nand U8612 (N_8612,N_8397,N_8395);
and U8613 (N_8613,N_8275,N_8380);
or U8614 (N_8614,N_8432,N_8362);
and U8615 (N_8615,N_8451,N_8354);
nand U8616 (N_8616,N_8355,N_8407);
and U8617 (N_8617,N_8426,N_8329);
or U8618 (N_8618,N_8371,N_8336);
or U8619 (N_8619,N_8470,N_8267);
nand U8620 (N_8620,N_8330,N_8253);
or U8621 (N_8621,N_8348,N_8328);
or U8622 (N_8622,N_8492,N_8346);
and U8623 (N_8623,N_8454,N_8481);
nor U8624 (N_8624,N_8403,N_8472);
nor U8625 (N_8625,N_8309,N_8428);
xor U8626 (N_8626,N_8456,N_8317);
and U8627 (N_8627,N_8441,N_8432);
or U8628 (N_8628,N_8441,N_8272);
xnor U8629 (N_8629,N_8476,N_8432);
nand U8630 (N_8630,N_8252,N_8270);
and U8631 (N_8631,N_8381,N_8332);
nor U8632 (N_8632,N_8459,N_8483);
and U8633 (N_8633,N_8348,N_8373);
or U8634 (N_8634,N_8253,N_8490);
nand U8635 (N_8635,N_8267,N_8327);
xnor U8636 (N_8636,N_8439,N_8251);
nand U8637 (N_8637,N_8379,N_8421);
or U8638 (N_8638,N_8454,N_8345);
nand U8639 (N_8639,N_8482,N_8356);
or U8640 (N_8640,N_8402,N_8426);
or U8641 (N_8641,N_8376,N_8377);
or U8642 (N_8642,N_8475,N_8484);
xnor U8643 (N_8643,N_8371,N_8287);
nand U8644 (N_8644,N_8352,N_8424);
nor U8645 (N_8645,N_8434,N_8344);
nor U8646 (N_8646,N_8465,N_8495);
nor U8647 (N_8647,N_8323,N_8270);
nand U8648 (N_8648,N_8492,N_8345);
nand U8649 (N_8649,N_8444,N_8421);
nand U8650 (N_8650,N_8300,N_8252);
and U8651 (N_8651,N_8412,N_8347);
nand U8652 (N_8652,N_8414,N_8424);
or U8653 (N_8653,N_8433,N_8355);
or U8654 (N_8654,N_8281,N_8319);
or U8655 (N_8655,N_8337,N_8332);
xor U8656 (N_8656,N_8398,N_8435);
or U8657 (N_8657,N_8490,N_8488);
or U8658 (N_8658,N_8371,N_8323);
xnor U8659 (N_8659,N_8303,N_8384);
or U8660 (N_8660,N_8343,N_8380);
nor U8661 (N_8661,N_8376,N_8485);
and U8662 (N_8662,N_8288,N_8481);
nand U8663 (N_8663,N_8402,N_8254);
or U8664 (N_8664,N_8425,N_8299);
and U8665 (N_8665,N_8369,N_8295);
or U8666 (N_8666,N_8321,N_8444);
or U8667 (N_8667,N_8369,N_8463);
and U8668 (N_8668,N_8469,N_8405);
xnor U8669 (N_8669,N_8449,N_8305);
or U8670 (N_8670,N_8341,N_8412);
xnor U8671 (N_8671,N_8456,N_8342);
or U8672 (N_8672,N_8283,N_8492);
nor U8673 (N_8673,N_8251,N_8286);
nor U8674 (N_8674,N_8365,N_8438);
or U8675 (N_8675,N_8302,N_8482);
and U8676 (N_8676,N_8482,N_8260);
and U8677 (N_8677,N_8431,N_8350);
nand U8678 (N_8678,N_8323,N_8421);
and U8679 (N_8679,N_8251,N_8289);
or U8680 (N_8680,N_8286,N_8365);
and U8681 (N_8681,N_8441,N_8263);
xor U8682 (N_8682,N_8489,N_8307);
nor U8683 (N_8683,N_8259,N_8476);
nor U8684 (N_8684,N_8308,N_8339);
or U8685 (N_8685,N_8316,N_8460);
nor U8686 (N_8686,N_8427,N_8340);
and U8687 (N_8687,N_8253,N_8353);
nor U8688 (N_8688,N_8250,N_8375);
nor U8689 (N_8689,N_8316,N_8324);
or U8690 (N_8690,N_8363,N_8345);
xnor U8691 (N_8691,N_8497,N_8360);
nand U8692 (N_8692,N_8406,N_8415);
and U8693 (N_8693,N_8314,N_8431);
or U8694 (N_8694,N_8459,N_8429);
nand U8695 (N_8695,N_8402,N_8394);
nor U8696 (N_8696,N_8271,N_8391);
nand U8697 (N_8697,N_8416,N_8462);
xnor U8698 (N_8698,N_8441,N_8486);
and U8699 (N_8699,N_8365,N_8331);
nand U8700 (N_8700,N_8432,N_8411);
or U8701 (N_8701,N_8498,N_8253);
or U8702 (N_8702,N_8381,N_8478);
or U8703 (N_8703,N_8317,N_8498);
nor U8704 (N_8704,N_8371,N_8447);
or U8705 (N_8705,N_8334,N_8287);
and U8706 (N_8706,N_8437,N_8329);
nor U8707 (N_8707,N_8448,N_8253);
and U8708 (N_8708,N_8452,N_8327);
and U8709 (N_8709,N_8318,N_8324);
nand U8710 (N_8710,N_8282,N_8320);
xor U8711 (N_8711,N_8304,N_8286);
and U8712 (N_8712,N_8348,N_8491);
nand U8713 (N_8713,N_8268,N_8432);
and U8714 (N_8714,N_8390,N_8374);
nand U8715 (N_8715,N_8318,N_8383);
or U8716 (N_8716,N_8466,N_8417);
nor U8717 (N_8717,N_8392,N_8284);
nor U8718 (N_8718,N_8459,N_8337);
nor U8719 (N_8719,N_8365,N_8472);
nand U8720 (N_8720,N_8474,N_8312);
or U8721 (N_8721,N_8289,N_8459);
nor U8722 (N_8722,N_8452,N_8284);
nor U8723 (N_8723,N_8317,N_8332);
nor U8724 (N_8724,N_8271,N_8307);
or U8725 (N_8725,N_8379,N_8487);
nor U8726 (N_8726,N_8454,N_8489);
and U8727 (N_8727,N_8394,N_8309);
nand U8728 (N_8728,N_8398,N_8457);
or U8729 (N_8729,N_8496,N_8446);
nor U8730 (N_8730,N_8360,N_8301);
or U8731 (N_8731,N_8451,N_8363);
or U8732 (N_8732,N_8348,N_8301);
or U8733 (N_8733,N_8408,N_8389);
nor U8734 (N_8734,N_8468,N_8442);
nor U8735 (N_8735,N_8344,N_8316);
nand U8736 (N_8736,N_8256,N_8336);
and U8737 (N_8737,N_8444,N_8378);
or U8738 (N_8738,N_8250,N_8292);
and U8739 (N_8739,N_8312,N_8289);
xnor U8740 (N_8740,N_8373,N_8446);
nor U8741 (N_8741,N_8291,N_8466);
nand U8742 (N_8742,N_8352,N_8443);
nor U8743 (N_8743,N_8312,N_8393);
and U8744 (N_8744,N_8495,N_8498);
nor U8745 (N_8745,N_8360,N_8363);
or U8746 (N_8746,N_8309,N_8488);
and U8747 (N_8747,N_8340,N_8481);
and U8748 (N_8748,N_8431,N_8325);
and U8749 (N_8749,N_8340,N_8293);
or U8750 (N_8750,N_8601,N_8715);
nor U8751 (N_8751,N_8548,N_8545);
or U8752 (N_8752,N_8625,N_8717);
nor U8753 (N_8753,N_8523,N_8580);
and U8754 (N_8754,N_8526,N_8515);
xnor U8755 (N_8755,N_8513,N_8655);
nor U8756 (N_8756,N_8719,N_8666);
nand U8757 (N_8757,N_8501,N_8564);
and U8758 (N_8758,N_8565,N_8691);
nor U8759 (N_8759,N_8516,N_8739);
or U8760 (N_8760,N_8631,N_8520);
nand U8761 (N_8761,N_8693,N_8543);
nand U8762 (N_8762,N_8728,N_8641);
or U8763 (N_8763,N_8542,N_8592);
nand U8764 (N_8764,N_8574,N_8714);
nand U8765 (N_8765,N_8658,N_8670);
xor U8766 (N_8766,N_8688,N_8649);
xor U8767 (N_8767,N_8698,N_8554);
and U8768 (N_8768,N_8732,N_8620);
and U8769 (N_8769,N_8558,N_8539);
or U8770 (N_8770,N_8503,N_8612);
nand U8771 (N_8771,N_8736,N_8629);
and U8772 (N_8772,N_8540,N_8737);
xnor U8773 (N_8773,N_8506,N_8725);
or U8774 (N_8774,N_8614,N_8703);
xor U8775 (N_8775,N_8579,N_8690);
xnor U8776 (N_8776,N_8514,N_8557);
nand U8777 (N_8777,N_8624,N_8602);
or U8778 (N_8778,N_8713,N_8561);
nand U8779 (N_8779,N_8528,N_8585);
nand U8780 (N_8780,N_8593,N_8595);
nor U8781 (N_8781,N_8529,N_8591);
or U8782 (N_8782,N_8550,N_8517);
and U8783 (N_8783,N_8672,N_8549);
and U8784 (N_8784,N_8748,N_8709);
and U8785 (N_8785,N_8696,N_8533);
or U8786 (N_8786,N_8570,N_8582);
or U8787 (N_8787,N_8747,N_8621);
and U8788 (N_8788,N_8664,N_8527);
xnor U8789 (N_8789,N_8563,N_8742);
and U8790 (N_8790,N_8692,N_8568);
or U8791 (N_8791,N_8507,N_8706);
or U8792 (N_8792,N_8560,N_8500);
nand U8793 (N_8793,N_8743,N_8668);
xor U8794 (N_8794,N_8589,N_8669);
and U8795 (N_8795,N_8642,N_8701);
or U8796 (N_8796,N_8610,N_8650);
xor U8797 (N_8797,N_8716,N_8578);
and U8798 (N_8798,N_8678,N_8673);
nor U8799 (N_8799,N_8685,N_8628);
nor U8800 (N_8800,N_8519,N_8617);
or U8801 (N_8801,N_8677,N_8600);
xor U8802 (N_8802,N_8594,N_8505);
and U8803 (N_8803,N_8608,N_8643);
and U8804 (N_8804,N_8731,N_8611);
or U8805 (N_8805,N_8730,N_8740);
nor U8806 (N_8806,N_8680,N_8738);
or U8807 (N_8807,N_8660,N_8615);
and U8808 (N_8808,N_8567,N_8534);
nand U8809 (N_8809,N_8577,N_8675);
xor U8810 (N_8810,N_8712,N_8687);
nand U8811 (N_8811,N_8575,N_8576);
and U8812 (N_8812,N_8735,N_8636);
and U8813 (N_8813,N_8679,N_8630);
or U8814 (N_8814,N_8722,N_8654);
xor U8815 (N_8815,N_8555,N_8697);
nor U8816 (N_8816,N_8613,N_8547);
nand U8817 (N_8817,N_8583,N_8559);
nor U8818 (N_8818,N_8535,N_8566);
nor U8819 (N_8819,N_8707,N_8647);
or U8820 (N_8820,N_8512,N_8606);
nand U8821 (N_8821,N_8635,N_8587);
and U8822 (N_8822,N_8708,N_8530);
or U8823 (N_8823,N_8531,N_8639);
or U8824 (N_8824,N_8700,N_8508);
nor U8825 (N_8825,N_8646,N_8683);
xor U8826 (N_8826,N_8599,N_8704);
or U8827 (N_8827,N_8727,N_8541);
nand U8828 (N_8828,N_8640,N_8699);
nand U8829 (N_8829,N_8588,N_8653);
or U8830 (N_8830,N_8537,N_8609);
nand U8831 (N_8831,N_8644,N_8681);
xnor U8832 (N_8832,N_8604,N_8590);
or U8833 (N_8833,N_8645,N_8552);
nor U8834 (N_8834,N_8525,N_8598);
and U8835 (N_8835,N_8584,N_8634);
or U8836 (N_8836,N_8510,N_8532);
nand U8837 (N_8837,N_8607,N_8749);
nor U8838 (N_8838,N_8729,N_8622);
and U8839 (N_8839,N_8652,N_8637);
nor U8840 (N_8840,N_8674,N_8605);
or U8841 (N_8841,N_8734,N_8682);
or U8842 (N_8842,N_8711,N_8745);
nor U8843 (N_8843,N_8511,N_8667);
nor U8844 (N_8844,N_8536,N_8741);
nor U8845 (N_8845,N_8538,N_8596);
xor U8846 (N_8846,N_8603,N_8569);
or U8847 (N_8847,N_8623,N_8581);
nand U8848 (N_8848,N_8695,N_8633);
or U8849 (N_8849,N_8638,N_8648);
and U8850 (N_8850,N_8733,N_8686);
and U8851 (N_8851,N_8702,N_8572);
and U8852 (N_8852,N_8618,N_8662);
and U8853 (N_8853,N_8710,N_8553);
nor U8854 (N_8854,N_8661,N_8651);
nor U8855 (N_8855,N_8556,N_8671);
or U8856 (N_8856,N_8522,N_8597);
nor U8857 (N_8857,N_8504,N_8626);
or U8858 (N_8858,N_8723,N_8718);
nand U8859 (N_8859,N_8509,N_8521);
nand U8860 (N_8860,N_8659,N_8721);
nor U8861 (N_8861,N_8656,N_8573);
or U8862 (N_8862,N_8724,N_8676);
and U8863 (N_8863,N_8544,N_8627);
nor U8864 (N_8864,N_8665,N_8726);
or U8865 (N_8865,N_8684,N_8746);
and U8866 (N_8866,N_8562,N_8632);
nor U8867 (N_8867,N_8663,N_8619);
nor U8868 (N_8868,N_8571,N_8551);
nand U8869 (N_8869,N_8546,N_8744);
xor U8870 (N_8870,N_8586,N_8657);
xnor U8871 (N_8871,N_8524,N_8689);
and U8872 (N_8872,N_8502,N_8705);
nand U8873 (N_8873,N_8694,N_8720);
nand U8874 (N_8874,N_8616,N_8518);
nand U8875 (N_8875,N_8661,N_8571);
and U8876 (N_8876,N_8511,N_8663);
nor U8877 (N_8877,N_8646,N_8633);
nor U8878 (N_8878,N_8718,N_8618);
and U8879 (N_8879,N_8559,N_8613);
and U8880 (N_8880,N_8684,N_8691);
or U8881 (N_8881,N_8664,N_8685);
nand U8882 (N_8882,N_8585,N_8666);
nor U8883 (N_8883,N_8540,N_8684);
nand U8884 (N_8884,N_8711,N_8677);
or U8885 (N_8885,N_8739,N_8657);
and U8886 (N_8886,N_8580,N_8615);
and U8887 (N_8887,N_8580,N_8718);
nand U8888 (N_8888,N_8585,N_8650);
nand U8889 (N_8889,N_8748,N_8610);
nor U8890 (N_8890,N_8646,N_8693);
or U8891 (N_8891,N_8690,N_8719);
and U8892 (N_8892,N_8632,N_8672);
or U8893 (N_8893,N_8619,N_8657);
or U8894 (N_8894,N_8599,N_8656);
and U8895 (N_8895,N_8705,N_8702);
and U8896 (N_8896,N_8579,N_8746);
or U8897 (N_8897,N_8734,N_8584);
and U8898 (N_8898,N_8690,N_8582);
nor U8899 (N_8899,N_8614,N_8633);
and U8900 (N_8900,N_8515,N_8505);
and U8901 (N_8901,N_8748,N_8712);
nor U8902 (N_8902,N_8686,N_8561);
or U8903 (N_8903,N_8742,N_8701);
or U8904 (N_8904,N_8597,N_8656);
nor U8905 (N_8905,N_8704,N_8653);
or U8906 (N_8906,N_8728,N_8700);
and U8907 (N_8907,N_8659,N_8671);
or U8908 (N_8908,N_8523,N_8615);
and U8909 (N_8909,N_8504,N_8569);
nor U8910 (N_8910,N_8628,N_8708);
nor U8911 (N_8911,N_8544,N_8548);
or U8912 (N_8912,N_8729,N_8512);
nor U8913 (N_8913,N_8740,N_8708);
nand U8914 (N_8914,N_8500,N_8566);
nor U8915 (N_8915,N_8510,N_8697);
or U8916 (N_8916,N_8693,N_8515);
nand U8917 (N_8917,N_8646,N_8628);
nor U8918 (N_8918,N_8623,N_8639);
nor U8919 (N_8919,N_8650,N_8526);
or U8920 (N_8920,N_8625,N_8632);
nand U8921 (N_8921,N_8681,N_8641);
or U8922 (N_8922,N_8640,N_8721);
and U8923 (N_8923,N_8618,N_8705);
xor U8924 (N_8924,N_8726,N_8715);
or U8925 (N_8925,N_8647,N_8543);
nor U8926 (N_8926,N_8593,N_8677);
nand U8927 (N_8927,N_8694,N_8596);
or U8928 (N_8928,N_8542,N_8562);
and U8929 (N_8929,N_8740,N_8592);
xnor U8930 (N_8930,N_8574,N_8703);
nor U8931 (N_8931,N_8532,N_8742);
and U8932 (N_8932,N_8709,N_8554);
nor U8933 (N_8933,N_8530,N_8613);
nor U8934 (N_8934,N_8600,N_8520);
nand U8935 (N_8935,N_8550,N_8682);
nand U8936 (N_8936,N_8558,N_8652);
nand U8937 (N_8937,N_8598,N_8518);
and U8938 (N_8938,N_8724,N_8641);
nor U8939 (N_8939,N_8516,N_8679);
nand U8940 (N_8940,N_8554,N_8547);
nand U8941 (N_8941,N_8558,N_8676);
nand U8942 (N_8942,N_8513,N_8571);
nand U8943 (N_8943,N_8549,N_8703);
nand U8944 (N_8944,N_8600,N_8558);
nor U8945 (N_8945,N_8601,N_8634);
or U8946 (N_8946,N_8674,N_8733);
xnor U8947 (N_8947,N_8671,N_8743);
nand U8948 (N_8948,N_8612,N_8638);
and U8949 (N_8949,N_8596,N_8748);
or U8950 (N_8950,N_8720,N_8575);
nand U8951 (N_8951,N_8657,N_8635);
nand U8952 (N_8952,N_8532,N_8563);
or U8953 (N_8953,N_8690,N_8506);
and U8954 (N_8954,N_8638,N_8516);
or U8955 (N_8955,N_8547,N_8582);
nand U8956 (N_8956,N_8504,N_8681);
nand U8957 (N_8957,N_8628,N_8730);
and U8958 (N_8958,N_8563,N_8575);
and U8959 (N_8959,N_8653,N_8730);
or U8960 (N_8960,N_8749,N_8579);
and U8961 (N_8961,N_8645,N_8703);
nand U8962 (N_8962,N_8667,N_8614);
and U8963 (N_8963,N_8738,N_8749);
nor U8964 (N_8964,N_8597,N_8588);
nor U8965 (N_8965,N_8628,N_8568);
and U8966 (N_8966,N_8601,N_8570);
nor U8967 (N_8967,N_8730,N_8569);
or U8968 (N_8968,N_8622,N_8639);
and U8969 (N_8969,N_8656,N_8561);
nor U8970 (N_8970,N_8502,N_8629);
or U8971 (N_8971,N_8516,N_8704);
nor U8972 (N_8972,N_8642,N_8721);
nand U8973 (N_8973,N_8587,N_8593);
and U8974 (N_8974,N_8613,N_8524);
xnor U8975 (N_8975,N_8694,N_8580);
nand U8976 (N_8976,N_8715,N_8682);
or U8977 (N_8977,N_8715,N_8627);
and U8978 (N_8978,N_8534,N_8607);
nor U8979 (N_8979,N_8552,N_8570);
nor U8980 (N_8980,N_8543,N_8578);
and U8981 (N_8981,N_8679,N_8533);
and U8982 (N_8982,N_8613,N_8694);
and U8983 (N_8983,N_8638,N_8716);
or U8984 (N_8984,N_8549,N_8547);
or U8985 (N_8985,N_8696,N_8746);
or U8986 (N_8986,N_8692,N_8749);
and U8987 (N_8987,N_8608,N_8625);
nand U8988 (N_8988,N_8736,N_8707);
and U8989 (N_8989,N_8704,N_8749);
nand U8990 (N_8990,N_8709,N_8519);
nand U8991 (N_8991,N_8518,N_8684);
nand U8992 (N_8992,N_8532,N_8610);
xor U8993 (N_8993,N_8573,N_8563);
nand U8994 (N_8994,N_8523,N_8550);
or U8995 (N_8995,N_8631,N_8744);
nand U8996 (N_8996,N_8616,N_8555);
nand U8997 (N_8997,N_8542,N_8571);
or U8998 (N_8998,N_8567,N_8641);
nand U8999 (N_8999,N_8693,N_8631);
nor U9000 (N_9000,N_8979,N_8800);
xor U9001 (N_9001,N_8975,N_8974);
and U9002 (N_9002,N_8833,N_8968);
and U9003 (N_9003,N_8980,N_8872);
nand U9004 (N_9004,N_8926,N_8981);
or U9005 (N_9005,N_8842,N_8865);
nor U9006 (N_9006,N_8900,N_8886);
nor U9007 (N_9007,N_8940,N_8766);
xnor U9008 (N_9008,N_8826,N_8985);
nor U9009 (N_9009,N_8901,N_8841);
and U9010 (N_9010,N_8783,N_8956);
nor U9011 (N_9011,N_8859,N_8753);
nor U9012 (N_9012,N_8768,N_8804);
nand U9013 (N_9013,N_8870,N_8948);
and U9014 (N_9014,N_8888,N_8908);
nand U9015 (N_9015,N_8879,N_8952);
nand U9016 (N_9016,N_8845,N_8993);
and U9017 (N_9017,N_8860,N_8871);
xnor U9018 (N_9018,N_8933,N_8792);
xnor U9019 (N_9019,N_8898,N_8772);
and U9020 (N_9020,N_8892,N_8893);
or U9021 (N_9021,N_8880,N_8784);
or U9022 (N_9022,N_8797,N_8942);
or U9023 (N_9023,N_8905,N_8799);
nand U9024 (N_9024,N_8978,N_8852);
nand U9025 (N_9025,N_8756,N_8881);
or U9026 (N_9026,N_8821,N_8781);
or U9027 (N_9027,N_8763,N_8820);
or U9028 (N_9028,N_8976,N_8838);
nor U9029 (N_9029,N_8932,N_8912);
and U9030 (N_9030,N_8970,N_8899);
or U9031 (N_9031,N_8996,N_8846);
and U9032 (N_9032,N_8946,N_8903);
nor U9033 (N_9033,N_8943,N_8759);
nor U9034 (N_9034,N_8798,N_8998);
and U9035 (N_9035,N_8844,N_8862);
and U9036 (N_9036,N_8913,N_8895);
or U9037 (N_9037,N_8780,N_8802);
and U9038 (N_9038,N_8855,N_8757);
or U9039 (N_9039,N_8839,N_8851);
nor U9040 (N_9040,N_8961,N_8819);
xor U9041 (N_9041,N_8857,N_8991);
xnor U9042 (N_9042,N_8929,N_8764);
or U9043 (N_9043,N_8779,N_8789);
nor U9044 (N_9044,N_8816,N_8917);
xor U9045 (N_9045,N_8951,N_8761);
or U9046 (N_9046,N_8868,N_8790);
or U9047 (N_9047,N_8924,N_8973);
and U9048 (N_9048,N_8812,N_8807);
nor U9049 (N_9049,N_8923,N_8873);
or U9050 (N_9050,N_8796,N_8752);
nand U9051 (N_9051,N_8849,N_8925);
and U9052 (N_9052,N_8914,N_8966);
and U9053 (N_9053,N_8861,N_8751);
nand U9054 (N_9054,N_8788,N_8863);
nor U9055 (N_9055,N_8941,N_8778);
or U9056 (N_9056,N_8967,N_8989);
nor U9057 (N_9057,N_8755,N_8953);
and U9058 (N_9058,N_8995,N_8769);
nor U9059 (N_9059,N_8896,N_8936);
and U9060 (N_9060,N_8918,N_8904);
nor U9061 (N_9061,N_8808,N_8986);
and U9062 (N_9062,N_8814,N_8824);
nor U9063 (N_9063,N_8876,N_8750);
and U9064 (N_9064,N_8916,N_8889);
nor U9065 (N_9065,N_8954,N_8882);
and U9066 (N_9066,N_8832,N_8960);
nand U9067 (N_9067,N_8885,N_8875);
or U9068 (N_9068,N_8878,N_8847);
nor U9069 (N_9069,N_8977,N_8866);
xor U9070 (N_9070,N_8843,N_8787);
nand U9071 (N_9071,N_8982,N_8958);
nand U9072 (N_9072,N_8915,N_8867);
xor U9073 (N_9073,N_8947,N_8969);
nor U9074 (N_9074,N_8853,N_8765);
and U9075 (N_9075,N_8939,N_8782);
nor U9076 (N_9076,N_8999,N_8927);
and U9077 (N_9077,N_8928,N_8988);
nor U9078 (N_9078,N_8822,N_8771);
xnor U9079 (N_9079,N_8987,N_8934);
nand U9080 (N_9080,N_8931,N_8869);
nand U9081 (N_9081,N_8962,N_8983);
and U9082 (N_9082,N_8754,N_8803);
and U9083 (N_9083,N_8950,N_8806);
nor U9084 (N_9084,N_8890,N_8801);
nand U9085 (N_9085,N_8919,N_8945);
nand U9086 (N_9086,N_8910,N_8937);
or U9087 (N_9087,N_8965,N_8776);
nand U9088 (N_9088,N_8850,N_8955);
nor U9089 (N_9089,N_8959,N_8795);
or U9090 (N_9090,N_8922,N_8840);
and U9091 (N_9091,N_8972,N_8894);
or U9092 (N_9092,N_8813,N_8794);
xnor U9093 (N_9093,N_8829,N_8891);
or U9094 (N_9094,N_8823,N_8774);
and U9095 (N_9095,N_8938,N_8992);
nor U9096 (N_9096,N_8902,N_8770);
and U9097 (N_9097,N_8963,N_8994);
and U9098 (N_9098,N_8836,N_8957);
nand U9099 (N_9099,N_8809,N_8793);
xor U9100 (N_9100,N_8758,N_8949);
or U9101 (N_9101,N_8828,N_8874);
xnor U9102 (N_9102,N_8964,N_8897);
and U9103 (N_9103,N_8935,N_8834);
nor U9104 (N_9104,N_8864,N_8920);
and U9105 (N_9105,N_8805,N_8921);
xnor U9106 (N_9106,N_8906,N_8786);
xnor U9107 (N_9107,N_8971,N_8911);
and U9108 (N_9108,N_8791,N_8831);
nor U9109 (N_9109,N_8810,N_8907);
nor U9110 (N_9110,N_8930,N_8835);
and U9111 (N_9111,N_8856,N_8854);
and U9112 (N_9112,N_8760,N_8909);
nor U9113 (N_9113,N_8811,N_8777);
and U9114 (N_9114,N_8825,N_8837);
nand U9115 (N_9115,N_8817,N_8762);
nor U9116 (N_9116,N_8818,N_8858);
nand U9117 (N_9117,N_8773,N_8990);
nand U9118 (N_9118,N_8887,N_8830);
nor U9119 (N_9119,N_8848,N_8884);
nand U9120 (N_9120,N_8767,N_8815);
nor U9121 (N_9121,N_8984,N_8944);
and U9122 (N_9122,N_8827,N_8785);
nor U9123 (N_9123,N_8883,N_8775);
or U9124 (N_9124,N_8877,N_8997);
xnor U9125 (N_9125,N_8812,N_8892);
xnor U9126 (N_9126,N_8854,N_8801);
nor U9127 (N_9127,N_8903,N_8909);
and U9128 (N_9128,N_8848,N_8812);
xor U9129 (N_9129,N_8929,N_8975);
nor U9130 (N_9130,N_8961,N_8977);
or U9131 (N_9131,N_8983,N_8984);
and U9132 (N_9132,N_8941,N_8992);
nand U9133 (N_9133,N_8799,N_8879);
and U9134 (N_9134,N_8781,N_8908);
xor U9135 (N_9135,N_8950,N_8824);
nand U9136 (N_9136,N_8981,N_8803);
and U9137 (N_9137,N_8956,N_8844);
nand U9138 (N_9138,N_8799,N_8758);
or U9139 (N_9139,N_8937,N_8951);
or U9140 (N_9140,N_8960,N_8800);
or U9141 (N_9141,N_8951,N_8874);
nor U9142 (N_9142,N_8891,N_8797);
or U9143 (N_9143,N_8776,N_8864);
and U9144 (N_9144,N_8820,N_8941);
nor U9145 (N_9145,N_8798,N_8852);
nor U9146 (N_9146,N_8942,N_8823);
nor U9147 (N_9147,N_8753,N_8940);
nor U9148 (N_9148,N_8991,N_8892);
and U9149 (N_9149,N_8930,N_8933);
and U9150 (N_9150,N_8842,N_8943);
nand U9151 (N_9151,N_8876,N_8754);
nand U9152 (N_9152,N_8913,N_8858);
nor U9153 (N_9153,N_8840,N_8930);
or U9154 (N_9154,N_8937,N_8844);
and U9155 (N_9155,N_8996,N_8987);
nand U9156 (N_9156,N_8985,N_8944);
and U9157 (N_9157,N_8846,N_8803);
or U9158 (N_9158,N_8903,N_8826);
or U9159 (N_9159,N_8813,N_8989);
and U9160 (N_9160,N_8997,N_8876);
nand U9161 (N_9161,N_8965,N_8981);
nand U9162 (N_9162,N_8944,N_8826);
nand U9163 (N_9163,N_8932,N_8792);
nor U9164 (N_9164,N_8935,N_8920);
or U9165 (N_9165,N_8896,N_8990);
nand U9166 (N_9166,N_8807,N_8996);
nor U9167 (N_9167,N_8881,N_8774);
nand U9168 (N_9168,N_8820,N_8759);
and U9169 (N_9169,N_8871,N_8988);
xnor U9170 (N_9170,N_8858,N_8875);
or U9171 (N_9171,N_8939,N_8900);
or U9172 (N_9172,N_8814,N_8996);
nor U9173 (N_9173,N_8967,N_8762);
nor U9174 (N_9174,N_8998,N_8779);
nand U9175 (N_9175,N_8924,N_8843);
and U9176 (N_9176,N_8853,N_8994);
nor U9177 (N_9177,N_8902,N_8801);
nor U9178 (N_9178,N_8896,N_8954);
xnor U9179 (N_9179,N_8859,N_8835);
xnor U9180 (N_9180,N_8930,N_8778);
and U9181 (N_9181,N_8878,N_8852);
nor U9182 (N_9182,N_8946,N_8828);
nand U9183 (N_9183,N_8934,N_8827);
or U9184 (N_9184,N_8900,N_8796);
nor U9185 (N_9185,N_8982,N_8831);
or U9186 (N_9186,N_8809,N_8828);
xnor U9187 (N_9187,N_8778,N_8924);
nand U9188 (N_9188,N_8871,N_8793);
and U9189 (N_9189,N_8854,N_8935);
nand U9190 (N_9190,N_8788,N_8834);
or U9191 (N_9191,N_8798,N_8977);
or U9192 (N_9192,N_8927,N_8857);
nor U9193 (N_9193,N_8862,N_8821);
nand U9194 (N_9194,N_8857,N_8762);
and U9195 (N_9195,N_8843,N_8912);
xnor U9196 (N_9196,N_8993,N_8943);
or U9197 (N_9197,N_8903,N_8906);
nor U9198 (N_9198,N_8866,N_8763);
nor U9199 (N_9199,N_8850,N_8945);
nor U9200 (N_9200,N_8798,N_8978);
or U9201 (N_9201,N_8805,N_8935);
nor U9202 (N_9202,N_8889,N_8867);
and U9203 (N_9203,N_8920,N_8858);
or U9204 (N_9204,N_8984,N_8758);
nor U9205 (N_9205,N_8846,N_8776);
nor U9206 (N_9206,N_8757,N_8991);
or U9207 (N_9207,N_8821,N_8859);
nor U9208 (N_9208,N_8890,N_8764);
nand U9209 (N_9209,N_8891,N_8816);
nand U9210 (N_9210,N_8946,N_8773);
xnor U9211 (N_9211,N_8915,N_8991);
or U9212 (N_9212,N_8965,N_8990);
nor U9213 (N_9213,N_8929,N_8928);
xnor U9214 (N_9214,N_8808,N_8920);
or U9215 (N_9215,N_8886,N_8959);
nor U9216 (N_9216,N_8801,N_8782);
and U9217 (N_9217,N_8868,N_8877);
nand U9218 (N_9218,N_8951,N_8794);
and U9219 (N_9219,N_8882,N_8879);
nor U9220 (N_9220,N_8755,N_8768);
nor U9221 (N_9221,N_8951,N_8876);
nor U9222 (N_9222,N_8961,N_8963);
and U9223 (N_9223,N_8988,N_8838);
and U9224 (N_9224,N_8909,N_8861);
or U9225 (N_9225,N_8892,N_8942);
or U9226 (N_9226,N_8954,N_8932);
nor U9227 (N_9227,N_8771,N_8827);
nor U9228 (N_9228,N_8780,N_8950);
nand U9229 (N_9229,N_8959,N_8767);
and U9230 (N_9230,N_8808,N_8990);
and U9231 (N_9231,N_8829,N_8903);
or U9232 (N_9232,N_8829,N_8831);
nor U9233 (N_9233,N_8818,N_8819);
or U9234 (N_9234,N_8968,N_8896);
nand U9235 (N_9235,N_8911,N_8998);
nand U9236 (N_9236,N_8999,N_8847);
and U9237 (N_9237,N_8811,N_8948);
or U9238 (N_9238,N_8887,N_8820);
or U9239 (N_9239,N_8802,N_8756);
and U9240 (N_9240,N_8884,N_8964);
or U9241 (N_9241,N_8896,N_8902);
nand U9242 (N_9242,N_8832,N_8951);
or U9243 (N_9243,N_8865,N_8828);
or U9244 (N_9244,N_8815,N_8783);
xor U9245 (N_9245,N_8902,N_8915);
nor U9246 (N_9246,N_8909,N_8859);
nor U9247 (N_9247,N_8775,N_8833);
and U9248 (N_9248,N_8772,N_8946);
or U9249 (N_9249,N_8984,N_8971);
and U9250 (N_9250,N_9060,N_9175);
and U9251 (N_9251,N_9165,N_9066);
or U9252 (N_9252,N_9015,N_9181);
nor U9253 (N_9253,N_9187,N_9176);
and U9254 (N_9254,N_9242,N_9231);
xor U9255 (N_9255,N_9012,N_9245);
and U9256 (N_9256,N_9133,N_9134);
xor U9257 (N_9257,N_9020,N_9006);
and U9258 (N_9258,N_9136,N_9026);
or U9259 (N_9259,N_9110,N_9170);
and U9260 (N_9260,N_9236,N_9099);
xor U9261 (N_9261,N_9159,N_9059);
xor U9262 (N_9262,N_9205,N_9149);
nand U9263 (N_9263,N_9085,N_9030);
nand U9264 (N_9264,N_9208,N_9228);
or U9265 (N_9265,N_9109,N_9115);
and U9266 (N_9266,N_9067,N_9218);
or U9267 (N_9267,N_9041,N_9064);
xnor U9268 (N_9268,N_9019,N_9162);
nand U9269 (N_9269,N_9166,N_9148);
nand U9270 (N_9270,N_9068,N_9077);
or U9271 (N_9271,N_9171,N_9223);
or U9272 (N_9272,N_9193,N_9211);
xor U9273 (N_9273,N_9210,N_9018);
nand U9274 (N_9274,N_9044,N_9103);
or U9275 (N_9275,N_9140,N_9076);
and U9276 (N_9276,N_9135,N_9038);
and U9277 (N_9277,N_9229,N_9070);
or U9278 (N_9278,N_9247,N_9189);
nor U9279 (N_9279,N_9074,N_9021);
and U9280 (N_9280,N_9122,N_9197);
nor U9281 (N_9281,N_9111,N_9052);
nand U9282 (N_9282,N_9198,N_9235);
or U9283 (N_9283,N_9057,N_9196);
and U9284 (N_9284,N_9040,N_9091);
nand U9285 (N_9285,N_9100,N_9105);
nor U9286 (N_9286,N_9054,N_9207);
nand U9287 (N_9287,N_9016,N_9062);
and U9288 (N_9288,N_9145,N_9084);
nor U9289 (N_9289,N_9154,N_9241);
and U9290 (N_9290,N_9119,N_9124);
or U9291 (N_9291,N_9232,N_9013);
or U9292 (N_9292,N_9129,N_9095);
and U9293 (N_9293,N_9220,N_9025);
and U9294 (N_9294,N_9024,N_9023);
nor U9295 (N_9295,N_9055,N_9209);
nor U9296 (N_9296,N_9072,N_9155);
nor U9297 (N_9297,N_9081,N_9083);
nand U9298 (N_9298,N_9017,N_9153);
nand U9299 (N_9299,N_9204,N_9001);
nand U9300 (N_9300,N_9195,N_9000);
xnor U9301 (N_9301,N_9061,N_9185);
nand U9302 (N_9302,N_9203,N_9009);
or U9303 (N_9303,N_9174,N_9219);
and U9304 (N_9304,N_9037,N_9182);
nor U9305 (N_9305,N_9128,N_9180);
nand U9306 (N_9306,N_9063,N_9143);
nor U9307 (N_9307,N_9011,N_9173);
and U9308 (N_9308,N_9082,N_9031);
or U9309 (N_9309,N_9049,N_9051);
nand U9310 (N_9310,N_9005,N_9075);
and U9311 (N_9311,N_9249,N_9113);
nand U9312 (N_9312,N_9144,N_9142);
nor U9313 (N_9313,N_9048,N_9169);
nand U9314 (N_9314,N_9215,N_9194);
or U9315 (N_9315,N_9131,N_9088);
and U9316 (N_9316,N_9121,N_9002);
or U9317 (N_9317,N_9087,N_9191);
or U9318 (N_9318,N_9058,N_9032);
and U9319 (N_9319,N_9098,N_9079);
nand U9320 (N_9320,N_9183,N_9114);
and U9321 (N_9321,N_9147,N_9192);
nand U9322 (N_9322,N_9199,N_9086);
nor U9323 (N_9323,N_9106,N_9080);
nand U9324 (N_9324,N_9233,N_9216);
nand U9325 (N_9325,N_9050,N_9188);
nand U9326 (N_9326,N_9108,N_9036);
nand U9327 (N_9327,N_9212,N_9168);
nand U9328 (N_9328,N_9101,N_9238);
nand U9329 (N_9329,N_9078,N_9164);
or U9330 (N_9330,N_9152,N_9008);
or U9331 (N_9331,N_9226,N_9150);
xor U9332 (N_9332,N_9248,N_9034);
nor U9333 (N_9333,N_9112,N_9116);
and U9334 (N_9334,N_9172,N_9027);
xnor U9335 (N_9335,N_9093,N_9132);
or U9336 (N_9336,N_9141,N_9158);
or U9337 (N_9337,N_9123,N_9167);
or U9338 (N_9338,N_9201,N_9222);
or U9339 (N_9339,N_9177,N_9156);
nor U9340 (N_9340,N_9102,N_9225);
and U9341 (N_9341,N_9120,N_9184);
or U9342 (N_9342,N_9043,N_9107);
and U9343 (N_9343,N_9117,N_9073);
and U9344 (N_9344,N_9094,N_9097);
or U9345 (N_9345,N_9039,N_9139);
nor U9346 (N_9346,N_9010,N_9096);
nor U9347 (N_9347,N_9186,N_9089);
nand U9348 (N_9348,N_9157,N_9230);
nand U9349 (N_9349,N_9227,N_9179);
and U9350 (N_9350,N_9178,N_9042);
or U9351 (N_9351,N_9071,N_9090);
nand U9352 (N_9352,N_9033,N_9246);
xor U9353 (N_9353,N_9127,N_9234);
and U9354 (N_9354,N_9007,N_9160);
and U9355 (N_9355,N_9161,N_9190);
nand U9356 (N_9356,N_9126,N_9104);
nor U9357 (N_9357,N_9028,N_9004);
xnor U9358 (N_9358,N_9053,N_9065);
and U9359 (N_9359,N_9224,N_9214);
nor U9360 (N_9360,N_9200,N_9146);
xnor U9361 (N_9361,N_9014,N_9137);
xnor U9362 (N_9362,N_9243,N_9092);
and U9363 (N_9363,N_9118,N_9217);
xor U9364 (N_9364,N_9035,N_9125);
or U9365 (N_9365,N_9151,N_9029);
nor U9366 (N_9366,N_9022,N_9138);
nand U9367 (N_9367,N_9047,N_9130);
and U9368 (N_9368,N_9221,N_9237);
and U9369 (N_9369,N_9239,N_9206);
and U9370 (N_9370,N_9213,N_9056);
and U9371 (N_9371,N_9240,N_9069);
nor U9372 (N_9372,N_9202,N_9046);
or U9373 (N_9373,N_9163,N_9003);
nor U9374 (N_9374,N_9045,N_9244);
and U9375 (N_9375,N_9009,N_9167);
nand U9376 (N_9376,N_9091,N_9203);
nand U9377 (N_9377,N_9111,N_9089);
nand U9378 (N_9378,N_9174,N_9218);
nor U9379 (N_9379,N_9066,N_9062);
and U9380 (N_9380,N_9238,N_9186);
and U9381 (N_9381,N_9095,N_9034);
and U9382 (N_9382,N_9193,N_9158);
or U9383 (N_9383,N_9086,N_9084);
and U9384 (N_9384,N_9017,N_9008);
nor U9385 (N_9385,N_9010,N_9079);
nand U9386 (N_9386,N_9155,N_9181);
nand U9387 (N_9387,N_9087,N_9156);
xnor U9388 (N_9388,N_9070,N_9150);
or U9389 (N_9389,N_9185,N_9225);
nand U9390 (N_9390,N_9043,N_9199);
nand U9391 (N_9391,N_9146,N_9136);
nor U9392 (N_9392,N_9212,N_9163);
xor U9393 (N_9393,N_9003,N_9123);
or U9394 (N_9394,N_9019,N_9054);
nand U9395 (N_9395,N_9154,N_9150);
nor U9396 (N_9396,N_9010,N_9180);
nand U9397 (N_9397,N_9014,N_9124);
and U9398 (N_9398,N_9195,N_9009);
or U9399 (N_9399,N_9046,N_9061);
nor U9400 (N_9400,N_9238,N_9217);
or U9401 (N_9401,N_9009,N_9176);
or U9402 (N_9402,N_9114,N_9034);
nor U9403 (N_9403,N_9141,N_9201);
nand U9404 (N_9404,N_9177,N_9141);
nand U9405 (N_9405,N_9220,N_9227);
or U9406 (N_9406,N_9083,N_9242);
or U9407 (N_9407,N_9024,N_9144);
xnor U9408 (N_9408,N_9154,N_9166);
and U9409 (N_9409,N_9236,N_9083);
and U9410 (N_9410,N_9029,N_9064);
xnor U9411 (N_9411,N_9010,N_9002);
xnor U9412 (N_9412,N_9230,N_9049);
xor U9413 (N_9413,N_9227,N_9032);
or U9414 (N_9414,N_9234,N_9178);
or U9415 (N_9415,N_9088,N_9221);
or U9416 (N_9416,N_9008,N_9103);
nor U9417 (N_9417,N_9163,N_9194);
nand U9418 (N_9418,N_9166,N_9093);
nor U9419 (N_9419,N_9162,N_9243);
nand U9420 (N_9420,N_9240,N_9131);
xnor U9421 (N_9421,N_9185,N_9014);
nand U9422 (N_9422,N_9150,N_9036);
and U9423 (N_9423,N_9065,N_9170);
or U9424 (N_9424,N_9239,N_9006);
and U9425 (N_9425,N_9114,N_9104);
nand U9426 (N_9426,N_9013,N_9045);
nand U9427 (N_9427,N_9018,N_9042);
nor U9428 (N_9428,N_9019,N_9155);
nand U9429 (N_9429,N_9090,N_9113);
nor U9430 (N_9430,N_9194,N_9218);
xnor U9431 (N_9431,N_9170,N_9091);
xnor U9432 (N_9432,N_9145,N_9048);
nor U9433 (N_9433,N_9056,N_9064);
and U9434 (N_9434,N_9162,N_9215);
xor U9435 (N_9435,N_9089,N_9173);
nor U9436 (N_9436,N_9187,N_9045);
nand U9437 (N_9437,N_9044,N_9034);
and U9438 (N_9438,N_9141,N_9166);
or U9439 (N_9439,N_9033,N_9020);
and U9440 (N_9440,N_9121,N_9174);
and U9441 (N_9441,N_9040,N_9206);
or U9442 (N_9442,N_9225,N_9132);
or U9443 (N_9443,N_9055,N_9012);
or U9444 (N_9444,N_9015,N_9243);
nand U9445 (N_9445,N_9241,N_9193);
and U9446 (N_9446,N_9031,N_9191);
nor U9447 (N_9447,N_9125,N_9054);
or U9448 (N_9448,N_9053,N_9060);
nor U9449 (N_9449,N_9238,N_9179);
and U9450 (N_9450,N_9135,N_9162);
or U9451 (N_9451,N_9163,N_9226);
or U9452 (N_9452,N_9202,N_9170);
or U9453 (N_9453,N_9230,N_9106);
and U9454 (N_9454,N_9120,N_9071);
xor U9455 (N_9455,N_9097,N_9061);
nand U9456 (N_9456,N_9085,N_9249);
nand U9457 (N_9457,N_9143,N_9220);
xnor U9458 (N_9458,N_9059,N_9092);
or U9459 (N_9459,N_9041,N_9093);
nor U9460 (N_9460,N_9217,N_9071);
or U9461 (N_9461,N_9081,N_9064);
nand U9462 (N_9462,N_9100,N_9134);
nand U9463 (N_9463,N_9067,N_9057);
xor U9464 (N_9464,N_9049,N_9184);
nand U9465 (N_9465,N_9220,N_9102);
and U9466 (N_9466,N_9079,N_9172);
or U9467 (N_9467,N_9174,N_9136);
and U9468 (N_9468,N_9025,N_9140);
or U9469 (N_9469,N_9166,N_9078);
nand U9470 (N_9470,N_9134,N_9020);
or U9471 (N_9471,N_9097,N_9164);
and U9472 (N_9472,N_9154,N_9053);
nand U9473 (N_9473,N_9153,N_9066);
and U9474 (N_9474,N_9108,N_9178);
xnor U9475 (N_9475,N_9118,N_9087);
or U9476 (N_9476,N_9068,N_9060);
nand U9477 (N_9477,N_9234,N_9041);
or U9478 (N_9478,N_9150,N_9224);
nand U9479 (N_9479,N_9030,N_9072);
or U9480 (N_9480,N_9178,N_9026);
nor U9481 (N_9481,N_9096,N_9166);
and U9482 (N_9482,N_9024,N_9177);
nor U9483 (N_9483,N_9222,N_9045);
nand U9484 (N_9484,N_9126,N_9107);
and U9485 (N_9485,N_9149,N_9104);
nor U9486 (N_9486,N_9089,N_9116);
and U9487 (N_9487,N_9038,N_9243);
nor U9488 (N_9488,N_9234,N_9098);
and U9489 (N_9489,N_9001,N_9075);
and U9490 (N_9490,N_9123,N_9069);
and U9491 (N_9491,N_9207,N_9034);
and U9492 (N_9492,N_9167,N_9195);
nor U9493 (N_9493,N_9170,N_9034);
and U9494 (N_9494,N_9085,N_9023);
nand U9495 (N_9495,N_9001,N_9224);
or U9496 (N_9496,N_9008,N_9237);
nor U9497 (N_9497,N_9135,N_9059);
nor U9498 (N_9498,N_9035,N_9110);
and U9499 (N_9499,N_9202,N_9156);
nor U9500 (N_9500,N_9465,N_9463);
and U9501 (N_9501,N_9278,N_9273);
and U9502 (N_9502,N_9424,N_9279);
nor U9503 (N_9503,N_9306,N_9254);
and U9504 (N_9504,N_9302,N_9420);
nor U9505 (N_9505,N_9417,N_9421);
nand U9506 (N_9506,N_9471,N_9360);
nand U9507 (N_9507,N_9371,N_9381);
nand U9508 (N_9508,N_9475,N_9378);
or U9509 (N_9509,N_9481,N_9297);
nor U9510 (N_9510,N_9310,N_9459);
or U9511 (N_9511,N_9335,N_9439);
and U9512 (N_9512,N_9358,N_9428);
and U9513 (N_9513,N_9396,N_9462);
or U9514 (N_9514,N_9489,N_9487);
and U9515 (N_9515,N_9313,N_9366);
nand U9516 (N_9516,N_9330,N_9458);
xnor U9517 (N_9517,N_9407,N_9447);
or U9518 (N_9518,N_9409,N_9474);
nor U9519 (N_9519,N_9392,N_9427);
xnor U9520 (N_9520,N_9291,N_9426);
and U9521 (N_9521,N_9425,N_9395);
xor U9522 (N_9522,N_9472,N_9325);
or U9523 (N_9523,N_9379,N_9478);
nand U9524 (N_9524,N_9466,N_9293);
xnor U9525 (N_9525,N_9285,N_9422);
nand U9526 (N_9526,N_9446,N_9256);
nand U9527 (N_9527,N_9494,N_9317);
or U9528 (N_9528,N_9434,N_9342);
or U9529 (N_9529,N_9389,N_9391);
nor U9530 (N_9530,N_9467,N_9349);
and U9531 (N_9531,N_9351,N_9345);
nor U9532 (N_9532,N_9418,N_9402);
nand U9533 (N_9533,N_9400,N_9315);
and U9534 (N_9534,N_9377,N_9367);
or U9535 (N_9535,N_9283,N_9333);
and U9536 (N_9536,N_9350,N_9398);
nand U9537 (N_9537,N_9403,N_9269);
and U9538 (N_9538,N_9264,N_9347);
xnor U9539 (N_9539,N_9486,N_9280);
nor U9540 (N_9540,N_9477,N_9271);
nand U9541 (N_9541,N_9448,N_9375);
nand U9542 (N_9542,N_9301,N_9479);
and U9543 (N_9543,N_9493,N_9263);
and U9544 (N_9544,N_9394,N_9414);
or U9545 (N_9545,N_9331,N_9384);
or U9546 (N_9546,N_9296,N_9382);
nor U9547 (N_9547,N_9388,N_9300);
nor U9548 (N_9548,N_9413,N_9326);
or U9549 (N_9549,N_9429,N_9294);
nor U9550 (N_9550,N_9348,N_9309);
or U9551 (N_9551,N_9499,N_9289);
nand U9552 (N_9552,N_9460,N_9488);
and U9553 (N_9553,N_9438,N_9406);
xnor U9554 (N_9554,N_9415,N_9374);
nor U9555 (N_9555,N_9255,N_9468);
nand U9556 (N_9556,N_9482,N_9356);
or U9557 (N_9557,N_9357,N_9383);
xnor U9558 (N_9558,N_9259,N_9364);
nand U9559 (N_9559,N_9473,N_9433);
or U9560 (N_9560,N_9496,N_9485);
nor U9561 (N_9561,N_9453,N_9476);
or U9562 (N_9562,N_9252,N_9292);
nor U9563 (N_9563,N_9362,N_9376);
nor U9564 (N_9564,N_9340,N_9483);
and U9565 (N_9565,N_9451,N_9308);
and U9566 (N_9566,N_9404,N_9265);
nand U9567 (N_9567,N_9341,N_9295);
and U9568 (N_9568,N_9430,N_9272);
nor U9569 (N_9569,N_9305,N_9435);
nor U9570 (N_9570,N_9286,N_9336);
nor U9571 (N_9571,N_9303,N_9282);
and U9572 (N_9572,N_9319,N_9361);
nand U9573 (N_9573,N_9470,N_9443);
nor U9574 (N_9574,N_9284,N_9250);
nor U9575 (N_9575,N_9311,N_9497);
nor U9576 (N_9576,N_9318,N_9492);
xnor U9577 (N_9577,N_9484,N_9346);
or U9578 (N_9578,N_9266,N_9281);
xor U9579 (N_9579,N_9321,N_9440);
nand U9580 (N_9580,N_9449,N_9253);
or U9581 (N_9581,N_9410,N_9495);
and U9582 (N_9582,N_9359,N_9363);
nand U9583 (N_9583,N_9436,N_9257);
and U9584 (N_9584,N_9490,N_9368);
xnor U9585 (N_9585,N_9464,N_9287);
and U9586 (N_9586,N_9299,N_9328);
or U9587 (N_9587,N_9298,N_9498);
nand U9588 (N_9588,N_9397,N_9369);
nor U9589 (N_9589,N_9304,N_9390);
or U9590 (N_9590,N_9314,N_9419);
nor U9591 (N_9591,N_9457,N_9412);
xor U9592 (N_9592,N_9373,N_9445);
or U9593 (N_9593,N_9320,N_9354);
nor U9594 (N_9594,N_9411,N_9260);
nand U9595 (N_9595,N_9307,N_9423);
nor U9596 (N_9596,N_9441,N_9437);
nand U9597 (N_9597,N_9316,N_9431);
nand U9598 (N_9598,N_9324,N_9332);
nand U9599 (N_9599,N_9327,N_9290);
nor U9600 (N_9600,N_9480,N_9416);
xnor U9601 (N_9601,N_9372,N_9393);
or U9602 (N_9602,N_9288,N_9261);
or U9603 (N_9603,N_9267,N_9270);
nor U9604 (N_9604,N_9258,N_9323);
or U9605 (N_9605,N_9405,N_9380);
or U9606 (N_9606,N_9268,N_9343);
nand U9607 (N_9607,N_9385,N_9455);
nand U9608 (N_9608,N_9452,N_9401);
and U9609 (N_9609,N_9275,N_9442);
and U9610 (N_9610,N_9491,N_9352);
and U9611 (N_9611,N_9276,N_9353);
xnor U9612 (N_9612,N_9334,N_9444);
or U9613 (N_9613,N_9344,N_9322);
nor U9614 (N_9614,N_9337,N_9251);
or U9615 (N_9615,N_9312,N_9274);
or U9616 (N_9616,N_9386,N_9262);
or U9617 (N_9617,N_9456,N_9355);
and U9618 (N_9618,N_9432,N_9370);
nor U9619 (N_9619,N_9461,N_9277);
nor U9620 (N_9620,N_9399,N_9365);
nor U9621 (N_9621,N_9469,N_9339);
nand U9622 (N_9622,N_9387,N_9338);
and U9623 (N_9623,N_9329,N_9454);
nand U9624 (N_9624,N_9408,N_9450);
nand U9625 (N_9625,N_9325,N_9347);
nor U9626 (N_9626,N_9324,N_9359);
and U9627 (N_9627,N_9294,N_9463);
nor U9628 (N_9628,N_9360,N_9318);
nor U9629 (N_9629,N_9261,N_9393);
and U9630 (N_9630,N_9450,N_9317);
and U9631 (N_9631,N_9286,N_9401);
nor U9632 (N_9632,N_9383,N_9378);
and U9633 (N_9633,N_9278,N_9488);
nor U9634 (N_9634,N_9258,N_9421);
nand U9635 (N_9635,N_9459,N_9267);
and U9636 (N_9636,N_9357,N_9495);
or U9637 (N_9637,N_9335,N_9387);
or U9638 (N_9638,N_9379,N_9318);
nand U9639 (N_9639,N_9383,N_9399);
nor U9640 (N_9640,N_9439,N_9333);
or U9641 (N_9641,N_9333,N_9463);
or U9642 (N_9642,N_9290,N_9364);
nand U9643 (N_9643,N_9391,N_9337);
nand U9644 (N_9644,N_9386,N_9265);
nand U9645 (N_9645,N_9254,N_9258);
nor U9646 (N_9646,N_9358,N_9380);
and U9647 (N_9647,N_9374,N_9436);
nor U9648 (N_9648,N_9336,N_9362);
or U9649 (N_9649,N_9322,N_9326);
nor U9650 (N_9650,N_9259,N_9387);
and U9651 (N_9651,N_9258,N_9385);
and U9652 (N_9652,N_9462,N_9392);
or U9653 (N_9653,N_9273,N_9261);
nor U9654 (N_9654,N_9497,N_9423);
nor U9655 (N_9655,N_9287,N_9447);
xnor U9656 (N_9656,N_9251,N_9320);
nand U9657 (N_9657,N_9376,N_9378);
nor U9658 (N_9658,N_9404,N_9286);
and U9659 (N_9659,N_9301,N_9409);
or U9660 (N_9660,N_9274,N_9414);
nand U9661 (N_9661,N_9449,N_9417);
nand U9662 (N_9662,N_9356,N_9400);
and U9663 (N_9663,N_9452,N_9250);
and U9664 (N_9664,N_9259,N_9357);
and U9665 (N_9665,N_9365,N_9369);
or U9666 (N_9666,N_9258,N_9280);
nand U9667 (N_9667,N_9389,N_9313);
xnor U9668 (N_9668,N_9282,N_9383);
nor U9669 (N_9669,N_9358,N_9343);
or U9670 (N_9670,N_9402,N_9299);
nor U9671 (N_9671,N_9415,N_9335);
xor U9672 (N_9672,N_9324,N_9277);
or U9673 (N_9673,N_9311,N_9409);
nor U9674 (N_9674,N_9422,N_9479);
or U9675 (N_9675,N_9435,N_9323);
nor U9676 (N_9676,N_9392,N_9273);
nand U9677 (N_9677,N_9446,N_9486);
nand U9678 (N_9678,N_9431,N_9322);
nand U9679 (N_9679,N_9398,N_9371);
nor U9680 (N_9680,N_9295,N_9392);
nor U9681 (N_9681,N_9378,N_9495);
nand U9682 (N_9682,N_9446,N_9436);
and U9683 (N_9683,N_9376,N_9421);
and U9684 (N_9684,N_9431,N_9467);
nand U9685 (N_9685,N_9424,N_9431);
and U9686 (N_9686,N_9487,N_9428);
and U9687 (N_9687,N_9377,N_9358);
and U9688 (N_9688,N_9423,N_9390);
nor U9689 (N_9689,N_9428,N_9412);
nor U9690 (N_9690,N_9341,N_9451);
or U9691 (N_9691,N_9268,N_9445);
nand U9692 (N_9692,N_9289,N_9481);
nand U9693 (N_9693,N_9269,N_9358);
xnor U9694 (N_9694,N_9412,N_9386);
nand U9695 (N_9695,N_9418,N_9320);
or U9696 (N_9696,N_9419,N_9399);
and U9697 (N_9697,N_9327,N_9492);
nand U9698 (N_9698,N_9437,N_9370);
nor U9699 (N_9699,N_9358,N_9267);
and U9700 (N_9700,N_9432,N_9332);
or U9701 (N_9701,N_9310,N_9448);
nor U9702 (N_9702,N_9386,N_9360);
and U9703 (N_9703,N_9422,N_9345);
or U9704 (N_9704,N_9384,N_9375);
nand U9705 (N_9705,N_9279,N_9380);
and U9706 (N_9706,N_9448,N_9467);
nor U9707 (N_9707,N_9347,N_9256);
xor U9708 (N_9708,N_9434,N_9343);
xnor U9709 (N_9709,N_9466,N_9440);
nand U9710 (N_9710,N_9470,N_9410);
nand U9711 (N_9711,N_9444,N_9288);
nor U9712 (N_9712,N_9311,N_9250);
nor U9713 (N_9713,N_9364,N_9275);
and U9714 (N_9714,N_9443,N_9260);
or U9715 (N_9715,N_9465,N_9290);
or U9716 (N_9716,N_9286,N_9258);
xor U9717 (N_9717,N_9437,N_9339);
xor U9718 (N_9718,N_9471,N_9484);
or U9719 (N_9719,N_9399,N_9422);
nor U9720 (N_9720,N_9498,N_9495);
and U9721 (N_9721,N_9344,N_9408);
and U9722 (N_9722,N_9363,N_9272);
xor U9723 (N_9723,N_9353,N_9378);
nand U9724 (N_9724,N_9269,N_9391);
nor U9725 (N_9725,N_9270,N_9309);
nand U9726 (N_9726,N_9495,N_9367);
nand U9727 (N_9727,N_9487,N_9344);
and U9728 (N_9728,N_9282,N_9418);
or U9729 (N_9729,N_9497,N_9388);
xor U9730 (N_9730,N_9372,N_9392);
and U9731 (N_9731,N_9405,N_9390);
nor U9732 (N_9732,N_9440,N_9318);
or U9733 (N_9733,N_9393,N_9389);
nand U9734 (N_9734,N_9288,N_9359);
and U9735 (N_9735,N_9321,N_9445);
or U9736 (N_9736,N_9255,N_9489);
nor U9737 (N_9737,N_9490,N_9373);
and U9738 (N_9738,N_9362,N_9262);
or U9739 (N_9739,N_9447,N_9451);
nor U9740 (N_9740,N_9311,N_9354);
nor U9741 (N_9741,N_9291,N_9469);
and U9742 (N_9742,N_9442,N_9307);
or U9743 (N_9743,N_9447,N_9440);
xor U9744 (N_9744,N_9486,N_9448);
or U9745 (N_9745,N_9337,N_9313);
nor U9746 (N_9746,N_9410,N_9296);
nand U9747 (N_9747,N_9335,N_9449);
and U9748 (N_9748,N_9431,N_9318);
nor U9749 (N_9749,N_9255,N_9351);
or U9750 (N_9750,N_9525,N_9575);
and U9751 (N_9751,N_9743,N_9725);
nand U9752 (N_9752,N_9501,N_9676);
and U9753 (N_9753,N_9744,N_9596);
xor U9754 (N_9754,N_9604,N_9644);
and U9755 (N_9755,N_9564,N_9640);
xor U9756 (N_9756,N_9556,N_9508);
nand U9757 (N_9757,N_9687,N_9610);
xor U9758 (N_9758,N_9648,N_9558);
nand U9759 (N_9759,N_9557,N_9568);
nor U9760 (N_9760,N_9590,N_9745);
xnor U9761 (N_9761,N_9576,N_9598);
nand U9762 (N_9762,N_9573,N_9519);
or U9763 (N_9763,N_9559,N_9711);
or U9764 (N_9764,N_9684,N_9584);
or U9765 (N_9765,N_9714,N_9555);
nor U9766 (N_9766,N_9692,N_9622);
and U9767 (N_9767,N_9732,N_9689);
xor U9768 (N_9768,N_9522,N_9628);
or U9769 (N_9769,N_9641,N_9599);
or U9770 (N_9770,N_9528,N_9589);
or U9771 (N_9771,N_9633,N_9665);
nor U9772 (N_9772,N_9603,N_9629);
and U9773 (N_9773,N_9550,N_9678);
nor U9774 (N_9774,N_9723,N_9693);
xor U9775 (N_9775,N_9746,N_9546);
and U9776 (N_9776,N_9695,N_9616);
or U9777 (N_9777,N_9702,N_9645);
and U9778 (N_9778,N_9668,N_9748);
and U9779 (N_9779,N_9592,N_9554);
nand U9780 (N_9780,N_9682,N_9652);
xnor U9781 (N_9781,N_9654,N_9516);
nor U9782 (N_9782,N_9619,N_9673);
and U9783 (N_9783,N_9587,N_9709);
nand U9784 (N_9784,N_9679,N_9642);
nand U9785 (N_9785,N_9726,N_9620);
nor U9786 (N_9786,N_9552,N_9542);
nand U9787 (N_9787,N_9520,N_9505);
nand U9788 (N_9788,N_9514,N_9515);
xnor U9789 (N_9789,N_9570,N_9696);
and U9790 (N_9790,N_9605,N_9588);
nand U9791 (N_9791,N_9591,N_9563);
and U9792 (N_9792,N_9541,N_9691);
nand U9793 (N_9793,N_9582,N_9722);
nor U9794 (N_9794,N_9670,N_9716);
nand U9795 (N_9795,N_9730,N_9607);
nor U9796 (N_9796,N_9708,N_9567);
xor U9797 (N_9797,N_9649,N_9712);
or U9798 (N_9798,N_9728,N_9735);
and U9799 (N_9799,N_9566,N_9513);
and U9800 (N_9800,N_9600,N_9583);
nand U9801 (N_9801,N_9660,N_9549);
nor U9802 (N_9802,N_9698,N_9710);
xor U9803 (N_9803,N_9720,N_9632);
nand U9804 (N_9804,N_9601,N_9545);
and U9805 (N_9805,N_9639,N_9608);
and U9806 (N_9806,N_9609,N_9635);
or U9807 (N_9807,N_9694,N_9544);
or U9808 (N_9808,N_9718,N_9602);
or U9809 (N_9809,N_9627,N_9580);
or U9810 (N_9810,N_9666,N_9749);
xor U9811 (N_9811,N_9672,N_9656);
or U9812 (N_9812,N_9659,N_9511);
nand U9813 (N_9813,N_9653,N_9675);
nand U9814 (N_9814,N_9500,N_9527);
and U9815 (N_9815,N_9548,N_9727);
nand U9816 (N_9816,N_9502,N_9506);
nand U9817 (N_9817,N_9700,N_9667);
nor U9818 (N_9818,N_9517,N_9724);
nand U9819 (N_9819,N_9569,N_9669);
nor U9820 (N_9820,N_9651,N_9634);
xor U9821 (N_9821,N_9581,N_9734);
or U9822 (N_9822,N_9638,N_9612);
nand U9823 (N_9823,N_9705,N_9657);
nand U9824 (N_9824,N_9621,N_9741);
and U9825 (N_9825,N_9731,N_9536);
or U9826 (N_9826,N_9637,N_9742);
and U9827 (N_9827,N_9613,N_9663);
and U9828 (N_9828,N_9685,N_9719);
or U9829 (N_9829,N_9646,N_9530);
or U9830 (N_9830,N_9717,N_9701);
xnor U9831 (N_9831,N_9579,N_9747);
and U9832 (N_9832,N_9737,N_9699);
nand U9833 (N_9833,N_9538,N_9521);
nand U9834 (N_9834,N_9553,N_9606);
and U9835 (N_9835,N_9560,N_9630);
nand U9836 (N_9836,N_9534,N_9585);
nor U9837 (N_9837,N_9510,N_9594);
or U9838 (N_9838,N_9626,N_9715);
and U9839 (N_9839,N_9540,N_9703);
xor U9840 (N_9840,N_9586,N_9611);
nand U9841 (N_9841,N_9503,N_9738);
nor U9842 (N_9842,N_9671,N_9704);
nand U9843 (N_9843,N_9578,N_9532);
nand U9844 (N_9844,N_9686,N_9680);
or U9845 (N_9845,N_9677,N_9664);
nand U9846 (N_9846,N_9577,N_9662);
xnor U9847 (N_9847,N_9683,N_9650);
nor U9848 (N_9848,N_9547,N_9565);
or U9849 (N_9849,N_9543,N_9661);
or U9850 (N_9850,N_9593,N_9572);
xnor U9851 (N_9851,N_9625,N_9674);
nor U9852 (N_9852,N_9643,N_9531);
nor U9853 (N_9853,N_9658,N_9636);
and U9854 (N_9854,N_9721,N_9507);
or U9855 (N_9855,N_9697,N_9740);
xor U9856 (N_9856,N_9504,N_9618);
nor U9857 (N_9857,N_9551,N_9533);
or U9858 (N_9858,N_9688,N_9733);
nand U9859 (N_9859,N_9707,N_9736);
and U9860 (N_9860,N_9512,N_9537);
xor U9861 (N_9861,N_9655,N_9518);
nor U9862 (N_9862,N_9615,N_9631);
or U9863 (N_9863,N_9523,N_9623);
xnor U9864 (N_9864,N_9561,N_9681);
nor U9865 (N_9865,N_9562,N_9729);
and U9866 (N_9866,N_9647,N_9526);
nor U9867 (N_9867,N_9571,N_9706);
nand U9868 (N_9868,N_9597,N_9539);
and U9869 (N_9869,N_9713,N_9624);
nor U9870 (N_9870,N_9574,N_9535);
or U9871 (N_9871,N_9509,N_9595);
and U9872 (N_9872,N_9524,N_9739);
or U9873 (N_9873,N_9690,N_9617);
nand U9874 (N_9874,N_9529,N_9614);
nand U9875 (N_9875,N_9596,N_9582);
and U9876 (N_9876,N_9591,N_9643);
nor U9877 (N_9877,N_9501,N_9554);
or U9878 (N_9878,N_9519,N_9656);
nor U9879 (N_9879,N_9601,N_9618);
and U9880 (N_9880,N_9631,N_9514);
xnor U9881 (N_9881,N_9664,N_9649);
or U9882 (N_9882,N_9748,N_9664);
nand U9883 (N_9883,N_9667,N_9737);
and U9884 (N_9884,N_9580,N_9592);
or U9885 (N_9885,N_9594,N_9523);
and U9886 (N_9886,N_9713,N_9708);
or U9887 (N_9887,N_9537,N_9536);
nand U9888 (N_9888,N_9733,N_9598);
and U9889 (N_9889,N_9690,N_9542);
nor U9890 (N_9890,N_9721,N_9613);
nor U9891 (N_9891,N_9633,N_9576);
nand U9892 (N_9892,N_9543,N_9734);
nand U9893 (N_9893,N_9637,N_9515);
nand U9894 (N_9894,N_9727,N_9593);
xor U9895 (N_9895,N_9634,N_9595);
or U9896 (N_9896,N_9659,N_9557);
xor U9897 (N_9897,N_9544,N_9556);
or U9898 (N_9898,N_9616,N_9714);
xnor U9899 (N_9899,N_9557,N_9549);
nand U9900 (N_9900,N_9746,N_9620);
and U9901 (N_9901,N_9729,N_9671);
nand U9902 (N_9902,N_9663,N_9694);
or U9903 (N_9903,N_9707,N_9742);
nand U9904 (N_9904,N_9558,N_9737);
nand U9905 (N_9905,N_9704,N_9668);
nor U9906 (N_9906,N_9688,N_9732);
nand U9907 (N_9907,N_9520,N_9540);
nand U9908 (N_9908,N_9568,N_9746);
or U9909 (N_9909,N_9692,N_9734);
xor U9910 (N_9910,N_9600,N_9607);
nand U9911 (N_9911,N_9603,N_9613);
or U9912 (N_9912,N_9630,N_9700);
and U9913 (N_9913,N_9649,N_9505);
nand U9914 (N_9914,N_9678,N_9537);
and U9915 (N_9915,N_9706,N_9730);
or U9916 (N_9916,N_9703,N_9736);
and U9917 (N_9917,N_9682,N_9638);
or U9918 (N_9918,N_9614,N_9735);
and U9919 (N_9919,N_9583,N_9628);
nor U9920 (N_9920,N_9603,N_9610);
xnor U9921 (N_9921,N_9540,N_9560);
nand U9922 (N_9922,N_9603,N_9649);
nor U9923 (N_9923,N_9537,N_9670);
and U9924 (N_9924,N_9711,N_9656);
or U9925 (N_9925,N_9702,N_9623);
nor U9926 (N_9926,N_9554,N_9724);
nor U9927 (N_9927,N_9724,N_9537);
nand U9928 (N_9928,N_9578,N_9559);
nand U9929 (N_9929,N_9740,N_9614);
nand U9930 (N_9930,N_9617,N_9584);
xnor U9931 (N_9931,N_9533,N_9704);
xnor U9932 (N_9932,N_9507,N_9515);
or U9933 (N_9933,N_9609,N_9520);
nand U9934 (N_9934,N_9640,N_9746);
or U9935 (N_9935,N_9640,N_9657);
nor U9936 (N_9936,N_9663,N_9616);
nand U9937 (N_9937,N_9589,N_9609);
and U9938 (N_9938,N_9653,N_9555);
nor U9939 (N_9939,N_9710,N_9740);
or U9940 (N_9940,N_9622,N_9625);
or U9941 (N_9941,N_9616,N_9547);
xnor U9942 (N_9942,N_9745,N_9575);
and U9943 (N_9943,N_9655,N_9730);
nand U9944 (N_9944,N_9721,N_9730);
and U9945 (N_9945,N_9514,N_9551);
xor U9946 (N_9946,N_9720,N_9593);
or U9947 (N_9947,N_9534,N_9711);
and U9948 (N_9948,N_9748,N_9597);
xnor U9949 (N_9949,N_9540,N_9737);
nand U9950 (N_9950,N_9732,N_9615);
nor U9951 (N_9951,N_9621,N_9510);
or U9952 (N_9952,N_9551,N_9691);
and U9953 (N_9953,N_9735,N_9661);
nor U9954 (N_9954,N_9557,N_9556);
xnor U9955 (N_9955,N_9623,N_9584);
xnor U9956 (N_9956,N_9581,N_9572);
nor U9957 (N_9957,N_9627,N_9549);
nand U9958 (N_9958,N_9555,N_9691);
nand U9959 (N_9959,N_9522,N_9615);
or U9960 (N_9960,N_9632,N_9631);
nor U9961 (N_9961,N_9738,N_9591);
nor U9962 (N_9962,N_9646,N_9675);
nor U9963 (N_9963,N_9562,N_9501);
and U9964 (N_9964,N_9512,N_9653);
nand U9965 (N_9965,N_9616,N_9645);
and U9966 (N_9966,N_9524,N_9566);
or U9967 (N_9967,N_9515,N_9573);
nor U9968 (N_9968,N_9628,N_9629);
and U9969 (N_9969,N_9714,N_9550);
or U9970 (N_9970,N_9698,N_9647);
nor U9971 (N_9971,N_9631,N_9691);
nor U9972 (N_9972,N_9546,N_9676);
or U9973 (N_9973,N_9554,N_9500);
nor U9974 (N_9974,N_9700,N_9566);
and U9975 (N_9975,N_9534,N_9685);
and U9976 (N_9976,N_9521,N_9737);
and U9977 (N_9977,N_9667,N_9625);
nor U9978 (N_9978,N_9532,N_9628);
nor U9979 (N_9979,N_9523,N_9566);
and U9980 (N_9980,N_9698,N_9513);
nand U9981 (N_9981,N_9526,N_9672);
nor U9982 (N_9982,N_9552,N_9648);
and U9983 (N_9983,N_9637,N_9562);
and U9984 (N_9984,N_9583,N_9677);
nand U9985 (N_9985,N_9510,N_9631);
and U9986 (N_9986,N_9639,N_9632);
nand U9987 (N_9987,N_9738,N_9560);
nand U9988 (N_9988,N_9728,N_9585);
or U9989 (N_9989,N_9600,N_9700);
and U9990 (N_9990,N_9505,N_9705);
nor U9991 (N_9991,N_9617,N_9716);
nand U9992 (N_9992,N_9611,N_9709);
nand U9993 (N_9993,N_9674,N_9726);
xor U9994 (N_9994,N_9591,N_9535);
xor U9995 (N_9995,N_9575,N_9726);
and U9996 (N_9996,N_9515,N_9693);
nor U9997 (N_9997,N_9573,N_9668);
nor U9998 (N_9998,N_9672,N_9732);
nor U9999 (N_9999,N_9652,N_9648);
or U10000 (N_10000,N_9881,N_9934);
nand U10001 (N_10001,N_9961,N_9972);
nand U10002 (N_10002,N_9774,N_9871);
xnor U10003 (N_10003,N_9791,N_9875);
nor U10004 (N_10004,N_9975,N_9806);
nor U10005 (N_10005,N_9950,N_9983);
and U10006 (N_10006,N_9942,N_9753);
nor U10007 (N_10007,N_9847,N_9785);
or U10008 (N_10008,N_9912,N_9816);
nand U10009 (N_10009,N_9865,N_9789);
nor U10010 (N_10010,N_9897,N_9922);
xor U10011 (N_10011,N_9913,N_9838);
xor U10012 (N_10012,N_9967,N_9958);
xor U10013 (N_10013,N_9925,N_9795);
nand U10014 (N_10014,N_9767,N_9834);
nand U10015 (N_10015,N_9794,N_9969);
nand U10016 (N_10016,N_9797,N_9927);
xor U10017 (N_10017,N_9994,N_9817);
nor U10018 (N_10018,N_9973,N_9829);
or U10019 (N_10019,N_9970,N_9869);
nand U10020 (N_10020,N_9798,N_9810);
nor U10021 (N_10021,N_9888,N_9991);
nor U10022 (N_10022,N_9860,N_9870);
and U10023 (N_10023,N_9779,N_9787);
nand U10024 (N_10024,N_9854,N_9914);
or U10025 (N_10025,N_9840,N_9805);
nand U10026 (N_10026,N_9812,N_9866);
nand U10027 (N_10027,N_9874,N_9986);
and U10028 (N_10028,N_9892,N_9773);
or U10029 (N_10029,N_9857,N_9793);
or U10030 (N_10030,N_9836,N_9832);
or U10031 (N_10031,N_9820,N_9886);
nand U10032 (N_10032,N_9943,N_9759);
and U10033 (N_10033,N_9880,N_9784);
or U10034 (N_10034,N_9781,N_9910);
or U10035 (N_10035,N_9852,N_9786);
nand U10036 (N_10036,N_9824,N_9878);
or U10037 (N_10037,N_9891,N_9826);
and U10038 (N_10038,N_9819,N_9955);
and U10039 (N_10039,N_9960,N_9978);
xor U10040 (N_10040,N_9889,N_9862);
and U10041 (N_10041,N_9867,N_9937);
or U10042 (N_10042,N_9872,N_9989);
nand U10043 (N_10043,N_9936,N_9901);
nand U10044 (N_10044,N_9764,N_9951);
and U10045 (N_10045,N_9837,N_9996);
and U10046 (N_10046,N_9974,N_9772);
or U10047 (N_10047,N_9903,N_9782);
nand U10048 (N_10048,N_9890,N_9775);
and U10049 (N_10049,N_9916,N_9949);
nor U10050 (N_10050,N_9845,N_9761);
xnor U10051 (N_10051,N_9771,N_9863);
and U10052 (N_10052,N_9964,N_9790);
and U10053 (N_10053,N_9939,N_9895);
nand U10054 (N_10054,N_9893,N_9769);
nor U10055 (N_10055,N_9887,N_9944);
and U10056 (N_10056,N_9911,N_9876);
nor U10057 (N_10057,N_9850,N_9777);
and U10058 (N_10058,N_9873,N_9899);
nor U10059 (N_10059,N_9923,N_9938);
nand U10060 (N_10060,N_9930,N_9858);
or U10061 (N_10061,N_9807,N_9990);
nor U10062 (N_10062,N_9956,N_9885);
nor U10063 (N_10063,N_9953,N_9813);
or U10064 (N_10064,N_9750,N_9844);
nor U10065 (N_10065,N_9906,N_9855);
xnor U10066 (N_10066,N_9754,N_9940);
nand U10067 (N_10067,N_9780,N_9999);
and U10068 (N_10068,N_9825,N_9859);
or U10069 (N_10069,N_9918,N_9921);
nand U10070 (N_10070,N_9988,N_9904);
or U10071 (N_10071,N_9846,N_9919);
or U10072 (N_10072,N_9755,N_9981);
xor U10073 (N_10073,N_9952,N_9751);
or U10074 (N_10074,N_9830,N_9868);
nor U10075 (N_10075,N_9997,N_9811);
nor U10076 (N_10076,N_9979,N_9962);
nor U10077 (N_10077,N_9948,N_9799);
nand U10078 (N_10078,N_9987,N_9947);
or U10079 (N_10079,N_9849,N_9941);
nand U10080 (N_10080,N_9915,N_9856);
nor U10081 (N_10081,N_9841,N_9800);
nor U10082 (N_10082,N_9851,N_9758);
nand U10083 (N_10083,N_9905,N_9843);
and U10084 (N_10084,N_9765,N_9926);
nand U10085 (N_10085,N_9877,N_9762);
nor U10086 (N_10086,N_9792,N_9833);
xnor U10087 (N_10087,N_9760,N_9884);
nand U10088 (N_10088,N_9928,N_9957);
or U10089 (N_10089,N_9965,N_9803);
and U10090 (N_10090,N_9931,N_9924);
nor U10091 (N_10091,N_9752,N_9900);
nand U10092 (N_10092,N_9823,N_9985);
or U10093 (N_10093,N_9776,N_9980);
xor U10094 (N_10094,N_9932,N_9842);
nand U10095 (N_10095,N_9963,N_9982);
or U10096 (N_10096,N_9818,N_9853);
and U10097 (N_10097,N_9883,N_9882);
xnor U10098 (N_10098,N_9766,N_9801);
or U10099 (N_10099,N_9796,N_9821);
xnor U10100 (N_10100,N_9768,N_9809);
xor U10101 (N_10101,N_9802,N_9822);
nor U10102 (N_10102,N_9839,N_9848);
nand U10103 (N_10103,N_9907,N_9946);
or U10104 (N_10104,N_9879,N_9827);
or U10105 (N_10105,N_9770,N_9971);
nand U10106 (N_10106,N_9917,N_9788);
or U10107 (N_10107,N_9783,N_9815);
xnor U10108 (N_10108,N_9976,N_9828);
and U10109 (N_10109,N_9808,N_9756);
nand U10110 (N_10110,N_9835,N_9757);
and U10111 (N_10111,N_9933,N_9992);
or U10112 (N_10112,N_9993,N_9763);
or U10113 (N_10113,N_9898,N_9909);
or U10114 (N_10114,N_9804,N_9908);
nand U10115 (N_10115,N_9814,N_9831);
nor U10116 (N_10116,N_9920,N_9959);
nand U10117 (N_10117,N_9778,N_9902);
nor U10118 (N_10118,N_9864,N_9977);
nor U10119 (N_10119,N_9998,N_9984);
nor U10120 (N_10120,N_9968,N_9935);
or U10121 (N_10121,N_9966,N_9945);
xnor U10122 (N_10122,N_9861,N_9896);
or U10123 (N_10123,N_9995,N_9894);
and U10124 (N_10124,N_9954,N_9929);
nor U10125 (N_10125,N_9911,N_9906);
nand U10126 (N_10126,N_9857,N_9827);
or U10127 (N_10127,N_9842,N_9874);
nor U10128 (N_10128,N_9942,N_9997);
or U10129 (N_10129,N_9772,N_9924);
and U10130 (N_10130,N_9766,N_9885);
nand U10131 (N_10131,N_9761,N_9916);
nor U10132 (N_10132,N_9936,N_9867);
xnor U10133 (N_10133,N_9797,N_9811);
or U10134 (N_10134,N_9939,N_9757);
nor U10135 (N_10135,N_9842,N_9817);
nand U10136 (N_10136,N_9967,N_9871);
and U10137 (N_10137,N_9986,N_9816);
and U10138 (N_10138,N_9819,N_9925);
and U10139 (N_10139,N_9932,N_9927);
nand U10140 (N_10140,N_9885,N_9973);
and U10141 (N_10141,N_9949,N_9924);
and U10142 (N_10142,N_9916,N_9977);
nand U10143 (N_10143,N_9982,N_9835);
and U10144 (N_10144,N_9999,N_9975);
xor U10145 (N_10145,N_9971,N_9906);
nor U10146 (N_10146,N_9991,N_9795);
nor U10147 (N_10147,N_9819,N_9764);
nand U10148 (N_10148,N_9934,N_9965);
nand U10149 (N_10149,N_9765,N_9780);
and U10150 (N_10150,N_9938,N_9979);
and U10151 (N_10151,N_9820,N_9878);
and U10152 (N_10152,N_9997,N_9774);
nand U10153 (N_10153,N_9883,N_9942);
nor U10154 (N_10154,N_9983,N_9770);
and U10155 (N_10155,N_9998,N_9873);
xnor U10156 (N_10156,N_9783,N_9968);
and U10157 (N_10157,N_9990,N_9853);
nor U10158 (N_10158,N_9763,N_9917);
nand U10159 (N_10159,N_9937,N_9968);
and U10160 (N_10160,N_9852,N_9913);
nor U10161 (N_10161,N_9831,N_9897);
nor U10162 (N_10162,N_9759,N_9890);
nand U10163 (N_10163,N_9941,N_9895);
nand U10164 (N_10164,N_9970,N_9901);
and U10165 (N_10165,N_9835,N_9934);
or U10166 (N_10166,N_9757,N_9982);
nor U10167 (N_10167,N_9868,N_9816);
and U10168 (N_10168,N_9837,N_9914);
and U10169 (N_10169,N_9807,N_9996);
nand U10170 (N_10170,N_9764,N_9989);
or U10171 (N_10171,N_9805,N_9821);
nor U10172 (N_10172,N_9821,N_9884);
nor U10173 (N_10173,N_9905,N_9962);
and U10174 (N_10174,N_9847,N_9826);
and U10175 (N_10175,N_9919,N_9817);
nor U10176 (N_10176,N_9825,N_9879);
nor U10177 (N_10177,N_9810,N_9894);
or U10178 (N_10178,N_9878,N_9943);
and U10179 (N_10179,N_9929,N_9827);
or U10180 (N_10180,N_9773,N_9781);
xnor U10181 (N_10181,N_9810,N_9880);
or U10182 (N_10182,N_9840,N_9972);
and U10183 (N_10183,N_9872,N_9878);
nor U10184 (N_10184,N_9793,N_9751);
nand U10185 (N_10185,N_9795,N_9993);
and U10186 (N_10186,N_9772,N_9914);
nand U10187 (N_10187,N_9847,N_9800);
and U10188 (N_10188,N_9750,N_9955);
or U10189 (N_10189,N_9787,N_9834);
and U10190 (N_10190,N_9910,N_9951);
nand U10191 (N_10191,N_9854,N_9941);
or U10192 (N_10192,N_9807,N_9898);
nand U10193 (N_10193,N_9847,N_9881);
or U10194 (N_10194,N_9788,N_9767);
nor U10195 (N_10195,N_9776,N_9920);
nand U10196 (N_10196,N_9857,N_9831);
or U10197 (N_10197,N_9834,N_9944);
nor U10198 (N_10198,N_9793,N_9846);
nand U10199 (N_10199,N_9801,N_9864);
or U10200 (N_10200,N_9980,N_9979);
or U10201 (N_10201,N_9846,N_9806);
nor U10202 (N_10202,N_9885,N_9752);
nor U10203 (N_10203,N_9822,N_9781);
or U10204 (N_10204,N_9905,N_9902);
or U10205 (N_10205,N_9901,N_9758);
and U10206 (N_10206,N_9944,N_9752);
xnor U10207 (N_10207,N_9809,N_9783);
nand U10208 (N_10208,N_9894,N_9848);
or U10209 (N_10209,N_9890,N_9812);
or U10210 (N_10210,N_9886,N_9985);
and U10211 (N_10211,N_9844,N_9992);
nor U10212 (N_10212,N_9932,N_9794);
xor U10213 (N_10213,N_9827,N_9753);
and U10214 (N_10214,N_9904,N_9854);
nor U10215 (N_10215,N_9833,N_9996);
or U10216 (N_10216,N_9952,N_9979);
or U10217 (N_10217,N_9831,N_9770);
xnor U10218 (N_10218,N_9776,N_9985);
nand U10219 (N_10219,N_9759,N_9827);
nor U10220 (N_10220,N_9963,N_9940);
or U10221 (N_10221,N_9937,N_9843);
nor U10222 (N_10222,N_9907,N_9756);
and U10223 (N_10223,N_9833,N_9900);
nand U10224 (N_10224,N_9974,N_9946);
nand U10225 (N_10225,N_9763,N_9890);
nor U10226 (N_10226,N_9803,N_9851);
or U10227 (N_10227,N_9990,N_9965);
or U10228 (N_10228,N_9948,N_9884);
or U10229 (N_10229,N_9954,N_9751);
nor U10230 (N_10230,N_9759,N_9965);
nand U10231 (N_10231,N_9961,N_9840);
xnor U10232 (N_10232,N_9921,N_9864);
nor U10233 (N_10233,N_9760,N_9861);
nand U10234 (N_10234,N_9849,N_9830);
and U10235 (N_10235,N_9892,N_9775);
nor U10236 (N_10236,N_9794,N_9940);
nand U10237 (N_10237,N_9960,N_9820);
nand U10238 (N_10238,N_9847,N_9860);
and U10239 (N_10239,N_9764,N_9900);
or U10240 (N_10240,N_9975,N_9974);
or U10241 (N_10241,N_9963,N_9911);
and U10242 (N_10242,N_9779,N_9808);
nor U10243 (N_10243,N_9762,N_9872);
or U10244 (N_10244,N_9938,N_9818);
nor U10245 (N_10245,N_9924,N_9778);
or U10246 (N_10246,N_9924,N_9919);
nor U10247 (N_10247,N_9958,N_9815);
or U10248 (N_10248,N_9919,N_9931);
and U10249 (N_10249,N_9929,N_9752);
nor U10250 (N_10250,N_10030,N_10123);
nand U10251 (N_10251,N_10152,N_10242);
xnor U10252 (N_10252,N_10246,N_10221);
and U10253 (N_10253,N_10230,N_10126);
or U10254 (N_10254,N_10228,N_10143);
nor U10255 (N_10255,N_10209,N_10102);
nor U10256 (N_10256,N_10089,N_10031);
xnor U10257 (N_10257,N_10138,N_10099);
or U10258 (N_10258,N_10176,N_10136);
nor U10259 (N_10259,N_10021,N_10182);
xnor U10260 (N_10260,N_10186,N_10225);
and U10261 (N_10261,N_10233,N_10129);
or U10262 (N_10262,N_10032,N_10160);
and U10263 (N_10263,N_10241,N_10144);
and U10264 (N_10264,N_10245,N_10148);
and U10265 (N_10265,N_10005,N_10055);
nor U10266 (N_10266,N_10057,N_10170);
and U10267 (N_10267,N_10014,N_10208);
nand U10268 (N_10268,N_10219,N_10147);
or U10269 (N_10269,N_10192,N_10217);
nor U10270 (N_10270,N_10153,N_10053);
nand U10271 (N_10271,N_10213,N_10082);
and U10272 (N_10272,N_10194,N_10211);
and U10273 (N_10273,N_10220,N_10068);
nor U10274 (N_10274,N_10066,N_10052);
nor U10275 (N_10275,N_10157,N_10028);
or U10276 (N_10276,N_10205,N_10218);
nor U10277 (N_10277,N_10238,N_10172);
and U10278 (N_10278,N_10222,N_10076);
nor U10279 (N_10279,N_10096,N_10134);
and U10280 (N_10280,N_10164,N_10146);
or U10281 (N_10281,N_10046,N_10008);
or U10282 (N_10282,N_10114,N_10229);
nor U10283 (N_10283,N_10119,N_10059);
and U10284 (N_10284,N_10034,N_10051);
or U10285 (N_10285,N_10110,N_10079);
nand U10286 (N_10286,N_10179,N_10072);
nor U10287 (N_10287,N_10124,N_10036);
nand U10288 (N_10288,N_10169,N_10161);
nand U10289 (N_10289,N_10120,N_10177);
and U10290 (N_10290,N_10127,N_10184);
nor U10291 (N_10291,N_10197,N_10084);
and U10292 (N_10292,N_10181,N_10216);
and U10293 (N_10293,N_10024,N_10029);
nor U10294 (N_10294,N_10044,N_10087);
xor U10295 (N_10295,N_10105,N_10166);
nor U10296 (N_10296,N_10163,N_10049);
nor U10297 (N_10297,N_10133,N_10188);
or U10298 (N_10298,N_10178,N_10113);
and U10299 (N_10299,N_10063,N_10204);
and U10300 (N_10300,N_10012,N_10131);
or U10301 (N_10301,N_10141,N_10198);
or U10302 (N_10302,N_10137,N_10065);
or U10303 (N_10303,N_10135,N_10060);
nand U10304 (N_10304,N_10115,N_10041);
nand U10305 (N_10305,N_10023,N_10185);
nand U10306 (N_10306,N_10097,N_10085);
or U10307 (N_10307,N_10202,N_10042);
nand U10308 (N_10308,N_10165,N_10022);
nor U10309 (N_10309,N_10103,N_10086);
nand U10310 (N_10310,N_10168,N_10003);
nand U10311 (N_10311,N_10104,N_10016);
nand U10312 (N_10312,N_10149,N_10158);
nor U10313 (N_10313,N_10173,N_10159);
and U10314 (N_10314,N_10155,N_10037);
and U10315 (N_10315,N_10234,N_10237);
nor U10316 (N_10316,N_10156,N_10154);
nor U10317 (N_10317,N_10027,N_10100);
nor U10318 (N_10318,N_10074,N_10018);
and U10319 (N_10319,N_10067,N_10017);
and U10320 (N_10320,N_10081,N_10191);
nor U10321 (N_10321,N_10092,N_10002);
and U10322 (N_10322,N_10019,N_10175);
and U10323 (N_10323,N_10050,N_10171);
nand U10324 (N_10324,N_10212,N_10224);
or U10325 (N_10325,N_10020,N_10078);
nand U10326 (N_10326,N_10232,N_10064);
nor U10327 (N_10327,N_10010,N_10247);
nor U10328 (N_10328,N_10062,N_10015);
or U10329 (N_10329,N_10145,N_10235);
and U10330 (N_10330,N_10132,N_10203);
nor U10331 (N_10331,N_10244,N_10004);
xor U10332 (N_10332,N_10201,N_10236);
or U10333 (N_10333,N_10026,N_10193);
nand U10334 (N_10334,N_10006,N_10118);
and U10335 (N_10335,N_10125,N_10071);
and U10336 (N_10336,N_10190,N_10095);
or U10337 (N_10337,N_10207,N_10174);
nand U10338 (N_10338,N_10223,N_10248);
xor U10339 (N_10339,N_10094,N_10199);
and U10340 (N_10340,N_10112,N_10226);
and U10341 (N_10341,N_10070,N_10195);
or U10342 (N_10342,N_10215,N_10206);
or U10343 (N_10343,N_10107,N_10054);
nor U10344 (N_10344,N_10239,N_10214);
nor U10345 (N_10345,N_10189,N_10128);
or U10346 (N_10346,N_10035,N_10000);
nor U10347 (N_10347,N_10162,N_10009);
xor U10348 (N_10348,N_10249,N_10243);
nor U10349 (N_10349,N_10069,N_10038);
or U10350 (N_10350,N_10098,N_10045);
or U10351 (N_10351,N_10196,N_10101);
nand U10352 (N_10352,N_10056,N_10040);
and U10353 (N_10353,N_10061,N_10077);
nand U10354 (N_10354,N_10075,N_10183);
or U10355 (N_10355,N_10043,N_10231);
xnor U10356 (N_10356,N_10058,N_10109);
nand U10357 (N_10357,N_10142,N_10073);
and U10358 (N_10358,N_10033,N_10150);
xnor U10359 (N_10359,N_10227,N_10106);
nand U10360 (N_10360,N_10151,N_10090);
nor U10361 (N_10361,N_10240,N_10140);
nand U10362 (N_10362,N_10083,N_10130);
and U10363 (N_10363,N_10111,N_10048);
nand U10364 (N_10364,N_10108,N_10025);
nand U10365 (N_10365,N_10091,N_10122);
and U10366 (N_10366,N_10047,N_10200);
and U10367 (N_10367,N_10093,N_10187);
nor U10368 (N_10368,N_10001,N_10039);
nand U10369 (N_10369,N_10088,N_10210);
and U10370 (N_10370,N_10167,N_10117);
or U10371 (N_10371,N_10116,N_10080);
nand U10372 (N_10372,N_10013,N_10121);
or U10373 (N_10373,N_10007,N_10180);
nor U10374 (N_10374,N_10139,N_10011);
and U10375 (N_10375,N_10212,N_10081);
nand U10376 (N_10376,N_10145,N_10233);
nand U10377 (N_10377,N_10063,N_10097);
nor U10378 (N_10378,N_10020,N_10199);
and U10379 (N_10379,N_10055,N_10020);
nand U10380 (N_10380,N_10228,N_10122);
xor U10381 (N_10381,N_10204,N_10247);
nor U10382 (N_10382,N_10014,N_10029);
and U10383 (N_10383,N_10167,N_10228);
and U10384 (N_10384,N_10009,N_10153);
and U10385 (N_10385,N_10121,N_10206);
and U10386 (N_10386,N_10156,N_10104);
nand U10387 (N_10387,N_10247,N_10196);
or U10388 (N_10388,N_10227,N_10161);
and U10389 (N_10389,N_10124,N_10235);
nor U10390 (N_10390,N_10143,N_10069);
xor U10391 (N_10391,N_10176,N_10108);
and U10392 (N_10392,N_10007,N_10223);
or U10393 (N_10393,N_10122,N_10106);
nand U10394 (N_10394,N_10119,N_10104);
nand U10395 (N_10395,N_10148,N_10055);
nand U10396 (N_10396,N_10146,N_10031);
nand U10397 (N_10397,N_10126,N_10184);
or U10398 (N_10398,N_10135,N_10096);
nand U10399 (N_10399,N_10182,N_10124);
or U10400 (N_10400,N_10232,N_10091);
and U10401 (N_10401,N_10135,N_10103);
nor U10402 (N_10402,N_10026,N_10135);
nand U10403 (N_10403,N_10045,N_10033);
nor U10404 (N_10404,N_10072,N_10224);
nand U10405 (N_10405,N_10064,N_10121);
or U10406 (N_10406,N_10107,N_10048);
nor U10407 (N_10407,N_10219,N_10114);
xnor U10408 (N_10408,N_10030,N_10037);
and U10409 (N_10409,N_10002,N_10248);
nand U10410 (N_10410,N_10152,N_10050);
xor U10411 (N_10411,N_10111,N_10131);
or U10412 (N_10412,N_10147,N_10052);
and U10413 (N_10413,N_10139,N_10138);
xor U10414 (N_10414,N_10156,N_10172);
and U10415 (N_10415,N_10209,N_10065);
or U10416 (N_10416,N_10036,N_10044);
and U10417 (N_10417,N_10131,N_10106);
and U10418 (N_10418,N_10000,N_10127);
and U10419 (N_10419,N_10029,N_10235);
nand U10420 (N_10420,N_10174,N_10021);
nor U10421 (N_10421,N_10180,N_10175);
nand U10422 (N_10422,N_10139,N_10140);
or U10423 (N_10423,N_10187,N_10177);
and U10424 (N_10424,N_10129,N_10046);
nor U10425 (N_10425,N_10125,N_10237);
xnor U10426 (N_10426,N_10230,N_10189);
xor U10427 (N_10427,N_10130,N_10116);
or U10428 (N_10428,N_10011,N_10103);
or U10429 (N_10429,N_10189,N_10022);
nand U10430 (N_10430,N_10239,N_10081);
or U10431 (N_10431,N_10040,N_10150);
nor U10432 (N_10432,N_10023,N_10243);
xor U10433 (N_10433,N_10178,N_10097);
and U10434 (N_10434,N_10217,N_10193);
and U10435 (N_10435,N_10167,N_10021);
and U10436 (N_10436,N_10102,N_10016);
nand U10437 (N_10437,N_10060,N_10196);
and U10438 (N_10438,N_10175,N_10091);
or U10439 (N_10439,N_10193,N_10135);
xnor U10440 (N_10440,N_10193,N_10030);
xor U10441 (N_10441,N_10194,N_10229);
nor U10442 (N_10442,N_10217,N_10060);
or U10443 (N_10443,N_10162,N_10064);
nor U10444 (N_10444,N_10202,N_10146);
or U10445 (N_10445,N_10151,N_10184);
xnor U10446 (N_10446,N_10166,N_10172);
nand U10447 (N_10447,N_10075,N_10021);
nor U10448 (N_10448,N_10144,N_10103);
nand U10449 (N_10449,N_10207,N_10057);
and U10450 (N_10450,N_10225,N_10153);
and U10451 (N_10451,N_10188,N_10061);
and U10452 (N_10452,N_10149,N_10037);
and U10453 (N_10453,N_10049,N_10065);
and U10454 (N_10454,N_10191,N_10072);
or U10455 (N_10455,N_10082,N_10119);
or U10456 (N_10456,N_10032,N_10187);
and U10457 (N_10457,N_10186,N_10188);
and U10458 (N_10458,N_10122,N_10192);
nor U10459 (N_10459,N_10238,N_10248);
nand U10460 (N_10460,N_10122,N_10243);
nand U10461 (N_10461,N_10144,N_10023);
or U10462 (N_10462,N_10019,N_10127);
nand U10463 (N_10463,N_10210,N_10221);
or U10464 (N_10464,N_10227,N_10000);
or U10465 (N_10465,N_10113,N_10067);
or U10466 (N_10466,N_10103,N_10247);
and U10467 (N_10467,N_10224,N_10002);
nand U10468 (N_10468,N_10066,N_10094);
nor U10469 (N_10469,N_10207,N_10242);
and U10470 (N_10470,N_10030,N_10240);
nand U10471 (N_10471,N_10191,N_10046);
nand U10472 (N_10472,N_10226,N_10125);
nor U10473 (N_10473,N_10248,N_10201);
and U10474 (N_10474,N_10215,N_10142);
or U10475 (N_10475,N_10052,N_10074);
xor U10476 (N_10476,N_10217,N_10178);
and U10477 (N_10477,N_10162,N_10105);
nor U10478 (N_10478,N_10013,N_10052);
and U10479 (N_10479,N_10165,N_10234);
nor U10480 (N_10480,N_10155,N_10099);
nand U10481 (N_10481,N_10186,N_10223);
xnor U10482 (N_10482,N_10155,N_10041);
nand U10483 (N_10483,N_10173,N_10109);
and U10484 (N_10484,N_10181,N_10076);
nand U10485 (N_10485,N_10011,N_10085);
and U10486 (N_10486,N_10104,N_10024);
and U10487 (N_10487,N_10197,N_10206);
and U10488 (N_10488,N_10086,N_10088);
and U10489 (N_10489,N_10054,N_10026);
and U10490 (N_10490,N_10010,N_10074);
nand U10491 (N_10491,N_10020,N_10119);
nor U10492 (N_10492,N_10202,N_10097);
and U10493 (N_10493,N_10130,N_10047);
xor U10494 (N_10494,N_10221,N_10178);
nor U10495 (N_10495,N_10079,N_10058);
or U10496 (N_10496,N_10192,N_10006);
xor U10497 (N_10497,N_10091,N_10161);
or U10498 (N_10498,N_10008,N_10049);
nor U10499 (N_10499,N_10200,N_10227);
nor U10500 (N_10500,N_10370,N_10489);
nor U10501 (N_10501,N_10371,N_10264);
xor U10502 (N_10502,N_10494,N_10275);
or U10503 (N_10503,N_10331,N_10480);
and U10504 (N_10504,N_10254,N_10394);
and U10505 (N_10505,N_10265,N_10399);
nor U10506 (N_10506,N_10352,N_10343);
nand U10507 (N_10507,N_10474,N_10281);
and U10508 (N_10508,N_10487,N_10409);
nor U10509 (N_10509,N_10391,N_10266);
or U10510 (N_10510,N_10448,N_10450);
nand U10511 (N_10511,N_10419,N_10303);
nor U10512 (N_10512,N_10460,N_10307);
nand U10513 (N_10513,N_10311,N_10459);
nor U10514 (N_10514,N_10478,N_10455);
or U10515 (N_10515,N_10288,N_10356);
or U10516 (N_10516,N_10403,N_10358);
and U10517 (N_10517,N_10386,N_10464);
nand U10518 (N_10518,N_10338,N_10385);
xor U10519 (N_10519,N_10492,N_10421);
nand U10520 (N_10520,N_10351,N_10317);
or U10521 (N_10521,N_10287,N_10484);
xnor U10522 (N_10522,N_10363,N_10458);
nor U10523 (N_10523,N_10270,N_10262);
xnor U10524 (N_10524,N_10446,N_10482);
or U10525 (N_10525,N_10252,N_10430);
or U10526 (N_10526,N_10420,N_10435);
nand U10527 (N_10527,N_10332,N_10250);
xor U10528 (N_10528,N_10471,N_10470);
and U10529 (N_10529,N_10289,N_10309);
nor U10530 (N_10530,N_10342,N_10360);
nor U10531 (N_10531,N_10441,N_10427);
and U10532 (N_10532,N_10497,N_10279);
and U10533 (N_10533,N_10490,N_10477);
xnor U10534 (N_10534,N_10318,N_10473);
nand U10535 (N_10535,N_10353,N_10326);
nor U10536 (N_10536,N_10321,N_10278);
nor U10537 (N_10537,N_10373,N_10268);
or U10538 (N_10538,N_10379,N_10443);
and U10539 (N_10539,N_10397,N_10453);
or U10540 (N_10540,N_10390,N_10447);
nor U10541 (N_10541,N_10328,N_10368);
nand U10542 (N_10542,N_10369,N_10322);
nand U10543 (N_10543,N_10323,N_10271);
or U10544 (N_10544,N_10407,N_10283);
and U10545 (N_10545,N_10451,N_10334);
nand U10546 (N_10546,N_10292,N_10260);
or U10547 (N_10547,N_10413,N_10395);
and U10548 (N_10548,N_10468,N_10344);
or U10549 (N_10549,N_10272,N_10364);
or U10550 (N_10550,N_10423,N_10383);
nand U10551 (N_10551,N_10357,N_10298);
nand U10552 (N_10552,N_10417,N_10434);
and U10553 (N_10553,N_10496,N_10336);
and U10554 (N_10554,N_10382,N_10469);
xor U10555 (N_10555,N_10428,N_10256);
or U10556 (N_10556,N_10493,N_10324);
nand U10557 (N_10557,N_10401,N_10274);
nor U10558 (N_10558,N_10315,N_10433);
or U10559 (N_10559,N_10376,N_10329);
or U10560 (N_10560,N_10426,N_10301);
nand U10561 (N_10561,N_10491,N_10257);
nand U10562 (N_10562,N_10296,N_10498);
nand U10563 (N_10563,N_10280,N_10365);
and U10564 (N_10564,N_10285,N_10463);
xor U10565 (N_10565,N_10346,N_10452);
and U10566 (N_10566,N_10359,N_10253);
nor U10567 (N_10567,N_10405,N_10400);
and U10568 (N_10568,N_10372,N_10442);
and U10569 (N_10569,N_10294,N_10313);
nand U10570 (N_10570,N_10389,N_10340);
nand U10571 (N_10571,N_10422,N_10415);
and U10572 (N_10572,N_10466,N_10263);
and U10573 (N_10573,N_10362,N_10416);
or U10574 (N_10574,N_10361,N_10472);
nand U10575 (N_10575,N_10412,N_10457);
or U10576 (N_10576,N_10374,N_10339);
nand U10577 (N_10577,N_10461,N_10402);
nor U10578 (N_10578,N_10377,N_10330);
or U10579 (N_10579,N_10411,N_10388);
nand U10580 (N_10580,N_10258,N_10485);
or U10581 (N_10581,N_10319,N_10424);
and U10582 (N_10582,N_10320,N_10345);
nand U10583 (N_10583,N_10341,N_10312);
and U10584 (N_10584,N_10425,N_10445);
nand U10585 (N_10585,N_10302,N_10436);
nor U10586 (N_10586,N_10380,N_10475);
nor U10587 (N_10587,N_10337,N_10290);
nand U10588 (N_10588,N_10483,N_10310);
nor U10589 (N_10589,N_10444,N_10387);
nand U10590 (N_10590,N_10308,N_10404);
nand U10591 (N_10591,N_10462,N_10479);
and U10592 (N_10592,N_10325,N_10261);
nand U10593 (N_10593,N_10454,N_10486);
nand U10594 (N_10594,N_10354,N_10476);
or U10595 (N_10595,N_10393,N_10297);
nor U10596 (N_10596,N_10384,N_10295);
or U10597 (N_10597,N_10282,N_10381);
xnor U10598 (N_10598,N_10286,N_10251);
or U10599 (N_10599,N_10437,N_10293);
xor U10600 (N_10600,N_10378,N_10366);
xor U10601 (N_10601,N_10429,N_10355);
or U10602 (N_10602,N_10255,N_10414);
and U10603 (N_10603,N_10299,N_10467);
and U10604 (N_10604,N_10488,N_10408);
nor U10605 (N_10605,N_10305,N_10335);
xnor U10606 (N_10606,N_10350,N_10277);
or U10607 (N_10607,N_10300,N_10398);
nand U10608 (N_10608,N_10269,N_10259);
and U10609 (N_10609,N_10284,N_10481);
or U10610 (N_10610,N_10327,N_10449);
nand U10611 (N_10611,N_10333,N_10316);
nand U10612 (N_10612,N_10273,N_10406);
nor U10613 (N_10613,N_10410,N_10314);
xnor U10614 (N_10614,N_10347,N_10349);
nand U10615 (N_10615,N_10375,N_10267);
nor U10616 (N_10616,N_10456,N_10438);
nand U10617 (N_10617,N_10465,N_10392);
or U10618 (N_10618,N_10495,N_10499);
and U10619 (N_10619,N_10367,N_10439);
nand U10620 (N_10620,N_10291,N_10418);
and U10621 (N_10621,N_10276,N_10396);
or U10622 (N_10622,N_10306,N_10304);
xor U10623 (N_10623,N_10432,N_10431);
and U10624 (N_10624,N_10440,N_10348);
xor U10625 (N_10625,N_10453,N_10416);
and U10626 (N_10626,N_10364,N_10398);
xnor U10627 (N_10627,N_10329,N_10352);
or U10628 (N_10628,N_10368,N_10358);
nor U10629 (N_10629,N_10436,N_10317);
nand U10630 (N_10630,N_10455,N_10364);
nor U10631 (N_10631,N_10312,N_10349);
and U10632 (N_10632,N_10491,N_10393);
or U10633 (N_10633,N_10362,N_10321);
or U10634 (N_10634,N_10472,N_10415);
nand U10635 (N_10635,N_10450,N_10327);
and U10636 (N_10636,N_10316,N_10298);
xor U10637 (N_10637,N_10429,N_10410);
or U10638 (N_10638,N_10348,N_10379);
and U10639 (N_10639,N_10357,N_10314);
or U10640 (N_10640,N_10266,N_10350);
nor U10641 (N_10641,N_10412,N_10444);
nand U10642 (N_10642,N_10329,N_10368);
or U10643 (N_10643,N_10436,N_10461);
nor U10644 (N_10644,N_10480,N_10305);
or U10645 (N_10645,N_10408,N_10280);
or U10646 (N_10646,N_10271,N_10341);
or U10647 (N_10647,N_10336,N_10400);
nand U10648 (N_10648,N_10399,N_10260);
or U10649 (N_10649,N_10315,N_10480);
nand U10650 (N_10650,N_10307,N_10318);
and U10651 (N_10651,N_10453,N_10419);
nor U10652 (N_10652,N_10373,N_10383);
nor U10653 (N_10653,N_10452,N_10351);
or U10654 (N_10654,N_10402,N_10278);
and U10655 (N_10655,N_10332,N_10340);
and U10656 (N_10656,N_10342,N_10350);
and U10657 (N_10657,N_10461,N_10463);
or U10658 (N_10658,N_10371,N_10364);
xor U10659 (N_10659,N_10355,N_10356);
nor U10660 (N_10660,N_10278,N_10251);
and U10661 (N_10661,N_10358,N_10488);
nor U10662 (N_10662,N_10492,N_10468);
and U10663 (N_10663,N_10326,N_10351);
nand U10664 (N_10664,N_10394,N_10307);
nand U10665 (N_10665,N_10484,N_10416);
or U10666 (N_10666,N_10382,N_10384);
and U10667 (N_10667,N_10393,N_10298);
and U10668 (N_10668,N_10341,N_10469);
or U10669 (N_10669,N_10338,N_10359);
nor U10670 (N_10670,N_10330,N_10479);
or U10671 (N_10671,N_10333,N_10353);
and U10672 (N_10672,N_10271,N_10497);
xnor U10673 (N_10673,N_10292,N_10333);
nand U10674 (N_10674,N_10376,N_10486);
and U10675 (N_10675,N_10396,N_10435);
nand U10676 (N_10676,N_10415,N_10414);
nor U10677 (N_10677,N_10488,N_10390);
nand U10678 (N_10678,N_10269,N_10393);
xnor U10679 (N_10679,N_10325,N_10435);
and U10680 (N_10680,N_10274,N_10329);
nor U10681 (N_10681,N_10256,N_10365);
nor U10682 (N_10682,N_10294,N_10465);
and U10683 (N_10683,N_10268,N_10277);
xor U10684 (N_10684,N_10374,N_10261);
and U10685 (N_10685,N_10432,N_10498);
nand U10686 (N_10686,N_10356,N_10255);
or U10687 (N_10687,N_10417,N_10294);
nand U10688 (N_10688,N_10303,N_10339);
nand U10689 (N_10689,N_10396,N_10258);
nor U10690 (N_10690,N_10329,N_10492);
and U10691 (N_10691,N_10274,N_10474);
or U10692 (N_10692,N_10481,N_10274);
nor U10693 (N_10693,N_10470,N_10478);
or U10694 (N_10694,N_10423,N_10397);
nor U10695 (N_10695,N_10276,N_10358);
and U10696 (N_10696,N_10487,N_10458);
or U10697 (N_10697,N_10284,N_10283);
and U10698 (N_10698,N_10304,N_10284);
nor U10699 (N_10699,N_10397,N_10345);
nand U10700 (N_10700,N_10286,N_10348);
nor U10701 (N_10701,N_10379,N_10409);
nand U10702 (N_10702,N_10459,N_10480);
and U10703 (N_10703,N_10474,N_10498);
nand U10704 (N_10704,N_10442,N_10411);
nand U10705 (N_10705,N_10469,N_10268);
and U10706 (N_10706,N_10487,N_10266);
nor U10707 (N_10707,N_10467,N_10319);
xnor U10708 (N_10708,N_10387,N_10412);
or U10709 (N_10709,N_10340,N_10401);
nor U10710 (N_10710,N_10266,N_10355);
nor U10711 (N_10711,N_10350,N_10484);
xor U10712 (N_10712,N_10286,N_10259);
and U10713 (N_10713,N_10251,N_10455);
and U10714 (N_10714,N_10406,N_10424);
xnor U10715 (N_10715,N_10489,N_10325);
xor U10716 (N_10716,N_10390,N_10366);
nand U10717 (N_10717,N_10432,N_10317);
nor U10718 (N_10718,N_10270,N_10453);
nand U10719 (N_10719,N_10324,N_10339);
and U10720 (N_10720,N_10327,N_10365);
or U10721 (N_10721,N_10487,N_10449);
nand U10722 (N_10722,N_10410,N_10265);
nand U10723 (N_10723,N_10487,N_10327);
or U10724 (N_10724,N_10446,N_10443);
nand U10725 (N_10725,N_10411,N_10301);
nand U10726 (N_10726,N_10421,N_10354);
nand U10727 (N_10727,N_10339,N_10265);
or U10728 (N_10728,N_10480,N_10441);
nand U10729 (N_10729,N_10250,N_10313);
nand U10730 (N_10730,N_10297,N_10472);
nor U10731 (N_10731,N_10416,N_10439);
nand U10732 (N_10732,N_10331,N_10406);
and U10733 (N_10733,N_10411,N_10419);
nor U10734 (N_10734,N_10324,N_10251);
nor U10735 (N_10735,N_10363,N_10488);
nor U10736 (N_10736,N_10261,N_10250);
xor U10737 (N_10737,N_10479,N_10494);
or U10738 (N_10738,N_10283,N_10378);
and U10739 (N_10739,N_10380,N_10371);
nand U10740 (N_10740,N_10386,N_10468);
or U10741 (N_10741,N_10357,N_10448);
xnor U10742 (N_10742,N_10311,N_10337);
nor U10743 (N_10743,N_10325,N_10403);
nor U10744 (N_10744,N_10447,N_10445);
nor U10745 (N_10745,N_10407,N_10483);
and U10746 (N_10746,N_10259,N_10355);
or U10747 (N_10747,N_10305,N_10308);
or U10748 (N_10748,N_10485,N_10353);
nand U10749 (N_10749,N_10349,N_10432);
nand U10750 (N_10750,N_10631,N_10623);
and U10751 (N_10751,N_10597,N_10652);
nand U10752 (N_10752,N_10533,N_10518);
and U10753 (N_10753,N_10744,N_10612);
nor U10754 (N_10754,N_10693,N_10526);
nand U10755 (N_10755,N_10588,N_10701);
or U10756 (N_10756,N_10564,N_10544);
nor U10757 (N_10757,N_10735,N_10747);
and U10758 (N_10758,N_10619,N_10705);
xnor U10759 (N_10759,N_10594,N_10503);
and U10760 (N_10760,N_10695,N_10749);
or U10761 (N_10761,N_10653,N_10713);
nand U10762 (N_10762,N_10629,N_10536);
and U10763 (N_10763,N_10674,N_10610);
nor U10764 (N_10764,N_10586,N_10531);
nor U10765 (N_10765,N_10616,N_10537);
xnor U10766 (N_10766,N_10504,N_10680);
and U10767 (N_10767,N_10549,N_10545);
xnor U10768 (N_10768,N_10525,N_10511);
nand U10769 (N_10769,N_10615,N_10719);
nand U10770 (N_10770,N_10581,N_10738);
or U10771 (N_10771,N_10611,N_10578);
nand U10772 (N_10772,N_10734,N_10563);
or U10773 (N_10773,N_10638,N_10643);
nand U10774 (N_10774,N_10649,N_10617);
and U10775 (N_10775,N_10607,N_10668);
and U10776 (N_10776,N_10727,N_10574);
xnor U10777 (N_10777,N_10609,N_10552);
or U10778 (N_10778,N_10625,N_10630);
nor U10779 (N_10779,N_10627,N_10534);
nor U10780 (N_10780,N_10570,N_10634);
and U10781 (N_10781,N_10515,N_10556);
and U10782 (N_10782,N_10672,N_10624);
nand U10783 (N_10783,N_10647,N_10679);
xnor U10784 (N_10784,N_10745,N_10746);
nor U10785 (N_10785,N_10725,N_10673);
and U10786 (N_10786,N_10710,N_10656);
nand U10787 (N_10787,N_10568,N_10614);
xor U10788 (N_10788,N_10626,N_10722);
and U10789 (N_10789,N_10553,N_10520);
or U10790 (N_10790,N_10642,N_10732);
or U10791 (N_10791,N_10692,N_10689);
nor U10792 (N_10792,N_10517,N_10714);
nand U10793 (N_10793,N_10528,N_10508);
xnor U10794 (N_10794,N_10726,N_10733);
nor U10795 (N_10795,N_10731,N_10605);
or U10796 (N_10796,N_10539,N_10524);
or U10797 (N_10797,N_10654,N_10620);
or U10798 (N_10798,N_10567,N_10579);
or U10799 (N_10799,N_10507,N_10576);
nor U10800 (N_10800,N_10669,N_10741);
and U10801 (N_10801,N_10593,N_10580);
or U10802 (N_10802,N_10635,N_10596);
and U10803 (N_10803,N_10748,N_10502);
nand U10804 (N_10804,N_10698,N_10509);
and U10805 (N_10805,N_10657,N_10548);
xor U10806 (N_10806,N_10583,N_10742);
and U10807 (N_10807,N_10685,N_10743);
nand U10808 (N_10808,N_10589,N_10648);
nor U10809 (N_10809,N_10683,N_10547);
xnor U10810 (N_10810,N_10501,N_10688);
or U10811 (N_10811,N_10723,N_10599);
or U10812 (N_10812,N_10637,N_10681);
nor U10813 (N_10813,N_10682,N_10711);
and U10814 (N_10814,N_10551,N_10558);
xnor U10815 (N_10815,N_10651,N_10591);
nor U10816 (N_10816,N_10529,N_10684);
xnor U10817 (N_10817,N_10587,N_10646);
and U10818 (N_10818,N_10641,N_10645);
nand U10819 (N_10819,N_10505,N_10696);
nor U10820 (N_10820,N_10557,N_10598);
and U10821 (N_10821,N_10707,N_10659);
and U10822 (N_10822,N_10699,N_10708);
nand U10823 (N_10823,N_10585,N_10535);
xor U10824 (N_10824,N_10527,N_10655);
and U10825 (N_10825,N_10514,N_10667);
and U10826 (N_10826,N_10640,N_10665);
and U10827 (N_10827,N_10715,N_10516);
nor U10828 (N_10828,N_10584,N_10561);
and U10829 (N_10829,N_10560,N_10729);
and U10830 (N_10830,N_10555,N_10632);
nand U10831 (N_10831,N_10554,N_10658);
nor U10832 (N_10832,N_10500,N_10540);
nor U10833 (N_10833,N_10690,N_10644);
and U10834 (N_10834,N_10532,N_10530);
nand U10835 (N_10835,N_10716,N_10739);
nor U10836 (N_10836,N_10592,N_10523);
and U10837 (N_10837,N_10694,N_10670);
and U10838 (N_10838,N_10572,N_10543);
or U10839 (N_10839,N_10541,N_10704);
nor U10840 (N_10840,N_10510,N_10671);
and U10841 (N_10841,N_10677,N_10724);
and U10842 (N_10842,N_10709,N_10675);
or U10843 (N_10843,N_10636,N_10602);
nand U10844 (N_10844,N_10661,N_10512);
nor U10845 (N_10845,N_10702,N_10676);
nor U10846 (N_10846,N_10550,N_10622);
nor U10847 (N_10847,N_10571,N_10559);
and U10848 (N_10848,N_10663,N_10562);
nand U10849 (N_10849,N_10595,N_10662);
nor U10850 (N_10850,N_10542,N_10600);
or U10851 (N_10851,N_10728,N_10687);
or U10852 (N_10852,N_10603,N_10628);
nor U10853 (N_10853,N_10703,N_10721);
or U10854 (N_10854,N_10633,N_10650);
nand U10855 (N_10855,N_10706,N_10606);
or U10856 (N_10856,N_10538,N_10519);
nand U10857 (N_10857,N_10660,N_10577);
nand U10858 (N_10858,N_10608,N_10740);
nand U10859 (N_10859,N_10522,N_10613);
nor U10860 (N_10860,N_10666,N_10546);
nor U10861 (N_10861,N_10506,N_10664);
nand U10862 (N_10862,N_10697,N_10686);
and U10863 (N_10863,N_10573,N_10639);
or U10864 (N_10864,N_10569,N_10737);
or U10865 (N_10865,N_10730,N_10618);
nor U10866 (N_10866,N_10601,N_10565);
and U10867 (N_10867,N_10736,N_10521);
or U10868 (N_10868,N_10575,N_10717);
nor U10869 (N_10869,N_10566,N_10700);
or U10870 (N_10870,N_10718,N_10621);
and U10871 (N_10871,N_10691,N_10720);
or U10872 (N_10872,N_10712,N_10513);
xor U10873 (N_10873,N_10604,N_10590);
or U10874 (N_10874,N_10582,N_10678);
nand U10875 (N_10875,N_10680,N_10699);
and U10876 (N_10876,N_10593,N_10646);
nand U10877 (N_10877,N_10571,N_10639);
nand U10878 (N_10878,N_10704,N_10691);
nor U10879 (N_10879,N_10554,N_10500);
nor U10880 (N_10880,N_10541,N_10633);
nor U10881 (N_10881,N_10668,N_10565);
and U10882 (N_10882,N_10691,N_10632);
xnor U10883 (N_10883,N_10551,N_10668);
or U10884 (N_10884,N_10677,N_10685);
nand U10885 (N_10885,N_10682,N_10654);
xor U10886 (N_10886,N_10517,N_10721);
and U10887 (N_10887,N_10680,N_10746);
nand U10888 (N_10888,N_10569,N_10525);
nor U10889 (N_10889,N_10544,N_10500);
nand U10890 (N_10890,N_10707,N_10650);
and U10891 (N_10891,N_10682,N_10741);
or U10892 (N_10892,N_10550,N_10712);
nor U10893 (N_10893,N_10532,N_10732);
or U10894 (N_10894,N_10744,N_10554);
nand U10895 (N_10895,N_10535,N_10576);
nand U10896 (N_10896,N_10646,N_10631);
xnor U10897 (N_10897,N_10707,N_10645);
or U10898 (N_10898,N_10743,N_10649);
nor U10899 (N_10899,N_10620,N_10511);
nand U10900 (N_10900,N_10636,N_10623);
or U10901 (N_10901,N_10523,N_10747);
and U10902 (N_10902,N_10533,N_10613);
nor U10903 (N_10903,N_10686,N_10689);
or U10904 (N_10904,N_10531,N_10553);
nand U10905 (N_10905,N_10631,N_10649);
and U10906 (N_10906,N_10590,N_10650);
or U10907 (N_10907,N_10667,N_10636);
xor U10908 (N_10908,N_10566,N_10533);
and U10909 (N_10909,N_10567,N_10500);
and U10910 (N_10910,N_10715,N_10735);
and U10911 (N_10911,N_10743,N_10519);
nand U10912 (N_10912,N_10536,N_10652);
xnor U10913 (N_10913,N_10700,N_10542);
and U10914 (N_10914,N_10700,N_10699);
nor U10915 (N_10915,N_10636,N_10638);
or U10916 (N_10916,N_10595,N_10661);
nand U10917 (N_10917,N_10635,N_10546);
xor U10918 (N_10918,N_10590,N_10527);
or U10919 (N_10919,N_10601,N_10703);
nor U10920 (N_10920,N_10656,N_10532);
and U10921 (N_10921,N_10542,N_10723);
nand U10922 (N_10922,N_10577,N_10710);
xor U10923 (N_10923,N_10574,N_10648);
and U10924 (N_10924,N_10526,N_10709);
nand U10925 (N_10925,N_10632,N_10726);
xor U10926 (N_10926,N_10643,N_10621);
or U10927 (N_10927,N_10670,N_10695);
and U10928 (N_10928,N_10529,N_10725);
nand U10929 (N_10929,N_10510,N_10578);
nor U10930 (N_10930,N_10582,N_10570);
or U10931 (N_10931,N_10604,N_10507);
or U10932 (N_10932,N_10522,N_10733);
and U10933 (N_10933,N_10542,N_10577);
and U10934 (N_10934,N_10661,N_10548);
nand U10935 (N_10935,N_10603,N_10617);
or U10936 (N_10936,N_10668,N_10577);
and U10937 (N_10937,N_10607,N_10562);
or U10938 (N_10938,N_10697,N_10665);
and U10939 (N_10939,N_10614,N_10630);
nor U10940 (N_10940,N_10513,N_10634);
and U10941 (N_10941,N_10504,N_10581);
nand U10942 (N_10942,N_10630,N_10667);
nand U10943 (N_10943,N_10624,N_10633);
or U10944 (N_10944,N_10705,N_10678);
nand U10945 (N_10945,N_10649,N_10572);
nor U10946 (N_10946,N_10748,N_10653);
and U10947 (N_10947,N_10698,N_10714);
and U10948 (N_10948,N_10724,N_10657);
nor U10949 (N_10949,N_10729,N_10595);
nor U10950 (N_10950,N_10592,N_10674);
xnor U10951 (N_10951,N_10696,N_10592);
nor U10952 (N_10952,N_10728,N_10507);
and U10953 (N_10953,N_10521,N_10705);
xnor U10954 (N_10954,N_10607,N_10708);
nand U10955 (N_10955,N_10748,N_10664);
or U10956 (N_10956,N_10681,N_10697);
nand U10957 (N_10957,N_10612,N_10556);
nand U10958 (N_10958,N_10552,N_10630);
nand U10959 (N_10959,N_10681,N_10698);
nor U10960 (N_10960,N_10743,N_10525);
or U10961 (N_10961,N_10583,N_10656);
nand U10962 (N_10962,N_10544,N_10723);
nor U10963 (N_10963,N_10554,N_10629);
or U10964 (N_10964,N_10745,N_10741);
or U10965 (N_10965,N_10646,N_10642);
or U10966 (N_10966,N_10603,N_10631);
xor U10967 (N_10967,N_10639,N_10645);
nand U10968 (N_10968,N_10719,N_10616);
or U10969 (N_10969,N_10616,N_10538);
nand U10970 (N_10970,N_10542,N_10733);
or U10971 (N_10971,N_10537,N_10701);
nor U10972 (N_10972,N_10542,N_10684);
xor U10973 (N_10973,N_10625,N_10617);
and U10974 (N_10974,N_10698,N_10712);
nand U10975 (N_10975,N_10696,N_10737);
and U10976 (N_10976,N_10521,N_10645);
and U10977 (N_10977,N_10632,N_10638);
nor U10978 (N_10978,N_10524,N_10518);
nor U10979 (N_10979,N_10628,N_10693);
and U10980 (N_10980,N_10567,N_10517);
or U10981 (N_10981,N_10675,N_10519);
xor U10982 (N_10982,N_10575,N_10556);
nor U10983 (N_10983,N_10596,N_10523);
nand U10984 (N_10984,N_10630,N_10555);
or U10985 (N_10985,N_10708,N_10502);
nand U10986 (N_10986,N_10500,N_10739);
nor U10987 (N_10987,N_10546,N_10655);
nor U10988 (N_10988,N_10713,N_10724);
xor U10989 (N_10989,N_10637,N_10518);
nand U10990 (N_10990,N_10549,N_10612);
or U10991 (N_10991,N_10596,N_10545);
xor U10992 (N_10992,N_10622,N_10649);
and U10993 (N_10993,N_10594,N_10637);
and U10994 (N_10994,N_10652,N_10544);
nand U10995 (N_10995,N_10671,N_10717);
nor U10996 (N_10996,N_10590,N_10511);
nand U10997 (N_10997,N_10597,N_10534);
nor U10998 (N_10998,N_10612,N_10738);
or U10999 (N_10999,N_10671,N_10728);
or U11000 (N_11000,N_10828,N_10992);
or U11001 (N_11001,N_10939,N_10956);
or U11002 (N_11002,N_10865,N_10875);
nor U11003 (N_11003,N_10868,N_10837);
nand U11004 (N_11004,N_10976,N_10794);
and U11005 (N_11005,N_10769,N_10781);
or U11006 (N_11006,N_10945,N_10783);
nor U11007 (N_11007,N_10898,N_10764);
and U11008 (N_11008,N_10827,N_10880);
or U11009 (N_11009,N_10754,N_10774);
nand U11010 (N_11010,N_10763,N_10829);
nand U11011 (N_11011,N_10947,N_10985);
and U11012 (N_11012,N_10864,N_10831);
and U11013 (N_11013,N_10784,N_10944);
nor U11014 (N_11014,N_10779,N_10917);
nor U11015 (N_11015,N_10772,N_10767);
or U11016 (N_11016,N_10757,N_10780);
and U11017 (N_11017,N_10942,N_10995);
or U11018 (N_11018,N_10792,N_10893);
nand U11019 (N_11019,N_10926,N_10921);
and U11020 (N_11020,N_10765,N_10884);
nand U11021 (N_11021,N_10869,N_10771);
nand U11022 (N_11022,N_10814,N_10907);
nand U11023 (N_11023,N_10925,N_10896);
or U11024 (N_11024,N_10873,N_10770);
and U11025 (N_11025,N_10988,N_10844);
and U11026 (N_11026,N_10891,N_10870);
nand U11027 (N_11027,N_10963,N_10800);
and U11028 (N_11028,N_10782,N_10803);
and U11029 (N_11029,N_10902,N_10820);
nand U11030 (N_11030,N_10804,N_10920);
and U11031 (N_11031,N_10801,N_10997);
or U11032 (N_11032,N_10959,N_10841);
nor U11033 (N_11033,N_10846,N_10847);
xnor U11034 (N_11034,N_10906,N_10924);
and U11035 (N_11035,N_10885,N_10979);
xnor U11036 (N_11036,N_10991,N_10759);
and U11037 (N_11037,N_10993,N_10855);
nand U11038 (N_11038,N_10861,N_10911);
and U11039 (N_11039,N_10857,N_10816);
nor U11040 (N_11040,N_10900,N_10927);
or U11041 (N_11041,N_10922,N_10912);
or U11042 (N_11042,N_10789,N_10830);
or U11043 (N_11043,N_10833,N_10928);
nor U11044 (N_11044,N_10984,N_10807);
nand U11045 (N_11045,N_10951,N_10903);
nor U11046 (N_11046,N_10834,N_10923);
nor U11047 (N_11047,N_10866,N_10753);
nor U11048 (N_11048,N_10845,N_10937);
nand U11049 (N_11049,N_10949,N_10823);
or U11050 (N_11050,N_10950,N_10969);
nor U11051 (N_11051,N_10788,N_10970);
nand U11052 (N_11052,N_10849,N_10972);
nand U11053 (N_11053,N_10766,N_10825);
or U11054 (N_11054,N_10961,N_10776);
nand U11055 (N_11055,N_10967,N_10863);
nand U11056 (N_11056,N_10876,N_10821);
nor U11057 (N_11057,N_10762,N_10892);
nor U11058 (N_11058,N_10839,N_10777);
or U11059 (N_11059,N_10796,N_10813);
and U11060 (N_11060,N_10994,N_10952);
and U11061 (N_11061,N_10879,N_10914);
and U11062 (N_11062,N_10895,N_10890);
nand U11063 (N_11063,N_10888,N_10860);
nand U11064 (N_11064,N_10878,N_10987);
or U11065 (N_11065,N_10808,N_10854);
nor U11066 (N_11066,N_10760,N_10981);
nor U11067 (N_11067,N_10802,N_10842);
nand U11068 (N_11068,N_10948,N_10982);
nand U11069 (N_11069,N_10983,N_10916);
or U11070 (N_11070,N_10971,N_10793);
nand U11071 (N_11071,N_10897,N_10953);
or U11072 (N_11072,N_10806,N_10930);
xnor U11073 (N_11073,N_10843,N_10932);
or U11074 (N_11074,N_10812,N_10955);
and U11075 (N_11075,N_10908,N_10797);
and U11076 (N_11076,N_10785,N_10968);
and U11077 (N_11077,N_10755,N_10974);
nor U11078 (N_11078,N_10929,N_10989);
or U11079 (N_11079,N_10874,N_10934);
nor U11080 (N_11080,N_10858,N_10931);
and U11081 (N_11081,N_10894,N_10965);
and U11082 (N_11082,N_10915,N_10935);
nand U11083 (N_11083,N_10957,N_10877);
and U11084 (N_11084,N_10835,N_10752);
xnor U11085 (N_11085,N_10838,N_10954);
or U11086 (N_11086,N_10901,N_10856);
nand U11087 (N_11087,N_10973,N_10990);
or U11088 (N_11088,N_10756,N_10905);
nor U11089 (N_11089,N_10853,N_10986);
nand U11090 (N_11090,N_10938,N_10882);
nor U11091 (N_11091,N_10946,N_10980);
xor U11092 (N_11092,N_10775,N_10811);
and U11093 (N_11093,N_10960,N_10818);
nand U11094 (N_11094,N_10848,N_10904);
and U11095 (N_11095,N_10791,N_10805);
nor U11096 (N_11096,N_10778,N_10881);
nand U11097 (N_11097,N_10850,N_10886);
nand U11098 (N_11098,N_10998,N_10872);
xor U11099 (N_11099,N_10799,N_10819);
xnor U11100 (N_11100,N_10798,N_10822);
nand U11101 (N_11101,N_10977,N_10910);
or U11102 (N_11102,N_10826,N_10978);
nand U11103 (N_11103,N_10809,N_10936);
or U11104 (N_11104,N_10975,N_10751);
xnor U11105 (N_11105,N_10824,N_10871);
or U11106 (N_11106,N_10909,N_10773);
nand U11107 (N_11107,N_10867,N_10795);
nor U11108 (N_11108,N_10790,N_10964);
nor U11109 (N_11109,N_10758,N_10918);
nor U11110 (N_11110,N_10962,N_10919);
nor U11111 (N_11111,N_10996,N_10832);
or U11112 (N_11112,N_10761,N_10958);
xor U11113 (N_11113,N_10851,N_10862);
or U11114 (N_11114,N_10859,N_10966);
or U11115 (N_11115,N_10887,N_10750);
or U11116 (N_11116,N_10883,N_10941);
nand U11117 (N_11117,N_10943,N_10933);
nor U11118 (N_11118,N_10940,N_10999);
xnor U11119 (N_11119,N_10840,N_10786);
nand U11120 (N_11120,N_10768,N_10817);
or U11121 (N_11121,N_10810,N_10889);
nor U11122 (N_11122,N_10836,N_10852);
or U11123 (N_11123,N_10815,N_10913);
or U11124 (N_11124,N_10899,N_10787);
xnor U11125 (N_11125,N_10837,N_10970);
xor U11126 (N_11126,N_10874,N_10760);
nor U11127 (N_11127,N_10935,N_10778);
or U11128 (N_11128,N_10865,N_10857);
and U11129 (N_11129,N_10865,N_10951);
and U11130 (N_11130,N_10956,N_10802);
and U11131 (N_11131,N_10840,N_10900);
nand U11132 (N_11132,N_10896,N_10776);
nor U11133 (N_11133,N_10985,N_10888);
and U11134 (N_11134,N_10767,N_10936);
and U11135 (N_11135,N_10839,N_10897);
nor U11136 (N_11136,N_10811,N_10961);
or U11137 (N_11137,N_10910,N_10898);
and U11138 (N_11138,N_10903,N_10964);
xor U11139 (N_11139,N_10781,N_10844);
or U11140 (N_11140,N_10993,N_10872);
or U11141 (N_11141,N_10962,N_10847);
nor U11142 (N_11142,N_10784,N_10984);
nor U11143 (N_11143,N_10974,N_10795);
or U11144 (N_11144,N_10952,N_10845);
nand U11145 (N_11145,N_10977,N_10901);
xnor U11146 (N_11146,N_10941,N_10755);
or U11147 (N_11147,N_10931,N_10889);
nand U11148 (N_11148,N_10843,N_10997);
xnor U11149 (N_11149,N_10799,N_10846);
nor U11150 (N_11150,N_10949,N_10757);
nor U11151 (N_11151,N_10984,N_10937);
and U11152 (N_11152,N_10873,N_10910);
or U11153 (N_11153,N_10757,N_10880);
nand U11154 (N_11154,N_10906,N_10817);
or U11155 (N_11155,N_10907,N_10797);
or U11156 (N_11156,N_10893,N_10935);
nand U11157 (N_11157,N_10803,N_10814);
or U11158 (N_11158,N_10771,N_10999);
and U11159 (N_11159,N_10798,N_10821);
or U11160 (N_11160,N_10990,N_10908);
and U11161 (N_11161,N_10871,N_10819);
or U11162 (N_11162,N_10797,N_10921);
or U11163 (N_11163,N_10981,N_10956);
nor U11164 (N_11164,N_10812,N_10863);
and U11165 (N_11165,N_10786,N_10948);
nor U11166 (N_11166,N_10947,N_10806);
nor U11167 (N_11167,N_10827,N_10987);
nor U11168 (N_11168,N_10780,N_10952);
or U11169 (N_11169,N_10855,N_10940);
or U11170 (N_11170,N_10791,N_10968);
or U11171 (N_11171,N_10881,N_10952);
nand U11172 (N_11172,N_10762,N_10920);
nor U11173 (N_11173,N_10966,N_10983);
nor U11174 (N_11174,N_10847,N_10991);
and U11175 (N_11175,N_10952,N_10904);
and U11176 (N_11176,N_10939,N_10989);
and U11177 (N_11177,N_10874,N_10850);
nor U11178 (N_11178,N_10894,N_10884);
and U11179 (N_11179,N_10988,N_10955);
nand U11180 (N_11180,N_10756,N_10785);
or U11181 (N_11181,N_10861,N_10929);
nand U11182 (N_11182,N_10960,N_10837);
and U11183 (N_11183,N_10839,N_10962);
or U11184 (N_11184,N_10758,N_10987);
or U11185 (N_11185,N_10763,N_10864);
or U11186 (N_11186,N_10761,N_10827);
and U11187 (N_11187,N_10925,N_10865);
nand U11188 (N_11188,N_10789,N_10875);
nor U11189 (N_11189,N_10819,N_10779);
and U11190 (N_11190,N_10940,N_10965);
xor U11191 (N_11191,N_10919,N_10823);
nand U11192 (N_11192,N_10951,N_10962);
nor U11193 (N_11193,N_10941,N_10928);
nand U11194 (N_11194,N_10996,N_10856);
nand U11195 (N_11195,N_10851,N_10813);
nand U11196 (N_11196,N_10962,N_10821);
nor U11197 (N_11197,N_10797,N_10997);
nor U11198 (N_11198,N_10997,N_10981);
nand U11199 (N_11199,N_10978,N_10982);
nor U11200 (N_11200,N_10784,N_10809);
xor U11201 (N_11201,N_10909,N_10870);
nor U11202 (N_11202,N_10993,N_10976);
nand U11203 (N_11203,N_10839,N_10862);
nand U11204 (N_11204,N_10889,N_10941);
or U11205 (N_11205,N_10831,N_10962);
and U11206 (N_11206,N_10848,N_10870);
nor U11207 (N_11207,N_10876,N_10826);
or U11208 (N_11208,N_10910,N_10823);
xnor U11209 (N_11209,N_10835,N_10965);
or U11210 (N_11210,N_10884,N_10825);
xor U11211 (N_11211,N_10917,N_10822);
nor U11212 (N_11212,N_10826,N_10867);
and U11213 (N_11213,N_10868,N_10890);
nor U11214 (N_11214,N_10855,N_10992);
or U11215 (N_11215,N_10832,N_10856);
or U11216 (N_11216,N_10915,N_10949);
and U11217 (N_11217,N_10969,N_10764);
and U11218 (N_11218,N_10810,N_10962);
and U11219 (N_11219,N_10804,N_10793);
nor U11220 (N_11220,N_10982,N_10892);
nor U11221 (N_11221,N_10788,N_10965);
and U11222 (N_11222,N_10947,N_10925);
nand U11223 (N_11223,N_10897,N_10962);
and U11224 (N_11224,N_10836,N_10859);
nor U11225 (N_11225,N_10999,N_10898);
nor U11226 (N_11226,N_10758,N_10959);
xnor U11227 (N_11227,N_10837,N_10798);
and U11228 (N_11228,N_10775,N_10940);
and U11229 (N_11229,N_10755,N_10868);
and U11230 (N_11230,N_10793,N_10816);
and U11231 (N_11231,N_10838,N_10788);
xnor U11232 (N_11232,N_10821,N_10830);
xor U11233 (N_11233,N_10762,N_10836);
nand U11234 (N_11234,N_10930,N_10918);
and U11235 (N_11235,N_10840,N_10960);
or U11236 (N_11236,N_10795,N_10973);
or U11237 (N_11237,N_10870,N_10928);
and U11238 (N_11238,N_10759,N_10874);
nor U11239 (N_11239,N_10843,N_10765);
nand U11240 (N_11240,N_10997,N_10796);
or U11241 (N_11241,N_10867,N_10835);
or U11242 (N_11242,N_10837,N_10909);
and U11243 (N_11243,N_10842,N_10824);
or U11244 (N_11244,N_10773,N_10877);
or U11245 (N_11245,N_10908,N_10867);
nor U11246 (N_11246,N_10962,N_10862);
nor U11247 (N_11247,N_10869,N_10933);
nor U11248 (N_11248,N_10957,N_10818);
nand U11249 (N_11249,N_10980,N_10987);
or U11250 (N_11250,N_11148,N_11077);
or U11251 (N_11251,N_11163,N_11110);
nand U11252 (N_11252,N_11119,N_11239);
and U11253 (N_11253,N_11207,N_11219);
nand U11254 (N_11254,N_11211,N_11111);
nand U11255 (N_11255,N_11043,N_11192);
and U11256 (N_11256,N_11059,N_11131);
and U11257 (N_11257,N_11039,N_11244);
nand U11258 (N_11258,N_11246,N_11008);
nor U11259 (N_11259,N_11231,N_11033);
or U11260 (N_11260,N_11159,N_11104);
nor U11261 (N_11261,N_11158,N_11050);
or U11262 (N_11262,N_11000,N_11180);
nand U11263 (N_11263,N_11206,N_11031);
nor U11264 (N_11264,N_11140,N_11145);
nor U11265 (N_11265,N_11221,N_11238);
and U11266 (N_11266,N_11025,N_11137);
or U11267 (N_11267,N_11210,N_11090);
nand U11268 (N_11268,N_11243,N_11197);
nand U11269 (N_11269,N_11103,N_11228);
xnor U11270 (N_11270,N_11213,N_11096);
nor U11271 (N_11271,N_11037,N_11012);
nor U11272 (N_11272,N_11247,N_11181);
nand U11273 (N_11273,N_11041,N_11193);
or U11274 (N_11274,N_11006,N_11068);
and U11275 (N_11275,N_11237,N_11182);
or U11276 (N_11276,N_11203,N_11030);
and U11277 (N_11277,N_11162,N_11015);
nand U11278 (N_11278,N_11184,N_11049);
xor U11279 (N_11279,N_11028,N_11116);
nand U11280 (N_11280,N_11010,N_11044);
xnor U11281 (N_11281,N_11241,N_11229);
nor U11282 (N_11282,N_11100,N_11153);
nor U11283 (N_11283,N_11017,N_11214);
and U11284 (N_11284,N_11105,N_11166);
or U11285 (N_11285,N_11106,N_11040);
and U11286 (N_11286,N_11136,N_11132);
nor U11287 (N_11287,N_11060,N_11141);
and U11288 (N_11288,N_11144,N_11075);
or U11289 (N_11289,N_11073,N_11069);
and U11290 (N_11290,N_11123,N_11078);
xnor U11291 (N_11291,N_11081,N_11005);
xor U11292 (N_11292,N_11091,N_11056);
and U11293 (N_11293,N_11095,N_11085);
nand U11294 (N_11294,N_11023,N_11194);
or U11295 (N_11295,N_11013,N_11127);
xnor U11296 (N_11296,N_11149,N_11045);
and U11297 (N_11297,N_11101,N_11208);
xnor U11298 (N_11298,N_11011,N_11058);
xnor U11299 (N_11299,N_11089,N_11191);
or U11300 (N_11300,N_11070,N_11034);
xor U11301 (N_11301,N_11165,N_11217);
nor U11302 (N_11302,N_11157,N_11086);
and U11303 (N_11303,N_11097,N_11155);
or U11304 (N_11304,N_11022,N_11220);
xor U11305 (N_11305,N_11186,N_11222);
or U11306 (N_11306,N_11019,N_11024);
nand U11307 (N_11307,N_11128,N_11076);
nor U11308 (N_11308,N_11133,N_11212);
xor U11309 (N_11309,N_11183,N_11062);
xor U11310 (N_11310,N_11021,N_11218);
and U11311 (N_11311,N_11199,N_11195);
or U11312 (N_11312,N_11249,N_11064);
or U11313 (N_11313,N_11160,N_11026);
nand U11314 (N_11314,N_11109,N_11168);
or U11315 (N_11315,N_11083,N_11138);
and U11316 (N_11316,N_11080,N_11233);
xor U11317 (N_11317,N_11240,N_11118);
or U11318 (N_11318,N_11014,N_11134);
nor U11319 (N_11319,N_11224,N_11171);
or U11320 (N_11320,N_11248,N_11169);
and U11321 (N_11321,N_11004,N_11230);
nor U11322 (N_11322,N_11072,N_11172);
and U11323 (N_11323,N_11121,N_11209);
and U11324 (N_11324,N_11066,N_11079);
nor U11325 (N_11325,N_11142,N_11055);
or U11326 (N_11326,N_11205,N_11174);
nand U11327 (N_11327,N_11236,N_11147);
nand U11328 (N_11328,N_11053,N_11232);
or U11329 (N_11329,N_11063,N_11176);
and U11330 (N_11330,N_11035,N_11223);
nand U11331 (N_11331,N_11225,N_11146);
nand U11332 (N_11332,N_11179,N_11001);
and U11333 (N_11333,N_11067,N_11087);
nor U11334 (N_11334,N_11234,N_11122);
and U11335 (N_11335,N_11143,N_11036);
and U11336 (N_11336,N_11130,N_11177);
and U11337 (N_11337,N_11188,N_11125);
nand U11338 (N_11338,N_11245,N_11108);
or U11339 (N_11339,N_11139,N_11027);
and U11340 (N_11340,N_11071,N_11092);
xnor U11341 (N_11341,N_11057,N_11046);
or U11342 (N_11342,N_11152,N_11115);
nand U11343 (N_11343,N_11175,N_11200);
nand U11344 (N_11344,N_11084,N_11242);
or U11345 (N_11345,N_11150,N_11112);
or U11346 (N_11346,N_11007,N_11201);
and U11347 (N_11347,N_11102,N_11178);
nand U11348 (N_11348,N_11202,N_11167);
xor U11349 (N_11349,N_11173,N_11018);
nand U11350 (N_11350,N_11204,N_11120);
and U11351 (N_11351,N_11051,N_11061);
xor U11352 (N_11352,N_11048,N_11235);
and U11353 (N_11353,N_11099,N_11114);
and U11354 (N_11354,N_11129,N_11029);
and U11355 (N_11355,N_11185,N_11126);
nand U11356 (N_11356,N_11164,N_11082);
nand U11357 (N_11357,N_11107,N_11198);
or U11358 (N_11358,N_11093,N_11226);
nand U11359 (N_11359,N_11154,N_11054);
nand U11360 (N_11360,N_11020,N_11156);
or U11361 (N_11361,N_11124,N_11113);
and U11362 (N_11362,N_11151,N_11032);
xor U11363 (N_11363,N_11215,N_11187);
and U11364 (N_11364,N_11117,N_11047);
nand U11365 (N_11365,N_11135,N_11052);
or U11366 (N_11366,N_11161,N_11002);
nand U11367 (N_11367,N_11190,N_11003);
or U11368 (N_11368,N_11038,N_11088);
and U11369 (N_11369,N_11196,N_11098);
or U11370 (N_11370,N_11042,N_11009);
and U11371 (N_11371,N_11094,N_11227);
and U11372 (N_11372,N_11189,N_11216);
and U11373 (N_11373,N_11016,N_11065);
and U11374 (N_11374,N_11074,N_11170);
nor U11375 (N_11375,N_11195,N_11003);
nand U11376 (N_11376,N_11053,N_11012);
and U11377 (N_11377,N_11012,N_11103);
nand U11378 (N_11378,N_11199,N_11111);
nand U11379 (N_11379,N_11196,N_11127);
nand U11380 (N_11380,N_11114,N_11246);
nand U11381 (N_11381,N_11072,N_11057);
nand U11382 (N_11382,N_11190,N_11211);
or U11383 (N_11383,N_11176,N_11014);
xnor U11384 (N_11384,N_11176,N_11123);
or U11385 (N_11385,N_11186,N_11065);
nor U11386 (N_11386,N_11101,N_11152);
or U11387 (N_11387,N_11219,N_11092);
nand U11388 (N_11388,N_11088,N_11015);
and U11389 (N_11389,N_11027,N_11229);
xnor U11390 (N_11390,N_11142,N_11173);
xor U11391 (N_11391,N_11235,N_11219);
or U11392 (N_11392,N_11082,N_11115);
and U11393 (N_11393,N_11075,N_11119);
and U11394 (N_11394,N_11219,N_11099);
nor U11395 (N_11395,N_11001,N_11232);
and U11396 (N_11396,N_11125,N_11243);
and U11397 (N_11397,N_11233,N_11134);
or U11398 (N_11398,N_11167,N_11102);
nor U11399 (N_11399,N_11160,N_11102);
nand U11400 (N_11400,N_11133,N_11150);
or U11401 (N_11401,N_11099,N_11180);
nand U11402 (N_11402,N_11021,N_11171);
or U11403 (N_11403,N_11085,N_11098);
nand U11404 (N_11404,N_11246,N_11018);
or U11405 (N_11405,N_11163,N_11196);
or U11406 (N_11406,N_11100,N_11216);
nand U11407 (N_11407,N_11147,N_11143);
or U11408 (N_11408,N_11126,N_11059);
nand U11409 (N_11409,N_11078,N_11214);
nand U11410 (N_11410,N_11065,N_11008);
nand U11411 (N_11411,N_11098,N_11151);
and U11412 (N_11412,N_11110,N_11018);
nand U11413 (N_11413,N_11057,N_11227);
nor U11414 (N_11414,N_11189,N_11109);
and U11415 (N_11415,N_11111,N_11148);
nand U11416 (N_11416,N_11147,N_11241);
or U11417 (N_11417,N_11000,N_11001);
xnor U11418 (N_11418,N_11193,N_11039);
nor U11419 (N_11419,N_11087,N_11103);
nor U11420 (N_11420,N_11197,N_11226);
xor U11421 (N_11421,N_11145,N_11005);
or U11422 (N_11422,N_11065,N_11086);
xor U11423 (N_11423,N_11072,N_11195);
and U11424 (N_11424,N_11054,N_11172);
and U11425 (N_11425,N_11092,N_11154);
and U11426 (N_11426,N_11027,N_11100);
nand U11427 (N_11427,N_11065,N_11055);
and U11428 (N_11428,N_11050,N_11076);
or U11429 (N_11429,N_11051,N_11019);
and U11430 (N_11430,N_11150,N_11002);
and U11431 (N_11431,N_11050,N_11215);
nor U11432 (N_11432,N_11089,N_11010);
nor U11433 (N_11433,N_11139,N_11048);
nand U11434 (N_11434,N_11199,N_11048);
nand U11435 (N_11435,N_11127,N_11058);
or U11436 (N_11436,N_11163,N_11037);
nand U11437 (N_11437,N_11107,N_11086);
nor U11438 (N_11438,N_11141,N_11046);
nand U11439 (N_11439,N_11221,N_11096);
nand U11440 (N_11440,N_11035,N_11125);
nand U11441 (N_11441,N_11116,N_11060);
nand U11442 (N_11442,N_11161,N_11241);
and U11443 (N_11443,N_11099,N_11184);
nand U11444 (N_11444,N_11133,N_11242);
or U11445 (N_11445,N_11088,N_11162);
nor U11446 (N_11446,N_11074,N_11018);
nor U11447 (N_11447,N_11174,N_11090);
or U11448 (N_11448,N_11158,N_11068);
xnor U11449 (N_11449,N_11167,N_11228);
nor U11450 (N_11450,N_11125,N_11045);
nand U11451 (N_11451,N_11237,N_11060);
nor U11452 (N_11452,N_11053,N_11148);
nor U11453 (N_11453,N_11220,N_11243);
nand U11454 (N_11454,N_11082,N_11005);
and U11455 (N_11455,N_11056,N_11230);
nand U11456 (N_11456,N_11109,N_11079);
or U11457 (N_11457,N_11040,N_11031);
nor U11458 (N_11458,N_11054,N_11106);
nand U11459 (N_11459,N_11211,N_11016);
nor U11460 (N_11460,N_11120,N_11216);
nand U11461 (N_11461,N_11214,N_11009);
xor U11462 (N_11462,N_11195,N_11218);
or U11463 (N_11463,N_11042,N_11244);
and U11464 (N_11464,N_11147,N_11161);
xor U11465 (N_11465,N_11080,N_11134);
nand U11466 (N_11466,N_11149,N_11074);
xnor U11467 (N_11467,N_11008,N_11115);
nand U11468 (N_11468,N_11004,N_11063);
or U11469 (N_11469,N_11019,N_11244);
and U11470 (N_11470,N_11055,N_11069);
and U11471 (N_11471,N_11036,N_11024);
and U11472 (N_11472,N_11220,N_11211);
and U11473 (N_11473,N_11235,N_11030);
or U11474 (N_11474,N_11147,N_11004);
xnor U11475 (N_11475,N_11185,N_11161);
nor U11476 (N_11476,N_11025,N_11167);
and U11477 (N_11477,N_11171,N_11199);
nand U11478 (N_11478,N_11218,N_11151);
and U11479 (N_11479,N_11224,N_11003);
nor U11480 (N_11480,N_11195,N_11114);
and U11481 (N_11481,N_11161,N_11167);
nor U11482 (N_11482,N_11072,N_11148);
or U11483 (N_11483,N_11235,N_11169);
and U11484 (N_11484,N_11181,N_11081);
and U11485 (N_11485,N_11191,N_11058);
nand U11486 (N_11486,N_11095,N_11132);
nand U11487 (N_11487,N_11246,N_11196);
and U11488 (N_11488,N_11100,N_11123);
or U11489 (N_11489,N_11062,N_11080);
and U11490 (N_11490,N_11048,N_11216);
or U11491 (N_11491,N_11239,N_11162);
or U11492 (N_11492,N_11216,N_11223);
or U11493 (N_11493,N_11107,N_11005);
and U11494 (N_11494,N_11091,N_11107);
and U11495 (N_11495,N_11216,N_11127);
or U11496 (N_11496,N_11124,N_11109);
or U11497 (N_11497,N_11117,N_11244);
or U11498 (N_11498,N_11100,N_11235);
nand U11499 (N_11499,N_11129,N_11093);
or U11500 (N_11500,N_11310,N_11391);
or U11501 (N_11501,N_11339,N_11463);
or U11502 (N_11502,N_11361,N_11259);
or U11503 (N_11503,N_11476,N_11400);
nor U11504 (N_11504,N_11274,N_11434);
xor U11505 (N_11505,N_11395,N_11304);
xnor U11506 (N_11506,N_11328,N_11253);
nand U11507 (N_11507,N_11416,N_11449);
and U11508 (N_11508,N_11473,N_11360);
nand U11509 (N_11509,N_11316,N_11357);
xnor U11510 (N_11510,N_11492,N_11260);
nor U11511 (N_11511,N_11427,N_11294);
and U11512 (N_11512,N_11439,N_11401);
xor U11513 (N_11513,N_11296,N_11290);
and U11514 (N_11514,N_11263,N_11444);
and U11515 (N_11515,N_11415,N_11338);
nor U11516 (N_11516,N_11309,N_11335);
or U11517 (N_11517,N_11433,N_11488);
and U11518 (N_11518,N_11337,N_11467);
and U11519 (N_11519,N_11451,N_11302);
nand U11520 (N_11520,N_11411,N_11375);
or U11521 (N_11521,N_11346,N_11409);
nor U11522 (N_11522,N_11251,N_11311);
and U11523 (N_11523,N_11490,N_11453);
or U11524 (N_11524,N_11368,N_11469);
xnor U11525 (N_11525,N_11455,N_11329);
nand U11526 (N_11526,N_11435,N_11266);
and U11527 (N_11527,N_11327,N_11317);
nor U11528 (N_11528,N_11265,N_11466);
or U11529 (N_11529,N_11477,N_11366);
xor U11530 (N_11530,N_11440,N_11422);
or U11531 (N_11531,N_11254,N_11282);
nor U11532 (N_11532,N_11355,N_11487);
nand U11533 (N_11533,N_11423,N_11273);
nand U11534 (N_11534,N_11456,N_11471);
nand U11535 (N_11535,N_11333,N_11499);
nand U11536 (N_11536,N_11464,N_11445);
or U11537 (N_11537,N_11478,N_11321);
or U11538 (N_11538,N_11402,N_11482);
nor U11539 (N_11539,N_11343,N_11480);
xnor U11540 (N_11540,N_11299,N_11326);
nand U11541 (N_11541,N_11381,N_11481);
and U11542 (N_11542,N_11475,N_11426);
nand U11543 (N_11543,N_11468,N_11261);
and U11544 (N_11544,N_11256,N_11275);
and U11545 (N_11545,N_11379,N_11356);
nand U11546 (N_11546,N_11363,N_11345);
nand U11547 (N_11547,N_11349,N_11407);
xnor U11548 (N_11548,N_11420,N_11399);
and U11549 (N_11549,N_11351,N_11396);
or U11550 (N_11550,N_11287,N_11472);
nand U11551 (N_11551,N_11308,N_11457);
nor U11552 (N_11552,N_11414,N_11257);
nand U11553 (N_11553,N_11285,N_11486);
or U11554 (N_11554,N_11271,N_11315);
or U11555 (N_11555,N_11276,N_11322);
nor U11556 (N_11556,N_11495,N_11268);
or U11557 (N_11557,N_11350,N_11278);
nor U11558 (N_11558,N_11384,N_11448);
and U11559 (N_11559,N_11280,N_11403);
and U11560 (N_11560,N_11485,N_11398);
or U11561 (N_11561,N_11295,N_11437);
nand U11562 (N_11562,N_11497,N_11313);
or U11563 (N_11563,N_11410,N_11293);
and U11564 (N_11564,N_11270,N_11470);
or U11565 (N_11565,N_11291,N_11341);
or U11566 (N_11566,N_11297,N_11412);
nand U11567 (N_11567,N_11306,N_11491);
nand U11568 (N_11568,N_11385,N_11496);
nand U11569 (N_11569,N_11320,N_11374);
nand U11570 (N_11570,N_11460,N_11377);
and U11571 (N_11571,N_11392,N_11283);
or U11572 (N_11572,N_11264,N_11388);
nand U11573 (N_11573,N_11454,N_11429);
or U11574 (N_11574,N_11354,N_11298);
or U11575 (N_11575,N_11277,N_11303);
nand U11576 (N_11576,N_11371,N_11314);
and U11577 (N_11577,N_11347,N_11250);
nor U11578 (N_11578,N_11359,N_11484);
or U11579 (N_11579,N_11408,N_11394);
xnor U11580 (N_11580,N_11438,N_11431);
or U11581 (N_11581,N_11336,N_11332);
nor U11582 (N_11582,N_11331,N_11292);
nor U11583 (N_11583,N_11312,N_11352);
and U11584 (N_11584,N_11413,N_11386);
and U11585 (N_11585,N_11446,N_11289);
and U11586 (N_11586,N_11382,N_11279);
nor U11587 (N_11587,N_11493,N_11325);
nor U11588 (N_11588,N_11380,N_11418);
and U11589 (N_11589,N_11462,N_11281);
or U11590 (N_11590,N_11348,N_11284);
nor U11591 (N_11591,N_11432,N_11483);
nor U11592 (N_11592,N_11334,N_11272);
or U11593 (N_11593,N_11479,N_11362);
or U11594 (N_11594,N_11353,N_11421);
or U11595 (N_11595,N_11269,N_11419);
xnor U11596 (N_11596,N_11404,N_11365);
and U11597 (N_11597,N_11393,N_11342);
nor U11598 (N_11598,N_11465,N_11430);
and U11599 (N_11599,N_11441,N_11425);
and U11600 (N_11600,N_11267,N_11305);
or U11601 (N_11601,N_11376,N_11364);
xnor U11602 (N_11602,N_11417,N_11344);
xor U11603 (N_11603,N_11498,N_11447);
and U11604 (N_11604,N_11340,N_11424);
xor U11605 (N_11605,N_11458,N_11450);
and U11606 (N_11606,N_11436,N_11370);
nor U11607 (N_11607,N_11442,N_11474);
and U11608 (N_11608,N_11369,N_11452);
or U11609 (N_11609,N_11397,N_11258);
or U11610 (N_11610,N_11390,N_11358);
xor U11611 (N_11611,N_11489,N_11405);
nor U11612 (N_11612,N_11286,N_11288);
nor U11613 (N_11613,N_11319,N_11383);
xor U11614 (N_11614,N_11324,N_11300);
or U11615 (N_11615,N_11301,N_11459);
nand U11616 (N_11616,N_11373,N_11378);
and U11617 (N_11617,N_11255,N_11387);
nand U11618 (N_11618,N_11330,N_11323);
nor U11619 (N_11619,N_11318,N_11461);
nand U11620 (N_11620,N_11307,N_11262);
or U11621 (N_11621,N_11428,N_11367);
nor U11622 (N_11622,N_11252,N_11494);
nand U11623 (N_11623,N_11443,N_11372);
and U11624 (N_11624,N_11389,N_11406);
xnor U11625 (N_11625,N_11451,N_11491);
and U11626 (N_11626,N_11299,N_11359);
nor U11627 (N_11627,N_11443,N_11472);
or U11628 (N_11628,N_11478,N_11303);
nand U11629 (N_11629,N_11414,N_11442);
xor U11630 (N_11630,N_11299,N_11350);
nor U11631 (N_11631,N_11377,N_11267);
xnor U11632 (N_11632,N_11412,N_11292);
and U11633 (N_11633,N_11470,N_11352);
nor U11634 (N_11634,N_11430,N_11321);
nand U11635 (N_11635,N_11432,N_11472);
and U11636 (N_11636,N_11284,N_11316);
or U11637 (N_11637,N_11329,N_11268);
or U11638 (N_11638,N_11481,N_11430);
nor U11639 (N_11639,N_11311,N_11394);
nand U11640 (N_11640,N_11263,N_11290);
or U11641 (N_11641,N_11309,N_11456);
nor U11642 (N_11642,N_11360,N_11390);
nor U11643 (N_11643,N_11332,N_11289);
nor U11644 (N_11644,N_11368,N_11364);
and U11645 (N_11645,N_11308,N_11318);
nand U11646 (N_11646,N_11474,N_11377);
nand U11647 (N_11647,N_11499,N_11267);
nor U11648 (N_11648,N_11256,N_11259);
and U11649 (N_11649,N_11353,N_11425);
and U11650 (N_11650,N_11254,N_11498);
and U11651 (N_11651,N_11446,N_11441);
and U11652 (N_11652,N_11433,N_11442);
or U11653 (N_11653,N_11462,N_11433);
nand U11654 (N_11654,N_11273,N_11320);
xor U11655 (N_11655,N_11303,N_11373);
nor U11656 (N_11656,N_11468,N_11453);
nand U11657 (N_11657,N_11494,N_11342);
and U11658 (N_11658,N_11463,N_11396);
xor U11659 (N_11659,N_11292,N_11410);
xor U11660 (N_11660,N_11404,N_11371);
nor U11661 (N_11661,N_11437,N_11359);
nand U11662 (N_11662,N_11390,N_11311);
nand U11663 (N_11663,N_11420,N_11473);
nand U11664 (N_11664,N_11453,N_11250);
or U11665 (N_11665,N_11338,N_11436);
nor U11666 (N_11666,N_11444,N_11276);
nor U11667 (N_11667,N_11498,N_11283);
and U11668 (N_11668,N_11334,N_11490);
nand U11669 (N_11669,N_11293,N_11255);
and U11670 (N_11670,N_11469,N_11265);
nand U11671 (N_11671,N_11452,N_11272);
nand U11672 (N_11672,N_11456,N_11276);
nand U11673 (N_11673,N_11275,N_11469);
and U11674 (N_11674,N_11464,N_11494);
and U11675 (N_11675,N_11424,N_11354);
nor U11676 (N_11676,N_11397,N_11420);
and U11677 (N_11677,N_11313,N_11274);
nand U11678 (N_11678,N_11308,N_11444);
or U11679 (N_11679,N_11324,N_11337);
or U11680 (N_11680,N_11480,N_11291);
nand U11681 (N_11681,N_11280,N_11433);
nor U11682 (N_11682,N_11388,N_11270);
and U11683 (N_11683,N_11293,N_11310);
nand U11684 (N_11684,N_11257,N_11405);
nor U11685 (N_11685,N_11447,N_11383);
or U11686 (N_11686,N_11353,N_11304);
and U11687 (N_11687,N_11395,N_11259);
and U11688 (N_11688,N_11458,N_11296);
or U11689 (N_11689,N_11489,N_11272);
or U11690 (N_11690,N_11408,N_11388);
or U11691 (N_11691,N_11384,N_11435);
xnor U11692 (N_11692,N_11487,N_11349);
nand U11693 (N_11693,N_11260,N_11373);
nor U11694 (N_11694,N_11465,N_11389);
or U11695 (N_11695,N_11339,N_11295);
nor U11696 (N_11696,N_11423,N_11404);
and U11697 (N_11697,N_11310,N_11335);
or U11698 (N_11698,N_11432,N_11453);
and U11699 (N_11699,N_11472,N_11276);
nand U11700 (N_11700,N_11434,N_11460);
or U11701 (N_11701,N_11361,N_11397);
and U11702 (N_11702,N_11479,N_11312);
xnor U11703 (N_11703,N_11279,N_11439);
or U11704 (N_11704,N_11281,N_11277);
nor U11705 (N_11705,N_11436,N_11296);
or U11706 (N_11706,N_11443,N_11325);
nand U11707 (N_11707,N_11424,N_11393);
nand U11708 (N_11708,N_11452,N_11391);
or U11709 (N_11709,N_11417,N_11431);
and U11710 (N_11710,N_11271,N_11477);
or U11711 (N_11711,N_11488,N_11271);
and U11712 (N_11712,N_11264,N_11266);
nor U11713 (N_11713,N_11278,N_11366);
or U11714 (N_11714,N_11332,N_11470);
xor U11715 (N_11715,N_11254,N_11477);
and U11716 (N_11716,N_11458,N_11334);
xnor U11717 (N_11717,N_11399,N_11480);
nor U11718 (N_11718,N_11402,N_11326);
nand U11719 (N_11719,N_11379,N_11257);
and U11720 (N_11720,N_11337,N_11489);
and U11721 (N_11721,N_11285,N_11414);
xor U11722 (N_11722,N_11334,N_11436);
nand U11723 (N_11723,N_11340,N_11277);
nand U11724 (N_11724,N_11275,N_11447);
nor U11725 (N_11725,N_11289,N_11348);
nor U11726 (N_11726,N_11490,N_11309);
nor U11727 (N_11727,N_11406,N_11297);
nor U11728 (N_11728,N_11345,N_11417);
nand U11729 (N_11729,N_11422,N_11476);
xnor U11730 (N_11730,N_11440,N_11488);
nand U11731 (N_11731,N_11474,N_11399);
nor U11732 (N_11732,N_11449,N_11315);
nor U11733 (N_11733,N_11425,N_11492);
nor U11734 (N_11734,N_11475,N_11383);
and U11735 (N_11735,N_11266,N_11433);
nor U11736 (N_11736,N_11407,N_11436);
nor U11737 (N_11737,N_11371,N_11445);
nand U11738 (N_11738,N_11478,N_11397);
or U11739 (N_11739,N_11341,N_11413);
nand U11740 (N_11740,N_11485,N_11419);
nor U11741 (N_11741,N_11413,N_11331);
and U11742 (N_11742,N_11365,N_11321);
or U11743 (N_11743,N_11348,N_11393);
and U11744 (N_11744,N_11453,N_11256);
nand U11745 (N_11745,N_11406,N_11475);
nand U11746 (N_11746,N_11435,N_11380);
nand U11747 (N_11747,N_11312,N_11452);
nand U11748 (N_11748,N_11464,N_11256);
nor U11749 (N_11749,N_11470,N_11347);
nand U11750 (N_11750,N_11617,N_11680);
and U11751 (N_11751,N_11517,N_11555);
or U11752 (N_11752,N_11591,N_11733);
nand U11753 (N_11753,N_11579,N_11737);
nand U11754 (N_11754,N_11572,N_11529);
nand U11755 (N_11755,N_11594,N_11660);
or U11756 (N_11756,N_11741,N_11723);
nand U11757 (N_11757,N_11585,N_11672);
or U11758 (N_11758,N_11716,N_11736);
xnor U11759 (N_11759,N_11726,N_11663);
nand U11760 (N_11760,N_11714,N_11512);
and U11761 (N_11761,N_11728,N_11653);
xor U11762 (N_11762,N_11735,N_11565);
and U11763 (N_11763,N_11605,N_11712);
nand U11764 (N_11764,N_11562,N_11639);
and U11765 (N_11765,N_11671,N_11532);
and U11766 (N_11766,N_11697,N_11646);
or U11767 (N_11767,N_11654,N_11701);
xor U11768 (N_11768,N_11560,N_11742);
or U11769 (N_11769,N_11541,N_11587);
nand U11770 (N_11770,N_11504,N_11502);
or U11771 (N_11771,N_11599,N_11643);
nor U11772 (N_11772,N_11515,N_11583);
and U11773 (N_11773,N_11527,N_11570);
nand U11774 (N_11774,N_11662,N_11530);
nand U11775 (N_11775,N_11507,N_11710);
nand U11776 (N_11776,N_11547,N_11553);
nand U11777 (N_11777,N_11718,N_11727);
nor U11778 (N_11778,N_11632,N_11729);
and U11779 (N_11779,N_11604,N_11719);
nand U11780 (N_11780,N_11650,N_11513);
and U11781 (N_11781,N_11689,N_11704);
nand U11782 (N_11782,N_11577,N_11644);
xor U11783 (N_11783,N_11679,N_11688);
nor U11784 (N_11784,N_11609,N_11593);
or U11785 (N_11785,N_11687,N_11596);
or U11786 (N_11786,N_11534,N_11709);
nor U11787 (N_11787,N_11576,N_11528);
or U11788 (N_11788,N_11563,N_11618);
or U11789 (N_11789,N_11700,N_11738);
and U11790 (N_11790,N_11702,N_11678);
xor U11791 (N_11791,N_11518,N_11721);
nor U11792 (N_11792,N_11612,N_11630);
or U11793 (N_11793,N_11580,N_11645);
nor U11794 (N_11794,N_11543,N_11588);
and U11795 (N_11795,N_11692,N_11717);
nor U11796 (N_11796,N_11656,N_11684);
or U11797 (N_11797,N_11720,N_11564);
and U11798 (N_11798,N_11525,N_11595);
or U11799 (N_11799,N_11607,N_11658);
xor U11800 (N_11800,N_11745,N_11624);
xor U11801 (N_11801,N_11670,N_11623);
nand U11802 (N_11802,N_11606,N_11748);
nor U11803 (N_11803,N_11651,N_11603);
or U11804 (N_11804,N_11707,N_11695);
and U11805 (N_11805,N_11676,N_11584);
or U11806 (N_11806,N_11664,N_11641);
and U11807 (N_11807,N_11608,N_11610);
nor U11808 (N_11808,N_11667,N_11682);
nor U11809 (N_11809,N_11567,N_11637);
xor U11810 (N_11810,N_11743,N_11511);
or U11811 (N_11811,N_11501,N_11559);
or U11812 (N_11812,N_11558,N_11746);
nor U11813 (N_11813,N_11681,N_11642);
nor U11814 (N_11814,N_11536,N_11731);
nand U11815 (N_11815,N_11744,N_11573);
nor U11816 (N_11816,N_11713,N_11524);
nand U11817 (N_11817,N_11503,N_11725);
xnor U11818 (N_11818,N_11626,N_11634);
nor U11819 (N_11819,N_11652,N_11677);
and U11820 (N_11820,N_11538,N_11602);
and U11821 (N_11821,N_11694,N_11699);
nor U11822 (N_11822,N_11581,N_11640);
or U11823 (N_11823,N_11620,N_11537);
nor U11824 (N_11824,N_11698,N_11566);
and U11825 (N_11825,N_11711,N_11522);
nand U11826 (N_11826,N_11638,N_11510);
nor U11827 (N_11827,N_11722,N_11520);
nor U11828 (N_11828,N_11597,N_11685);
nand U11829 (N_11829,N_11589,N_11542);
and U11830 (N_11830,N_11708,N_11552);
nand U11831 (N_11831,N_11519,N_11615);
and U11832 (N_11832,N_11619,N_11673);
xor U11833 (N_11833,N_11613,N_11622);
or U11834 (N_11834,N_11683,N_11705);
nand U11835 (N_11835,N_11732,N_11556);
nand U11836 (N_11836,N_11648,N_11531);
or U11837 (N_11837,N_11533,N_11614);
or U11838 (N_11838,N_11561,N_11675);
or U11839 (N_11839,N_11539,N_11633);
or U11840 (N_11840,N_11516,N_11724);
and U11841 (N_11841,N_11526,N_11569);
and U11842 (N_11842,N_11546,N_11616);
or U11843 (N_11843,N_11739,N_11657);
xor U11844 (N_11844,N_11540,N_11568);
xor U11845 (N_11845,N_11669,N_11600);
xnor U11846 (N_11846,N_11590,N_11635);
nor U11847 (N_11847,N_11575,N_11535);
nand U11848 (N_11848,N_11668,N_11548);
nand U11849 (N_11849,N_11740,N_11598);
and U11850 (N_11850,N_11592,N_11554);
nor U11851 (N_11851,N_11734,N_11523);
and U11852 (N_11852,N_11611,N_11506);
and U11853 (N_11853,N_11747,N_11691);
nor U11854 (N_11854,N_11627,N_11715);
or U11855 (N_11855,N_11549,N_11574);
and U11856 (N_11856,N_11550,N_11508);
and U11857 (N_11857,N_11730,N_11749);
or U11858 (N_11858,N_11690,N_11625);
nand U11859 (N_11859,N_11544,N_11647);
nand U11860 (N_11860,N_11686,N_11514);
nor U11861 (N_11861,N_11557,N_11601);
nor U11862 (N_11862,N_11628,N_11649);
or U11863 (N_11863,N_11655,N_11509);
nor U11864 (N_11864,N_11578,N_11693);
nand U11865 (N_11865,N_11500,N_11706);
nor U11866 (N_11866,N_11661,N_11659);
and U11867 (N_11867,N_11666,N_11621);
and U11868 (N_11868,N_11586,N_11665);
nand U11869 (N_11869,N_11629,N_11505);
or U11870 (N_11870,N_11545,N_11631);
nand U11871 (N_11871,N_11521,N_11674);
nand U11872 (N_11872,N_11582,N_11636);
and U11873 (N_11873,N_11571,N_11696);
xnor U11874 (N_11874,N_11551,N_11703);
nand U11875 (N_11875,N_11697,N_11737);
and U11876 (N_11876,N_11678,N_11657);
or U11877 (N_11877,N_11662,N_11669);
and U11878 (N_11878,N_11650,N_11617);
and U11879 (N_11879,N_11655,N_11623);
or U11880 (N_11880,N_11526,N_11609);
and U11881 (N_11881,N_11536,N_11637);
and U11882 (N_11882,N_11656,N_11710);
nor U11883 (N_11883,N_11565,N_11647);
nor U11884 (N_11884,N_11570,N_11725);
and U11885 (N_11885,N_11596,N_11591);
nor U11886 (N_11886,N_11525,N_11746);
nand U11887 (N_11887,N_11571,N_11644);
nor U11888 (N_11888,N_11689,N_11615);
and U11889 (N_11889,N_11683,N_11570);
and U11890 (N_11890,N_11730,N_11610);
and U11891 (N_11891,N_11726,N_11671);
nor U11892 (N_11892,N_11712,N_11642);
nand U11893 (N_11893,N_11736,N_11605);
and U11894 (N_11894,N_11747,N_11743);
xor U11895 (N_11895,N_11611,N_11641);
nor U11896 (N_11896,N_11594,N_11532);
and U11897 (N_11897,N_11602,N_11603);
nand U11898 (N_11898,N_11579,N_11516);
and U11899 (N_11899,N_11572,N_11530);
and U11900 (N_11900,N_11611,N_11553);
nand U11901 (N_11901,N_11518,N_11643);
nand U11902 (N_11902,N_11570,N_11530);
or U11903 (N_11903,N_11625,N_11643);
nand U11904 (N_11904,N_11727,N_11699);
nor U11905 (N_11905,N_11650,N_11607);
nand U11906 (N_11906,N_11746,N_11734);
and U11907 (N_11907,N_11515,N_11543);
or U11908 (N_11908,N_11514,N_11639);
or U11909 (N_11909,N_11639,N_11699);
nand U11910 (N_11910,N_11604,N_11730);
and U11911 (N_11911,N_11570,N_11738);
nand U11912 (N_11912,N_11730,N_11559);
xnor U11913 (N_11913,N_11679,N_11644);
nor U11914 (N_11914,N_11628,N_11664);
nand U11915 (N_11915,N_11530,N_11666);
xor U11916 (N_11916,N_11525,N_11715);
nor U11917 (N_11917,N_11542,N_11609);
nand U11918 (N_11918,N_11744,N_11612);
or U11919 (N_11919,N_11536,N_11555);
nand U11920 (N_11920,N_11633,N_11561);
nor U11921 (N_11921,N_11741,N_11608);
nor U11922 (N_11922,N_11603,N_11716);
nand U11923 (N_11923,N_11669,N_11714);
and U11924 (N_11924,N_11613,N_11504);
and U11925 (N_11925,N_11610,N_11578);
nor U11926 (N_11926,N_11551,N_11729);
and U11927 (N_11927,N_11734,N_11625);
or U11928 (N_11928,N_11733,N_11631);
nand U11929 (N_11929,N_11519,N_11582);
nand U11930 (N_11930,N_11638,N_11571);
nand U11931 (N_11931,N_11516,N_11675);
or U11932 (N_11932,N_11514,N_11554);
or U11933 (N_11933,N_11648,N_11566);
and U11934 (N_11934,N_11526,N_11574);
and U11935 (N_11935,N_11505,N_11732);
nand U11936 (N_11936,N_11722,N_11537);
nor U11937 (N_11937,N_11534,N_11698);
or U11938 (N_11938,N_11618,N_11559);
nor U11939 (N_11939,N_11670,N_11535);
nor U11940 (N_11940,N_11571,N_11717);
nor U11941 (N_11941,N_11748,N_11719);
and U11942 (N_11942,N_11653,N_11703);
and U11943 (N_11943,N_11623,N_11695);
or U11944 (N_11944,N_11527,N_11708);
and U11945 (N_11945,N_11605,N_11697);
xor U11946 (N_11946,N_11506,N_11615);
and U11947 (N_11947,N_11511,N_11654);
nand U11948 (N_11948,N_11744,N_11504);
nor U11949 (N_11949,N_11721,N_11746);
or U11950 (N_11950,N_11514,N_11615);
nor U11951 (N_11951,N_11527,N_11673);
and U11952 (N_11952,N_11663,N_11534);
nand U11953 (N_11953,N_11655,N_11654);
nand U11954 (N_11954,N_11711,N_11536);
or U11955 (N_11955,N_11580,N_11644);
nand U11956 (N_11956,N_11711,N_11530);
or U11957 (N_11957,N_11551,N_11679);
nor U11958 (N_11958,N_11609,N_11551);
and U11959 (N_11959,N_11554,N_11598);
nor U11960 (N_11960,N_11601,N_11608);
or U11961 (N_11961,N_11629,N_11630);
nor U11962 (N_11962,N_11708,N_11671);
or U11963 (N_11963,N_11599,N_11694);
nand U11964 (N_11964,N_11592,N_11591);
and U11965 (N_11965,N_11542,N_11648);
or U11966 (N_11966,N_11625,N_11527);
nand U11967 (N_11967,N_11505,N_11518);
and U11968 (N_11968,N_11693,N_11590);
and U11969 (N_11969,N_11525,N_11605);
nand U11970 (N_11970,N_11570,N_11661);
or U11971 (N_11971,N_11515,N_11743);
or U11972 (N_11972,N_11743,N_11738);
or U11973 (N_11973,N_11673,N_11571);
nor U11974 (N_11974,N_11651,N_11645);
nand U11975 (N_11975,N_11549,N_11745);
nor U11976 (N_11976,N_11555,N_11560);
nor U11977 (N_11977,N_11504,N_11734);
or U11978 (N_11978,N_11671,N_11636);
or U11979 (N_11979,N_11684,N_11546);
nand U11980 (N_11980,N_11639,N_11540);
or U11981 (N_11981,N_11646,N_11575);
or U11982 (N_11982,N_11524,N_11531);
and U11983 (N_11983,N_11612,N_11737);
nand U11984 (N_11984,N_11685,N_11562);
and U11985 (N_11985,N_11592,N_11593);
or U11986 (N_11986,N_11731,N_11609);
nand U11987 (N_11987,N_11747,N_11648);
or U11988 (N_11988,N_11717,N_11562);
xnor U11989 (N_11989,N_11690,N_11548);
nand U11990 (N_11990,N_11647,N_11668);
xor U11991 (N_11991,N_11691,N_11647);
xnor U11992 (N_11992,N_11680,N_11747);
nor U11993 (N_11993,N_11713,N_11622);
or U11994 (N_11994,N_11590,N_11595);
and U11995 (N_11995,N_11702,N_11745);
and U11996 (N_11996,N_11728,N_11541);
or U11997 (N_11997,N_11731,N_11707);
nor U11998 (N_11998,N_11580,N_11530);
and U11999 (N_11999,N_11587,N_11713);
nor U12000 (N_12000,N_11823,N_11975);
and U12001 (N_12001,N_11919,N_11961);
nor U12002 (N_12002,N_11798,N_11787);
nor U12003 (N_12003,N_11928,N_11771);
xnor U12004 (N_12004,N_11865,N_11825);
nand U12005 (N_12005,N_11855,N_11756);
nor U12006 (N_12006,N_11805,N_11984);
or U12007 (N_12007,N_11964,N_11988);
and U12008 (N_12008,N_11889,N_11973);
nor U12009 (N_12009,N_11772,N_11884);
and U12010 (N_12010,N_11894,N_11819);
nor U12011 (N_12011,N_11836,N_11930);
or U12012 (N_12012,N_11862,N_11763);
or U12013 (N_12013,N_11985,N_11751);
xor U12014 (N_12014,N_11801,N_11790);
or U12015 (N_12015,N_11870,N_11824);
nor U12016 (N_12016,N_11864,N_11886);
nor U12017 (N_12017,N_11812,N_11814);
nor U12018 (N_12018,N_11911,N_11942);
nor U12019 (N_12019,N_11969,N_11829);
nor U12020 (N_12020,N_11784,N_11817);
nand U12021 (N_12021,N_11827,N_11998);
and U12022 (N_12022,N_11932,N_11811);
nor U12023 (N_12023,N_11958,N_11800);
nor U12024 (N_12024,N_11776,N_11978);
nor U12025 (N_12025,N_11910,N_11873);
nor U12026 (N_12026,N_11979,N_11781);
or U12027 (N_12027,N_11766,N_11878);
nand U12028 (N_12028,N_11991,N_11788);
and U12029 (N_12029,N_11774,N_11752);
or U12030 (N_12030,N_11770,N_11931);
or U12031 (N_12031,N_11996,N_11980);
nand U12032 (N_12032,N_11757,N_11780);
or U12033 (N_12033,N_11885,N_11778);
and U12034 (N_12034,N_11833,N_11990);
and U12035 (N_12035,N_11842,N_11891);
or U12036 (N_12036,N_11773,N_11807);
nor U12037 (N_12037,N_11904,N_11963);
or U12038 (N_12038,N_11959,N_11835);
and U12039 (N_12039,N_11848,N_11793);
nand U12040 (N_12040,N_11943,N_11915);
nor U12041 (N_12041,N_11896,N_11949);
and U12042 (N_12042,N_11899,N_11765);
and U12043 (N_12043,N_11857,N_11952);
xor U12044 (N_12044,N_11871,N_11892);
and U12045 (N_12045,N_11913,N_11923);
and U12046 (N_12046,N_11921,N_11883);
or U12047 (N_12047,N_11818,N_11900);
or U12048 (N_12048,N_11982,N_11914);
or U12049 (N_12049,N_11852,N_11951);
nor U12050 (N_12050,N_11834,N_11925);
nor U12051 (N_12051,N_11839,N_11957);
xnor U12052 (N_12052,N_11768,N_11796);
or U12053 (N_12053,N_11755,N_11846);
or U12054 (N_12054,N_11916,N_11926);
nor U12055 (N_12055,N_11820,N_11905);
or U12056 (N_12056,N_11840,N_11940);
nor U12057 (N_12057,N_11950,N_11944);
nand U12058 (N_12058,N_11861,N_11859);
and U12059 (N_12059,N_11815,N_11753);
nand U12060 (N_12060,N_11999,N_11821);
xnor U12061 (N_12061,N_11762,N_11983);
and U12062 (N_12062,N_11795,N_11863);
and U12063 (N_12063,N_11898,N_11809);
nand U12064 (N_12064,N_11803,N_11858);
and U12065 (N_12065,N_11888,N_11764);
or U12066 (N_12066,N_11997,N_11813);
nor U12067 (N_12067,N_11804,N_11927);
nor U12068 (N_12068,N_11956,N_11901);
nand U12069 (N_12069,N_11936,N_11879);
and U12070 (N_12070,N_11977,N_11856);
and U12071 (N_12071,N_11783,N_11989);
and U12072 (N_12072,N_11881,N_11939);
or U12073 (N_12073,N_11994,N_11906);
or U12074 (N_12074,N_11831,N_11971);
and U12075 (N_12075,N_11777,N_11924);
nand U12076 (N_12076,N_11877,N_11887);
xnor U12077 (N_12077,N_11791,N_11967);
nand U12078 (N_12078,N_11941,N_11830);
and U12079 (N_12079,N_11847,N_11938);
and U12080 (N_12080,N_11920,N_11761);
and U12081 (N_12081,N_11841,N_11860);
and U12082 (N_12082,N_11767,N_11785);
and U12083 (N_12083,N_11789,N_11869);
nor U12084 (N_12084,N_11955,N_11912);
and U12085 (N_12085,N_11909,N_11868);
xnor U12086 (N_12086,N_11769,N_11947);
and U12087 (N_12087,N_11972,N_11968);
nor U12088 (N_12088,N_11822,N_11850);
nand U12089 (N_12089,N_11851,N_11876);
and U12090 (N_12090,N_11797,N_11962);
xor U12091 (N_12091,N_11960,N_11775);
or U12092 (N_12092,N_11937,N_11987);
or U12093 (N_12093,N_11872,N_11882);
and U12094 (N_12094,N_11849,N_11837);
nor U12095 (N_12095,N_11945,N_11929);
and U12096 (N_12096,N_11895,N_11953);
nand U12097 (N_12097,N_11810,N_11806);
and U12098 (N_12098,N_11832,N_11802);
and U12099 (N_12099,N_11875,N_11993);
nor U12100 (N_12100,N_11974,N_11897);
nor U12101 (N_12101,N_11792,N_11786);
xor U12102 (N_12102,N_11754,N_11948);
nand U12103 (N_12103,N_11838,N_11907);
and U12104 (N_12104,N_11976,N_11908);
or U12105 (N_12105,N_11760,N_11893);
or U12106 (N_12106,N_11854,N_11808);
nand U12107 (N_12107,N_11965,N_11867);
nand U12108 (N_12108,N_11794,N_11981);
nor U12109 (N_12109,N_11759,N_11954);
xnor U12110 (N_12110,N_11750,N_11917);
nand U12111 (N_12111,N_11992,N_11903);
or U12112 (N_12112,N_11933,N_11866);
and U12113 (N_12113,N_11970,N_11902);
xor U12114 (N_12114,N_11826,N_11779);
or U12115 (N_12115,N_11782,N_11986);
nand U12116 (N_12116,N_11844,N_11995);
nor U12117 (N_12117,N_11874,N_11934);
and U12118 (N_12118,N_11890,N_11816);
nor U12119 (N_12119,N_11799,N_11853);
nor U12120 (N_12120,N_11843,N_11935);
or U12121 (N_12121,N_11918,N_11922);
and U12122 (N_12122,N_11845,N_11946);
nor U12123 (N_12123,N_11828,N_11966);
nor U12124 (N_12124,N_11758,N_11880);
nand U12125 (N_12125,N_11972,N_11875);
xnor U12126 (N_12126,N_11773,N_11847);
nor U12127 (N_12127,N_11803,N_11882);
nand U12128 (N_12128,N_11832,N_11964);
nand U12129 (N_12129,N_11840,N_11934);
and U12130 (N_12130,N_11877,N_11929);
xnor U12131 (N_12131,N_11926,N_11975);
xor U12132 (N_12132,N_11832,N_11817);
or U12133 (N_12133,N_11955,N_11867);
nand U12134 (N_12134,N_11981,N_11882);
and U12135 (N_12135,N_11798,N_11756);
nand U12136 (N_12136,N_11867,N_11953);
or U12137 (N_12137,N_11811,N_11984);
nor U12138 (N_12138,N_11960,N_11805);
and U12139 (N_12139,N_11877,N_11822);
xnor U12140 (N_12140,N_11956,N_11926);
xnor U12141 (N_12141,N_11961,N_11773);
nand U12142 (N_12142,N_11794,N_11983);
or U12143 (N_12143,N_11841,N_11996);
and U12144 (N_12144,N_11928,N_11865);
nor U12145 (N_12145,N_11927,N_11955);
and U12146 (N_12146,N_11849,N_11950);
and U12147 (N_12147,N_11880,N_11906);
nor U12148 (N_12148,N_11769,N_11768);
or U12149 (N_12149,N_11988,N_11887);
and U12150 (N_12150,N_11824,N_11863);
nor U12151 (N_12151,N_11817,N_11934);
nand U12152 (N_12152,N_11756,N_11768);
nor U12153 (N_12153,N_11892,N_11868);
and U12154 (N_12154,N_11943,N_11786);
nand U12155 (N_12155,N_11800,N_11930);
or U12156 (N_12156,N_11790,N_11817);
nand U12157 (N_12157,N_11996,N_11899);
nand U12158 (N_12158,N_11931,N_11984);
nand U12159 (N_12159,N_11816,N_11770);
and U12160 (N_12160,N_11832,N_11822);
nand U12161 (N_12161,N_11894,N_11961);
nor U12162 (N_12162,N_11825,N_11802);
and U12163 (N_12163,N_11951,N_11900);
nand U12164 (N_12164,N_11762,N_11979);
nand U12165 (N_12165,N_11848,N_11925);
and U12166 (N_12166,N_11825,N_11801);
and U12167 (N_12167,N_11970,N_11954);
nor U12168 (N_12168,N_11976,N_11972);
xor U12169 (N_12169,N_11800,N_11871);
and U12170 (N_12170,N_11880,N_11950);
nor U12171 (N_12171,N_11787,N_11882);
and U12172 (N_12172,N_11831,N_11807);
and U12173 (N_12173,N_11757,N_11953);
nand U12174 (N_12174,N_11989,N_11915);
and U12175 (N_12175,N_11856,N_11836);
and U12176 (N_12176,N_11914,N_11881);
or U12177 (N_12177,N_11785,N_11956);
nor U12178 (N_12178,N_11914,N_11853);
nor U12179 (N_12179,N_11759,N_11796);
nand U12180 (N_12180,N_11890,N_11787);
nor U12181 (N_12181,N_11849,N_11904);
or U12182 (N_12182,N_11825,N_11819);
or U12183 (N_12183,N_11893,N_11946);
nand U12184 (N_12184,N_11906,N_11962);
nor U12185 (N_12185,N_11852,N_11793);
or U12186 (N_12186,N_11920,N_11971);
nand U12187 (N_12187,N_11795,N_11784);
nand U12188 (N_12188,N_11880,N_11840);
xnor U12189 (N_12189,N_11903,N_11886);
and U12190 (N_12190,N_11750,N_11768);
or U12191 (N_12191,N_11883,N_11794);
nor U12192 (N_12192,N_11871,N_11897);
xnor U12193 (N_12193,N_11988,N_11994);
or U12194 (N_12194,N_11830,N_11879);
nor U12195 (N_12195,N_11909,N_11750);
nand U12196 (N_12196,N_11861,N_11855);
or U12197 (N_12197,N_11791,N_11952);
nor U12198 (N_12198,N_11761,N_11862);
nand U12199 (N_12199,N_11979,N_11944);
and U12200 (N_12200,N_11997,N_11985);
or U12201 (N_12201,N_11911,N_11874);
nand U12202 (N_12202,N_11949,N_11969);
xor U12203 (N_12203,N_11929,N_11909);
nor U12204 (N_12204,N_11770,N_11927);
nand U12205 (N_12205,N_11771,N_11770);
nor U12206 (N_12206,N_11860,N_11767);
nand U12207 (N_12207,N_11891,N_11952);
xnor U12208 (N_12208,N_11893,N_11896);
nor U12209 (N_12209,N_11976,N_11819);
nor U12210 (N_12210,N_11762,N_11921);
and U12211 (N_12211,N_11874,N_11837);
xnor U12212 (N_12212,N_11911,N_11877);
nor U12213 (N_12213,N_11785,N_11968);
xor U12214 (N_12214,N_11833,N_11937);
nand U12215 (N_12215,N_11795,N_11802);
or U12216 (N_12216,N_11891,N_11968);
nor U12217 (N_12217,N_11794,N_11873);
nand U12218 (N_12218,N_11880,N_11830);
or U12219 (N_12219,N_11933,N_11848);
nand U12220 (N_12220,N_11861,N_11822);
or U12221 (N_12221,N_11820,N_11931);
nor U12222 (N_12222,N_11838,N_11893);
nand U12223 (N_12223,N_11854,N_11951);
xor U12224 (N_12224,N_11867,N_11768);
nor U12225 (N_12225,N_11790,N_11992);
nor U12226 (N_12226,N_11845,N_11950);
and U12227 (N_12227,N_11927,N_11801);
or U12228 (N_12228,N_11929,N_11898);
nor U12229 (N_12229,N_11889,N_11761);
nor U12230 (N_12230,N_11910,N_11957);
nor U12231 (N_12231,N_11822,N_11757);
xnor U12232 (N_12232,N_11769,N_11954);
or U12233 (N_12233,N_11812,N_11839);
nand U12234 (N_12234,N_11953,N_11878);
xor U12235 (N_12235,N_11822,N_11808);
or U12236 (N_12236,N_11925,N_11772);
nor U12237 (N_12237,N_11983,N_11921);
and U12238 (N_12238,N_11835,N_11826);
xnor U12239 (N_12239,N_11996,N_11966);
nand U12240 (N_12240,N_11758,N_11962);
or U12241 (N_12241,N_11881,N_11947);
nand U12242 (N_12242,N_11790,N_11966);
and U12243 (N_12243,N_11856,N_11759);
nor U12244 (N_12244,N_11824,N_11774);
nor U12245 (N_12245,N_11918,N_11996);
xor U12246 (N_12246,N_11782,N_11851);
or U12247 (N_12247,N_11800,N_11917);
and U12248 (N_12248,N_11921,N_11953);
or U12249 (N_12249,N_11959,N_11872);
and U12250 (N_12250,N_12115,N_12172);
or U12251 (N_12251,N_12061,N_12162);
nor U12252 (N_12252,N_12049,N_12021);
nor U12253 (N_12253,N_12089,N_12034);
or U12254 (N_12254,N_12016,N_12243);
nand U12255 (N_12255,N_12093,N_12195);
and U12256 (N_12256,N_12134,N_12232);
nor U12257 (N_12257,N_12221,N_12094);
or U12258 (N_12258,N_12113,N_12000);
nand U12259 (N_12259,N_12152,N_12236);
nor U12260 (N_12260,N_12097,N_12110);
nor U12261 (N_12261,N_12025,N_12071);
or U12262 (N_12262,N_12167,N_12099);
nor U12263 (N_12263,N_12011,N_12072);
nor U12264 (N_12264,N_12193,N_12092);
and U12265 (N_12265,N_12129,N_12111);
nand U12266 (N_12266,N_12009,N_12233);
nand U12267 (N_12267,N_12154,N_12015);
nor U12268 (N_12268,N_12048,N_12216);
and U12269 (N_12269,N_12032,N_12155);
nand U12270 (N_12270,N_12051,N_12191);
nor U12271 (N_12271,N_12106,N_12181);
or U12272 (N_12272,N_12143,N_12166);
or U12273 (N_12273,N_12098,N_12230);
and U12274 (N_12274,N_12180,N_12248);
or U12275 (N_12275,N_12074,N_12184);
nand U12276 (N_12276,N_12133,N_12065);
nor U12277 (N_12277,N_12102,N_12220);
nor U12278 (N_12278,N_12022,N_12038);
and U12279 (N_12279,N_12249,N_12207);
or U12280 (N_12280,N_12068,N_12130);
nor U12281 (N_12281,N_12204,N_12215);
nor U12282 (N_12282,N_12079,N_12235);
and U12283 (N_12283,N_12142,N_12205);
xor U12284 (N_12284,N_12023,N_12218);
or U12285 (N_12285,N_12096,N_12153);
nor U12286 (N_12286,N_12187,N_12137);
xnor U12287 (N_12287,N_12138,N_12222);
nor U12288 (N_12288,N_12241,N_12037);
and U12289 (N_12289,N_12003,N_12202);
nand U12290 (N_12290,N_12196,N_12024);
and U12291 (N_12291,N_12198,N_12183);
nand U12292 (N_12292,N_12045,N_12170);
xor U12293 (N_12293,N_12036,N_12147);
nand U12294 (N_12294,N_12225,N_12064);
nor U12295 (N_12295,N_12059,N_12017);
and U12296 (N_12296,N_12040,N_12151);
nand U12297 (N_12297,N_12208,N_12161);
xnor U12298 (N_12298,N_12116,N_12186);
nor U12299 (N_12299,N_12063,N_12246);
and U12300 (N_12300,N_12135,N_12044);
and U12301 (N_12301,N_12242,N_12231);
xnor U12302 (N_12302,N_12132,N_12131);
and U12303 (N_12303,N_12120,N_12090);
xnor U12304 (N_12304,N_12179,N_12054);
nor U12305 (N_12305,N_12042,N_12041);
xnor U12306 (N_12306,N_12005,N_12101);
nor U12307 (N_12307,N_12019,N_12157);
nand U12308 (N_12308,N_12105,N_12082);
and U12309 (N_12309,N_12095,N_12212);
and U12310 (N_12310,N_12226,N_12109);
and U12311 (N_12311,N_12052,N_12239);
and U12312 (N_12312,N_12006,N_12123);
and U12313 (N_12313,N_12237,N_12192);
nor U12314 (N_12314,N_12209,N_12104);
nor U12315 (N_12315,N_12199,N_12146);
nor U12316 (N_12316,N_12014,N_12211);
and U12317 (N_12317,N_12066,N_12141);
or U12318 (N_12318,N_12185,N_12083);
or U12319 (N_12319,N_12112,N_12050);
xor U12320 (N_12320,N_12013,N_12190);
nor U12321 (N_12321,N_12165,N_12008);
or U12322 (N_12322,N_12245,N_12001);
or U12323 (N_12323,N_12247,N_12229);
or U12324 (N_12324,N_12228,N_12018);
xor U12325 (N_12325,N_12140,N_12163);
nor U12326 (N_12326,N_12053,N_12122);
or U12327 (N_12327,N_12168,N_12121);
or U12328 (N_12328,N_12182,N_12149);
nand U12329 (N_12329,N_12081,N_12035);
or U12330 (N_12330,N_12159,N_12127);
or U12331 (N_12331,N_12238,N_12060);
or U12332 (N_12332,N_12114,N_12224);
nand U12333 (N_12333,N_12136,N_12171);
or U12334 (N_12334,N_12057,N_12164);
nand U12335 (N_12335,N_12145,N_12084);
nor U12336 (N_12336,N_12108,N_12070);
nand U12337 (N_12337,N_12002,N_12177);
nor U12338 (N_12338,N_12214,N_12158);
and U12339 (N_12339,N_12091,N_12088);
xor U12340 (N_12340,N_12128,N_12028);
xor U12341 (N_12341,N_12062,N_12213);
or U12342 (N_12342,N_12039,N_12026);
and U12343 (N_12343,N_12056,N_12124);
xor U12344 (N_12344,N_12139,N_12240);
or U12345 (N_12345,N_12194,N_12103);
nand U12346 (N_12346,N_12227,N_12007);
and U12347 (N_12347,N_12085,N_12033);
nor U12348 (N_12348,N_12169,N_12077);
or U12349 (N_12349,N_12203,N_12117);
nand U12350 (N_12350,N_12118,N_12027);
xor U12351 (N_12351,N_12189,N_12201);
nand U12352 (N_12352,N_12178,N_12075);
nor U12353 (N_12353,N_12217,N_12197);
and U12354 (N_12354,N_12188,N_12029);
nand U12355 (N_12355,N_12156,N_12175);
and U12356 (N_12356,N_12150,N_12030);
or U12357 (N_12357,N_12058,N_12223);
and U12358 (N_12358,N_12047,N_12100);
nor U12359 (N_12359,N_12043,N_12010);
and U12360 (N_12360,N_12012,N_12031);
nand U12361 (N_12361,N_12174,N_12076);
xor U12362 (N_12362,N_12087,N_12176);
and U12363 (N_12363,N_12219,N_12004);
xnor U12364 (N_12364,N_12119,N_12126);
and U12365 (N_12365,N_12210,N_12148);
or U12366 (N_12366,N_12020,N_12055);
nand U12367 (N_12367,N_12160,N_12173);
xnor U12368 (N_12368,N_12125,N_12107);
nor U12369 (N_12369,N_12046,N_12080);
nor U12370 (N_12370,N_12069,N_12234);
and U12371 (N_12371,N_12200,N_12073);
and U12372 (N_12372,N_12086,N_12144);
xor U12373 (N_12373,N_12067,N_12244);
xor U12374 (N_12374,N_12206,N_12078);
or U12375 (N_12375,N_12233,N_12103);
or U12376 (N_12376,N_12181,N_12000);
and U12377 (N_12377,N_12238,N_12128);
nand U12378 (N_12378,N_12069,N_12131);
nand U12379 (N_12379,N_12216,N_12008);
nor U12380 (N_12380,N_12078,N_12192);
and U12381 (N_12381,N_12147,N_12214);
nand U12382 (N_12382,N_12028,N_12110);
and U12383 (N_12383,N_12073,N_12244);
nand U12384 (N_12384,N_12059,N_12196);
nand U12385 (N_12385,N_12225,N_12203);
nand U12386 (N_12386,N_12054,N_12198);
and U12387 (N_12387,N_12174,N_12241);
xnor U12388 (N_12388,N_12037,N_12095);
or U12389 (N_12389,N_12219,N_12039);
nand U12390 (N_12390,N_12006,N_12120);
or U12391 (N_12391,N_12201,N_12144);
or U12392 (N_12392,N_12166,N_12202);
or U12393 (N_12393,N_12017,N_12093);
or U12394 (N_12394,N_12104,N_12103);
nand U12395 (N_12395,N_12104,N_12188);
nor U12396 (N_12396,N_12118,N_12181);
or U12397 (N_12397,N_12110,N_12165);
and U12398 (N_12398,N_12232,N_12009);
nand U12399 (N_12399,N_12064,N_12041);
or U12400 (N_12400,N_12065,N_12220);
nand U12401 (N_12401,N_12017,N_12192);
or U12402 (N_12402,N_12006,N_12105);
xor U12403 (N_12403,N_12018,N_12196);
nand U12404 (N_12404,N_12218,N_12155);
nor U12405 (N_12405,N_12071,N_12165);
nor U12406 (N_12406,N_12228,N_12002);
nor U12407 (N_12407,N_12219,N_12217);
and U12408 (N_12408,N_12165,N_12075);
nand U12409 (N_12409,N_12249,N_12061);
or U12410 (N_12410,N_12093,N_12243);
and U12411 (N_12411,N_12158,N_12130);
and U12412 (N_12412,N_12138,N_12046);
nor U12413 (N_12413,N_12194,N_12200);
and U12414 (N_12414,N_12228,N_12184);
nor U12415 (N_12415,N_12113,N_12001);
nor U12416 (N_12416,N_12190,N_12141);
xor U12417 (N_12417,N_12158,N_12108);
and U12418 (N_12418,N_12154,N_12117);
xnor U12419 (N_12419,N_12195,N_12135);
nor U12420 (N_12420,N_12229,N_12147);
and U12421 (N_12421,N_12171,N_12149);
or U12422 (N_12422,N_12103,N_12102);
or U12423 (N_12423,N_12118,N_12149);
nand U12424 (N_12424,N_12002,N_12089);
nand U12425 (N_12425,N_12133,N_12179);
or U12426 (N_12426,N_12205,N_12236);
nand U12427 (N_12427,N_12215,N_12213);
nand U12428 (N_12428,N_12148,N_12052);
and U12429 (N_12429,N_12212,N_12210);
nand U12430 (N_12430,N_12082,N_12114);
or U12431 (N_12431,N_12175,N_12130);
and U12432 (N_12432,N_12186,N_12084);
nor U12433 (N_12433,N_12226,N_12186);
and U12434 (N_12434,N_12111,N_12103);
and U12435 (N_12435,N_12112,N_12135);
or U12436 (N_12436,N_12099,N_12136);
nand U12437 (N_12437,N_12248,N_12217);
nor U12438 (N_12438,N_12056,N_12189);
and U12439 (N_12439,N_12156,N_12065);
and U12440 (N_12440,N_12084,N_12133);
or U12441 (N_12441,N_12172,N_12122);
xnor U12442 (N_12442,N_12069,N_12006);
xor U12443 (N_12443,N_12013,N_12107);
nor U12444 (N_12444,N_12001,N_12249);
nor U12445 (N_12445,N_12184,N_12248);
nand U12446 (N_12446,N_12166,N_12038);
xor U12447 (N_12447,N_12135,N_12036);
nor U12448 (N_12448,N_12035,N_12145);
nor U12449 (N_12449,N_12237,N_12214);
and U12450 (N_12450,N_12149,N_12227);
nand U12451 (N_12451,N_12115,N_12241);
nand U12452 (N_12452,N_12062,N_12034);
or U12453 (N_12453,N_12170,N_12188);
nor U12454 (N_12454,N_12051,N_12086);
nand U12455 (N_12455,N_12194,N_12011);
and U12456 (N_12456,N_12177,N_12156);
nand U12457 (N_12457,N_12159,N_12017);
xor U12458 (N_12458,N_12027,N_12115);
or U12459 (N_12459,N_12243,N_12069);
nand U12460 (N_12460,N_12009,N_12057);
or U12461 (N_12461,N_12010,N_12047);
nand U12462 (N_12462,N_12150,N_12117);
or U12463 (N_12463,N_12012,N_12186);
nor U12464 (N_12464,N_12242,N_12175);
nor U12465 (N_12465,N_12063,N_12061);
and U12466 (N_12466,N_12127,N_12186);
nor U12467 (N_12467,N_12086,N_12246);
or U12468 (N_12468,N_12248,N_12207);
or U12469 (N_12469,N_12018,N_12192);
nand U12470 (N_12470,N_12100,N_12168);
or U12471 (N_12471,N_12001,N_12152);
and U12472 (N_12472,N_12011,N_12041);
or U12473 (N_12473,N_12038,N_12063);
nor U12474 (N_12474,N_12149,N_12069);
and U12475 (N_12475,N_12208,N_12103);
nand U12476 (N_12476,N_12070,N_12189);
and U12477 (N_12477,N_12073,N_12054);
nor U12478 (N_12478,N_12113,N_12050);
nand U12479 (N_12479,N_12077,N_12143);
nor U12480 (N_12480,N_12142,N_12079);
and U12481 (N_12481,N_12189,N_12034);
and U12482 (N_12482,N_12053,N_12032);
or U12483 (N_12483,N_12169,N_12200);
nand U12484 (N_12484,N_12060,N_12088);
nor U12485 (N_12485,N_12110,N_12176);
or U12486 (N_12486,N_12085,N_12014);
nor U12487 (N_12487,N_12013,N_12134);
nor U12488 (N_12488,N_12134,N_12180);
nand U12489 (N_12489,N_12053,N_12235);
nor U12490 (N_12490,N_12161,N_12152);
or U12491 (N_12491,N_12107,N_12074);
and U12492 (N_12492,N_12003,N_12186);
and U12493 (N_12493,N_12065,N_12014);
and U12494 (N_12494,N_12215,N_12228);
or U12495 (N_12495,N_12056,N_12147);
xor U12496 (N_12496,N_12127,N_12189);
nor U12497 (N_12497,N_12080,N_12036);
xnor U12498 (N_12498,N_12198,N_12017);
and U12499 (N_12499,N_12235,N_12049);
nand U12500 (N_12500,N_12411,N_12495);
and U12501 (N_12501,N_12391,N_12333);
or U12502 (N_12502,N_12463,N_12478);
nand U12503 (N_12503,N_12387,N_12383);
or U12504 (N_12504,N_12279,N_12328);
nand U12505 (N_12505,N_12355,N_12461);
or U12506 (N_12506,N_12464,N_12470);
nand U12507 (N_12507,N_12353,N_12298);
and U12508 (N_12508,N_12402,N_12462);
or U12509 (N_12509,N_12288,N_12335);
and U12510 (N_12510,N_12423,N_12334);
nor U12511 (N_12511,N_12418,N_12499);
or U12512 (N_12512,N_12251,N_12339);
nand U12513 (N_12513,N_12483,N_12290);
nand U12514 (N_12514,N_12451,N_12262);
xnor U12515 (N_12515,N_12364,N_12489);
or U12516 (N_12516,N_12349,N_12322);
or U12517 (N_12517,N_12385,N_12346);
nor U12518 (N_12518,N_12250,N_12321);
and U12519 (N_12519,N_12417,N_12376);
nand U12520 (N_12520,N_12331,N_12413);
nor U12521 (N_12521,N_12458,N_12394);
nand U12522 (N_12522,N_12257,N_12379);
nor U12523 (N_12523,N_12273,N_12443);
or U12524 (N_12524,N_12481,N_12332);
nor U12525 (N_12525,N_12450,N_12432);
and U12526 (N_12526,N_12371,N_12253);
nor U12527 (N_12527,N_12404,N_12338);
and U12528 (N_12528,N_12330,N_12284);
xnor U12529 (N_12529,N_12358,N_12313);
or U12530 (N_12530,N_12434,N_12325);
nor U12531 (N_12531,N_12449,N_12398);
nor U12532 (N_12532,N_12380,N_12366);
nor U12533 (N_12533,N_12405,N_12341);
xor U12534 (N_12534,N_12367,N_12390);
and U12535 (N_12535,N_12302,N_12282);
and U12536 (N_12536,N_12430,N_12269);
nor U12537 (N_12537,N_12497,N_12424);
or U12538 (N_12538,N_12441,N_12280);
or U12539 (N_12539,N_12484,N_12309);
or U12540 (N_12540,N_12392,N_12435);
xor U12541 (N_12541,N_12403,N_12479);
nand U12542 (N_12542,N_12274,N_12293);
nor U12543 (N_12543,N_12393,N_12261);
xor U12544 (N_12544,N_12277,N_12406);
or U12545 (N_12545,N_12471,N_12488);
nor U12546 (N_12546,N_12336,N_12351);
nand U12547 (N_12547,N_12456,N_12347);
and U12548 (N_12548,N_12315,N_12460);
nand U12549 (N_12549,N_12278,N_12490);
nor U12550 (N_12550,N_12276,N_12303);
nor U12551 (N_12551,N_12327,N_12427);
or U12552 (N_12552,N_12452,N_12281);
and U12553 (N_12553,N_12375,N_12305);
nand U12554 (N_12554,N_12388,N_12348);
nand U12555 (N_12555,N_12373,N_12306);
and U12556 (N_12556,N_12421,N_12440);
and U12557 (N_12557,N_12326,N_12468);
and U12558 (N_12558,N_12399,N_12295);
nand U12559 (N_12559,N_12397,N_12473);
and U12560 (N_12560,N_12420,N_12268);
nand U12561 (N_12561,N_12289,N_12267);
nor U12562 (N_12562,N_12485,N_12258);
nand U12563 (N_12563,N_12272,N_12360);
nand U12564 (N_12564,N_12422,N_12363);
nand U12565 (N_12565,N_12439,N_12415);
nor U12566 (N_12566,N_12414,N_12287);
and U12567 (N_12567,N_12445,N_12454);
nor U12568 (N_12568,N_12378,N_12359);
or U12569 (N_12569,N_12476,N_12300);
nand U12570 (N_12570,N_12426,N_12340);
nand U12571 (N_12571,N_12448,N_12386);
xnor U12572 (N_12572,N_12377,N_12316);
nand U12573 (N_12573,N_12304,N_12487);
or U12574 (N_12574,N_12477,N_12362);
or U12575 (N_12575,N_12465,N_12492);
nor U12576 (N_12576,N_12350,N_12264);
nand U12577 (N_12577,N_12395,N_12260);
and U12578 (N_12578,N_12266,N_12354);
and U12579 (N_12579,N_12344,N_12370);
or U12580 (N_12580,N_12412,N_12292);
nand U12581 (N_12581,N_12365,N_12270);
nand U12582 (N_12582,N_12345,N_12431);
or U12583 (N_12583,N_12318,N_12337);
or U12584 (N_12584,N_12283,N_12401);
or U12585 (N_12585,N_12286,N_12444);
and U12586 (N_12586,N_12372,N_12259);
nor U12587 (N_12587,N_12474,N_12410);
or U12588 (N_12588,N_12496,N_12407);
and U12589 (N_12589,N_12312,N_12342);
xnor U12590 (N_12590,N_12408,N_12428);
xor U12591 (N_12591,N_12459,N_12433);
and U12592 (N_12592,N_12447,N_12455);
nor U12593 (N_12593,N_12299,N_12425);
nand U12594 (N_12594,N_12311,N_12466);
nor U12595 (N_12595,N_12446,N_12429);
nor U12596 (N_12596,N_12475,N_12437);
nor U12597 (N_12597,N_12493,N_12482);
and U12598 (N_12598,N_12301,N_12416);
nand U12599 (N_12599,N_12357,N_12494);
nand U12600 (N_12600,N_12369,N_12396);
and U12601 (N_12601,N_12291,N_12419);
nor U12602 (N_12602,N_12384,N_12356);
xor U12603 (N_12603,N_12310,N_12486);
nor U12604 (N_12604,N_12255,N_12480);
and U12605 (N_12605,N_12491,N_12457);
or U12606 (N_12606,N_12314,N_12294);
and U12607 (N_12607,N_12307,N_12498);
xor U12608 (N_12608,N_12368,N_12374);
or U12609 (N_12609,N_12409,N_12469);
nand U12610 (N_12610,N_12275,N_12352);
nor U12611 (N_12611,N_12297,N_12323);
and U12612 (N_12612,N_12453,N_12382);
nor U12613 (N_12613,N_12265,N_12254);
xnor U12614 (N_12614,N_12442,N_12320);
nor U12615 (N_12615,N_12438,N_12308);
nand U12616 (N_12616,N_12285,N_12324);
nand U12617 (N_12617,N_12317,N_12329);
and U12618 (N_12618,N_12319,N_12467);
nor U12619 (N_12619,N_12271,N_12263);
or U12620 (N_12620,N_12296,N_12252);
and U12621 (N_12621,N_12472,N_12381);
nand U12622 (N_12622,N_12436,N_12400);
nor U12623 (N_12623,N_12361,N_12256);
nor U12624 (N_12624,N_12389,N_12343);
and U12625 (N_12625,N_12268,N_12385);
nand U12626 (N_12626,N_12499,N_12402);
nand U12627 (N_12627,N_12462,N_12329);
or U12628 (N_12628,N_12329,N_12324);
and U12629 (N_12629,N_12413,N_12265);
xor U12630 (N_12630,N_12458,N_12353);
and U12631 (N_12631,N_12333,N_12497);
or U12632 (N_12632,N_12488,N_12400);
nor U12633 (N_12633,N_12446,N_12494);
nand U12634 (N_12634,N_12277,N_12313);
nand U12635 (N_12635,N_12482,N_12364);
and U12636 (N_12636,N_12499,N_12257);
xor U12637 (N_12637,N_12387,N_12421);
or U12638 (N_12638,N_12261,N_12381);
nor U12639 (N_12639,N_12486,N_12462);
nor U12640 (N_12640,N_12441,N_12267);
nand U12641 (N_12641,N_12412,N_12433);
nor U12642 (N_12642,N_12269,N_12452);
or U12643 (N_12643,N_12252,N_12366);
nor U12644 (N_12644,N_12455,N_12256);
nand U12645 (N_12645,N_12366,N_12271);
and U12646 (N_12646,N_12270,N_12285);
and U12647 (N_12647,N_12337,N_12356);
and U12648 (N_12648,N_12283,N_12414);
xor U12649 (N_12649,N_12497,N_12319);
nor U12650 (N_12650,N_12481,N_12462);
nand U12651 (N_12651,N_12294,N_12458);
and U12652 (N_12652,N_12258,N_12418);
and U12653 (N_12653,N_12496,N_12255);
nor U12654 (N_12654,N_12430,N_12271);
nand U12655 (N_12655,N_12321,N_12387);
and U12656 (N_12656,N_12496,N_12421);
nand U12657 (N_12657,N_12398,N_12466);
xor U12658 (N_12658,N_12432,N_12351);
or U12659 (N_12659,N_12488,N_12340);
nand U12660 (N_12660,N_12257,N_12437);
nand U12661 (N_12661,N_12425,N_12449);
nor U12662 (N_12662,N_12410,N_12359);
or U12663 (N_12663,N_12362,N_12317);
xnor U12664 (N_12664,N_12340,N_12475);
xnor U12665 (N_12665,N_12322,N_12421);
or U12666 (N_12666,N_12312,N_12261);
xor U12667 (N_12667,N_12250,N_12254);
or U12668 (N_12668,N_12469,N_12472);
nor U12669 (N_12669,N_12495,N_12287);
and U12670 (N_12670,N_12472,N_12255);
and U12671 (N_12671,N_12316,N_12447);
or U12672 (N_12672,N_12464,N_12315);
nand U12673 (N_12673,N_12370,N_12264);
nand U12674 (N_12674,N_12324,N_12411);
or U12675 (N_12675,N_12353,N_12356);
nor U12676 (N_12676,N_12419,N_12394);
or U12677 (N_12677,N_12340,N_12345);
xor U12678 (N_12678,N_12382,N_12430);
nor U12679 (N_12679,N_12393,N_12317);
and U12680 (N_12680,N_12294,N_12499);
nor U12681 (N_12681,N_12376,N_12378);
nor U12682 (N_12682,N_12438,N_12309);
nand U12683 (N_12683,N_12361,N_12460);
or U12684 (N_12684,N_12475,N_12492);
nand U12685 (N_12685,N_12454,N_12429);
xor U12686 (N_12686,N_12457,N_12497);
and U12687 (N_12687,N_12426,N_12489);
nor U12688 (N_12688,N_12412,N_12429);
nand U12689 (N_12689,N_12454,N_12384);
nor U12690 (N_12690,N_12473,N_12491);
and U12691 (N_12691,N_12473,N_12267);
nand U12692 (N_12692,N_12423,N_12405);
nand U12693 (N_12693,N_12494,N_12381);
and U12694 (N_12694,N_12354,N_12369);
nand U12695 (N_12695,N_12495,N_12296);
nor U12696 (N_12696,N_12324,N_12497);
and U12697 (N_12697,N_12440,N_12492);
nand U12698 (N_12698,N_12471,N_12481);
and U12699 (N_12699,N_12351,N_12387);
nor U12700 (N_12700,N_12391,N_12319);
nor U12701 (N_12701,N_12259,N_12462);
or U12702 (N_12702,N_12478,N_12373);
or U12703 (N_12703,N_12445,N_12349);
nor U12704 (N_12704,N_12433,N_12468);
nand U12705 (N_12705,N_12270,N_12499);
xor U12706 (N_12706,N_12323,N_12370);
xnor U12707 (N_12707,N_12283,N_12334);
and U12708 (N_12708,N_12279,N_12294);
and U12709 (N_12709,N_12268,N_12455);
nand U12710 (N_12710,N_12267,N_12427);
and U12711 (N_12711,N_12254,N_12321);
and U12712 (N_12712,N_12252,N_12463);
or U12713 (N_12713,N_12444,N_12431);
or U12714 (N_12714,N_12400,N_12360);
nor U12715 (N_12715,N_12304,N_12295);
nor U12716 (N_12716,N_12271,N_12404);
nor U12717 (N_12717,N_12377,N_12473);
xnor U12718 (N_12718,N_12329,N_12399);
nor U12719 (N_12719,N_12471,N_12474);
nor U12720 (N_12720,N_12320,N_12380);
or U12721 (N_12721,N_12286,N_12284);
xnor U12722 (N_12722,N_12303,N_12369);
nand U12723 (N_12723,N_12391,N_12471);
or U12724 (N_12724,N_12486,N_12484);
and U12725 (N_12725,N_12387,N_12432);
nor U12726 (N_12726,N_12464,N_12460);
nor U12727 (N_12727,N_12453,N_12441);
nor U12728 (N_12728,N_12370,N_12346);
nand U12729 (N_12729,N_12262,N_12327);
or U12730 (N_12730,N_12463,N_12383);
or U12731 (N_12731,N_12342,N_12498);
nor U12732 (N_12732,N_12384,N_12301);
or U12733 (N_12733,N_12347,N_12326);
or U12734 (N_12734,N_12428,N_12371);
and U12735 (N_12735,N_12346,N_12485);
and U12736 (N_12736,N_12268,N_12264);
and U12737 (N_12737,N_12306,N_12415);
or U12738 (N_12738,N_12279,N_12259);
nor U12739 (N_12739,N_12389,N_12455);
nand U12740 (N_12740,N_12337,N_12340);
nand U12741 (N_12741,N_12478,N_12299);
or U12742 (N_12742,N_12258,N_12335);
nor U12743 (N_12743,N_12491,N_12448);
nor U12744 (N_12744,N_12479,N_12415);
and U12745 (N_12745,N_12303,N_12455);
or U12746 (N_12746,N_12375,N_12285);
nand U12747 (N_12747,N_12441,N_12316);
and U12748 (N_12748,N_12256,N_12465);
or U12749 (N_12749,N_12305,N_12254);
and U12750 (N_12750,N_12686,N_12669);
or U12751 (N_12751,N_12697,N_12588);
or U12752 (N_12752,N_12574,N_12571);
nand U12753 (N_12753,N_12609,N_12516);
nor U12754 (N_12754,N_12711,N_12740);
and U12755 (N_12755,N_12533,N_12628);
nor U12756 (N_12756,N_12612,N_12714);
or U12757 (N_12757,N_12739,N_12723);
or U12758 (N_12758,N_12617,N_12730);
nor U12759 (N_12759,N_12576,N_12643);
nand U12760 (N_12760,N_12598,N_12635);
nor U12761 (N_12761,N_12512,N_12713);
nor U12762 (N_12762,N_12554,N_12508);
nor U12763 (N_12763,N_12705,N_12620);
and U12764 (N_12764,N_12606,N_12679);
and U12765 (N_12765,N_12544,N_12710);
nor U12766 (N_12766,N_12636,N_12657);
and U12767 (N_12767,N_12535,N_12590);
nor U12768 (N_12768,N_12532,N_12547);
nor U12769 (N_12769,N_12735,N_12642);
nand U12770 (N_12770,N_12591,N_12717);
or U12771 (N_12771,N_12629,N_12542);
or U12772 (N_12772,N_12649,N_12559);
or U12773 (N_12773,N_12600,N_12731);
or U12774 (N_12774,N_12659,N_12682);
xnor U12775 (N_12775,N_12691,N_12602);
nor U12776 (N_12776,N_12593,N_12651);
xor U12777 (N_12777,N_12644,N_12551);
xor U12778 (N_12778,N_12672,N_12561);
or U12779 (N_12779,N_12673,N_12560);
and U12780 (N_12780,N_12661,N_12652);
and U12781 (N_12781,N_12663,N_12616);
nand U12782 (N_12782,N_12577,N_12684);
nor U12783 (N_12783,N_12678,N_12623);
and U12784 (N_12784,N_12634,N_12614);
and U12785 (N_12785,N_12747,N_12685);
or U12786 (N_12786,N_12683,N_12507);
nand U12787 (N_12787,N_12513,N_12668);
nand U12788 (N_12788,N_12658,N_12514);
or U12789 (N_12789,N_12690,N_12563);
and U12790 (N_12790,N_12648,N_12749);
nand U12791 (N_12791,N_12601,N_12580);
and U12792 (N_12792,N_12693,N_12582);
nand U12793 (N_12793,N_12568,N_12521);
and U12794 (N_12794,N_12696,N_12650);
and U12795 (N_12795,N_12724,N_12646);
nor U12796 (N_12796,N_12564,N_12728);
and U12797 (N_12797,N_12525,N_12587);
xor U12798 (N_12798,N_12742,N_12562);
and U12799 (N_12799,N_12529,N_12708);
nor U12800 (N_12800,N_12594,N_12503);
nor U12801 (N_12801,N_12570,N_12569);
or U12802 (N_12802,N_12639,N_12622);
nand U12803 (N_12803,N_12706,N_12726);
or U12804 (N_12804,N_12527,N_12712);
xnor U12805 (N_12805,N_12611,N_12703);
or U12806 (N_12806,N_12737,N_12545);
or U12807 (N_12807,N_12566,N_12733);
or U12808 (N_12808,N_12548,N_12677);
or U12809 (N_12809,N_12510,N_12653);
nand U12810 (N_12810,N_12715,N_12736);
nand U12811 (N_12811,N_12523,N_12707);
and U12812 (N_12812,N_12665,N_12689);
or U12813 (N_12813,N_12627,N_12725);
and U12814 (N_12814,N_12556,N_12699);
nand U12815 (N_12815,N_12501,N_12667);
nand U12816 (N_12816,N_12505,N_12519);
or U12817 (N_12817,N_12608,N_12709);
or U12818 (N_12818,N_12660,N_12656);
nor U12819 (N_12819,N_12546,N_12687);
nand U12820 (N_12820,N_12702,N_12567);
or U12821 (N_12821,N_12543,N_12654);
or U12822 (N_12822,N_12597,N_12578);
or U12823 (N_12823,N_12721,N_12741);
xor U12824 (N_12824,N_12540,N_12727);
and U12825 (N_12825,N_12671,N_12509);
nor U12826 (N_12826,N_12732,N_12664);
nand U12827 (N_12827,N_12537,N_12719);
and U12828 (N_12828,N_12641,N_12575);
and U12829 (N_12829,N_12729,N_12662);
and U12830 (N_12830,N_12701,N_12638);
nor U12831 (N_12831,N_12655,N_12698);
and U12832 (N_12832,N_12675,N_12637);
or U12833 (N_12833,N_12704,N_12599);
and U12834 (N_12834,N_12688,N_12502);
nand U12835 (N_12835,N_12716,N_12541);
and U12836 (N_12836,N_12674,N_12584);
nor U12837 (N_12837,N_12504,N_12692);
xor U12838 (N_12838,N_12555,N_12645);
and U12839 (N_12839,N_12586,N_12625);
and U12840 (N_12840,N_12557,N_12676);
or U12841 (N_12841,N_12605,N_12734);
nand U12842 (N_12842,N_12518,N_12624);
or U12843 (N_12843,N_12621,N_12500);
xor U12844 (N_12844,N_12630,N_12536);
and U12845 (N_12845,N_12748,N_12528);
nand U12846 (N_12846,N_12596,N_12720);
nand U12847 (N_12847,N_12632,N_12633);
and U12848 (N_12848,N_12680,N_12522);
or U12849 (N_12849,N_12583,N_12613);
and U12850 (N_12850,N_12539,N_12524);
and U12851 (N_12851,N_12681,N_12517);
or U12852 (N_12852,N_12530,N_12534);
nand U12853 (N_12853,N_12552,N_12647);
nor U12854 (N_12854,N_12531,N_12618);
nor U12855 (N_12855,N_12722,N_12589);
nor U12856 (N_12856,N_12515,N_12718);
nor U12857 (N_12857,N_12610,N_12603);
or U12858 (N_12858,N_12549,N_12626);
and U12859 (N_12859,N_12553,N_12666);
nor U12860 (N_12860,N_12670,N_12565);
or U12861 (N_12861,N_12550,N_12595);
or U12862 (N_12862,N_12615,N_12604);
or U12863 (N_12863,N_12694,N_12585);
nor U12864 (N_12864,N_12506,N_12573);
or U12865 (N_12865,N_12607,N_12631);
nor U12866 (N_12866,N_12745,N_12619);
or U12867 (N_12867,N_12640,N_12700);
nand U12868 (N_12868,N_12581,N_12572);
and U12869 (N_12869,N_12526,N_12520);
nor U12870 (N_12870,N_12743,N_12744);
nand U12871 (N_12871,N_12511,N_12746);
xnor U12872 (N_12872,N_12579,N_12558);
xor U12873 (N_12873,N_12538,N_12738);
or U12874 (N_12874,N_12592,N_12695);
nor U12875 (N_12875,N_12726,N_12560);
or U12876 (N_12876,N_12686,N_12665);
nor U12877 (N_12877,N_12613,N_12571);
nor U12878 (N_12878,N_12684,N_12536);
xnor U12879 (N_12879,N_12702,N_12642);
nor U12880 (N_12880,N_12694,N_12680);
xnor U12881 (N_12881,N_12737,N_12745);
nor U12882 (N_12882,N_12513,N_12669);
or U12883 (N_12883,N_12517,N_12621);
xor U12884 (N_12884,N_12502,N_12715);
nand U12885 (N_12885,N_12713,N_12591);
and U12886 (N_12886,N_12721,N_12601);
nand U12887 (N_12887,N_12583,N_12615);
or U12888 (N_12888,N_12516,N_12584);
nor U12889 (N_12889,N_12730,N_12506);
xor U12890 (N_12890,N_12552,N_12544);
nand U12891 (N_12891,N_12698,N_12611);
or U12892 (N_12892,N_12568,N_12507);
and U12893 (N_12893,N_12634,N_12600);
nor U12894 (N_12894,N_12720,N_12669);
and U12895 (N_12895,N_12500,N_12557);
nor U12896 (N_12896,N_12510,N_12635);
nand U12897 (N_12897,N_12519,N_12579);
and U12898 (N_12898,N_12635,N_12693);
and U12899 (N_12899,N_12660,N_12513);
nand U12900 (N_12900,N_12653,N_12716);
nor U12901 (N_12901,N_12527,N_12721);
nand U12902 (N_12902,N_12616,N_12514);
nand U12903 (N_12903,N_12592,N_12616);
or U12904 (N_12904,N_12668,N_12584);
nand U12905 (N_12905,N_12655,N_12523);
and U12906 (N_12906,N_12510,N_12533);
nor U12907 (N_12907,N_12502,N_12555);
or U12908 (N_12908,N_12674,N_12643);
nor U12909 (N_12909,N_12522,N_12735);
nand U12910 (N_12910,N_12697,N_12541);
or U12911 (N_12911,N_12506,N_12582);
and U12912 (N_12912,N_12605,N_12511);
nor U12913 (N_12913,N_12536,N_12702);
or U12914 (N_12914,N_12696,N_12538);
nand U12915 (N_12915,N_12559,N_12612);
or U12916 (N_12916,N_12554,N_12600);
nor U12917 (N_12917,N_12743,N_12579);
or U12918 (N_12918,N_12712,N_12710);
nor U12919 (N_12919,N_12514,N_12668);
nand U12920 (N_12920,N_12537,N_12572);
nand U12921 (N_12921,N_12559,N_12705);
and U12922 (N_12922,N_12723,N_12508);
nor U12923 (N_12923,N_12660,N_12556);
nor U12924 (N_12924,N_12700,N_12669);
or U12925 (N_12925,N_12645,N_12564);
nand U12926 (N_12926,N_12739,N_12695);
or U12927 (N_12927,N_12634,N_12641);
or U12928 (N_12928,N_12578,N_12663);
or U12929 (N_12929,N_12727,N_12596);
nor U12930 (N_12930,N_12665,N_12537);
nor U12931 (N_12931,N_12711,N_12675);
or U12932 (N_12932,N_12702,N_12623);
nor U12933 (N_12933,N_12722,N_12732);
or U12934 (N_12934,N_12638,N_12554);
and U12935 (N_12935,N_12655,N_12552);
xnor U12936 (N_12936,N_12657,N_12509);
xnor U12937 (N_12937,N_12630,N_12743);
and U12938 (N_12938,N_12709,N_12685);
xnor U12939 (N_12939,N_12652,N_12636);
and U12940 (N_12940,N_12743,N_12614);
and U12941 (N_12941,N_12712,N_12601);
or U12942 (N_12942,N_12652,N_12607);
nor U12943 (N_12943,N_12578,N_12509);
nor U12944 (N_12944,N_12707,N_12637);
and U12945 (N_12945,N_12668,N_12617);
xnor U12946 (N_12946,N_12594,N_12635);
and U12947 (N_12947,N_12559,N_12715);
or U12948 (N_12948,N_12747,N_12522);
nor U12949 (N_12949,N_12696,N_12549);
or U12950 (N_12950,N_12536,N_12621);
or U12951 (N_12951,N_12637,N_12666);
and U12952 (N_12952,N_12581,N_12612);
and U12953 (N_12953,N_12655,N_12532);
xor U12954 (N_12954,N_12520,N_12608);
nand U12955 (N_12955,N_12556,N_12670);
or U12956 (N_12956,N_12655,N_12635);
xnor U12957 (N_12957,N_12747,N_12558);
or U12958 (N_12958,N_12621,N_12560);
or U12959 (N_12959,N_12644,N_12646);
and U12960 (N_12960,N_12509,N_12602);
nor U12961 (N_12961,N_12679,N_12517);
or U12962 (N_12962,N_12599,N_12594);
nand U12963 (N_12963,N_12656,N_12659);
nand U12964 (N_12964,N_12607,N_12504);
nand U12965 (N_12965,N_12669,N_12511);
or U12966 (N_12966,N_12604,N_12505);
nor U12967 (N_12967,N_12669,N_12683);
nand U12968 (N_12968,N_12730,N_12557);
or U12969 (N_12969,N_12538,N_12594);
xnor U12970 (N_12970,N_12699,N_12610);
nor U12971 (N_12971,N_12561,N_12690);
xor U12972 (N_12972,N_12595,N_12743);
nor U12973 (N_12973,N_12563,N_12631);
and U12974 (N_12974,N_12579,N_12540);
nand U12975 (N_12975,N_12738,N_12529);
nor U12976 (N_12976,N_12561,N_12659);
nor U12977 (N_12977,N_12621,N_12719);
nand U12978 (N_12978,N_12564,N_12527);
and U12979 (N_12979,N_12653,N_12694);
xor U12980 (N_12980,N_12583,N_12710);
nand U12981 (N_12981,N_12674,N_12594);
xor U12982 (N_12982,N_12546,N_12729);
and U12983 (N_12983,N_12606,N_12702);
nand U12984 (N_12984,N_12523,N_12594);
nor U12985 (N_12985,N_12695,N_12508);
nor U12986 (N_12986,N_12626,N_12530);
and U12987 (N_12987,N_12516,N_12562);
and U12988 (N_12988,N_12568,N_12645);
or U12989 (N_12989,N_12713,N_12596);
or U12990 (N_12990,N_12673,N_12534);
nand U12991 (N_12991,N_12694,N_12541);
nand U12992 (N_12992,N_12692,N_12665);
nor U12993 (N_12993,N_12632,N_12610);
or U12994 (N_12994,N_12542,N_12582);
nand U12995 (N_12995,N_12741,N_12688);
or U12996 (N_12996,N_12667,N_12543);
and U12997 (N_12997,N_12502,N_12634);
or U12998 (N_12998,N_12583,N_12684);
nor U12999 (N_12999,N_12749,N_12707);
or U13000 (N_13000,N_12990,N_12809);
or U13001 (N_13001,N_12754,N_12880);
or U13002 (N_13002,N_12875,N_12854);
nor U13003 (N_13003,N_12763,N_12975);
or U13004 (N_13004,N_12773,N_12852);
nor U13005 (N_13005,N_12891,N_12766);
or U13006 (N_13006,N_12853,N_12983);
nor U13007 (N_13007,N_12834,N_12783);
nand U13008 (N_13008,N_12966,N_12985);
nor U13009 (N_13009,N_12930,N_12770);
or U13010 (N_13010,N_12866,N_12776);
nor U13011 (N_13011,N_12786,N_12845);
or U13012 (N_13012,N_12810,N_12860);
nor U13013 (N_13013,N_12818,N_12937);
nor U13014 (N_13014,N_12806,N_12790);
nor U13015 (N_13015,N_12795,N_12992);
nand U13016 (N_13016,N_12752,N_12898);
and U13017 (N_13017,N_12914,N_12904);
nand U13018 (N_13018,N_12791,N_12878);
nand U13019 (N_13019,N_12807,N_12986);
and U13020 (N_13020,N_12855,N_12824);
nor U13021 (N_13021,N_12906,N_12826);
nor U13022 (N_13022,N_12756,N_12915);
and U13023 (N_13023,N_12829,N_12760);
nor U13024 (N_13024,N_12989,N_12903);
nand U13025 (N_13025,N_12831,N_12902);
nand U13026 (N_13026,N_12982,N_12821);
nor U13027 (N_13027,N_12883,N_12832);
and U13028 (N_13028,N_12941,N_12779);
nor U13029 (N_13029,N_12792,N_12888);
nand U13030 (N_13030,N_12976,N_12830);
or U13031 (N_13031,N_12996,N_12957);
xnor U13032 (N_13032,N_12840,N_12789);
and U13033 (N_13033,N_12784,N_12774);
or U13034 (N_13034,N_12936,N_12965);
or U13035 (N_13035,N_12884,N_12961);
or U13036 (N_13036,N_12767,N_12970);
and U13037 (N_13037,N_12950,N_12951);
and U13038 (N_13038,N_12920,N_12839);
xnor U13039 (N_13039,N_12939,N_12847);
nor U13040 (N_13040,N_12843,N_12799);
and U13041 (N_13041,N_12999,N_12935);
nand U13042 (N_13042,N_12922,N_12775);
xor U13043 (N_13043,N_12900,N_12955);
or U13044 (N_13044,N_12962,N_12988);
or U13045 (N_13045,N_12872,N_12960);
nand U13046 (N_13046,N_12871,N_12850);
and U13047 (N_13047,N_12894,N_12828);
nor U13048 (N_13048,N_12817,N_12924);
and U13049 (N_13049,N_12921,N_12816);
and U13050 (N_13050,N_12946,N_12814);
nor U13051 (N_13051,N_12858,N_12907);
nand U13052 (N_13052,N_12943,N_12812);
xnor U13053 (N_13053,N_12971,N_12905);
or U13054 (N_13054,N_12833,N_12873);
nand U13055 (N_13055,N_12750,N_12893);
xor U13056 (N_13056,N_12849,N_12802);
nor U13057 (N_13057,N_12808,N_12993);
or U13058 (N_13058,N_12972,N_12815);
and U13059 (N_13059,N_12846,N_12864);
nor U13060 (N_13060,N_12890,N_12781);
nand U13061 (N_13061,N_12796,N_12822);
nand U13062 (N_13062,N_12956,N_12811);
and U13063 (N_13063,N_12844,N_12753);
nand U13064 (N_13064,N_12889,N_12793);
nor U13065 (N_13065,N_12819,N_12994);
or U13066 (N_13066,N_12835,N_12798);
nand U13067 (N_13067,N_12868,N_12899);
or U13068 (N_13068,N_12842,N_12895);
or U13069 (N_13069,N_12954,N_12948);
and U13070 (N_13070,N_12979,N_12967);
and U13071 (N_13071,N_12977,N_12931);
and U13072 (N_13072,N_12813,N_12757);
and U13073 (N_13073,N_12919,N_12928);
nand U13074 (N_13074,N_12938,N_12780);
nand U13075 (N_13075,N_12927,N_12772);
and U13076 (N_13076,N_12778,N_12803);
xor U13077 (N_13077,N_12874,N_12917);
or U13078 (N_13078,N_12765,N_12925);
nand U13079 (N_13079,N_12908,N_12859);
or U13080 (N_13080,N_12952,N_12885);
or U13081 (N_13081,N_12998,N_12877);
nand U13082 (N_13082,N_12973,N_12929);
or U13083 (N_13083,N_12782,N_12947);
nand U13084 (N_13084,N_12823,N_12837);
or U13085 (N_13085,N_12879,N_12851);
nor U13086 (N_13086,N_12794,N_12987);
nand U13087 (N_13087,N_12882,N_12926);
nor U13088 (N_13088,N_12755,N_12841);
or U13089 (N_13089,N_12887,N_12969);
nor U13090 (N_13090,N_12838,N_12861);
xor U13091 (N_13091,N_12945,N_12862);
and U13092 (N_13092,N_12964,N_12827);
nand U13093 (N_13093,N_12892,N_12764);
and U13094 (N_13094,N_12916,N_12785);
and U13095 (N_13095,N_12881,N_12953);
and U13096 (N_13096,N_12801,N_12857);
and U13097 (N_13097,N_12804,N_12869);
or U13098 (N_13098,N_12797,N_12771);
nor U13099 (N_13099,N_12949,N_12896);
or U13100 (N_13100,N_12758,N_12913);
and U13101 (N_13101,N_12867,N_12805);
and U13102 (N_13102,N_12912,N_12968);
or U13103 (N_13103,N_12777,N_12787);
nor U13104 (N_13104,N_12769,N_12980);
or U13105 (N_13105,N_12958,N_12768);
nand U13106 (N_13106,N_12911,N_12909);
or U13107 (N_13107,N_12856,N_12978);
or U13108 (N_13108,N_12981,N_12933);
and U13109 (N_13109,N_12910,N_12901);
nor U13110 (N_13110,N_12940,N_12886);
nand U13111 (N_13111,N_12974,N_12942);
and U13112 (N_13112,N_12932,N_12865);
xnor U13113 (N_13113,N_12997,N_12800);
nor U13114 (N_13114,N_12820,N_12836);
nor U13115 (N_13115,N_12963,N_12934);
or U13116 (N_13116,N_12918,N_12959);
nor U13117 (N_13117,N_12863,N_12788);
or U13118 (N_13118,N_12870,N_12944);
or U13119 (N_13119,N_12991,N_12984);
and U13120 (N_13120,N_12825,N_12897);
and U13121 (N_13121,N_12751,N_12848);
xor U13122 (N_13122,N_12995,N_12923);
xor U13123 (N_13123,N_12761,N_12759);
and U13124 (N_13124,N_12762,N_12876);
nand U13125 (N_13125,N_12788,N_12777);
and U13126 (N_13126,N_12804,N_12750);
nor U13127 (N_13127,N_12868,N_12948);
and U13128 (N_13128,N_12938,N_12891);
xor U13129 (N_13129,N_12945,N_12986);
and U13130 (N_13130,N_12890,N_12902);
or U13131 (N_13131,N_12963,N_12943);
nor U13132 (N_13132,N_12795,N_12750);
and U13133 (N_13133,N_12786,N_12793);
nor U13134 (N_13134,N_12888,N_12795);
xor U13135 (N_13135,N_12809,N_12938);
or U13136 (N_13136,N_12887,N_12815);
nand U13137 (N_13137,N_12821,N_12894);
nor U13138 (N_13138,N_12960,N_12888);
nand U13139 (N_13139,N_12922,N_12899);
and U13140 (N_13140,N_12842,N_12820);
xor U13141 (N_13141,N_12858,N_12797);
nand U13142 (N_13142,N_12966,N_12930);
or U13143 (N_13143,N_12808,N_12909);
and U13144 (N_13144,N_12777,N_12853);
nand U13145 (N_13145,N_12768,N_12976);
and U13146 (N_13146,N_12892,N_12818);
and U13147 (N_13147,N_12932,N_12761);
nor U13148 (N_13148,N_12910,N_12877);
and U13149 (N_13149,N_12989,N_12971);
and U13150 (N_13150,N_12921,N_12941);
or U13151 (N_13151,N_12929,N_12792);
nand U13152 (N_13152,N_12811,N_12906);
nand U13153 (N_13153,N_12951,N_12900);
nor U13154 (N_13154,N_12789,N_12956);
nand U13155 (N_13155,N_12979,N_12857);
xor U13156 (N_13156,N_12809,N_12860);
or U13157 (N_13157,N_12770,N_12988);
and U13158 (N_13158,N_12832,N_12946);
or U13159 (N_13159,N_12933,N_12799);
and U13160 (N_13160,N_12866,N_12881);
xor U13161 (N_13161,N_12808,N_12786);
and U13162 (N_13162,N_12858,N_12810);
nor U13163 (N_13163,N_12982,N_12971);
nor U13164 (N_13164,N_12836,N_12974);
and U13165 (N_13165,N_12822,N_12927);
nand U13166 (N_13166,N_12927,N_12784);
nor U13167 (N_13167,N_12986,N_12768);
nor U13168 (N_13168,N_12784,N_12766);
and U13169 (N_13169,N_12845,N_12963);
nand U13170 (N_13170,N_12931,N_12916);
nor U13171 (N_13171,N_12986,N_12755);
nand U13172 (N_13172,N_12881,N_12967);
or U13173 (N_13173,N_12935,N_12991);
and U13174 (N_13174,N_12764,N_12933);
and U13175 (N_13175,N_12752,N_12810);
and U13176 (N_13176,N_12983,N_12776);
nor U13177 (N_13177,N_12981,N_12998);
and U13178 (N_13178,N_12927,N_12945);
nor U13179 (N_13179,N_12979,N_12894);
and U13180 (N_13180,N_12834,N_12936);
nand U13181 (N_13181,N_12829,N_12821);
or U13182 (N_13182,N_12906,N_12951);
nor U13183 (N_13183,N_12828,N_12983);
xnor U13184 (N_13184,N_12832,N_12863);
or U13185 (N_13185,N_12977,N_12968);
nor U13186 (N_13186,N_12965,N_12759);
nor U13187 (N_13187,N_12959,N_12992);
nand U13188 (N_13188,N_12858,N_12958);
xnor U13189 (N_13189,N_12986,N_12884);
xor U13190 (N_13190,N_12939,N_12768);
or U13191 (N_13191,N_12940,N_12800);
and U13192 (N_13192,N_12887,N_12997);
and U13193 (N_13193,N_12821,N_12928);
nand U13194 (N_13194,N_12787,N_12778);
nand U13195 (N_13195,N_12940,N_12912);
or U13196 (N_13196,N_12757,N_12933);
nand U13197 (N_13197,N_12792,N_12761);
or U13198 (N_13198,N_12872,N_12785);
nand U13199 (N_13199,N_12805,N_12974);
and U13200 (N_13200,N_12804,N_12935);
or U13201 (N_13201,N_12919,N_12995);
nand U13202 (N_13202,N_12779,N_12757);
or U13203 (N_13203,N_12897,N_12816);
nand U13204 (N_13204,N_12935,N_12771);
nor U13205 (N_13205,N_12841,N_12978);
nor U13206 (N_13206,N_12788,N_12999);
and U13207 (N_13207,N_12756,N_12911);
and U13208 (N_13208,N_12990,N_12798);
or U13209 (N_13209,N_12946,N_12840);
or U13210 (N_13210,N_12798,N_12795);
and U13211 (N_13211,N_12998,N_12815);
or U13212 (N_13212,N_12991,N_12961);
and U13213 (N_13213,N_12776,N_12913);
nor U13214 (N_13214,N_12907,N_12932);
and U13215 (N_13215,N_12906,N_12910);
and U13216 (N_13216,N_12767,N_12803);
and U13217 (N_13217,N_12929,N_12978);
nor U13218 (N_13218,N_12814,N_12970);
nor U13219 (N_13219,N_12773,N_12944);
nand U13220 (N_13220,N_12784,N_12825);
or U13221 (N_13221,N_12954,N_12800);
and U13222 (N_13222,N_12945,N_12771);
nor U13223 (N_13223,N_12799,N_12898);
or U13224 (N_13224,N_12937,N_12925);
and U13225 (N_13225,N_12981,N_12918);
or U13226 (N_13226,N_12762,N_12790);
nor U13227 (N_13227,N_12915,N_12831);
nand U13228 (N_13228,N_12968,N_12859);
or U13229 (N_13229,N_12756,N_12822);
nand U13230 (N_13230,N_12964,N_12887);
and U13231 (N_13231,N_12919,N_12751);
or U13232 (N_13232,N_12765,N_12892);
or U13233 (N_13233,N_12845,N_12921);
xor U13234 (N_13234,N_12876,N_12786);
or U13235 (N_13235,N_12828,N_12888);
or U13236 (N_13236,N_12904,N_12841);
nor U13237 (N_13237,N_12815,N_12857);
nor U13238 (N_13238,N_12874,N_12855);
xor U13239 (N_13239,N_12928,N_12981);
nor U13240 (N_13240,N_12966,N_12998);
nand U13241 (N_13241,N_12955,N_12792);
nor U13242 (N_13242,N_12987,N_12770);
or U13243 (N_13243,N_12958,N_12972);
nor U13244 (N_13244,N_12879,N_12771);
nor U13245 (N_13245,N_12891,N_12932);
and U13246 (N_13246,N_12923,N_12848);
nor U13247 (N_13247,N_12892,N_12796);
or U13248 (N_13248,N_12796,N_12869);
xnor U13249 (N_13249,N_12868,N_12820);
or U13250 (N_13250,N_13044,N_13229);
nand U13251 (N_13251,N_13064,N_13002);
or U13252 (N_13252,N_13100,N_13206);
nor U13253 (N_13253,N_13190,N_13033);
or U13254 (N_13254,N_13234,N_13209);
nor U13255 (N_13255,N_13088,N_13056);
or U13256 (N_13256,N_13014,N_13141);
nor U13257 (N_13257,N_13243,N_13222);
and U13258 (N_13258,N_13197,N_13115);
or U13259 (N_13259,N_13000,N_13245);
or U13260 (N_13260,N_13193,N_13099);
or U13261 (N_13261,N_13181,N_13173);
xor U13262 (N_13262,N_13031,N_13246);
xnor U13263 (N_13263,N_13248,N_13108);
xor U13264 (N_13264,N_13066,N_13138);
or U13265 (N_13265,N_13109,N_13172);
nor U13266 (N_13266,N_13210,N_13208);
nand U13267 (N_13267,N_13244,N_13156);
nor U13268 (N_13268,N_13140,N_13231);
nand U13269 (N_13269,N_13089,N_13082);
nand U13270 (N_13270,N_13015,N_13105);
xnor U13271 (N_13271,N_13101,N_13226);
and U13272 (N_13272,N_13004,N_13154);
nand U13273 (N_13273,N_13071,N_13011);
and U13274 (N_13274,N_13084,N_13073);
and U13275 (N_13275,N_13152,N_13218);
and U13276 (N_13276,N_13185,N_13035);
nand U13277 (N_13277,N_13180,N_13125);
and U13278 (N_13278,N_13155,N_13060);
nor U13279 (N_13279,N_13232,N_13238);
or U13280 (N_13280,N_13239,N_13079);
and U13281 (N_13281,N_13047,N_13030);
or U13282 (N_13282,N_13203,N_13070);
nor U13283 (N_13283,N_13083,N_13116);
xor U13284 (N_13284,N_13114,N_13055);
nor U13285 (N_13285,N_13147,N_13110);
and U13286 (N_13286,N_13215,N_13166);
xnor U13287 (N_13287,N_13168,N_13098);
xnor U13288 (N_13288,N_13202,N_13205);
nand U13289 (N_13289,N_13135,N_13150);
nor U13290 (N_13290,N_13103,N_13224);
or U13291 (N_13291,N_13176,N_13221);
nand U13292 (N_13292,N_13167,N_13007);
and U13293 (N_13293,N_13001,N_13008);
xor U13294 (N_13294,N_13050,N_13042);
and U13295 (N_13295,N_13131,N_13249);
or U13296 (N_13296,N_13021,N_13187);
nor U13297 (N_13297,N_13092,N_13217);
xor U13298 (N_13298,N_13093,N_13120);
and U13299 (N_13299,N_13069,N_13183);
and U13300 (N_13300,N_13123,N_13024);
nor U13301 (N_13301,N_13113,N_13121);
or U13302 (N_13302,N_13219,N_13195);
xnor U13303 (N_13303,N_13143,N_13199);
or U13304 (N_13304,N_13170,N_13177);
nor U13305 (N_13305,N_13133,N_13171);
or U13306 (N_13306,N_13091,N_13200);
or U13307 (N_13307,N_13020,N_13028);
nor U13308 (N_13308,N_13142,N_13151);
and U13309 (N_13309,N_13097,N_13068);
nand U13310 (N_13310,N_13159,N_13049);
nand U13311 (N_13311,N_13085,N_13111);
or U13312 (N_13312,N_13204,N_13130);
xor U13313 (N_13313,N_13017,N_13240);
and U13314 (N_13314,N_13016,N_13037);
nor U13315 (N_13315,N_13201,N_13126);
and U13316 (N_13316,N_13189,N_13134);
nand U13317 (N_13317,N_13019,N_13074);
and U13318 (N_13318,N_13128,N_13160);
and U13319 (N_13319,N_13146,N_13072);
or U13320 (N_13320,N_13078,N_13077);
nor U13321 (N_13321,N_13026,N_13090);
nor U13322 (N_13322,N_13059,N_13118);
and U13323 (N_13323,N_13198,N_13018);
nor U13324 (N_13324,N_13003,N_13153);
and U13325 (N_13325,N_13043,N_13162);
and U13326 (N_13326,N_13212,N_13122);
nor U13327 (N_13327,N_13235,N_13242);
nor U13328 (N_13328,N_13196,N_13223);
and U13329 (N_13329,N_13048,N_13006);
and U13330 (N_13330,N_13192,N_13013);
nor U13331 (N_13331,N_13054,N_13080);
or U13332 (N_13332,N_13136,N_13061);
or U13333 (N_13333,N_13157,N_13076);
nor U13334 (N_13334,N_13023,N_13102);
and U13335 (N_13335,N_13241,N_13225);
nor U13336 (N_13336,N_13165,N_13233);
or U13337 (N_13337,N_13075,N_13194);
and U13338 (N_13338,N_13032,N_13036);
nand U13339 (N_13339,N_13164,N_13216);
xor U13340 (N_13340,N_13087,N_13041);
and U13341 (N_13341,N_13247,N_13058);
and U13342 (N_13342,N_13228,N_13094);
or U13343 (N_13343,N_13174,N_13038);
nand U13344 (N_13344,N_13095,N_13179);
or U13345 (N_13345,N_13186,N_13107);
or U13346 (N_13346,N_13149,N_13227);
nand U13347 (N_13347,N_13034,N_13057);
and U13348 (N_13348,N_13139,N_13161);
and U13349 (N_13349,N_13175,N_13052);
nor U13350 (N_13350,N_13022,N_13096);
and U13351 (N_13351,N_13065,N_13067);
nand U13352 (N_13352,N_13039,N_13040);
nand U13353 (N_13353,N_13112,N_13062);
nand U13354 (N_13354,N_13005,N_13163);
xnor U13355 (N_13355,N_13027,N_13051);
nor U13356 (N_13356,N_13188,N_13009);
xnor U13357 (N_13357,N_13220,N_13086);
nor U13358 (N_13358,N_13063,N_13211);
nand U13359 (N_13359,N_13129,N_13137);
or U13360 (N_13360,N_13045,N_13207);
nor U13361 (N_13361,N_13132,N_13237);
nand U13362 (N_13362,N_13010,N_13119);
nor U13363 (N_13363,N_13158,N_13104);
nand U13364 (N_13364,N_13117,N_13127);
and U13365 (N_13365,N_13213,N_13029);
or U13366 (N_13366,N_13145,N_13148);
or U13367 (N_13367,N_13012,N_13182);
or U13368 (N_13368,N_13230,N_13124);
nand U13369 (N_13369,N_13081,N_13144);
and U13370 (N_13370,N_13025,N_13214);
and U13371 (N_13371,N_13184,N_13053);
nand U13372 (N_13372,N_13191,N_13046);
nor U13373 (N_13373,N_13178,N_13169);
nor U13374 (N_13374,N_13106,N_13236);
and U13375 (N_13375,N_13235,N_13202);
nor U13376 (N_13376,N_13021,N_13056);
xor U13377 (N_13377,N_13044,N_13118);
nand U13378 (N_13378,N_13047,N_13180);
nor U13379 (N_13379,N_13219,N_13041);
and U13380 (N_13380,N_13070,N_13228);
nand U13381 (N_13381,N_13070,N_13231);
nor U13382 (N_13382,N_13196,N_13076);
and U13383 (N_13383,N_13242,N_13143);
nor U13384 (N_13384,N_13148,N_13207);
or U13385 (N_13385,N_13078,N_13049);
and U13386 (N_13386,N_13092,N_13093);
nand U13387 (N_13387,N_13180,N_13202);
nor U13388 (N_13388,N_13101,N_13033);
nor U13389 (N_13389,N_13095,N_13076);
or U13390 (N_13390,N_13208,N_13085);
or U13391 (N_13391,N_13079,N_13169);
nor U13392 (N_13392,N_13095,N_13121);
and U13393 (N_13393,N_13171,N_13184);
nand U13394 (N_13394,N_13241,N_13202);
nor U13395 (N_13395,N_13160,N_13009);
xnor U13396 (N_13396,N_13111,N_13175);
and U13397 (N_13397,N_13128,N_13165);
nand U13398 (N_13398,N_13123,N_13107);
nor U13399 (N_13399,N_13220,N_13196);
nand U13400 (N_13400,N_13052,N_13151);
nor U13401 (N_13401,N_13149,N_13231);
nand U13402 (N_13402,N_13137,N_13143);
and U13403 (N_13403,N_13225,N_13193);
and U13404 (N_13404,N_13094,N_13234);
nor U13405 (N_13405,N_13191,N_13162);
and U13406 (N_13406,N_13055,N_13144);
nor U13407 (N_13407,N_13132,N_13022);
nor U13408 (N_13408,N_13158,N_13185);
or U13409 (N_13409,N_13060,N_13059);
and U13410 (N_13410,N_13152,N_13170);
and U13411 (N_13411,N_13088,N_13203);
xor U13412 (N_13412,N_13229,N_13083);
nand U13413 (N_13413,N_13021,N_13165);
xnor U13414 (N_13414,N_13232,N_13202);
nor U13415 (N_13415,N_13011,N_13245);
xor U13416 (N_13416,N_13039,N_13082);
and U13417 (N_13417,N_13197,N_13153);
nor U13418 (N_13418,N_13074,N_13042);
or U13419 (N_13419,N_13159,N_13193);
nand U13420 (N_13420,N_13215,N_13155);
or U13421 (N_13421,N_13049,N_13149);
nand U13422 (N_13422,N_13069,N_13117);
nand U13423 (N_13423,N_13183,N_13075);
and U13424 (N_13424,N_13240,N_13179);
xor U13425 (N_13425,N_13019,N_13083);
nor U13426 (N_13426,N_13078,N_13101);
xor U13427 (N_13427,N_13106,N_13055);
nor U13428 (N_13428,N_13036,N_13133);
or U13429 (N_13429,N_13194,N_13101);
nand U13430 (N_13430,N_13093,N_13037);
and U13431 (N_13431,N_13216,N_13133);
nor U13432 (N_13432,N_13083,N_13122);
and U13433 (N_13433,N_13057,N_13032);
and U13434 (N_13434,N_13241,N_13154);
and U13435 (N_13435,N_13181,N_13148);
nor U13436 (N_13436,N_13169,N_13031);
nor U13437 (N_13437,N_13099,N_13022);
or U13438 (N_13438,N_13032,N_13196);
xnor U13439 (N_13439,N_13055,N_13139);
xor U13440 (N_13440,N_13027,N_13079);
or U13441 (N_13441,N_13073,N_13172);
or U13442 (N_13442,N_13013,N_13014);
nor U13443 (N_13443,N_13144,N_13099);
nand U13444 (N_13444,N_13109,N_13054);
nor U13445 (N_13445,N_13123,N_13109);
nor U13446 (N_13446,N_13235,N_13198);
nor U13447 (N_13447,N_13139,N_13217);
nor U13448 (N_13448,N_13140,N_13122);
nor U13449 (N_13449,N_13052,N_13098);
or U13450 (N_13450,N_13203,N_13191);
nor U13451 (N_13451,N_13080,N_13043);
and U13452 (N_13452,N_13105,N_13163);
nand U13453 (N_13453,N_13114,N_13049);
nand U13454 (N_13454,N_13073,N_13009);
and U13455 (N_13455,N_13110,N_13220);
nor U13456 (N_13456,N_13142,N_13025);
nor U13457 (N_13457,N_13235,N_13164);
nand U13458 (N_13458,N_13090,N_13228);
and U13459 (N_13459,N_13236,N_13223);
or U13460 (N_13460,N_13190,N_13055);
and U13461 (N_13461,N_13043,N_13172);
or U13462 (N_13462,N_13070,N_13092);
or U13463 (N_13463,N_13116,N_13157);
nand U13464 (N_13464,N_13198,N_13004);
and U13465 (N_13465,N_13049,N_13071);
nand U13466 (N_13466,N_13130,N_13157);
or U13467 (N_13467,N_13210,N_13227);
nor U13468 (N_13468,N_13183,N_13081);
and U13469 (N_13469,N_13042,N_13198);
or U13470 (N_13470,N_13007,N_13008);
nor U13471 (N_13471,N_13157,N_13141);
and U13472 (N_13472,N_13119,N_13093);
and U13473 (N_13473,N_13068,N_13096);
nor U13474 (N_13474,N_13186,N_13004);
nand U13475 (N_13475,N_13226,N_13055);
or U13476 (N_13476,N_13236,N_13151);
or U13477 (N_13477,N_13149,N_13163);
nor U13478 (N_13478,N_13231,N_13118);
nand U13479 (N_13479,N_13157,N_13077);
or U13480 (N_13480,N_13174,N_13177);
and U13481 (N_13481,N_13060,N_13201);
or U13482 (N_13482,N_13211,N_13230);
and U13483 (N_13483,N_13176,N_13104);
nand U13484 (N_13484,N_13097,N_13154);
nand U13485 (N_13485,N_13079,N_13095);
nor U13486 (N_13486,N_13121,N_13169);
or U13487 (N_13487,N_13130,N_13115);
or U13488 (N_13488,N_13158,N_13210);
and U13489 (N_13489,N_13235,N_13160);
nor U13490 (N_13490,N_13064,N_13222);
or U13491 (N_13491,N_13205,N_13079);
or U13492 (N_13492,N_13088,N_13017);
nand U13493 (N_13493,N_13106,N_13168);
nand U13494 (N_13494,N_13118,N_13152);
or U13495 (N_13495,N_13169,N_13115);
xor U13496 (N_13496,N_13205,N_13000);
nor U13497 (N_13497,N_13128,N_13107);
nand U13498 (N_13498,N_13154,N_13068);
nand U13499 (N_13499,N_13158,N_13184);
nand U13500 (N_13500,N_13271,N_13422);
or U13501 (N_13501,N_13385,N_13416);
nand U13502 (N_13502,N_13310,N_13414);
or U13503 (N_13503,N_13328,N_13429);
and U13504 (N_13504,N_13363,N_13255);
nand U13505 (N_13505,N_13365,N_13484);
nand U13506 (N_13506,N_13267,N_13307);
nand U13507 (N_13507,N_13457,N_13330);
or U13508 (N_13508,N_13460,N_13486);
and U13509 (N_13509,N_13398,N_13437);
or U13510 (N_13510,N_13364,N_13344);
and U13511 (N_13511,N_13270,N_13407);
xor U13512 (N_13512,N_13280,N_13458);
nor U13513 (N_13513,N_13298,N_13288);
nor U13514 (N_13514,N_13435,N_13260);
or U13515 (N_13515,N_13356,N_13475);
and U13516 (N_13516,N_13321,N_13281);
or U13517 (N_13517,N_13371,N_13284);
xnor U13518 (N_13518,N_13473,N_13411);
or U13519 (N_13519,N_13444,N_13353);
nand U13520 (N_13520,N_13285,N_13468);
nor U13521 (N_13521,N_13256,N_13439);
and U13522 (N_13522,N_13495,N_13292);
nor U13523 (N_13523,N_13431,N_13463);
nor U13524 (N_13524,N_13262,N_13372);
nand U13525 (N_13525,N_13480,N_13393);
nand U13526 (N_13526,N_13254,N_13391);
or U13527 (N_13527,N_13327,N_13478);
or U13528 (N_13528,N_13423,N_13474);
xnor U13529 (N_13529,N_13388,N_13370);
and U13530 (N_13530,N_13419,N_13490);
or U13531 (N_13531,N_13358,N_13461);
nand U13532 (N_13532,N_13433,N_13263);
nor U13533 (N_13533,N_13389,N_13438);
or U13534 (N_13534,N_13311,N_13415);
xor U13535 (N_13535,N_13346,N_13387);
or U13536 (N_13536,N_13336,N_13287);
nor U13537 (N_13537,N_13317,N_13485);
xor U13538 (N_13538,N_13487,N_13343);
nor U13539 (N_13539,N_13335,N_13402);
xnor U13540 (N_13540,N_13338,N_13420);
or U13541 (N_13541,N_13290,N_13282);
or U13542 (N_13542,N_13275,N_13483);
nor U13543 (N_13543,N_13496,N_13384);
or U13544 (N_13544,N_13312,N_13305);
or U13545 (N_13545,N_13339,N_13297);
nor U13546 (N_13546,N_13395,N_13251);
and U13547 (N_13547,N_13452,N_13477);
and U13548 (N_13548,N_13257,N_13441);
or U13549 (N_13549,N_13471,N_13379);
or U13550 (N_13550,N_13482,N_13410);
or U13551 (N_13551,N_13324,N_13465);
nor U13552 (N_13552,N_13319,N_13352);
and U13553 (N_13553,N_13369,N_13318);
nor U13554 (N_13554,N_13403,N_13476);
nor U13555 (N_13555,N_13313,N_13382);
or U13556 (N_13556,N_13294,N_13467);
or U13557 (N_13557,N_13302,N_13396);
and U13558 (N_13558,N_13481,N_13424);
or U13559 (N_13559,N_13491,N_13394);
nor U13560 (N_13560,N_13445,N_13308);
nand U13561 (N_13561,N_13283,N_13268);
and U13562 (N_13562,N_13274,N_13377);
nor U13563 (N_13563,N_13265,N_13334);
nor U13564 (N_13564,N_13462,N_13325);
xor U13565 (N_13565,N_13266,N_13259);
or U13566 (N_13566,N_13426,N_13383);
nand U13567 (N_13567,N_13320,N_13314);
and U13568 (N_13568,N_13442,N_13432);
nand U13569 (N_13569,N_13303,N_13373);
nand U13570 (N_13570,N_13326,N_13451);
or U13571 (N_13571,N_13472,N_13332);
nand U13572 (N_13572,N_13340,N_13376);
nor U13573 (N_13573,N_13295,N_13447);
nor U13574 (N_13574,N_13425,N_13408);
or U13575 (N_13575,N_13299,N_13404);
nand U13576 (N_13576,N_13306,N_13291);
and U13577 (N_13577,N_13479,N_13406);
nor U13578 (N_13578,N_13455,N_13349);
nor U13579 (N_13579,N_13492,N_13417);
and U13580 (N_13580,N_13497,N_13440);
nor U13581 (N_13581,N_13378,N_13331);
or U13582 (N_13582,N_13357,N_13309);
nor U13583 (N_13583,N_13253,N_13374);
nor U13584 (N_13584,N_13296,N_13493);
nand U13585 (N_13585,N_13354,N_13392);
or U13586 (N_13586,N_13273,N_13413);
or U13587 (N_13587,N_13401,N_13386);
nand U13588 (N_13588,N_13397,N_13341);
or U13589 (N_13589,N_13470,N_13277);
nand U13590 (N_13590,N_13390,N_13367);
nand U13591 (N_13591,N_13488,N_13355);
nand U13592 (N_13592,N_13469,N_13368);
nor U13593 (N_13593,N_13449,N_13466);
xor U13594 (N_13594,N_13412,N_13252);
and U13595 (N_13595,N_13464,N_13342);
nor U13596 (N_13596,N_13286,N_13366);
nand U13597 (N_13597,N_13436,N_13278);
nand U13598 (N_13598,N_13453,N_13261);
nor U13599 (N_13599,N_13333,N_13329);
nor U13600 (N_13600,N_13375,N_13446);
nor U13601 (N_13601,N_13418,N_13360);
or U13602 (N_13602,N_13489,N_13399);
or U13603 (N_13603,N_13421,N_13293);
and U13604 (N_13604,N_13459,N_13400);
nand U13605 (N_13605,N_13405,N_13380);
and U13606 (N_13606,N_13276,N_13323);
xor U13607 (N_13607,N_13428,N_13347);
nand U13608 (N_13608,N_13362,N_13450);
or U13609 (N_13609,N_13359,N_13430);
nor U13610 (N_13610,N_13448,N_13381);
nand U13611 (N_13611,N_13264,N_13443);
nand U13612 (N_13612,N_13269,N_13494);
and U13613 (N_13613,N_13304,N_13272);
and U13614 (N_13614,N_13300,N_13456);
and U13615 (N_13615,N_13498,N_13345);
or U13616 (N_13616,N_13301,N_13322);
or U13617 (N_13617,N_13499,N_13351);
xor U13618 (N_13618,N_13316,N_13409);
nor U13619 (N_13619,N_13250,N_13361);
and U13620 (N_13620,N_13427,N_13454);
xor U13621 (N_13621,N_13258,N_13289);
nand U13622 (N_13622,N_13315,N_13337);
and U13623 (N_13623,N_13434,N_13348);
and U13624 (N_13624,N_13350,N_13279);
or U13625 (N_13625,N_13360,N_13397);
xor U13626 (N_13626,N_13334,N_13352);
nand U13627 (N_13627,N_13364,N_13395);
nand U13628 (N_13628,N_13392,N_13286);
nand U13629 (N_13629,N_13254,N_13455);
nor U13630 (N_13630,N_13496,N_13322);
and U13631 (N_13631,N_13494,N_13387);
nor U13632 (N_13632,N_13292,N_13304);
and U13633 (N_13633,N_13292,N_13256);
or U13634 (N_13634,N_13359,N_13333);
and U13635 (N_13635,N_13357,N_13297);
nor U13636 (N_13636,N_13419,N_13497);
nand U13637 (N_13637,N_13457,N_13490);
and U13638 (N_13638,N_13290,N_13457);
xor U13639 (N_13639,N_13286,N_13499);
nor U13640 (N_13640,N_13415,N_13357);
and U13641 (N_13641,N_13313,N_13302);
nor U13642 (N_13642,N_13257,N_13404);
nand U13643 (N_13643,N_13345,N_13373);
nor U13644 (N_13644,N_13322,N_13308);
or U13645 (N_13645,N_13325,N_13452);
and U13646 (N_13646,N_13288,N_13384);
or U13647 (N_13647,N_13327,N_13286);
xor U13648 (N_13648,N_13252,N_13394);
and U13649 (N_13649,N_13406,N_13274);
nor U13650 (N_13650,N_13401,N_13409);
nand U13651 (N_13651,N_13474,N_13266);
nor U13652 (N_13652,N_13290,N_13461);
nor U13653 (N_13653,N_13291,N_13308);
xor U13654 (N_13654,N_13470,N_13296);
nand U13655 (N_13655,N_13285,N_13337);
and U13656 (N_13656,N_13327,N_13295);
xnor U13657 (N_13657,N_13457,N_13446);
or U13658 (N_13658,N_13268,N_13322);
nor U13659 (N_13659,N_13353,N_13469);
nand U13660 (N_13660,N_13407,N_13306);
xor U13661 (N_13661,N_13348,N_13415);
nor U13662 (N_13662,N_13319,N_13431);
nand U13663 (N_13663,N_13415,N_13342);
and U13664 (N_13664,N_13367,N_13310);
and U13665 (N_13665,N_13252,N_13395);
xor U13666 (N_13666,N_13430,N_13315);
and U13667 (N_13667,N_13253,N_13301);
nand U13668 (N_13668,N_13455,N_13379);
and U13669 (N_13669,N_13300,N_13496);
or U13670 (N_13670,N_13365,N_13260);
or U13671 (N_13671,N_13266,N_13346);
xor U13672 (N_13672,N_13449,N_13457);
and U13673 (N_13673,N_13479,N_13405);
or U13674 (N_13674,N_13319,N_13277);
or U13675 (N_13675,N_13477,N_13291);
nor U13676 (N_13676,N_13369,N_13348);
xnor U13677 (N_13677,N_13441,N_13396);
nand U13678 (N_13678,N_13344,N_13423);
or U13679 (N_13679,N_13371,N_13251);
nand U13680 (N_13680,N_13338,N_13310);
nand U13681 (N_13681,N_13347,N_13340);
and U13682 (N_13682,N_13304,N_13326);
nor U13683 (N_13683,N_13439,N_13379);
or U13684 (N_13684,N_13281,N_13441);
and U13685 (N_13685,N_13492,N_13317);
nor U13686 (N_13686,N_13319,N_13490);
nor U13687 (N_13687,N_13304,N_13368);
or U13688 (N_13688,N_13412,N_13311);
and U13689 (N_13689,N_13275,N_13407);
or U13690 (N_13690,N_13297,N_13401);
and U13691 (N_13691,N_13374,N_13316);
and U13692 (N_13692,N_13459,N_13475);
nand U13693 (N_13693,N_13466,N_13288);
nand U13694 (N_13694,N_13422,N_13266);
xnor U13695 (N_13695,N_13281,N_13301);
nand U13696 (N_13696,N_13488,N_13481);
nor U13697 (N_13697,N_13368,N_13493);
and U13698 (N_13698,N_13488,N_13367);
nand U13699 (N_13699,N_13372,N_13399);
or U13700 (N_13700,N_13267,N_13296);
and U13701 (N_13701,N_13492,N_13292);
nand U13702 (N_13702,N_13423,N_13309);
or U13703 (N_13703,N_13437,N_13275);
or U13704 (N_13704,N_13400,N_13346);
nor U13705 (N_13705,N_13301,N_13429);
or U13706 (N_13706,N_13369,N_13306);
xor U13707 (N_13707,N_13369,N_13339);
nand U13708 (N_13708,N_13303,N_13367);
or U13709 (N_13709,N_13451,N_13328);
nor U13710 (N_13710,N_13269,N_13385);
and U13711 (N_13711,N_13284,N_13299);
and U13712 (N_13712,N_13426,N_13302);
nor U13713 (N_13713,N_13381,N_13401);
nor U13714 (N_13714,N_13367,N_13449);
nor U13715 (N_13715,N_13451,N_13426);
nand U13716 (N_13716,N_13259,N_13485);
and U13717 (N_13717,N_13368,N_13353);
or U13718 (N_13718,N_13478,N_13472);
and U13719 (N_13719,N_13326,N_13413);
nor U13720 (N_13720,N_13285,N_13336);
nor U13721 (N_13721,N_13450,N_13277);
and U13722 (N_13722,N_13479,N_13421);
and U13723 (N_13723,N_13450,N_13283);
nand U13724 (N_13724,N_13447,N_13495);
nand U13725 (N_13725,N_13495,N_13435);
nor U13726 (N_13726,N_13256,N_13455);
and U13727 (N_13727,N_13396,N_13456);
nand U13728 (N_13728,N_13499,N_13426);
and U13729 (N_13729,N_13383,N_13375);
nand U13730 (N_13730,N_13453,N_13465);
or U13731 (N_13731,N_13316,N_13498);
and U13732 (N_13732,N_13449,N_13355);
nor U13733 (N_13733,N_13336,N_13303);
and U13734 (N_13734,N_13294,N_13464);
nor U13735 (N_13735,N_13345,N_13477);
or U13736 (N_13736,N_13334,N_13403);
or U13737 (N_13737,N_13442,N_13389);
and U13738 (N_13738,N_13380,N_13450);
and U13739 (N_13739,N_13272,N_13340);
nand U13740 (N_13740,N_13273,N_13284);
and U13741 (N_13741,N_13265,N_13373);
xnor U13742 (N_13742,N_13479,N_13392);
nor U13743 (N_13743,N_13428,N_13261);
nor U13744 (N_13744,N_13442,N_13434);
nor U13745 (N_13745,N_13340,N_13412);
or U13746 (N_13746,N_13250,N_13313);
nand U13747 (N_13747,N_13403,N_13288);
nor U13748 (N_13748,N_13412,N_13436);
and U13749 (N_13749,N_13319,N_13492);
nor U13750 (N_13750,N_13729,N_13601);
and U13751 (N_13751,N_13518,N_13566);
nor U13752 (N_13752,N_13620,N_13623);
and U13753 (N_13753,N_13569,N_13737);
or U13754 (N_13754,N_13543,N_13742);
and U13755 (N_13755,N_13593,N_13663);
xnor U13756 (N_13756,N_13656,N_13688);
nand U13757 (N_13757,N_13727,N_13536);
nor U13758 (N_13758,N_13733,N_13607);
and U13759 (N_13759,N_13724,N_13707);
nand U13760 (N_13760,N_13686,N_13626);
xnor U13761 (N_13761,N_13554,N_13500);
or U13762 (N_13762,N_13628,N_13710);
and U13763 (N_13763,N_13571,N_13602);
and U13764 (N_13764,N_13680,N_13615);
or U13765 (N_13765,N_13638,N_13735);
nor U13766 (N_13766,N_13552,N_13563);
and U13767 (N_13767,N_13624,N_13722);
nor U13768 (N_13768,N_13644,N_13517);
xnor U13769 (N_13769,N_13502,N_13698);
nand U13770 (N_13770,N_13587,N_13622);
nor U13771 (N_13771,N_13661,N_13514);
nand U13772 (N_13772,N_13654,N_13702);
and U13773 (N_13773,N_13515,N_13549);
nand U13774 (N_13774,N_13540,N_13556);
nand U13775 (N_13775,N_13504,N_13558);
xnor U13776 (N_13776,N_13512,N_13676);
and U13777 (N_13777,N_13511,N_13719);
or U13778 (N_13778,N_13604,N_13618);
or U13779 (N_13779,N_13651,N_13667);
nand U13780 (N_13780,N_13613,N_13709);
and U13781 (N_13781,N_13521,N_13508);
and U13782 (N_13782,N_13541,N_13665);
or U13783 (N_13783,N_13526,N_13546);
nor U13784 (N_13784,N_13542,N_13568);
xnor U13785 (N_13785,N_13599,N_13744);
and U13786 (N_13786,N_13561,N_13690);
nor U13787 (N_13787,N_13695,N_13575);
nor U13788 (N_13788,N_13528,N_13678);
nor U13789 (N_13789,N_13625,N_13582);
nand U13790 (N_13790,N_13637,N_13712);
nand U13791 (N_13791,N_13642,N_13588);
nand U13792 (N_13792,N_13633,N_13681);
or U13793 (N_13793,N_13657,N_13714);
and U13794 (N_13794,N_13529,N_13736);
nand U13795 (N_13795,N_13648,N_13720);
nand U13796 (N_13796,N_13603,N_13718);
nor U13797 (N_13797,N_13745,N_13592);
nand U13798 (N_13798,N_13619,N_13595);
or U13799 (N_13799,N_13574,N_13721);
xor U13800 (N_13800,N_13564,N_13723);
or U13801 (N_13801,N_13562,N_13666);
or U13802 (N_13802,N_13610,N_13594);
xnor U13803 (N_13803,N_13725,N_13635);
and U13804 (N_13804,N_13658,N_13509);
nor U13805 (N_13805,N_13598,N_13522);
or U13806 (N_13806,N_13584,N_13649);
nand U13807 (N_13807,N_13576,N_13501);
nand U13808 (N_13808,N_13664,N_13660);
nor U13809 (N_13809,N_13747,N_13559);
and U13810 (N_13810,N_13506,N_13730);
nand U13811 (N_13811,N_13748,N_13672);
nor U13812 (N_13812,N_13694,N_13550);
nand U13813 (N_13813,N_13567,N_13643);
or U13814 (N_13814,N_13674,N_13706);
or U13815 (N_13815,N_13617,N_13697);
or U13816 (N_13816,N_13662,N_13641);
nand U13817 (N_13817,N_13537,N_13749);
or U13818 (N_13818,N_13734,N_13606);
nand U13819 (N_13819,N_13557,N_13590);
nor U13820 (N_13820,N_13668,N_13539);
nand U13821 (N_13821,N_13596,N_13591);
nand U13822 (N_13822,N_13731,N_13728);
nor U13823 (N_13823,N_13673,N_13685);
and U13824 (N_13824,N_13560,N_13503);
nand U13825 (N_13825,N_13530,N_13645);
and U13826 (N_13826,N_13715,N_13655);
and U13827 (N_13827,N_13650,N_13646);
and U13828 (N_13828,N_13732,N_13614);
or U13829 (N_13829,N_13671,N_13533);
nor U13830 (N_13830,N_13589,N_13516);
or U13831 (N_13831,N_13684,N_13581);
or U13832 (N_13832,N_13682,N_13565);
or U13833 (N_13833,N_13519,N_13621);
or U13834 (N_13834,N_13585,N_13640);
and U13835 (N_13835,N_13700,N_13687);
and U13836 (N_13836,N_13545,N_13534);
or U13837 (N_13837,N_13743,N_13693);
nand U13838 (N_13838,N_13551,N_13739);
and U13839 (N_13839,N_13675,N_13669);
xor U13840 (N_13840,N_13634,N_13741);
and U13841 (N_13841,N_13583,N_13555);
or U13842 (N_13842,N_13580,N_13647);
nor U13843 (N_13843,N_13713,N_13716);
xnor U13844 (N_13844,N_13746,N_13573);
nor U13845 (N_13845,N_13578,N_13726);
xnor U13846 (N_13846,N_13600,N_13548);
and U13847 (N_13847,N_13505,N_13740);
and U13848 (N_13848,N_13670,N_13523);
and U13849 (N_13849,N_13738,N_13544);
and U13850 (N_13850,N_13609,N_13524);
nor U13851 (N_13851,N_13627,N_13535);
nor U13852 (N_13852,N_13705,N_13696);
nand U13853 (N_13853,N_13683,N_13639);
nor U13854 (N_13854,N_13691,N_13570);
and U13855 (N_13855,N_13527,N_13701);
or U13856 (N_13856,N_13636,N_13708);
and U13857 (N_13857,N_13612,N_13630);
or U13858 (N_13858,N_13611,N_13572);
xor U13859 (N_13859,N_13520,N_13513);
xor U13860 (N_13860,N_13659,N_13692);
nor U13861 (N_13861,N_13531,N_13677);
xor U13862 (N_13862,N_13553,N_13679);
nand U13863 (N_13863,N_13532,N_13652);
or U13864 (N_13864,N_13653,N_13579);
or U13865 (N_13865,N_13608,N_13538);
and U13866 (N_13866,N_13507,N_13629);
nor U13867 (N_13867,N_13689,N_13704);
or U13868 (N_13868,N_13597,N_13605);
and U13869 (N_13869,N_13586,N_13577);
or U13870 (N_13870,N_13510,N_13699);
or U13871 (N_13871,N_13616,N_13547);
and U13872 (N_13872,N_13525,N_13717);
nor U13873 (N_13873,N_13632,N_13711);
nand U13874 (N_13874,N_13631,N_13703);
nor U13875 (N_13875,N_13563,N_13691);
nor U13876 (N_13876,N_13703,N_13524);
or U13877 (N_13877,N_13526,N_13514);
xnor U13878 (N_13878,N_13666,N_13622);
nor U13879 (N_13879,N_13627,N_13547);
or U13880 (N_13880,N_13685,N_13633);
nor U13881 (N_13881,N_13561,N_13556);
nand U13882 (N_13882,N_13515,N_13698);
and U13883 (N_13883,N_13682,N_13563);
or U13884 (N_13884,N_13713,N_13651);
or U13885 (N_13885,N_13691,N_13729);
xnor U13886 (N_13886,N_13622,N_13584);
and U13887 (N_13887,N_13633,N_13507);
nand U13888 (N_13888,N_13587,N_13639);
nand U13889 (N_13889,N_13515,N_13574);
and U13890 (N_13890,N_13501,N_13599);
or U13891 (N_13891,N_13650,N_13645);
nand U13892 (N_13892,N_13546,N_13709);
and U13893 (N_13893,N_13561,N_13584);
or U13894 (N_13894,N_13539,N_13720);
nand U13895 (N_13895,N_13531,N_13540);
nand U13896 (N_13896,N_13602,N_13565);
and U13897 (N_13897,N_13616,N_13664);
nor U13898 (N_13898,N_13557,N_13624);
nand U13899 (N_13899,N_13713,N_13637);
nand U13900 (N_13900,N_13615,N_13527);
and U13901 (N_13901,N_13592,N_13558);
nand U13902 (N_13902,N_13530,N_13566);
and U13903 (N_13903,N_13573,N_13501);
or U13904 (N_13904,N_13516,N_13500);
and U13905 (N_13905,N_13692,N_13611);
nand U13906 (N_13906,N_13505,N_13515);
and U13907 (N_13907,N_13618,N_13565);
nand U13908 (N_13908,N_13730,N_13646);
or U13909 (N_13909,N_13556,N_13580);
nand U13910 (N_13910,N_13596,N_13659);
nand U13911 (N_13911,N_13559,N_13555);
or U13912 (N_13912,N_13720,N_13666);
or U13913 (N_13913,N_13578,N_13556);
nor U13914 (N_13914,N_13681,N_13701);
nor U13915 (N_13915,N_13727,N_13648);
and U13916 (N_13916,N_13640,N_13503);
or U13917 (N_13917,N_13508,N_13721);
or U13918 (N_13918,N_13506,N_13546);
nor U13919 (N_13919,N_13747,N_13700);
or U13920 (N_13920,N_13575,N_13744);
nor U13921 (N_13921,N_13649,N_13521);
nand U13922 (N_13922,N_13559,N_13637);
or U13923 (N_13923,N_13504,N_13577);
xor U13924 (N_13924,N_13633,N_13735);
or U13925 (N_13925,N_13595,N_13509);
and U13926 (N_13926,N_13602,N_13745);
nand U13927 (N_13927,N_13641,N_13744);
nand U13928 (N_13928,N_13709,N_13720);
nand U13929 (N_13929,N_13506,N_13690);
and U13930 (N_13930,N_13568,N_13603);
nand U13931 (N_13931,N_13522,N_13511);
nand U13932 (N_13932,N_13639,N_13660);
xor U13933 (N_13933,N_13620,N_13671);
nand U13934 (N_13934,N_13593,N_13509);
nor U13935 (N_13935,N_13558,N_13619);
or U13936 (N_13936,N_13692,N_13566);
or U13937 (N_13937,N_13665,N_13654);
and U13938 (N_13938,N_13570,N_13575);
nor U13939 (N_13939,N_13541,N_13668);
and U13940 (N_13940,N_13635,N_13717);
or U13941 (N_13941,N_13566,N_13543);
nand U13942 (N_13942,N_13642,N_13537);
nor U13943 (N_13943,N_13501,N_13697);
or U13944 (N_13944,N_13700,N_13621);
nor U13945 (N_13945,N_13592,N_13604);
nand U13946 (N_13946,N_13657,N_13504);
and U13947 (N_13947,N_13508,N_13685);
nand U13948 (N_13948,N_13725,N_13716);
nand U13949 (N_13949,N_13634,N_13563);
and U13950 (N_13950,N_13722,N_13550);
or U13951 (N_13951,N_13571,N_13730);
and U13952 (N_13952,N_13703,N_13509);
and U13953 (N_13953,N_13645,N_13622);
nand U13954 (N_13954,N_13674,N_13682);
and U13955 (N_13955,N_13592,N_13665);
nand U13956 (N_13956,N_13548,N_13564);
nand U13957 (N_13957,N_13734,N_13693);
nand U13958 (N_13958,N_13592,N_13634);
nand U13959 (N_13959,N_13573,N_13684);
xor U13960 (N_13960,N_13635,N_13648);
and U13961 (N_13961,N_13559,N_13634);
and U13962 (N_13962,N_13540,N_13647);
or U13963 (N_13963,N_13581,N_13656);
and U13964 (N_13964,N_13547,N_13558);
nor U13965 (N_13965,N_13542,N_13684);
and U13966 (N_13966,N_13567,N_13629);
nor U13967 (N_13967,N_13715,N_13706);
nand U13968 (N_13968,N_13696,N_13630);
xor U13969 (N_13969,N_13605,N_13642);
and U13970 (N_13970,N_13541,N_13717);
and U13971 (N_13971,N_13595,N_13522);
nor U13972 (N_13972,N_13526,N_13507);
or U13973 (N_13973,N_13547,N_13651);
nand U13974 (N_13974,N_13700,N_13516);
nor U13975 (N_13975,N_13609,N_13520);
nand U13976 (N_13976,N_13575,N_13673);
or U13977 (N_13977,N_13524,N_13679);
nor U13978 (N_13978,N_13546,N_13683);
nand U13979 (N_13979,N_13589,N_13635);
nor U13980 (N_13980,N_13689,N_13721);
xor U13981 (N_13981,N_13535,N_13734);
xnor U13982 (N_13982,N_13715,N_13620);
nand U13983 (N_13983,N_13680,N_13593);
nand U13984 (N_13984,N_13579,N_13638);
or U13985 (N_13985,N_13530,N_13586);
or U13986 (N_13986,N_13671,N_13636);
or U13987 (N_13987,N_13701,N_13727);
nor U13988 (N_13988,N_13742,N_13598);
or U13989 (N_13989,N_13503,N_13624);
nor U13990 (N_13990,N_13626,N_13567);
nand U13991 (N_13991,N_13642,N_13687);
or U13992 (N_13992,N_13648,N_13738);
nand U13993 (N_13993,N_13693,N_13673);
nor U13994 (N_13994,N_13645,N_13603);
or U13995 (N_13995,N_13565,N_13683);
nand U13996 (N_13996,N_13548,N_13711);
nor U13997 (N_13997,N_13672,N_13624);
and U13998 (N_13998,N_13675,N_13533);
nand U13999 (N_13999,N_13708,N_13553);
nor U14000 (N_14000,N_13921,N_13829);
nor U14001 (N_14001,N_13761,N_13997);
nor U14002 (N_14002,N_13898,N_13854);
xor U14003 (N_14003,N_13964,N_13792);
and U14004 (N_14004,N_13920,N_13950);
or U14005 (N_14005,N_13817,N_13773);
nand U14006 (N_14006,N_13840,N_13808);
or U14007 (N_14007,N_13990,N_13986);
and U14008 (N_14008,N_13873,N_13752);
or U14009 (N_14009,N_13899,N_13767);
nor U14010 (N_14010,N_13935,N_13960);
nand U14011 (N_14011,N_13769,N_13895);
nor U14012 (N_14012,N_13778,N_13903);
nand U14013 (N_14013,N_13813,N_13844);
nand U14014 (N_14014,N_13883,N_13956);
or U14015 (N_14015,N_13993,N_13849);
or U14016 (N_14016,N_13926,N_13803);
nor U14017 (N_14017,N_13830,N_13762);
or U14018 (N_14018,N_13901,N_13868);
and U14019 (N_14019,N_13824,N_13969);
nor U14020 (N_14020,N_13764,N_13765);
or U14021 (N_14021,N_13911,N_13794);
and U14022 (N_14022,N_13980,N_13947);
and U14023 (N_14023,N_13820,N_13800);
and U14024 (N_14024,N_13798,N_13835);
nor U14025 (N_14025,N_13755,N_13793);
or U14026 (N_14026,N_13856,N_13771);
or U14027 (N_14027,N_13788,N_13968);
and U14028 (N_14028,N_13836,N_13825);
and U14029 (N_14029,N_13860,N_13970);
xnor U14030 (N_14030,N_13959,N_13878);
nor U14031 (N_14031,N_13858,N_13861);
and U14032 (N_14032,N_13904,N_13996);
nor U14033 (N_14033,N_13910,N_13987);
or U14034 (N_14034,N_13823,N_13949);
xnor U14035 (N_14035,N_13859,N_13984);
or U14036 (N_14036,N_13971,N_13790);
and U14037 (N_14037,N_13916,N_13811);
nand U14038 (N_14038,N_13795,N_13754);
nor U14039 (N_14039,N_13757,N_13966);
and U14040 (N_14040,N_13967,N_13924);
nand U14041 (N_14041,N_13892,N_13822);
or U14042 (N_14042,N_13938,N_13838);
and U14043 (N_14043,N_13994,N_13982);
or U14044 (N_14044,N_13880,N_13891);
or U14045 (N_14045,N_13770,N_13818);
nor U14046 (N_14046,N_13827,N_13962);
nor U14047 (N_14047,N_13974,N_13922);
and U14048 (N_14048,N_13846,N_13884);
nand U14049 (N_14049,N_13936,N_13985);
nand U14050 (N_14050,N_13907,N_13785);
or U14051 (N_14051,N_13981,N_13954);
nand U14052 (N_14052,N_13851,N_13925);
nor U14053 (N_14053,N_13976,N_13796);
nor U14054 (N_14054,N_13995,N_13882);
or U14055 (N_14055,N_13957,N_13945);
or U14056 (N_14056,N_13992,N_13801);
and U14057 (N_14057,N_13784,N_13821);
and U14058 (N_14058,N_13831,N_13782);
and U14059 (N_14059,N_13937,N_13870);
or U14060 (N_14060,N_13912,N_13975);
nor U14061 (N_14061,N_13948,N_13963);
or U14062 (N_14062,N_13760,N_13841);
xnor U14063 (N_14063,N_13802,N_13988);
or U14064 (N_14064,N_13750,N_13864);
and U14065 (N_14065,N_13852,N_13958);
nor U14066 (N_14066,N_13890,N_13906);
xor U14067 (N_14067,N_13874,N_13972);
xor U14068 (N_14068,N_13776,N_13917);
and U14069 (N_14069,N_13815,N_13872);
or U14070 (N_14070,N_13863,N_13914);
or U14071 (N_14071,N_13928,N_13900);
nand U14072 (N_14072,N_13918,N_13845);
nand U14073 (N_14073,N_13833,N_13961);
nand U14074 (N_14074,N_13826,N_13983);
and U14075 (N_14075,N_13828,N_13832);
or U14076 (N_14076,N_13929,N_13881);
and U14077 (N_14077,N_13867,N_13989);
or U14078 (N_14078,N_13991,N_13923);
and U14079 (N_14079,N_13893,N_13941);
or U14080 (N_14080,N_13809,N_13876);
nand U14081 (N_14081,N_13889,N_13804);
xor U14082 (N_14082,N_13886,N_13812);
xor U14083 (N_14083,N_13953,N_13763);
nor U14084 (N_14084,N_13805,N_13857);
nand U14085 (N_14085,N_13894,N_13806);
or U14086 (N_14086,N_13853,N_13816);
nand U14087 (N_14087,N_13998,N_13839);
nor U14088 (N_14088,N_13939,N_13759);
xnor U14089 (N_14089,N_13869,N_13887);
nand U14090 (N_14090,N_13753,N_13834);
nand U14091 (N_14091,N_13837,N_13942);
nor U14092 (N_14092,N_13946,N_13940);
or U14093 (N_14093,N_13774,N_13965);
or U14094 (N_14094,N_13933,N_13797);
and U14095 (N_14095,N_13930,N_13842);
or U14096 (N_14096,N_13766,N_13877);
nand U14097 (N_14097,N_13850,N_13919);
and U14098 (N_14098,N_13955,N_13848);
and U14099 (N_14099,N_13973,N_13814);
and U14100 (N_14100,N_13847,N_13908);
nor U14101 (N_14101,N_13934,N_13913);
and U14102 (N_14102,N_13978,N_13943);
xnor U14103 (N_14103,N_13927,N_13783);
nand U14104 (N_14104,N_13779,N_13751);
xor U14105 (N_14105,N_13897,N_13768);
nor U14106 (N_14106,N_13979,N_13871);
nand U14107 (N_14107,N_13758,N_13931);
and U14108 (N_14108,N_13875,N_13885);
nand U14109 (N_14109,N_13977,N_13944);
or U14110 (N_14110,N_13896,N_13952);
and U14111 (N_14111,N_13866,N_13843);
and U14112 (N_14112,N_13999,N_13879);
and U14113 (N_14113,N_13807,N_13819);
nor U14114 (N_14114,N_13780,N_13855);
and U14115 (N_14115,N_13787,N_13932);
or U14116 (N_14116,N_13902,N_13786);
nor U14117 (N_14117,N_13915,N_13789);
and U14118 (N_14118,N_13865,N_13756);
and U14119 (N_14119,N_13772,N_13810);
and U14120 (N_14120,N_13799,N_13781);
nand U14121 (N_14121,N_13951,N_13888);
or U14122 (N_14122,N_13791,N_13775);
or U14123 (N_14123,N_13862,N_13905);
or U14124 (N_14124,N_13909,N_13777);
nand U14125 (N_14125,N_13910,N_13839);
or U14126 (N_14126,N_13994,N_13990);
and U14127 (N_14127,N_13774,N_13828);
or U14128 (N_14128,N_13804,N_13838);
nand U14129 (N_14129,N_13914,N_13797);
and U14130 (N_14130,N_13813,N_13882);
or U14131 (N_14131,N_13787,N_13829);
nand U14132 (N_14132,N_13840,N_13857);
nand U14133 (N_14133,N_13990,N_13947);
or U14134 (N_14134,N_13792,N_13813);
and U14135 (N_14135,N_13962,N_13825);
and U14136 (N_14136,N_13825,N_13916);
xnor U14137 (N_14137,N_13783,N_13768);
or U14138 (N_14138,N_13935,N_13817);
or U14139 (N_14139,N_13933,N_13842);
and U14140 (N_14140,N_13986,N_13808);
and U14141 (N_14141,N_13896,N_13994);
xnor U14142 (N_14142,N_13904,N_13929);
nor U14143 (N_14143,N_13836,N_13858);
and U14144 (N_14144,N_13885,N_13947);
and U14145 (N_14145,N_13951,N_13879);
xnor U14146 (N_14146,N_13999,N_13895);
or U14147 (N_14147,N_13885,N_13840);
nand U14148 (N_14148,N_13792,N_13775);
and U14149 (N_14149,N_13815,N_13983);
or U14150 (N_14150,N_13894,N_13776);
and U14151 (N_14151,N_13908,N_13821);
nand U14152 (N_14152,N_13784,N_13840);
and U14153 (N_14153,N_13895,N_13966);
nand U14154 (N_14154,N_13824,N_13944);
and U14155 (N_14155,N_13890,N_13815);
nand U14156 (N_14156,N_13772,N_13940);
and U14157 (N_14157,N_13921,N_13887);
and U14158 (N_14158,N_13780,N_13880);
nor U14159 (N_14159,N_13966,N_13897);
and U14160 (N_14160,N_13751,N_13936);
nand U14161 (N_14161,N_13980,N_13836);
and U14162 (N_14162,N_13845,N_13783);
and U14163 (N_14163,N_13812,N_13827);
and U14164 (N_14164,N_13950,N_13848);
nor U14165 (N_14165,N_13978,N_13969);
nor U14166 (N_14166,N_13917,N_13857);
nor U14167 (N_14167,N_13773,N_13967);
and U14168 (N_14168,N_13769,N_13945);
nand U14169 (N_14169,N_13798,N_13771);
or U14170 (N_14170,N_13924,N_13822);
xnor U14171 (N_14171,N_13803,N_13832);
nor U14172 (N_14172,N_13975,N_13955);
xnor U14173 (N_14173,N_13808,N_13906);
nor U14174 (N_14174,N_13867,N_13801);
and U14175 (N_14175,N_13955,N_13874);
nor U14176 (N_14176,N_13752,N_13907);
nand U14177 (N_14177,N_13834,N_13952);
nand U14178 (N_14178,N_13753,N_13883);
nand U14179 (N_14179,N_13842,N_13887);
and U14180 (N_14180,N_13761,N_13963);
nor U14181 (N_14181,N_13753,N_13826);
or U14182 (N_14182,N_13879,N_13777);
nand U14183 (N_14183,N_13991,N_13857);
or U14184 (N_14184,N_13873,N_13928);
and U14185 (N_14185,N_13985,N_13805);
nor U14186 (N_14186,N_13865,N_13988);
or U14187 (N_14187,N_13843,N_13857);
xor U14188 (N_14188,N_13783,N_13911);
nor U14189 (N_14189,N_13992,N_13921);
and U14190 (N_14190,N_13860,N_13841);
nand U14191 (N_14191,N_13776,N_13759);
nor U14192 (N_14192,N_13773,N_13899);
or U14193 (N_14193,N_13881,N_13815);
nor U14194 (N_14194,N_13990,N_13946);
or U14195 (N_14195,N_13928,N_13790);
nand U14196 (N_14196,N_13856,N_13832);
and U14197 (N_14197,N_13797,N_13830);
xor U14198 (N_14198,N_13967,N_13870);
nand U14199 (N_14199,N_13997,N_13874);
nand U14200 (N_14200,N_13866,N_13780);
nand U14201 (N_14201,N_13991,N_13970);
xor U14202 (N_14202,N_13930,N_13973);
and U14203 (N_14203,N_13789,N_13982);
nor U14204 (N_14204,N_13802,N_13831);
nor U14205 (N_14205,N_13791,N_13997);
nor U14206 (N_14206,N_13883,N_13815);
nor U14207 (N_14207,N_13852,N_13933);
or U14208 (N_14208,N_13753,N_13758);
xnor U14209 (N_14209,N_13878,N_13951);
nand U14210 (N_14210,N_13823,N_13974);
nor U14211 (N_14211,N_13807,N_13919);
nor U14212 (N_14212,N_13895,N_13971);
nand U14213 (N_14213,N_13905,N_13793);
xnor U14214 (N_14214,N_13799,N_13849);
nand U14215 (N_14215,N_13863,N_13927);
nand U14216 (N_14216,N_13811,N_13836);
nand U14217 (N_14217,N_13938,N_13994);
xnor U14218 (N_14218,N_13781,N_13955);
and U14219 (N_14219,N_13756,N_13786);
xnor U14220 (N_14220,N_13846,N_13985);
and U14221 (N_14221,N_13933,N_13878);
nor U14222 (N_14222,N_13914,N_13803);
nor U14223 (N_14223,N_13956,N_13763);
or U14224 (N_14224,N_13779,N_13984);
xnor U14225 (N_14225,N_13876,N_13784);
nor U14226 (N_14226,N_13863,N_13753);
nand U14227 (N_14227,N_13907,N_13920);
xnor U14228 (N_14228,N_13751,N_13871);
and U14229 (N_14229,N_13870,N_13894);
nand U14230 (N_14230,N_13790,N_13985);
nor U14231 (N_14231,N_13974,N_13964);
nand U14232 (N_14232,N_13898,N_13866);
and U14233 (N_14233,N_13938,N_13850);
nor U14234 (N_14234,N_13961,N_13963);
xnor U14235 (N_14235,N_13919,N_13958);
and U14236 (N_14236,N_13996,N_13814);
nand U14237 (N_14237,N_13980,N_13868);
nor U14238 (N_14238,N_13765,N_13879);
nor U14239 (N_14239,N_13828,N_13758);
or U14240 (N_14240,N_13851,N_13912);
nand U14241 (N_14241,N_13922,N_13775);
or U14242 (N_14242,N_13764,N_13843);
nand U14243 (N_14243,N_13781,N_13790);
nor U14244 (N_14244,N_13819,N_13767);
nand U14245 (N_14245,N_13756,N_13787);
nor U14246 (N_14246,N_13958,N_13782);
nor U14247 (N_14247,N_13945,N_13802);
nand U14248 (N_14248,N_13960,N_13765);
nand U14249 (N_14249,N_13891,N_13866);
or U14250 (N_14250,N_14136,N_14060);
xor U14251 (N_14251,N_14050,N_14088);
nor U14252 (N_14252,N_14047,N_14230);
and U14253 (N_14253,N_14203,N_14196);
nand U14254 (N_14254,N_14000,N_14124);
nand U14255 (N_14255,N_14023,N_14046);
nor U14256 (N_14256,N_14036,N_14140);
and U14257 (N_14257,N_14211,N_14226);
nor U14258 (N_14258,N_14242,N_14214);
and U14259 (N_14259,N_14123,N_14195);
nor U14260 (N_14260,N_14122,N_14161);
nand U14261 (N_14261,N_14021,N_14058);
or U14262 (N_14262,N_14182,N_14162);
nor U14263 (N_14263,N_14144,N_14110);
or U14264 (N_14264,N_14139,N_14163);
nor U14265 (N_14265,N_14133,N_14084);
xnor U14266 (N_14266,N_14237,N_14033);
nor U14267 (N_14267,N_14020,N_14238);
nor U14268 (N_14268,N_14146,N_14044);
nor U14269 (N_14269,N_14151,N_14028);
nand U14270 (N_14270,N_14248,N_14216);
and U14271 (N_14271,N_14164,N_14007);
nand U14272 (N_14272,N_14108,N_14170);
and U14273 (N_14273,N_14006,N_14165);
or U14274 (N_14274,N_14131,N_14159);
nor U14275 (N_14275,N_14045,N_14002);
nor U14276 (N_14276,N_14068,N_14116);
nand U14277 (N_14277,N_14208,N_14075);
and U14278 (N_14278,N_14077,N_14143);
xnor U14279 (N_14279,N_14115,N_14041);
nand U14280 (N_14280,N_14065,N_14086);
or U14281 (N_14281,N_14079,N_14071);
nand U14282 (N_14282,N_14245,N_14022);
nand U14283 (N_14283,N_14099,N_14193);
nand U14284 (N_14284,N_14149,N_14184);
and U14285 (N_14285,N_14119,N_14016);
nand U14286 (N_14286,N_14180,N_14246);
nor U14287 (N_14287,N_14055,N_14073);
or U14288 (N_14288,N_14176,N_14094);
or U14289 (N_14289,N_14096,N_14104);
nor U14290 (N_14290,N_14090,N_14109);
nor U14291 (N_14291,N_14040,N_14014);
and U14292 (N_14292,N_14153,N_14039);
nor U14293 (N_14293,N_14142,N_14015);
or U14294 (N_14294,N_14168,N_14220);
or U14295 (N_14295,N_14158,N_14137);
and U14296 (N_14296,N_14236,N_14064);
nor U14297 (N_14297,N_14054,N_14197);
nor U14298 (N_14298,N_14082,N_14191);
and U14299 (N_14299,N_14222,N_14138);
or U14300 (N_14300,N_14097,N_14154);
or U14301 (N_14301,N_14053,N_14025);
and U14302 (N_14302,N_14061,N_14009);
or U14303 (N_14303,N_14240,N_14056);
and U14304 (N_14304,N_14187,N_14098);
nand U14305 (N_14305,N_14037,N_14171);
and U14306 (N_14306,N_14003,N_14189);
nor U14307 (N_14307,N_14147,N_14231);
and U14308 (N_14308,N_14188,N_14031);
nand U14309 (N_14309,N_14114,N_14118);
and U14310 (N_14310,N_14186,N_14190);
nand U14311 (N_14311,N_14232,N_14092);
xor U14312 (N_14312,N_14224,N_14004);
and U14313 (N_14313,N_14239,N_14194);
and U14314 (N_14314,N_14048,N_14113);
and U14315 (N_14315,N_14013,N_14057);
nor U14316 (N_14316,N_14038,N_14201);
nor U14317 (N_14317,N_14218,N_14229);
or U14318 (N_14318,N_14233,N_14063);
or U14319 (N_14319,N_14095,N_14204);
nor U14320 (N_14320,N_14102,N_14129);
nand U14321 (N_14321,N_14029,N_14235);
and U14322 (N_14322,N_14083,N_14241);
or U14323 (N_14323,N_14217,N_14173);
or U14324 (N_14324,N_14125,N_14127);
nor U14325 (N_14325,N_14166,N_14062);
nand U14326 (N_14326,N_14132,N_14209);
nor U14327 (N_14327,N_14052,N_14049);
and U14328 (N_14328,N_14042,N_14121);
nand U14329 (N_14329,N_14223,N_14177);
nand U14330 (N_14330,N_14005,N_14091);
and U14331 (N_14331,N_14010,N_14072);
nand U14332 (N_14332,N_14078,N_14145);
nor U14333 (N_14333,N_14174,N_14179);
or U14334 (N_14334,N_14192,N_14034);
or U14335 (N_14335,N_14080,N_14212);
nand U14336 (N_14336,N_14181,N_14215);
and U14337 (N_14337,N_14249,N_14018);
xor U14338 (N_14338,N_14105,N_14152);
nor U14339 (N_14339,N_14030,N_14093);
or U14340 (N_14340,N_14234,N_14059);
nor U14341 (N_14341,N_14070,N_14178);
xor U14342 (N_14342,N_14244,N_14167);
or U14343 (N_14343,N_14156,N_14227);
xnor U14344 (N_14344,N_14221,N_14101);
and U14345 (N_14345,N_14205,N_14027);
and U14346 (N_14346,N_14134,N_14150);
xnor U14347 (N_14347,N_14111,N_14069);
nor U14348 (N_14348,N_14117,N_14200);
nor U14349 (N_14349,N_14112,N_14213);
or U14350 (N_14350,N_14207,N_14128);
nor U14351 (N_14351,N_14012,N_14087);
or U14352 (N_14352,N_14141,N_14076);
and U14353 (N_14353,N_14017,N_14219);
and U14354 (N_14354,N_14024,N_14001);
nor U14355 (N_14355,N_14155,N_14148);
or U14356 (N_14356,N_14228,N_14066);
nand U14357 (N_14357,N_14135,N_14008);
nor U14358 (N_14358,N_14126,N_14051);
xnor U14359 (N_14359,N_14011,N_14175);
xor U14360 (N_14360,N_14043,N_14157);
or U14361 (N_14361,N_14243,N_14199);
nor U14362 (N_14362,N_14172,N_14103);
and U14363 (N_14363,N_14183,N_14247);
or U14364 (N_14364,N_14019,N_14107);
nor U14365 (N_14365,N_14067,N_14120);
xnor U14366 (N_14366,N_14225,N_14210);
nor U14367 (N_14367,N_14100,N_14074);
and U14368 (N_14368,N_14169,N_14026);
and U14369 (N_14369,N_14130,N_14202);
or U14370 (N_14370,N_14085,N_14160);
nor U14371 (N_14371,N_14106,N_14206);
nand U14372 (N_14372,N_14198,N_14185);
xor U14373 (N_14373,N_14089,N_14035);
and U14374 (N_14374,N_14032,N_14081);
or U14375 (N_14375,N_14071,N_14104);
nor U14376 (N_14376,N_14027,N_14192);
nor U14377 (N_14377,N_14180,N_14201);
nor U14378 (N_14378,N_14073,N_14164);
nand U14379 (N_14379,N_14028,N_14182);
nor U14380 (N_14380,N_14227,N_14244);
nand U14381 (N_14381,N_14002,N_14200);
nor U14382 (N_14382,N_14033,N_14036);
and U14383 (N_14383,N_14153,N_14009);
nand U14384 (N_14384,N_14114,N_14231);
nor U14385 (N_14385,N_14239,N_14220);
nor U14386 (N_14386,N_14023,N_14022);
and U14387 (N_14387,N_14038,N_14008);
or U14388 (N_14388,N_14192,N_14121);
and U14389 (N_14389,N_14206,N_14212);
or U14390 (N_14390,N_14052,N_14007);
and U14391 (N_14391,N_14014,N_14192);
and U14392 (N_14392,N_14181,N_14154);
nor U14393 (N_14393,N_14034,N_14195);
nand U14394 (N_14394,N_14220,N_14159);
xor U14395 (N_14395,N_14204,N_14050);
nor U14396 (N_14396,N_14095,N_14000);
nand U14397 (N_14397,N_14009,N_14092);
nand U14398 (N_14398,N_14069,N_14208);
and U14399 (N_14399,N_14032,N_14192);
nor U14400 (N_14400,N_14133,N_14139);
nand U14401 (N_14401,N_14089,N_14033);
nand U14402 (N_14402,N_14120,N_14162);
or U14403 (N_14403,N_14010,N_14029);
and U14404 (N_14404,N_14156,N_14151);
xor U14405 (N_14405,N_14210,N_14195);
nor U14406 (N_14406,N_14122,N_14105);
and U14407 (N_14407,N_14089,N_14229);
or U14408 (N_14408,N_14071,N_14073);
nor U14409 (N_14409,N_14187,N_14115);
xnor U14410 (N_14410,N_14049,N_14043);
and U14411 (N_14411,N_14170,N_14161);
nor U14412 (N_14412,N_14224,N_14181);
and U14413 (N_14413,N_14249,N_14165);
nand U14414 (N_14414,N_14149,N_14192);
or U14415 (N_14415,N_14177,N_14096);
nor U14416 (N_14416,N_14005,N_14022);
nor U14417 (N_14417,N_14032,N_14243);
nor U14418 (N_14418,N_14111,N_14015);
xor U14419 (N_14419,N_14240,N_14188);
nand U14420 (N_14420,N_14039,N_14227);
nor U14421 (N_14421,N_14227,N_14004);
and U14422 (N_14422,N_14122,N_14245);
and U14423 (N_14423,N_14094,N_14038);
nand U14424 (N_14424,N_14178,N_14241);
and U14425 (N_14425,N_14167,N_14156);
and U14426 (N_14426,N_14198,N_14238);
nand U14427 (N_14427,N_14178,N_14114);
or U14428 (N_14428,N_14234,N_14125);
and U14429 (N_14429,N_14218,N_14231);
or U14430 (N_14430,N_14051,N_14120);
nand U14431 (N_14431,N_14100,N_14059);
nor U14432 (N_14432,N_14126,N_14016);
nor U14433 (N_14433,N_14141,N_14043);
nand U14434 (N_14434,N_14159,N_14040);
and U14435 (N_14435,N_14181,N_14115);
and U14436 (N_14436,N_14053,N_14188);
or U14437 (N_14437,N_14206,N_14066);
nor U14438 (N_14438,N_14203,N_14030);
or U14439 (N_14439,N_14038,N_14199);
nor U14440 (N_14440,N_14184,N_14244);
or U14441 (N_14441,N_14103,N_14035);
and U14442 (N_14442,N_14237,N_14057);
nand U14443 (N_14443,N_14062,N_14228);
or U14444 (N_14444,N_14106,N_14199);
nor U14445 (N_14445,N_14114,N_14025);
or U14446 (N_14446,N_14169,N_14195);
or U14447 (N_14447,N_14124,N_14196);
or U14448 (N_14448,N_14082,N_14150);
nand U14449 (N_14449,N_14064,N_14140);
nor U14450 (N_14450,N_14131,N_14135);
nor U14451 (N_14451,N_14084,N_14229);
nor U14452 (N_14452,N_14063,N_14097);
nor U14453 (N_14453,N_14004,N_14143);
nor U14454 (N_14454,N_14108,N_14163);
or U14455 (N_14455,N_14241,N_14020);
or U14456 (N_14456,N_14186,N_14017);
nor U14457 (N_14457,N_14093,N_14180);
nand U14458 (N_14458,N_14117,N_14013);
and U14459 (N_14459,N_14015,N_14098);
nor U14460 (N_14460,N_14000,N_14170);
and U14461 (N_14461,N_14061,N_14081);
or U14462 (N_14462,N_14130,N_14093);
nand U14463 (N_14463,N_14103,N_14093);
or U14464 (N_14464,N_14110,N_14219);
nor U14465 (N_14465,N_14012,N_14187);
nand U14466 (N_14466,N_14196,N_14234);
and U14467 (N_14467,N_14088,N_14041);
xnor U14468 (N_14468,N_14189,N_14018);
nand U14469 (N_14469,N_14210,N_14185);
nand U14470 (N_14470,N_14224,N_14151);
nor U14471 (N_14471,N_14024,N_14062);
nor U14472 (N_14472,N_14045,N_14222);
nor U14473 (N_14473,N_14153,N_14233);
nand U14474 (N_14474,N_14210,N_14009);
nand U14475 (N_14475,N_14206,N_14233);
nor U14476 (N_14476,N_14093,N_14211);
nor U14477 (N_14477,N_14192,N_14151);
nor U14478 (N_14478,N_14160,N_14236);
or U14479 (N_14479,N_14106,N_14025);
and U14480 (N_14480,N_14088,N_14161);
nor U14481 (N_14481,N_14094,N_14033);
nand U14482 (N_14482,N_14060,N_14045);
nor U14483 (N_14483,N_14094,N_14057);
and U14484 (N_14484,N_14183,N_14152);
and U14485 (N_14485,N_14007,N_14094);
nand U14486 (N_14486,N_14170,N_14021);
nor U14487 (N_14487,N_14098,N_14122);
or U14488 (N_14488,N_14070,N_14103);
or U14489 (N_14489,N_14245,N_14148);
or U14490 (N_14490,N_14007,N_14166);
xor U14491 (N_14491,N_14116,N_14137);
and U14492 (N_14492,N_14003,N_14211);
and U14493 (N_14493,N_14104,N_14091);
nor U14494 (N_14494,N_14054,N_14114);
nand U14495 (N_14495,N_14153,N_14191);
nand U14496 (N_14496,N_14111,N_14079);
nor U14497 (N_14497,N_14022,N_14126);
nor U14498 (N_14498,N_14075,N_14039);
or U14499 (N_14499,N_14178,N_14011);
nor U14500 (N_14500,N_14471,N_14368);
and U14501 (N_14501,N_14280,N_14260);
nand U14502 (N_14502,N_14311,N_14296);
nor U14503 (N_14503,N_14343,N_14393);
or U14504 (N_14504,N_14415,N_14364);
nand U14505 (N_14505,N_14365,N_14372);
nor U14506 (N_14506,N_14265,N_14403);
nand U14507 (N_14507,N_14346,N_14470);
or U14508 (N_14508,N_14307,N_14392);
or U14509 (N_14509,N_14273,N_14310);
or U14510 (N_14510,N_14384,N_14448);
xnor U14511 (N_14511,N_14254,N_14308);
nand U14512 (N_14512,N_14333,N_14405);
or U14513 (N_14513,N_14450,N_14295);
xnor U14514 (N_14514,N_14477,N_14290);
nor U14515 (N_14515,N_14267,N_14465);
nor U14516 (N_14516,N_14467,N_14386);
nor U14517 (N_14517,N_14288,N_14257);
and U14518 (N_14518,N_14278,N_14447);
xnor U14519 (N_14519,N_14395,N_14277);
or U14520 (N_14520,N_14313,N_14420);
nor U14521 (N_14521,N_14391,N_14256);
nand U14522 (N_14522,N_14468,N_14371);
or U14523 (N_14523,N_14418,N_14279);
and U14524 (N_14524,N_14414,N_14266);
or U14525 (N_14525,N_14359,N_14322);
nand U14526 (N_14526,N_14457,N_14432);
nor U14527 (N_14527,N_14453,N_14426);
nor U14528 (N_14528,N_14408,N_14360);
xnor U14529 (N_14529,N_14258,N_14251);
or U14530 (N_14530,N_14250,N_14422);
xor U14531 (N_14531,N_14319,N_14263);
nor U14532 (N_14532,N_14373,N_14487);
nor U14533 (N_14533,N_14276,N_14361);
nor U14534 (N_14534,N_14321,N_14261);
or U14535 (N_14535,N_14340,N_14462);
nor U14536 (N_14536,N_14452,N_14349);
nor U14537 (N_14537,N_14388,N_14486);
xor U14538 (N_14538,N_14375,N_14379);
nand U14539 (N_14539,N_14406,N_14402);
or U14540 (N_14540,N_14433,N_14301);
and U14541 (N_14541,N_14429,N_14304);
xnor U14542 (N_14542,N_14347,N_14382);
nor U14543 (N_14543,N_14376,N_14456);
nor U14544 (N_14544,N_14445,N_14297);
nor U14545 (N_14545,N_14374,N_14412);
or U14546 (N_14546,N_14454,N_14305);
or U14547 (N_14547,N_14272,N_14460);
nor U14548 (N_14548,N_14337,N_14383);
xor U14549 (N_14549,N_14317,N_14396);
xor U14550 (N_14550,N_14427,N_14262);
nand U14551 (N_14551,N_14355,N_14293);
nor U14552 (N_14552,N_14281,N_14320);
xor U14553 (N_14553,N_14463,N_14303);
or U14554 (N_14554,N_14252,N_14345);
nand U14555 (N_14555,N_14430,N_14394);
nor U14556 (N_14556,N_14271,N_14398);
xor U14557 (N_14557,N_14299,N_14356);
and U14558 (N_14558,N_14341,N_14275);
or U14559 (N_14559,N_14397,N_14302);
xor U14560 (N_14560,N_14323,N_14497);
xor U14561 (N_14561,N_14409,N_14440);
xnor U14562 (N_14562,N_14259,N_14464);
nor U14563 (N_14563,N_14357,N_14475);
nand U14564 (N_14564,N_14270,N_14421);
and U14565 (N_14565,N_14329,N_14253);
or U14566 (N_14566,N_14424,N_14435);
and U14567 (N_14567,N_14300,N_14411);
nor U14568 (N_14568,N_14439,N_14351);
or U14569 (N_14569,N_14327,N_14385);
xnor U14570 (N_14570,N_14399,N_14413);
or U14571 (N_14571,N_14315,N_14476);
xnor U14572 (N_14572,N_14331,N_14268);
or U14573 (N_14573,N_14335,N_14472);
xnor U14574 (N_14574,N_14494,N_14255);
xnor U14575 (N_14575,N_14401,N_14342);
or U14576 (N_14576,N_14498,N_14483);
or U14577 (N_14577,N_14469,N_14489);
nor U14578 (N_14578,N_14478,N_14442);
xor U14579 (N_14579,N_14474,N_14285);
nand U14580 (N_14580,N_14289,N_14325);
and U14581 (N_14581,N_14479,N_14284);
or U14582 (N_14582,N_14370,N_14423);
nand U14583 (N_14583,N_14380,N_14283);
nand U14584 (N_14584,N_14490,N_14328);
nand U14585 (N_14585,N_14353,N_14496);
or U14586 (N_14586,N_14390,N_14344);
nand U14587 (N_14587,N_14458,N_14377);
and U14588 (N_14588,N_14488,N_14264);
and U14589 (N_14589,N_14428,N_14416);
or U14590 (N_14590,N_14298,N_14358);
nand U14591 (N_14591,N_14389,N_14438);
nor U14592 (N_14592,N_14334,N_14348);
nor U14593 (N_14593,N_14352,N_14367);
xor U14594 (N_14594,N_14437,N_14354);
or U14595 (N_14595,N_14436,N_14292);
or U14596 (N_14596,N_14291,N_14446);
nand U14597 (N_14597,N_14407,N_14484);
or U14598 (N_14598,N_14366,N_14434);
nor U14599 (N_14599,N_14330,N_14449);
or U14600 (N_14600,N_14318,N_14419);
nand U14601 (N_14601,N_14410,N_14482);
and U14602 (N_14602,N_14400,N_14495);
nor U14603 (N_14603,N_14339,N_14294);
or U14604 (N_14604,N_14274,N_14441);
nand U14605 (N_14605,N_14480,N_14369);
or U14606 (N_14606,N_14431,N_14481);
and U14607 (N_14607,N_14417,N_14444);
nor U14608 (N_14608,N_14332,N_14363);
and U14609 (N_14609,N_14381,N_14485);
nor U14610 (N_14610,N_14378,N_14306);
nand U14611 (N_14611,N_14404,N_14309);
nand U14612 (N_14612,N_14336,N_14499);
nand U14613 (N_14613,N_14350,N_14338);
nor U14614 (N_14614,N_14459,N_14286);
and U14615 (N_14615,N_14387,N_14425);
xor U14616 (N_14616,N_14455,N_14287);
or U14617 (N_14617,N_14451,N_14493);
and U14618 (N_14618,N_14473,N_14314);
and U14619 (N_14619,N_14491,N_14466);
nor U14620 (N_14620,N_14362,N_14324);
xnor U14621 (N_14621,N_14443,N_14312);
or U14622 (N_14622,N_14492,N_14282);
nor U14623 (N_14623,N_14269,N_14461);
nand U14624 (N_14624,N_14326,N_14316);
nor U14625 (N_14625,N_14390,N_14323);
nand U14626 (N_14626,N_14417,N_14436);
nand U14627 (N_14627,N_14274,N_14385);
or U14628 (N_14628,N_14433,N_14343);
or U14629 (N_14629,N_14294,N_14427);
nor U14630 (N_14630,N_14257,N_14379);
nor U14631 (N_14631,N_14397,N_14390);
and U14632 (N_14632,N_14361,N_14431);
or U14633 (N_14633,N_14405,N_14432);
or U14634 (N_14634,N_14263,N_14455);
nand U14635 (N_14635,N_14310,N_14280);
xnor U14636 (N_14636,N_14258,N_14274);
and U14637 (N_14637,N_14300,N_14366);
nor U14638 (N_14638,N_14388,N_14358);
or U14639 (N_14639,N_14480,N_14291);
xor U14640 (N_14640,N_14356,N_14283);
nor U14641 (N_14641,N_14384,N_14326);
or U14642 (N_14642,N_14481,N_14443);
and U14643 (N_14643,N_14459,N_14318);
nand U14644 (N_14644,N_14325,N_14462);
or U14645 (N_14645,N_14409,N_14287);
nor U14646 (N_14646,N_14313,N_14378);
nand U14647 (N_14647,N_14349,N_14315);
or U14648 (N_14648,N_14358,N_14267);
nand U14649 (N_14649,N_14386,N_14356);
and U14650 (N_14650,N_14269,N_14312);
nor U14651 (N_14651,N_14497,N_14457);
nor U14652 (N_14652,N_14434,N_14271);
and U14653 (N_14653,N_14260,N_14353);
or U14654 (N_14654,N_14353,N_14400);
nor U14655 (N_14655,N_14420,N_14338);
and U14656 (N_14656,N_14428,N_14410);
and U14657 (N_14657,N_14464,N_14250);
nand U14658 (N_14658,N_14297,N_14318);
or U14659 (N_14659,N_14414,N_14412);
xnor U14660 (N_14660,N_14378,N_14407);
and U14661 (N_14661,N_14427,N_14252);
and U14662 (N_14662,N_14314,N_14368);
nand U14663 (N_14663,N_14460,N_14271);
nor U14664 (N_14664,N_14351,N_14353);
and U14665 (N_14665,N_14397,N_14393);
and U14666 (N_14666,N_14372,N_14352);
xor U14667 (N_14667,N_14485,N_14283);
xor U14668 (N_14668,N_14288,N_14307);
nand U14669 (N_14669,N_14260,N_14360);
or U14670 (N_14670,N_14252,N_14451);
or U14671 (N_14671,N_14285,N_14469);
nor U14672 (N_14672,N_14484,N_14314);
and U14673 (N_14673,N_14398,N_14383);
or U14674 (N_14674,N_14482,N_14463);
nor U14675 (N_14675,N_14456,N_14379);
nor U14676 (N_14676,N_14453,N_14322);
or U14677 (N_14677,N_14334,N_14316);
nor U14678 (N_14678,N_14470,N_14402);
or U14679 (N_14679,N_14277,N_14463);
or U14680 (N_14680,N_14253,N_14375);
or U14681 (N_14681,N_14388,N_14369);
nor U14682 (N_14682,N_14412,N_14387);
nor U14683 (N_14683,N_14279,N_14469);
nand U14684 (N_14684,N_14307,N_14262);
nor U14685 (N_14685,N_14290,N_14268);
nor U14686 (N_14686,N_14266,N_14399);
and U14687 (N_14687,N_14460,N_14497);
nor U14688 (N_14688,N_14413,N_14301);
or U14689 (N_14689,N_14282,N_14497);
nor U14690 (N_14690,N_14494,N_14303);
and U14691 (N_14691,N_14473,N_14339);
nor U14692 (N_14692,N_14277,N_14367);
nand U14693 (N_14693,N_14497,N_14379);
and U14694 (N_14694,N_14346,N_14279);
and U14695 (N_14695,N_14292,N_14463);
or U14696 (N_14696,N_14418,N_14262);
or U14697 (N_14697,N_14312,N_14387);
nor U14698 (N_14698,N_14467,N_14455);
nand U14699 (N_14699,N_14288,N_14340);
or U14700 (N_14700,N_14455,N_14291);
nand U14701 (N_14701,N_14419,N_14438);
or U14702 (N_14702,N_14424,N_14483);
nor U14703 (N_14703,N_14495,N_14412);
nand U14704 (N_14704,N_14496,N_14464);
and U14705 (N_14705,N_14400,N_14369);
and U14706 (N_14706,N_14451,N_14393);
or U14707 (N_14707,N_14277,N_14366);
nand U14708 (N_14708,N_14293,N_14396);
nor U14709 (N_14709,N_14354,N_14308);
nand U14710 (N_14710,N_14293,N_14413);
or U14711 (N_14711,N_14408,N_14402);
or U14712 (N_14712,N_14407,N_14394);
nand U14713 (N_14713,N_14317,N_14431);
and U14714 (N_14714,N_14493,N_14340);
nand U14715 (N_14715,N_14327,N_14278);
nand U14716 (N_14716,N_14476,N_14414);
nor U14717 (N_14717,N_14381,N_14285);
or U14718 (N_14718,N_14372,N_14388);
and U14719 (N_14719,N_14293,N_14313);
and U14720 (N_14720,N_14276,N_14377);
nand U14721 (N_14721,N_14409,N_14486);
nand U14722 (N_14722,N_14335,N_14357);
nand U14723 (N_14723,N_14300,N_14312);
nand U14724 (N_14724,N_14486,N_14407);
and U14725 (N_14725,N_14415,N_14379);
or U14726 (N_14726,N_14313,N_14259);
and U14727 (N_14727,N_14456,N_14306);
xnor U14728 (N_14728,N_14341,N_14390);
or U14729 (N_14729,N_14479,N_14253);
or U14730 (N_14730,N_14393,N_14372);
nor U14731 (N_14731,N_14270,N_14378);
and U14732 (N_14732,N_14406,N_14327);
or U14733 (N_14733,N_14336,N_14355);
or U14734 (N_14734,N_14316,N_14435);
nor U14735 (N_14735,N_14484,N_14300);
nand U14736 (N_14736,N_14443,N_14465);
or U14737 (N_14737,N_14288,N_14255);
or U14738 (N_14738,N_14416,N_14363);
and U14739 (N_14739,N_14377,N_14494);
or U14740 (N_14740,N_14443,N_14396);
and U14741 (N_14741,N_14367,N_14374);
nand U14742 (N_14742,N_14488,N_14463);
or U14743 (N_14743,N_14372,N_14271);
nand U14744 (N_14744,N_14452,N_14325);
or U14745 (N_14745,N_14327,N_14494);
or U14746 (N_14746,N_14342,N_14421);
or U14747 (N_14747,N_14280,N_14319);
and U14748 (N_14748,N_14287,N_14310);
or U14749 (N_14749,N_14442,N_14384);
xor U14750 (N_14750,N_14595,N_14612);
or U14751 (N_14751,N_14626,N_14680);
and U14752 (N_14752,N_14731,N_14539);
xnor U14753 (N_14753,N_14651,N_14535);
and U14754 (N_14754,N_14698,N_14544);
xnor U14755 (N_14755,N_14510,N_14693);
nor U14756 (N_14756,N_14649,N_14563);
nor U14757 (N_14757,N_14660,N_14537);
or U14758 (N_14758,N_14621,N_14507);
nor U14759 (N_14759,N_14548,N_14723);
nand U14760 (N_14760,N_14691,N_14591);
nor U14761 (N_14761,N_14629,N_14619);
nand U14762 (N_14762,N_14589,N_14526);
or U14763 (N_14763,N_14650,N_14711);
nor U14764 (N_14764,N_14538,N_14746);
and U14765 (N_14765,N_14594,N_14632);
nand U14766 (N_14766,N_14631,N_14547);
and U14767 (N_14767,N_14610,N_14648);
xnor U14768 (N_14768,N_14713,N_14639);
and U14769 (N_14769,N_14509,N_14505);
and U14770 (N_14770,N_14551,N_14502);
or U14771 (N_14771,N_14749,N_14607);
nor U14772 (N_14772,N_14617,N_14721);
nand U14773 (N_14773,N_14730,N_14670);
and U14774 (N_14774,N_14733,N_14618);
or U14775 (N_14775,N_14518,N_14641);
xnor U14776 (N_14776,N_14716,N_14704);
nor U14777 (N_14777,N_14702,N_14673);
nor U14778 (N_14778,N_14569,N_14598);
xor U14779 (N_14779,N_14703,N_14732);
nand U14780 (N_14780,N_14655,N_14748);
and U14781 (N_14781,N_14540,N_14735);
nand U14782 (N_14782,N_14678,N_14728);
nor U14783 (N_14783,N_14644,N_14636);
or U14784 (N_14784,N_14599,N_14506);
and U14785 (N_14785,N_14688,N_14571);
nor U14786 (N_14786,N_14508,N_14683);
xor U14787 (N_14787,N_14593,N_14564);
and U14788 (N_14788,N_14581,N_14533);
xor U14789 (N_14789,N_14685,N_14675);
nand U14790 (N_14790,N_14582,N_14602);
and U14791 (N_14791,N_14725,N_14737);
or U14792 (N_14792,N_14729,N_14630);
nand U14793 (N_14793,N_14714,N_14664);
and U14794 (N_14794,N_14718,N_14740);
and U14795 (N_14795,N_14623,N_14640);
or U14796 (N_14796,N_14739,N_14588);
nand U14797 (N_14797,N_14604,N_14567);
nor U14798 (N_14798,N_14738,N_14661);
nand U14799 (N_14799,N_14642,N_14500);
and U14800 (N_14800,N_14541,N_14565);
or U14801 (N_14801,N_14719,N_14579);
nand U14802 (N_14802,N_14734,N_14580);
and U14803 (N_14803,N_14592,N_14558);
nand U14804 (N_14804,N_14634,N_14628);
nand U14805 (N_14805,N_14549,N_14705);
nor U14806 (N_14806,N_14727,N_14695);
nand U14807 (N_14807,N_14736,N_14679);
xor U14808 (N_14808,N_14674,N_14609);
nand U14809 (N_14809,N_14536,N_14552);
and U14810 (N_14810,N_14543,N_14525);
or U14811 (N_14811,N_14597,N_14521);
nand U14812 (N_14812,N_14692,N_14656);
xor U14813 (N_14813,N_14556,N_14722);
or U14814 (N_14814,N_14585,N_14701);
xnor U14815 (N_14815,N_14653,N_14530);
nand U14816 (N_14816,N_14577,N_14687);
nand U14817 (N_14817,N_14646,N_14720);
or U14818 (N_14818,N_14625,N_14570);
nor U14819 (N_14819,N_14643,N_14635);
nand U14820 (N_14820,N_14501,N_14503);
and U14821 (N_14821,N_14613,N_14645);
xnor U14822 (N_14822,N_14696,N_14712);
nor U14823 (N_14823,N_14677,N_14668);
and U14824 (N_14824,N_14504,N_14710);
nor U14825 (N_14825,N_14647,N_14513);
or U14826 (N_14826,N_14605,N_14559);
nor U14827 (N_14827,N_14534,N_14574);
xor U14828 (N_14828,N_14554,N_14608);
nand U14829 (N_14829,N_14708,N_14615);
nand U14830 (N_14830,N_14747,N_14614);
and U14831 (N_14831,N_14700,N_14524);
nand U14832 (N_14832,N_14663,N_14568);
nor U14833 (N_14833,N_14743,N_14527);
nor U14834 (N_14834,N_14652,N_14633);
or U14835 (N_14835,N_14516,N_14697);
nor U14836 (N_14836,N_14709,N_14726);
and U14837 (N_14837,N_14522,N_14627);
or U14838 (N_14838,N_14745,N_14699);
and U14839 (N_14839,N_14694,N_14603);
nand U14840 (N_14840,N_14690,N_14658);
and U14841 (N_14841,N_14555,N_14715);
nor U14842 (N_14842,N_14511,N_14662);
nor U14843 (N_14843,N_14666,N_14572);
xor U14844 (N_14844,N_14573,N_14596);
nor U14845 (N_14845,N_14672,N_14657);
or U14846 (N_14846,N_14566,N_14560);
nor U14847 (N_14847,N_14744,N_14590);
nand U14848 (N_14848,N_14584,N_14682);
and U14849 (N_14849,N_14724,N_14638);
nor U14850 (N_14850,N_14586,N_14553);
or U14851 (N_14851,N_14557,N_14611);
nor U14852 (N_14852,N_14706,N_14545);
nor U14853 (N_14853,N_14616,N_14671);
or U14854 (N_14854,N_14514,N_14717);
nand U14855 (N_14855,N_14575,N_14659);
and U14856 (N_14856,N_14519,N_14561);
and U14857 (N_14857,N_14689,N_14523);
or U14858 (N_14858,N_14532,N_14546);
nand U14859 (N_14859,N_14669,N_14562);
and U14860 (N_14860,N_14531,N_14667);
or U14861 (N_14861,N_14606,N_14542);
nand U14862 (N_14862,N_14654,N_14601);
nor U14863 (N_14863,N_14550,N_14681);
xnor U14864 (N_14864,N_14620,N_14665);
or U14865 (N_14865,N_14600,N_14707);
or U14866 (N_14866,N_14676,N_14583);
nand U14867 (N_14867,N_14742,N_14622);
and U14868 (N_14868,N_14637,N_14520);
nor U14869 (N_14869,N_14686,N_14578);
and U14870 (N_14870,N_14512,N_14587);
nand U14871 (N_14871,N_14684,N_14741);
and U14872 (N_14872,N_14528,N_14624);
xor U14873 (N_14873,N_14529,N_14517);
nand U14874 (N_14874,N_14576,N_14515);
and U14875 (N_14875,N_14611,N_14748);
nand U14876 (N_14876,N_14503,N_14551);
and U14877 (N_14877,N_14659,N_14558);
nor U14878 (N_14878,N_14729,N_14575);
or U14879 (N_14879,N_14576,N_14572);
or U14880 (N_14880,N_14591,N_14638);
nor U14881 (N_14881,N_14530,N_14721);
or U14882 (N_14882,N_14639,N_14650);
or U14883 (N_14883,N_14628,N_14528);
or U14884 (N_14884,N_14551,N_14586);
nor U14885 (N_14885,N_14667,N_14600);
and U14886 (N_14886,N_14608,N_14726);
nor U14887 (N_14887,N_14598,N_14661);
nand U14888 (N_14888,N_14613,N_14674);
or U14889 (N_14889,N_14695,N_14732);
xor U14890 (N_14890,N_14592,N_14671);
or U14891 (N_14891,N_14684,N_14564);
or U14892 (N_14892,N_14588,N_14586);
nand U14893 (N_14893,N_14633,N_14746);
nand U14894 (N_14894,N_14530,N_14733);
nor U14895 (N_14895,N_14629,N_14535);
nor U14896 (N_14896,N_14646,N_14516);
nor U14897 (N_14897,N_14511,N_14542);
and U14898 (N_14898,N_14623,N_14576);
nor U14899 (N_14899,N_14520,N_14705);
xor U14900 (N_14900,N_14574,N_14609);
and U14901 (N_14901,N_14527,N_14611);
or U14902 (N_14902,N_14742,N_14706);
and U14903 (N_14903,N_14536,N_14567);
and U14904 (N_14904,N_14638,N_14746);
and U14905 (N_14905,N_14546,N_14648);
and U14906 (N_14906,N_14635,N_14502);
xnor U14907 (N_14907,N_14544,N_14712);
or U14908 (N_14908,N_14669,N_14530);
nor U14909 (N_14909,N_14600,N_14711);
or U14910 (N_14910,N_14740,N_14513);
nand U14911 (N_14911,N_14548,N_14712);
and U14912 (N_14912,N_14659,N_14726);
and U14913 (N_14913,N_14641,N_14671);
or U14914 (N_14914,N_14534,N_14722);
nor U14915 (N_14915,N_14605,N_14706);
nor U14916 (N_14916,N_14654,N_14547);
and U14917 (N_14917,N_14643,N_14594);
nor U14918 (N_14918,N_14653,N_14554);
and U14919 (N_14919,N_14598,N_14736);
nor U14920 (N_14920,N_14611,N_14694);
nor U14921 (N_14921,N_14598,N_14514);
nor U14922 (N_14922,N_14642,N_14559);
nand U14923 (N_14923,N_14516,N_14575);
xor U14924 (N_14924,N_14728,N_14731);
and U14925 (N_14925,N_14689,N_14622);
and U14926 (N_14926,N_14524,N_14624);
nor U14927 (N_14927,N_14728,N_14522);
and U14928 (N_14928,N_14727,N_14511);
nand U14929 (N_14929,N_14673,N_14712);
nor U14930 (N_14930,N_14635,N_14566);
and U14931 (N_14931,N_14556,N_14549);
and U14932 (N_14932,N_14698,N_14562);
nand U14933 (N_14933,N_14726,N_14555);
xor U14934 (N_14934,N_14532,N_14564);
nand U14935 (N_14935,N_14508,N_14588);
nand U14936 (N_14936,N_14633,N_14707);
nor U14937 (N_14937,N_14671,N_14648);
and U14938 (N_14938,N_14648,N_14557);
and U14939 (N_14939,N_14636,N_14502);
nand U14940 (N_14940,N_14608,N_14595);
nor U14941 (N_14941,N_14603,N_14658);
and U14942 (N_14942,N_14566,N_14727);
xnor U14943 (N_14943,N_14501,N_14580);
nand U14944 (N_14944,N_14521,N_14524);
xnor U14945 (N_14945,N_14659,N_14512);
nand U14946 (N_14946,N_14553,N_14504);
nor U14947 (N_14947,N_14736,N_14686);
or U14948 (N_14948,N_14646,N_14685);
and U14949 (N_14949,N_14606,N_14562);
and U14950 (N_14950,N_14653,N_14515);
nand U14951 (N_14951,N_14608,N_14667);
nand U14952 (N_14952,N_14671,N_14621);
or U14953 (N_14953,N_14561,N_14650);
nand U14954 (N_14954,N_14694,N_14507);
or U14955 (N_14955,N_14565,N_14669);
nand U14956 (N_14956,N_14516,N_14547);
or U14957 (N_14957,N_14506,N_14603);
and U14958 (N_14958,N_14692,N_14623);
or U14959 (N_14959,N_14733,N_14537);
nor U14960 (N_14960,N_14623,N_14646);
and U14961 (N_14961,N_14634,N_14701);
nor U14962 (N_14962,N_14565,N_14647);
and U14963 (N_14963,N_14653,N_14717);
and U14964 (N_14964,N_14745,N_14626);
nor U14965 (N_14965,N_14506,N_14633);
and U14966 (N_14966,N_14673,N_14520);
xnor U14967 (N_14967,N_14583,N_14714);
or U14968 (N_14968,N_14714,N_14636);
nand U14969 (N_14969,N_14638,N_14555);
or U14970 (N_14970,N_14573,N_14660);
and U14971 (N_14971,N_14698,N_14601);
and U14972 (N_14972,N_14541,N_14736);
nand U14973 (N_14973,N_14651,N_14720);
or U14974 (N_14974,N_14565,N_14576);
and U14975 (N_14975,N_14626,N_14590);
nand U14976 (N_14976,N_14664,N_14641);
xnor U14977 (N_14977,N_14590,N_14530);
and U14978 (N_14978,N_14601,N_14694);
nand U14979 (N_14979,N_14534,N_14514);
nand U14980 (N_14980,N_14547,N_14742);
and U14981 (N_14981,N_14706,N_14529);
and U14982 (N_14982,N_14728,N_14707);
or U14983 (N_14983,N_14581,N_14604);
nand U14984 (N_14984,N_14555,N_14655);
nor U14985 (N_14985,N_14661,N_14586);
and U14986 (N_14986,N_14570,N_14735);
nor U14987 (N_14987,N_14551,N_14544);
nor U14988 (N_14988,N_14694,N_14595);
nand U14989 (N_14989,N_14686,N_14582);
nand U14990 (N_14990,N_14641,N_14714);
nor U14991 (N_14991,N_14636,N_14673);
nor U14992 (N_14992,N_14717,N_14561);
nor U14993 (N_14993,N_14517,N_14546);
nand U14994 (N_14994,N_14626,N_14733);
and U14995 (N_14995,N_14604,N_14646);
and U14996 (N_14996,N_14561,N_14634);
and U14997 (N_14997,N_14518,N_14626);
and U14998 (N_14998,N_14511,N_14650);
and U14999 (N_14999,N_14710,N_14658);
nand U15000 (N_15000,N_14865,N_14794);
nor U15001 (N_15001,N_14925,N_14762);
nor U15002 (N_15002,N_14864,N_14960);
nand U15003 (N_15003,N_14752,N_14991);
or U15004 (N_15004,N_14847,N_14940);
xnor U15005 (N_15005,N_14935,N_14826);
nor U15006 (N_15006,N_14905,N_14822);
nand U15007 (N_15007,N_14763,N_14926);
and U15008 (N_15008,N_14915,N_14963);
or U15009 (N_15009,N_14813,N_14814);
xor U15010 (N_15010,N_14977,N_14758);
nor U15011 (N_15011,N_14850,N_14823);
and U15012 (N_15012,N_14992,N_14891);
or U15013 (N_15013,N_14927,N_14999);
and U15014 (N_15014,N_14831,N_14860);
nand U15015 (N_15015,N_14945,N_14978);
xnor U15016 (N_15016,N_14983,N_14810);
and U15017 (N_15017,N_14791,N_14824);
or U15018 (N_15018,N_14816,N_14759);
or U15019 (N_15019,N_14884,N_14760);
and U15020 (N_15020,N_14754,N_14937);
nor U15021 (N_15021,N_14876,N_14962);
nand U15022 (N_15022,N_14885,N_14751);
nor U15023 (N_15023,N_14873,N_14859);
and U15024 (N_15024,N_14781,N_14775);
nor U15025 (N_15025,N_14782,N_14829);
nor U15026 (N_15026,N_14818,N_14770);
and U15027 (N_15027,N_14870,N_14966);
nor U15028 (N_15028,N_14776,N_14879);
nor U15029 (N_15029,N_14954,N_14750);
xnor U15030 (N_15030,N_14936,N_14808);
xor U15031 (N_15031,N_14863,N_14929);
xnor U15032 (N_15032,N_14861,N_14820);
nor U15033 (N_15033,N_14806,N_14947);
nor U15034 (N_15034,N_14757,N_14874);
nand U15035 (N_15035,N_14877,N_14792);
and U15036 (N_15036,N_14838,N_14788);
or U15037 (N_15037,N_14778,N_14812);
or U15038 (N_15038,N_14890,N_14867);
nor U15039 (N_15039,N_14761,N_14817);
or U15040 (N_15040,N_14968,N_14986);
or U15041 (N_15041,N_14881,N_14796);
or U15042 (N_15042,N_14793,N_14943);
xnor U15043 (N_15043,N_14857,N_14779);
nor U15044 (N_15044,N_14883,N_14953);
nand U15045 (N_15045,N_14755,N_14842);
nand U15046 (N_15046,N_14786,N_14764);
nand U15047 (N_15047,N_14771,N_14912);
nand U15048 (N_15048,N_14866,N_14923);
or U15049 (N_15049,N_14853,N_14997);
nand U15050 (N_15050,N_14783,N_14787);
or U15051 (N_15051,N_14875,N_14913);
nand U15052 (N_15052,N_14920,N_14766);
or U15053 (N_15053,N_14897,N_14805);
or U15054 (N_15054,N_14839,N_14854);
and U15055 (N_15055,N_14959,N_14888);
and U15056 (N_15056,N_14955,N_14941);
nor U15057 (N_15057,N_14772,N_14828);
and U15058 (N_15058,N_14996,N_14811);
nor U15059 (N_15059,N_14952,N_14894);
or U15060 (N_15060,N_14969,N_14918);
nand U15061 (N_15061,N_14834,N_14893);
or U15062 (N_15062,N_14949,N_14895);
or U15063 (N_15063,N_14835,N_14848);
or U15064 (N_15064,N_14851,N_14973);
and U15065 (N_15065,N_14769,N_14956);
xnor U15066 (N_15066,N_14798,N_14934);
nor U15067 (N_15067,N_14804,N_14914);
or U15068 (N_15068,N_14872,N_14980);
nand U15069 (N_15069,N_14801,N_14836);
nor U15070 (N_15070,N_14887,N_14768);
xor U15071 (N_15071,N_14832,N_14821);
nor U15072 (N_15072,N_14800,N_14948);
nand U15073 (N_15073,N_14880,N_14773);
xnor U15074 (N_15074,N_14930,N_14789);
and U15075 (N_15075,N_14998,N_14987);
nor U15076 (N_15076,N_14971,N_14931);
or U15077 (N_15077,N_14901,N_14862);
nor U15078 (N_15078,N_14827,N_14974);
and U15079 (N_15079,N_14855,N_14837);
nand U15080 (N_15080,N_14845,N_14988);
or U15081 (N_15081,N_14932,N_14904);
nand U15082 (N_15082,N_14922,N_14833);
nor U15083 (N_15083,N_14868,N_14843);
nor U15084 (N_15084,N_14964,N_14967);
and U15085 (N_15085,N_14858,N_14939);
and U15086 (N_15086,N_14938,N_14902);
xnor U15087 (N_15087,N_14797,N_14795);
or U15088 (N_15088,N_14957,N_14993);
xnor U15089 (N_15089,N_14976,N_14889);
or U15090 (N_15090,N_14911,N_14906);
or U15091 (N_15091,N_14970,N_14830);
or U15092 (N_15092,N_14944,N_14882);
or U15093 (N_15093,N_14753,N_14946);
nand U15094 (N_15094,N_14907,N_14765);
and U15095 (N_15095,N_14756,N_14958);
nand U15096 (N_15096,N_14989,N_14802);
nor U15097 (N_15097,N_14844,N_14965);
nand U15098 (N_15098,N_14908,N_14886);
xor U15099 (N_15099,N_14950,N_14928);
or U15100 (N_15100,N_14985,N_14990);
or U15101 (N_15101,N_14919,N_14899);
nand U15102 (N_15102,N_14924,N_14841);
nand U15103 (N_15103,N_14981,N_14979);
nand U15104 (N_15104,N_14780,N_14807);
and U15105 (N_15105,N_14921,N_14916);
and U15106 (N_15106,N_14825,N_14819);
xnor U15107 (N_15107,N_14917,N_14961);
nand U15108 (N_15108,N_14790,N_14910);
nor U15109 (N_15109,N_14774,N_14984);
nor U15110 (N_15110,N_14900,N_14846);
or U15111 (N_15111,N_14995,N_14849);
nor U15112 (N_15112,N_14975,N_14869);
or U15113 (N_15113,N_14815,N_14903);
and U15114 (N_15114,N_14785,N_14871);
and U15115 (N_15115,N_14852,N_14972);
nor U15116 (N_15116,N_14878,N_14892);
or U15117 (N_15117,N_14994,N_14982);
nand U15118 (N_15118,N_14803,N_14896);
nand U15119 (N_15119,N_14951,N_14856);
xor U15120 (N_15120,N_14909,N_14840);
or U15121 (N_15121,N_14809,N_14898);
nor U15122 (N_15122,N_14799,N_14777);
or U15123 (N_15123,N_14784,N_14942);
xnor U15124 (N_15124,N_14933,N_14767);
or U15125 (N_15125,N_14789,N_14780);
nand U15126 (N_15126,N_14978,N_14902);
nor U15127 (N_15127,N_14807,N_14806);
nand U15128 (N_15128,N_14751,N_14858);
nor U15129 (N_15129,N_14876,N_14864);
or U15130 (N_15130,N_14779,N_14963);
nor U15131 (N_15131,N_14922,N_14779);
nand U15132 (N_15132,N_14805,N_14924);
xnor U15133 (N_15133,N_14903,N_14926);
or U15134 (N_15134,N_14763,N_14865);
or U15135 (N_15135,N_14977,N_14943);
xor U15136 (N_15136,N_14871,N_14817);
xor U15137 (N_15137,N_14920,N_14997);
and U15138 (N_15138,N_14872,N_14933);
xnor U15139 (N_15139,N_14805,N_14849);
nor U15140 (N_15140,N_14859,N_14847);
or U15141 (N_15141,N_14954,N_14827);
nor U15142 (N_15142,N_14880,N_14987);
nand U15143 (N_15143,N_14996,N_14837);
nand U15144 (N_15144,N_14993,N_14917);
or U15145 (N_15145,N_14891,N_14782);
nand U15146 (N_15146,N_14847,N_14907);
xor U15147 (N_15147,N_14871,N_14998);
or U15148 (N_15148,N_14920,N_14790);
and U15149 (N_15149,N_14835,N_14759);
nor U15150 (N_15150,N_14814,N_14762);
nor U15151 (N_15151,N_14868,N_14929);
nor U15152 (N_15152,N_14971,N_14832);
or U15153 (N_15153,N_14788,N_14801);
nand U15154 (N_15154,N_14976,N_14810);
xnor U15155 (N_15155,N_14929,N_14961);
or U15156 (N_15156,N_14911,N_14932);
nand U15157 (N_15157,N_14969,N_14954);
and U15158 (N_15158,N_14789,N_14872);
nor U15159 (N_15159,N_14899,N_14750);
xor U15160 (N_15160,N_14758,N_14783);
nor U15161 (N_15161,N_14788,N_14970);
nand U15162 (N_15162,N_14946,N_14824);
or U15163 (N_15163,N_14885,N_14899);
and U15164 (N_15164,N_14954,N_14978);
or U15165 (N_15165,N_14839,N_14890);
or U15166 (N_15166,N_14872,N_14828);
nor U15167 (N_15167,N_14947,N_14838);
nand U15168 (N_15168,N_14808,N_14861);
and U15169 (N_15169,N_14890,N_14816);
nor U15170 (N_15170,N_14801,N_14908);
or U15171 (N_15171,N_14844,N_14853);
nand U15172 (N_15172,N_14761,N_14992);
nor U15173 (N_15173,N_14915,N_14927);
nor U15174 (N_15174,N_14798,N_14835);
nor U15175 (N_15175,N_14870,N_14760);
nand U15176 (N_15176,N_14907,N_14934);
nor U15177 (N_15177,N_14819,N_14763);
or U15178 (N_15178,N_14771,N_14831);
or U15179 (N_15179,N_14923,N_14779);
or U15180 (N_15180,N_14949,N_14914);
nand U15181 (N_15181,N_14854,N_14753);
or U15182 (N_15182,N_14851,N_14853);
nand U15183 (N_15183,N_14841,N_14986);
and U15184 (N_15184,N_14809,N_14753);
or U15185 (N_15185,N_14789,N_14822);
nand U15186 (N_15186,N_14952,N_14772);
or U15187 (N_15187,N_14780,N_14966);
or U15188 (N_15188,N_14933,N_14946);
and U15189 (N_15189,N_14750,N_14880);
or U15190 (N_15190,N_14825,N_14776);
xnor U15191 (N_15191,N_14820,N_14781);
nor U15192 (N_15192,N_14962,N_14893);
or U15193 (N_15193,N_14949,N_14971);
nor U15194 (N_15194,N_14902,N_14969);
nor U15195 (N_15195,N_14983,N_14990);
nor U15196 (N_15196,N_14874,N_14970);
nand U15197 (N_15197,N_14773,N_14874);
or U15198 (N_15198,N_14800,N_14772);
nand U15199 (N_15199,N_14816,N_14992);
nand U15200 (N_15200,N_14838,N_14912);
or U15201 (N_15201,N_14949,N_14840);
xnor U15202 (N_15202,N_14771,N_14819);
and U15203 (N_15203,N_14986,N_14858);
and U15204 (N_15204,N_14868,N_14899);
nand U15205 (N_15205,N_14989,N_14773);
nand U15206 (N_15206,N_14919,N_14948);
nor U15207 (N_15207,N_14786,N_14969);
nand U15208 (N_15208,N_14866,N_14946);
and U15209 (N_15209,N_14754,N_14953);
nand U15210 (N_15210,N_14894,N_14973);
xor U15211 (N_15211,N_14863,N_14873);
xnor U15212 (N_15212,N_14862,N_14861);
nand U15213 (N_15213,N_14848,N_14999);
and U15214 (N_15214,N_14980,N_14916);
or U15215 (N_15215,N_14997,N_14881);
xnor U15216 (N_15216,N_14925,N_14844);
nand U15217 (N_15217,N_14892,N_14903);
nand U15218 (N_15218,N_14981,N_14911);
and U15219 (N_15219,N_14962,N_14957);
xnor U15220 (N_15220,N_14792,N_14795);
and U15221 (N_15221,N_14752,N_14777);
nand U15222 (N_15222,N_14988,N_14853);
nand U15223 (N_15223,N_14792,N_14762);
and U15224 (N_15224,N_14986,N_14788);
nor U15225 (N_15225,N_14832,N_14894);
or U15226 (N_15226,N_14973,N_14977);
nor U15227 (N_15227,N_14972,N_14857);
or U15228 (N_15228,N_14916,N_14986);
xnor U15229 (N_15229,N_14917,N_14984);
and U15230 (N_15230,N_14906,N_14832);
or U15231 (N_15231,N_14973,N_14818);
or U15232 (N_15232,N_14975,N_14855);
nand U15233 (N_15233,N_14934,N_14884);
or U15234 (N_15234,N_14870,N_14952);
or U15235 (N_15235,N_14860,N_14875);
nand U15236 (N_15236,N_14992,N_14795);
or U15237 (N_15237,N_14798,N_14969);
xor U15238 (N_15238,N_14828,N_14932);
or U15239 (N_15239,N_14851,N_14902);
or U15240 (N_15240,N_14947,N_14954);
or U15241 (N_15241,N_14931,N_14801);
nand U15242 (N_15242,N_14865,N_14885);
xnor U15243 (N_15243,N_14973,N_14865);
and U15244 (N_15244,N_14948,N_14828);
nand U15245 (N_15245,N_14761,N_14766);
nand U15246 (N_15246,N_14851,N_14797);
nand U15247 (N_15247,N_14903,N_14989);
nand U15248 (N_15248,N_14763,N_14933);
and U15249 (N_15249,N_14855,N_14958);
xnor U15250 (N_15250,N_15063,N_15036);
nand U15251 (N_15251,N_15126,N_15231);
nor U15252 (N_15252,N_15054,N_15176);
nor U15253 (N_15253,N_15027,N_15028);
nand U15254 (N_15254,N_15211,N_15012);
or U15255 (N_15255,N_15050,N_15216);
nor U15256 (N_15256,N_15144,N_15142);
or U15257 (N_15257,N_15242,N_15114);
nand U15258 (N_15258,N_15119,N_15112);
nor U15259 (N_15259,N_15009,N_15210);
nand U15260 (N_15260,N_15171,N_15059);
or U15261 (N_15261,N_15104,N_15090);
and U15262 (N_15262,N_15219,N_15020);
nor U15263 (N_15263,N_15046,N_15130);
nand U15264 (N_15264,N_15241,N_15209);
and U15265 (N_15265,N_15147,N_15083);
nand U15266 (N_15266,N_15017,N_15151);
or U15267 (N_15267,N_15014,N_15096);
nand U15268 (N_15268,N_15071,N_15229);
nand U15269 (N_15269,N_15178,N_15057);
nor U15270 (N_15270,N_15196,N_15105);
and U15271 (N_15271,N_15115,N_15010);
and U15272 (N_15272,N_15111,N_15032);
or U15273 (N_15273,N_15035,N_15238);
or U15274 (N_15274,N_15169,N_15011);
or U15275 (N_15275,N_15019,N_15204);
or U15276 (N_15276,N_15002,N_15086);
nand U15277 (N_15277,N_15234,N_15110);
nor U15278 (N_15278,N_15179,N_15199);
and U15279 (N_15279,N_15088,N_15116);
or U15280 (N_15280,N_15207,N_15053);
and U15281 (N_15281,N_15038,N_15079);
and U15282 (N_15282,N_15099,N_15021);
nor U15283 (N_15283,N_15244,N_15190);
and U15284 (N_15284,N_15180,N_15093);
nor U15285 (N_15285,N_15158,N_15015);
nor U15286 (N_15286,N_15206,N_15137);
nand U15287 (N_15287,N_15198,N_15228);
and U15288 (N_15288,N_15183,N_15163);
or U15289 (N_15289,N_15201,N_15120);
or U15290 (N_15290,N_15108,N_15162);
and U15291 (N_15291,N_15165,N_15177);
nand U15292 (N_15292,N_15166,N_15107);
nor U15293 (N_15293,N_15246,N_15194);
and U15294 (N_15294,N_15000,N_15016);
or U15295 (N_15295,N_15221,N_15058);
nor U15296 (N_15296,N_15202,N_15129);
nor U15297 (N_15297,N_15157,N_15139);
or U15298 (N_15298,N_15133,N_15066);
and U15299 (N_15299,N_15153,N_15131);
nor U15300 (N_15300,N_15239,N_15005);
xnor U15301 (N_15301,N_15067,N_15042);
nor U15302 (N_15302,N_15001,N_15217);
and U15303 (N_15303,N_15135,N_15127);
and U15304 (N_15304,N_15152,N_15249);
xor U15305 (N_15305,N_15212,N_15245);
nand U15306 (N_15306,N_15182,N_15013);
nand U15307 (N_15307,N_15047,N_15055);
nor U15308 (N_15308,N_15215,N_15026);
and U15309 (N_15309,N_15225,N_15154);
or U15310 (N_15310,N_15213,N_15006);
and U15311 (N_15311,N_15197,N_15173);
xnor U15312 (N_15312,N_15195,N_15024);
nand U15313 (N_15313,N_15193,N_15175);
xnor U15314 (N_15314,N_15069,N_15168);
or U15315 (N_15315,N_15141,N_15061);
or U15316 (N_15316,N_15188,N_15072);
xor U15317 (N_15317,N_15200,N_15117);
and U15318 (N_15318,N_15094,N_15164);
nand U15319 (N_15319,N_15121,N_15143);
nand U15320 (N_15320,N_15167,N_15076);
xor U15321 (N_15321,N_15078,N_15159);
nor U15322 (N_15322,N_15003,N_15233);
and U15323 (N_15323,N_15146,N_15034);
and U15324 (N_15324,N_15227,N_15084);
or U15325 (N_15325,N_15172,N_15237);
or U15326 (N_15326,N_15134,N_15186);
nand U15327 (N_15327,N_15208,N_15040);
or U15328 (N_15328,N_15161,N_15075);
nor U15329 (N_15329,N_15243,N_15087);
and U15330 (N_15330,N_15248,N_15041);
nor U15331 (N_15331,N_15073,N_15030);
and U15332 (N_15332,N_15102,N_15123);
and U15333 (N_15333,N_15223,N_15140);
or U15334 (N_15334,N_15174,N_15220);
nor U15335 (N_15335,N_15185,N_15095);
and U15336 (N_15336,N_15118,N_15004);
nor U15337 (N_15337,N_15214,N_15037);
nand U15338 (N_15338,N_15065,N_15189);
and U15339 (N_15339,N_15008,N_15044);
nand U15340 (N_15340,N_15064,N_15160);
and U15341 (N_15341,N_15007,N_15224);
xnor U15342 (N_15342,N_15022,N_15018);
nor U15343 (N_15343,N_15049,N_15222);
and U15344 (N_15344,N_15128,N_15136);
nor U15345 (N_15345,N_15149,N_15106);
and U15346 (N_15346,N_15125,N_15150);
and U15347 (N_15347,N_15051,N_15098);
xor U15348 (N_15348,N_15235,N_15045);
nand U15349 (N_15349,N_15033,N_15060);
xnor U15350 (N_15350,N_15080,N_15025);
and U15351 (N_15351,N_15048,N_15247);
or U15352 (N_15352,N_15056,N_15155);
and U15353 (N_15353,N_15122,N_15132);
or U15354 (N_15354,N_15023,N_15101);
or U15355 (N_15355,N_15230,N_15236);
nor U15356 (N_15356,N_15097,N_15109);
or U15357 (N_15357,N_15091,N_15138);
or U15358 (N_15358,N_15043,N_15187);
nor U15359 (N_15359,N_15031,N_15240);
nand U15360 (N_15360,N_15077,N_15205);
nor U15361 (N_15361,N_15181,N_15145);
nand U15362 (N_15362,N_15070,N_15124);
and U15363 (N_15363,N_15100,N_15148);
nand U15364 (N_15364,N_15089,N_15184);
xor U15365 (N_15365,N_15103,N_15082);
nand U15366 (N_15366,N_15062,N_15192);
or U15367 (N_15367,N_15052,N_15074);
or U15368 (N_15368,N_15191,N_15226);
and U15369 (N_15369,N_15068,N_15156);
nand U15370 (N_15370,N_15085,N_15170);
or U15371 (N_15371,N_15218,N_15081);
nand U15372 (N_15372,N_15092,N_15203);
and U15373 (N_15373,N_15113,N_15232);
or U15374 (N_15374,N_15039,N_15029);
and U15375 (N_15375,N_15034,N_15028);
or U15376 (N_15376,N_15191,N_15083);
nand U15377 (N_15377,N_15024,N_15090);
nor U15378 (N_15378,N_15028,N_15105);
nor U15379 (N_15379,N_15121,N_15235);
xor U15380 (N_15380,N_15039,N_15151);
or U15381 (N_15381,N_15113,N_15207);
nor U15382 (N_15382,N_15202,N_15109);
xnor U15383 (N_15383,N_15032,N_15064);
nand U15384 (N_15384,N_15151,N_15236);
and U15385 (N_15385,N_15160,N_15040);
and U15386 (N_15386,N_15000,N_15222);
and U15387 (N_15387,N_15227,N_15222);
nand U15388 (N_15388,N_15063,N_15101);
xnor U15389 (N_15389,N_15240,N_15170);
and U15390 (N_15390,N_15028,N_15158);
nand U15391 (N_15391,N_15038,N_15210);
nor U15392 (N_15392,N_15019,N_15138);
nand U15393 (N_15393,N_15195,N_15097);
and U15394 (N_15394,N_15091,N_15177);
nor U15395 (N_15395,N_15148,N_15082);
nand U15396 (N_15396,N_15118,N_15119);
nor U15397 (N_15397,N_15092,N_15064);
nor U15398 (N_15398,N_15019,N_15163);
and U15399 (N_15399,N_15201,N_15195);
or U15400 (N_15400,N_15149,N_15016);
xor U15401 (N_15401,N_15058,N_15232);
and U15402 (N_15402,N_15183,N_15249);
and U15403 (N_15403,N_15079,N_15102);
or U15404 (N_15404,N_15211,N_15174);
and U15405 (N_15405,N_15249,N_15205);
nand U15406 (N_15406,N_15040,N_15235);
xor U15407 (N_15407,N_15099,N_15200);
and U15408 (N_15408,N_15039,N_15208);
nor U15409 (N_15409,N_15072,N_15050);
nand U15410 (N_15410,N_15126,N_15172);
xnor U15411 (N_15411,N_15137,N_15035);
and U15412 (N_15412,N_15200,N_15120);
and U15413 (N_15413,N_15100,N_15230);
or U15414 (N_15414,N_15179,N_15024);
nor U15415 (N_15415,N_15077,N_15131);
and U15416 (N_15416,N_15249,N_15207);
xor U15417 (N_15417,N_15209,N_15082);
nor U15418 (N_15418,N_15121,N_15028);
nand U15419 (N_15419,N_15125,N_15065);
and U15420 (N_15420,N_15145,N_15237);
or U15421 (N_15421,N_15107,N_15223);
nand U15422 (N_15422,N_15243,N_15189);
and U15423 (N_15423,N_15200,N_15017);
or U15424 (N_15424,N_15083,N_15127);
nor U15425 (N_15425,N_15201,N_15129);
or U15426 (N_15426,N_15108,N_15099);
and U15427 (N_15427,N_15189,N_15163);
nand U15428 (N_15428,N_15079,N_15013);
or U15429 (N_15429,N_15082,N_15139);
or U15430 (N_15430,N_15198,N_15112);
and U15431 (N_15431,N_15219,N_15166);
or U15432 (N_15432,N_15100,N_15241);
nor U15433 (N_15433,N_15221,N_15220);
or U15434 (N_15434,N_15053,N_15130);
xnor U15435 (N_15435,N_15164,N_15004);
or U15436 (N_15436,N_15059,N_15146);
nor U15437 (N_15437,N_15236,N_15004);
or U15438 (N_15438,N_15143,N_15103);
xor U15439 (N_15439,N_15181,N_15020);
nor U15440 (N_15440,N_15245,N_15152);
nor U15441 (N_15441,N_15026,N_15001);
or U15442 (N_15442,N_15081,N_15085);
xnor U15443 (N_15443,N_15218,N_15060);
or U15444 (N_15444,N_15155,N_15082);
and U15445 (N_15445,N_15179,N_15226);
or U15446 (N_15446,N_15098,N_15213);
nand U15447 (N_15447,N_15124,N_15189);
nor U15448 (N_15448,N_15126,N_15038);
or U15449 (N_15449,N_15116,N_15174);
nand U15450 (N_15450,N_15053,N_15059);
or U15451 (N_15451,N_15194,N_15093);
nand U15452 (N_15452,N_15193,N_15134);
nand U15453 (N_15453,N_15160,N_15124);
and U15454 (N_15454,N_15244,N_15014);
or U15455 (N_15455,N_15109,N_15198);
nor U15456 (N_15456,N_15228,N_15018);
and U15457 (N_15457,N_15112,N_15126);
or U15458 (N_15458,N_15069,N_15092);
xnor U15459 (N_15459,N_15149,N_15165);
and U15460 (N_15460,N_15077,N_15031);
nor U15461 (N_15461,N_15029,N_15136);
nor U15462 (N_15462,N_15124,N_15045);
nor U15463 (N_15463,N_15099,N_15019);
nor U15464 (N_15464,N_15043,N_15205);
or U15465 (N_15465,N_15113,N_15189);
and U15466 (N_15466,N_15234,N_15014);
nor U15467 (N_15467,N_15070,N_15206);
nor U15468 (N_15468,N_15210,N_15002);
or U15469 (N_15469,N_15175,N_15085);
xor U15470 (N_15470,N_15207,N_15046);
nand U15471 (N_15471,N_15017,N_15113);
xnor U15472 (N_15472,N_15047,N_15073);
and U15473 (N_15473,N_15153,N_15203);
nand U15474 (N_15474,N_15168,N_15116);
nand U15475 (N_15475,N_15172,N_15122);
and U15476 (N_15476,N_15185,N_15218);
nor U15477 (N_15477,N_15239,N_15130);
nand U15478 (N_15478,N_15122,N_15144);
nand U15479 (N_15479,N_15103,N_15232);
or U15480 (N_15480,N_15132,N_15063);
nand U15481 (N_15481,N_15011,N_15165);
nor U15482 (N_15482,N_15138,N_15217);
nor U15483 (N_15483,N_15040,N_15162);
nand U15484 (N_15484,N_15033,N_15100);
nand U15485 (N_15485,N_15118,N_15165);
nor U15486 (N_15486,N_15183,N_15052);
nand U15487 (N_15487,N_15155,N_15080);
or U15488 (N_15488,N_15097,N_15171);
nand U15489 (N_15489,N_15191,N_15091);
nand U15490 (N_15490,N_15181,N_15168);
and U15491 (N_15491,N_15161,N_15089);
xor U15492 (N_15492,N_15232,N_15107);
or U15493 (N_15493,N_15235,N_15144);
or U15494 (N_15494,N_15028,N_15249);
and U15495 (N_15495,N_15076,N_15146);
nor U15496 (N_15496,N_15164,N_15230);
nor U15497 (N_15497,N_15173,N_15248);
nand U15498 (N_15498,N_15099,N_15158);
nor U15499 (N_15499,N_15027,N_15194);
and U15500 (N_15500,N_15276,N_15329);
nor U15501 (N_15501,N_15326,N_15307);
or U15502 (N_15502,N_15366,N_15297);
or U15503 (N_15503,N_15474,N_15430);
and U15504 (N_15504,N_15396,N_15417);
nor U15505 (N_15505,N_15360,N_15389);
nor U15506 (N_15506,N_15291,N_15495);
nor U15507 (N_15507,N_15472,N_15385);
nand U15508 (N_15508,N_15344,N_15295);
xor U15509 (N_15509,N_15395,N_15491);
nor U15510 (N_15510,N_15321,N_15447);
nor U15511 (N_15511,N_15342,N_15299);
nor U15512 (N_15512,N_15282,N_15384);
nor U15513 (N_15513,N_15328,N_15335);
or U15514 (N_15514,N_15442,N_15457);
nor U15515 (N_15515,N_15313,N_15273);
nand U15516 (N_15516,N_15425,N_15353);
and U15517 (N_15517,N_15399,N_15306);
nand U15518 (N_15518,N_15263,N_15439);
or U15519 (N_15519,N_15316,N_15429);
and U15520 (N_15520,N_15293,N_15484);
nor U15521 (N_15521,N_15289,N_15435);
and U15522 (N_15522,N_15304,N_15317);
nor U15523 (N_15523,N_15336,N_15437);
or U15524 (N_15524,N_15333,N_15287);
nor U15525 (N_15525,N_15413,N_15266);
nand U15526 (N_15526,N_15422,N_15372);
nor U15527 (N_15527,N_15378,N_15332);
or U15528 (N_15528,N_15477,N_15486);
nand U15529 (N_15529,N_15368,N_15462);
or U15530 (N_15530,N_15444,N_15479);
nor U15531 (N_15531,N_15402,N_15432);
nand U15532 (N_15532,N_15408,N_15351);
or U15533 (N_15533,N_15339,N_15473);
and U15534 (N_15534,N_15460,N_15356);
nand U15535 (N_15535,N_15456,N_15301);
or U15536 (N_15536,N_15449,N_15303);
or U15537 (N_15537,N_15373,N_15364);
nor U15538 (N_15538,N_15250,N_15265);
or U15539 (N_15539,N_15355,N_15327);
and U15540 (N_15540,N_15397,N_15374);
nand U15541 (N_15541,N_15275,N_15280);
or U15542 (N_15542,N_15443,N_15390);
nor U15543 (N_15543,N_15255,N_15369);
and U15544 (N_15544,N_15286,N_15466);
and U15545 (N_15545,N_15464,N_15322);
or U15546 (N_15546,N_15404,N_15296);
and U15547 (N_15547,N_15411,N_15285);
or U15548 (N_15548,N_15278,N_15310);
or U15549 (N_15549,N_15434,N_15259);
nor U15550 (N_15550,N_15488,N_15423);
nand U15551 (N_15551,N_15338,N_15309);
nand U15552 (N_15552,N_15468,N_15334);
nand U15553 (N_15553,N_15412,N_15270);
nand U15554 (N_15554,N_15382,N_15256);
xnor U15555 (N_15555,N_15451,N_15331);
nand U15556 (N_15556,N_15314,N_15469);
and U15557 (N_15557,N_15290,N_15325);
or U15558 (N_15558,N_15380,N_15418);
nand U15559 (N_15559,N_15386,N_15489);
and U15560 (N_15560,N_15281,N_15337);
nor U15561 (N_15561,N_15267,N_15420);
or U15562 (N_15562,N_15414,N_15377);
and U15563 (N_15563,N_15343,N_15375);
nand U15564 (N_15564,N_15305,N_15323);
nor U15565 (N_15565,N_15478,N_15379);
or U15566 (N_15566,N_15340,N_15401);
nor U15567 (N_15567,N_15403,N_15485);
xnor U15568 (N_15568,N_15268,N_15279);
and U15569 (N_15569,N_15312,N_15405);
xnor U15570 (N_15570,N_15454,N_15357);
and U15571 (N_15571,N_15352,N_15490);
or U15572 (N_15572,N_15450,N_15427);
nand U15573 (N_15573,N_15440,N_15428);
or U15574 (N_15574,N_15480,N_15387);
xor U15575 (N_15575,N_15453,N_15358);
xor U15576 (N_15576,N_15493,N_15363);
xnor U15577 (N_15577,N_15251,N_15496);
nor U15578 (N_15578,N_15475,N_15349);
nand U15579 (N_15579,N_15371,N_15407);
nor U15580 (N_15580,N_15283,N_15367);
nor U15581 (N_15581,N_15274,N_15436);
nor U15582 (N_15582,N_15406,N_15277);
or U15583 (N_15583,N_15459,N_15361);
and U15584 (N_15584,N_15497,N_15467);
nor U15585 (N_15585,N_15398,N_15448);
nand U15586 (N_15586,N_15257,N_15320);
nand U15587 (N_15587,N_15264,N_15260);
xor U15588 (N_15588,N_15292,N_15254);
nor U15589 (N_15589,N_15300,N_15471);
nand U15590 (N_15590,N_15308,N_15483);
xnor U15591 (N_15591,N_15492,N_15341);
nand U15592 (N_15592,N_15481,N_15394);
and U15593 (N_15593,N_15381,N_15476);
nor U15594 (N_15594,N_15391,N_15271);
nand U15595 (N_15595,N_15383,N_15294);
and U15596 (N_15596,N_15470,N_15359);
and U15597 (N_15597,N_15494,N_15269);
or U15598 (N_15598,N_15347,N_15419);
and U15599 (N_15599,N_15272,N_15258);
nand U15600 (N_15600,N_15298,N_15441);
and U15601 (N_15601,N_15350,N_15487);
or U15602 (N_15602,N_15288,N_15446);
nor U15603 (N_15603,N_15424,N_15253);
xor U15604 (N_15604,N_15431,N_15410);
nand U15605 (N_15605,N_15455,N_15499);
nor U15606 (N_15606,N_15330,N_15302);
and U15607 (N_15607,N_15376,N_15482);
and U15608 (N_15608,N_15348,N_15262);
or U15609 (N_15609,N_15370,N_15426);
or U15610 (N_15610,N_15452,N_15392);
nand U15611 (N_15611,N_15445,N_15393);
nand U15612 (N_15612,N_15463,N_15438);
nor U15613 (N_15613,N_15409,N_15388);
and U15614 (N_15614,N_15458,N_15324);
and U15615 (N_15615,N_15315,N_15415);
nand U15616 (N_15616,N_15400,N_15261);
or U15617 (N_15617,N_15318,N_15354);
nand U15618 (N_15618,N_15498,N_15319);
nand U15619 (N_15619,N_15362,N_15365);
nand U15620 (N_15620,N_15461,N_15346);
or U15621 (N_15621,N_15416,N_15345);
nand U15622 (N_15622,N_15465,N_15433);
nand U15623 (N_15623,N_15421,N_15311);
nand U15624 (N_15624,N_15284,N_15252);
and U15625 (N_15625,N_15302,N_15335);
nand U15626 (N_15626,N_15350,N_15386);
or U15627 (N_15627,N_15273,N_15260);
and U15628 (N_15628,N_15251,N_15367);
nand U15629 (N_15629,N_15314,N_15490);
or U15630 (N_15630,N_15312,N_15401);
and U15631 (N_15631,N_15290,N_15450);
nor U15632 (N_15632,N_15267,N_15332);
nand U15633 (N_15633,N_15340,N_15416);
nand U15634 (N_15634,N_15450,N_15261);
nand U15635 (N_15635,N_15269,N_15293);
nand U15636 (N_15636,N_15425,N_15398);
and U15637 (N_15637,N_15497,N_15256);
and U15638 (N_15638,N_15392,N_15323);
or U15639 (N_15639,N_15273,N_15410);
or U15640 (N_15640,N_15325,N_15316);
nor U15641 (N_15641,N_15385,N_15473);
nor U15642 (N_15642,N_15327,N_15252);
or U15643 (N_15643,N_15256,N_15337);
and U15644 (N_15644,N_15459,N_15348);
xor U15645 (N_15645,N_15375,N_15294);
or U15646 (N_15646,N_15293,N_15445);
and U15647 (N_15647,N_15275,N_15300);
and U15648 (N_15648,N_15394,N_15355);
or U15649 (N_15649,N_15279,N_15344);
xnor U15650 (N_15650,N_15302,N_15498);
nand U15651 (N_15651,N_15257,N_15362);
nor U15652 (N_15652,N_15481,N_15427);
nand U15653 (N_15653,N_15287,N_15438);
nor U15654 (N_15654,N_15424,N_15266);
xnor U15655 (N_15655,N_15339,N_15464);
nor U15656 (N_15656,N_15372,N_15387);
and U15657 (N_15657,N_15329,N_15439);
nor U15658 (N_15658,N_15350,N_15367);
and U15659 (N_15659,N_15410,N_15289);
and U15660 (N_15660,N_15438,N_15335);
or U15661 (N_15661,N_15338,N_15423);
or U15662 (N_15662,N_15365,N_15350);
nor U15663 (N_15663,N_15478,N_15488);
nand U15664 (N_15664,N_15464,N_15460);
or U15665 (N_15665,N_15332,N_15255);
nor U15666 (N_15666,N_15335,N_15414);
nand U15667 (N_15667,N_15305,N_15285);
nand U15668 (N_15668,N_15391,N_15406);
nand U15669 (N_15669,N_15351,N_15365);
nor U15670 (N_15670,N_15277,N_15261);
nor U15671 (N_15671,N_15281,N_15262);
nor U15672 (N_15672,N_15294,N_15398);
and U15673 (N_15673,N_15442,N_15438);
nand U15674 (N_15674,N_15382,N_15283);
and U15675 (N_15675,N_15335,N_15405);
nor U15676 (N_15676,N_15268,N_15479);
xor U15677 (N_15677,N_15417,N_15268);
or U15678 (N_15678,N_15290,N_15405);
xnor U15679 (N_15679,N_15301,N_15310);
xnor U15680 (N_15680,N_15471,N_15493);
or U15681 (N_15681,N_15429,N_15397);
and U15682 (N_15682,N_15389,N_15301);
or U15683 (N_15683,N_15462,N_15391);
or U15684 (N_15684,N_15375,N_15300);
nor U15685 (N_15685,N_15437,N_15292);
and U15686 (N_15686,N_15414,N_15477);
or U15687 (N_15687,N_15440,N_15492);
and U15688 (N_15688,N_15412,N_15438);
and U15689 (N_15689,N_15255,N_15443);
xnor U15690 (N_15690,N_15455,N_15434);
xor U15691 (N_15691,N_15371,N_15280);
nor U15692 (N_15692,N_15493,N_15312);
or U15693 (N_15693,N_15395,N_15460);
or U15694 (N_15694,N_15350,N_15274);
nand U15695 (N_15695,N_15269,N_15449);
or U15696 (N_15696,N_15319,N_15367);
and U15697 (N_15697,N_15402,N_15332);
xnor U15698 (N_15698,N_15401,N_15369);
nand U15699 (N_15699,N_15480,N_15311);
or U15700 (N_15700,N_15431,N_15335);
and U15701 (N_15701,N_15432,N_15311);
nor U15702 (N_15702,N_15267,N_15341);
and U15703 (N_15703,N_15396,N_15405);
xor U15704 (N_15704,N_15265,N_15478);
xor U15705 (N_15705,N_15424,N_15419);
nor U15706 (N_15706,N_15319,N_15467);
nor U15707 (N_15707,N_15426,N_15333);
and U15708 (N_15708,N_15265,N_15281);
nand U15709 (N_15709,N_15289,N_15252);
nand U15710 (N_15710,N_15282,N_15394);
nand U15711 (N_15711,N_15451,N_15414);
nand U15712 (N_15712,N_15426,N_15334);
xor U15713 (N_15713,N_15252,N_15377);
nand U15714 (N_15714,N_15389,N_15289);
nor U15715 (N_15715,N_15317,N_15474);
and U15716 (N_15716,N_15467,N_15365);
or U15717 (N_15717,N_15379,N_15306);
or U15718 (N_15718,N_15268,N_15272);
nor U15719 (N_15719,N_15391,N_15356);
or U15720 (N_15720,N_15405,N_15442);
nand U15721 (N_15721,N_15345,N_15311);
nand U15722 (N_15722,N_15333,N_15498);
and U15723 (N_15723,N_15367,N_15420);
xnor U15724 (N_15724,N_15446,N_15407);
and U15725 (N_15725,N_15479,N_15497);
nand U15726 (N_15726,N_15257,N_15392);
or U15727 (N_15727,N_15297,N_15417);
nor U15728 (N_15728,N_15413,N_15327);
or U15729 (N_15729,N_15397,N_15489);
nand U15730 (N_15730,N_15264,N_15423);
or U15731 (N_15731,N_15498,N_15306);
nand U15732 (N_15732,N_15317,N_15406);
nor U15733 (N_15733,N_15327,N_15254);
xnor U15734 (N_15734,N_15291,N_15399);
or U15735 (N_15735,N_15341,N_15398);
nor U15736 (N_15736,N_15357,N_15494);
and U15737 (N_15737,N_15395,N_15366);
nor U15738 (N_15738,N_15388,N_15446);
nor U15739 (N_15739,N_15273,N_15360);
nor U15740 (N_15740,N_15360,N_15495);
or U15741 (N_15741,N_15255,N_15415);
nor U15742 (N_15742,N_15409,N_15444);
and U15743 (N_15743,N_15301,N_15324);
xnor U15744 (N_15744,N_15300,N_15462);
or U15745 (N_15745,N_15395,N_15271);
nor U15746 (N_15746,N_15465,N_15436);
and U15747 (N_15747,N_15337,N_15437);
nand U15748 (N_15748,N_15429,N_15445);
xor U15749 (N_15749,N_15262,N_15445);
or U15750 (N_15750,N_15655,N_15504);
nor U15751 (N_15751,N_15622,N_15533);
nand U15752 (N_15752,N_15551,N_15539);
and U15753 (N_15753,N_15574,N_15611);
and U15754 (N_15754,N_15594,N_15575);
nor U15755 (N_15755,N_15693,N_15708);
nand U15756 (N_15756,N_15546,N_15564);
xor U15757 (N_15757,N_15627,N_15563);
and U15758 (N_15758,N_15542,N_15628);
nand U15759 (N_15759,N_15745,N_15608);
nor U15760 (N_15760,N_15601,N_15560);
nor U15761 (N_15761,N_15573,N_15713);
xnor U15762 (N_15762,N_15570,N_15537);
nand U15763 (N_15763,N_15653,N_15636);
nor U15764 (N_15764,N_15562,N_15721);
nand U15765 (N_15765,N_15508,N_15675);
or U15766 (N_15766,N_15672,N_15669);
or U15767 (N_15767,N_15589,N_15722);
and U15768 (N_15768,N_15707,N_15626);
xor U15769 (N_15769,N_15614,N_15699);
nor U15770 (N_15770,N_15686,N_15748);
nor U15771 (N_15771,N_15746,N_15665);
nor U15772 (N_15772,N_15531,N_15730);
nor U15773 (N_15773,N_15616,N_15631);
xor U15774 (N_15774,N_15676,N_15577);
nor U15775 (N_15775,N_15662,N_15618);
nand U15776 (N_15776,N_15650,N_15732);
nor U15777 (N_15777,N_15599,N_15718);
and U15778 (N_15778,N_15603,N_15696);
and U15779 (N_15779,N_15617,N_15625);
and U15780 (N_15780,N_15717,N_15526);
or U15781 (N_15781,N_15744,N_15540);
or U15782 (N_15782,N_15667,N_15641);
and U15783 (N_15783,N_15691,N_15595);
and U15784 (N_15784,N_15630,N_15688);
or U15785 (N_15785,N_15685,N_15710);
nand U15786 (N_15786,N_15511,N_15668);
and U15787 (N_15787,N_15505,N_15644);
and U15788 (N_15788,N_15525,N_15552);
and U15789 (N_15789,N_15687,N_15606);
nand U15790 (N_15790,N_15523,N_15532);
and U15791 (N_15791,N_15649,N_15637);
or U15792 (N_15792,N_15666,N_15547);
xnor U15793 (N_15793,N_15664,N_15646);
and U15794 (N_15794,N_15576,N_15731);
nor U15795 (N_15795,N_15583,N_15528);
or U15796 (N_15796,N_15638,N_15677);
nor U15797 (N_15797,N_15507,N_15682);
or U15798 (N_15798,N_15600,N_15648);
or U15799 (N_15799,N_15612,N_15538);
or U15800 (N_15800,N_15736,N_15561);
and U15801 (N_15801,N_15515,N_15679);
nand U15802 (N_15802,N_15520,N_15705);
and U15803 (N_15803,N_15527,N_15517);
nand U15804 (N_15804,N_15529,N_15720);
nor U15805 (N_15805,N_15697,N_15536);
nand U15806 (N_15806,N_15654,N_15739);
nand U15807 (N_15807,N_15579,N_15559);
and U15808 (N_15808,N_15738,N_15500);
nand U15809 (N_15809,N_15639,N_15543);
nor U15810 (N_15810,N_15545,N_15632);
nor U15811 (N_15811,N_15597,N_15554);
xnor U15812 (N_15812,N_15728,N_15714);
xnor U15813 (N_15813,N_15716,N_15521);
or U15814 (N_15814,N_15590,N_15660);
and U15815 (N_15815,N_15541,N_15678);
nand U15816 (N_15816,N_15510,N_15742);
and U15817 (N_15817,N_15689,N_15535);
or U15818 (N_15818,N_15733,N_15629);
nand U15819 (N_15819,N_15723,N_15702);
or U15820 (N_15820,N_15503,N_15591);
or U15821 (N_15821,N_15567,N_15613);
or U15822 (N_15822,N_15727,N_15555);
nor U15823 (N_15823,N_15624,N_15619);
and U15824 (N_15824,N_15719,N_15700);
nand U15825 (N_15825,N_15524,N_15509);
nand U15826 (N_15826,N_15704,N_15661);
nor U15827 (N_15827,N_15725,N_15605);
and U15828 (N_15828,N_15544,N_15569);
nand U15829 (N_15829,N_15580,N_15729);
or U15830 (N_15830,N_15530,N_15749);
or U15831 (N_15831,N_15706,N_15610);
nand U15832 (N_15832,N_15651,N_15645);
nor U15833 (N_15833,N_15703,N_15587);
or U15834 (N_15834,N_15514,N_15596);
nand U15835 (N_15835,N_15516,N_15643);
nor U15836 (N_15836,N_15673,N_15747);
and U15837 (N_15837,N_15598,N_15534);
nand U15838 (N_15838,N_15620,N_15657);
or U15839 (N_15839,N_15671,N_15726);
nand U15840 (N_15840,N_15711,N_15680);
and U15841 (N_15841,N_15585,N_15647);
and U15842 (N_15842,N_15522,N_15656);
and U15843 (N_15843,N_15690,N_15615);
nand U15844 (N_15844,N_15588,N_15735);
or U15845 (N_15845,N_15642,N_15556);
nor U15846 (N_15846,N_15586,N_15506);
nor U15847 (N_15847,N_15681,N_15501);
or U15848 (N_15848,N_15712,N_15715);
or U15849 (N_15849,N_15578,N_15633);
or U15850 (N_15850,N_15695,N_15584);
or U15851 (N_15851,N_15621,N_15652);
or U15852 (N_15852,N_15568,N_15694);
or U15853 (N_15853,N_15684,N_15698);
or U15854 (N_15854,N_15549,N_15674);
nor U15855 (N_15855,N_15592,N_15607);
nor U15856 (N_15856,N_15623,N_15692);
xor U15857 (N_15857,N_15659,N_15737);
and U15858 (N_15858,N_15743,N_15558);
or U15859 (N_15859,N_15565,N_15553);
nand U15860 (N_15860,N_15709,N_15740);
nor U15861 (N_15861,N_15502,N_15593);
xnor U15862 (N_15862,N_15566,N_15512);
and U15863 (N_15863,N_15635,N_15683);
xor U15864 (N_15864,N_15604,N_15581);
and U15865 (N_15865,N_15548,N_15701);
or U15866 (N_15866,N_15550,N_15513);
and U15867 (N_15867,N_15582,N_15609);
or U15868 (N_15868,N_15557,N_15663);
and U15869 (N_15869,N_15724,N_15741);
nand U15870 (N_15870,N_15571,N_15640);
nand U15871 (N_15871,N_15658,N_15634);
and U15872 (N_15872,N_15518,N_15734);
xnor U15873 (N_15873,N_15602,N_15519);
and U15874 (N_15874,N_15572,N_15670);
nand U15875 (N_15875,N_15606,N_15724);
and U15876 (N_15876,N_15696,N_15517);
xnor U15877 (N_15877,N_15515,N_15578);
or U15878 (N_15878,N_15711,N_15587);
and U15879 (N_15879,N_15624,N_15661);
and U15880 (N_15880,N_15695,N_15551);
and U15881 (N_15881,N_15504,N_15520);
and U15882 (N_15882,N_15654,N_15581);
and U15883 (N_15883,N_15717,N_15517);
nand U15884 (N_15884,N_15570,N_15708);
nor U15885 (N_15885,N_15749,N_15549);
nand U15886 (N_15886,N_15676,N_15520);
and U15887 (N_15887,N_15646,N_15726);
and U15888 (N_15888,N_15516,N_15553);
nor U15889 (N_15889,N_15522,N_15570);
or U15890 (N_15890,N_15546,N_15502);
and U15891 (N_15891,N_15706,N_15737);
or U15892 (N_15892,N_15504,N_15581);
or U15893 (N_15893,N_15528,N_15712);
nand U15894 (N_15894,N_15676,N_15594);
nand U15895 (N_15895,N_15529,N_15664);
and U15896 (N_15896,N_15623,N_15535);
nor U15897 (N_15897,N_15569,N_15723);
or U15898 (N_15898,N_15705,N_15503);
xor U15899 (N_15899,N_15545,N_15671);
or U15900 (N_15900,N_15542,N_15605);
nor U15901 (N_15901,N_15722,N_15686);
and U15902 (N_15902,N_15733,N_15608);
nor U15903 (N_15903,N_15618,N_15671);
nor U15904 (N_15904,N_15600,N_15711);
nand U15905 (N_15905,N_15717,N_15552);
or U15906 (N_15906,N_15643,N_15656);
or U15907 (N_15907,N_15673,N_15560);
and U15908 (N_15908,N_15629,N_15559);
and U15909 (N_15909,N_15695,N_15717);
or U15910 (N_15910,N_15712,N_15512);
nand U15911 (N_15911,N_15692,N_15578);
nor U15912 (N_15912,N_15704,N_15588);
and U15913 (N_15913,N_15652,N_15622);
or U15914 (N_15914,N_15509,N_15646);
or U15915 (N_15915,N_15506,N_15717);
or U15916 (N_15916,N_15549,N_15733);
and U15917 (N_15917,N_15588,N_15652);
nor U15918 (N_15918,N_15673,N_15705);
nand U15919 (N_15919,N_15567,N_15576);
xnor U15920 (N_15920,N_15657,N_15580);
xnor U15921 (N_15921,N_15730,N_15737);
nand U15922 (N_15922,N_15729,N_15657);
and U15923 (N_15923,N_15747,N_15744);
and U15924 (N_15924,N_15518,N_15730);
or U15925 (N_15925,N_15516,N_15505);
and U15926 (N_15926,N_15728,N_15545);
nor U15927 (N_15927,N_15728,N_15589);
nand U15928 (N_15928,N_15579,N_15740);
and U15929 (N_15929,N_15544,N_15591);
nand U15930 (N_15930,N_15545,N_15524);
nor U15931 (N_15931,N_15585,N_15683);
nand U15932 (N_15932,N_15742,N_15620);
xor U15933 (N_15933,N_15553,N_15578);
nand U15934 (N_15934,N_15638,N_15659);
nor U15935 (N_15935,N_15742,N_15671);
nand U15936 (N_15936,N_15677,N_15724);
or U15937 (N_15937,N_15528,N_15552);
nand U15938 (N_15938,N_15707,N_15533);
or U15939 (N_15939,N_15594,N_15532);
nand U15940 (N_15940,N_15707,N_15615);
or U15941 (N_15941,N_15592,N_15613);
or U15942 (N_15942,N_15548,N_15507);
xor U15943 (N_15943,N_15748,N_15692);
or U15944 (N_15944,N_15738,N_15637);
nor U15945 (N_15945,N_15701,N_15727);
and U15946 (N_15946,N_15599,N_15700);
and U15947 (N_15947,N_15510,N_15745);
and U15948 (N_15948,N_15717,N_15612);
nor U15949 (N_15949,N_15635,N_15634);
nand U15950 (N_15950,N_15709,N_15606);
nor U15951 (N_15951,N_15622,N_15714);
or U15952 (N_15952,N_15633,N_15550);
nand U15953 (N_15953,N_15720,N_15585);
nor U15954 (N_15954,N_15605,N_15598);
nor U15955 (N_15955,N_15624,N_15709);
nor U15956 (N_15956,N_15656,N_15680);
nor U15957 (N_15957,N_15670,N_15518);
and U15958 (N_15958,N_15629,N_15511);
nor U15959 (N_15959,N_15662,N_15573);
or U15960 (N_15960,N_15732,N_15713);
xor U15961 (N_15961,N_15706,N_15509);
nand U15962 (N_15962,N_15602,N_15533);
and U15963 (N_15963,N_15603,N_15507);
and U15964 (N_15964,N_15530,N_15557);
or U15965 (N_15965,N_15582,N_15620);
nand U15966 (N_15966,N_15635,N_15656);
nand U15967 (N_15967,N_15748,N_15644);
xnor U15968 (N_15968,N_15672,N_15697);
or U15969 (N_15969,N_15668,N_15529);
nor U15970 (N_15970,N_15654,N_15593);
nand U15971 (N_15971,N_15592,N_15683);
nor U15972 (N_15972,N_15637,N_15583);
nand U15973 (N_15973,N_15561,N_15748);
and U15974 (N_15974,N_15668,N_15677);
and U15975 (N_15975,N_15590,N_15541);
nand U15976 (N_15976,N_15563,N_15574);
and U15977 (N_15977,N_15632,N_15532);
and U15978 (N_15978,N_15732,N_15579);
nor U15979 (N_15979,N_15542,N_15521);
nor U15980 (N_15980,N_15575,N_15694);
and U15981 (N_15981,N_15537,N_15530);
nand U15982 (N_15982,N_15652,N_15568);
nand U15983 (N_15983,N_15679,N_15675);
nor U15984 (N_15984,N_15673,N_15520);
nor U15985 (N_15985,N_15719,N_15735);
nor U15986 (N_15986,N_15576,N_15577);
nor U15987 (N_15987,N_15503,N_15644);
or U15988 (N_15988,N_15595,N_15677);
nor U15989 (N_15989,N_15570,N_15702);
or U15990 (N_15990,N_15580,N_15721);
nor U15991 (N_15991,N_15574,N_15653);
nor U15992 (N_15992,N_15519,N_15727);
or U15993 (N_15993,N_15686,N_15647);
nand U15994 (N_15994,N_15580,N_15510);
and U15995 (N_15995,N_15590,N_15676);
nand U15996 (N_15996,N_15631,N_15706);
xor U15997 (N_15997,N_15590,N_15539);
or U15998 (N_15998,N_15611,N_15669);
or U15999 (N_15999,N_15691,N_15580);
and U16000 (N_16000,N_15779,N_15861);
or U16001 (N_16001,N_15798,N_15990);
nor U16002 (N_16002,N_15936,N_15966);
xor U16003 (N_16003,N_15805,N_15882);
or U16004 (N_16004,N_15840,N_15775);
or U16005 (N_16005,N_15785,N_15995);
xnor U16006 (N_16006,N_15915,N_15946);
nor U16007 (N_16007,N_15949,N_15884);
nand U16008 (N_16008,N_15802,N_15807);
or U16009 (N_16009,N_15824,N_15985);
or U16010 (N_16010,N_15790,N_15832);
and U16011 (N_16011,N_15846,N_15976);
nor U16012 (N_16012,N_15797,N_15765);
or U16013 (N_16013,N_15883,N_15770);
xnor U16014 (N_16014,N_15787,N_15784);
or U16015 (N_16015,N_15893,N_15923);
nand U16016 (N_16016,N_15930,N_15842);
nor U16017 (N_16017,N_15828,N_15862);
nor U16018 (N_16018,N_15845,N_15788);
nor U16019 (N_16019,N_15868,N_15947);
nand U16020 (N_16020,N_15937,N_15789);
or U16021 (N_16021,N_15847,N_15863);
xnor U16022 (N_16022,N_15927,N_15953);
and U16023 (N_16023,N_15950,N_15928);
and U16024 (N_16024,N_15815,N_15909);
nand U16025 (N_16025,N_15849,N_15996);
and U16026 (N_16026,N_15929,N_15829);
or U16027 (N_16027,N_15834,N_15892);
xor U16028 (N_16028,N_15757,N_15945);
nand U16029 (N_16029,N_15974,N_15848);
nor U16030 (N_16030,N_15806,N_15877);
nor U16031 (N_16031,N_15766,N_15767);
and U16032 (N_16032,N_15854,N_15837);
xor U16033 (N_16033,N_15955,N_15954);
or U16034 (N_16034,N_15850,N_15869);
nand U16035 (N_16035,N_15980,N_15918);
xor U16036 (N_16036,N_15859,N_15926);
nand U16037 (N_16037,N_15920,N_15763);
nand U16038 (N_16038,N_15856,N_15780);
or U16039 (N_16039,N_15800,N_15759);
nor U16040 (N_16040,N_15777,N_15948);
and U16041 (N_16041,N_15817,N_15857);
or U16042 (N_16042,N_15899,N_15897);
nand U16043 (N_16043,N_15755,N_15890);
xor U16044 (N_16044,N_15917,N_15822);
and U16045 (N_16045,N_15760,N_15752);
nor U16046 (N_16046,N_15879,N_15764);
and U16047 (N_16047,N_15914,N_15997);
and U16048 (N_16048,N_15988,N_15794);
or U16049 (N_16049,N_15870,N_15751);
and U16050 (N_16050,N_15906,N_15811);
nand U16051 (N_16051,N_15992,N_15872);
and U16052 (N_16052,N_15783,N_15762);
or U16053 (N_16053,N_15820,N_15903);
and U16054 (N_16054,N_15907,N_15982);
or U16055 (N_16055,N_15924,N_15981);
or U16056 (N_16056,N_15833,N_15853);
nor U16057 (N_16057,N_15964,N_15812);
or U16058 (N_16058,N_15855,N_15962);
or U16059 (N_16059,N_15801,N_15919);
or U16060 (N_16060,N_15836,N_15968);
and U16061 (N_16061,N_15838,N_15881);
and U16062 (N_16062,N_15852,N_15750);
and U16063 (N_16063,N_15808,N_15971);
or U16064 (N_16064,N_15814,N_15942);
or U16065 (N_16065,N_15804,N_15977);
and U16066 (N_16066,N_15774,N_15809);
or U16067 (N_16067,N_15792,N_15758);
nand U16068 (N_16068,N_15835,N_15894);
or U16069 (N_16069,N_15813,N_15876);
nand U16070 (N_16070,N_15773,N_15944);
nand U16071 (N_16071,N_15819,N_15895);
nor U16072 (N_16072,N_15978,N_15867);
or U16073 (N_16073,N_15796,N_15889);
and U16074 (N_16074,N_15998,N_15943);
xor U16075 (N_16075,N_15756,N_15776);
or U16076 (N_16076,N_15973,N_15984);
xor U16077 (N_16077,N_15791,N_15825);
or U16078 (N_16078,N_15908,N_15873);
nor U16079 (N_16079,N_15858,N_15781);
and U16080 (N_16080,N_15799,N_15898);
nand U16081 (N_16081,N_15951,N_15963);
nor U16082 (N_16082,N_15911,N_15831);
nand U16083 (N_16083,N_15989,N_15778);
nand U16084 (N_16084,N_15933,N_15865);
or U16085 (N_16085,N_15994,N_15826);
nor U16086 (N_16086,N_15782,N_15916);
nor U16087 (N_16087,N_15941,N_15875);
or U16088 (N_16088,N_15761,N_15910);
xor U16089 (N_16089,N_15905,N_15866);
or U16090 (N_16090,N_15880,N_15972);
or U16091 (N_16091,N_15904,N_15754);
xor U16092 (N_16092,N_15816,N_15769);
xor U16093 (N_16093,N_15940,N_15961);
or U16094 (N_16094,N_15969,N_15839);
xor U16095 (N_16095,N_15887,N_15901);
nor U16096 (N_16096,N_15902,N_15925);
or U16097 (N_16097,N_15965,N_15970);
and U16098 (N_16098,N_15772,N_15888);
nand U16099 (N_16099,N_15771,N_15896);
and U16100 (N_16100,N_15932,N_15768);
nand U16101 (N_16101,N_15957,N_15913);
and U16102 (N_16102,N_15939,N_15864);
xor U16103 (N_16103,N_15871,N_15987);
or U16104 (N_16104,N_15986,N_15891);
nor U16105 (N_16105,N_15960,N_15922);
nand U16106 (N_16106,N_15900,N_15860);
or U16107 (N_16107,N_15983,N_15967);
nand U16108 (N_16108,N_15878,N_15958);
and U16109 (N_16109,N_15979,N_15803);
nor U16110 (N_16110,N_15956,N_15843);
nand U16111 (N_16111,N_15934,N_15818);
xnor U16112 (N_16112,N_15975,N_15844);
and U16113 (N_16113,N_15952,N_15821);
or U16114 (N_16114,N_15810,N_15921);
and U16115 (N_16115,N_15959,N_15886);
or U16116 (N_16116,N_15823,N_15793);
or U16117 (N_16117,N_15999,N_15993);
nor U16118 (N_16118,N_15786,N_15991);
and U16119 (N_16119,N_15912,N_15885);
nor U16120 (N_16120,N_15935,N_15874);
or U16121 (N_16121,N_15938,N_15851);
nand U16122 (N_16122,N_15830,N_15841);
nand U16123 (N_16123,N_15931,N_15753);
and U16124 (N_16124,N_15827,N_15795);
and U16125 (N_16125,N_15842,N_15920);
and U16126 (N_16126,N_15796,N_15957);
or U16127 (N_16127,N_15837,N_15760);
nor U16128 (N_16128,N_15971,N_15790);
or U16129 (N_16129,N_15797,N_15796);
or U16130 (N_16130,N_15763,N_15832);
xor U16131 (N_16131,N_15750,N_15764);
or U16132 (N_16132,N_15948,N_15859);
nor U16133 (N_16133,N_15911,N_15799);
nand U16134 (N_16134,N_15934,N_15995);
or U16135 (N_16135,N_15902,N_15875);
nor U16136 (N_16136,N_15974,N_15995);
nand U16137 (N_16137,N_15813,N_15975);
nor U16138 (N_16138,N_15854,N_15881);
or U16139 (N_16139,N_15964,N_15757);
or U16140 (N_16140,N_15879,N_15967);
or U16141 (N_16141,N_15943,N_15894);
xnor U16142 (N_16142,N_15891,N_15923);
xor U16143 (N_16143,N_15797,N_15912);
nand U16144 (N_16144,N_15881,N_15974);
xor U16145 (N_16145,N_15881,N_15953);
and U16146 (N_16146,N_15772,N_15843);
nor U16147 (N_16147,N_15814,N_15848);
or U16148 (N_16148,N_15782,N_15960);
xnor U16149 (N_16149,N_15786,N_15984);
or U16150 (N_16150,N_15864,N_15962);
and U16151 (N_16151,N_15909,N_15964);
and U16152 (N_16152,N_15943,N_15786);
nand U16153 (N_16153,N_15866,N_15904);
nor U16154 (N_16154,N_15900,N_15774);
or U16155 (N_16155,N_15872,N_15753);
and U16156 (N_16156,N_15957,N_15791);
and U16157 (N_16157,N_15823,N_15820);
nand U16158 (N_16158,N_15968,N_15801);
nor U16159 (N_16159,N_15985,N_15945);
xnor U16160 (N_16160,N_15840,N_15809);
nor U16161 (N_16161,N_15810,N_15879);
or U16162 (N_16162,N_15916,N_15994);
nor U16163 (N_16163,N_15925,N_15962);
and U16164 (N_16164,N_15867,N_15944);
or U16165 (N_16165,N_15890,N_15822);
nor U16166 (N_16166,N_15978,N_15895);
nor U16167 (N_16167,N_15771,N_15974);
and U16168 (N_16168,N_15859,N_15782);
and U16169 (N_16169,N_15911,N_15815);
or U16170 (N_16170,N_15996,N_15993);
and U16171 (N_16171,N_15771,N_15965);
nand U16172 (N_16172,N_15785,N_15824);
and U16173 (N_16173,N_15903,N_15860);
nand U16174 (N_16174,N_15795,N_15828);
or U16175 (N_16175,N_15755,N_15914);
nor U16176 (N_16176,N_15750,N_15779);
nor U16177 (N_16177,N_15918,N_15913);
or U16178 (N_16178,N_15984,N_15795);
xnor U16179 (N_16179,N_15902,N_15830);
xor U16180 (N_16180,N_15916,N_15874);
nand U16181 (N_16181,N_15825,N_15974);
and U16182 (N_16182,N_15753,N_15790);
nor U16183 (N_16183,N_15917,N_15936);
nand U16184 (N_16184,N_15926,N_15818);
and U16185 (N_16185,N_15755,N_15879);
or U16186 (N_16186,N_15967,N_15848);
and U16187 (N_16187,N_15902,N_15922);
and U16188 (N_16188,N_15939,N_15917);
or U16189 (N_16189,N_15942,N_15866);
and U16190 (N_16190,N_15870,N_15832);
and U16191 (N_16191,N_15781,N_15832);
nand U16192 (N_16192,N_15923,N_15770);
and U16193 (N_16193,N_15806,N_15959);
or U16194 (N_16194,N_15930,N_15753);
xor U16195 (N_16195,N_15769,N_15758);
and U16196 (N_16196,N_15793,N_15835);
nor U16197 (N_16197,N_15947,N_15927);
or U16198 (N_16198,N_15932,N_15906);
nor U16199 (N_16199,N_15792,N_15769);
and U16200 (N_16200,N_15889,N_15814);
or U16201 (N_16201,N_15884,N_15965);
or U16202 (N_16202,N_15773,N_15862);
nand U16203 (N_16203,N_15885,N_15840);
or U16204 (N_16204,N_15991,N_15763);
and U16205 (N_16205,N_15962,N_15814);
xnor U16206 (N_16206,N_15848,N_15987);
xor U16207 (N_16207,N_15946,N_15864);
nor U16208 (N_16208,N_15853,N_15819);
and U16209 (N_16209,N_15965,N_15756);
or U16210 (N_16210,N_15888,N_15835);
nand U16211 (N_16211,N_15917,N_15762);
nor U16212 (N_16212,N_15791,N_15867);
and U16213 (N_16213,N_15912,N_15881);
nor U16214 (N_16214,N_15945,N_15848);
nand U16215 (N_16215,N_15900,N_15941);
nand U16216 (N_16216,N_15996,N_15966);
or U16217 (N_16217,N_15875,N_15954);
or U16218 (N_16218,N_15952,N_15970);
or U16219 (N_16219,N_15890,N_15807);
nand U16220 (N_16220,N_15963,N_15758);
nand U16221 (N_16221,N_15922,N_15865);
nand U16222 (N_16222,N_15979,N_15774);
nor U16223 (N_16223,N_15877,N_15759);
nor U16224 (N_16224,N_15843,N_15912);
nor U16225 (N_16225,N_15820,N_15766);
nor U16226 (N_16226,N_15803,N_15769);
xnor U16227 (N_16227,N_15799,N_15909);
or U16228 (N_16228,N_15979,N_15923);
or U16229 (N_16229,N_15991,N_15919);
or U16230 (N_16230,N_15838,N_15899);
xnor U16231 (N_16231,N_15951,N_15924);
or U16232 (N_16232,N_15902,N_15872);
xor U16233 (N_16233,N_15966,N_15838);
xnor U16234 (N_16234,N_15841,N_15931);
xor U16235 (N_16235,N_15855,N_15947);
nand U16236 (N_16236,N_15763,N_15986);
xnor U16237 (N_16237,N_15929,N_15758);
or U16238 (N_16238,N_15767,N_15765);
or U16239 (N_16239,N_15898,N_15802);
nor U16240 (N_16240,N_15934,N_15839);
and U16241 (N_16241,N_15837,N_15868);
or U16242 (N_16242,N_15975,N_15875);
and U16243 (N_16243,N_15971,N_15801);
xor U16244 (N_16244,N_15758,N_15917);
nand U16245 (N_16245,N_15754,N_15798);
and U16246 (N_16246,N_15997,N_15754);
xor U16247 (N_16247,N_15898,N_15808);
nand U16248 (N_16248,N_15908,N_15937);
and U16249 (N_16249,N_15927,N_15907);
nor U16250 (N_16250,N_16097,N_16051);
and U16251 (N_16251,N_16092,N_16134);
or U16252 (N_16252,N_16149,N_16129);
or U16253 (N_16253,N_16182,N_16003);
and U16254 (N_16254,N_16185,N_16198);
nor U16255 (N_16255,N_16172,N_16009);
nor U16256 (N_16256,N_16019,N_16024);
nand U16257 (N_16257,N_16152,N_16062);
xnor U16258 (N_16258,N_16156,N_16140);
nand U16259 (N_16259,N_16007,N_16157);
and U16260 (N_16260,N_16099,N_16011);
nor U16261 (N_16261,N_16073,N_16133);
and U16262 (N_16262,N_16096,N_16032);
nand U16263 (N_16263,N_16059,N_16022);
or U16264 (N_16264,N_16033,N_16141);
xor U16265 (N_16265,N_16166,N_16014);
or U16266 (N_16266,N_16178,N_16114);
nor U16267 (N_16267,N_16146,N_16148);
or U16268 (N_16268,N_16091,N_16087);
or U16269 (N_16269,N_16113,N_16176);
nand U16270 (N_16270,N_16162,N_16081);
nor U16271 (N_16271,N_16232,N_16004);
nor U16272 (N_16272,N_16021,N_16023);
nand U16273 (N_16273,N_16168,N_16240);
nor U16274 (N_16274,N_16042,N_16184);
nand U16275 (N_16275,N_16052,N_16135);
nand U16276 (N_16276,N_16050,N_16206);
nand U16277 (N_16277,N_16001,N_16218);
xor U16278 (N_16278,N_16125,N_16196);
and U16279 (N_16279,N_16237,N_16201);
xnor U16280 (N_16280,N_16054,N_16035);
and U16281 (N_16281,N_16199,N_16236);
and U16282 (N_16282,N_16153,N_16057);
and U16283 (N_16283,N_16018,N_16160);
nor U16284 (N_16284,N_16205,N_16034);
and U16285 (N_16285,N_16233,N_16098);
xor U16286 (N_16286,N_16060,N_16038);
nor U16287 (N_16287,N_16090,N_16249);
nand U16288 (N_16288,N_16223,N_16213);
or U16289 (N_16289,N_16025,N_16136);
nor U16290 (N_16290,N_16246,N_16002);
nor U16291 (N_16291,N_16179,N_16226);
or U16292 (N_16292,N_16040,N_16221);
or U16293 (N_16293,N_16143,N_16144);
and U16294 (N_16294,N_16122,N_16008);
and U16295 (N_16295,N_16217,N_16055);
nor U16296 (N_16296,N_16071,N_16006);
nor U16297 (N_16297,N_16147,N_16102);
nand U16298 (N_16298,N_16164,N_16074);
and U16299 (N_16299,N_16077,N_16208);
or U16300 (N_16300,N_16126,N_16078);
or U16301 (N_16301,N_16121,N_16220);
and U16302 (N_16302,N_16186,N_16171);
and U16303 (N_16303,N_16085,N_16242);
nor U16304 (N_16304,N_16244,N_16190);
and U16305 (N_16305,N_16028,N_16193);
xnor U16306 (N_16306,N_16131,N_16120);
nand U16307 (N_16307,N_16159,N_16241);
or U16308 (N_16308,N_16013,N_16031);
nand U16309 (N_16309,N_16111,N_16106);
nor U16310 (N_16310,N_16197,N_16044);
xnor U16311 (N_16311,N_16058,N_16219);
and U16312 (N_16312,N_16247,N_16000);
nand U16313 (N_16313,N_16067,N_16215);
and U16314 (N_16314,N_16089,N_16245);
nor U16315 (N_16315,N_16248,N_16118);
nor U16316 (N_16316,N_16104,N_16175);
and U16317 (N_16317,N_16155,N_16243);
nand U16318 (N_16318,N_16015,N_16211);
or U16319 (N_16319,N_16203,N_16010);
xor U16320 (N_16320,N_16066,N_16026);
and U16321 (N_16321,N_16228,N_16239);
nor U16322 (N_16322,N_16093,N_16229);
or U16323 (N_16323,N_16167,N_16030);
nor U16324 (N_16324,N_16195,N_16139);
nand U16325 (N_16325,N_16072,N_16115);
nor U16326 (N_16326,N_16142,N_16173);
nor U16327 (N_16327,N_16177,N_16174);
and U16328 (N_16328,N_16227,N_16123);
and U16329 (N_16329,N_16235,N_16082);
xnor U16330 (N_16330,N_16047,N_16101);
xnor U16331 (N_16331,N_16225,N_16061);
nor U16332 (N_16332,N_16127,N_16105);
or U16333 (N_16333,N_16154,N_16194);
and U16334 (N_16334,N_16188,N_16036);
nor U16335 (N_16335,N_16180,N_16063);
or U16336 (N_16336,N_16187,N_16016);
nor U16337 (N_16337,N_16224,N_16183);
nor U16338 (N_16338,N_16070,N_16210);
or U16339 (N_16339,N_16017,N_16107);
nand U16340 (N_16340,N_16189,N_16012);
and U16341 (N_16341,N_16238,N_16079);
and U16342 (N_16342,N_16109,N_16191);
nand U16343 (N_16343,N_16209,N_16039);
and U16344 (N_16344,N_16110,N_16069);
or U16345 (N_16345,N_16045,N_16234);
nand U16346 (N_16346,N_16161,N_16151);
nand U16347 (N_16347,N_16088,N_16231);
and U16348 (N_16348,N_16170,N_16132);
nand U16349 (N_16349,N_16137,N_16124);
or U16350 (N_16350,N_16112,N_16165);
xnor U16351 (N_16351,N_16103,N_16075);
nor U16352 (N_16352,N_16138,N_16065);
nand U16353 (N_16353,N_16094,N_16083);
or U16354 (N_16354,N_16064,N_16100);
and U16355 (N_16355,N_16005,N_16192);
nor U16356 (N_16356,N_16212,N_16108);
nor U16357 (N_16357,N_16222,N_16116);
or U16358 (N_16358,N_16119,N_16076);
nand U16359 (N_16359,N_16086,N_16117);
and U16360 (N_16360,N_16056,N_16150);
or U16361 (N_16361,N_16029,N_16169);
nor U16362 (N_16362,N_16163,N_16041);
nand U16363 (N_16363,N_16084,N_16202);
nor U16364 (N_16364,N_16216,N_16230);
xnor U16365 (N_16365,N_16130,N_16046);
or U16366 (N_16366,N_16020,N_16068);
nand U16367 (N_16367,N_16145,N_16095);
nor U16368 (N_16368,N_16027,N_16128);
xor U16369 (N_16369,N_16200,N_16204);
xnor U16370 (N_16370,N_16181,N_16080);
nor U16371 (N_16371,N_16053,N_16207);
or U16372 (N_16372,N_16049,N_16043);
or U16373 (N_16373,N_16037,N_16214);
and U16374 (N_16374,N_16048,N_16158);
or U16375 (N_16375,N_16069,N_16152);
xnor U16376 (N_16376,N_16060,N_16010);
and U16377 (N_16377,N_16066,N_16128);
and U16378 (N_16378,N_16208,N_16037);
nor U16379 (N_16379,N_16244,N_16237);
or U16380 (N_16380,N_16035,N_16039);
or U16381 (N_16381,N_16102,N_16188);
or U16382 (N_16382,N_16032,N_16216);
and U16383 (N_16383,N_16209,N_16075);
xnor U16384 (N_16384,N_16004,N_16245);
or U16385 (N_16385,N_16058,N_16047);
nor U16386 (N_16386,N_16181,N_16108);
or U16387 (N_16387,N_16240,N_16154);
nor U16388 (N_16388,N_16230,N_16127);
or U16389 (N_16389,N_16133,N_16228);
xor U16390 (N_16390,N_16062,N_16192);
or U16391 (N_16391,N_16005,N_16046);
and U16392 (N_16392,N_16037,N_16190);
nor U16393 (N_16393,N_16033,N_16223);
nand U16394 (N_16394,N_16196,N_16176);
xnor U16395 (N_16395,N_16039,N_16184);
nor U16396 (N_16396,N_16109,N_16232);
or U16397 (N_16397,N_16223,N_16066);
nor U16398 (N_16398,N_16100,N_16184);
and U16399 (N_16399,N_16129,N_16011);
nand U16400 (N_16400,N_16007,N_16005);
xnor U16401 (N_16401,N_16238,N_16012);
nor U16402 (N_16402,N_16169,N_16233);
and U16403 (N_16403,N_16043,N_16027);
and U16404 (N_16404,N_16117,N_16101);
and U16405 (N_16405,N_16043,N_16181);
or U16406 (N_16406,N_16172,N_16000);
nand U16407 (N_16407,N_16072,N_16222);
nand U16408 (N_16408,N_16239,N_16222);
nor U16409 (N_16409,N_16067,N_16093);
and U16410 (N_16410,N_16235,N_16159);
xor U16411 (N_16411,N_16058,N_16105);
nand U16412 (N_16412,N_16006,N_16107);
nor U16413 (N_16413,N_16247,N_16064);
xor U16414 (N_16414,N_16047,N_16010);
or U16415 (N_16415,N_16141,N_16209);
nand U16416 (N_16416,N_16226,N_16134);
nand U16417 (N_16417,N_16069,N_16203);
and U16418 (N_16418,N_16063,N_16024);
and U16419 (N_16419,N_16128,N_16236);
and U16420 (N_16420,N_16018,N_16044);
nor U16421 (N_16421,N_16043,N_16204);
and U16422 (N_16422,N_16244,N_16054);
and U16423 (N_16423,N_16049,N_16072);
nor U16424 (N_16424,N_16019,N_16044);
xor U16425 (N_16425,N_16126,N_16010);
and U16426 (N_16426,N_16212,N_16040);
xor U16427 (N_16427,N_16018,N_16211);
nand U16428 (N_16428,N_16051,N_16217);
or U16429 (N_16429,N_16070,N_16021);
nand U16430 (N_16430,N_16076,N_16186);
nand U16431 (N_16431,N_16157,N_16242);
nand U16432 (N_16432,N_16153,N_16049);
nand U16433 (N_16433,N_16247,N_16115);
and U16434 (N_16434,N_16167,N_16081);
xor U16435 (N_16435,N_16071,N_16027);
xor U16436 (N_16436,N_16157,N_16164);
nand U16437 (N_16437,N_16005,N_16200);
or U16438 (N_16438,N_16248,N_16008);
or U16439 (N_16439,N_16198,N_16103);
xor U16440 (N_16440,N_16047,N_16112);
xnor U16441 (N_16441,N_16218,N_16107);
or U16442 (N_16442,N_16062,N_16039);
nand U16443 (N_16443,N_16022,N_16161);
xor U16444 (N_16444,N_16153,N_16139);
and U16445 (N_16445,N_16099,N_16026);
nand U16446 (N_16446,N_16076,N_16030);
or U16447 (N_16447,N_16164,N_16052);
or U16448 (N_16448,N_16153,N_16210);
and U16449 (N_16449,N_16121,N_16030);
or U16450 (N_16450,N_16019,N_16092);
nand U16451 (N_16451,N_16094,N_16022);
nor U16452 (N_16452,N_16243,N_16241);
nor U16453 (N_16453,N_16088,N_16029);
and U16454 (N_16454,N_16198,N_16240);
nand U16455 (N_16455,N_16117,N_16052);
or U16456 (N_16456,N_16107,N_16143);
nand U16457 (N_16457,N_16142,N_16124);
and U16458 (N_16458,N_16162,N_16176);
nor U16459 (N_16459,N_16002,N_16071);
xor U16460 (N_16460,N_16236,N_16010);
xor U16461 (N_16461,N_16158,N_16000);
or U16462 (N_16462,N_16064,N_16107);
xor U16463 (N_16463,N_16115,N_16019);
and U16464 (N_16464,N_16168,N_16200);
or U16465 (N_16465,N_16215,N_16165);
nor U16466 (N_16466,N_16067,N_16159);
nor U16467 (N_16467,N_16175,N_16015);
nor U16468 (N_16468,N_16135,N_16070);
nor U16469 (N_16469,N_16243,N_16235);
or U16470 (N_16470,N_16088,N_16213);
and U16471 (N_16471,N_16032,N_16229);
nand U16472 (N_16472,N_16072,N_16197);
nand U16473 (N_16473,N_16228,N_16154);
nand U16474 (N_16474,N_16027,N_16015);
nand U16475 (N_16475,N_16113,N_16063);
and U16476 (N_16476,N_16060,N_16093);
nand U16477 (N_16477,N_16143,N_16046);
nor U16478 (N_16478,N_16031,N_16041);
or U16479 (N_16479,N_16074,N_16122);
nor U16480 (N_16480,N_16133,N_16067);
and U16481 (N_16481,N_16088,N_16133);
nor U16482 (N_16482,N_16051,N_16206);
or U16483 (N_16483,N_16118,N_16152);
or U16484 (N_16484,N_16050,N_16140);
nor U16485 (N_16485,N_16144,N_16111);
or U16486 (N_16486,N_16030,N_16117);
xnor U16487 (N_16487,N_16184,N_16029);
nor U16488 (N_16488,N_16002,N_16234);
and U16489 (N_16489,N_16128,N_16045);
nand U16490 (N_16490,N_16047,N_16242);
nand U16491 (N_16491,N_16174,N_16054);
nand U16492 (N_16492,N_16083,N_16136);
xnor U16493 (N_16493,N_16061,N_16243);
nand U16494 (N_16494,N_16189,N_16001);
or U16495 (N_16495,N_16140,N_16003);
nor U16496 (N_16496,N_16027,N_16197);
or U16497 (N_16497,N_16211,N_16019);
nand U16498 (N_16498,N_16105,N_16229);
xor U16499 (N_16499,N_16010,N_16239);
and U16500 (N_16500,N_16342,N_16439);
and U16501 (N_16501,N_16380,N_16357);
and U16502 (N_16502,N_16353,N_16309);
or U16503 (N_16503,N_16464,N_16328);
and U16504 (N_16504,N_16320,N_16422);
nor U16505 (N_16505,N_16266,N_16433);
or U16506 (N_16506,N_16445,N_16428);
nand U16507 (N_16507,N_16420,N_16360);
nor U16508 (N_16508,N_16415,N_16308);
nand U16509 (N_16509,N_16440,N_16267);
and U16510 (N_16510,N_16379,N_16306);
or U16511 (N_16511,N_16284,N_16273);
nor U16512 (N_16512,N_16251,N_16381);
nor U16513 (N_16513,N_16389,N_16408);
xnor U16514 (N_16514,N_16326,N_16329);
or U16515 (N_16515,N_16423,N_16252);
nor U16516 (N_16516,N_16369,N_16335);
or U16517 (N_16517,N_16290,N_16259);
xor U16518 (N_16518,N_16463,N_16377);
and U16519 (N_16519,N_16414,N_16449);
and U16520 (N_16520,N_16318,N_16429);
nand U16521 (N_16521,N_16270,N_16358);
nand U16522 (N_16522,N_16395,N_16253);
or U16523 (N_16523,N_16289,N_16368);
xnor U16524 (N_16524,N_16340,N_16283);
nand U16525 (N_16525,N_16456,N_16452);
nand U16526 (N_16526,N_16364,N_16269);
or U16527 (N_16527,N_16454,N_16467);
and U16528 (N_16528,N_16301,N_16255);
nor U16529 (N_16529,N_16258,N_16388);
or U16530 (N_16530,N_16485,N_16453);
or U16531 (N_16531,N_16393,N_16278);
and U16532 (N_16532,N_16332,N_16490);
or U16533 (N_16533,N_16483,N_16406);
nand U16534 (N_16534,N_16469,N_16375);
or U16535 (N_16535,N_16480,N_16392);
or U16536 (N_16536,N_16257,N_16391);
and U16537 (N_16537,N_16446,N_16465);
or U16538 (N_16538,N_16384,N_16313);
or U16539 (N_16539,N_16495,N_16302);
or U16540 (N_16540,N_16402,N_16396);
and U16541 (N_16541,N_16298,N_16441);
nand U16542 (N_16542,N_16323,N_16494);
nand U16543 (N_16543,N_16344,N_16272);
xor U16544 (N_16544,N_16333,N_16442);
xnor U16545 (N_16545,N_16427,N_16443);
nand U16546 (N_16546,N_16496,N_16482);
and U16547 (N_16547,N_16386,N_16451);
nor U16548 (N_16548,N_16492,N_16387);
or U16549 (N_16549,N_16277,N_16321);
nor U16550 (N_16550,N_16421,N_16472);
or U16551 (N_16551,N_16330,N_16411);
nand U16552 (N_16552,N_16274,N_16474);
and U16553 (N_16553,N_16322,N_16304);
or U16554 (N_16554,N_16437,N_16460);
nor U16555 (N_16555,N_16432,N_16383);
nor U16556 (N_16556,N_16405,N_16281);
or U16557 (N_16557,N_16286,N_16425);
xnor U16558 (N_16558,N_16305,N_16316);
xor U16559 (N_16559,N_16361,N_16497);
nand U16560 (N_16560,N_16307,N_16418);
or U16561 (N_16561,N_16412,N_16296);
and U16562 (N_16562,N_16498,N_16457);
and U16563 (N_16563,N_16324,N_16417);
or U16564 (N_16564,N_16435,N_16374);
xor U16565 (N_16565,N_16285,N_16426);
nor U16566 (N_16566,N_16250,N_16473);
nand U16567 (N_16567,N_16331,N_16303);
nor U16568 (N_16568,N_16484,N_16292);
nor U16569 (N_16569,N_16314,N_16294);
or U16570 (N_16570,N_16488,N_16327);
nor U16571 (N_16571,N_16399,N_16410);
nor U16572 (N_16572,N_16487,N_16350);
and U16573 (N_16573,N_16419,N_16352);
or U16574 (N_16574,N_16450,N_16373);
and U16575 (N_16575,N_16459,N_16404);
xor U16576 (N_16576,N_16493,N_16343);
nor U16577 (N_16577,N_16416,N_16462);
nand U16578 (N_16578,N_16299,N_16293);
and U16579 (N_16579,N_16471,N_16458);
nor U16580 (N_16580,N_16346,N_16268);
nand U16581 (N_16581,N_16295,N_16264);
or U16582 (N_16582,N_16300,N_16362);
nor U16583 (N_16583,N_16491,N_16363);
xor U16584 (N_16584,N_16262,N_16436);
nand U16585 (N_16585,N_16261,N_16434);
or U16586 (N_16586,N_16397,N_16351);
or U16587 (N_16587,N_16401,N_16486);
nor U16588 (N_16588,N_16297,N_16390);
and U16589 (N_16589,N_16477,N_16376);
or U16590 (N_16590,N_16339,N_16385);
nor U16591 (N_16591,N_16430,N_16382);
and U16592 (N_16592,N_16347,N_16279);
nand U16593 (N_16593,N_16478,N_16407);
and U16594 (N_16594,N_16319,N_16365);
or U16595 (N_16595,N_16312,N_16489);
nand U16596 (N_16596,N_16348,N_16359);
xnor U16597 (N_16597,N_16499,N_16468);
nor U16598 (N_16598,N_16371,N_16317);
and U16599 (N_16599,N_16349,N_16275);
and U16600 (N_16600,N_16288,N_16479);
nor U16601 (N_16601,N_16413,N_16345);
or U16602 (N_16602,N_16341,N_16431);
nand U16603 (N_16603,N_16476,N_16400);
nor U16604 (N_16604,N_16265,N_16481);
and U16605 (N_16605,N_16263,N_16315);
and U16606 (N_16606,N_16254,N_16378);
nor U16607 (N_16607,N_16372,N_16455);
or U16608 (N_16608,N_16356,N_16282);
nand U16609 (N_16609,N_16409,N_16276);
or U16610 (N_16610,N_16355,N_16334);
or U16611 (N_16611,N_16311,N_16310);
nand U16612 (N_16612,N_16438,N_16366);
nand U16613 (N_16613,N_16466,N_16444);
xnor U16614 (N_16614,N_16394,N_16291);
and U16615 (N_16615,N_16447,N_16367);
nand U16616 (N_16616,N_16337,N_16260);
and U16617 (N_16617,N_16398,N_16336);
nor U16618 (N_16618,N_16325,N_16338);
or U16619 (N_16619,N_16461,N_16256);
or U16620 (N_16620,N_16287,N_16424);
and U16621 (N_16621,N_16470,N_16403);
nor U16622 (N_16622,N_16475,N_16370);
or U16623 (N_16623,N_16271,N_16354);
or U16624 (N_16624,N_16448,N_16280);
and U16625 (N_16625,N_16469,N_16326);
and U16626 (N_16626,N_16496,N_16324);
or U16627 (N_16627,N_16472,N_16363);
nand U16628 (N_16628,N_16421,N_16435);
or U16629 (N_16629,N_16253,N_16344);
or U16630 (N_16630,N_16374,N_16314);
and U16631 (N_16631,N_16393,N_16295);
nor U16632 (N_16632,N_16257,N_16275);
nor U16633 (N_16633,N_16490,N_16267);
or U16634 (N_16634,N_16376,N_16414);
nor U16635 (N_16635,N_16272,N_16456);
nand U16636 (N_16636,N_16404,N_16462);
or U16637 (N_16637,N_16401,N_16357);
or U16638 (N_16638,N_16335,N_16465);
and U16639 (N_16639,N_16356,N_16298);
nand U16640 (N_16640,N_16375,N_16448);
and U16641 (N_16641,N_16330,N_16321);
nor U16642 (N_16642,N_16396,N_16260);
or U16643 (N_16643,N_16343,N_16377);
nand U16644 (N_16644,N_16400,N_16402);
and U16645 (N_16645,N_16254,N_16356);
nor U16646 (N_16646,N_16256,N_16465);
and U16647 (N_16647,N_16325,N_16365);
or U16648 (N_16648,N_16448,N_16442);
xor U16649 (N_16649,N_16492,N_16306);
nor U16650 (N_16650,N_16317,N_16363);
and U16651 (N_16651,N_16476,N_16261);
nor U16652 (N_16652,N_16426,N_16420);
nor U16653 (N_16653,N_16319,N_16364);
nand U16654 (N_16654,N_16327,N_16436);
or U16655 (N_16655,N_16278,N_16484);
or U16656 (N_16656,N_16325,N_16410);
and U16657 (N_16657,N_16269,N_16381);
or U16658 (N_16658,N_16300,N_16395);
nor U16659 (N_16659,N_16464,N_16331);
nor U16660 (N_16660,N_16349,N_16331);
and U16661 (N_16661,N_16286,N_16414);
and U16662 (N_16662,N_16358,N_16405);
and U16663 (N_16663,N_16427,N_16341);
xor U16664 (N_16664,N_16432,N_16330);
nand U16665 (N_16665,N_16277,N_16269);
nand U16666 (N_16666,N_16311,N_16300);
and U16667 (N_16667,N_16482,N_16362);
nand U16668 (N_16668,N_16298,N_16470);
nand U16669 (N_16669,N_16450,N_16480);
nor U16670 (N_16670,N_16295,N_16427);
and U16671 (N_16671,N_16391,N_16437);
nor U16672 (N_16672,N_16464,N_16272);
nor U16673 (N_16673,N_16440,N_16478);
nor U16674 (N_16674,N_16373,N_16255);
nand U16675 (N_16675,N_16422,N_16291);
and U16676 (N_16676,N_16488,N_16268);
or U16677 (N_16677,N_16454,N_16424);
nand U16678 (N_16678,N_16293,N_16436);
and U16679 (N_16679,N_16413,N_16341);
xor U16680 (N_16680,N_16499,N_16284);
xnor U16681 (N_16681,N_16453,N_16491);
xor U16682 (N_16682,N_16322,N_16446);
nor U16683 (N_16683,N_16313,N_16470);
nor U16684 (N_16684,N_16359,N_16294);
or U16685 (N_16685,N_16435,N_16465);
nand U16686 (N_16686,N_16282,N_16419);
nor U16687 (N_16687,N_16316,N_16428);
nor U16688 (N_16688,N_16305,N_16291);
and U16689 (N_16689,N_16291,N_16343);
or U16690 (N_16690,N_16304,N_16259);
or U16691 (N_16691,N_16380,N_16430);
and U16692 (N_16692,N_16299,N_16373);
or U16693 (N_16693,N_16320,N_16390);
or U16694 (N_16694,N_16335,N_16366);
nor U16695 (N_16695,N_16453,N_16499);
nor U16696 (N_16696,N_16441,N_16361);
nand U16697 (N_16697,N_16274,N_16498);
nor U16698 (N_16698,N_16420,N_16414);
and U16699 (N_16699,N_16483,N_16347);
nor U16700 (N_16700,N_16331,N_16334);
or U16701 (N_16701,N_16493,N_16300);
xnor U16702 (N_16702,N_16488,N_16431);
or U16703 (N_16703,N_16440,N_16491);
and U16704 (N_16704,N_16417,N_16355);
nand U16705 (N_16705,N_16311,N_16464);
nor U16706 (N_16706,N_16345,N_16360);
or U16707 (N_16707,N_16331,N_16451);
nand U16708 (N_16708,N_16330,N_16417);
xnor U16709 (N_16709,N_16400,N_16458);
xnor U16710 (N_16710,N_16463,N_16388);
and U16711 (N_16711,N_16472,N_16400);
nor U16712 (N_16712,N_16369,N_16283);
or U16713 (N_16713,N_16481,N_16325);
or U16714 (N_16714,N_16405,N_16496);
nand U16715 (N_16715,N_16308,N_16297);
nor U16716 (N_16716,N_16374,N_16439);
and U16717 (N_16717,N_16397,N_16251);
or U16718 (N_16718,N_16303,N_16354);
nor U16719 (N_16719,N_16472,N_16456);
nor U16720 (N_16720,N_16444,N_16265);
or U16721 (N_16721,N_16438,N_16480);
and U16722 (N_16722,N_16495,N_16438);
xor U16723 (N_16723,N_16284,N_16381);
and U16724 (N_16724,N_16432,N_16307);
nand U16725 (N_16725,N_16286,N_16447);
and U16726 (N_16726,N_16337,N_16391);
nand U16727 (N_16727,N_16351,N_16275);
or U16728 (N_16728,N_16297,N_16354);
and U16729 (N_16729,N_16341,N_16367);
nor U16730 (N_16730,N_16464,N_16441);
xnor U16731 (N_16731,N_16290,N_16450);
or U16732 (N_16732,N_16278,N_16437);
or U16733 (N_16733,N_16314,N_16443);
xnor U16734 (N_16734,N_16283,N_16254);
nor U16735 (N_16735,N_16264,N_16337);
nand U16736 (N_16736,N_16276,N_16331);
and U16737 (N_16737,N_16326,N_16380);
nor U16738 (N_16738,N_16491,N_16374);
or U16739 (N_16739,N_16418,N_16354);
xnor U16740 (N_16740,N_16316,N_16264);
or U16741 (N_16741,N_16295,N_16428);
nor U16742 (N_16742,N_16437,N_16381);
nor U16743 (N_16743,N_16331,N_16336);
nor U16744 (N_16744,N_16313,N_16486);
or U16745 (N_16745,N_16263,N_16394);
and U16746 (N_16746,N_16276,N_16428);
and U16747 (N_16747,N_16489,N_16272);
and U16748 (N_16748,N_16449,N_16492);
and U16749 (N_16749,N_16420,N_16359);
or U16750 (N_16750,N_16690,N_16504);
nor U16751 (N_16751,N_16634,N_16571);
or U16752 (N_16752,N_16675,N_16554);
and U16753 (N_16753,N_16654,N_16535);
xor U16754 (N_16754,N_16505,N_16596);
nand U16755 (N_16755,N_16702,N_16600);
and U16756 (N_16756,N_16614,N_16689);
and U16757 (N_16757,N_16575,N_16644);
nor U16758 (N_16758,N_16706,N_16549);
nand U16759 (N_16759,N_16522,N_16602);
or U16760 (N_16760,N_16550,N_16532);
and U16761 (N_16761,N_16525,N_16703);
and U16762 (N_16762,N_16607,N_16520);
nand U16763 (N_16763,N_16743,N_16728);
or U16764 (N_16764,N_16727,N_16611);
or U16765 (N_16765,N_16649,N_16552);
or U16766 (N_16766,N_16618,N_16686);
xor U16767 (N_16767,N_16632,N_16544);
or U16768 (N_16768,N_16709,N_16734);
nand U16769 (N_16769,N_16601,N_16529);
and U16770 (N_16770,N_16643,N_16513);
and U16771 (N_16771,N_16569,N_16674);
and U16772 (N_16772,N_16722,N_16630);
and U16773 (N_16773,N_16666,N_16555);
and U16774 (N_16774,N_16588,N_16567);
or U16775 (N_16775,N_16700,N_16633);
and U16776 (N_16776,N_16723,N_16534);
nand U16777 (N_16777,N_16669,N_16506);
nor U16778 (N_16778,N_16545,N_16629);
and U16779 (N_16779,N_16548,N_16578);
nor U16780 (N_16780,N_16647,N_16608);
and U16781 (N_16781,N_16655,N_16673);
nor U16782 (N_16782,N_16694,N_16711);
or U16783 (N_16783,N_16605,N_16665);
xor U16784 (N_16784,N_16697,N_16540);
nor U16785 (N_16785,N_16720,N_16736);
nor U16786 (N_16786,N_16667,N_16716);
nand U16787 (N_16787,N_16682,N_16719);
nor U16788 (N_16788,N_16714,N_16586);
nand U16789 (N_16789,N_16565,N_16701);
nor U16790 (N_16790,N_16536,N_16515);
xnor U16791 (N_16791,N_16585,N_16672);
or U16792 (N_16792,N_16599,N_16574);
or U16793 (N_16793,N_16712,N_16748);
and U16794 (N_16794,N_16635,N_16645);
xor U16795 (N_16795,N_16528,N_16713);
and U16796 (N_16796,N_16636,N_16721);
nor U16797 (N_16797,N_16501,N_16741);
nand U16798 (N_16798,N_16546,N_16509);
xnor U16799 (N_16799,N_16622,N_16747);
nand U16800 (N_16800,N_16559,N_16742);
and U16801 (N_16801,N_16612,N_16749);
nand U16802 (N_16802,N_16729,N_16652);
or U16803 (N_16803,N_16537,N_16597);
or U16804 (N_16804,N_16651,N_16648);
nand U16805 (N_16805,N_16606,N_16561);
or U16806 (N_16806,N_16609,N_16676);
nand U16807 (N_16807,N_16510,N_16604);
or U16808 (N_16808,N_16646,N_16507);
and U16809 (N_16809,N_16625,N_16627);
or U16810 (N_16810,N_16512,N_16572);
nand U16811 (N_16811,N_16542,N_16725);
and U16812 (N_16812,N_16637,N_16615);
or U16813 (N_16813,N_16500,N_16718);
or U16814 (N_16814,N_16731,N_16590);
nor U16815 (N_16815,N_16623,N_16710);
xor U16816 (N_16816,N_16558,N_16613);
nand U16817 (N_16817,N_16735,N_16527);
xor U16818 (N_16818,N_16530,N_16547);
or U16819 (N_16819,N_16740,N_16705);
and U16820 (N_16820,N_16661,N_16587);
nand U16821 (N_16821,N_16603,N_16591);
or U16822 (N_16822,N_16678,N_16662);
nor U16823 (N_16823,N_16557,N_16650);
nor U16824 (N_16824,N_16564,N_16579);
nor U16825 (N_16825,N_16692,N_16685);
nand U16826 (N_16826,N_16539,N_16626);
and U16827 (N_16827,N_16593,N_16670);
nor U16828 (N_16828,N_16733,N_16715);
nand U16829 (N_16829,N_16659,N_16553);
nand U16830 (N_16830,N_16511,N_16744);
and U16831 (N_16831,N_16533,N_16704);
xor U16832 (N_16832,N_16680,N_16589);
and U16833 (N_16833,N_16624,N_16562);
or U16834 (N_16834,N_16642,N_16502);
nand U16835 (N_16835,N_16566,N_16683);
or U16836 (N_16836,N_16573,N_16679);
or U16837 (N_16837,N_16707,N_16577);
nor U16838 (N_16838,N_16746,N_16580);
nand U16839 (N_16839,N_16583,N_16738);
nor U16840 (N_16840,N_16668,N_16677);
and U16841 (N_16841,N_16737,N_16508);
xor U16842 (N_16842,N_16556,N_16628);
nand U16843 (N_16843,N_16517,N_16518);
nand U16844 (N_16844,N_16581,N_16663);
and U16845 (N_16845,N_16598,N_16730);
and U16846 (N_16846,N_16687,N_16732);
nand U16847 (N_16847,N_16592,N_16568);
or U16848 (N_16848,N_16671,N_16576);
nand U16849 (N_16849,N_16631,N_16524);
and U16850 (N_16850,N_16541,N_16739);
and U16851 (N_16851,N_16519,N_16516);
or U16852 (N_16852,N_16745,N_16695);
and U16853 (N_16853,N_16621,N_16620);
nor U16854 (N_16854,N_16619,N_16657);
or U16855 (N_16855,N_16639,N_16664);
nor U16856 (N_16856,N_16616,N_16543);
nor U16857 (N_16857,N_16521,N_16688);
or U16858 (N_16858,N_16523,N_16724);
nand U16859 (N_16859,N_16681,N_16595);
or U16860 (N_16860,N_16641,N_16640);
nor U16861 (N_16861,N_16514,N_16691);
and U16862 (N_16862,N_16594,N_16526);
nor U16863 (N_16863,N_16538,N_16658);
nand U16864 (N_16864,N_16563,N_16696);
and U16865 (N_16865,N_16560,N_16699);
and U16866 (N_16866,N_16708,N_16698);
and U16867 (N_16867,N_16717,N_16551);
or U16868 (N_16868,N_16582,N_16653);
xnor U16869 (N_16869,N_16584,N_16503);
nand U16870 (N_16870,N_16656,N_16617);
nor U16871 (N_16871,N_16570,N_16638);
nor U16872 (N_16872,N_16660,N_16610);
or U16873 (N_16873,N_16726,N_16684);
or U16874 (N_16874,N_16531,N_16693);
nand U16875 (N_16875,N_16673,N_16675);
or U16876 (N_16876,N_16637,N_16646);
or U16877 (N_16877,N_16641,N_16542);
and U16878 (N_16878,N_16551,N_16558);
nor U16879 (N_16879,N_16614,N_16508);
or U16880 (N_16880,N_16525,N_16668);
and U16881 (N_16881,N_16679,N_16649);
xnor U16882 (N_16882,N_16602,N_16640);
and U16883 (N_16883,N_16521,N_16619);
and U16884 (N_16884,N_16671,N_16679);
nand U16885 (N_16885,N_16722,N_16687);
or U16886 (N_16886,N_16740,N_16512);
nor U16887 (N_16887,N_16555,N_16624);
nor U16888 (N_16888,N_16511,N_16703);
xnor U16889 (N_16889,N_16578,N_16737);
or U16890 (N_16890,N_16592,N_16718);
nor U16891 (N_16891,N_16747,N_16573);
and U16892 (N_16892,N_16511,N_16645);
nor U16893 (N_16893,N_16595,N_16688);
and U16894 (N_16894,N_16566,N_16641);
nor U16895 (N_16895,N_16513,N_16663);
nand U16896 (N_16896,N_16669,N_16501);
and U16897 (N_16897,N_16710,N_16573);
xnor U16898 (N_16898,N_16539,N_16659);
nor U16899 (N_16899,N_16629,N_16674);
and U16900 (N_16900,N_16585,N_16575);
nand U16901 (N_16901,N_16608,N_16628);
nand U16902 (N_16902,N_16588,N_16598);
nor U16903 (N_16903,N_16580,N_16726);
nand U16904 (N_16904,N_16633,N_16733);
or U16905 (N_16905,N_16517,N_16529);
and U16906 (N_16906,N_16649,N_16684);
and U16907 (N_16907,N_16555,N_16508);
or U16908 (N_16908,N_16526,N_16716);
or U16909 (N_16909,N_16544,N_16608);
nor U16910 (N_16910,N_16557,N_16621);
and U16911 (N_16911,N_16663,N_16520);
or U16912 (N_16912,N_16638,N_16529);
xor U16913 (N_16913,N_16597,N_16576);
or U16914 (N_16914,N_16625,N_16531);
nand U16915 (N_16915,N_16625,N_16689);
or U16916 (N_16916,N_16680,N_16585);
and U16917 (N_16917,N_16552,N_16531);
nor U16918 (N_16918,N_16551,N_16727);
nor U16919 (N_16919,N_16719,N_16535);
or U16920 (N_16920,N_16551,N_16606);
and U16921 (N_16921,N_16505,N_16613);
xor U16922 (N_16922,N_16600,N_16741);
or U16923 (N_16923,N_16590,N_16666);
or U16924 (N_16924,N_16621,N_16535);
xor U16925 (N_16925,N_16578,N_16575);
xnor U16926 (N_16926,N_16516,N_16580);
nand U16927 (N_16927,N_16574,N_16548);
and U16928 (N_16928,N_16560,N_16725);
nand U16929 (N_16929,N_16542,N_16716);
nand U16930 (N_16930,N_16667,N_16552);
nor U16931 (N_16931,N_16681,N_16691);
xnor U16932 (N_16932,N_16711,N_16729);
nand U16933 (N_16933,N_16713,N_16735);
and U16934 (N_16934,N_16645,N_16681);
and U16935 (N_16935,N_16656,N_16715);
xor U16936 (N_16936,N_16661,N_16685);
nand U16937 (N_16937,N_16730,N_16581);
nor U16938 (N_16938,N_16615,N_16539);
xnor U16939 (N_16939,N_16632,N_16698);
xor U16940 (N_16940,N_16511,N_16556);
and U16941 (N_16941,N_16684,N_16588);
nor U16942 (N_16942,N_16735,N_16656);
nor U16943 (N_16943,N_16631,N_16564);
and U16944 (N_16944,N_16610,N_16577);
nor U16945 (N_16945,N_16603,N_16514);
or U16946 (N_16946,N_16670,N_16570);
nand U16947 (N_16947,N_16745,N_16704);
nor U16948 (N_16948,N_16700,N_16677);
and U16949 (N_16949,N_16519,N_16529);
nand U16950 (N_16950,N_16610,N_16640);
or U16951 (N_16951,N_16529,N_16541);
or U16952 (N_16952,N_16748,N_16624);
and U16953 (N_16953,N_16531,N_16689);
nand U16954 (N_16954,N_16666,N_16560);
nand U16955 (N_16955,N_16681,N_16529);
nor U16956 (N_16956,N_16591,N_16740);
or U16957 (N_16957,N_16554,N_16703);
and U16958 (N_16958,N_16690,N_16510);
xor U16959 (N_16959,N_16690,N_16571);
or U16960 (N_16960,N_16541,N_16628);
nand U16961 (N_16961,N_16666,N_16696);
or U16962 (N_16962,N_16650,N_16580);
or U16963 (N_16963,N_16677,N_16559);
nand U16964 (N_16964,N_16563,N_16564);
xnor U16965 (N_16965,N_16618,N_16542);
and U16966 (N_16966,N_16562,N_16682);
nor U16967 (N_16967,N_16584,N_16668);
nand U16968 (N_16968,N_16567,N_16563);
nand U16969 (N_16969,N_16579,N_16522);
nand U16970 (N_16970,N_16636,N_16686);
xor U16971 (N_16971,N_16744,N_16527);
or U16972 (N_16972,N_16589,N_16522);
or U16973 (N_16973,N_16733,N_16736);
or U16974 (N_16974,N_16651,N_16671);
nor U16975 (N_16975,N_16636,N_16509);
and U16976 (N_16976,N_16688,N_16501);
and U16977 (N_16977,N_16628,N_16502);
and U16978 (N_16978,N_16572,N_16681);
nand U16979 (N_16979,N_16588,N_16674);
nor U16980 (N_16980,N_16719,N_16521);
and U16981 (N_16981,N_16638,N_16552);
nand U16982 (N_16982,N_16627,N_16705);
or U16983 (N_16983,N_16694,N_16624);
and U16984 (N_16984,N_16617,N_16641);
or U16985 (N_16985,N_16549,N_16559);
and U16986 (N_16986,N_16663,N_16518);
nand U16987 (N_16987,N_16672,N_16714);
or U16988 (N_16988,N_16558,N_16659);
nand U16989 (N_16989,N_16561,N_16683);
nand U16990 (N_16990,N_16644,N_16500);
nor U16991 (N_16991,N_16727,N_16558);
nand U16992 (N_16992,N_16735,N_16622);
nor U16993 (N_16993,N_16571,N_16706);
nand U16994 (N_16994,N_16526,N_16503);
nand U16995 (N_16995,N_16514,N_16732);
xor U16996 (N_16996,N_16597,N_16560);
nor U16997 (N_16997,N_16602,N_16665);
nor U16998 (N_16998,N_16727,N_16681);
xor U16999 (N_16999,N_16670,N_16641);
or U17000 (N_17000,N_16981,N_16941);
or U17001 (N_17001,N_16977,N_16863);
or U17002 (N_17002,N_16838,N_16996);
or U17003 (N_17003,N_16766,N_16908);
nor U17004 (N_17004,N_16982,N_16866);
xnor U17005 (N_17005,N_16767,N_16752);
nand U17006 (N_17006,N_16761,N_16760);
xor U17007 (N_17007,N_16844,N_16913);
or U17008 (N_17008,N_16832,N_16876);
or U17009 (N_17009,N_16872,N_16772);
or U17010 (N_17010,N_16971,N_16785);
or U17011 (N_17011,N_16815,N_16823);
or U17012 (N_17012,N_16993,N_16888);
nand U17013 (N_17013,N_16972,N_16892);
and U17014 (N_17014,N_16789,N_16847);
nand U17015 (N_17015,N_16975,N_16919);
or U17016 (N_17016,N_16841,N_16895);
or U17017 (N_17017,N_16867,N_16936);
nand U17018 (N_17018,N_16950,N_16860);
nor U17019 (N_17019,N_16927,N_16986);
xor U17020 (N_17020,N_16859,N_16764);
nand U17021 (N_17021,N_16973,N_16791);
xnor U17022 (N_17022,N_16976,N_16902);
nand U17023 (N_17023,N_16934,N_16962);
nand U17024 (N_17024,N_16937,N_16834);
nand U17025 (N_17025,N_16978,N_16850);
nand U17026 (N_17026,N_16904,N_16935);
or U17027 (N_17027,N_16906,N_16967);
xor U17028 (N_17028,N_16826,N_16958);
nand U17029 (N_17029,N_16756,N_16802);
nor U17030 (N_17030,N_16883,N_16852);
xnor U17031 (N_17031,N_16818,N_16956);
and U17032 (N_17032,N_16920,N_16991);
xor U17033 (N_17033,N_16942,N_16851);
and U17034 (N_17034,N_16944,N_16914);
and U17035 (N_17035,N_16911,N_16932);
nor U17036 (N_17036,N_16763,N_16905);
or U17037 (N_17037,N_16759,N_16819);
xor U17038 (N_17038,N_16984,N_16994);
nand U17039 (N_17039,N_16774,N_16943);
nand U17040 (N_17040,N_16786,N_16870);
or U17041 (N_17041,N_16762,N_16881);
and U17042 (N_17042,N_16813,N_16931);
nand U17043 (N_17043,N_16947,N_16821);
nor U17044 (N_17044,N_16897,N_16829);
nand U17045 (N_17045,N_16926,N_16960);
nand U17046 (N_17046,N_16896,N_16801);
nand U17047 (N_17047,N_16803,N_16778);
nand U17048 (N_17048,N_16854,N_16957);
and U17049 (N_17049,N_16768,N_16753);
nand U17050 (N_17050,N_16833,N_16842);
or U17051 (N_17051,N_16800,N_16884);
nor U17052 (N_17052,N_16946,N_16938);
and U17053 (N_17053,N_16828,N_16792);
nor U17054 (N_17054,N_16900,N_16755);
nor U17055 (N_17055,N_16979,N_16835);
and U17056 (N_17056,N_16865,N_16848);
xor U17057 (N_17057,N_16775,N_16793);
and U17058 (N_17058,N_16930,N_16916);
or U17059 (N_17059,N_16794,N_16809);
nor U17060 (N_17060,N_16907,N_16857);
or U17061 (N_17061,N_16757,N_16814);
and U17062 (N_17062,N_16776,N_16773);
nor U17063 (N_17063,N_16827,N_16945);
and U17064 (N_17064,N_16806,N_16771);
or U17065 (N_17065,N_16893,N_16990);
or U17066 (N_17066,N_16878,N_16940);
or U17067 (N_17067,N_16923,N_16846);
or U17068 (N_17068,N_16858,N_16825);
or U17069 (N_17069,N_16751,N_16784);
or U17070 (N_17070,N_16843,N_16961);
nor U17071 (N_17071,N_16782,N_16929);
xnor U17072 (N_17072,N_16915,N_16985);
or U17073 (N_17073,N_16822,N_16820);
nor U17074 (N_17074,N_16951,N_16839);
or U17075 (N_17075,N_16777,N_16901);
nor U17076 (N_17076,N_16995,N_16816);
nor U17077 (N_17077,N_16871,N_16918);
nor U17078 (N_17078,N_16840,N_16894);
nand U17079 (N_17079,N_16868,N_16799);
or U17080 (N_17080,N_16817,N_16890);
nor U17081 (N_17081,N_16925,N_16965);
and U17082 (N_17082,N_16966,N_16928);
nand U17083 (N_17083,N_16989,N_16810);
nand U17084 (N_17084,N_16998,N_16797);
and U17085 (N_17085,N_16889,N_16770);
nand U17086 (N_17086,N_16811,N_16952);
and U17087 (N_17087,N_16974,N_16855);
nand U17088 (N_17088,N_16765,N_16917);
and U17089 (N_17089,N_16922,N_16798);
or U17090 (N_17090,N_16836,N_16963);
nand U17091 (N_17091,N_16861,N_16970);
and U17092 (N_17092,N_16796,N_16783);
nand U17093 (N_17093,N_16808,N_16795);
and U17094 (N_17094,N_16869,N_16912);
nor U17095 (N_17095,N_16987,N_16877);
xnor U17096 (N_17096,N_16910,N_16831);
and U17097 (N_17097,N_16909,N_16837);
xnor U17098 (N_17098,N_16999,N_16824);
or U17099 (N_17099,N_16880,N_16864);
or U17100 (N_17100,N_16862,N_16879);
and U17101 (N_17101,N_16886,N_16921);
and U17102 (N_17102,N_16875,N_16845);
or U17103 (N_17103,N_16754,N_16853);
and U17104 (N_17104,N_16924,N_16882);
and U17105 (N_17105,N_16788,N_16769);
and U17106 (N_17106,N_16830,N_16885);
xnor U17107 (N_17107,N_16898,N_16887);
nand U17108 (N_17108,N_16849,N_16949);
nor U17109 (N_17109,N_16983,N_16968);
and U17110 (N_17110,N_16969,N_16954);
and U17111 (N_17111,N_16780,N_16903);
xor U17112 (N_17112,N_16953,N_16891);
or U17113 (N_17113,N_16959,N_16787);
nand U17114 (N_17114,N_16750,N_16804);
and U17115 (N_17115,N_16781,N_16933);
nand U17116 (N_17116,N_16758,N_16805);
nor U17117 (N_17117,N_16899,N_16790);
nand U17118 (N_17118,N_16997,N_16812);
or U17119 (N_17119,N_16992,N_16939);
nand U17120 (N_17120,N_16779,N_16988);
nor U17121 (N_17121,N_16980,N_16874);
or U17122 (N_17122,N_16856,N_16948);
nor U17123 (N_17123,N_16807,N_16964);
nor U17124 (N_17124,N_16873,N_16955);
nand U17125 (N_17125,N_16838,N_16932);
xor U17126 (N_17126,N_16829,N_16961);
xnor U17127 (N_17127,N_16786,N_16752);
and U17128 (N_17128,N_16946,N_16869);
and U17129 (N_17129,N_16770,N_16778);
xor U17130 (N_17130,N_16852,N_16989);
nor U17131 (N_17131,N_16845,N_16910);
and U17132 (N_17132,N_16882,N_16818);
nand U17133 (N_17133,N_16905,N_16890);
nor U17134 (N_17134,N_16921,N_16888);
nor U17135 (N_17135,N_16891,N_16761);
nand U17136 (N_17136,N_16957,N_16938);
or U17137 (N_17137,N_16800,N_16801);
or U17138 (N_17138,N_16899,N_16891);
and U17139 (N_17139,N_16919,N_16944);
xor U17140 (N_17140,N_16831,N_16788);
and U17141 (N_17141,N_16773,N_16985);
xor U17142 (N_17142,N_16939,N_16856);
nand U17143 (N_17143,N_16912,N_16903);
or U17144 (N_17144,N_16830,N_16775);
nand U17145 (N_17145,N_16919,N_16883);
nor U17146 (N_17146,N_16755,N_16917);
or U17147 (N_17147,N_16793,N_16858);
nor U17148 (N_17148,N_16962,N_16774);
nor U17149 (N_17149,N_16753,N_16981);
nor U17150 (N_17150,N_16886,N_16813);
nor U17151 (N_17151,N_16752,N_16983);
nand U17152 (N_17152,N_16818,N_16804);
nor U17153 (N_17153,N_16803,N_16970);
or U17154 (N_17154,N_16796,N_16934);
nand U17155 (N_17155,N_16898,N_16928);
or U17156 (N_17156,N_16911,N_16865);
xnor U17157 (N_17157,N_16813,N_16863);
nand U17158 (N_17158,N_16943,N_16773);
or U17159 (N_17159,N_16768,N_16773);
and U17160 (N_17160,N_16882,N_16915);
nor U17161 (N_17161,N_16984,N_16956);
nand U17162 (N_17162,N_16787,N_16920);
and U17163 (N_17163,N_16974,N_16945);
and U17164 (N_17164,N_16794,N_16913);
nor U17165 (N_17165,N_16789,N_16942);
nand U17166 (N_17166,N_16939,N_16794);
nand U17167 (N_17167,N_16908,N_16965);
nand U17168 (N_17168,N_16981,N_16972);
or U17169 (N_17169,N_16955,N_16916);
or U17170 (N_17170,N_16926,N_16975);
nor U17171 (N_17171,N_16950,N_16943);
and U17172 (N_17172,N_16900,N_16840);
and U17173 (N_17173,N_16759,N_16945);
nand U17174 (N_17174,N_16892,N_16851);
or U17175 (N_17175,N_16961,N_16761);
nor U17176 (N_17176,N_16858,N_16946);
or U17177 (N_17177,N_16847,N_16827);
nand U17178 (N_17178,N_16751,N_16884);
or U17179 (N_17179,N_16881,N_16898);
nor U17180 (N_17180,N_16811,N_16930);
or U17181 (N_17181,N_16936,N_16763);
nand U17182 (N_17182,N_16959,N_16848);
nor U17183 (N_17183,N_16995,N_16966);
nand U17184 (N_17184,N_16886,N_16827);
nand U17185 (N_17185,N_16983,N_16955);
or U17186 (N_17186,N_16953,N_16833);
and U17187 (N_17187,N_16840,N_16830);
and U17188 (N_17188,N_16814,N_16989);
or U17189 (N_17189,N_16855,N_16847);
or U17190 (N_17190,N_16825,N_16904);
nor U17191 (N_17191,N_16991,N_16763);
nand U17192 (N_17192,N_16964,N_16813);
xnor U17193 (N_17193,N_16807,N_16892);
and U17194 (N_17194,N_16942,N_16929);
nor U17195 (N_17195,N_16904,N_16838);
or U17196 (N_17196,N_16832,N_16768);
nand U17197 (N_17197,N_16797,N_16921);
nand U17198 (N_17198,N_16750,N_16862);
nand U17199 (N_17199,N_16790,N_16881);
or U17200 (N_17200,N_16808,N_16811);
or U17201 (N_17201,N_16971,N_16784);
xor U17202 (N_17202,N_16920,N_16997);
or U17203 (N_17203,N_16828,N_16998);
and U17204 (N_17204,N_16886,N_16907);
nor U17205 (N_17205,N_16854,N_16823);
nor U17206 (N_17206,N_16890,N_16954);
nor U17207 (N_17207,N_16832,N_16900);
nand U17208 (N_17208,N_16857,N_16968);
and U17209 (N_17209,N_16924,N_16834);
nand U17210 (N_17210,N_16943,N_16963);
xor U17211 (N_17211,N_16939,N_16875);
and U17212 (N_17212,N_16841,N_16976);
nor U17213 (N_17213,N_16953,N_16750);
or U17214 (N_17214,N_16814,N_16969);
or U17215 (N_17215,N_16979,N_16911);
and U17216 (N_17216,N_16843,N_16982);
or U17217 (N_17217,N_16909,N_16900);
nand U17218 (N_17218,N_16756,N_16806);
nor U17219 (N_17219,N_16822,N_16870);
nor U17220 (N_17220,N_16821,N_16780);
and U17221 (N_17221,N_16854,N_16820);
nand U17222 (N_17222,N_16991,N_16908);
nor U17223 (N_17223,N_16900,N_16923);
nor U17224 (N_17224,N_16988,N_16823);
xor U17225 (N_17225,N_16807,N_16766);
nor U17226 (N_17226,N_16834,N_16854);
or U17227 (N_17227,N_16999,N_16857);
and U17228 (N_17228,N_16850,N_16752);
xnor U17229 (N_17229,N_16923,N_16959);
nand U17230 (N_17230,N_16952,N_16804);
and U17231 (N_17231,N_16936,N_16809);
nand U17232 (N_17232,N_16784,N_16837);
or U17233 (N_17233,N_16987,N_16968);
nor U17234 (N_17234,N_16777,N_16834);
nand U17235 (N_17235,N_16907,N_16963);
nor U17236 (N_17236,N_16923,N_16985);
and U17237 (N_17237,N_16751,N_16904);
nand U17238 (N_17238,N_16951,N_16933);
nor U17239 (N_17239,N_16972,N_16876);
nor U17240 (N_17240,N_16933,N_16980);
and U17241 (N_17241,N_16811,N_16992);
and U17242 (N_17242,N_16874,N_16752);
nor U17243 (N_17243,N_16944,N_16921);
and U17244 (N_17244,N_16782,N_16868);
and U17245 (N_17245,N_16849,N_16916);
and U17246 (N_17246,N_16918,N_16869);
and U17247 (N_17247,N_16995,N_16991);
xnor U17248 (N_17248,N_16837,N_16798);
nor U17249 (N_17249,N_16847,N_16882);
and U17250 (N_17250,N_17142,N_17005);
xor U17251 (N_17251,N_17034,N_17062);
nor U17252 (N_17252,N_17087,N_17052);
and U17253 (N_17253,N_17233,N_17159);
nor U17254 (N_17254,N_17056,N_17079);
or U17255 (N_17255,N_17118,N_17019);
or U17256 (N_17256,N_17100,N_17096);
and U17257 (N_17257,N_17182,N_17082);
or U17258 (N_17258,N_17149,N_17178);
nor U17259 (N_17259,N_17176,N_17048);
nor U17260 (N_17260,N_17055,N_17217);
or U17261 (N_17261,N_17141,N_17059);
nor U17262 (N_17262,N_17058,N_17115);
or U17263 (N_17263,N_17084,N_17161);
nor U17264 (N_17264,N_17114,N_17077);
nand U17265 (N_17265,N_17071,N_17249);
nand U17266 (N_17266,N_17125,N_17183);
and U17267 (N_17267,N_17037,N_17074);
and U17268 (N_17268,N_17193,N_17234);
nand U17269 (N_17269,N_17136,N_17007);
or U17270 (N_17270,N_17085,N_17145);
nor U17271 (N_17271,N_17002,N_17154);
nand U17272 (N_17272,N_17091,N_17033);
xnor U17273 (N_17273,N_17194,N_17102);
nor U17274 (N_17274,N_17119,N_17137);
xnor U17275 (N_17275,N_17029,N_17143);
or U17276 (N_17276,N_17127,N_17173);
and U17277 (N_17277,N_17185,N_17057);
nor U17278 (N_17278,N_17101,N_17032);
or U17279 (N_17279,N_17236,N_17230);
nor U17280 (N_17280,N_17139,N_17020);
nor U17281 (N_17281,N_17109,N_17080);
nand U17282 (N_17282,N_17014,N_17140);
or U17283 (N_17283,N_17174,N_17244);
nor U17284 (N_17284,N_17012,N_17078);
nor U17285 (N_17285,N_17171,N_17120);
and U17286 (N_17286,N_17105,N_17049);
nor U17287 (N_17287,N_17006,N_17025);
and U17288 (N_17288,N_17117,N_17218);
and U17289 (N_17289,N_17069,N_17245);
or U17290 (N_17290,N_17061,N_17221);
xnor U17291 (N_17291,N_17163,N_17206);
nand U17292 (N_17292,N_17042,N_17197);
or U17293 (N_17293,N_17108,N_17131);
nand U17294 (N_17294,N_17072,N_17044);
nor U17295 (N_17295,N_17093,N_17162);
and U17296 (N_17296,N_17111,N_17207);
or U17297 (N_17297,N_17051,N_17065);
and U17298 (N_17298,N_17144,N_17248);
nand U17299 (N_17299,N_17150,N_17081);
nand U17300 (N_17300,N_17215,N_17135);
nor U17301 (N_17301,N_17168,N_17238);
nor U17302 (N_17302,N_17041,N_17024);
nand U17303 (N_17303,N_17021,N_17121);
or U17304 (N_17304,N_17022,N_17177);
or U17305 (N_17305,N_17098,N_17018);
or U17306 (N_17306,N_17172,N_17152);
nand U17307 (N_17307,N_17153,N_17158);
or U17308 (N_17308,N_17148,N_17112);
nand U17309 (N_17309,N_17190,N_17211);
or U17310 (N_17310,N_17130,N_17202);
nand U17311 (N_17311,N_17040,N_17205);
and U17312 (N_17312,N_17195,N_17103);
nor U17313 (N_17313,N_17170,N_17070);
nand U17314 (N_17314,N_17128,N_17229);
or U17315 (N_17315,N_17023,N_17189);
or U17316 (N_17316,N_17180,N_17209);
nand U17317 (N_17317,N_17222,N_17090);
nor U17318 (N_17318,N_17030,N_17063);
nor U17319 (N_17319,N_17126,N_17179);
nor U17320 (N_17320,N_17167,N_17165);
nor U17321 (N_17321,N_17247,N_17129);
or U17322 (N_17322,N_17017,N_17210);
nor U17323 (N_17323,N_17242,N_17060);
and U17324 (N_17324,N_17246,N_17031);
or U17325 (N_17325,N_17160,N_17035);
nand U17326 (N_17326,N_17232,N_17198);
nand U17327 (N_17327,N_17146,N_17075);
or U17328 (N_17328,N_17009,N_17054);
nand U17329 (N_17329,N_17187,N_17192);
nor U17330 (N_17330,N_17157,N_17036);
nor U17331 (N_17331,N_17116,N_17122);
and U17332 (N_17332,N_17201,N_17004);
and U17333 (N_17333,N_17235,N_17068);
nor U17334 (N_17334,N_17104,N_17099);
xnor U17335 (N_17335,N_17000,N_17151);
or U17336 (N_17336,N_17097,N_17067);
nand U17337 (N_17337,N_17133,N_17164);
nand U17338 (N_17338,N_17231,N_17203);
and U17339 (N_17339,N_17200,N_17223);
nor U17340 (N_17340,N_17110,N_17124);
and U17341 (N_17341,N_17132,N_17086);
and U17342 (N_17342,N_17216,N_17191);
nor U17343 (N_17343,N_17188,N_17220);
and U17344 (N_17344,N_17239,N_17066);
or U17345 (N_17345,N_17008,N_17196);
or U17346 (N_17346,N_17106,N_17240);
or U17347 (N_17347,N_17199,N_17046);
or U17348 (N_17348,N_17003,N_17001);
nor U17349 (N_17349,N_17010,N_17226);
nor U17350 (N_17350,N_17092,N_17073);
nor U17351 (N_17351,N_17013,N_17045);
nor U17352 (N_17352,N_17243,N_17213);
and U17353 (N_17353,N_17237,N_17241);
nand U17354 (N_17354,N_17186,N_17175);
or U17355 (N_17355,N_17123,N_17088);
xnor U17356 (N_17356,N_17214,N_17181);
nor U17357 (N_17357,N_17027,N_17016);
xor U17358 (N_17358,N_17047,N_17039);
and U17359 (N_17359,N_17095,N_17064);
and U17360 (N_17360,N_17026,N_17011);
or U17361 (N_17361,N_17043,N_17107);
and U17362 (N_17362,N_17155,N_17227);
xnor U17363 (N_17363,N_17166,N_17212);
or U17364 (N_17364,N_17083,N_17204);
and U17365 (N_17365,N_17028,N_17053);
and U17366 (N_17366,N_17156,N_17050);
or U17367 (N_17367,N_17134,N_17169);
or U17368 (N_17368,N_17089,N_17038);
nand U17369 (N_17369,N_17219,N_17094);
or U17370 (N_17370,N_17138,N_17225);
nor U17371 (N_17371,N_17208,N_17224);
xor U17372 (N_17372,N_17076,N_17113);
nand U17373 (N_17373,N_17184,N_17147);
nor U17374 (N_17374,N_17015,N_17228);
and U17375 (N_17375,N_17187,N_17084);
nand U17376 (N_17376,N_17162,N_17096);
xor U17377 (N_17377,N_17176,N_17157);
xnor U17378 (N_17378,N_17219,N_17205);
nor U17379 (N_17379,N_17076,N_17039);
or U17380 (N_17380,N_17108,N_17057);
nor U17381 (N_17381,N_17036,N_17071);
nand U17382 (N_17382,N_17241,N_17131);
and U17383 (N_17383,N_17056,N_17070);
and U17384 (N_17384,N_17217,N_17171);
xor U17385 (N_17385,N_17073,N_17193);
and U17386 (N_17386,N_17188,N_17056);
and U17387 (N_17387,N_17076,N_17091);
xnor U17388 (N_17388,N_17062,N_17189);
or U17389 (N_17389,N_17026,N_17166);
nor U17390 (N_17390,N_17246,N_17139);
nor U17391 (N_17391,N_17095,N_17130);
and U17392 (N_17392,N_17081,N_17044);
xor U17393 (N_17393,N_17129,N_17069);
and U17394 (N_17394,N_17130,N_17049);
or U17395 (N_17395,N_17123,N_17045);
nor U17396 (N_17396,N_17122,N_17114);
and U17397 (N_17397,N_17217,N_17124);
or U17398 (N_17398,N_17118,N_17247);
and U17399 (N_17399,N_17213,N_17019);
nor U17400 (N_17400,N_17011,N_17081);
nand U17401 (N_17401,N_17176,N_17160);
nor U17402 (N_17402,N_17123,N_17030);
and U17403 (N_17403,N_17193,N_17155);
and U17404 (N_17404,N_17185,N_17112);
nor U17405 (N_17405,N_17055,N_17046);
or U17406 (N_17406,N_17088,N_17073);
xnor U17407 (N_17407,N_17177,N_17127);
nor U17408 (N_17408,N_17065,N_17102);
and U17409 (N_17409,N_17127,N_17230);
nor U17410 (N_17410,N_17099,N_17249);
or U17411 (N_17411,N_17223,N_17184);
or U17412 (N_17412,N_17228,N_17233);
and U17413 (N_17413,N_17226,N_17022);
nor U17414 (N_17414,N_17128,N_17221);
nor U17415 (N_17415,N_17045,N_17049);
nor U17416 (N_17416,N_17078,N_17130);
nand U17417 (N_17417,N_17013,N_17187);
xor U17418 (N_17418,N_17164,N_17216);
nor U17419 (N_17419,N_17020,N_17151);
nand U17420 (N_17420,N_17220,N_17059);
xor U17421 (N_17421,N_17009,N_17219);
nor U17422 (N_17422,N_17137,N_17045);
and U17423 (N_17423,N_17051,N_17115);
nand U17424 (N_17424,N_17239,N_17138);
nor U17425 (N_17425,N_17042,N_17192);
or U17426 (N_17426,N_17074,N_17161);
or U17427 (N_17427,N_17033,N_17171);
xor U17428 (N_17428,N_17118,N_17222);
or U17429 (N_17429,N_17095,N_17038);
and U17430 (N_17430,N_17236,N_17232);
and U17431 (N_17431,N_17171,N_17193);
nand U17432 (N_17432,N_17003,N_17242);
or U17433 (N_17433,N_17031,N_17146);
or U17434 (N_17434,N_17157,N_17230);
nand U17435 (N_17435,N_17188,N_17123);
xnor U17436 (N_17436,N_17109,N_17204);
nand U17437 (N_17437,N_17138,N_17028);
or U17438 (N_17438,N_17193,N_17020);
and U17439 (N_17439,N_17077,N_17123);
and U17440 (N_17440,N_17161,N_17070);
nand U17441 (N_17441,N_17197,N_17229);
and U17442 (N_17442,N_17198,N_17028);
and U17443 (N_17443,N_17020,N_17120);
and U17444 (N_17444,N_17012,N_17089);
or U17445 (N_17445,N_17195,N_17139);
nand U17446 (N_17446,N_17213,N_17229);
and U17447 (N_17447,N_17176,N_17167);
nand U17448 (N_17448,N_17088,N_17201);
nor U17449 (N_17449,N_17073,N_17173);
and U17450 (N_17450,N_17087,N_17181);
nand U17451 (N_17451,N_17181,N_17138);
or U17452 (N_17452,N_17175,N_17031);
nor U17453 (N_17453,N_17031,N_17210);
or U17454 (N_17454,N_17090,N_17219);
and U17455 (N_17455,N_17095,N_17086);
nand U17456 (N_17456,N_17192,N_17008);
nor U17457 (N_17457,N_17091,N_17188);
and U17458 (N_17458,N_17201,N_17230);
or U17459 (N_17459,N_17197,N_17239);
nor U17460 (N_17460,N_17005,N_17004);
xor U17461 (N_17461,N_17135,N_17031);
or U17462 (N_17462,N_17142,N_17175);
nand U17463 (N_17463,N_17185,N_17191);
nor U17464 (N_17464,N_17183,N_17083);
and U17465 (N_17465,N_17099,N_17026);
and U17466 (N_17466,N_17037,N_17000);
and U17467 (N_17467,N_17242,N_17155);
or U17468 (N_17468,N_17028,N_17238);
nor U17469 (N_17469,N_17115,N_17245);
or U17470 (N_17470,N_17092,N_17111);
nor U17471 (N_17471,N_17033,N_17071);
or U17472 (N_17472,N_17154,N_17056);
nor U17473 (N_17473,N_17235,N_17029);
xor U17474 (N_17474,N_17138,N_17187);
or U17475 (N_17475,N_17008,N_17112);
nand U17476 (N_17476,N_17185,N_17148);
nor U17477 (N_17477,N_17135,N_17033);
xnor U17478 (N_17478,N_17068,N_17011);
xnor U17479 (N_17479,N_17087,N_17043);
nor U17480 (N_17480,N_17040,N_17033);
nand U17481 (N_17481,N_17037,N_17154);
or U17482 (N_17482,N_17165,N_17209);
nand U17483 (N_17483,N_17017,N_17010);
and U17484 (N_17484,N_17067,N_17076);
or U17485 (N_17485,N_17240,N_17143);
nand U17486 (N_17486,N_17147,N_17046);
and U17487 (N_17487,N_17171,N_17242);
or U17488 (N_17488,N_17151,N_17079);
or U17489 (N_17489,N_17009,N_17240);
nor U17490 (N_17490,N_17094,N_17177);
nand U17491 (N_17491,N_17017,N_17088);
and U17492 (N_17492,N_17096,N_17214);
and U17493 (N_17493,N_17120,N_17240);
nand U17494 (N_17494,N_17048,N_17117);
and U17495 (N_17495,N_17138,N_17111);
and U17496 (N_17496,N_17219,N_17245);
xnor U17497 (N_17497,N_17249,N_17129);
nor U17498 (N_17498,N_17164,N_17121);
nand U17499 (N_17499,N_17142,N_17112);
nand U17500 (N_17500,N_17399,N_17272);
and U17501 (N_17501,N_17306,N_17390);
nor U17502 (N_17502,N_17350,N_17447);
xor U17503 (N_17503,N_17470,N_17253);
nor U17504 (N_17504,N_17268,N_17326);
nand U17505 (N_17505,N_17285,N_17356);
or U17506 (N_17506,N_17265,N_17331);
xor U17507 (N_17507,N_17444,N_17277);
xor U17508 (N_17508,N_17415,N_17389);
nor U17509 (N_17509,N_17370,N_17305);
xor U17510 (N_17510,N_17347,N_17290);
and U17511 (N_17511,N_17288,N_17320);
nor U17512 (N_17512,N_17273,N_17448);
and U17513 (N_17513,N_17426,N_17413);
nand U17514 (N_17514,N_17318,N_17383);
or U17515 (N_17515,N_17374,N_17276);
or U17516 (N_17516,N_17365,N_17393);
and U17517 (N_17517,N_17418,N_17269);
and U17518 (N_17518,N_17385,N_17372);
nand U17519 (N_17519,N_17280,N_17464);
or U17520 (N_17520,N_17299,N_17352);
or U17521 (N_17521,N_17258,N_17403);
xor U17522 (N_17522,N_17298,N_17495);
nand U17523 (N_17523,N_17455,N_17349);
or U17524 (N_17524,N_17364,N_17338);
nand U17525 (N_17525,N_17345,N_17420);
or U17526 (N_17526,N_17437,N_17395);
nor U17527 (N_17527,N_17262,N_17377);
xnor U17528 (N_17528,N_17300,N_17375);
xor U17529 (N_17529,N_17497,N_17368);
and U17530 (N_17530,N_17401,N_17283);
and U17531 (N_17531,N_17266,N_17316);
nand U17532 (N_17532,N_17303,N_17434);
nand U17533 (N_17533,N_17438,N_17348);
and U17534 (N_17534,N_17473,N_17257);
or U17535 (N_17535,N_17427,N_17432);
nand U17536 (N_17536,N_17481,N_17419);
or U17537 (N_17537,N_17446,N_17479);
nor U17538 (N_17538,N_17452,N_17296);
xnor U17539 (N_17539,N_17477,N_17263);
nor U17540 (N_17540,N_17330,N_17400);
nand U17541 (N_17541,N_17450,N_17260);
or U17542 (N_17542,N_17367,N_17471);
nand U17543 (N_17543,N_17256,N_17468);
or U17544 (N_17544,N_17414,N_17484);
or U17545 (N_17545,N_17482,N_17284);
or U17546 (N_17546,N_17371,N_17435);
nand U17547 (N_17547,N_17398,N_17463);
and U17548 (N_17548,N_17255,N_17381);
and U17549 (N_17549,N_17421,N_17328);
or U17550 (N_17550,N_17379,N_17363);
or U17551 (N_17551,N_17384,N_17355);
xnor U17552 (N_17552,N_17281,N_17422);
xor U17553 (N_17553,N_17360,N_17496);
nand U17554 (N_17554,N_17341,N_17394);
or U17555 (N_17555,N_17297,N_17402);
nor U17556 (N_17556,N_17252,N_17287);
nand U17557 (N_17557,N_17357,N_17295);
and U17558 (N_17558,N_17322,N_17314);
nor U17559 (N_17559,N_17325,N_17334);
and U17560 (N_17560,N_17431,N_17445);
or U17561 (N_17561,N_17301,N_17430);
nor U17562 (N_17562,N_17443,N_17472);
or U17563 (N_17563,N_17312,N_17286);
xor U17564 (N_17564,N_17270,N_17485);
xor U17565 (N_17565,N_17336,N_17488);
or U17566 (N_17566,N_17321,N_17441);
or U17567 (N_17567,N_17397,N_17457);
or U17568 (N_17568,N_17289,N_17396);
nor U17569 (N_17569,N_17494,N_17254);
nand U17570 (N_17570,N_17267,N_17456);
and U17571 (N_17571,N_17359,N_17346);
and U17572 (N_17572,N_17311,N_17309);
and U17573 (N_17573,N_17410,N_17475);
nor U17574 (N_17574,N_17264,N_17342);
and U17575 (N_17575,N_17428,N_17308);
nand U17576 (N_17576,N_17275,N_17340);
or U17577 (N_17577,N_17271,N_17492);
nand U17578 (N_17578,N_17442,N_17291);
and U17579 (N_17579,N_17453,N_17404);
or U17580 (N_17580,N_17474,N_17462);
or U17581 (N_17581,N_17467,N_17476);
or U17582 (N_17582,N_17250,N_17391);
nand U17583 (N_17583,N_17405,N_17424);
or U17584 (N_17584,N_17489,N_17292);
nand U17585 (N_17585,N_17408,N_17361);
xor U17586 (N_17586,N_17333,N_17324);
nand U17587 (N_17587,N_17387,N_17366);
or U17588 (N_17588,N_17466,N_17433);
and U17589 (N_17589,N_17440,N_17458);
or U17590 (N_17590,N_17460,N_17351);
or U17591 (N_17591,N_17388,N_17332);
or U17592 (N_17592,N_17353,N_17373);
or U17593 (N_17593,N_17449,N_17259);
nand U17594 (N_17594,N_17327,N_17382);
nor U17595 (N_17595,N_17490,N_17412);
or U17596 (N_17596,N_17251,N_17411);
nand U17597 (N_17597,N_17282,N_17323);
nor U17598 (N_17598,N_17465,N_17354);
nor U17599 (N_17599,N_17469,N_17362);
nand U17600 (N_17600,N_17459,N_17278);
or U17601 (N_17601,N_17343,N_17358);
or U17602 (N_17602,N_17429,N_17416);
or U17603 (N_17603,N_17380,N_17392);
nor U17604 (N_17604,N_17439,N_17313);
and U17605 (N_17605,N_17478,N_17302);
nor U17606 (N_17606,N_17406,N_17261);
or U17607 (N_17607,N_17409,N_17307);
nand U17608 (N_17608,N_17339,N_17317);
nand U17609 (N_17609,N_17378,N_17425);
nand U17610 (N_17610,N_17294,N_17451);
and U17611 (N_17611,N_17376,N_17344);
and U17612 (N_17612,N_17417,N_17436);
nor U17613 (N_17613,N_17369,N_17319);
nor U17614 (N_17614,N_17491,N_17274);
nor U17615 (N_17615,N_17293,N_17461);
nor U17616 (N_17616,N_17480,N_17304);
nand U17617 (N_17617,N_17483,N_17454);
or U17618 (N_17618,N_17329,N_17486);
and U17619 (N_17619,N_17407,N_17335);
or U17620 (N_17620,N_17498,N_17337);
and U17621 (N_17621,N_17310,N_17423);
nand U17622 (N_17622,N_17487,N_17499);
xor U17623 (N_17623,N_17386,N_17279);
nand U17624 (N_17624,N_17315,N_17493);
and U17625 (N_17625,N_17482,N_17330);
or U17626 (N_17626,N_17456,N_17349);
or U17627 (N_17627,N_17459,N_17324);
nor U17628 (N_17628,N_17331,N_17303);
nand U17629 (N_17629,N_17428,N_17407);
nand U17630 (N_17630,N_17314,N_17354);
nor U17631 (N_17631,N_17423,N_17267);
and U17632 (N_17632,N_17480,N_17399);
nand U17633 (N_17633,N_17377,N_17381);
and U17634 (N_17634,N_17342,N_17390);
and U17635 (N_17635,N_17314,N_17447);
nand U17636 (N_17636,N_17401,N_17323);
or U17637 (N_17637,N_17379,N_17365);
and U17638 (N_17638,N_17489,N_17311);
xnor U17639 (N_17639,N_17341,N_17373);
nor U17640 (N_17640,N_17260,N_17411);
or U17641 (N_17641,N_17319,N_17480);
xnor U17642 (N_17642,N_17478,N_17481);
and U17643 (N_17643,N_17383,N_17437);
and U17644 (N_17644,N_17352,N_17375);
or U17645 (N_17645,N_17429,N_17464);
nor U17646 (N_17646,N_17406,N_17450);
nand U17647 (N_17647,N_17269,N_17472);
nand U17648 (N_17648,N_17256,N_17319);
nor U17649 (N_17649,N_17480,N_17409);
or U17650 (N_17650,N_17487,N_17360);
nor U17651 (N_17651,N_17310,N_17419);
and U17652 (N_17652,N_17298,N_17303);
and U17653 (N_17653,N_17265,N_17284);
nor U17654 (N_17654,N_17498,N_17437);
and U17655 (N_17655,N_17326,N_17369);
or U17656 (N_17656,N_17330,N_17305);
xor U17657 (N_17657,N_17492,N_17368);
and U17658 (N_17658,N_17294,N_17495);
and U17659 (N_17659,N_17486,N_17268);
or U17660 (N_17660,N_17258,N_17294);
and U17661 (N_17661,N_17355,N_17412);
nor U17662 (N_17662,N_17321,N_17367);
nand U17663 (N_17663,N_17373,N_17442);
nor U17664 (N_17664,N_17402,N_17426);
and U17665 (N_17665,N_17277,N_17466);
or U17666 (N_17666,N_17390,N_17368);
nand U17667 (N_17667,N_17436,N_17443);
and U17668 (N_17668,N_17254,N_17315);
nand U17669 (N_17669,N_17438,N_17430);
and U17670 (N_17670,N_17329,N_17466);
or U17671 (N_17671,N_17283,N_17264);
and U17672 (N_17672,N_17461,N_17350);
nor U17673 (N_17673,N_17425,N_17426);
or U17674 (N_17674,N_17280,N_17421);
nand U17675 (N_17675,N_17252,N_17344);
nand U17676 (N_17676,N_17498,N_17370);
nor U17677 (N_17677,N_17483,N_17427);
nand U17678 (N_17678,N_17330,N_17437);
or U17679 (N_17679,N_17446,N_17467);
or U17680 (N_17680,N_17376,N_17428);
or U17681 (N_17681,N_17398,N_17317);
xnor U17682 (N_17682,N_17283,N_17479);
nor U17683 (N_17683,N_17276,N_17280);
nor U17684 (N_17684,N_17464,N_17381);
or U17685 (N_17685,N_17356,N_17274);
xnor U17686 (N_17686,N_17294,N_17250);
xnor U17687 (N_17687,N_17453,N_17318);
or U17688 (N_17688,N_17475,N_17478);
or U17689 (N_17689,N_17461,N_17377);
nand U17690 (N_17690,N_17468,N_17314);
nand U17691 (N_17691,N_17311,N_17254);
or U17692 (N_17692,N_17486,N_17321);
nor U17693 (N_17693,N_17255,N_17389);
nand U17694 (N_17694,N_17284,N_17376);
nor U17695 (N_17695,N_17466,N_17458);
or U17696 (N_17696,N_17267,N_17327);
xor U17697 (N_17697,N_17352,N_17404);
xnor U17698 (N_17698,N_17310,N_17305);
nand U17699 (N_17699,N_17331,N_17257);
and U17700 (N_17700,N_17378,N_17254);
nand U17701 (N_17701,N_17493,N_17368);
or U17702 (N_17702,N_17319,N_17412);
xnor U17703 (N_17703,N_17417,N_17471);
and U17704 (N_17704,N_17267,N_17291);
and U17705 (N_17705,N_17377,N_17308);
or U17706 (N_17706,N_17291,N_17412);
or U17707 (N_17707,N_17375,N_17499);
nor U17708 (N_17708,N_17396,N_17389);
or U17709 (N_17709,N_17426,N_17336);
and U17710 (N_17710,N_17387,N_17469);
nand U17711 (N_17711,N_17304,N_17305);
nor U17712 (N_17712,N_17290,N_17478);
nand U17713 (N_17713,N_17447,N_17334);
nor U17714 (N_17714,N_17489,N_17476);
and U17715 (N_17715,N_17282,N_17450);
nand U17716 (N_17716,N_17331,N_17274);
xnor U17717 (N_17717,N_17429,N_17257);
nor U17718 (N_17718,N_17444,N_17299);
and U17719 (N_17719,N_17385,N_17353);
nor U17720 (N_17720,N_17486,N_17276);
nand U17721 (N_17721,N_17478,N_17394);
and U17722 (N_17722,N_17420,N_17383);
xor U17723 (N_17723,N_17263,N_17405);
and U17724 (N_17724,N_17486,N_17255);
or U17725 (N_17725,N_17391,N_17318);
or U17726 (N_17726,N_17463,N_17266);
nor U17727 (N_17727,N_17409,N_17411);
nand U17728 (N_17728,N_17354,N_17415);
nor U17729 (N_17729,N_17372,N_17388);
and U17730 (N_17730,N_17344,N_17359);
and U17731 (N_17731,N_17372,N_17252);
nor U17732 (N_17732,N_17327,N_17409);
nor U17733 (N_17733,N_17496,N_17371);
and U17734 (N_17734,N_17466,N_17450);
and U17735 (N_17735,N_17478,N_17375);
xor U17736 (N_17736,N_17255,N_17318);
nor U17737 (N_17737,N_17489,N_17426);
or U17738 (N_17738,N_17330,N_17393);
and U17739 (N_17739,N_17333,N_17286);
or U17740 (N_17740,N_17340,N_17446);
xor U17741 (N_17741,N_17320,N_17325);
nand U17742 (N_17742,N_17283,N_17351);
or U17743 (N_17743,N_17452,N_17444);
and U17744 (N_17744,N_17425,N_17484);
or U17745 (N_17745,N_17422,N_17442);
nand U17746 (N_17746,N_17344,N_17385);
and U17747 (N_17747,N_17437,N_17274);
nand U17748 (N_17748,N_17454,N_17445);
nor U17749 (N_17749,N_17365,N_17449);
nand U17750 (N_17750,N_17715,N_17682);
nand U17751 (N_17751,N_17728,N_17610);
nor U17752 (N_17752,N_17620,N_17617);
and U17753 (N_17753,N_17675,N_17714);
and U17754 (N_17754,N_17723,N_17525);
and U17755 (N_17755,N_17697,N_17710);
nand U17756 (N_17756,N_17543,N_17551);
nor U17757 (N_17757,N_17571,N_17588);
nand U17758 (N_17758,N_17535,N_17604);
xnor U17759 (N_17759,N_17672,N_17623);
and U17760 (N_17760,N_17502,N_17522);
and U17761 (N_17761,N_17555,N_17547);
and U17762 (N_17762,N_17685,N_17716);
or U17763 (N_17763,N_17625,N_17702);
nor U17764 (N_17764,N_17626,N_17667);
xor U17765 (N_17765,N_17698,N_17506);
xnor U17766 (N_17766,N_17513,N_17524);
or U17767 (N_17767,N_17615,N_17738);
nor U17768 (N_17768,N_17662,N_17735);
and U17769 (N_17769,N_17589,N_17600);
and U17770 (N_17770,N_17621,N_17520);
nand U17771 (N_17771,N_17542,N_17654);
and U17772 (N_17772,N_17597,N_17678);
xnor U17773 (N_17773,N_17544,N_17657);
and U17774 (N_17774,N_17612,N_17700);
nand U17775 (N_17775,N_17648,N_17596);
or U17776 (N_17776,N_17550,N_17580);
or U17777 (N_17777,N_17701,N_17521);
and U17778 (N_17778,N_17512,N_17507);
nor U17779 (N_17779,N_17745,N_17699);
and U17780 (N_17780,N_17640,N_17603);
and U17781 (N_17781,N_17721,N_17691);
xor U17782 (N_17782,N_17684,N_17646);
and U17783 (N_17783,N_17650,N_17594);
and U17784 (N_17784,N_17633,N_17739);
or U17785 (N_17785,N_17537,N_17712);
or U17786 (N_17786,N_17539,N_17747);
nor U17787 (N_17787,N_17643,N_17511);
nor U17788 (N_17788,N_17705,N_17687);
xnor U17789 (N_17789,N_17634,N_17541);
and U17790 (N_17790,N_17618,N_17583);
nand U17791 (N_17791,N_17674,N_17622);
xnor U17792 (N_17792,N_17593,N_17567);
nor U17793 (N_17793,N_17549,N_17530);
xnor U17794 (N_17794,N_17627,N_17501);
or U17795 (N_17795,N_17532,N_17632);
and U17796 (N_17796,N_17740,N_17516);
nor U17797 (N_17797,N_17717,N_17628);
nand U17798 (N_17798,N_17713,N_17693);
nor U17799 (N_17799,N_17584,N_17658);
nand U17800 (N_17800,N_17649,N_17679);
and U17801 (N_17801,N_17565,N_17592);
or U17802 (N_17802,N_17722,N_17686);
nand U17803 (N_17803,N_17670,N_17742);
and U17804 (N_17804,N_17671,N_17732);
or U17805 (N_17805,N_17538,N_17609);
and U17806 (N_17806,N_17585,N_17659);
nand U17807 (N_17807,N_17529,N_17526);
xnor U17808 (N_17808,N_17587,N_17656);
nor U17809 (N_17809,N_17606,N_17719);
nand U17810 (N_17810,N_17653,N_17602);
or U17811 (N_17811,N_17611,N_17720);
xnor U17812 (N_17812,N_17504,N_17639);
or U17813 (N_17813,N_17500,N_17680);
and U17814 (N_17814,N_17560,N_17569);
nor U17815 (N_17815,N_17531,N_17730);
xnor U17816 (N_17816,N_17707,N_17545);
nor U17817 (N_17817,N_17515,N_17665);
nand U17818 (N_17818,N_17737,N_17718);
or U17819 (N_17819,N_17556,N_17708);
nand U17820 (N_17820,N_17561,N_17527);
and U17821 (N_17821,N_17661,N_17651);
xor U17822 (N_17822,N_17688,N_17616);
and U17823 (N_17823,N_17690,N_17505);
nor U17824 (N_17824,N_17663,N_17607);
or U17825 (N_17825,N_17729,N_17562);
nand U17826 (N_17826,N_17553,N_17676);
and U17827 (N_17827,N_17566,N_17608);
nor U17828 (N_17828,N_17664,N_17548);
and U17829 (N_17829,N_17591,N_17647);
or U17830 (N_17830,N_17668,N_17629);
and U17831 (N_17831,N_17533,N_17694);
nand U17832 (N_17832,N_17711,N_17636);
or U17833 (N_17833,N_17637,N_17605);
and U17834 (N_17834,N_17568,N_17540);
nand U17835 (N_17835,N_17695,N_17546);
nand U17836 (N_17836,N_17614,N_17572);
and U17837 (N_17837,N_17576,N_17578);
and U17838 (N_17838,N_17564,N_17523);
nor U17839 (N_17839,N_17724,N_17734);
nand U17840 (N_17840,N_17630,N_17638);
and U17841 (N_17841,N_17704,N_17514);
nand U17842 (N_17842,N_17613,N_17509);
nor U17843 (N_17843,N_17517,N_17631);
and U17844 (N_17844,N_17519,N_17510);
and U17845 (N_17845,N_17645,N_17536);
and U17846 (N_17846,N_17703,N_17641);
nor U17847 (N_17847,N_17534,N_17579);
xor U17848 (N_17848,N_17727,N_17642);
and U17849 (N_17849,N_17528,N_17689);
or U17850 (N_17850,N_17683,N_17744);
nor U17851 (N_17851,N_17660,N_17575);
nor U17852 (N_17852,N_17590,N_17574);
nand U17853 (N_17853,N_17558,N_17552);
nor U17854 (N_17854,N_17673,N_17669);
nor U17855 (N_17855,N_17741,N_17709);
nor U17856 (N_17856,N_17582,N_17746);
nand U17857 (N_17857,N_17559,N_17624);
nand U17858 (N_17858,N_17598,N_17731);
and U17859 (N_17859,N_17554,N_17518);
nor U17860 (N_17860,N_17743,N_17573);
and U17861 (N_17861,N_17503,N_17557);
xnor U17862 (N_17862,N_17749,N_17577);
xor U17863 (N_17863,N_17666,N_17599);
nor U17864 (N_17864,N_17736,N_17696);
and U17865 (N_17865,N_17581,N_17692);
nand U17866 (N_17866,N_17748,N_17725);
nand U17867 (N_17867,N_17570,N_17681);
or U17868 (N_17868,N_17595,N_17619);
nor U17869 (N_17869,N_17635,N_17706);
nor U17870 (N_17870,N_17677,N_17733);
xnor U17871 (N_17871,N_17508,N_17563);
nor U17872 (N_17872,N_17726,N_17655);
or U17873 (N_17873,N_17652,N_17644);
nor U17874 (N_17874,N_17586,N_17601);
nor U17875 (N_17875,N_17510,N_17725);
nand U17876 (N_17876,N_17525,N_17591);
nand U17877 (N_17877,N_17545,N_17682);
nor U17878 (N_17878,N_17557,N_17649);
nand U17879 (N_17879,N_17631,N_17704);
or U17880 (N_17880,N_17646,N_17645);
or U17881 (N_17881,N_17645,N_17609);
or U17882 (N_17882,N_17539,N_17606);
nand U17883 (N_17883,N_17508,N_17740);
nor U17884 (N_17884,N_17748,N_17625);
xor U17885 (N_17885,N_17697,N_17675);
nand U17886 (N_17886,N_17635,N_17516);
and U17887 (N_17887,N_17554,N_17661);
nor U17888 (N_17888,N_17598,N_17727);
nor U17889 (N_17889,N_17542,N_17553);
xnor U17890 (N_17890,N_17606,N_17698);
and U17891 (N_17891,N_17594,N_17620);
xor U17892 (N_17892,N_17576,N_17681);
and U17893 (N_17893,N_17647,N_17563);
or U17894 (N_17894,N_17746,N_17607);
and U17895 (N_17895,N_17696,N_17742);
nor U17896 (N_17896,N_17570,N_17575);
or U17897 (N_17897,N_17542,N_17554);
nor U17898 (N_17898,N_17740,N_17720);
or U17899 (N_17899,N_17682,N_17527);
nand U17900 (N_17900,N_17627,N_17569);
and U17901 (N_17901,N_17703,N_17574);
nand U17902 (N_17902,N_17552,N_17727);
nand U17903 (N_17903,N_17594,N_17666);
nor U17904 (N_17904,N_17563,N_17567);
or U17905 (N_17905,N_17729,N_17730);
and U17906 (N_17906,N_17716,N_17523);
xnor U17907 (N_17907,N_17579,N_17545);
nand U17908 (N_17908,N_17576,N_17732);
or U17909 (N_17909,N_17725,N_17567);
and U17910 (N_17910,N_17710,N_17678);
nor U17911 (N_17911,N_17502,N_17701);
nor U17912 (N_17912,N_17557,N_17585);
nand U17913 (N_17913,N_17514,N_17696);
or U17914 (N_17914,N_17678,N_17682);
xor U17915 (N_17915,N_17650,N_17733);
nand U17916 (N_17916,N_17566,N_17570);
nand U17917 (N_17917,N_17524,N_17561);
xor U17918 (N_17918,N_17699,N_17574);
nor U17919 (N_17919,N_17613,N_17559);
and U17920 (N_17920,N_17728,N_17533);
nand U17921 (N_17921,N_17738,N_17643);
or U17922 (N_17922,N_17679,N_17588);
nor U17923 (N_17923,N_17534,N_17583);
or U17924 (N_17924,N_17671,N_17663);
nand U17925 (N_17925,N_17725,N_17676);
and U17926 (N_17926,N_17628,N_17716);
nor U17927 (N_17927,N_17539,N_17534);
nand U17928 (N_17928,N_17608,N_17714);
nand U17929 (N_17929,N_17504,N_17642);
or U17930 (N_17930,N_17601,N_17518);
and U17931 (N_17931,N_17528,N_17728);
or U17932 (N_17932,N_17633,N_17568);
nor U17933 (N_17933,N_17635,N_17615);
xnor U17934 (N_17934,N_17607,N_17662);
and U17935 (N_17935,N_17504,N_17619);
nor U17936 (N_17936,N_17577,N_17558);
nand U17937 (N_17937,N_17594,N_17612);
or U17938 (N_17938,N_17615,N_17703);
and U17939 (N_17939,N_17686,N_17695);
and U17940 (N_17940,N_17612,N_17731);
and U17941 (N_17941,N_17665,N_17667);
nor U17942 (N_17942,N_17536,N_17641);
and U17943 (N_17943,N_17674,N_17522);
and U17944 (N_17944,N_17535,N_17687);
and U17945 (N_17945,N_17719,N_17627);
nor U17946 (N_17946,N_17589,N_17551);
xnor U17947 (N_17947,N_17569,N_17578);
xnor U17948 (N_17948,N_17674,N_17730);
and U17949 (N_17949,N_17630,N_17601);
or U17950 (N_17950,N_17581,N_17712);
or U17951 (N_17951,N_17640,N_17515);
and U17952 (N_17952,N_17626,N_17523);
nor U17953 (N_17953,N_17510,N_17500);
nor U17954 (N_17954,N_17547,N_17742);
or U17955 (N_17955,N_17687,N_17619);
or U17956 (N_17956,N_17733,N_17679);
and U17957 (N_17957,N_17620,N_17674);
and U17958 (N_17958,N_17657,N_17659);
nand U17959 (N_17959,N_17698,N_17666);
and U17960 (N_17960,N_17594,N_17548);
and U17961 (N_17961,N_17619,N_17749);
or U17962 (N_17962,N_17552,N_17732);
and U17963 (N_17963,N_17591,N_17532);
nor U17964 (N_17964,N_17743,N_17673);
nand U17965 (N_17965,N_17698,N_17596);
xnor U17966 (N_17966,N_17729,N_17644);
and U17967 (N_17967,N_17512,N_17730);
or U17968 (N_17968,N_17678,N_17730);
or U17969 (N_17969,N_17641,N_17635);
or U17970 (N_17970,N_17571,N_17643);
and U17971 (N_17971,N_17584,N_17606);
nor U17972 (N_17972,N_17691,N_17633);
xor U17973 (N_17973,N_17538,N_17549);
or U17974 (N_17974,N_17740,N_17544);
or U17975 (N_17975,N_17700,N_17610);
nand U17976 (N_17976,N_17574,N_17530);
nor U17977 (N_17977,N_17691,N_17603);
nor U17978 (N_17978,N_17595,N_17740);
nor U17979 (N_17979,N_17588,N_17662);
nand U17980 (N_17980,N_17659,N_17678);
xor U17981 (N_17981,N_17696,N_17558);
or U17982 (N_17982,N_17527,N_17648);
xor U17983 (N_17983,N_17624,N_17669);
nor U17984 (N_17984,N_17654,N_17744);
and U17985 (N_17985,N_17599,N_17578);
nor U17986 (N_17986,N_17589,N_17720);
nor U17987 (N_17987,N_17748,N_17516);
xnor U17988 (N_17988,N_17724,N_17606);
or U17989 (N_17989,N_17646,N_17660);
xor U17990 (N_17990,N_17604,N_17595);
and U17991 (N_17991,N_17581,N_17628);
and U17992 (N_17992,N_17689,N_17739);
nand U17993 (N_17993,N_17605,N_17613);
nor U17994 (N_17994,N_17599,N_17589);
or U17995 (N_17995,N_17523,N_17644);
xnor U17996 (N_17996,N_17670,N_17599);
or U17997 (N_17997,N_17583,N_17721);
nand U17998 (N_17998,N_17548,N_17577);
xnor U17999 (N_17999,N_17724,N_17696);
nand U18000 (N_18000,N_17810,N_17880);
and U18001 (N_18001,N_17755,N_17847);
nor U18002 (N_18002,N_17989,N_17835);
nor U18003 (N_18003,N_17815,N_17837);
and U18004 (N_18004,N_17924,N_17881);
xor U18005 (N_18005,N_17927,N_17788);
and U18006 (N_18006,N_17859,N_17852);
nor U18007 (N_18007,N_17857,N_17777);
nand U18008 (N_18008,N_17874,N_17932);
or U18009 (N_18009,N_17866,N_17809);
xor U18010 (N_18010,N_17780,N_17955);
xnor U18011 (N_18011,N_17772,N_17831);
or U18012 (N_18012,N_17877,N_17919);
nor U18013 (N_18013,N_17790,N_17757);
nand U18014 (N_18014,N_17851,N_17762);
xor U18015 (N_18015,N_17822,N_17830);
xor U18016 (N_18016,N_17984,N_17952);
and U18017 (N_18017,N_17977,N_17970);
nor U18018 (N_18018,N_17792,N_17871);
and U18019 (N_18019,N_17933,N_17827);
nor U18020 (N_18020,N_17950,N_17858);
or U18021 (N_18021,N_17825,N_17785);
or U18022 (N_18022,N_17850,N_17818);
and U18023 (N_18023,N_17945,N_17972);
and U18024 (N_18024,N_17943,N_17861);
and U18025 (N_18025,N_17786,N_17946);
or U18026 (N_18026,N_17836,N_17860);
nand U18027 (N_18027,N_17899,N_17969);
nor U18028 (N_18028,N_17968,N_17900);
and U18029 (N_18029,N_17803,N_17804);
or U18030 (N_18030,N_17844,N_17800);
nor U18031 (N_18031,N_17854,N_17855);
nand U18032 (N_18032,N_17940,N_17751);
or U18033 (N_18033,N_17928,N_17816);
nor U18034 (N_18034,N_17795,N_17921);
nor U18035 (N_18035,N_17895,N_17781);
or U18036 (N_18036,N_17753,N_17833);
or U18037 (N_18037,N_17988,N_17886);
xor U18038 (N_18038,N_17965,N_17776);
xor U18039 (N_18039,N_17956,N_17992);
and U18040 (N_18040,N_17962,N_17875);
or U18041 (N_18041,N_17750,N_17820);
nor U18042 (N_18042,N_17996,N_17845);
nor U18043 (N_18043,N_17774,N_17849);
and U18044 (N_18044,N_17915,N_17868);
nand U18045 (N_18045,N_17896,N_17796);
nand U18046 (N_18046,N_17973,N_17769);
xor U18047 (N_18047,N_17913,N_17798);
or U18048 (N_18048,N_17981,N_17839);
or U18049 (N_18049,N_17975,N_17889);
xor U18050 (N_18050,N_17765,N_17791);
or U18051 (N_18051,N_17824,N_17901);
and U18052 (N_18052,N_17879,N_17941);
xnor U18053 (N_18053,N_17997,N_17767);
and U18054 (N_18054,N_17961,N_17812);
nor U18055 (N_18055,N_17920,N_17905);
nor U18056 (N_18056,N_17821,N_17954);
nand U18057 (N_18057,N_17853,N_17906);
nand U18058 (N_18058,N_17763,N_17864);
or U18059 (N_18059,N_17912,N_17971);
nor U18060 (N_18060,N_17843,N_17892);
nor U18061 (N_18061,N_17951,N_17890);
nor U18062 (N_18062,N_17814,N_17967);
nor U18063 (N_18063,N_17957,N_17856);
or U18064 (N_18064,N_17993,N_17797);
and U18065 (N_18065,N_17960,N_17778);
or U18066 (N_18066,N_17888,N_17907);
or U18067 (N_18067,N_17935,N_17916);
and U18068 (N_18068,N_17867,N_17953);
nand U18069 (N_18069,N_17938,N_17817);
nand U18070 (N_18070,N_17761,N_17801);
nand U18071 (N_18071,N_17937,N_17869);
nor U18072 (N_18072,N_17768,N_17841);
xnor U18073 (N_18073,N_17966,N_17991);
nor U18074 (N_18074,N_17986,N_17982);
nand U18075 (N_18075,N_17862,N_17775);
nand U18076 (N_18076,N_17987,N_17829);
nor U18077 (N_18077,N_17995,N_17909);
or U18078 (N_18078,N_17942,N_17799);
or U18079 (N_18079,N_17959,N_17828);
or U18080 (N_18080,N_17936,N_17926);
nand U18081 (N_18081,N_17832,N_17998);
nand U18082 (N_18082,N_17771,N_17923);
nand U18083 (N_18083,N_17902,N_17793);
or U18084 (N_18084,N_17873,N_17976);
or U18085 (N_18085,N_17811,N_17910);
xor U18086 (N_18086,N_17897,N_17949);
or U18087 (N_18087,N_17846,N_17848);
or U18088 (N_18088,N_17948,N_17898);
or U18089 (N_18089,N_17934,N_17783);
and U18090 (N_18090,N_17787,N_17760);
and U18091 (N_18091,N_17929,N_17964);
nor U18092 (N_18092,N_17806,N_17842);
nand U18093 (N_18093,N_17805,N_17930);
or U18094 (N_18094,N_17872,N_17939);
or U18095 (N_18095,N_17882,N_17782);
nor U18096 (N_18096,N_17773,N_17931);
nand U18097 (N_18097,N_17980,N_17887);
nor U18098 (N_18098,N_17994,N_17807);
xor U18099 (N_18099,N_17974,N_17891);
nand U18100 (N_18100,N_17759,N_17802);
xor U18101 (N_18101,N_17983,N_17999);
or U18102 (N_18102,N_17922,N_17978);
or U18103 (N_18103,N_17840,N_17893);
nand U18104 (N_18104,N_17752,N_17764);
or U18105 (N_18105,N_17826,N_17789);
nand U18106 (N_18106,N_17784,N_17770);
xor U18107 (N_18107,N_17838,N_17947);
nor U18108 (N_18108,N_17779,N_17944);
nand U18109 (N_18109,N_17925,N_17894);
or U18110 (N_18110,N_17904,N_17914);
or U18111 (N_18111,N_17903,N_17979);
xnor U18112 (N_18112,N_17758,N_17990);
nand U18113 (N_18113,N_17834,N_17908);
nor U18114 (N_18114,N_17963,N_17884);
xnor U18115 (N_18115,N_17756,N_17918);
or U18116 (N_18116,N_17911,N_17863);
and U18117 (N_18117,N_17878,N_17794);
nor U18118 (N_18118,N_17766,N_17883);
and U18119 (N_18119,N_17917,N_17823);
and U18120 (N_18120,N_17958,N_17813);
nand U18121 (N_18121,N_17808,N_17985);
or U18122 (N_18122,N_17754,N_17819);
xor U18123 (N_18123,N_17870,N_17865);
xor U18124 (N_18124,N_17885,N_17876);
xor U18125 (N_18125,N_17954,N_17792);
nor U18126 (N_18126,N_17957,N_17777);
nor U18127 (N_18127,N_17961,N_17810);
nor U18128 (N_18128,N_17822,N_17929);
or U18129 (N_18129,N_17866,N_17776);
and U18130 (N_18130,N_17972,N_17927);
and U18131 (N_18131,N_17758,N_17813);
nand U18132 (N_18132,N_17946,N_17860);
nand U18133 (N_18133,N_17974,N_17895);
and U18134 (N_18134,N_17798,N_17967);
nor U18135 (N_18135,N_17878,N_17994);
nand U18136 (N_18136,N_17918,N_17852);
and U18137 (N_18137,N_17820,N_17812);
xnor U18138 (N_18138,N_17880,N_17955);
nor U18139 (N_18139,N_17796,N_17952);
nor U18140 (N_18140,N_17879,N_17932);
nor U18141 (N_18141,N_17782,N_17862);
xor U18142 (N_18142,N_17816,N_17955);
or U18143 (N_18143,N_17981,N_17987);
or U18144 (N_18144,N_17895,N_17855);
nand U18145 (N_18145,N_17969,N_17854);
and U18146 (N_18146,N_17939,N_17858);
and U18147 (N_18147,N_17779,N_17810);
nor U18148 (N_18148,N_17931,N_17759);
xnor U18149 (N_18149,N_17817,N_17886);
and U18150 (N_18150,N_17941,N_17959);
or U18151 (N_18151,N_17878,N_17834);
xor U18152 (N_18152,N_17993,N_17812);
or U18153 (N_18153,N_17770,N_17775);
and U18154 (N_18154,N_17754,N_17766);
nand U18155 (N_18155,N_17855,N_17907);
or U18156 (N_18156,N_17969,N_17931);
nor U18157 (N_18157,N_17943,N_17757);
or U18158 (N_18158,N_17818,N_17924);
and U18159 (N_18159,N_17841,N_17968);
and U18160 (N_18160,N_17907,N_17868);
nand U18161 (N_18161,N_17839,N_17760);
nand U18162 (N_18162,N_17899,N_17932);
or U18163 (N_18163,N_17944,N_17881);
or U18164 (N_18164,N_17770,N_17957);
nand U18165 (N_18165,N_17978,N_17885);
and U18166 (N_18166,N_17950,N_17976);
and U18167 (N_18167,N_17934,N_17931);
nor U18168 (N_18168,N_17897,N_17843);
nand U18169 (N_18169,N_17823,N_17843);
or U18170 (N_18170,N_17767,N_17851);
and U18171 (N_18171,N_17751,N_17886);
and U18172 (N_18172,N_17770,N_17857);
or U18173 (N_18173,N_17907,N_17799);
nor U18174 (N_18174,N_17794,N_17830);
and U18175 (N_18175,N_17886,N_17941);
nand U18176 (N_18176,N_17924,N_17878);
nor U18177 (N_18177,N_17948,N_17803);
nor U18178 (N_18178,N_17999,N_17952);
or U18179 (N_18179,N_17950,N_17841);
and U18180 (N_18180,N_17971,N_17882);
and U18181 (N_18181,N_17852,N_17987);
xnor U18182 (N_18182,N_17855,N_17843);
nand U18183 (N_18183,N_17978,N_17848);
nand U18184 (N_18184,N_17895,N_17857);
or U18185 (N_18185,N_17766,N_17887);
nor U18186 (N_18186,N_17925,N_17772);
nor U18187 (N_18187,N_17996,N_17788);
nor U18188 (N_18188,N_17843,N_17816);
nor U18189 (N_18189,N_17803,N_17793);
or U18190 (N_18190,N_17916,N_17943);
and U18191 (N_18191,N_17928,N_17830);
or U18192 (N_18192,N_17909,N_17991);
nor U18193 (N_18193,N_17863,N_17953);
or U18194 (N_18194,N_17794,N_17774);
nor U18195 (N_18195,N_17934,N_17828);
xnor U18196 (N_18196,N_17790,N_17808);
nor U18197 (N_18197,N_17974,N_17859);
and U18198 (N_18198,N_17800,N_17950);
nand U18199 (N_18199,N_17785,N_17919);
xor U18200 (N_18200,N_17821,N_17841);
nand U18201 (N_18201,N_17952,N_17998);
or U18202 (N_18202,N_17764,N_17820);
or U18203 (N_18203,N_17909,N_17839);
nor U18204 (N_18204,N_17958,N_17880);
nor U18205 (N_18205,N_17916,N_17827);
nand U18206 (N_18206,N_17999,N_17896);
or U18207 (N_18207,N_17757,N_17880);
xnor U18208 (N_18208,N_17937,N_17815);
and U18209 (N_18209,N_17922,N_17986);
and U18210 (N_18210,N_17866,N_17934);
xor U18211 (N_18211,N_17906,N_17914);
or U18212 (N_18212,N_17906,N_17784);
nand U18213 (N_18213,N_17916,N_17818);
and U18214 (N_18214,N_17793,N_17844);
nand U18215 (N_18215,N_17785,N_17865);
nand U18216 (N_18216,N_17912,N_17867);
nand U18217 (N_18217,N_17923,N_17775);
or U18218 (N_18218,N_17980,N_17932);
and U18219 (N_18219,N_17990,N_17831);
nor U18220 (N_18220,N_17799,N_17982);
or U18221 (N_18221,N_17860,N_17827);
nor U18222 (N_18222,N_17862,N_17949);
nand U18223 (N_18223,N_17858,N_17807);
and U18224 (N_18224,N_17864,N_17872);
and U18225 (N_18225,N_17854,N_17968);
nor U18226 (N_18226,N_17910,N_17882);
nand U18227 (N_18227,N_17778,N_17822);
and U18228 (N_18228,N_17853,N_17967);
nor U18229 (N_18229,N_17857,N_17883);
or U18230 (N_18230,N_17945,N_17961);
xnor U18231 (N_18231,N_17900,N_17811);
or U18232 (N_18232,N_17880,N_17935);
or U18233 (N_18233,N_17923,N_17784);
and U18234 (N_18234,N_17779,N_17847);
and U18235 (N_18235,N_17888,N_17791);
or U18236 (N_18236,N_17779,N_17835);
nand U18237 (N_18237,N_17855,N_17779);
nand U18238 (N_18238,N_17862,N_17886);
or U18239 (N_18239,N_17848,N_17968);
xor U18240 (N_18240,N_17948,N_17959);
nand U18241 (N_18241,N_17822,N_17932);
nand U18242 (N_18242,N_17995,N_17777);
and U18243 (N_18243,N_17880,N_17783);
nor U18244 (N_18244,N_17954,N_17811);
or U18245 (N_18245,N_17811,N_17932);
or U18246 (N_18246,N_17942,N_17995);
xnor U18247 (N_18247,N_17830,N_17774);
nor U18248 (N_18248,N_17767,N_17883);
and U18249 (N_18249,N_17903,N_17852);
or U18250 (N_18250,N_18221,N_18099);
and U18251 (N_18251,N_18092,N_18117);
nor U18252 (N_18252,N_18125,N_18104);
nor U18253 (N_18253,N_18155,N_18045);
nand U18254 (N_18254,N_18244,N_18066);
nor U18255 (N_18255,N_18138,N_18132);
nand U18256 (N_18256,N_18174,N_18048);
and U18257 (N_18257,N_18004,N_18051);
nor U18258 (N_18258,N_18195,N_18114);
nor U18259 (N_18259,N_18075,N_18223);
nand U18260 (N_18260,N_18178,N_18215);
or U18261 (N_18261,N_18067,N_18192);
xor U18262 (N_18262,N_18007,N_18096);
or U18263 (N_18263,N_18000,N_18231);
and U18264 (N_18264,N_18175,N_18081);
nand U18265 (N_18265,N_18173,N_18182);
nand U18266 (N_18266,N_18163,N_18208);
or U18267 (N_18267,N_18033,N_18124);
and U18268 (N_18268,N_18167,N_18018);
and U18269 (N_18269,N_18006,N_18180);
nor U18270 (N_18270,N_18184,N_18198);
nand U18271 (N_18271,N_18166,N_18013);
nor U18272 (N_18272,N_18064,N_18227);
xnor U18273 (N_18273,N_18226,N_18108);
nor U18274 (N_18274,N_18187,N_18152);
or U18275 (N_18275,N_18194,N_18249);
nor U18276 (N_18276,N_18135,N_18210);
and U18277 (N_18277,N_18070,N_18097);
and U18278 (N_18278,N_18055,N_18023);
nand U18279 (N_18279,N_18188,N_18127);
and U18280 (N_18280,N_18179,N_18161);
and U18281 (N_18281,N_18142,N_18058);
nand U18282 (N_18282,N_18079,N_18086);
or U18283 (N_18283,N_18074,N_18020);
nor U18284 (N_18284,N_18145,N_18060);
and U18285 (N_18285,N_18089,N_18243);
nand U18286 (N_18286,N_18078,N_18168);
nor U18287 (N_18287,N_18091,N_18128);
or U18288 (N_18288,N_18032,N_18062);
and U18289 (N_18289,N_18016,N_18053);
xnor U18290 (N_18290,N_18120,N_18201);
xor U18291 (N_18291,N_18037,N_18131);
nor U18292 (N_18292,N_18042,N_18147);
xnor U18293 (N_18293,N_18030,N_18123);
nand U18294 (N_18294,N_18217,N_18009);
or U18295 (N_18295,N_18071,N_18199);
and U18296 (N_18296,N_18186,N_18214);
and U18297 (N_18297,N_18109,N_18112);
nor U18298 (N_18298,N_18200,N_18111);
or U18299 (N_18299,N_18043,N_18121);
or U18300 (N_18300,N_18100,N_18082);
nand U18301 (N_18301,N_18025,N_18136);
and U18302 (N_18302,N_18151,N_18090);
xor U18303 (N_18303,N_18213,N_18177);
nor U18304 (N_18304,N_18196,N_18130);
nand U18305 (N_18305,N_18170,N_18156);
or U18306 (N_18306,N_18034,N_18229);
nand U18307 (N_18307,N_18176,N_18069);
nand U18308 (N_18308,N_18050,N_18241);
or U18309 (N_18309,N_18087,N_18035);
nor U18310 (N_18310,N_18165,N_18134);
or U18311 (N_18311,N_18040,N_18001);
xnor U18312 (N_18312,N_18218,N_18026);
nor U18313 (N_18313,N_18202,N_18101);
or U18314 (N_18314,N_18206,N_18242);
and U18315 (N_18315,N_18068,N_18028);
nor U18316 (N_18316,N_18162,N_18228);
or U18317 (N_18317,N_18103,N_18240);
and U18318 (N_18318,N_18056,N_18220);
or U18319 (N_18319,N_18005,N_18116);
or U18320 (N_18320,N_18118,N_18222);
nor U18321 (N_18321,N_18185,N_18157);
and U18322 (N_18322,N_18012,N_18015);
nor U18323 (N_18323,N_18235,N_18189);
or U18324 (N_18324,N_18225,N_18137);
or U18325 (N_18325,N_18072,N_18140);
and U18326 (N_18326,N_18230,N_18193);
nand U18327 (N_18327,N_18149,N_18148);
nor U18328 (N_18328,N_18203,N_18164);
and U18329 (N_18329,N_18234,N_18083);
nand U18330 (N_18330,N_18247,N_18139);
nand U18331 (N_18331,N_18224,N_18065);
and U18332 (N_18332,N_18238,N_18047);
or U18333 (N_18333,N_18044,N_18141);
nor U18334 (N_18334,N_18144,N_18031);
and U18335 (N_18335,N_18246,N_18204);
nor U18336 (N_18336,N_18052,N_18098);
nand U18337 (N_18337,N_18014,N_18160);
nand U18338 (N_18338,N_18080,N_18143);
and U18339 (N_18339,N_18190,N_18039);
and U18340 (N_18340,N_18085,N_18245);
nand U18341 (N_18341,N_18094,N_18106);
nand U18342 (N_18342,N_18232,N_18150);
xnor U18343 (N_18343,N_18041,N_18063);
nand U18344 (N_18344,N_18237,N_18054);
nor U18345 (N_18345,N_18146,N_18077);
or U18346 (N_18346,N_18129,N_18107);
nand U18347 (N_18347,N_18236,N_18248);
xor U18348 (N_18348,N_18017,N_18159);
or U18349 (N_18349,N_18171,N_18019);
and U18350 (N_18350,N_18191,N_18183);
or U18351 (N_18351,N_18073,N_18181);
nor U18352 (N_18352,N_18088,N_18084);
nor U18353 (N_18353,N_18126,N_18153);
and U18354 (N_18354,N_18197,N_18057);
xnor U18355 (N_18355,N_18209,N_18022);
nand U18356 (N_18356,N_18095,N_18038);
and U18357 (N_18357,N_18212,N_18002);
or U18358 (N_18358,N_18046,N_18122);
nand U18359 (N_18359,N_18172,N_18211);
and U18360 (N_18360,N_18110,N_18003);
nor U18361 (N_18361,N_18158,N_18219);
nor U18362 (N_18362,N_18115,N_18207);
xor U18363 (N_18363,N_18105,N_18233);
nand U18364 (N_18364,N_18061,N_18113);
nor U18365 (N_18365,N_18029,N_18239);
nand U18366 (N_18366,N_18008,N_18119);
or U18367 (N_18367,N_18024,N_18205);
xor U18368 (N_18368,N_18169,N_18059);
or U18369 (N_18369,N_18021,N_18076);
nand U18370 (N_18370,N_18216,N_18049);
or U18371 (N_18371,N_18093,N_18011);
and U18372 (N_18372,N_18027,N_18102);
or U18373 (N_18373,N_18010,N_18154);
nand U18374 (N_18374,N_18133,N_18036);
or U18375 (N_18375,N_18180,N_18002);
nor U18376 (N_18376,N_18016,N_18215);
nor U18377 (N_18377,N_18107,N_18200);
and U18378 (N_18378,N_18183,N_18066);
or U18379 (N_18379,N_18005,N_18082);
or U18380 (N_18380,N_18092,N_18228);
nor U18381 (N_18381,N_18052,N_18166);
nand U18382 (N_18382,N_18037,N_18064);
and U18383 (N_18383,N_18141,N_18185);
nand U18384 (N_18384,N_18038,N_18193);
nor U18385 (N_18385,N_18034,N_18091);
nand U18386 (N_18386,N_18241,N_18058);
or U18387 (N_18387,N_18000,N_18191);
nand U18388 (N_18388,N_18246,N_18165);
and U18389 (N_18389,N_18175,N_18020);
nor U18390 (N_18390,N_18047,N_18185);
and U18391 (N_18391,N_18016,N_18171);
nor U18392 (N_18392,N_18143,N_18159);
nor U18393 (N_18393,N_18055,N_18002);
and U18394 (N_18394,N_18139,N_18228);
nand U18395 (N_18395,N_18190,N_18060);
nor U18396 (N_18396,N_18224,N_18049);
and U18397 (N_18397,N_18059,N_18164);
xor U18398 (N_18398,N_18010,N_18052);
nand U18399 (N_18399,N_18112,N_18089);
and U18400 (N_18400,N_18231,N_18086);
nand U18401 (N_18401,N_18022,N_18131);
nand U18402 (N_18402,N_18142,N_18226);
or U18403 (N_18403,N_18071,N_18238);
or U18404 (N_18404,N_18063,N_18097);
or U18405 (N_18405,N_18012,N_18135);
nand U18406 (N_18406,N_18023,N_18116);
xor U18407 (N_18407,N_18199,N_18186);
xor U18408 (N_18408,N_18008,N_18069);
xor U18409 (N_18409,N_18210,N_18155);
nor U18410 (N_18410,N_18167,N_18233);
or U18411 (N_18411,N_18249,N_18146);
nand U18412 (N_18412,N_18070,N_18047);
xor U18413 (N_18413,N_18070,N_18233);
or U18414 (N_18414,N_18014,N_18126);
nor U18415 (N_18415,N_18095,N_18249);
or U18416 (N_18416,N_18101,N_18022);
and U18417 (N_18417,N_18034,N_18111);
nand U18418 (N_18418,N_18053,N_18155);
and U18419 (N_18419,N_18204,N_18046);
or U18420 (N_18420,N_18048,N_18123);
or U18421 (N_18421,N_18249,N_18159);
nand U18422 (N_18422,N_18106,N_18018);
xor U18423 (N_18423,N_18229,N_18078);
nand U18424 (N_18424,N_18008,N_18065);
or U18425 (N_18425,N_18020,N_18205);
and U18426 (N_18426,N_18064,N_18094);
and U18427 (N_18427,N_18241,N_18060);
or U18428 (N_18428,N_18170,N_18185);
nor U18429 (N_18429,N_18124,N_18170);
and U18430 (N_18430,N_18053,N_18094);
xnor U18431 (N_18431,N_18208,N_18177);
nor U18432 (N_18432,N_18099,N_18128);
and U18433 (N_18433,N_18036,N_18224);
nor U18434 (N_18434,N_18192,N_18044);
nor U18435 (N_18435,N_18027,N_18208);
and U18436 (N_18436,N_18141,N_18082);
and U18437 (N_18437,N_18193,N_18170);
nand U18438 (N_18438,N_18120,N_18147);
or U18439 (N_18439,N_18130,N_18013);
xnor U18440 (N_18440,N_18166,N_18160);
and U18441 (N_18441,N_18090,N_18207);
or U18442 (N_18442,N_18127,N_18177);
nor U18443 (N_18443,N_18150,N_18031);
nand U18444 (N_18444,N_18146,N_18049);
nor U18445 (N_18445,N_18028,N_18201);
nor U18446 (N_18446,N_18194,N_18239);
or U18447 (N_18447,N_18005,N_18063);
and U18448 (N_18448,N_18049,N_18018);
xor U18449 (N_18449,N_18169,N_18206);
nand U18450 (N_18450,N_18003,N_18195);
or U18451 (N_18451,N_18189,N_18200);
or U18452 (N_18452,N_18018,N_18249);
nor U18453 (N_18453,N_18026,N_18115);
or U18454 (N_18454,N_18149,N_18213);
nand U18455 (N_18455,N_18170,N_18003);
nor U18456 (N_18456,N_18228,N_18246);
and U18457 (N_18457,N_18170,N_18174);
nor U18458 (N_18458,N_18247,N_18109);
nor U18459 (N_18459,N_18031,N_18047);
nor U18460 (N_18460,N_18145,N_18201);
xnor U18461 (N_18461,N_18125,N_18150);
nor U18462 (N_18462,N_18227,N_18010);
or U18463 (N_18463,N_18044,N_18225);
and U18464 (N_18464,N_18147,N_18181);
and U18465 (N_18465,N_18185,N_18182);
xor U18466 (N_18466,N_18065,N_18147);
nor U18467 (N_18467,N_18115,N_18071);
or U18468 (N_18468,N_18057,N_18032);
or U18469 (N_18469,N_18032,N_18137);
xnor U18470 (N_18470,N_18220,N_18180);
xor U18471 (N_18471,N_18050,N_18147);
nand U18472 (N_18472,N_18210,N_18247);
and U18473 (N_18473,N_18028,N_18219);
nand U18474 (N_18474,N_18224,N_18043);
xnor U18475 (N_18475,N_18141,N_18098);
nor U18476 (N_18476,N_18042,N_18170);
and U18477 (N_18477,N_18114,N_18115);
or U18478 (N_18478,N_18195,N_18150);
xor U18479 (N_18479,N_18021,N_18004);
and U18480 (N_18480,N_18032,N_18017);
nand U18481 (N_18481,N_18157,N_18137);
or U18482 (N_18482,N_18173,N_18194);
and U18483 (N_18483,N_18111,N_18175);
nor U18484 (N_18484,N_18242,N_18192);
nand U18485 (N_18485,N_18197,N_18247);
nor U18486 (N_18486,N_18218,N_18236);
or U18487 (N_18487,N_18236,N_18103);
and U18488 (N_18488,N_18213,N_18217);
and U18489 (N_18489,N_18084,N_18110);
and U18490 (N_18490,N_18234,N_18088);
nand U18491 (N_18491,N_18170,N_18012);
and U18492 (N_18492,N_18116,N_18104);
nand U18493 (N_18493,N_18020,N_18241);
nand U18494 (N_18494,N_18163,N_18181);
or U18495 (N_18495,N_18192,N_18200);
nand U18496 (N_18496,N_18072,N_18037);
nand U18497 (N_18497,N_18222,N_18216);
or U18498 (N_18498,N_18075,N_18200);
or U18499 (N_18499,N_18053,N_18123);
and U18500 (N_18500,N_18255,N_18342);
nor U18501 (N_18501,N_18406,N_18370);
and U18502 (N_18502,N_18454,N_18286);
or U18503 (N_18503,N_18392,N_18345);
and U18504 (N_18504,N_18250,N_18312);
xnor U18505 (N_18505,N_18279,N_18377);
nor U18506 (N_18506,N_18446,N_18496);
nor U18507 (N_18507,N_18266,N_18379);
and U18508 (N_18508,N_18398,N_18321);
xor U18509 (N_18509,N_18395,N_18252);
nor U18510 (N_18510,N_18492,N_18347);
nor U18511 (N_18511,N_18360,N_18257);
nand U18512 (N_18512,N_18290,N_18383);
and U18513 (N_18513,N_18339,N_18283);
nand U18514 (N_18514,N_18357,N_18302);
nor U18515 (N_18515,N_18385,N_18336);
or U18516 (N_18516,N_18415,N_18325);
nor U18517 (N_18517,N_18378,N_18344);
nor U18518 (N_18518,N_18437,N_18268);
or U18519 (N_18519,N_18317,N_18326);
nor U18520 (N_18520,N_18396,N_18284);
nor U18521 (N_18521,N_18292,N_18369);
or U18522 (N_18522,N_18341,N_18427);
nand U18523 (N_18523,N_18265,N_18289);
nor U18524 (N_18524,N_18447,N_18306);
or U18525 (N_18525,N_18382,N_18470);
xor U18526 (N_18526,N_18333,N_18424);
nor U18527 (N_18527,N_18494,N_18272);
nor U18528 (N_18528,N_18411,N_18429);
or U18529 (N_18529,N_18493,N_18423);
nor U18530 (N_18530,N_18460,N_18376);
and U18531 (N_18531,N_18480,N_18295);
nor U18532 (N_18532,N_18461,N_18416);
nand U18533 (N_18533,N_18452,N_18335);
nand U18534 (N_18534,N_18439,N_18402);
or U18535 (N_18535,N_18456,N_18485);
nor U18536 (N_18536,N_18418,N_18412);
or U18537 (N_18537,N_18450,N_18403);
or U18538 (N_18538,N_18466,N_18278);
nand U18539 (N_18539,N_18261,N_18404);
and U18540 (N_18540,N_18274,N_18414);
and U18541 (N_18541,N_18401,N_18331);
nor U18542 (N_18542,N_18388,N_18288);
and U18543 (N_18543,N_18354,N_18374);
nor U18544 (N_18544,N_18459,N_18353);
nand U18545 (N_18545,N_18386,N_18256);
or U18546 (N_18546,N_18408,N_18371);
nor U18547 (N_18547,N_18430,N_18313);
or U18548 (N_18548,N_18343,N_18359);
nor U18549 (N_18549,N_18328,N_18293);
and U18550 (N_18550,N_18294,N_18332);
nand U18551 (N_18551,N_18356,N_18267);
or U18552 (N_18552,N_18463,N_18348);
nor U18553 (N_18553,N_18434,N_18445);
and U18554 (N_18554,N_18276,N_18413);
nor U18555 (N_18555,N_18490,N_18471);
nand U18556 (N_18556,N_18375,N_18472);
nor U18557 (N_18557,N_18393,N_18462);
nor U18558 (N_18558,N_18428,N_18489);
nand U18559 (N_18559,N_18482,N_18422);
or U18560 (N_18560,N_18327,N_18330);
or U18561 (N_18561,N_18491,N_18442);
nand U18562 (N_18562,N_18270,N_18253);
nor U18563 (N_18563,N_18475,N_18373);
or U18564 (N_18564,N_18487,N_18458);
nand U18565 (N_18565,N_18483,N_18363);
or U18566 (N_18566,N_18259,N_18387);
nor U18567 (N_18567,N_18477,N_18469);
xor U18568 (N_18568,N_18320,N_18337);
and U18569 (N_18569,N_18441,N_18263);
or U18570 (N_18570,N_18285,N_18486);
nand U18571 (N_18571,N_18417,N_18419);
nand U18572 (N_18572,N_18298,N_18262);
nor U18573 (N_18573,N_18291,N_18425);
xor U18574 (N_18574,N_18399,N_18436);
and U18575 (N_18575,N_18304,N_18323);
and U18576 (N_18576,N_18432,N_18346);
nand U18577 (N_18577,N_18473,N_18449);
nor U18578 (N_18578,N_18394,N_18340);
and U18579 (N_18579,N_18438,N_18364);
nand U18580 (N_18580,N_18451,N_18301);
xnor U18581 (N_18581,N_18499,N_18440);
nor U18582 (N_18582,N_18431,N_18453);
nand U18583 (N_18583,N_18433,N_18297);
xnor U18584 (N_18584,N_18300,N_18350);
nor U18585 (N_18585,N_18361,N_18315);
nand U18586 (N_18586,N_18352,N_18384);
and U18587 (N_18587,N_18366,N_18324);
nor U18588 (N_18588,N_18319,N_18264);
nand U18589 (N_18589,N_18474,N_18421);
nor U18590 (N_18590,N_18381,N_18351);
nand U18591 (N_18591,N_18380,N_18362);
nor U18592 (N_18592,N_18355,N_18299);
or U18593 (N_18593,N_18467,N_18251);
nor U18594 (N_18594,N_18281,N_18308);
or U18595 (N_18595,N_18254,N_18495);
nand U18596 (N_18596,N_18296,N_18368);
nor U18597 (N_18597,N_18271,N_18329);
and U18598 (N_18598,N_18407,N_18307);
nand U18599 (N_18599,N_18468,N_18318);
and U18600 (N_18600,N_18465,N_18273);
or U18601 (N_18601,N_18479,N_18338);
and U18602 (N_18602,N_18372,N_18277);
nand U18603 (N_18603,N_18310,N_18334);
xnor U18604 (N_18604,N_18309,N_18269);
or U18605 (N_18605,N_18275,N_18457);
and U18606 (N_18606,N_18280,N_18409);
nand U18607 (N_18607,N_18311,N_18455);
or U18608 (N_18608,N_18484,N_18405);
nand U18609 (N_18609,N_18367,N_18488);
xnor U18610 (N_18610,N_18358,N_18481);
nand U18611 (N_18611,N_18389,N_18497);
nand U18612 (N_18612,N_18303,N_18365);
and U18613 (N_18613,N_18316,N_18478);
nor U18614 (N_18614,N_18322,N_18443);
and U18615 (N_18615,N_18287,N_18426);
nor U18616 (N_18616,N_18390,N_18314);
nor U18617 (N_18617,N_18349,N_18444);
and U18618 (N_18618,N_18420,N_18435);
xnor U18619 (N_18619,N_18282,N_18498);
nand U18620 (N_18620,N_18476,N_18391);
nor U18621 (N_18621,N_18400,N_18258);
and U18622 (N_18622,N_18464,N_18448);
nor U18623 (N_18623,N_18410,N_18305);
nand U18624 (N_18624,N_18260,N_18397);
or U18625 (N_18625,N_18368,N_18340);
nor U18626 (N_18626,N_18332,N_18368);
nor U18627 (N_18627,N_18491,N_18251);
or U18628 (N_18628,N_18449,N_18435);
nand U18629 (N_18629,N_18403,N_18446);
nand U18630 (N_18630,N_18439,N_18455);
nand U18631 (N_18631,N_18392,N_18449);
nor U18632 (N_18632,N_18462,N_18390);
and U18633 (N_18633,N_18376,N_18428);
and U18634 (N_18634,N_18325,N_18291);
xor U18635 (N_18635,N_18421,N_18400);
nor U18636 (N_18636,N_18277,N_18286);
or U18637 (N_18637,N_18458,N_18336);
nand U18638 (N_18638,N_18498,N_18382);
xnor U18639 (N_18639,N_18387,N_18451);
nand U18640 (N_18640,N_18271,N_18458);
nand U18641 (N_18641,N_18483,N_18346);
or U18642 (N_18642,N_18460,N_18332);
nand U18643 (N_18643,N_18390,N_18367);
and U18644 (N_18644,N_18408,N_18459);
nand U18645 (N_18645,N_18252,N_18331);
nor U18646 (N_18646,N_18308,N_18443);
nand U18647 (N_18647,N_18417,N_18496);
and U18648 (N_18648,N_18496,N_18364);
nand U18649 (N_18649,N_18302,N_18476);
or U18650 (N_18650,N_18488,N_18429);
xnor U18651 (N_18651,N_18444,N_18272);
nor U18652 (N_18652,N_18451,N_18275);
nor U18653 (N_18653,N_18428,N_18492);
and U18654 (N_18654,N_18404,N_18447);
xor U18655 (N_18655,N_18350,N_18370);
nand U18656 (N_18656,N_18385,N_18484);
nor U18657 (N_18657,N_18366,N_18255);
nor U18658 (N_18658,N_18383,N_18440);
xnor U18659 (N_18659,N_18477,N_18384);
or U18660 (N_18660,N_18352,N_18288);
or U18661 (N_18661,N_18433,N_18319);
or U18662 (N_18662,N_18371,N_18469);
nor U18663 (N_18663,N_18473,N_18307);
nor U18664 (N_18664,N_18324,N_18281);
or U18665 (N_18665,N_18263,N_18322);
nand U18666 (N_18666,N_18450,N_18269);
xor U18667 (N_18667,N_18487,N_18350);
xor U18668 (N_18668,N_18289,N_18497);
or U18669 (N_18669,N_18368,N_18258);
or U18670 (N_18670,N_18463,N_18331);
nor U18671 (N_18671,N_18388,N_18464);
and U18672 (N_18672,N_18349,N_18337);
nand U18673 (N_18673,N_18496,N_18343);
and U18674 (N_18674,N_18391,N_18298);
or U18675 (N_18675,N_18311,N_18255);
nor U18676 (N_18676,N_18378,N_18440);
nor U18677 (N_18677,N_18282,N_18447);
and U18678 (N_18678,N_18349,N_18288);
and U18679 (N_18679,N_18409,N_18484);
and U18680 (N_18680,N_18254,N_18348);
nand U18681 (N_18681,N_18443,N_18409);
nand U18682 (N_18682,N_18345,N_18393);
xnor U18683 (N_18683,N_18388,N_18483);
and U18684 (N_18684,N_18478,N_18292);
nor U18685 (N_18685,N_18280,N_18404);
and U18686 (N_18686,N_18466,N_18379);
and U18687 (N_18687,N_18378,N_18360);
nand U18688 (N_18688,N_18466,N_18342);
or U18689 (N_18689,N_18457,N_18263);
nand U18690 (N_18690,N_18426,N_18425);
and U18691 (N_18691,N_18385,N_18276);
and U18692 (N_18692,N_18395,N_18306);
and U18693 (N_18693,N_18426,N_18358);
nor U18694 (N_18694,N_18332,N_18342);
nand U18695 (N_18695,N_18289,N_18446);
nor U18696 (N_18696,N_18495,N_18462);
xor U18697 (N_18697,N_18376,N_18489);
nor U18698 (N_18698,N_18257,N_18454);
nor U18699 (N_18699,N_18289,N_18366);
or U18700 (N_18700,N_18490,N_18358);
nor U18701 (N_18701,N_18462,N_18420);
or U18702 (N_18702,N_18399,N_18453);
and U18703 (N_18703,N_18447,N_18349);
nor U18704 (N_18704,N_18271,N_18457);
nor U18705 (N_18705,N_18485,N_18454);
or U18706 (N_18706,N_18334,N_18273);
xnor U18707 (N_18707,N_18271,N_18311);
nor U18708 (N_18708,N_18367,N_18418);
nand U18709 (N_18709,N_18485,N_18433);
and U18710 (N_18710,N_18382,N_18406);
and U18711 (N_18711,N_18324,N_18315);
nor U18712 (N_18712,N_18397,N_18251);
or U18713 (N_18713,N_18381,N_18356);
or U18714 (N_18714,N_18349,N_18498);
or U18715 (N_18715,N_18464,N_18428);
nand U18716 (N_18716,N_18463,N_18400);
nand U18717 (N_18717,N_18359,N_18391);
nor U18718 (N_18718,N_18340,N_18250);
and U18719 (N_18719,N_18436,N_18268);
and U18720 (N_18720,N_18362,N_18425);
nand U18721 (N_18721,N_18412,N_18292);
nor U18722 (N_18722,N_18295,N_18357);
nand U18723 (N_18723,N_18487,N_18345);
nand U18724 (N_18724,N_18453,N_18472);
nand U18725 (N_18725,N_18323,N_18496);
and U18726 (N_18726,N_18402,N_18396);
nor U18727 (N_18727,N_18451,N_18336);
nand U18728 (N_18728,N_18407,N_18415);
xor U18729 (N_18729,N_18276,N_18272);
nor U18730 (N_18730,N_18472,N_18471);
nor U18731 (N_18731,N_18423,N_18337);
and U18732 (N_18732,N_18334,N_18437);
or U18733 (N_18733,N_18263,N_18290);
nor U18734 (N_18734,N_18301,N_18304);
nor U18735 (N_18735,N_18394,N_18320);
and U18736 (N_18736,N_18499,N_18353);
nor U18737 (N_18737,N_18316,N_18317);
nand U18738 (N_18738,N_18279,N_18330);
nand U18739 (N_18739,N_18352,N_18287);
and U18740 (N_18740,N_18259,N_18430);
nand U18741 (N_18741,N_18374,N_18342);
nor U18742 (N_18742,N_18349,N_18321);
nor U18743 (N_18743,N_18403,N_18267);
nand U18744 (N_18744,N_18343,N_18440);
nor U18745 (N_18745,N_18456,N_18310);
nand U18746 (N_18746,N_18301,N_18422);
and U18747 (N_18747,N_18289,N_18293);
xor U18748 (N_18748,N_18255,N_18322);
nor U18749 (N_18749,N_18438,N_18334);
xor U18750 (N_18750,N_18706,N_18616);
nand U18751 (N_18751,N_18739,N_18705);
nor U18752 (N_18752,N_18684,N_18698);
nand U18753 (N_18753,N_18552,N_18649);
nand U18754 (N_18754,N_18663,N_18590);
nand U18755 (N_18755,N_18719,N_18716);
or U18756 (N_18756,N_18650,N_18559);
or U18757 (N_18757,N_18621,N_18626);
nor U18758 (N_18758,N_18516,N_18712);
and U18759 (N_18759,N_18628,N_18566);
and U18760 (N_18760,N_18581,N_18704);
nand U18761 (N_18761,N_18667,N_18583);
or U18762 (N_18762,N_18724,N_18518);
or U18763 (N_18763,N_18665,N_18611);
nand U18764 (N_18764,N_18620,N_18553);
or U18765 (N_18765,N_18609,N_18554);
nand U18766 (N_18766,N_18722,N_18575);
and U18767 (N_18767,N_18668,N_18652);
or U18768 (N_18768,N_18746,N_18714);
and U18769 (N_18769,N_18571,N_18504);
xnor U18770 (N_18770,N_18721,N_18735);
nand U18771 (N_18771,N_18588,N_18658);
or U18772 (N_18772,N_18615,N_18531);
nand U18773 (N_18773,N_18744,N_18550);
xnor U18774 (N_18774,N_18634,N_18689);
xor U18775 (N_18775,N_18709,N_18597);
nand U18776 (N_18776,N_18748,N_18688);
and U18777 (N_18777,N_18717,N_18514);
or U18778 (N_18778,N_18501,N_18521);
xnor U18779 (N_18779,N_18573,N_18731);
nand U18780 (N_18780,N_18636,N_18745);
nand U18781 (N_18781,N_18655,N_18738);
nor U18782 (N_18782,N_18619,N_18586);
nor U18783 (N_18783,N_18508,N_18700);
or U18784 (N_18784,N_18557,N_18677);
nand U18785 (N_18785,N_18718,N_18682);
nor U18786 (N_18786,N_18733,N_18506);
or U18787 (N_18787,N_18708,N_18728);
or U18788 (N_18788,N_18568,N_18535);
nor U18789 (N_18789,N_18533,N_18574);
and U18790 (N_18790,N_18690,N_18502);
and U18791 (N_18791,N_18599,N_18605);
nand U18792 (N_18792,N_18522,N_18529);
or U18793 (N_18793,N_18530,N_18577);
or U18794 (N_18794,N_18743,N_18528);
and U18795 (N_18795,N_18676,N_18653);
or U18796 (N_18796,N_18726,N_18725);
nand U18797 (N_18797,N_18623,N_18582);
or U18798 (N_18798,N_18596,N_18641);
or U18799 (N_18799,N_18657,N_18606);
nand U18800 (N_18800,N_18694,N_18610);
or U18801 (N_18801,N_18699,N_18526);
nor U18802 (N_18802,N_18720,N_18578);
nor U18803 (N_18803,N_18618,N_18622);
or U18804 (N_18804,N_18598,N_18512);
xnor U18805 (N_18805,N_18685,N_18642);
nand U18806 (N_18806,N_18584,N_18695);
and U18807 (N_18807,N_18569,N_18587);
or U18808 (N_18808,N_18540,N_18555);
nor U18809 (N_18809,N_18683,N_18696);
nand U18810 (N_18810,N_18643,N_18702);
nor U18811 (N_18811,N_18585,N_18503);
or U18812 (N_18812,N_18637,N_18507);
nand U18813 (N_18813,N_18707,N_18551);
nor U18814 (N_18814,N_18638,N_18669);
nand U18815 (N_18815,N_18564,N_18654);
and U18816 (N_18816,N_18513,N_18670);
or U18817 (N_18817,N_18749,N_18693);
or U18818 (N_18818,N_18567,N_18608);
nand U18819 (N_18819,N_18659,N_18520);
nand U18820 (N_18820,N_18539,N_18523);
nor U18821 (N_18821,N_18664,N_18614);
nor U18822 (N_18822,N_18730,N_18524);
nor U18823 (N_18823,N_18612,N_18644);
and U18824 (N_18824,N_18736,N_18661);
or U18825 (N_18825,N_18589,N_18572);
nor U18826 (N_18826,N_18701,N_18673);
nor U18827 (N_18827,N_18604,N_18660);
xor U18828 (N_18828,N_18505,N_18633);
xnor U18829 (N_18829,N_18556,N_18687);
nor U18830 (N_18830,N_18629,N_18713);
xor U18831 (N_18831,N_18625,N_18692);
and U18832 (N_18832,N_18500,N_18647);
nor U18833 (N_18833,N_18675,N_18635);
xor U18834 (N_18834,N_18576,N_18517);
nor U18835 (N_18835,N_18681,N_18729);
nand U18836 (N_18836,N_18594,N_18562);
or U18837 (N_18837,N_18640,N_18666);
or U18838 (N_18838,N_18563,N_18593);
and U18839 (N_18839,N_18710,N_18648);
nor U18840 (N_18840,N_18591,N_18607);
or U18841 (N_18841,N_18561,N_18645);
nand U18842 (N_18842,N_18727,N_18541);
or U18843 (N_18843,N_18543,N_18715);
and U18844 (N_18844,N_18509,N_18592);
nand U18845 (N_18845,N_18536,N_18532);
nand U18846 (N_18846,N_18601,N_18651);
xnor U18847 (N_18847,N_18519,N_18613);
and U18848 (N_18848,N_18680,N_18742);
nor U18849 (N_18849,N_18617,N_18525);
nand U18850 (N_18850,N_18595,N_18627);
nand U18851 (N_18851,N_18737,N_18734);
or U18852 (N_18852,N_18631,N_18630);
and U18853 (N_18853,N_18741,N_18678);
or U18854 (N_18854,N_18679,N_18639);
xor U18855 (N_18855,N_18686,N_18671);
xor U18856 (N_18856,N_18542,N_18548);
nand U18857 (N_18857,N_18534,N_18602);
nor U18858 (N_18858,N_18674,N_18703);
nand U18859 (N_18859,N_18632,N_18656);
or U18860 (N_18860,N_18515,N_18527);
nand U18861 (N_18861,N_18697,N_18580);
and U18862 (N_18862,N_18538,N_18570);
or U18863 (N_18863,N_18547,N_18723);
xnor U18864 (N_18864,N_18545,N_18662);
or U18865 (N_18865,N_18511,N_18603);
nand U18866 (N_18866,N_18546,N_18565);
or U18867 (N_18867,N_18579,N_18740);
and U18868 (N_18868,N_18560,N_18747);
and U18869 (N_18869,N_18732,N_18600);
xor U18870 (N_18870,N_18510,N_18691);
nand U18871 (N_18871,N_18646,N_18711);
nand U18872 (N_18872,N_18672,N_18537);
xor U18873 (N_18873,N_18549,N_18558);
xnor U18874 (N_18874,N_18544,N_18624);
nand U18875 (N_18875,N_18593,N_18614);
nor U18876 (N_18876,N_18666,N_18585);
or U18877 (N_18877,N_18662,N_18710);
xor U18878 (N_18878,N_18698,N_18521);
and U18879 (N_18879,N_18629,N_18609);
nor U18880 (N_18880,N_18743,N_18679);
or U18881 (N_18881,N_18699,N_18586);
nor U18882 (N_18882,N_18702,N_18642);
xor U18883 (N_18883,N_18734,N_18667);
or U18884 (N_18884,N_18693,N_18709);
nor U18885 (N_18885,N_18530,N_18629);
xnor U18886 (N_18886,N_18625,N_18633);
nand U18887 (N_18887,N_18725,N_18744);
nand U18888 (N_18888,N_18723,N_18509);
and U18889 (N_18889,N_18680,N_18728);
and U18890 (N_18890,N_18701,N_18615);
and U18891 (N_18891,N_18569,N_18609);
and U18892 (N_18892,N_18666,N_18650);
nand U18893 (N_18893,N_18710,N_18615);
nor U18894 (N_18894,N_18510,N_18644);
and U18895 (N_18895,N_18622,N_18700);
and U18896 (N_18896,N_18730,N_18699);
nand U18897 (N_18897,N_18664,N_18507);
nor U18898 (N_18898,N_18713,N_18510);
and U18899 (N_18899,N_18586,N_18583);
nand U18900 (N_18900,N_18713,N_18705);
and U18901 (N_18901,N_18513,N_18574);
nand U18902 (N_18902,N_18568,N_18554);
or U18903 (N_18903,N_18723,N_18719);
or U18904 (N_18904,N_18625,N_18503);
nor U18905 (N_18905,N_18621,N_18652);
nand U18906 (N_18906,N_18703,N_18684);
and U18907 (N_18907,N_18544,N_18564);
and U18908 (N_18908,N_18749,N_18587);
and U18909 (N_18909,N_18672,N_18600);
nor U18910 (N_18910,N_18632,N_18589);
nand U18911 (N_18911,N_18660,N_18729);
xnor U18912 (N_18912,N_18706,N_18737);
nand U18913 (N_18913,N_18519,N_18697);
nor U18914 (N_18914,N_18743,N_18533);
and U18915 (N_18915,N_18538,N_18660);
or U18916 (N_18916,N_18588,N_18546);
and U18917 (N_18917,N_18636,N_18603);
nand U18918 (N_18918,N_18582,N_18741);
or U18919 (N_18919,N_18624,N_18727);
xnor U18920 (N_18920,N_18679,N_18509);
and U18921 (N_18921,N_18656,N_18500);
and U18922 (N_18922,N_18739,N_18699);
nor U18923 (N_18923,N_18502,N_18685);
nor U18924 (N_18924,N_18503,N_18718);
xnor U18925 (N_18925,N_18543,N_18580);
nand U18926 (N_18926,N_18560,N_18568);
nor U18927 (N_18927,N_18666,N_18592);
xor U18928 (N_18928,N_18580,N_18512);
nand U18929 (N_18929,N_18537,N_18556);
and U18930 (N_18930,N_18592,N_18676);
nand U18931 (N_18931,N_18521,N_18696);
nor U18932 (N_18932,N_18506,N_18566);
nand U18933 (N_18933,N_18624,N_18519);
or U18934 (N_18934,N_18521,N_18646);
and U18935 (N_18935,N_18747,N_18507);
and U18936 (N_18936,N_18501,N_18657);
and U18937 (N_18937,N_18602,N_18563);
and U18938 (N_18938,N_18586,N_18616);
nor U18939 (N_18939,N_18747,N_18527);
nand U18940 (N_18940,N_18594,N_18699);
nand U18941 (N_18941,N_18548,N_18618);
and U18942 (N_18942,N_18582,N_18693);
nand U18943 (N_18943,N_18625,N_18561);
nand U18944 (N_18944,N_18665,N_18673);
or U18945 (N_18945,N_18638,N_18528);
nor U18946 (N_18946,N_18666,N_18655);
xnor U18947 (N_18947,N_18502,N_18615);
or U18948 (N_18948,N_18730,N_18577);
or U18949 (N_18949,N_18703,N_18504);
nor U18950 (N_18950,N_18507,N_18640);
nand U18951 (N_18951,N_18662,N_18742);
or U18952 (N_18952,N_18505,N_18724);
and U18953 (N_18953,N_18643,N_18503);
and U18954 (N_18954,N_18533,N_18706);
nand U18955 (N_18955,N_18525,N_18556);
and U18956 (N_18956,N_18651,N_18540);
nor U18957 (N_18957,N_18607,N_18604);
or U18958 (N_18958,N_18619,N_18674);
nand U18959 (N_18959,N_18732,N_18548);
and U18960 (N_18960,N_18685,N_18527);
xor U18961 (N_18961,N_18539,N_18719);
nor U18962 (N_18962,N_18510,N_18509);
or U18963 (N_18963,N_18547,N_18711);
xor U18964 (N_18964,N_18556,N_18630);
nand U18965 (N_18965,N_18693,N_18520);
and U18966 (N_18966,N_18595,N_18571);
or U18967 (N_18967,N_18516,N_18550);
or U18968 (N_18968,N_18544,N_18575);
and U18969 (N_18969,N_18618,N_18691);
nor U18970 (N_18970,N_18563,N_18553);
nand U18971 (N_18971,N_18528,N_18538);
nand U18972 (N_18972,N_18714,N_18736);
nand U18973 (N_18973,N_18606,N_18594);
or U18974 (N_18974,N_18556,N_18677);
or U18975 (N_18975,N_18745,N_18510);
nand U18976 (N_18976,N_18518,N_18500);
nor U18977 (N_18977,N_18714,N_18544);
or U18978 (N_18978,N_18651,N_18512);
nor U18979 (N_18979,N_18656,N_18674);
nor U18980 (N_18980,N_18580,N_18668);
and U18981 (N_18981,N_18676,N_18518);
nand U18982 (N_18982,N_18695,N_18688);
nor U18983 (N_18983,N_18525,N_18635);
or U18984 (N_18984,N_18733,N_18522);
nor U18985 (N_18985,N_18627,N_18515);
or U18986 (N_18986,N_18718,N_18613);
nor U18987 (N_18987,N_18749,N_18545);
or U18988 (N_18988,N_18672,N_18519);
xor U18989 (N_18989,N_18700,N_18684);
nand U18990 (N_18990,N_18706,N_18511);
and U18991 (N_18991,N_18576,N_18610);
and U18992 (N_18992,N_18722,N_18534);
or U18993 (N_18993,N_18588,N_18729);
nand U18994 (N_18994,N_18745,N_18686);
xnor U18995 (N_18995,N_18639,N_18525);
nor U18996 (N_18996,N_18688,N_18653);
nor U18997 (N_18997,N_18568,N_18587);
and U18998 (N_18998,N_18744,N_18569);
or U18999 (N_18999,N_18662,N_18613);
xor U19000 (N_19000,N_18759,N_18955);
or U19001 (N_19001,N_18842,N_18905);
nor U19002 (N_19002,N_18962,N_18879);
or U19003 (N_19003,N_18979,N_18788);
and U19004 (N_19004,N_18907,N_18755);
xnor U19005 (N_19005,N_18976,N_18901);
and U19006 (N_19006,N_18806,N_18751);
nor U19007 (N_19007,N_18822,N_18963);
nand U19008 (N_19008,N_18969,N_18951);
and U19009 (N_19009,N_18770,N_18990);
xor U19010 (N_19010,N_18884,N_18880);
nand U19011 (N_19011,N_18872,N_18996);
nor U19012 (N_19012,N_18787,N_18946);
and U19013 (N_19013,N_18863,N_18851);
or U19014 (N_19014,N_18906,N_18839);
or U19015 (N_19015,N_18950,N_18958);
and U19016 (N_19016,N_18892,N_18853);
nand U19017 (N_19017,N_18888,N_18940);
or U19018 (N_19018,N_18846,N_18778);
or U19019 (N_19019,N_18840,N_18970);
nor U19020 (N_19020,N_18924,N_18843);
and U19021 (N_19021,N_18855,N_18952);
nand U19022 (N_19022,N_18966,N_18804);
nand U19023 (N_19023,N_18761,N_18774);
nor U19024 (N_19024,N_18868,N_18988);
nor U19025 (N_19025,N_18753,N_18783);
xor U19026 (N_19026,N_18964,N_18781);
xor U19027 (N_19027,N_18800,N_18847);
and U19028 (N_19028,N_18827,N_18848);
and U19029 (N_19029,N_18998,N_18796);
nor U19030 (N_19030,N_18815,N_18967);
or U19031 (N_19031,N_18866,N_18959);
nand U19032 (N_19032,N_18895,N_18993);
and U19033 (N_19033,N_18826,N_18914);
nor U19034 (N_19034,N_18909,N_18776);
nand U19035 (N_19035,N_18797,N_18831);
nor U19036 (N_19036,N_18999,N_18852);
or U19037 (N_19037,N_18937,N_18771);
or U19038 (N_19038,N_18881,N_18968);
and U19039 (N_19039,N_18792,N_18899);
or U19040 (N_19040,N_18793,N_18981);
xor U19041 (N_19041,N_18938,N_18798);
or U19042 (N_19042,N_18786,N_18816);
xnor U19043 (N_19043,N_18911,N_18760);
or U19044 (N_19044,N_18859,N_18809);
nor U19045 (N_19045,N_18942,N_18886);
xnor U19046 (N_19046,N_18954,N_18849);
and U19047 (N_19047,N_18874,N_18875);
and U19048 (N_19048,N_18823,N_18864);
or U19049 (N_19049,N_18908,N_18972);
or U19050 (N_19050,N_18975,N_18926);
and U19051 (N_19051,N_18763,N_18936);
and U19052 (N_19052,N_18844,N_18889);
nor U19053 (N_19053,N_18769,N_18836);
nor U19054 (N_19054,N_18768,N_18834);
nor U19055 (N_19055,N_18887,N_18820);
nand U19056 (N_19056,N_18939,N_18845);
nand U19057 (N_19057,N_18803,N_18752);
xnor U19058 (N_19058,N_18949,N_18865);
xnor U19059 (N_19059,N_18807,N_18986);
nand U19060 (N_19060,N_18904,N_18854);
or U19061 (N_19061,N_18789,N_18775);
or U19062 (N_19062,N_18971,N_18945);
nand U19063 (N_19063,N_18877,N_18919);
nor U19064 (N_19064,N_18883,N_18858);
nor U19065 (N_19065,N_18921,N_18982);
and U19066 (N_19066,N_18782,N_18817);
nand U19067 (N_19067,N_18856,N_18861);
or U19068 (N_19068,N_18898,N_18978);
and U19069 (N_19069,N_18873,N_18814);
or U19070 (N_19070,N_18754,N_18857);
and U19071 (N_19071,N_18828,N_18935);
and U19072 (N_19072,N_18891,N_18766);
xnor U19073 (N_19073,N_18762,N_18933);
nor U19074 (N_19074,N_18910,N_18987);
nor U19075 (N_19075,N_18890,N_18902);
or U19076 (N_19076,N_18984,N_18830);
nor U19077 (N_19077,N_18934,N_18994);
nor U19078 (N_19078,N_18767,N_18824);
xor U19079 (N_19079,N_18923,N_18862);
or U19080 (N_19080,N_18810,N_18784);
nor U19081 (N_19081,N_18912,N_18885);
xnor U19082 (N_19082,N_18870,N_18896);
nor U19083 (N_19083,N_18876,N_18801);
and U19084 (N_19084,N_18779,N_18947);
or U19085 (N_19085,N_18821,N_18925);
and U19086 (N_19086,N_18841,N_18882);
or U19087 (N_19087,N_18871,N_18974);
and U19088 (N_19088,N_18785,N_18931);
xor U19089 (N_19089,N_18811,N_18825);
or U19090 (N_19090,N_18928,N_18900);
or U19091 (N_19091,N_18985,N_18819);
and U19092 (N_19092,N_18780,N_18960);
nor U19093 (N_19093,N_18922,N_18750);
nand U19094 (N_19094,N_18869,N_18764);
nor U19095 (N_19095,N_18989,N_18957);
nand U19096 (N_19096,N_18927,N_18773);
or U19097 (N_19097,N_18860,N_18867);
xnor U19098 (N_19098,N_18757,N_18916);
nand U19099 (N_19099,N_18795,N_18878);
nand U19100 (N_19100,N_18992,N_18956);
nor U19101 (N_19101,N_18756,N_18812);
nand U19102 (N_19102,N_18977,N_18838);
nor U19103 (N_19103,N_18965,N_18917);
nand U19104 (N_19104,N_18997,N_18833);
nor U19105 (N_19105,N_18932,N_18777);
nand U19106 (N_19106,N_18813,N_18913);
nand U19107 (N_19107,N_18808,N_18802);
nor U19108 (N_19108,N_18805,N_18772);
nand U19109 (N_19109,N_18929,N_18791);
or U19110 (N_19110,N_18973,N_18897);
and U19111 (N_19111,N_18894,N_18829);
nand U19112 (N_19112,N_18995,N_18835);
and U19113 (N_19113,N_18799,N_18920);
or U19114 (N_19114,N_18948,N_18961);
or U19115 (N_19115,N_18943,N_18991);
nand U19116 (N_19116,N_18941,N_18818);
nand U19117 (N_19117,N_18893,N_18953);
or U19118 (N_19118,N_18980,N_18758);
or U19119 (N_19119,N_18850,N_18794);
nand U19120 (N_19120,N_18918,N_18837);
and U19121 (N_19121,N_18983,N_18930);
or U19122 (N_19122,N_18903,N_18832);
nor U19123 (N_19123,N_18790,N_18944);
nand U19124 (N_19124,N_18765,N_18915);
nor U19125 (N_19125,N_18756,N_18885);
and U19126 (N_19126,N_18822,N_18846);
and U19127 (N_19127,N_18913,N_18858);
nand U19128 (N_19128,N_18798,N_18859);
or U19129 (N_19129,N_18963,N_18791);
nor U19130 (N_19130,N_18752,N_18986);
xnor U19131 (N_19131,N_18785,N_18779);
nor U19132 (N_19132,N_18948,N_18814);
nand U19133 (N_19133,N_18943,N_18901);
and U19134 (N_19134,N_18952,N_18966);
xor U19135 (N_19135,N_18765,N_18966);
or U19136 (N_19136,N_18991,N_18915);
nor U19137 (N_19137,N_18889,N_18983);
nor U19138 (N_19138,N_18840,N_18994);
nor U19139 (N_19139,N_18769,N_18917);
nor U19140 (N_19140,N_18874,N_18767);
or U19141 (N_19141,N_18872,N_18925);
and U19142 (N_19142,N_18832,N_18856);
or U19143 (N_19143,N_18783,N_18852);
xor U19144 (N_19144,N_18790,N_18832);
xnor U19145 (N_19145,N_18879,N_18908);
nor U19146 (N_19146,N_18924,N_18879);
nand U19147 (N_19147,N_18786,N_18873);
or U19148 (N_19148,N_18915,N_18910);
xor U19149 (N_19149,N_18781,N_18802);
or U19150 (N_19150,N_18810,N_18867);
or U19151 (N_19151,N_18928,N_18884);
nand U19152 (N_19152,N_18953,N_18823);
xor U19153 (N_19153,N_18805,N_18925);
nand U19154 (N_19154,N_18990,N_18963);
or U19155 (N_19155,N_18768,N_18976);
or U19156 (N_19156,N_18809,N_18944);
or U19157 (N_19157,N_18791,N_18887);
and U19158 (N_19158,N_18766,N_18941);
and U19159 (N_19159,N_18754,N_18985);
xor U19160 (N_19160,N_18865,N_18755);
nor U19161 (N_19161,N_18863,N_18881);
nor U19162 (N_19162,N_18819,N_18763);
and U19163 (N_19163,N_18890,N_18820);
or U19164 (N_19164,N_18920,N_18892);
nand U19165 (N_19165,N_18820,N_18787);
nand U19166 (N_19166,N_18998,N_18972);
nor U19167 (N_19167,N_18869,N_18981);
nor U19168 (N_19168,N_18761,N_18807);
nand U19169 (N_19169,N_18778,N_18853);
nand U19170 (N_19170,N_18789,N_18848);
xnor U19171 (N_19171,N_18996,N_18885);
and U19172 (N_19172,N_18937,N_18842);
nor U19173 (N_19173,N_18997,N_18844);
and U19174 (N_19174,N_18821,N_18874);
nor U19175 (N_19175,N_18925,N_18803);
xor U19176 (N_19176,N_18845,N_18887);
or U19177 (N_19177,N_18981,N_18848);
nor U19178 (N_19178,N_18879,N_18946);
and U19179 (N_19179,N_18935,N_18847);
nor U19180 (N_19180,N_18941,N_18792);
nand U19181 (N_19181,N_18973,N_18756);
or U19182 (N_19182,N_18789,N_18891);
nor U19183 (N_19183,N_18845,N_18753);
nand U19184 (N_19184,N_18919,N_18850);
nand U19185 (N_19185,N_18814,N_18970);
and U19186 (N_19186,N_18796,N_18880);
and U19187 (N_19187,N_18961,N_18854);
nor U19188 (N_19188,N_18856,N_18843);
or U19189 (N_19189,N_18818,N_18787);
nor U19190 (N_19190,N_18935,N_18911);
or U19191 (N_19191,N_18940,N_18828);
or U19192 (N_19192,N_18987,N_18892);
xnor U19193 (N_19193,N_18819,N_18845);
nor U19194 (N_19194,N_18925,N_18957);
nand U19195 (N_19195,N_18996,N_18757);
xnor U19196 (N_19196,N_18947,N_18848);
nor U19197 (N_19197,N_18925,N_18780);
nor U19198 (N_19198,N_18805,N_18808);
or U19199 (N_19199,N_18841,N_18834);
nand U19200 (N_19200,N_18769,N_18826);
or U19201 (N_19201,N_18881,N_18759);
nor U19202 (N_19202,N_18893,N_18990);
nand U19203 (N_19203,N_18764,N_18959);
xor U19204 (N_19204,N_18835,N_18972);
or U19205 (N_19205,N_18955,N_18972);
xnor U19206 (N_19206,N_18953,N_18807);
nand U19207 (N_19207,N_18952,N_18931);
and U19208 (N_19208,N_18985,N_18841);
or U19209 (N_19209,N_18969,N_18995);
nand U19210 (N_19210,N_18957,N_18798);
nand U19211 (N_19211,N_18926,N_18857);
or U19212 (N_19212,N_18839,N_18759);
and U19213 (N_19213,N_18929,N_18796);
or U19214 (N_19214,N_18883,N_18875);
xnor U19215 (N_19215,N_18904,N_18901);
nand U19216 (N_19216,N_18842,N_18794);
or U19217 (N_19217,N_18991,N_18989);
nor U19218 (N_19218,N_18960,N_18947);
or U19219 (N_19219,N_18943,N_18903);
and U19220 (N_19220,N_18914,N_18783);
nor U19221 (N_19221,N_18996,N_18859);
and U19222 (N_19222,N_18829,N_18986);
and U19223 (N_19223,N_18785,N_18821);
or U19224 (N_19224,N_18964,N_18983);
and U19225 (N_19225,N_18994,N_18773);
or U19226 (N_19226,N_18873,N_18959);
and U19227 (N_19227,N_18938,N_18779);
nor U19228 (N_19228,N_18915,N_18899);
or U19229 (N_19229,N_18961,N_18951);
nor U19230 (N_19230,N_18816,N_18878);
nor U19231 (N_19231,N_18865,N_18798);
and U19232 (N_19232,N_18873,N_18965);
or U19233 (N_19233,N_18864,N_18983);
nor U19234 (N_19234,N_18786,N_18853);
and U19235 (N_19235,N_18793,N_18894);
and U19236 (N_19236,N_18767,N_18845);
and U19237 (N_19237,N_18818,N_18813);
and U19238 (N_19238,N_18755,N_18754);
nand U19239 (N_19239,N_18852,N_18871);
nand U19240 (N_19240,N_18980,N_18957);
nor U19241 (N_19241,N_18933,N_18915);
or U19242 (N_19242,N_18800,N_18828);
nor U19243 (N_19243,N_18875,N_18959);
or U19244 (N_19244,N_18766,N_18860);
nand U19245 (N_19245,N_18948,N_18906);
or U19246 (N_19246,N_18910,N_18828);
xnor U19247 (N_19247,N_18896,N_18917);
and U19248 (N_19248,N_18950,N_18998);
and U19249 (N_19249,N_18779,N_18814);
xor U19250 (N_19250,N_19059,N_19179);
and U19251 (N_19251,N_19084,N_19184);
and U19252 (N_19252,N_19122,N_19237);
nand U19253 (N_19253,N_19029,N_19174);
and U19254 (N_19254,N_19111,N_19074);
or U19255 (N_19255,N_19039,N_19138);
or U19256 (N_19256,N_19054,N_19093);
nand U19257 (N_19257,N_19119,N_19090);
and U19258 (N_19258,N_19200,N_19225);
or U19259 (N_19259,N_19035,N_19183);
nand U19260 (N_19260,N_19246,N_19025);
xnor U19261 (N_19261,N_19129,N_19095);
nor U19262 (N_19262,N_19005,N_19133);
and U19263 (N_19263,N_19128,N_19102);
nor U19264 (N_19264,N_19069,N_19242);
nor U19265 (N_19265,N_19023,N_19240);
nand U19266 (N_19266,N_19165,N_19064);
and U19267 (N_19267,N_19034,N_19002);
or U19268 (N_19268,N_19062,N_19190);
and U19269 (N_19269,N_19003,N_19234);
nand U19270 (N_19270,N_19121,N_19016);
or U19271 (N_19271,N_19141,N_19143);
or U19272 (N_19272,N_19108,N_19080);
or U19273 (N_19273,N_19157,N_19088);
nand U19274 (N_19274,N_19092,N_19186);
nor U19275 (N_19275,N_19065,N_19169);
and U19276 (N_19276,N_19154,N_19032);
or U19277 (N_19277,N_19203,N_19006);
xnor U19278 (N_19278,N_19118,N_19137);
and U19279 (N_19279,N_19012,N_19040);
nor U19280 (N_19280,N_19055,N_19087);
nor U19281 (N_19281,N_19124,N_19209);
nor U19282 (N_19282,N_19170,N_19221);
and U19283 (N_19283,N_19213,N_19191);
and U19284 (N_19284,N_19053,N_19175);
xor U19285 (N_19285,N_19049,N_19127);
or U19286 (N_19286,N_19142,N_19104);
or U19287 (N_19287,N_19113,N_19197);
nor U19288 (N_19288,N_19027,N_19238);
and U19289 (N_19289,N_19105,N_19130);
nor U19290 (N_19290,N_19222,N_19231);
and U19291 (N_19291,N_19145,N_19163);
nand U19292 (N_19292,N_19063,N_19009);
nand U19293 (N_19293,N_19230,N_19198);
nand U19294 (N_19294,N_19178,N_19004);
and U19295 (N_19295,N_19192,N_19233);
nand U19296 (N_19296,N_19245,N_19199);
xor U19297 (N_19297,N_19236,N_19140);
nor U19298 (N_19298,N_19126,N_19151);
nor U19299 (N_19299,N_19239,N_19132);
xnor U19300 (N_19300,N_19116,N_19217);
nor U19301 (N_19301,N_19048,N_19147);
or U19302 (N_19302,N_19103,N_19135);
nor U19303 (N_19303,N_19187,N_19071);
and U19304 (N_19304,N_19086,N_19070);
or U19305 (N_19305,N_19038,N_19114);
or U19306 (N_19306,N_19153,N_19218);
and U19307 (N_19307,N_19101,N_19219);
nand U19308 (N_19308,N_19037,N_19017);
and U19309 (N_19309,N_19073,N_19216);
and U19310 (N_19310,N_19232,N_19161);
nand U19311 (N_19311,N_19195,N_19176);
and U19312 (N_19312,N_19051,N_19189);
xnor U19313 (N_19313,N_19028,N_19208);
or U19314 (N_19314,N_19041,N_19000);
nor U19315 (N_19315,N_19204,N_19146);
nand U19316 (N_19316,N_19120,N_19223);
and U19317 (N_19317,N_19019,N_19010);
nand U19318 (N_19318,N_19097,N_19091);
nor U19319 (N_19319,N_19125,N_19043);
and U19320 (N_19320,N_19085,N_19008);
nor U19321 (N_19321,N_19220,N_19036);
nand U19322 (N_19322,N_19030,N_19158);
or U19323 (N_19323,N_19248,N_19079);
or U19324 (N_19324,N_19033,N_19112);
nand U19325 (N_19325,N_19226,N_19060);
nor U19326 (N_19326,N_19056,N_19107);
nor U19327 (N_19327,N_19235,N_19244);
and U19328 (N_19328,N_19021,N_19068);
nand U19329 (N_19329,N_19177,N_19078);
nand U19330 (N_19330,N_19099,N_19182);
nor U19331 (N_19331,N_19148,N_19052);
nand U19332 (N_19332,N_19045,N_19188);
and U19333 (N_19333,N_19098,N_19160);
nor U19334 (N_19334,N_19058,N_19083);
and U19335 (N_19335,N_19047,N_19013);
nand U19336 (N_19336,N_19022,N_19202);
nor U19337 (N_19337,N_19089,N_19150);
nand U19338 (N_19338,N_19007,N_19094);
and U19339 (N_19339,N_19057,N_19211);
xnor U19340 (N_19340,N_19046,N_19224);
xnor U19341 (N_19341,N_19156,N_19072);
and U19342 (N_19342,N_19172,N_19131);
or U19343 (N_19343,N_19144,N_19193);
nor U19344 (N_19344,N_19166,N_19066);
or U19345 (N_19345,N_19075,N_19044);
and U19346 (N_19346,N_19162,N_19115);
xnor U19347 (N_19347,N_19159,N_19139);
nor U19348 (N_19348,N_19228,N_19229);
or U19349 (N_19349,N_19206,N_19212);
nand U19350 (N_19350,N_19136,N_19210);
nor U19351 (N_19351,N_19185,N_19082);
and U19352 (N_19352,N_19020,N_19109);
or U19353 (N_19353,N_19001,N_19077);
and U19354 (N_19354,N_19123,N_19015);
nor U19355 (N_19355,N_19031,N_19081);
or U19356 (N_19356,N_19011,N_19205);
and U19357 (N_19357,N_19096,N_19173);
nand U19358 (N_19358,N_19180,N_19110);
and U19359 (N_19359,N_19241,N_19168);
or U19360 (N_19360,N_19042,N_19152);
or U19361 (N_19361,N_19024,N_19194);
nand U19362 (N_19362,N_19201,N_19171);
nor U19363 (N_19363,N_19247,N_19061);
and U19364 (N_19364,N_19134,N_19018);
or U19365 (N_19365,N_19249,N_19076);
and U19366 (N_19366,N_19243,N_19196);
xor U19367 (N_19367,N_19155,N_19227);
and U19368 (N_19368,N_19215,N_19167);
or U19369 (N_19369,N_19100,N_19181);
and U19370 (N_19370,N_19207,N_19117);
nor U19371 (N_19371,N_19050,N_19026);
and U19372 (N_19372,N_19106,N_19149);
or U19373 (N_19373,N_19067,N_19214);
nor U19374 (N_19374,N_19014,N_19164);
xor U19375 (N_19375,N_19177,N_19105);
nor U19376 (N_19376,N_19132,N_19241);
nor U19377 (N_19377,N_19212,N_19103);
nand U19378 (N_19378,N_19057,N_19131);
and U19379 (N_19379,N_19210,N_19000);
nor U19380 (N_19380,N_19112,N_19018);
nor U19381 (N_19381,N_19113,N_19198);
or U19382 (N_19382,N_19216,N_19222);
or U19383 (N_19383,N_19136,N_19220);
xnor U19384 (N_19384,N_19133,N_19051);
and U19385 (N_19385,N_19171,N_19200);
or U19386 (N_19386,N_19048,N_19198);
nand U19387 (N_19387,N_19223,N_19081);
and U19388 (N_19388,N_19178,N_19101);
or U19389 (N_19389,N_19120,N_19056);
nor U19390 (N_19390,N_19196,N_19092);
and U19391 (N_19391,N_19144,N_19248);
or U19392 (N_19392,N_19047,N_19200);
and U19393 (N_19393,N_19087,N_19152);
xor U19394 (N_19394,N_19031,N_19177);
nor U19395 (N_19395,N_19146,N_19084);
xor U19396 (N_19396,N_19118,N_19026);
nor U19397 (N_19397,N_19126,N_19142);
nand U19398 (N_19398,N_19066,N_19243);
and U19399 (N_19399,N_19073,N_19031);
and U19400 (N_19400,N_19186,N_19160);
and U19401 (N_19401,N_19133,N_19163);
nand U19402 (N_19402,N_19234,N_19164);
nor U19403 (N_19403,N_19089,N_19137);
nand U19404 (N_19404,N_19100,N_19200);
and U19405 (N_19405,N_19124,N_19007);
nand U19406 (N_19406,N_19167,N_19082);
and U19407 (N_19407,N_19053,N_19014);
nand U19408 (N_19408,N_19007,N_19075);
nand U19409 (N_19409,N_19103,N_19085);
nand U19410 (N_19410,N_19078,N_19231);
and U19411 (N_19411,N_19245,N_19229);
or U19412 (N_19412,N_19035,N_19244);
nand U19413 (N_19413,N_19079,N_19175);
and U19414 (N_19414,N_19001,N_19172);
and U19415 (N_19415,N_19202,N_19198);
and U19416 (N_19416,N_19002,N_19160);
and U19417 (N_19417,N_19063,N_19198);
nor U19418 (N_19418,N_19032,N_19207);
or U19419 (N_19419,N_19126,N_19080);
nor U19420 (N_19420,N_19089,N_19174);
or U19421 (N_19421,N_19186,N_19178);
nand U19422 (N_19422,N_19037,N_19182);
or U19423 (N_19423,N_19023,N_19160);
and U19424 (N_19424,N_19199,N_19166);
nor U19425 (N_19425,N_19195,N_19220);
xnor U19426 (N_19426,N_19105,N_19058);
and U19427 (N_19427,N_19027,N_19229);
nor U19428 (N_19428,N_19156,N_19146);
nand U19429 (N_19429,N_19071,N_19106);
nand U19430 (N_19430,N_19033,N_19052);
nor U19431 (N_19431,N_19223,N_19211);
nor U19432 (N_19432,N_19248,N_19204);
or U19433 (N_19433,N_19225,N_19149);
or U19434 (N_19434,N_19081,N_19051);
nand U19435 (N_19435,N_19022,N_19159);
nor U19436 (N_19436,N_19169,N_19135);
or U19437 (N_19437,N_19121,N_19221);
or U19438 (N_19438,N_19001,N_19220);
nand U19439 (N_19439,N_19132,N_19077);
and U19440 (N_19440,N_19216,N_19238);
nand U19441 (N_19441,N_19046,N_19118);
nand U19442 (N_19442,N_19073,N_19189);
nand U19443 (N_19443,N_19178,N_19059);
and U19444 (N_19444,N_19106,N_19042);
or U19445 (N_19445,N_19036,N_19239);
nor U19446 (N_19446,N_19056,N_19192);
xor U19447 (N_19447,N_19028,N_19140);
nor U19448 (N_19448,N_19080,N_19110);
or U19449 (N_19449,N_19093,N_19068);
nand U19450 (N_19450,N_19121,N_19165);
or U19451 (N_19451,N_19057,N_19147);
and U19452 (N_19452,N_19045,N_19092);
nor U19453 (N_19453,N_19093,N_19218);
nand U19454 (N_19454,N_19001,N_19175);
nand U19455 (N_19455,N_19093,N_19083);
and U19456 (N_19456,N_19171,N_19093);
nor U19457 (N_19457,N_19047,N_19127);
nor U19458 (N_19458,N_19078,N_19062);
and U19459 (N_19459,N_19172,N_19088);
nand U19460 (N_19460,N_19024,N_19076);
nor U19461 (N_19461,N_19157,N_19173);
xnor U19462 (N_19462,N_19063,N_19194);
xor U19463 (N_19463,N_19126,N_19072);
and U19464 (N_19464,N_19139,N_19241);
nand U19465 (N_19465,N_19187,N_19190);
nor U19466 (N_19466,N_19073,N_19027);
and U19467 (N_19467,N_19157,N_19136);
or U19468 (N_19468,N_19202,N_19228);
xor U19469 (N_19469,N_19018,N_19163);
xnor U19470 (N_19470,N_19180,N_19065);
or U19471 (N_19471,N_19206,N_19142);
nand U19472 (N_19472,N_19246,N_19105);
nand U19473 (N_19473,N_19037,N_19124);
xnor U19474 (N_19474,N_19166,N_19136);
or U19475 (N_19475,N_19003,N_19188);
nand U19476 (N_19476,N_19139,N_19095);
nand U19477 (N_19477,N_19132,N_19091);
nand U19478 (N_19478,N_19008,N_19235);
xor U19479 (N_19479,N_19199,N_19021);
and U19480 (N_19480,N_19191,N_19153);
and U19481 (N_19481,N_19053,N_19150);
and U19482 (N_19482,N_19149,N_19062);
and U19483 (N_19483,N_19069,N_19018);
nand U19484 (N_19484,N_19179,N_19151);
and U19485 (N_19485,N_19026,N_19017);
and U19486 (N_19486,N_19123,N_19120);
or U19487 (N_19487,N_19177,N_19168);
or U19488 (N_19488,N_19132,N_19111);
xnor U19489 (N_19489,N_19062,N_19072);
xnor U19490 (N_19490,N_19236,N_19086);
nand U19491 (N_19491,N_19132,N_19018);
nand U19492 (N_19492,N_19155,N_19238);
and U19493 (N_19493,N_19035,N_19193);
nand U19494 (N_19494,N_19160,N_19007);
and U19495 (N_19495,N_19021,N_19028);
or U19496 (N_19496,N_19198,N_19213);
or U19497 (N_19497,N_19139,N_19118);
or U19498 (N_19498,N_19027,N_19172);
nor U19499 (N_19499,N_19070,N_19080);
and U19500 (N_19500,N_19261,N_19424);
or U19501 (N_19501,N_19298,N_19254);
or U19502 (N_19502,N_19339,N_19275);
nand U19503 (N_19503,N_19406,N_19445);
xnor U19504 (N_19504,N_19310,N_19335);
nand U19505 (N_19505,N_19460,N_19475);
nand U19506 (N_19506,N_19472,N_19269);
nor U19507 (N_19507,N_19377,N_19267);
and U19508 (N_19508,N_19444,N_19262);
or U19509 (N_19509,N_19497,N_19312);
nor U19510 (N_19510,N_19354,N_19255);
nor U19511 (N_19511,N_19471,N_19495);
or U19512 (N_19512,N_19401,N_19399);
or U19513 (N_19513,N_19389,N_19301);
xor U19514 (N_19514,N_19321,N_19392);
xor U19515 (N_19515,N_19333,N_19348);
and U19516 (N_19516,N_19429,N_19409);
nor U19517 (N_19517,N_19430,N_19338);
nor U19518 (N_19518,N_19415,N_19371);
nor U19519 (N_19519,N_19258,N_19367);
and U19520 (N_19520,N_19324,N_19400);
or U19521 (N_19521,N_19363,N_19426);
or U19522 (N_19522,N_19441,N_19366);
nor U19523 (N_19523,N_19281,N_19420);
xor U19524 (N_19524,N_19264,N_19470);
and U19525 (N_19525,N_19271,N_19385);
nor U19526 (N_19526,N_19250,N_19266);
nor U19527 (N_19527,N_19467,N_19292);
and U19528 (N_19528,N_19357,N_19300);
nor U19529 (N_19529,N_19439,N_19370);
nor U19530 (N_19530,N_19422,N_19345);
or U19531 (N_19531,N_19440,N_19365);
and U19532 (N_19532,N_19252,N_19364);
nand U19533 (N_19533,N_19316,N_19383);
nand U19534 (N_19534,N_19373,N_19465);
or U19535 (N_19535,N_19270,N_19427);
nor U19536 (N_19536,N_19448,N_19265);
nor U19537 (N_19537,N_19280,N_19489);
nor U19538 (N_19538,N_19342,N_19311);
and U19539 (N_19539,N_19478,N_19408);
and U19540 (N_19540,N_19278,N_19332);
nand U19541 (N_19541,N_19337,N_19463);
and U19542 (N_19542,N_19378,N_19484);
nand U19543 (N_19543,N_19344,N_19251);
and U19544 (N_19544,N_19263,N_19381);
nor U19545 (N_19545,N_19346,N_19313);
or U19546 (N_19546,N_19368,N_19453);
nor U19547 (N_19547,N_19375,N_19395);
or U19548 (N_19548,N_19286,N_19274);
or U19549 (N_19549,N_19493,N_19474);
nor U19550 (N_19550,N_19343,N_19412);
or U19551 (N_19551,N_19355,N_19257);
nand U19552 (N_19552,N_19358,N_19442);
nand U19553 (N_19553,N_19486,N_19290);
or U19554 (N_19554,N_19432,N_19396);
nand U19555 (N_19555,N_19287,N_19329);
nor U19556 (N_19556,N_19410,N_19293);
and U19557 (N_19557,N_19386,N_19302);
nand U19558 (N_19558,N_19289,N_19323);
and U19559 (N_19559,N_19256,N_19380);
nor U19560 (N_19560,N_19319,N_19379);
nor U19561 (N_19561,N_19417,N_19499);
nand U19562 (N_19562,N_19359,N_19416);
and U19563 (N_19563,N_19374,N_19288);
or U19564 (N_19564,N_19382,N_19282);
xnor U19565 (N_19565,N_19330,N_19443);
xnor U19566 (N_19566,N_19414,N_19259);
nand U19567 (N_19567,N_19455,N_19483);
or U19568 (N_19568,N_19434,N_19352);
nand U19569 (N_19569,N_19418,N_19279);
and U19570 (N_19570,N_19277,N_19404);
and U19571 (N_19571,N_19309,N_19435);
or U19572 (N_19572,N_19260,N_19423);
or U19573 (N_19573,N_19303,N_19268);
or U19574 (N_19574,N_19306,N_19491);
xor U19575 (N_19575,N_19433,N_19446);
nor U19576 (N_19576,N_19314,N_19360);
or U19577 (N_19577,N_19391,N_19459);
or U19578 (N_19578,N_19384,N_19327);
and U19579 (N_19579,N_19253,N_19437);
and U19580 (N_19580,N_19295,N_19353);
or U19581 (N_19581,N_19450,N_19449);
or U19582 (N_19582,N_19403,N_19487);
nor U19583 (N_19583,N_19390,N_19494);
and U19584 (N_19584,N_19480,N_19369);
and U19585 (N_19585,N_19473,N_19468);
or U19586 (N_19586,N_19461,N_19376);
nor U19587 (N_19587,N_19347,N_19304);
nor U19588 (N_19588,N_19485,N_19421);
nor U19589 (N_19589,N_19297,N_19305);
nor U19590 (N_19590,N_19413,N_19356);
or U19591 (N_19591,N_19498,N_19388);
xor U19592 (N_19592,N_19393,N_19447);
or U19593 (N_19593,N_19462,N_19331);
or U19594 (N_19594,N_19431,N_19496);
and U19595 (N_19595,N_19362,N_19372);
nand U19596 (N_19596,N_19349,N_19488);
nand U19597 (N_19597,N_19325,N_19456);
nor U19598 (N_19598,N_19272,N_19328);
nand U19599 (N_19599,N_19308,N_19464);
or U19600 (N_19600,N_19284,N_19340);
nor U19601 (N_19601,N_19457,N_19438);
nor U19602 (N_19602,N_19482,N_19322);
nand U19603 (N_19603,N_19466,N_19458);
nand U19604 (N_19604,N_19411,N_19405);
nand U19605 (N_19605,N_19387,N_19336);
or U19606 (N_19606,N_19476,N_19285);
or U19607 (N_19607,N_19398,N_19318);
or U19608 (N_19608,N_19407,N_19452);
or U19609 (N_19609,N_19397,N_19436);
nor U19610 (N_19610,N_19394,N_19315);
xnor U19611 (N_19611,N_19273,N_19320);
nand U19612 (N_19612,N_19454,N_19341);
nand U19613 (N_19613,N_19481,N_19317);
and U19614 (N_19614,N_19326,N_19490);
or U19615 (N_19615,N_19477,N_19294);
nand U19616 (N_19616,N_19350,N_19351);
and U19617 (N_19617,N_19361,N_19299);
or U19618 (N_19618,N_19428,N_19334);
nor U19619 (N_19619,N_19276,N_19479);
xor U19620 (N_19620,N_19492,N_19296);
nand U19621 (N_19621,N_19425,N_19307);
nand U19622 (N_19622,N_19451,N_19419);
or U19623 (N_19623,N_19291,N_19283);
and U19624 (N_19624,N_19469,N_19402);
or U19625 (N_19625,N_19301,N_19443);
and U19626 (N_19626,N_19371,N_19331);
xor U19627 (N_19627,N_19271,N_19430);
nand U19628 (N_19628,N_19389,N_19443);
or U19629 (N_19629,N_19444,N_19438);
or U19630 (N_19630,N_19316,N_19425);
nand U19631 (N_19631,N_19452,N_19314);
and U19632 (N_19632,N_19456,N_19404);
or U19633 (N_19633,N_19486,N_19269);
and U19634 (N_19634,N_19425,N_19381);
nand U19635 (N_19635,N_19290,N_19429);
xnor U19636 (N_19636,N_19278,N_19313);
and U19637 (N_19637,N_19429,N_19332);
nand U19638 (N_19638,N_19319,N_19448);
nand U19639 (N_19639,N_19423,N_19351);
or U19640 (N_19640,N_19417,N_19387);
nor U19641 (N_19641,N_19300,N_19331);
xor U19642 (N_19642,N_19332,N_19474);
nor U19643 (N_19643,N_19442,N_19259);
nand U19644 (N_19644,N_19408,N_19293);
or U19645 (N_19645,N_19295,N_19371);
nand U19646 (N_19646,N_19418,N_19436);
and U19647 (N_19647,N_19277,N_19310);
nor U19648 (N_19648,N_19433,N_19428);
nor U19649 (N_19649,N_19252,N_19299);
nor U19650 (N_19650,N_19402,N_19261);
nor U19651 (N_19651,N_19373,N_19371);
nor U19652 (N_19652,N_19493,N_19308);
nand U19653 (N_19653,N_19406,N_19305);
or U19654 (N_19654,N_19283,N_19303);
nand U19655 (N_19655,N_19338,N_19280);
and U19656 (N_19656,N_19337,N_19397);
nor U19657 (N_19657,N_19340,N_19470);
xor U19658 (N_19658,N_19344,N_19331);
nand U19659 (N_19659,N_19362,N_19446);
or U19660 (N_19660,N_19438,N_19470);
nand U19661 (N_19661,N_19356,N_19254);
nor U19662 (N_19662,N_19482,N_19297);
or U19663 (N_19663,N_19462,N_19313);
nand U19664 (N_19664,N_19403,N_19483);
or U19665 (N_19665,N_19313,N_19445);
or U19666 (N_19666,N_19344,N_19418);
nor U19667 (N_19667,N_19271,N_19321);
or U19668 (N_19668,N_19398,N_19438);
nor U19669 (N_19669,N_19498,N_19382);
or U19670 (N_19670,N_19387,N_19285);
nand U19671 (N_19671,N_19456,N_19422);
or U19672 (N_19672,N_19309,N_19414);
or U19673 (N_19673,N_19357,N_19489);
or U19674 (N_19674,N_19392,N_19330);
and U19675 (N_19675,N_19275,N_19385);
or U19676 (N_19676,N_19382,N_19299);
and U19677 (N_19677,N_19351,N_19368);
or U19678 (N_19678,N_19358,N_19352);
and U19679 (N_19679,N_19404,N_19442);
and U19680 (N_19680,N_19373,N_19497);
nor U19681 (N_19681,N_19463,N_19423);
and U19682 (N_19682,N_19406,N_19472);
nand U19683 (N_19683,N_19393,N_19268);
and U19684 (N_19684,N_19291,N_19389);
nand U19685 (N_19685,N_19388,N_19306);
and U19686 (N_19686,N_19354,N_19457);
nand U19687 (N_19687,N_19486,N_19496);
or U19688 (N_19688,N_19352,N_19443);
and U19689 (N_19689,N_19462,N_19422);
xor U19690 (N_19690,N_19284,N_19341);
nor U19691 (N_19691,N_19442,N_19377);
and U19692 (N_19692,N_19397,N_19456);
nor U19693 (N_19693,N_19457,N_19371);
nor U19694 (N_19694,N_19439,N_19414);
or U19695 (N_19695,N_19405,N_19441);
nand U19696 (N_19696,N_19324,N_19424);
nand U19697 (N_19697,N_19369,N_19463);
xor U19698 (N_19698,N_19350,N_19420);
nand U19699 (N_19699,N_19356,N_19380);
nand U19700 (N_19700,N_19416,N_19474);
or U19701 (N_19701,N_19336,N_19266);
nand U19702 (N_19702,N_19453,N_19277);
and U19703 (N_19703,N_19488,N_19401);
nor U19704 (N_19704,N_19495,N_19425);
nor U19705 (N_19705,N_19274,N_19425);
nor U19706 (N_19706,N_19437,N_19395);
xor U19707 (N_19707,N_19490,N_19298);
nand U19708 (N_19708,N_19281,N_19427);
nand U19709 (N_19709,N_19461,N_19285);
nor U19710 (N_19710,N_19461,N_19297);
and U19711 (N_19711,N_19271,N_19488);
nor U19712 (N_19712,N_19281,N_19383);
nor U19713 (N_19713,N_19431,N_19479);
nand U19714 (N_19714,N_19306,N_19351);
or U19715 (N_19715,N_19366,N_19294);
or U19716 (N_19716,N_19256,N_19299);
or U19717 (N_19717,N_19485,N_19284);
nand U19718 (N_19718,N_19484,N_19493);
and U19719 (N_19719,N_19400,N_19368);
and U19720 (N_19720,N_19314,N_19260);
and U19721 (N_19721,N_19319,N_19418);
and U19722 (N_19722,N_19340,N_19423);
and U19723 (N_19723,N_19339,N_19382);
xnor U19724 (N_19724,N_19383,N_19389);
or U19725 (N_19725,N_19282,N_19392);
xor U19726 (N_19726,N_19260,N_19252);
nor U19727 (N_19727,N_19481,N_19492);
and U19728 (N_19728,N_19428,N_19496);
or U19729 (N_19729,N_19374,N_19451);
or U19730 (N_19730,N_19250,N_19325);
nand U19731 (N_19731,N_19432,N_19497);
or U19732 (N_19732,N_19378,N_19487);
or U19733 (N_19733,N_19279,N_19432);
or U19734 (N_19734,N_19463,N_19327);
or U19735 (N_19735,N_19362,N_19436);
or U19736 (N_19736,N_19397,N_19309);
or U19737 (N_19737,N_19376,N_19418);
or U19738 (N_19738,N_19378,N_19269);
and U19739 (N_19739,N_19306,N_19369);
nand U19740 (N_19740,N_19319,N_19467);
or U19741 (N_19741,N_19343,N_19304);
or U19742 (N_19742,N_19468,N_19440);
and U19743 (N_19743,N_19457,N_19315);
nand U19744 (N_19744,N_19311,N_19276);
and U19745 (N_19745,N_19412,N_19250);
or U19746 (N_19746,N_19309,N_19359);
and U19747 (N_19747,N_19328,N_19478);
nor U19748 (N_19748,N_19323,N_19494);
and U19749 (N_19749,N_19395,N_19388);
nor U19750 (N_19750,N_19566,N_19520);
nand U19751 (N_19751,N_19734,N_19556);
nand U19752 (N_19752,N_19705,N_19604);
and U19753 (N_19753,N_19699,N_19632);
xor U19754 (N_19754,N_19693,N_19550);
xnor U19755 (N_19755,N_19679,N_19542);
and U19756 (N_19756,N_19683,N_19514);
nor U19757 (N_19757,N_19560,N_19587);
or U19758 (N_19758,N_19685,N_19538);
and U19759 (N_19759,N_19638,N_19649);
nand U19760 (N_19760,N_19633,N_19681);
xor U19761 (N_19761,N_19745,N_19674);
and U19762 (N_19762,N_19531,N_19618);
or U19763 (N_19763,N_19664,N_19748);
or U19764 (N_19764,N_19534,N_19720);
nand U19765 (N_19765,N_19673,N_19564);
nand U19766 (N_19766,N_19608,N_19606);
nand U19767 (N_19767,N_19594,N_19529);
nor U19768 (N_19768,N_19688,N_19667);
or U19769 (N_19769,N_19635,N_19581);
nand U19770 (N_19770,N_19503,N_19569);
and U19771 (N_19771,N_19710,N_19694);
nand U19772 (N_19772,N_19665,N_19675);
and U19773 (N_19773,N_19509,N_19640);
nor U19774 (N_19774,N_19714,N_19631);
and U19775 (N_19775,N_19661,N_19735);
nor U19776 (N_19776,N_19702,N_19582);
nor U19777 (N_19777,N_19506,N_19590);
or U19778 (N_19778,N_19572,N_19712);
nand U19779 (N_19779,N_19684,N_19639);
xor U19780 (N_19780,N_19553,N_19613);
and U19781 (N_19781,N_19519,N_19744);
nand U19782 (N_19782,N_19727,N_19525);
nand U19783 (N_19783,N_19657,N_19703);
nand U19784 (N_19784,N_19636,N_19687);
nand U19785 (N_19785,N_19588,N_19725);
or U19786 (N_19786,N_19648,N_19521);
nor U19787 (N_19787,N_19616,N_19709);
nor U19788 (N_19788,N_19686,N_19620);
and U19789 (N_19789,N_19698,N_19697);
nor U19790 (N_19790,N_19577,N_19585);
and U19791 (N_19791,N_19523,N_19637);
or U19792 (N_19792,N_19568,N_19549);
nand U19793 (N_19793,N_19733,N_19557);
and U19794 (N_19794,N_19539,N_19610);
nor U19795 (N_19795,N_19645,N_19626);
or U19796 (N_19796,N_19600,N_19641);
and U19797 (N_19797,N_19644,N_19736);
nor U19798 (N_19798,N_19695,N_19548);
and U19799 (N_19799,N_19551,N_19724);
xor U19800 (N_19800,N_19715,N_19743);
nor U19801 (N_19801,N_19722,N_19691);
or U19802 (N_19802,N_19669,N_19670);
nor U19803 (N_19803,N_19532,N_19562);
xnor U19804 (N_19804,N_19502,N_19629);
or U19805 (N_19805,N_19563,N_19627);
and U19806 (N_19806,N_19574,N_19742);
nor U19807 (N_19807,N_19711,N_19614);
nand U19808 (N_19808,N_19729,N_19630);
or U19809 (N_19809,N_19654,N_19653);
nand U19810 (N_19810,N_19628,N_19612);
nor U19811 (N_19811,N_19545,N_19652);
or U19812 (N_19812,N_19676,N_19726);
and U19813 (N_19813,N_19597,N_19561);
nand U19814 (N_19814,N_19501,N_19619);
or U19815 (N_19815,N_19515,N_19718);
nand U19816 (N_19816,N_19730,N_19536);
and U19817 (N_19817,N_19728,N_19598);
xor U19818 (N_19818,N_19552,N_19659);
and U19819 (N_19819,N_19500,N_19625);
or U19820 (N_19820,N_19599,N_19747);
nor U19821 (N_19821,N_19739,N_19646);
xnor U19822 (N_19822,N_19655,N_19690);
and U19823 (N_19823,N_19555,N_19576);
nor U19824 (N_19824,N_19544,N_19541);
or U19825 (N_19825,N_19680,N_19660);
nand U19826 (N_19826,N_19731,N_19701);
nor U19827 (N_19827,N_19708,N_19516);
xnor U19828 (N_19828,N_19622,N_19706);
xor U19829 (N_19829,N_19603,N_19647);
nand U19830 (N_19830,N_19666,N_19584);
nor U19831 (N_19831,N_19696,N_19672);
or U19832 (N_19832,N_19634,N_19578);
or U19833 (N_19833,N_19740,N_19573);
and U19834 (N_19834,N_19716,N_19554);
nand U19835 (N_19835,N_19513,N_19583);
nor U19836 (N_19836,N_19677,N_19526);
and U19837 (N_19837,N_19596,N_19591);
or U19838 (N_19838,N_19546,N_19707);
xnor U19839 (N_19839,N_19540,N_19528);
nor U19840 (N_19840,N_19537,N_19579);
or U19841 (N_19841,N_19678,N_19558);
nand U19842 (N_19842,N_19723,N_19504);
nor U19843 (N_19843,N_19671,N_19530);
nand U19844 (N_19844,N_19533,N_19607);
xor U19845 (N_19845,N_19592,N_19656);
nand U19846 (N_19846,N_19524,N_19611);
nor U19847 (N_19847,N_19589,N_19580);
nor U19848 (N_19848,N_19567,N_19700);
nand U19849 (N_19849,N_19713,N_19651);
nand U19850 (N_19850,N_19737,N_19593);
and U19851 (N_19851,N_19623,N_19559);
nand U19852 (N_19852,N_19575,N_19662);
or U19853 (N_19853,N_19642,N_19602);
and U19854 (N_19854,N_19522,N_19650);
xnor U19855 (N_19855,N_19738,N_19527);
nand U19856 (N_19856,N_19511,N_19689);
and U19857 (N_19857,N_19609,N_19658);
nand U19858 (N_19858,N_19605,N_19565);
nor U19859 (N_19859,N_19547,N_19663);
and U19860 (N_19860,N_19746,N_19518);
or U19861 (N_19861,N_19749,N_19543);
or U19862 (N_19862,N_19624,N_19732);
and U19863 (N_19863,N_19741,N_19668);
and U19864 (N_19864,N_19682,N_19621);
or U19865 (N_19865,N_19601,N_19721);
nand U19866 (N_19866,N_19507,N_19505);
and U19867 (N_19867,N_19719,N_19571);
nor U19868 (N_19868,N_19617,N_19704);
and U19869 (N_19869,N_19517,N_19595);
or U19870 (N_19870,N_19643,N_19717);
and U19871 (N_19871,N_19586,N_19615);
and U19872 (N_19872,N_19510,N_19692);
nand U19873 (N_19873,N_19570,N_19535);
nand U19874 (N_19874,N_19508,N_19512);
nand U19875 (N_19875,N_19523,N_19616);
and U19876 (N_19876,N_19590,N_19718);
and U19877 (N_19877,N_19706,N_19524);
nand U19878 (N_19878,N_19534,N_19518);
xnor U19879 (N_19879,N_19690,N_19680);
or U19880 (N_19880,N_19710,N_19678);
or U19881 (N_19881,N_19639,N_19536);
or U19882 (N_19882,N_19697,N_19748);
xnor U19883 (N_19883,N_19666,N_19700);
xor U19884 (N_19884,N_19644,N_19512);
or U19885 (N_19885,N_19718,N_19707);
nand U19886 (N_19886,N_19601,N_19662);
and U19887 (N_19887,N_19680,N_19747);
and U19888 (N_19888,N_19522,N_19595);
nand U19889 (N_19889,N_19591,N_19743);
xor U19890 (N_19890,N_19650,N_19648);
nand U19891 (N_19891,N_19744,N_19575);
nor U19892 (N_19892,N_19629,N_19518);
or U19893 (N_19893,N_19649,N_19539);
xnor U19894 (N_19894,N_19555,N_19613);
xnor U19895 (N_19895,N_19710,N_19748);
and U19896 (N_19896,N_19749,N_19642);
and U19897 (N_19897,N_19508,N_19746);
nor U19898 (N_19898,N_19610,N_19737);
xor U19899 (N_19899,N_19559,N_19735);
xnor U19900 (N_19900,N_19658,N_19639);
nor U19901 (N_19901,N_19619,N_19642);
nand U19902 (N_19902,N_19719,N_19556);
nor U19903 (N_19903,N_19583,N_19613);
or U19904 (N_19904,N_19560,N_19605);
nor U19905 (N_19905,N_19709,N_19683);
nand U19906 (N_19906,N_19537,N_19534);
and U19907 (N_19907,N_19615,N_19713);
and U19908 (N_19908,N_19516,N_19554);
nand U19909 (N_19909,N_19693,N_19747);
nand U19910 (N_19910,N_19508,N_19619);
nand U19911 (N_19911,N_19643,N_19553);
nor U19912 (N_19912,N_19692,N_19542);
nor U19913 (N_19913,N_19576,N_19650);
nor U19914 (N_19914,N_19716,N_19563);
xnor U19915 (N_19915,N_19563,N_19727);
and U19916 (N_19916,N_19679,N_19680);
or U19917 (N_19917,N_19721,N_19591);
or U19918 (N_19918,N_19649,N_19603);
or U19919 (N_19919,N_19655,N_19539);
nand U19920 (N_19920,N_19537,N_19726);
or U19921 (N_19921,N_19741,N_19729);
or U19922 (N_19922,N_19729,N_19602);
and U19923 (N_19923,N_19748,N_19723);
or U19924 (N_19924,N_19578,N_19702);
xnor U19925 (N_19925,N_19569,N_19737);
and U19926 (N_19926,N_19694,N_19659);
and U19927 (N_19927,N_19668,N_19524);
or U19928 (N_19928,N_19610,N_19501);
or U19929 (N_19929,N_19722,N_19675);
and U19930 (N_19930,N_19631,N_19727);
nor U19931 (N_19931,N_19698,N_19582);
or U19932 (N_19932,N_19675,N_19689);
and U19933 (N_19933,N_19554,N_19531);
nor U19934 (N_19934,N_19664,N_19699);
nor U19935 (N_19935,N_19581,N_19740);
nor U19936 (N_19936,N_19542,N_19522);
or U19937 (N_19937,N_19637,N_19500);
or U19938 (N_19938,N_19602,N_19542);
or U19939 (N_19939,N_19605,N_19640);
and U19940 (N_19940,N_19730,N_19562);
nand U19941 (N_19941,N_19570,N_19730);
or U19942 (N_19942,N_19560,N_19707);
nor U19943 (N_19943,N_19709,N_19575);
and U19944 (N_19944,N_19730,N_19539);
or U19945 (N_19945,N_19543,N_19567);
and U19946 (N_19946,N_19558,N_19741);
or U19947 (N_19947,N_19698,N_19549);
or U19948 (N_19948,N_19608,N_19604);
xor U19949 (N_19949,N_19722,N_19670);
nand U19950 (N_19950,N_19551,N_19533);
xor U19951 (N_19951,N_19601,N_19501);
nand U19952 (N_19952,N_19620,N_19524);
or U19953 (N_19953,N_19502,N_19690);
nand U19954 (N_19954,N_19667,N_19631);
xor U19955 (N_19955,N_19504,N_19592);
or U19956 (N_19956,N_19567,N_19654);
or U19957 (N_19957,N_19623,N_19722);
and U19958 (N_19958,N_19582,N_19660);
or U19959 (N_19959,N_19717,N_19664);
and U19960 (N_19960,N_19609,N_19663);
nand U19961 (N_19961,N_19653,N_19684);
and U19962 (N_19962,N_19522,N_19518);
or U19963 (N_19963,N_19741,N_19744);
xnor U19964 (N_19964,N_19542,N_19707);
or U19965 (N_19965,N_19662,N_19569);
and U19966 (N_19966,N_19544,N_19580);
or U19967 (N_19967,N_19526,N_19672);
and U19968 (N_19968,N_19554,N_19739);
nand U19969 (N_19969,N_19594,N_19553);
xor U19970 (N_19970,N_19566,N_19640);
and U19971 (N_19971,N_19606,N_19717);
and U19972 (N_19972,N_19734,N_19587);
and U19973 (N_19973,N_19526,N_19700);
or U19974 (N_19974,N_19625,N_19723);
and U19975 (N_19975,N_19573,N_19502);
xor U19976 (N_19976,N_19518,N_19610);
nor U19977 (N_19977,N_19528,N_19534);
and U19978 (N_19978,N_19591,N_19513);
nand U19979 (N_19979,N_19597,N_19571);
nand U19980 (N_19980,N_19673,N_19665);
nand U19981 (N_19981,N_19733,N_19700);
or U19982 (N_19982,N_19546,N_19660);
or U19983 (N_19983,N_19706,N_19637);
or U19984 (N_19984,N_19735,N_19660);
nor U19985 (N_19985,N_19724,N_19710);
and U19986 (N_19986,N_19731,N_19678);
and U19987 (N_19987,N_19515,N_19632);
or U19988 (N_19988,N_19601,N_19638);
nand U19989 (N_19989,N_19686,N_19580);
nor U19990 (N_19990,N_19552,N_19662);
nand U19991 (N_19991,N_19612,N_19623);
nand U19992 (N_19992,N_19730,N_19606);
and U19993 (N_19993,N_19516,N_19520);
nor U19994 (N_19994,N_19696,N_19562);
xnor U19995 (N_19995,N_19730,N_19599);
or U19996 (N_19996,N_19606,N_19535);
and U19997 (N_19997,N_19529,N_19704);
xnor U19998 (N_19998,N_19632,N_19593);
nand U19999 (N_19999,N_19565,N_19571);
and U20000 (N_20000,N_19929,N_19800);
and U20001 (N_20001,N_19906,N_19888);
nor U20002 (N_20002,N_19933,N_19856);
and U20003 (N_20003,N_19814,N_19945);
and U20004 (N_20004,N_19910,N_19980);
or U20005 (N_20005,N_19836,N_19838);
nand U20006 (N_20006,N_19843,N_19771);
or U20007 (N_20007,N_19818,N_19764);
or U20008 (N_20008,N_19950,N_19878);
or U20009 (N_20009,N_19908,N_19953);
and U20010 (N_20010,N_19979,N_19847);
and U20011 (N_20011,N_19808,N_19880);
or U20012 (N_20012,N_19909,N_19799);
nor U20013 (N_20013,N_19751,N_19896);
nor U20014 (N_20014,N_19840,N_19887);
nor U20015 (N_20015,N_19999,N_19823);
or U20016 (N_20016,N_19901,N_19826);
or U20017 (N_20017,N_19892,N_19768);
or U20018 (N_20018,N_19873,N_19855);
or U20019 (N_20019,N_19867,N_19796);
nand U20020 (N_20020,N_19996,N_19778);
nor U20021 (N_20021,N_19951,N_19824);
xor U20022 (N_20022,N_19852,N_19981);
or U20023 (N_20023,N_19988,N_19825);
or U20024 (N_20024,N_19829,N_19923);
nand U20025 (N_20025,N_19932,N_19756);
xnor U20026 (N_20026,N_19822,N_19970);
or U20027 (N_20027,N_19889,N_19767);
nand U20028 (N_20028,N_19957,N_19915);
xor U20029 (N_20029,N_19968,N_19962);
and U20030 (N_20030,N_19890,N_19786);
nor U20031 (N_20031,N_19986,N_19955);
or U20032 (N_20032,N_19788,N_19918);
xor U20033 (N_20033,N_19922,N_19914);
xnor U20034 (N_20034,N_19937,N_19921);
or U20035 (N_20035,N_19780,N_19924);
xor U20036 (N_20036,N_19973,N_19900);
and U20037 (N_20037,N_19985,N_19883);
or U20038 (N_20038,N_19812,N_19787);
or U20039 (N_20039,N_19763,N_19903);
xor U20040 (N_20040,N_19833,N_19783);
or U20041 (N_20041,N_19998,N_19835);
and U20042 (N_20042,N_19958,N_19765);
nor U20043 (N_20043,N_19804,N_19948);
xor U20044 (N_20044,N_19877,N_19895);
nand U20045 (N_20045,N_19960,N_19819);
and U20046 (N_20046,N_19795,N_19934);
or U20047 (N_20047,N_19874,N_19758);
nand U20048 (N_20048,N_19911,N_19966);
and U20049 (N_20049,N_19854,N_19961);
and U20050 (N_20050,N_19801,N_19991);
or U20051 (N_20051,N_19941,N_19884);
nor U20052 (N_20052,N_19817,N_19913);
or U20053 (N_20053,N_19912,N_19893);
nand U20054 (N_20054,N_19789,N_19875);
nand U20055 (N_20055,N_19757,N_19885);
nor U20056 (N_20056,N_19978,N_19997);
and U20057 (N_20057,N_19865,N_19868);
nand U20058 (N_20058,N_19956,N_19927);
nand U20059 (N_20059,N_19831,N_19853);
nand U20060 (N_20060,N_19790,N_19940);
and U20061 (N_20061,N_19839,N_19754);
and U20062 (N_20062,N_19907,N_19841);
xnor U20063 (N_20063,N_19827,N_19784);
and U20064 (N_20064,N_19936,N_19872);
nand U20065 (N_20065,N_19864,N_19845);
xor U20066 (N_20066,N_19811,N_19870);
and U20067 (N_20067,N_19776,N_19886);
nand U20068 (N_20068,N_19777,N_19965);
or U20069 (N_20069,N_19769,N_19994);
nor U20070 (N_20070,N_19871,N_19820);
nor U20071 (N_20071,N_19946,N_19898);
and U20072 (N_20072,N_19809,N_19815);
or U20073 (N_20073,N_19926,N_19976);
nor U20074 (N_20074,N_19916,N_19938);
nor U20075 (N_20075,N_19806,N_19935);
or U20076 (N_20076,N_19813,N_19925);
nor U20077 (N_20077,N_19990,N_19860);
xnor U20078 (N_20078,N_19761,N_19802);
and U20079 (N_20079,N_19995,N_19770);
and U20080 (N_20080,N_19897,N_19905);
or U20081 (N_20081,N_19832,N_19848);
or U20082 (N_20082,N_19899,N_19807);
and U20083 (N_20083,N_19882,N_19821);
xor U20084 (N_20084,N_19891,N_19775);
nor U20085 (N_20085,N_19837,N_19942);
nor U20086 (N_20086,N_19952,N_19857);
nand U20087 (N_20087,N_19944,N_19816);
and U20088 (N_20088,N_19851,N_19774);
and U20089 (N_20089,N_19850,N_19928);
or U20090 (N_20090,N_19773,N_19869);
xnor U20091 (N_20091,N_19989,N_19977);
or U20092 (N_20092,N_19861,N_19943);
nor U20093 (N_20093,N_19752,N_19959);
nor U20094 (N_20094,N_19766,N_19930);
nor U20095 (N_20095,N_19793,N_19931);
nor U20096 (N_20096,N_19830,N_19805);
or U20097 (N_20097,N_19785,N_19834);
and U20098 (N_20098,N_19920,N_19964);
nor U20099 (N_20099,N_19772,N_19760);
xor U20100 (N_20100,N_19987,N_19967);
and U20101 (N_20101,N_19803,N_19863);
nor U20102 (N_20102,N_19750,N_19879);
nand U20103 (N_20103,N_19939,N_19992);
and U20104 (N_20104,N_19794,N_19762);
nand U20105 (N_20105,N_19791,N_19902);
nor U20106 (N_20106,N_19917,N_19759);
nor U20107 (N_20107,N_19842,N_19963);
nor U20108 (N_20108,N_19858,N_19881);
nand U20109 (N_20109,N_19810,N_19982);
and U20110 (N_20110,N_19993,N_19797);
nand U20111 (N_20111,N_19866,N_19954);
or U20112 (N_20112,N_19782,N_19984);
xor U20113 (N_20113,N_19844,N_19969);
or U20114 (N_20114,N_19894,N_19971);
or U20115 (N_20115,N_19753,N_19876);
and U20116 (N_20116,N_19972,N_19846);
or U20117 (N_20117,N_19919,N_19779);
and U20118 (N_20118,N_19947,N_19781);
nor U20119 (N_20119,N_19975,N_19849);
nor U20120 (N_20120,N_19792,N_19983);
or U20121 (N_20121,N_19862,N_19755);
and U20122 (N_20122,N_19828,N_19798);
nor U20123 (N_20123,N_19974,N_19904);
or U20124 (N_20124,N_19859,N_19949);
nor U20125 (N_20125,N_19768,N_19873);
nand U20126 (N_20126,N_19871,N_19857);
or U20127 (N_20127,N_19753,N_19899);
nor U20128 (N_20128,N_19985,N_19806);
nand U20129 (N_20129,N_19826,N_19977);
nor U20130 (N_20130,N_19867,N_19775);
or U20131 (N_20131,N_19960,N_19805);
or U20132 (N_20132,N_19977,N_19908);
xnor U20133 (N_20133,N_19985,N_19823);
and U20134 (N_20134,N_19794,N_19793);
or U20135 (N_20135,N_19995,N_19877);
and U20136 (N_20136,N_19922,N_19980);
nand U20137 (N_20137,N_19774,N_19997);
nand U20138 (N_20138,N_19932,N_19906);
and U20139 (N_20139,N_19878,N_19956);
or U20140 (N_20140,N_19754,N_19991);
nand U20141 (N_20141,N_19964,N_19787);
nor U20142 (N_20142,N_19775,N_19918);
and U20143 (N_20143,N_19930,N_19966);
and U20144 (N_20144,N_19861,N_19894);
nand U20145 (N_20145,N_19877,N_19843);
nand U20146 (N_20146,N_19993,N_19933);
and U20147 (N_20147,N_19861,N_19868);
and U20148 (N_20148,N_19825,N_19859);
nor U20149 (N_20149,N_19762,N_19842);
nor U20150 (N_20150,N_19998,N_19887);
xor U20151 (N_20151,N_19808,N_19751);
nand U20152 (N_20152,N_19803,N_19784);
xor U20153 (N_20153,N_19754,N_19964);
or U20154 (N_20154,N_19760,N_19827);
nor U20155 (N_20155,N_19868,N_19992);
and U20156 (N_20156,N_19894,N_19964);
nor U20157 (N_20157,N_19788,N_19832);
nand U20158 (N_20158,N_19958,N_19955);
nor U20159 (N_20159,N_19762,N_19788);
or U20160 (N_20160,N_19914,N_19838);
and U20161 (N_20161,N_19776,N_19858);
nand U20162 (N_20162,N_19750,N_19897);
or U20163 (N_20163,N_19977,N_19877);
and U20164 (N_20164,N_19815,N_19853);
nand U20165 (N_20165,N_19912,N_19963);
or U20166 (N_20166,N_19951,N_19949);
and U20167 (N_20167,N_19759,N_19895);
or U20168 (N_20168,N_19882,N_19788);
xor U20169 (N_20169,N_19935,N_19786);
and U20170 (N_20170,N_19866,N_19791);
nor U20171 (N_20171,N_19915,N_19809);
and U20172 (N_20172,N_19785,N_19842);
and U20173 (N_20173,N_19855,N_19941);
and U20174 (N_20174,N_19921,N_19986);
nor U20175 (N_20175,N_19969,N_19908);
or U20176 (N_20176,N_19914,N_19995);
nand U20177 (N_20177,N_19989,N_19879);
and U20178 (N_20178,N_19906,N_19750);
or U20179 (N_20179,N_19972,N_19856);
nand U20180 (N_20180,N_19962,N_19821);
and U20181 (N_20181,N_19960,N_19962);
and U20182 (N_20182,N_19836,N_19821);
nor U20183 (N_20183,N_19986,N_19974);
nand U20184 (N_20184,N_19756,N_19776);
nand U20185 (N_20185,N_19970,N_19957);
nor U20186 (N_20186,N_19943,N_19892);
nor U20187 (N_20187,N_19758,N_19762);
and U20188 (N_20188,N_19829,N_19771);
and U20189 (N_20189,N_19757,N_19994);
nand U20190 (N_20190,N_19919,N_19837);
nand U20191 (N_20191,N_19833,N_19929);
and U20192 (N_20192,N_19807,N_19764);
nor U20193 (N_20193,N_19910,N_19952);
nor U20194 (N_20194,N_19774,N_19816);
or U20195 (N_20195,N_19932,N_19859);
or U20196 (N_20196,N_19991,N_19872);
or U20197 (N_20197,N_19959,N_19965);
nor U20198 (N_20198,N_19767,N_19894);
nor U20199 (N_20199,N_19802,N_19870);
and U20200 (N_20200,N_19769,N_19956);
nand U20201 (N_20201,N_19790,N_19975);
nor U20202 (N_20202,N_19755,N_19830);
and U20203 (N_20203,N_19915,N_19970);
or U20204 (N_20204,N_19884,N_19873);
or U20205 (N_20205,N_19836,N_19990);
xor U20206 (N_20206,N_19831,N_19936);
or U20207 (N_20207,N_19944,N_19797);
nor U20208 (N_20208,N_19872,N_19993);
xor U20209 (N_20209,N_19857,N_19861);
or U20210 (N_20210,N_19913,N_19789);
nor U20211 (N_20211,N_19904,N_19772);
xnor U20212 (N_20212,N_19851,N_19866);
and U20213 (N_20213,N_19916,N_19796);
and U20214 (N_20214,N_19957,N_19893);
nor U20215 (N_20215,N_19780,N_19925);
or U20216 (N_20216,N_19831,N_19910);
nand U20217 (N_20217,N_19798,N_19952);
nor U20218 (N_20218,N_19854,N_19846);
or U20219 (N_20219,N_19925,N_19818);
and U20220 (N_20220,N_19760,N_19923);
nor U20221 (N_20221,N_19847,N_19855);
nor U20222 (N_20222,N_19849,N_19964);
nor U20223 (N_20223,N_19923,N_19908);
xor U20224 (N_20224,N_19905,N_19788);
nand U20225 (N_20225,N_19967,N_19792);
nand U20226 (N_20226,N_19806,N_19983);
nor U20227 (N_20227,N_19773,N_19751);
and U20228 (N_20228,N_19990,N_19960);
and U20229 (N_20229,N_19777,N_19792);
or U20230 (N_20230,N_19868,N_19850);
nor U20231 (N_20231,N_19826,N_19964);
or U20232 (N_20232,N_19762,N_19838);
and U20233 (N_20233,N_19978,N_19981);
nand U20234 (N_20234,N_19884,N_19782);
xor U20235 (N_20235,N_19755,N_19761);
xor U20236 (N_20236,N_19793,N_19951);
nor U20237 (N_20237,N_19967,N_19915);
nor U20238 (N_20238,N_19991,N_19900);
xor U20239 (N_20239,N_19926,N_19785);
or U20240 (N_20240,N_19904,N_19758);
nand U20241 (N_20241,N_19822,N_19952);
and U20242 (N_20242,N_19774,N_19974);
xnor U20243 (N_20243,N_19850,N_19893);
and U20244 (N_20244,N_19924,N_19883);
nand U20245 (N_20245,N_19786,N_19920);
nand U20246 (N_20246,N_19821,N_19953);
nand U20247 (N_20247,N_19830,N_19992);
nor U20248 (N_20248,N_19765,N_19927);
nor U20249 (N_20249,N_19810,N_19912);
or U20250 (N_20250,N_20247,N_20236);
and U20251 (N_20251,N_20178,N_20158);
nor U20252 (N_20252,N_20095,N_20148);
and U20253 (N_20253,N_20223,N_20219);
nand U20254 (N_20254,N_20221,N_20090);
nand U20255 (N_20255,N_20170,N_20103);
nand U20256 (N_20256,N_20101,N_20084);
or U20257 (N_20257,N_20194,N_20150);
nor U20258 (N_20258,N_20065,N_20210);
and U20259 (N_20259,N_20208,N_20098);
or U20260 (N_20260,N_20079,N_20193);
and U20261 (N_20261,N_20238,N_20243);
and U20262 (N_20262,N_20212,N_20138);
and U20263 (N_20263,N_20032,N_20112);
nand U20264 (N_20264,N_20015,N_20056);
xnor U20265 (N_20265,N_20020,N_20126);
nand U20266 (N_20266,N_20190,N_20191);
nor U20267 (N_20267,N_20063,N_20043);
or U20268 (N_20268,N_20041,N_20174);
nor U20269 (N_20269,N_20017,N_20083);
and U20270 (N_20270,N_20025,N_20048);
nor U20271 (N_20271,N_20038,N_20012);
and U20272 (N_20272,N_20100,N_20119);
nand U20273 (N_20273,N_20022,N_20155);
nor U20274 (N_20274,N_20124,N_20143);
and U20275 (N_20275,N_20147,N_20152);
and U20276 (N_20276,N_20005,N_20241);
and U20277 (N_20277,N_20206,N_20185);
or U20278 (N_20278,N_20078,N_20107);
and U20279 (N_20279,N_20237,N_20102);
or U20280 (N_20280,N_20245,N_20196);
nor U20281 (N_20281,N_20077,N_20044);
or U20282 (N_20282,N_20004,N_20104);
nand U20283 (N_20283,N_20207,N_20091);
or U20284 (N_20284,N_20156,N_20135);
nand U20285 (N_20285,N_20199,N_20085);
nand U20286 (N_20286,N_20159,N_20074);
nand U20287 (N_20287,N_20042,N_20113);
nand U20288 (N_20288,N_20198,N_20233);
xnor U20289 (N_20289,N_20209,N_20172);
or U20290 (N_20290,N_20202,N_20160);
nand U20291 (N_20291,N_20062,N_20034);
or U20292 (N_20292,N_20176,N_20000);
nand U20293 (N_20293,N_20059,N_20087);
nor U20294 (N_20294,N_20089,N_20018);
or U20295 (N_20295,N_20184,N_20224);
nor U20296 (N_20296,N_20030,N_20167);
nand U20297 (N_20297,N_20016,N_20248);
or U20298 (N_20298,N_20227,N_20175);
or U20299 (N_20299,N_20226,N_20029);
or U20300 (N_20300,N_20009,N_20076);
nand U20301 (N_20301,N_20118,N_20021);
nor U20302 (N_20302,N_20144,N_20181);
and U20303 (N_20303,N_20055,N_20123);
nor U20304 (N_20304,N_20067,N_20052);
nand U20305 (N_20305,N_20211,N_20186);
or U20306 (N_20306,N_20234,N_20114);
and U20307 (N_20307,N_20070,N_20080);
and U20308 (N_20308,N_20157,N_20109);
and U20309 (N_20309,N_20133,N_20036);
and U20310 (N_20310,N_20249,N_20235);
and U20311 (N_20311,N_20239,N_20180);
nor U20312 (N_20312,N_20242,N_20068);
nor U20313 (N_20313,N_20115,N_20128);
and U20314 (N_20314,N_20117,N_20131);
or U20315 (N_20315,N_20195,N_20140);
nor U20316 (N_20316,N_20086,N_20240);
and U20317 (N_20317,N_20137,N_20028);
nand U20318 (N_20318,N_20054,N_20228);
and U20319 (N_20319,N_20058,N_20153);
nand U20320 (N_20320,N_20040,N_20183);
nor U20321 (N_20321,N_20057,N_20099);
or U20322 (N_20322,N_20106,N_20244);
nand U20323 (N_20323,N_20035,N_20093);
and U20324 (N_20324,N_20069,N_20072);
nor U20325 (N_20325,N_20121,N_20229);
xor U20326 (N_20326,N_20007,N_20051);
or U20327 (N_20327,N_20218,N_20164);
nand U20328 (N_20328,N_20033,N_20073);
nor U20329 (N_20329,N_20066,N_20116);
nand U20330 (N_20330,N_20203,N_20081);
nand U20331 (N_20331,N_20154,N_20162);
nor U20332 (N_20332,N_20097,N_20142);
nand U20333 (N_20333,N_20061,N_20125);
nand U20334 (N_20334,N_20204,N_20075);
or U20335 (N_20335,N_20166,N_20096);
nor U20336 (N_20336,N_20039,N_20006);
nand U20337 (N_20337,N_20037,N_20111);
or U20338 (N_20338,N_20214,N_20047);
nor U20339 (N_20339,N_20187,N_20008);
nor U20340 (N_20340,N_20002,N_20171);
nand U20341 (N_20341,N_20088,N_20082);
and U20342 (N_20342,N_20134,N_20094);
nor U20343 (N_20343,N_20023,N_20231);
nand U20344 (N_20344,N_20192,N_20188);
or U20345 (N_20345,N_20136,N_20139);
nor U20346 (N_20346,N_20230,N_20060);
and U20347 (N_20347,N_20163,N_20011);
nand U20348 (N_20348,N_20216,N_20013);
nor U20349 (N_20349,N_20014,N_20046);
and U20350 (N_20350,N_20177,N_20129);
nor U20351 (N_20351,N_20132,N_20092);
or U20352 (N_20352,N_20003,N_20105);
or U20353 (N_20353,N_20049,N_20165);
or U20354 (N_20354,N_20120,N_20026);
or U20355 (N_20355,N_20168,N_20189);
or U20356 (N_20356,N_20045,N_20031);
nand U20357 (N_20357,N_20161,N_20232);
xor U20358 (N_20358,N_20200,N_20217);
or U20359 (N_20359,N_20225,N_20053);
or U20360 (N_20360,N_20205,N_20169);
nor U20361 (N_20361,N_20215,N_20149);
or U20362 (N_20362,N_20130,N_20122);
xnor U20363 (N_20363,N_20213,N_20071);
and U20364 (N_20364,N_20019,N_20182);
or U20365 (N_20365,N_20201,N_20024);
nor U20366 (N_20366,N_20127,N_20108);
nand U20367 (N_20367,N_20001,N_20010);
and U20368 (N_20368,N_20050,N_20064);
or U20369 (N_20369,N_20179,N_20027);
xor U20370 (N_20370,N_20110,N_20220);
nor U20371 (N_20371,N_20173,N_20222);
nor U20372 (N_20372,N_20141,N_20146);
and U20373 (N_20373,N_20246,N_20145);
or U20374 (N_20374,N_20197,N_20151);
or U20375 (N_20375,N_20024,N_20220);
and U20376 (N_20376,N_20040,N_20091);
nand U20377 (N_20377,N_20093,N_20246);
xor U20378 (N_20378,N_20140,N_20201);
nand U20379 (N_20379,N_20107,N_20226);
or U20380 (N_20380,N_20199,N_20219);
or U20381 (N_20381,N_20073,N_20199);
nor U20382 (N_20382,N_20205,N_20193);
nor U20383 (N_20383,N_20001,N_20113);
nor U20384 (N_20384,N_20226,N_20137);
nor U20385 (N_20385,N_20105,N_20160);
or U20386 (N_20386,N_20248,N_20184);
nand U20387 (N_20387,N_20013,N_20042);
nor U20388 (N_20388,N_20181,N_20172);
nand U20389 (N_20389,N_20107,N_20166);
or U20390 (N_20390,N_20108,N_20137);
nand U20391 (N_20391,N_20087,N_20155);
nand U20392 (N_20392,N_20183,N_20015);
or U20393 (N_20393,N_20247,N_20091);
and U20394 (N_20394,N_20024,N_20130);
nor U20395 (N_20395,N_20223,N_20214);
and U20396 (N_20396,N_20154,N_20057);
nand U20397 (N_20397,N_20074,N_20175);
nor U20398 (N_20398,N_20183,N_20132);
nand U20399 (N_20399,N_20246,N_20094);
nor U20400 (N_20400,N_20010,N_20184);
nand U20401 (N_20401,N_20148,N_20131);
nand U20402 (N_20402,N_20232,N_20060);
nor U20403 (N_20403,N_20165,N_20196);
xnor U20404 (N_20404,N_20175,N_20206);
nand U20405 (N_20405,N_20156,N_20070);
and U20406 (N_20406,N_20239,N_20166);
nand U20407 (N_20407,N_20034,N_20199);
and U20408 (N_20408,N_20021,N_20017);
nand U20409 (N_20409,N_20092,N_20212);
or U20410 (N_20410,N_20030,N_20187);
nand U20411 (N_20411,N_20026,N_20165);
xnor U20412 (N_20412,N_20052,N_20238);
or U20413 (N_20413,N_20011,N_20233);
or U20414 (N_20414,N_20046,N_20010);
nor U20415 (N_20415,N_20204,N_20244);
nand U20416 (N_20416,N_20159,N_20053);
or U20417 (N_20417,N_20091,N_20249);
nand U20418 (N_20418,N_20001,N_20025);
nor U20419 (N_20419,N_20178,N_20013);
and U20420 (N_20420,N_20200,N_20102);
nor U20421 (N_20421,N_20086,N_20149);
nand U20422 (N_20422,N_20223,N_20242);
nor U20423 (N_20423,N_20195,N_20248);
nand U20424 (N_20424,N_20126,N_20121);
or U20425 (N_20425,N_20082,N_20018);
and U20426 (N_20426,N_20215,N_20194);
and U20427 (N_20427,N_20023,N_20162);
nand U20428 (N_20428,N_20080,N_20037);
nand U20429 (N_20429,N_20096,N_20032);
nand U20430 (N_20430,N_20194,N_20014);
nand U20431 (N_20431,N_20225,N_20167);
or U20432 (N_20432,N_20090,N_20193);
or U20433 (N_20433,N_20110,N_20223);
xnor U20434 (N_20434,N_20005,N_20004);
and U20435 (N_20435,N_20023,N_20095);
or U20436 (N_20436,N_20140,N_20026);
and U20437 (N_20437,N_20232,N_20044);
and U20438 (N_20438,N_20109,N_20183);
xor U20439 (N_20439,N_20206,N_20013);
or U20440 (N_20440,N_20014,N_20211);
and U20441 (N_20441,N_20075,N_20235);
nand U20442 (N_20442,N_20228,N_20109);
nor U20443 (N_20443,N_20061,N_20229);
and U20444 (N_20444,N_20030,N_20171);
nor U20445 (N_20445,N_20070,N_20149);
and U20446 (N_20446,N_20013,N_20054);
nor U20447 (N_20447,N_20153,N_20003);
nand U20448 (N_20448,N_20225,N_20029);
and U20449 (N_20449,N_20158,N_20142);
nand U20450 (N_20450,N_20191,N_20056);
nor U20451 (N_20451,N_20160,N_20052);
and U20452 (N_20452,N_20167,N_20065);
xnor U20453 (N_20453,N_20240,N_20197);
nor U20454 (N_20454,N_20032,N_20144);
or U20455 (N_20455,N_20031,N_20010);
nor U20456 (N_20456,N_20077,N_20014);
or U20457 (N_20457,N_20064,N_20153);
nand U20458 (N_20458,N_20164,N_20191);
and U20459 (N_20459,N_20079,N_20197);
nand U20460 (N_20460,N_20200,N_20012);
nand U20461 (N_20461,N_20169,N_20131);
nor U20462 (N_20462,N_20012,N_20212);
nor U20463 (N_20463,N_20158,N_20224);
or U20464 (N_20464,N_20154,N_20010);
and U20465 (N_20465,N_20017,N_20143);
and U20466 (N_20466,N_20149,N_20239);
nand U20467 (N_20467,N_20233,N_20098);
and U20468 (N_20468,N_20075,N_20096);
and U20469 (N_20469,N_20216,N_20101);
nor U20470 (N_20470,N_20170,N_20038);
nand U20471 (N_20471,N_20156,N_20019);
nand U20472 (N_20472,N_20049,N_20013);
and U20473 (N_20473,N_20070,N_20147);
nand U20474 (N_20474,N_20098,N_20226);
nor U20475 (N_20475,N_20221,N_20123);
nand U20476 (N_20476,N_20232,N_20081);
xnor U20477 (N_20477,N_20201,N_20105);
or U20478 (N_20478,N_20219,N_20041);
nor U20479 (N_20479,N_20040,N_20142);
or U20480 (N_20480,N_20032,N_20099);
and U20481 (N_20481,N_20153,N_20171);
and U20482 (N_20482,N_20097,N_20010);
or U20483 (N_20483,N_20124,N_20110);
or U20484 (N_20484,N_20010,N_20038);
and U20485 (N_20485,N_20011,N_20199);
nor U20486 (N_20486,N_20210,N_20023);
nor U20487 (N_20487,N_20207,N_20028);
nand U20488 (N_20488,N_20099,N_20159);
nor U20489 (N_20489,N_20131,N_20173);
nor U20490 (N_20490,N_20032,N_20014);
nand U20491 (N_20491,N_20162,N_20239);
or U20492 (N_20492,N_20179,N_20127);
nor U20493 (N_20493,N_20217,N_20144);
or U20494 (N_20494,N_20240,N_20068);
and U20495 (N_20495,N_20237,N_20008);
nor U20496 (N_20496,N_20188,N_20133);
nor U20497 (N_20497,N_20062,N_20116);
or U20498 (N_20498,N_20184,N_20078);
nor U20499 (N_20499,N_20162,N_20090);
nor U20500 (N_20500,N_20383,N_20331);
nor U20501 (N_20501,N_20439,N_20353);
xnor U20502 (N_20502,N_20250,N_20339);
and U20503 (N_20503,N_20387,N_20262);
nor U20504 (N_20504,N_20451,N_20254);
xnor U20505 (N_20505,N_20462,N_20269);
nand U20506 (N_20506,N_20258,N_20295);
nand U20507 (N_20507,N_20329,N_20290);
nand U20508 (N_20508,N_20322,N_20311);
or U20509 (N_20509,N_20412,N_20498);
or U20510 (N_20510,N_20417,N_20463);
nand U20511 (N_20511,N_20313,N_20285);
xnor U20512 (N_20512,N_20281,N_20493);
or U20513 (N_20513,N_20264,N_20275);
nor U20514 (N_20514,N_20409,N_20489);
nor U20515 (N_20515,N_20482,N_20459);
or U20516 (N_20516,N_20455,N_20468);
and U20517 (N_20517,N_20450,N_20461);
and U20518 (N_20518,N_20321,N_20346);
nand U20519 (N_20519,N_20465,N_20328);
nor U20520 (N_20520,N_20305,N_20288);
or U20521 (N_20521,N_20298,N_20272);
and U20522 (N_20522,N_20415,N_20314);
nand U20523 (N_20523,N_20278,N_20271);
and U20524 (N_20524,N_20361,N_20429);
nor U20525 (N_20525,N_20408,N_20471);
xor U20526 (N_20526,N_20464,N_20484);
nor U20527 (N_20527,N_20304,N_20357);
nand U20528 (N_20528,N_20384,N_20293);
and U20529 (N_20529,N_20265,N_20467);
xnor U20530 (N_20530,N_20418,N_20443);
and U20531 (N_20531,N_20347,N_20479);
nand U20532 (N_20532,N_20359,N_20444);
nand U20533 (N_20533,N_20323,N_20385);
nand U20534 (N_20534,N_20363,N_20472);
xor U20535 (N_20535,N_20381,N_20326);
nand U20536 (N_20536,N_20488,N_20277);
or U20537 (N_20537,N_20431,N_20343);
and U20538 (N_20538,N_20406,N_20414);
or U20539 (N_20539,N_20376,N_20327);
xor U20540 (N_20540,N_20342,N_20437);
nor U20541 (N_20541,N_20452,N_20380);
nand U20542 (N_20542,N_20396,N_20394);
xor U20543 (N_20543,N_20318,N_20338);
and U20544 (N_20544,N_20286,N_20393);
and U20545 (N_20545,N_20485,N_20320);
and U20546 (N_20546,N_20292,N_20370);
and U20547 (N_20547,N_20354,N_20345);
and U20548 (N_20548,N_20411,N_20299);
nand U20549 (N_20549,N_20268,N_20270);
or U20550 (N_20550,N_20274,N_20495);
or U20551 (N_20551,N_20497,N_20438);
xnor U20552 (N_20552,N_20366,N_20340);
or U20553 (N_20553,N_20282,N_20392);
xnor U20554 (N_20554,N_20317,N_20373);
nor U20555 (N_20555,N_20441,N_20294);
or U20556 (N_20556,N_20424,N_20447);
nand U20557 (N_20557,N_20445,N_20350);
nand U20558 (N_20558,N_20413,N_20255);
or U20559 (N_20559,N_20378,N_20432);
nor U20560 (N_20560,N_20422,N_20263);
and U20561 (N_20561,N_20352,N_20430);
and U20562 (N_20562,N_20435,N_20402);
or U20563 (N_20563,N_20391,N_20351);
xnor U20564 (N_20564,N_20344,N_20404);
nor U20565 (N_20565,N_20315,N_20284);
xnor U20566 (N_20566,N_20316,N_20401);
nand U20567 (N_20567,N_20266,N_20349);
nand U20568 (N_20568,N_20480,N_20446);
nor U20569 (N_20569,N_20454,N_20300);
nand U20570 (N_20570,N_20436,N_20466);
or U20571 (N_20571,N_20302,N_20358);
and U20572 (N_20572,N_20458,N_20460);
nand U20573 (N_20573,N_20390,N_20473);
and U20574 (N_20574,N_20306,N_20478);
nand U20575 (N_20575,N_20389,N_20253);
and U20576 (N_20576,N_20362,N_20388);
and U20577 (N_20577,N_20379,N_20279);
and U20578 (N_20578,N_20453,N_20457);
or U20579 (N_20579,N_20371,N_20470);
nor U20580 (N_20580,N_20398,N_20334);
xnor U20581 (N_20581,N_20260,N_20407);
nand U20582 (N_20582,N_20337,N_20309);
nor U20583 (N_20583,N_20487,N_20368);
or U20584 (N_20584,N_20369,N_20259);
and U20585 (N_20585,N_20427,N_20297);
nor U20586 (N_20586,N_20419,N_20301);
nand U20587 (N_20587,N_20416,N_20367);
and U20588 (N_20588,N_20426,N_20377);
nand U20589 (N_20589,N_20421,N_20335);
and U20590 (N_20590,N_20273,N_20499);
nand U20591 (N_20591,N_20423,N_20481);
nand U20592 (N_20592,N_20486,N_20490);
nand U20593 (N_20593,N_20375,N_20374);
or U20594 (N_20594,N_20397,N_20469);
or U20595 (N_20595,N_20434,N_20356);
nor U20596 (N_20596,N_20477,N_20496);
nand U20597 (N_20597,N_20448,N_20494);
or U20598 (N_20598,N_20251,N_20324);
xor U20599 (N_20599,N_20330,N_20425);
and U20600 (N_20600,N_20267,N_20355);
or U20601 (N_20601,N_20325,N_20476);
and U20602 (N_20602,N_20372,N_20483);
xnor U20603 (N_20603,N_20308,N_20287);
xnor U20604 (N_20604,N_20283,N_20310);
nand U20605 (N_20605,N_20365,N_20410);
and U20606 (N_20606,N_20492,N_20399);
nor U20607 (N_20607,N_20348,N_20261);
or U20608 (N_20608,N_20395,N_20307);
nand U20609 (N_20609,N_20341,N_20440);
nand U20610 (N_20610,N_20475,N_20420);
or U20611 (N_20611,N_20296,N_20289);
xor U20612 (N_20612,N_20386,N_20291);
and U20613 (N_20613,N_20428,N_20491);
or U20614 (N_20614,N_20360,N_20364);
or U20615 (N_20615,N_20280,N_20257);
and U20616 (N_20616,N_20403,N_20332);
nand U20617 (N_20617,N_20319,N_20256);
and U20618 (N_20618,N_20400,N_20442);
nand U20619 (N_20619,N_20252,N_20449);
nand U20620 (N_20620,N_20433,N_20336);
nor U20621 (N_20621,N_20312,N_20405);
nand U20622 (N_20622,N_20333,N_20276);
xor U20623 (N_20623,N_20382,N_20456);
xnor U20624 (N_20624,N_20303,N_20474);
or U20625 (N_20625,N_20370,N_20407);
or U20626 (N_20626,N_20356,N_20282);
or U20627 (N_20627,N_20292,N_20435);
and U20628 (N_20628,N_20476,N_20458);
nor U20629 (N_20629,N_20367,N_20342);
nand U20630 (N_20630,N_20430,N_20374);
nor U20631 (N_20631,N_20415,N_20408);
or U20632 (N_20632,N_20376,N_20449);
or U20633 (N_20633,N_20445,N_20286);
or U20634 (N_20634,N_20392,N_20426);
and U20635 (N_20635,N_20340,N_20423);
or U20636 (N_20636,N_20496,N_20317);
xnor U20637 (N_20637,N_20492,N_20290);
or U20638 (N_20638,N_20494,N_20386);
and U20639 (N_20639,N_20396,N_20418);
xor U20640 (N_20640,N_20385,N_20380);
nand U20641 (N_20641,N_20491,N_20421);
or U20642 (N_20642,N_20343,N_20419);
xor U20643 (N_20643,N_20288,N_20499);
nand U20644 (N_20644,N_20292,N_20461);
nor U20645 (N_20645,N_20441,N_20283);
and U20646 (N_20646,N_20331,N_20461);
and U20647 (N_20647,N_20283,N_20253);
nor U20648 (N_20648,N_20262,N_20428);
nor U20649 (N_20649,N_20323,N_20431);
nor U20650 (N_20650,N_20359,N_20396);
nand U20651 (N_20651,N_20396,N_20256);
xnor U20652 (N_20652,N_20409,N_20396);
or U20653 (N_20653,N_20436,N_20291);
xnor U20654 (N_20654,N_20299,N_20341);
nand U20655 (N_20655,N_20331,N_20480);
and U20656 (N_20656,N_20446,N_20468);
or U20657 (N_20657,N_20377,N_20393);
or U20658 (N_20658,N_20305,N_20477);
nand U20659 (N_20659,N_20316,N_20373);
and U20660 (N_20660,N_20346,N_20306);
or U20661 (N_20661,N_20407,N_20326);
or U20662 (N_20662,N_20298,N_20269);
nand U20663 (N_20663,N_20352,N_20305);
nand U20664 (N_20664,N_20402,N_20389);
and U20665 (N_20665,N_20491,N_20436);
and U20666 (N_20666,N_20381,N_20416);
or U20667 (N_20667,N_20443,N_20337);
nor U20668 (N_20668,N_20434,N_20288);
nand U20669 (N_20669,N_20447,N_20286);
and U20670 (N_20670,N_20369,N_20436);
nand U20671 (N_20671,N_20315,N_20448);
or U20672 (N_20672,N_20253,N_20401);
xor U20673 (N_20673,N_20335,N_20345);
and U20674 (N_20674,N_20266,N_20466);
and U20675 (N_20675,N_20450,N_20267);
nor U20676 (N_20676,N_20295,N_20333);
and U20677 (N_20677,N_20280,N_20290);
or U20678 (N_20678,N_20460,N_20408);
xor U20679 (N_20679,N_20300,N_20321);
nand U20680 (N_20680,N_20492,N_20421);
or U20681 (N_20681,N_20347,N_20459);
or U20682 (N_20682,N_20324,N_20264);
nand U20683 (N_20683,N_20416,N_20290);
nor U20684 (N_20684,N_20382,N_20481);
or U20685 (N_20685,N_20451,N_20436);
nand U20686 (N_20686,N_20370,N_20339);
nand U20687 (N_20687,N_20439,N_20254);
or U20688 (N_20688,N_20348,N_20475);
nor U20689 (N_20689,N_20296,N_20342);
or U20690 (N_20690,N_20469,N_20499);
nand U20691 (N_20691,N_20495,N_20257);
or U20692 (N_20692,N_20350,N_20462);
and U20693 (N_20693,N_20291,N_20277);
or U20694 (N_20694,N_20377,N_20321);
nand U20695 (N_20695,N_20380,N_20494);
nand U20696 (N_20696,N_20440,N_20256);
or U20697 (N_20697,N_20258,N_20418);
nor U20698 (N_20698,N_20432,N_20334);
xnor U20699 (N_20699,N_20359,N_20303);
and U20700 (N_20700,N_20339,N_20303);
and U20701 (N_20701,N_20382,N_20375);
or U20702 (N_20702,N_20310,N_20445);
nor U20703 (N_20703,N_20434,N_20404);
or U20704 (N_20704,N_20378,N_20466);
and U20705 (N_20705,N_20429,N_20404);
nand U20706 (N_20706,N_20479,N_20331);
nand U20707 (N_20707,N_20258,N_20496);
xor U20708 (N_20708,N_20449,N_20425);
or U20709 (N_20709,N_20397,N_20379);
and U20710 (N_20710,N_20430,N_20423);
and U20711 (N_20711,N_20314,N_20322);
nor U20712 (N_20712,N_20393,N_20363);
or U20713 (N_20713,N_20411,N_20387);
nand U20714 (N_20714,N_20497,N_20393);
nor U20715 (N_20715,N_20269,N_20367);
xor U20716 (N_20716,N_20259,N_20427);
nand U20717 (N_20717,N_20382,N_20430);
and U20718 (N_20718,N_20253,N_20337);
xnor U20719 (N_20719,N_20357,N_20303);
nand U20720 (N_20720,N_20360,N_20497);
or U20721 (N_20721,N_20339,N_20381);
nand U20722 (N_20722,N_20462,N_20490);
and U20723 (N_20723,N_20320,N_20417);
xnor U20724 (N_20724,N_20401,N_20351);
xor U20725 (N_20725,N_20276,N_20437);
nor U20726 (N_20726,N_20443,N_20312);
xor U20727 (N_20727,N_20432,N_20358);
nor U20728 (N_20728,N_20431,N_20314);
or U20729 (N_20729,N_20368,N_20254);
and U20730 (N_20730,N_20360,N_20460);
nand U20731 (N_20731,N_20450,N_20418);
or U20732 (N_20732,N_20382,N_20462);
and U20733 (N_20733,N_20491,N_20269);
xnor U20734 (N_20734,N_20260,N_20459);
and U20735 (N_20735,N_20270,N_20427);
xnor U20736 (N_20736,N_20461,N_20350);
and U20737 (N_20737,N_20361,N_20309);
nor U20738 (N_20738,N_20265,N_20432);
nand U20739 (N_20739,N_20463,N_20427);
and U20740 (N_20740,N_20378,N_20383);
or U20741 (N_20741,N_20400,N_20342);
nand U20742 (N_20742,N_20480,N_20379);
nor U20743 (N_20743,N_20269,N_20492);
and U20744 (N_20744,N_20460,N_20465);
nor U20745 (N_20745,N_20442,N_20459);
nand U20746 (N_20746,N_20378,N_20414);
nand U20747 (N_20747,N_20493,N_20259);
and U20748 (N_20748,N_20255,N_20456);
xor U20749 (N_20749,N_20261,N_20293);
or U20750 (N_20750,N_20646,N_20508);
xnor U20751 (N_20751,N_20665,N_20577);
or U20752 (N_20752,N_20651,N_20582);
nand U20753 (N_20753,N_20562,N_20624);
nor U20754 (N_20754,N_20587,N_20679);
nand U20755 (N_20755,N_20553,N_20689);
xor U20756 (N_20756,N_20736,N_20653);
nand U20757 (N_20757,N_20709,N_20571);
and U20758 (N_20758,N_20724,N_20563);
or U20759 (N_20759,N_20639,N_20732);
nor U20760 (N_20760,N_20513,N_20502);
or U20761 (N_20761,N_20666,N_20680);
nor U20762 (N_20762,N_20602,N_20578);
and U20763 (N_20763,N_20550,N_20500);
or U20764 (N_20764,N_20717,N_20668);
or U20765 (N_20765,N_20609,N_20641);
nand U20766 (N_20766,N_20711,N_20735);
nand U20767 (N_20767,N_20524,N_20740);
nor U20768 (N_20768,N_20628,N_20659);
nor U20769 (N_20769,N_20600,N_20565);
nand U20770 (N_20770,N_20688,N_20716);
xor U20771 (N_20771,N_20597,N_20517);
and U20772 (N_20772,N_20743,N_20595);
nor U20773 (N_20773,N_20621,N_20534);
nand U20774 (N_20774,N_20612,N_20503);
nand U20775 (N_20775,N_20625,N_20521);
nor U20776 (N_20776,N_20674,N_20672);
or U20777 (N_20777,N_20731,N_20685);
nand U20778 (N_20778,N_20719,N_20615);
nor U20779 (N_20779,N_20616,N_20580);
nor U20780 (N_20780,N_20671,N_20722);
nor U20781 (N_20781,N_20699,N_20585);
and U20782 (N_20782,N_20686,N_20648);
and U20783 (N_20783,N_20566,N_20569);
and U20784 (N_20784,N_20710,N_20739);
nor U20785 (N_20785,N_20538,N_20734);
xnor U20786 (N_20786,N_20670,N_20726);
nand U20787 (N_20787,N_20532,N_20526);
or U20788 (N_20788,N_20638,N_20733);
nand U20789 (N_20789,N_20525,N_20505);
nor U20790 (N_20790,N_20515,N_20748);
xnor U20791 (N_20791,N_20570,N_20511);
xnor U20792 (N_20792,N_20558,N_20682);
or U20793 (N_20793,N_20542,N_20703);
nand U20794 (N_20794,N_20541,N_20554);
nor U20795 (N_20795,N_20634,N_20694);
and U20796 (N_20796,N_20529,N_20676);
nand U20797 (N_20797,N_20627,N_20539);
or U20798 (N_20798,N_20608,N_20592);
and U20799 (N_20799,N_20512,N_20556);
nand U20800 (N_20800,N_20697,N_20714);
and U20801 (N_20801,N_20528,N_20746);
nor U20802 (N_20802,N_20619,N_20579);
nand U20803 (N_20803,N_20728,N_20663);
nor U20804 (N_20804,N_20721,N_20533);
and U20805 (N_20805,N_20509,N_20588);
or U20806 (N_20806,N_20667,N_20705);
and U20807 (N_20807,N_20557,N_20604);
and U20808 (N_20808,N_20530,N_20594);
or U20809 (N_20809,N_20544,N_20702);
and U20810 (N_20810,N_20549,N_20729);
or U20811 (N_20811,N_20637,N_20575);
nor U20812 (N_20812,N_20555,N_20738);
nand U20813 (N_20813,N_20617,N_20650);
nand U20814 (N_20814,N_20715,N_20560);
and U20815 (N_20815,N_20684,N_20572);
or U20816 (N_20816,N_20603,N_20633);
or U20817 (N_20817,N_20713,N_20626);
and U20818 (N_20818,N_20654,N_20547);
nand U20819 (N_20819,N_20606,N_20573);
nand U20820 (N_20820,N_20708,N_20749);
nand U20821 (N_20821,N_20652,N_20581);
nor U20822 (N_20822,N_20723,N_20744);
nand U20823 (N_20823,N_20546,N_20564);
xor U20824 (N_20824,N_20683,N_20506);
nor U20825 (N_20825,N_20501,N_20656);
nand U20826 (N_20826,N_20605,N_20593);
nand U20827 (N_20827,N_20681,N_20698);
nor U20828 (N_20828,N_20640,N_20507);
or U20829 (N_20829,N_20536,N_20718);
nor U20830 (N_20830,N_20618,N_20590);
xnor U20831 (N_20831,N_20601,N_20559);
nor U20832 (N_20832,N_20631,N_20504);
xnor U20833 (N_20833,N_20518,N_20620);
nand U20834 (N_20834,N_20540,N_20584);
nand U20835 (N_20835,N_20636,N_20707);
xor U20836 (N_20836,N_20704,N_20576);
and U20837 (N_20837,N_20516,N_20531);
or U20838 (N_20838,N_20611,N_20589);
nor U20839 (N_20839,N_20664,N_20690);
and U20840 (N_20840,N_20586,N_20527);
and U20841 (N_20841,N_20693,N_20510);
nor U20842 (N_20842,N_20645,N_20519);
nor U20843 (N_20843,N_20630,N_20742);
nand U20844 (N_20844,N_20523,N_20548);
or U20845 (N_20845,N_20535,N_20658);
or U20846 (N_20846,N_20644,N_20552);
nand U20847 (N_20847,N_20632,N_20675);
nand U20848 (N_20848,N_20591,N_20720);
nor U20849 (N_20849,N_20706,N_20561);
nor U20850 (N_20850,N_20545,N_20551);
nor U20851 (N_20851,N_20730,N_20607);
nor U20852 (N_20852,N_20747,N_20522);
and U20853 (N_20853,N_20691,N_20655);
xor U20854 (N_20854,N_20673,N_20614);
nor U20855 (N_20855,N_20622,N_20568);
nand U20856 (N_20856,N_20635,N_20647);
and U20857 (N_20857,N_20537,N_20649);
nor U20858 (N_20858,N_20701,N_20613);
nand U20859 (N_20859,N_20629,N_20737);
and U20860 (N_20860,N_20574,N_20662);
nand U20861 (N_20861,N_20700,N_20583);
nand U20862 (N_20862,N_20543,N_20623);
nand U20863 (N_20863,N_20661,N_20669);
nor U20864 (N_20864,N_20695,N_20696);
nor U20865 (N_20865,N_20596,N_20727);
xnor U20866 (N_20866,N_20610,N_20567);
nand U20867 (N_20867,N_20677,N_20657);
or U20868 (N_20868,N_20712,N_20692);
xnor U20869 (N_20869,N_20643,N_20642);
or U20870 (N_20870,N_20678,N_20687);
nor U20871 (N_20871,N_20660,N_20598);
nor U20872 (N_20872,N_20520,N_20741);
nor U20873 (N_20873,N_20725,N_20745);
nor U20874 (N_20874,N_20599,N_20514);
nor U20875 (N_20875,N_20666,N_20716);
nand U20876 (N_20876,N_20706,N_20730);
or U20877 (N_20877,N_20724,N_20605);
or U20878 (N_20878,N_20658,N_20578);
and U20879 (N_20879,N_20704,N_20625);
nand U20880 (N_20880,N_20639,N_20721);
nor U20881 (N_20881,N_20558,N_20727);
or U20882 (N_20882,N_20573,N_20597);
nor U20883 (N_20883,N_20639,N_20567);
nand U20884 (N_20884,N_20528,N_20521);
nand U20885 (N_20885,N_20514,N_20738);
nor U20886 (N_20886,N_20602,N_20554);
and U20887 (N_20887,N_20507,N_20683);
nand U20888 (N_20888,N_20559,N_20573);
or U20889 (N_20889,N_20685,N_20536);
nand U20890 (N_20890,N_20522,N_20737);
nand U20891 (N_20891,N_20501,N_20531);
nor U20892 (N_20892,N_20561,N_20641);
or U20893 (N_20893,N_20595,N_20584);
or U20894 (N_20894,N_20516,N_20525);
or U20895 (N_20895,N_20561,N_20688);
nand U20896 (N_20896,N_20504,N_20577);
nand U20897 (N_20897,N_20546,N_20645);
or U20898 (N_20898,N_20687,N_20532);
nand U20899 (N_20899,N_20523,N_20671);
and U20900 (N_20900,N_20749,N_20510);
nand U20901 (N_20901,N_20749,N_20529);
nor U20902 (N_20902,N_20634,N_20528);
and U20903 (N_20903,N_20540,N_20599);
and U20904 (N_20904,N_20541,N_20532);
and U20905 (N_20905,N_20731,N_20584);
nor U20906 (N_20906,N_20601,N_20704);
nand U20907 (N_20907,N_20546,N_20737);
nor U20908 (N_20908,N_20741,N_20510);
nand U20909 (N_20909,N_20540,N_20588);
or U20910 (N_20910,N_20585,N_20548);
nor U20911 (N_20911,N_20690,N_20714);
nor U20912 (N_20912,N_20671,N_20543);
or U20913 (N_20913,N_20661,N_20716);
xor U20914 (N_20914,N_20682,N_20699);
nand U20915 (N_20915,N_20571,N_20614);
nor U20916 (N_20916,N_20736,N_20665);
nand U20917 (N_20917,N_20636,N_20534);
and U20918 (N_20918,N_20609,N_20688);
nand U20919 (N_20919,N_20550,N_20663);
nor U20920 (N_20920,N_20510,N_20540);
or U20921 (N_20921,N_20705,N_20690);
nor U20922 (N_20922,N_20559,N_20670);
nand U20923 (N_20923,N_20695,N_20700);
nand U20924 (N_20924,N_20686,N_20664);
or U20925 (N_20925,N_20667,N_20567);
nand U20926 (N_20926,N_20535,N_20630);
nor U20927 (N_20927,N_20508,N_20643);
and U20928 (N_20928,N_20745,N_20672);
nor U20929 (N_20929,N_20718,N_20546);
nand U20930 (N_20930,N_20614,N_20501);
or U20931 (N_20931,N_20647,N_20628);
nor U20932 (N_20932,N_20628,N_20624);
nor U20933 (N_20933,N_20659,N_20558);
or U20934 (N_20934,N_20698,N_20741);
and U20935 (N_20935,N_20745,N_20583);
xor U20936 (N_20936,N_20652,N_20720);
or U20937 (N_20937,N_20564,N_20686);
or U20938 (N_20938,N_20502,N_20628);
nand U20939 (N_20939,N_20666,N_20531);
nor U20940 (N_20940,N_20599,N_20582);
and U20941 (N_20941,N_20565,N_20574);
nand U20942 (N_20942,N_20547,N_20609);
nand U20943 (N_20943,N_20596,N_20518);
and U20944 (N_20944,N_20602,N_20728);
or U20945 (N_20945,N_20584,N_20587);
nor U20946 (N_20946,N_20596,N_20503);
nand U20947 (N_20947,N_20731,N_20675);
and U20948 (N_20948,N_20623,N_20610);
nand U20949 (N_20949,N_20554,N_20580);
nor U20950 (N_20950,N_20674,N_20591);
and U20951 (N_20951,N_20539,N_20597);
and U20952 (N_20952,N_20572,N_20691);
xnor U20953 (N_20953,N_20639,N_20600);
xnor U20954 (N_20954,N_20617,N_20551);
or U20955 (N_20955,N_20563,N_20682);
nand U20956 (N_20956,N_20723,N_20635);
nand U20957 (N_20957,N_20705,N_20661);
nand U20958 (N_20958,N_20536,N_20714);
and U20959 (N_20959,N_20603,N_20707);
xnor U20960 (N_20960,N_20685,N_20559);
nand U20961 (N_20961,N_20639,N_20653);
and U20962 (N_20962,N_20534,N_20729);
or U20963 (N_20963,N_20593,N_20548);
nand U20964 (N_20964,N_20553,N_20622);
nor U20965 (N_20965,N_20652,N_20659);
nor U20966 (N_20966,N_20502,N_20718);
and U20967 (N_20967,N_20683,N_20716);
nor U20968 (N_20968,N_20711,N_20714);
nand U20969 (N_20969,N_20622,N_20636);
and U20970 (N_20970,N_20596,N_20640);
xor U20971 (N_20971,N_20583,N_20635);
nand U20972 (N_20972,N_20678,N_20629);
nand U20973 (N_20973,N_20694,N_20675);
or U20974 (N_20974,N_20641,N_20631);
and U20975 (N_20975,N_20650,N_20588);
nand U20976 (N_20976,N_20679,N_20505);
or U20977 (N_20977,N_20653,N_20741);
xnor U20978 (N_20978,N_20613,N_20500);
and U20979 (N_20979,N_20510,N_20592);
and U20980 (N_20980,N_20523,N_20738);
and U20981 (N_20981,N_20545,N_20522);
and U20982 (N_20982,N_20537,N_20579);
and U20983 (N_20983,N_20668,N_20519);
or U20984 (N_20984,N_20534,N_20569);
nand U20985 (N_20985,N_20665,N_20643);
nand U20986 (N_20986,N_20535,N_20551);
or U20987 (N_20987,N_20503,N_20704);
nor U20988 (N_20988,N_20613,N_20531);
or U20989 (N_20989,N_20661,N_20531);
nor U20990 (N_20990,N_20502,N_20749);
nand U20991 (N_20991,N_20697,N_20557);
and U20992 (N_20992,N_20537,N_20722);
and U20993 (N_20993,N_20572,N_20643);
or U20994 (N_20994,N_20713,N_20720);
nor U20995 (N_20995,N_20539,N_20715);
xor U20996 (N_20996,N_20749,N_20601);
and U20997 (N_20997,N_20503,N_20599);
and U20998 (N_20998,N_20586,N_20711);
and U20999 (N_20999,N_20615,N_20653);
nand U21000 (N_21000,N_20828,N_20966);
nor U21001 (N_21001,N_20953,N_20803);
nand U21002 (N_21002,N_20792,N_20939);
or U21003 (N_21003,N_20863,N_20936);
and U21004 (N_21004,N_20945,N_20901);
nor U21005 (N_21005,N_20868,N_20820);
nor U21006 (N_21006,N_20970,N_20914);
nand U21007 (N_21007,N_20765,N_20899);
nand U21008 (N_21008,N_20922,N_20844);
nor U21009 (N_21009,N_20769,N_20791);
nand U21010 (N_21010,N_20923,N_20790);
xnor U21011 (N_21011,N_20960,N_20916);
nand U21012 (N_21012,N_20772,N_20834);
nor U21013 (N_21013,N_20987,N_20858);
or U21014 (N_21014,N_20956,N_20823);
and U21015 (N_21015,N_20891,N_20937);
or U21016 (N_21016,N_20979,N_20821);
nor U21017 (N_21017,N_20782,N_20997);
nor U21018 (N_21018,N_20962,N_20940);
nand U21019 (N_21019,N_20985,N_20872);
and U21020 (N_21020,N_20827,N_20885);
xnor U21021 (N_21021,N_20757,N_20959);
nand U21022 (N_21022,N_20919,N_20942);
nand U21023 (N_21023,N_20935,N_20780);
and U21024 (N_21024,N_20944,N_20927);
or U21025 (N_21025,N_20915,N_20992);
nand U21026 (N_21026,N_20795,N_20850);
or U21027 (N_21027,N_20829,N_20907);
and U21028 (N_21028,N_20948,N_20855);
nand U21029 (N_21029,N_20837,N_20952);
and U21030 (N_21030,N_20958,N_20893);
nand U21031 (N_21031,N_20993,N_20892);
or U21032 (N_21032,N_20882,N_20760);
or U21033 (N_21033,N_20943,N_20869);
nor U21034 (N_21034,N_20813,N_20975);
and U21035 (N_21035,N_20900,N_20890);
nand U21036 (N_21036,N_20968,N_20951);
and U21037 (N_21037,N_20920,N_20750);
or U21038 (N_21038,N_20807,N_20859);
or U21039 (N_21039,N_20978,N_20811);
and U21040 (N_21040,N_20866,N_20832);
nand U21041 (N_21041,N_20840,N_20789);
and U21042 (N_21042,N_20822,N_20902);
or U21043 (N_21043,N_20895,N_20836);
nor U21044 (N_21044,N_20818,N_20843);
and U21045 (N_21045,N_20846,N_20949);
nand U21046 (N_21046,N_20857,N_20759);
xor U21047 (N_21047,N_20826,N_20861);
or U21048 (N_21048,N_20982,N_20774);
nor U21049 (N_21049,N_20810,N_20877);
or U21050 (N_21050,N_20842,N_20998);
and U21051 (N_21051,N_20931,N_20947);
xor U21052 (N_21052,N_20785,N_20963);
or U21053 (N_21053,N_20876,N_20875);
or U21054 (N_21054,N_20853,N_20908);
or U21055 (N_21055,N_20996,N_20870);
or U21056 (N_21056,N_20917,N_20903);
and U21057 (N_21057,N_20905,N_20833);
nor U21058 (N_21058,N_20887,N_20897);
and U21059 (N_21059,N_20886,N_20938);
xnor U21060 (N_21060,N_20786,N_20972);
nor U21061 (N_21061,N_20924,N_20809);
nor U21062 (N_21062,N_20812,N_20773);
and U21063 (N_21063,N_20753,N_20961);
nor U21064 (N_21064,N_20969,N_20814);
and U21065 (N_21065,N_20845,N_20880);
and U21066 (N_21066,N_20831,N_20934);
nor U21067 (N_21067,N_20751,N_20994);
nor U21068 (N_21068,N_20838,N_20841);
nand U21069 (N_21069,N_20766,N_20796);
nor U21070 (N_21070,N_20787,N_20763);
or U21071 (N_21071,N_20851,N_20848);
nor U21072 (N_21072,N_20824,N_20889);
or U21073 (N_21073,N_20913,N_20894);
nor U21074 (N_21074,N_20847,N_20925);
nor U21075 (N_21075,N_20898,N_20921);
nand U21076 (N_21076,N_20804,N_20999);
nor U21077 (N_21077,N_20761,N_20865);
and U21078 (N_21078,N_20930,N_20878);
and U21079 (N_21079,N_20867,N_20794);
and U21080 (N_21080,N_20802,N_20941);
or U21081 (N_21081,N_20817,N_20797);
nor U21082 (N_21082,N_20779,N_20758);
and U21083 (N_21083,N_20778,N_20819);
and U21084 (N_21084,N_20946,N_20871);
and U21085 (N_21085,N_20755,N_20860);
nor U21086 (N_21086,N_20783,N_20988);
xor U21087 (N_21087,N_20767,N_20874);
or U21088 (N_21088,N_20967,N_20762);
and U21089 (N_21089,N_20756,N_20775);
or U21090 (N_21090,N_20904,N_20906);
and U21091 (N_21091,N_20801,N_20784);
and U21092 (N_21092,N_20799,N_20825);
nor U21093 (N_21093,N_20918,N_20856);
xnor U21094 (N_21094,N_20768,N_20771);
nor U21095 (N_21095,N_20888,N_20764);
nor U21096 (N_21096,N_20879,N_20781);
nand U21097 (N_21097,N_20933,N_20911);
and U21098 (N_21098,N_20929,N_20770);
nor U21099 (N_21099,N_20950,N_20984);
nand U21100 (N_21100,N_20835,N_20981);
or U21101 (N_21101,N_20881,N_20862);
nand U21102 (N_21102,N_20976,N_20990);
nand U21103 (N_21103,N_20986,N_20816);
and U21104 (N_21104,N_20954,N_20883);
nand U21105 (N_21105,N_20896,N_20989);
nand U21106 (N_21106,N_20912,N_20854);
nor U21107 (N_21107,N_20839,N_20788);
nand U21108 (N_21108,N_20864,N_20973);
nand U21109 (N_21109,N_20777,N_20928);
or U21110 (N_21110,N_20955,N_20991);
xor U21111 (N_21111,N_20957,N_20806);
nor U21112 (N_21112,N_20805,N_20852);
nor U21113 (N_21113,N_20910,N_20815);
xor U21114 (N_21114,N_20926,N_20909);
or U21115 (N_21115,N_20971,N_20980);
nor U21116 (N_21116,N_20776,N_20932);
nand U21117 (N_21117,N_20884,N_20983);
nand U21118 (N_21118,N_20808,N_20830);
and U21119 (N_21119,N_20873,N_20974);
xor U21120 (N_21120,N_20800,N_20977);
and U21121 (N_21121,N_20793,N_20964);
or U21122 (N_21122,N_20965,N_20849);
nor U21123 (N_21123,N_20995,N_20752);
nor U21124 (N_21124,N_20754,N_20798);
xnor U21125 (N_21125,N_20908,N_20989);
xnor U21126 (N_21126,N_20901,N_20782);
nand U21127 (N_21127,N_20906,N_20870);
xnor U21128 (N_21128,N_20771,N_20963);
nor U21129 (N_21129,N_20983,N_20929);
or U21130 (N_21130,N_20987,N_20795);
nor U21131 (N_21131,N_20858,N_20810);
nor U21132 (N_21132,N_20836,N_20786);
and U21133 (N_21133,N_20786,N_20938);
nand U21134 (N_21134,N_20799,N_20998);
and U21135 (N_21135,N_20901,N_20971);
and U21136 (N_21136,N_20882,N_20792);
nor U21137 (N_21137,N_20939,N_20769);
or U21138 (N_21138,N_20851,N_20964);
nor U21139 (N_21139,N_20761,N_20789);
and U21140 (N_21140,N_20864,N_20821);
or U21141 (N_21141,N_20983,N_20998);
and U21142 (N_21142,N_20950,N_20771);
and U21143 (N_21143,N_20937,N_20999);
or U21144 (N_21144,N_20855,N_20754);
nor U21145 (N_21145,N_20830,N_20767);
nand U21146 (N_21146,N_20892,N_20846);
nand U21147 (N_21147,N_20890,N_20881);
and U21148 (N_21148,N_20777,N_20934);
nor U21149 (N_21149,N_20949,N_20936);
nor U21150 (N_21150,N_20974,N_20926);
nor U21151 (N_21151,N_20912,N_20960);
nand U21152 (N_21152,N_20896,N_20836);
nand U21153 (N_21153,N_20888,N_20810);
and U21154 (N_21154,N_20923,N_20844);
and U21155 (N_21155,N_20932,N_20913);
nor U21156 (N_21156,N_20870,N_20833);
nor U21157 (N_21157,N_20860,N_20779);
nand U21158 (N_21158,N_20832,N_20788);
and U21159 (N_21159,N_20882,N_20823);
and U21160 (N_21160,N_20790,N_20755);
xnor U21161 (N_21161,N_20891,N_20777);
xor U21162 (N_21162,N_20968,N_20905);
nand U21163 (N_21163,N_20965,N_20912);
or U21164 (N_21164,N_20938,N_20940);
nand U21165 (N_21165,N_20945,N_20843);
or U21166 (N_21166,N_20813,N_20880);
or U21167 (N_21167,N_20854,N_20902);
nor U21168 (N_21168,N_20876,N_20989);
nand U21169 (N_21169,N_20778,N_20979);
nor U21170 (N_21170,N_20819,N_20868);
nor U21171 (N_21171,N_20944,N_20929);
nand U21172 (N_21172,N_20964,N_20879);
nand U21173 (N_21173,N_20890,N_20924);
and U21174 (N_21174,N_20851,N_20825);
nor U21175 (N_21175,N_20860,N_20865);
or U21176 (N_21176,N_20939,N_20979);
and U21177 (N_21177,N_20902,N_20928);
or U21178 (N_21178,N_20982,N_20787);
nor U21179 (N_21179,N_20760,N_20821);
nand U21180 (N_21180,N_20935,N_20953);
nor U21181 (N_21181,N_20915,N_20943);
nand U21182 (N_21182,N_20805,N_20821);
and U21183 (N_21183,N_20760,N_20931);
nor U21184 (N_21184,N_20871,N_20920);
or U21185 (N_21185,N_20927,N_20991);
nand U21186 (N_21186,N_20904,N_20889);
and U21187 (N_21187,N_20836,N_20977);
nand U21188 (N_21188,N_20830,N_20858);
xnor U21189 (N_21189,N_20882,N_20811);
or U21190 (N_21190,N_20884,N_20828);
or U21191 (N_21191,N_20879,N_20939);
nor U21192 (N_21192,N_20961,N_20882);
nand U21193 (N_21193,N_20983,N_20773);
and U21194 (N_21194,N_20910,N_20907);
or U21195 (N_21195,N_20992,N_20847);
or U21196 (N_21196,N_20985,N_20808);
xnor U21197 (N_21197,N_20852,N_20810);
nand U21198 (N_21198,N_20778,N_20821);
nand U21199 (N_21199,N_20904,N_20854);
nor U21200 (N_21200,N_20975,N_20860);
xor U21201 (N_21201,N_20817,N_20941);
and U21202 (N_21202,N_20963,N_20788);
nand U21203 (N_21203,N_20911,N_20803);
and U21204 (N_21204,N_20897,N_20935);
nor U21205 (N_21205,N_20756,N_20924);
nand U21206 (N_21206,N_20908,N_20828);
or U21207 (N_21207,N_20754,N_20933);
nor U21208 (N_21208,N_20769,N_20852);
nor U21209 (N_21209,N_20929,N_20788);
nand U21210 (N_21210,N_20774,N_20873);
nand U21211 (N_21211,N_20868,N_20871);
and U21212 (N_21212,N_20900,N_20859);
or U21213 (N_21213,N_20963,N_20799);
or U21214 (N_21214,N_20751,N_20764);
or U21215 (N_21215,N_20862,N_20782);
or U21216 (N_21216,N_20949,N_20873);
and U21217 (N_21217,N_20750,N_20835);
nor U21218 (N_21218,N_20906,N_20829);
and U21219 (N_21219,N_20781,N_20927);
or U21220 (N_21220,N_20951,N_20898);
nor U21221 (N_21221,N_20903,N_20848);
nor U21222 (N_21222,N_20975,N_20942);
nor U21223 (N_21223,N_20866,N_20884);
nor U21224 (N_21224,N_20928,N_20954);
or U21225 (N_21225,N_20789,N_20872);
nor U21226 (N_21226,N_20973,N_20877);
or U21227 (N_21227,N_20867,N_20832);
nand U21228 (N_21228,N_20955,N_20894);
nand U21229 (N_21229,N_20976,N_20833);
nor U21230 (N_21230,N_20836,N_20762);
and U21231 (N_21231,N_20827,N_20853);
or U21232 (N_21232,N_20817,N_20762);
xnor U21233 (N_21233,N_20977,N_20906);
nand U21234 (N_21234,N_20979,N_20830);
xor U21235 (N_21235,N_20916,N_20995);
or U21236 (N_21236,N_20869,N_20832);
nor U21237 (N_21237,N_20956,N_20991);
nor U21238 (N_21238,N_20965,N_20776);
or U21239 (N_21239,N_20783,N_20895);
or U21240 (N_21240,N_20797,N_20770);
xnor U21241 (N_21241,N_20975,N_20764);
nand U21242 (N_21242,N_20800,N_20765);
nand U21243 (N_21243,N_20980,N_20823);
and U21244 (N_21244,N_20904,N_20771);
and U21245 (N_21245,N_20828,N_20859);
and U21246 (N_21246,N_20782,N_20859);
xor U21247 (N_21247,N_20905,N_20810);
nor U21248 (N_21248,N_20792,N_20925);
nor U21249 (N_21249,N_20976,N_20764);
nand U21250 (N_21250,N_21187,N_21084);
and U21251 (N_21251,N_21088,N_21140);
nor U21252 (N_21252,N_21011,N_21208);
or U21253 (N_21253,N_21128,N_21051);
or U21254 (N_21254,N_21061,N_21171);
or U21255 (N_21255,N_21151,N_21113);
nand U21256 (N_21256,N_21137,N_21127);
xor U21257 (N_21257,N_21062,N_21207);
nor U21258 (N_21258,N_21203,N_21010);
or U21259 (N_21259,N_21042,N_21013);
nand U21260 (N_21260,N_21068,N_21043);
and U21261 (N_21261,N_21135,N_21122);
nand U21262 (N_21262,N_21035,N_21060);
and U21263 (N_21263,N_21094,N_21149);
nor U21264 (N_21264,N_21235,N_21064);
xor U21265 (N_21265,N_21097,N_21161);
xnor U21266 (N_21266,N_21226,N_21000);
nand U21267 (N_21267,N_21195,N_21220);
and U21268 (N_21268,N_21031,N_21157);
or U21269 (N_21269,N_21102,N_21192);
or U21270 (N_21270,N_21019,N_21188);
nor U21271 (N_21271,N_21210,N_21212);
nor U21272 (N_21272,N_21152,N_21052);
nor U21273 (N_21273,N_21156,N_21003);
and U21274 (N_21274,N_21050,N_21092);
nor U21275 (N_21275,N_21083,N_21246);
xor U21276 (N_21276,N_21146,N_21144);
or U21277 (N_21277,N_21100,N_21016);
and U21278 (N_21278,N_21045,N_21225);
and U21279 (N_21279,N_21026,N_21181);
or U21280 (N_21280,N_21160,N_21008);
xor U21281 (N_21281,N_21239,N_21240);
nor U21282 (N_21282,N_21227,N_21023);
nand U21283 (N_21283,N_21070,N_21086);
and U21284 (N_21284,N_21184,N_21096);
xor U21285 (N_21285,N_21036,N_21107);
and U21286 (N_21286,N_21038,N_21154);
nand U21287 (N_21287,N_21054,N_21124);
xnor U21288 (N_21288,N_21034,N_21230);
or U21289 (N_21289,N_21029,N_21028);
nand U21290 (N_21290,N_21224,N_21180);
nand U21291 (N_21291,N_21001,N_21002);
nand U21292 (N_21292,N_21056,N_21053);
nor U21293 (N_21293,N_21039,N_21098);
nor U21294 (N_21294,N_21211,N_21205);
nor U21295 (N_21295,N_21093,N_21147);
nand U21296 (N_21296,N_21085,N_21164);
nor U21297 (N_21297,N_21020,N_21167);
or U21298 (N_21298,N_21072,N_21223);
nor U21299 (N_21299,N_21080,N_21063);
or U21300 (N_21300,N_21229,N_21216);
or U21301 (N_21301,N_21129,N_21006);
nand U21302 (N_21302,N_21197,N_21118);
or U21303 (N_21303,N_21109,N_21130);
nand U21304 (N_21304,N_21081,N_21055);
and U21305 (N_21305,N_21091,N_21131);
nor U21306 (N_21306,N_21231,N_21159);
nor U21307 (N_21307,N_21133,N_21241);
or U21308 (N_21308,N_21243,N_21047);
and U21309 (N_21309,N_21079,N_21082);
nor U21310 (N_21310,N_21136,N_21125);
nand U21311 (N_21311,N_21204,N_21110);
or U21312 (N_21312,N_21044,N_21027);
or U21313 (N_21313,N_21066,N_21142);
or U21314 (N_21314,N_21190,N_21065);
and U21315 (N_21315,N_21089,N_21170);
and U21316 (N_21316,N_21025,N_21134);
nor U21317 (N_21317,N_21057,N_21214);
or U21318 (N_21318,N_21015,N_21067);
nor U21319 (N_21319,N_21032,N_21219);
or U21320 (N_21320,N_21169,N_21059);
or U21321 (N_21321,N_21155,N_21014);
or U21322 (N_21322,N_21114,N_21221);
xnor U21323 (N_21323,N_21087,N_21004);
or U21324 (N_21324,N_21215,N_21162);
nor U21325 (N_21325,N_21049,N_21017);
nand U21326 (N_21326,N_21007,N_21021);
nor U21327 (N_21327,N_21126,N_21116);
xor U21328 (N_21328,N_21244,N_21105);
nor U21329 (N_21329,N_21117,N_21012);
or U21330 (N_21330,N_21168,N_21236);
xnor U21331 (N_21331,N_21058,N_21234);
nand U21332 (N_21332,N_21148,N_21106);
or U21333 (N_21333,N_21075,N_21018);
or U21334 (N_21334,N_21121,N_21248);
nand U21335 (N_21335,N_21217,N_21233);
xor U21336 (N_21336,N_21249,N_21175);
nand U21337 (N_21337,N_21022,N_21206);
nor U21338 (N_21338,N_21048,N_21153);
and U21339 (N_21339,N_21009,N_21090);
nor U21340 (N_21340,N_21196,N_21099);
or U21341 (N_21341,N_21041,N_21218);
nand U21342 (N_21342,N_21119,N_21037);
nand U21343 (N_21343,N_21115,N_21076);
nor U21344 (N_21344,N_21199,N_21242);
or U21345 (N_21345,N_21139,N_21201);
nand U21346 (N_21346,N_21166,N_21120);
nand U21347 (N_21347,N_21183,N_21237);
nand U21348 (N_21348,N_21158,N_21173);
nor U21349 (N_21349,N_21222,N_21172);
nor U21350 (N_21350,N_21200,N_21030);
and U21351 (N_21351,N_21194,N_21005);
nor U21352 (N_21352,N_21185,N_21245);
or U21353 (N_21353,N_21141,N_21189);
nor U21354 (N_21354,N_21143,N_21179);
nand U21355 (N_21355,N_21108,N_21178);
and U21356 (N_21356,N_21071,N_21074);
nor U21357 (N_21357,N_21123,N_21138);
nor U21358 (N_21358,N_21073,N_21198);
nor U21359 (N_21359,N_21213,N_21104);
and U21360 (N_21360,N_21077,N_21112);
and U21361 (N_21361,N_21191,N_21238);
nand U21362 (N_21362,N_21046,N_21033);
or U21363 (N_21363,N_21145,N_21228);
and U21364 (N_21364,N_21101,N_21202);
and U21365 (N_21365,N_21132,N_21024);
nand U21366 (N_21366,N_21111,N_21177);
nor U21367 (N_21367,N_21232,N_21150);
or U21368 (N_21368,N_21069,N_21095);
nand U21369 (N_21369,N_21247,N_21209);
nor U21370 (N_21370,N_21186,N_21176);
nand U21371 (N_21371,N_21163,N_21103);
nand U21372 (N_21372,N_21174,N_21193);
nand U21373 (N_21373,N_21078,N_21182);
or U21374 (N_21374,N_21040,N_21165);
nor U21375 (N_21375,N_21217,N_21062);
or U21376 (N_21376,N_21242,N_21103);
nand U21377 (N_21377,N_21012,N_21094);
or U21378 (N_21378,N_21129,N_21090);
and U21379 (N_21379,N_21048,N_21044);
nand U21380 (N_21380,N_21154,N_21108);
nor U21381 (N_21381,N_21241,N_21199);
xnor U21382 (N_21382,N_21094,N_21225);
or U21383 (N_21383,N_21170,N_21102);
or U21384 (N_21384,N_21117,N_21064);
nor U21385 (N_21385,N_21219,N_21244);
xnor U21386 (N_21386,N_21119,N_21202);
nand U21387 (N_21387,N_21028,N_21087);
or U21388 (N_21388,N_21172,N_21247);
nor U21389 (N_21389,N_21197,N_21110);
nand U21390 (N_21390,N_21013,N_21079);
nor U21391 (N_21391,N_21140,N_21189);
or U21392 (N_21392,N_21022,N_21246);
and U21393 (N_21393,N_21050,N_21134);
or U21394 (N_21394,N_21243,N_21073);
nor U21395 (N_21395,N_21027,N_21207);
and U21396 (N_21396,N_21244,N_21163);
nor U21397 (N_21397,N_21114,N_21073);
and U21398 (N_21398,N_21009,N_21199);
nand U21399 (N_21399,N_21035,N_21019);
and U21400 (N_21400,N_21246,N_21076);
nand U21401 (N_21401,N_21168,N_21048);
nand U21402 (N_21402,N_21079,N_21213);
and U21403 (N_21403,N_21217,N_21065);
and U21404 (N_21404,N_21043,N_21237);
or U21405 (N_21405,N_21056,N_21002);
xnor U21406 (N_21406,N_21098,N_21087);
and U21407 (N_21407,N_21007,N_21110);
nand U21408 (N_21408,N_21150,N_21196);
and U21409 (N_21409,N_21124,N_21065);
nand U21410 (N_21410,N_21227,N_21116);
nor U21411 (N_21411,N_21043,N_21062);
or U21412 (N_21412,N_21160,N_21015);
and U21413 (N_21413,N_21102,N_21186);
nor U21414 (N_21414,N_21146,N_21243);
and U21415 (N_21415,N_21139,N_21103);
or U21416 (N_21416,N_21198,N_21221);
or U21417 (N_21417,N_21009,N_21140);
nor U21418 (N_21418,N_21018,N_21249);
and U21419 (N_21419,N_21110,N_21234);
xor U21420 (N_21420,N_21145,N_21235);
xnor U21421 (N_21421,N_21151,N_21023);
nor U21422 (N_21422,N_21079,N_21062);
or U21423 (N_21423,N_21099,N_21117);
xnor U21424 (N_21424,N_21215,N_21184);
nand U21425 (N_21425,N_21227,N_21019);
or U21426 (N_21426,N_21177,N_21162);
and U21427 (N_21427,N_21145,N_21008);
nor U21428 (N_21428,N_21003,N_21096);
and U21429 (N_21429,N_21133,N_21230);
and U21430 (N_21430,N_21092,N_21122);
nand U21431 (N_21431,N_21017,N_21144);
nor U21432 (N_21432,N_21143,N_21215);
or U21433 (N_21433,N_21222,N_21185);
xor U21434 (N_21434,N_21246,N_21066);
nor U21435 (N_21435,N_21191,N_21135);
nand U21436 (N_21436,N_21152,N_21142);
and U21437 (N_21437,N_21095,N_21233);
or U21438 (N_21438,N_21180,N_21203);
or U21439 (N_21439,N_21245,N_21237);
and U21440 (N_21440,N_21209,N_21218);
nor U21441 (N_21441,N_21080,N_21235);
and U21442 (N_21442,N_21247,N_21135);
or U21443 (N_21443,N_21014,N_21109);
or U21444 (N_21444,N_21046,N_21113);
nor U21445 (N_21445,N_21175,N_21087);
or U21446 (N_21446,N_21127,N_21171);
and U21447 (N_21447,N_21003,N_21221);
or U21448 (N_21448,N_21221,N_21082);
or U21449 (N_21449,N_21056,N_21075);
and U21450 (N_21450,N_21002,N_21222);
or U21451 (N_21451,N_21108,N_21064);
nand U21452 (N_21452,N_21233,N_21000);
nand U21453 (N_21453,N_21089,N_21025);
nor U21454 (N_21454,N_21079,N_21163);
and U21455 (N_21455,N_21199,N_21224);
xnor U21456 (N_21456,N_21053,N_21243);
and U21457 (N_21457,N_21116,N_21028);
xnor U21458 (N_21458,N_21179,N_21121);
or U21459 (N_21459,N_21060,N_21033);
or U21460 (N_21460,N_21156,N_21199);
and U21461 (N_21461,N_21101,N_21179);
or U21462 (N_21462,N_21142,N_21245);
and U21463 (N_21463,N_21242,N_21145);
or U21464 (N_21464,N_21156,N_21150);
nand U21465 (N_21465,N_21206,N_21048);
nor U21466 (N_21466,N_21064,N_21129);
and U21467 (N_21467,N_21231,N_21143);
nand U21468 (N_21468,N_21235,N_21020);
and U21469 (N_21469,N_21153,N_21064);
or U21470 (N_21470,N_21006,N_21166);
and U21471 (N_21471,N_21145,N_21132);
nand U21472 (N_21472,N_21213,N_21169);
nand U21473 (N_21473,N_21022,N_21228);
xor U21474 (N_21474,N_21219,N_21236);
or U21475 (N_21475,N_21061,N_21165);
nor U21476 (N_21476,N_21137,N_21181);
and U21477 (N_21477,N_21013,N_21063);
or U21478 (N_21478,N_21058,N_21018);
nor U21479 (N_21479,N_21158,N_21199);
nor U21480 (N_21480,N_21102,N_21132);
nor U21481 (N_21481,N_21116,N_21095);
xor U21482 (N_21482,N_21135,N_21099);
nand U21483 (N_21483,N_21137,N_21059);
nor U21484 (N_21484,N_21093,N_21136);
nor U21485 (N_21485,N_21063,N_21153);
nor U21486 (N_21486,N_21231,N_21084);
nand U21487 (N_21487,N_21227,N_21089);
xor U21488 (N_21488,N_21116,N_21173);
and U21489 (N_21489,N_21176,N_21021);
nor U21490 (N_21490,N_21032,N_21200);
xor U21491 (N_21491,N_21196,N_21111);
and U21492 (N_21492,N_21050,N_21201);
nor U21493 (N_21493,N_21149,N_21189);
nor U21494 (N_21494,N_21025,N_21182);
xnor U21495 (N_21495,N_21041,N_21045);
and U21496 (N_21496,N_21229,N_21133);
nand U21497 (N_21497,N_21134,N_21243);
and U21498 (N_21498,N_21211,N_21128);
or U21499 (N_21499,N_21214,N_21026);
or U21500 (N_21500,N_21363,N_21470);
nand U21501 (N_21501,N_21498,N_21274);
xnor U21502 (N_21502,N_21250,N_21359);
or U21503 (N_21503,N_21352,N_21454);
or U21504 (N_21504,N_21407,N_21329);
xnor U21505 (N_21505,N_21287,N_21305);
nor U21506 (N_21506,N_21499,N_21429);
and U21507 (N_21507,N_21448,N_21330);
and U21508 (N_21508,N_21477,N_21424);
nand U21509 (N_21509,N_21387,N_21426);
and U21510 (N_21510,N_21441,N_21260);
or U21511 (N_21511,N_21483,N_21374);
and U21512 (N_21512,N_21464,N_21345);
xnor U21513 (N_21513,N_21447,N_21372);
nand U21514 (N_21514,N_21295,N_21421);
and U21515 (N_21515,N_21254,N_21405);
nand U21516 (N_21516,N_21416,N_21268);
nand U21517 (N_21517,N_21257,N_21453);
xor U21518 (N_21518,N_21388,N_21435);
nor U21519 (N_21519,N_21475,N_21315);
and U21520 (N_21520,N_21450,N_21458);
nand U21521 (N_21521,N_21273,N_21456);
nand U21522 (N_21522,N_21382,N_21288);
xnor U21523 (N_21523,N_21313,N_21482);
nor U21524 (N_21524,N_21495,N_21394);
or U21525 (N_21525,N_21439,N_21338);
and U21526 (N_21526,N_21466,N_21402);
and U21527 (N_21527,N_21357,N_21266);
and U21528 (N_21528,N_21370,N_21391);
xnor U21529 (N_21529,N_21479,N_21281);
nor U21530 (N_21530,N_21320,N_21304);
and U21531 (N_21531,N_21444,N_21472);
nand U21532 (N_21532,N_21377,N_21280);
xnor U21533 (N_21533,N_21327,N_21425);
or U21534 (N_21534,N_21310,N_21368);
and U21535 (N_21535,N_21417,N_21346);
or U21536 (N_21536,N_21399,N_21414);
nor U21537 (N_21537,N_21271,N_21440);
nor U21538 (N_21538,N_21361,N_21390);
nor U21539 (N_21539,N_21321,N_21264);
nor U21540 (N_21540,N_21471,N_21270);
xnor U21541 (N_21541,N_21344,N_21339);
nand U21542 (N_21542,N_21303,N_21398);
nor U21543 (N_21543,N_21400,N_21443);
nand U21544 (N_21544,N_21319,N_21316);
and U21545 (N_21545,N_21384,N_21393);
and U21546 (N_21546,N_21297,N_21465);
nor U21547 (N_21547,N_21301,N_21350);
or U21548 (N_21548,N_21341,N_21434);
xnor U21549 (N_21549,N_21348,N_21497);
and U21550 (N_21550,N_21252,N_21331);
xnor U21551 (N_21551,N_21298,N_21251);
or U21552 (N_21552,N_21397,N_21317);
nor U21553 (N_21553,N_21311,N_21360);
or U21554 (N_21554,N_21406,N_21463);
and U21555 (N_21555,N_21415,N_21476);
and U21556 (N_21556,N_21267,N_21496);
nor U21557 (N_21557,N_21309,N_21326);
nand U21558 (N_21558,N_21437,N_21409);
nand U21559 (N_21559,N_21473,N_21299);
and U21560 (N_21560,N_21308,N_21282);
nand U21561 (N_21561,N_21375,N_21389);
nor U21562 (N_21562,N_21428,N_21446);
and U21563 (N_21563,N_21334,N_21486);
nor U21564 (N_21564,N_21460,N_21478);
and U21565 (N_21565,N_21379,N_21380);
xnor U21566 (N_21566,N_21291,N_21278);
and U21567 (N_21567,N_21449,N_21353);
or U21568 (N_21568,N_21276,N_21365);
nand U21569 (N_21569,N_21294,N_21392);
and U21570 (N_21570,N_21355,N_21459);
nor U21571 (N_21571,N_21277,N_21481);
nor U21572 (N_21572,N_21488,N_21369);
and U21573 (N_21573,N_21494,N_21323);
nor U21574 (N_21574,N_21457,N_21351);
and U21575 (N_21575,N_21306,N_21354);
nand U21576 (N_21576,N_21296,N_21364);
nor U21577 (N_21577,N_21358,N_21445);
xnor U21578 (N_21578,N_21436,N_21283);
nand U21579 (N_21579,N_21340,N_21462);
nor U21580 (N_21580,N_21403,N_21401);
or U21581 (N_21581,N_21427,N_21376);
or U21582 (N_21582,N_21461,N_21279);
nand U21583 (N_21583,N_21259,N_21256);
or U21584 (N_21584,N_21493,N_21312);
nand U21585 (N_21585,N_21333,N_21255);
and U21586 (N_21586,N_21442,N_21289);
or U21587 (N_21587,N_21302,N_21285);
or U21588 (N_21588,N_21335,N_21366);
or U21589 (N_21589,N_21284,N_21385);
nor U21590 (N_21590,N_21336,N_21485);
or U21591 (N_21591,N_21325,N_21419);
nand U21592 (N_21592,N_21432,N_21418);
nor U21593 (N_21593,N_21293,N_21300);
nand U21594 (N_21594,N_21318,N_21420);
and U21595 (N_21595,N_21322,N_21314);
or U21596 (N_21596,N_21337,N_21342);
xnor U21597 (N_21597,N_21286,N_21491);
nand U21598 (N_21598,N_21343,N_21253);
nor U21599 (N_21599,N_21262,N_21469);
or U21600 (N_21600,N_21258,N_21396);
nand U21601 (N_21601,N_21349,N_21452);
or U21602 (N_21602,N_21272,N_21408);
xor U21603 (N_21603,N_21433,N_21324);
or U21604 (N_21604,N_21468,N_21484);
nor U21605 (N_21605,N_21307,N_21378);
or U21606 (N_21606,N_21381,N_21474);
nand U21607 (N_21607,N_21404,N_21290);
and U21608 (N_21608,N_21367,N_21490);
and U21609 (N_21609,N_21269,N_21328);
nor U21610 (N_21610,N_21412,N_21410);
xnor U21611 (N_21611,N_21430,N_21362);
xnor U21612 (N_21612,N_21383,N_21487);
and U21613 (N_21613,N_21356,N_21423);
nand U21614 (N_21614,N_21413,N_21347);
nand U21615 (N_21615,N_21492,N_21480);
nand U21616 (N_21616,N_21455,N_21373);
nor U21617 (N_21617,N_21411,N_21489);
nor U21618 (N_21618,N_21451,N_21467);
and U21619 (N_21619,N_21292,N_21261);
and U21620 (N_21620,N_21371,N_21438);
or U21621 (N_21621,N_21275,N_21422);
nor U21622 (N_21622,N_21263,N_21386);
nand U21623 (N_21623,N_21265,N_21332);
xnor U21624 (N_21624,N_21395,N_21431);
and U21625 (N_21625,N_21376,N_21406);
nor U21626 (N_21626,N_21434,N_21481);
nor U21627 (N_21627,N_21493,N_21422);
or U21628 (N_21628,N_21290,N_21258);
nand U21629 (N_21629,N_21345,N_21393);
nand U21630 (N_21630,N_21406,N_21392);
nor U21631 (N_21631,N_21486,N_21315);
nand U21632 (N_21632,N_21337,N_21254);
and U21633 (N_21633,N_21352,N_21496);
and U21634 (N_21634,N_21492,N_21307);
and U21635 (N_21635,N_21487,N_21287);
or U21636 (N_21636,N_21432,N_21328);
and U21637 (N_21637,N_21443,N_21477);
nand U21638 (N_21638,N_21350,N_21277);
and U21639 (N_21639,N_21423,N_21278);
and U21640 (N_21640,N_21297,N_21253);
or U21641 (N_21641,N_21410,N_21484);
and U21642 (N_21642,N_21480,N_21455);
nor U21643 (N_21643,N_21404,N_21354);
nor U21644 (N_21644,N_21267,N_21292);
nor U21645 (N_21645,N_21273,N_21332);
xor U21646 (N_21646,N_21282,N_21437);
nor U21647 (N_21647,N_21345,N_21447);
or U21648 (N_21648,N_21376,N_21441);
nor U21649 (N_21649,N_21252,N_21312);
and U21650 (N_21650,N_21284,N_21478);
or U21651 (N_21651,N_21340,N_21291);
nor U21652 (N_21652,N_21453,N_21268);
or U21653 (N_21653,N_21448,N_21476);
or U21654 (N_21654,N_21475,N_21387);
and U21655 (N_21655,N_21475,N_21402);
xor U21656 (N_21656,N_21362,N_21306);
or U21657 (N_21657,N_21385,N_21437);
or U21658 (N_21658,N_21307,N_21410);
nor U21659 (N_21659,N_21257,N_21365);
or U21660 (N_21660,N_21373,N_21274);
or U21661 (N_21661,N_21256,N_21305);
nor U21662 (N_21662,N_21326,N_21320);
nor U21663 (N_21663,N_21281,N_21407);
or U21664 (N_21664,N_21310,N_21349);
nor U21665 (N_21665,N_21273,N_21253);
or U21666 (N_21666,N_21395,N_21375);
or U21667 (N_21667,N_21282,N_21396);
and U21668 (N_21668,N_21251,N_21440);
or U21669 (N_21669,N_21476,N_21485);
nand U21670 (N_21670,N_21382,N_21380);
xnor U21671 (N_21671,N_21308,N_21498);
nor U21672 (N_21672,N_21268,N_21251);
nand U21673 (N_21673,N_21315,N_21360);
nor U21674 (N_21674,N_21321,N_21285);
and U21675 (N_21675,N_21275,N_21376);
or U21676 (N_21676,N_21449,N_21468);
nand U21677 (N_21677,N_21276,N_21297);
nand U21678 (N_21678,N_21426,N_21458);
or U21679 (N_21679,N_21441,N_21290);
xnor U21680 (N_21680,N_21332,N_21381);
nand U21681 (N_21681,N_21309,N_21306);
and U21682 (N_21682,N_21449,N_21459);
and U21683 (N_21683,N_21311,N_21363);
nor U21684 (N_21684,N_21490,N_21422);
or U21685 (N_21685,N_21343,N_21446);
nand U21686 (N_21686,N_21330,N_21353);
or U21687 (N_21687,N_21446,N_21377);
or U21688 (N_21688,N_21308,N_21261);
or U21689 (N_21689,N_21287,N_21364);
xnor U21690 (N_21690,N_21462,N_21285);
or U21691 (N_21691,N_21330,N_21472);
nand U21692 (N_21692,N_21394,N_21473);
nor U21693 (N_21693,N_21386,N_21309);
nand U21694 (N_21694,N_21486,N_21320);
or U21695 (N_21695,N_21403,N_21354);
nand U21696 (N_21696,N_21283,N_21425);
nor U21697 (N_21697,N_21428,N_21354);
nor U21698 (N_21698,N_21409,N_21360);
xnor U21699 (N_21699,N_21478,N_21453);
nand U21700 (N_21700,N_21267,N_21439);
or U21701 (N_21701,N_21281,N_21341);
and U21702 (N_21702,N_21343,N_21260);
nor U21703 (N_21703,N_21368,N_21422);
nor U21704 (N_21704,N_21377,N_21491);
and U21705 (N_21705,N_21346,N_21478);
nand U21706 (N_21706,N_21278,N_21396);
nand U21707 (N_21707,N_21405,N_21308);
nand U21708 (N_21708,N_21384,N_21371);
nor U21709 (N_21709,N_21302,N_21348);
nand U21710 (N_21710,N_21333,N_21461);
nor U21711 (N_21711,N_21259,N_21273);
nor U21712 (N_21712,N_21282,N_21258);
and U21713 (N_21713,N_21271,N_21495);
and U21714 (N_21714,N_21471,N_21408);
nand U21715 (N_21715,N_21475,N_21294);
nand U21716 (N_21716,N_21403,N_21418);
nor U21717 (N_21717,N_21447,N_21279);
nor U21718 (N_21718,N_21498,N_21448);
or U21719 (N_21719,N_21331,N_21290);
nor U21720 (N_21720,N_21390,N_21256);
nor U21721 (N_21721,N_21387,N_21296);
nand U21722 (N_21722,N_21312,N_21303);
nor U21723 (N_21723,N_21409,N_21264);
nand U21724 (N_21724,N_21386,N_21294);
nand U21725 (N_21725,N_21336,N_21369);
nand U21726 (N_21726,N_21494,N_21358);
nand U21727 (N_21727,N_21301,N_21308);
nand U21728 (N_21728,N_21338,N_21370);
nand U21729 (N_21729,N_21311,N_21272);
nand U21730 (N_21730,N_21317,N_21361);
nand U21731 (N_21731,N_21352,N_21423);
or U21732 (N_21732,N_21278,N_21407);
nor U21733 (N_21733,N_21459,N_21352);
nand U21734 (N_21734,N_21374,N_21269);
or U21735 (N_21735,N_21287,N_21296);
and U21736 (N_21736,N_21280,N_21365);
nor U21737 (N_21737,N_21292,N_21456);
and U21738 (N_21738,N_21268,N_21364);
nand U21739 (N_21739,N_21457,N_21365);
or U21740 (N_21740,N_21411,N_21478);
nor U21741 (N_21741,N_21359,N_21395);
or U21742 (N_21742,N_21259,N_21318);
xor U21743 (N_21743,N_21490,N_21458);
xor U21744 (N_21744,N_21322,N_21369);
nor U21745 (N_21745,N_21363,N_21303);
and U21746 (N_21746,N_21352,N_21493);
or U21747 (N_21747,N_21251,N_21392);
nor U21748 (N_21748,N_21462,N_21479);
xor U21749 (N_21749,N_21454,N_21467);
nand U21750 (N_21750,N_21534,N_21657);
nand U21751 (N_21751,N_21553,N_21623);
or U21752 (N_21752,N_21702,N_21564);
xor U21753 (N_21753,N_21630,N_21629);
or U21754 (N_21754,N_21527,N_21699);
xor U21755 (N_21755,N_21594,N_21710);
and U21756 (N_21756,N_21730,N_21679);
nand U21757 (N_21757,N_21646,N_21524);
or U21758 (N_21758,N_21715,N_21732);
nand U21759 (N_21759,N_21525,N_21705);
nor U21760 (N_21760,N_21691,N_21675);
nand U21761 (N_21761,N_21543,N_21516);
nor U21762 (N_21762,N_21625,N_21743);
nand U21763 (N_21763,N_21648,N_21502);
nand U21764 (N_21764,N_21568,N_21592);
nand U21765 (N_21765,N_21550,N_21503);
nand U21766 (N_21766,N_21624,N_21749);
nor U21767 (N_21767,N_21717,N_21682);
nor U21768 (N_21768,N_21612,N_21662);
nand U21769 (N_21769,N_21703,N_21532);
nor U21770 (N_21770,N_21554,N_21620);
or U21771 (N_21771,N_21667,N_21688);
or U21772 (N_21772,N_21570,N_21601);
nand U21773 (N_21773,N_21610,N_21513);
xor U21774 (N_21774,N_21747,N_21638);
nand U21775 (N_21775,N_21724,N_21668);
xnor U21776 (N_21776,N_21511,N_21678);
xor U21777 (N_21777,N_21714,N_21509);
and U21778 (N_21778,N_21510,N_21693);
nand U21779 (N_21779,N_21653,N_21671);
nand U21780 (N_21780,N_21697,N_21566);
or U21781 (N_21781,N_21613,N_21698);
nor U21782 (N_21782,N_21636,N_21522);
nor U21783 (N_21783,N_21549,N_21645);
or U21784 (N_21784,N_21582,N_21631);
or U21785 (N_21785,N_21606,N_21716);
nor U21786 (N_21786,N_21512,N_21571);
nor U21787 (N_21787,N_21580,N_21692);
or U21788 (N_21788,N_21655,N_21713);
nor U21789 (N_21789,N_21587,N_21731);
nand U21790 (N_21790,N_21514,N_21595);
nor U21791 (N_21791,N_21650,N_21628);
and U21792 (N_21792,N_21721,N_21530);
nand U21793 (N_21793,N_21538,N_21683);
nor U21794 (N_21794,N_21643,N_21729);
nand U21795 (N_21795,N_21515,N_21674);
or U21796 (N_21796,N_21575,N_21621);
and U21797 (N_21797,N_21569,N_21586);
and U21798 (N_21798,N_21540,N_21618);
and U21799 (N_21799,N_21720,N_21644);
nor U21800 (N_21800,N_21508,N_21607);
or U21801 (N_21801,N_21573,N_21526);
and U21802 (N_21802,N_21589,N_21633);
nor U21803 (N_21803,N_21739,N_21632);
nand U21804 (N_21804,N_21658,N_21647);
and U21805 (N_21805,N_21560,N_21727);
xnor U21806 (N_21806,N_21615,N_21725);
and U21807 (N_21807,N_21616,N_21637);
or U21808 (N_21808,N_21562,N_21673);
and U21809 (N_21809,N_21583,N_21742);
or U21810 (N_21810,N_21689,N_21617);
nand U21811 (N_21811,N_21622,N_21608);
or U21812 (N_21812,N_21572,N_21519);
nand U21813 (N_21813,N_21701,N_21561);
and U21814 (N_21814,N_21545,N_21709);
nand U21815 (N_21815,N_21627,N_21591);
or U21816 (N_21816,N_21507,N_21558);
xor U21817 (N_21817,N_21556,N_21733);
or U21818 (N_21818,N_21664,N_21563);
and U21819 (N_21819,N_21711,N_21734);
nor U21820 (N_21820,N_21619,N_21719);
or U21821 (N_21821,N_21567,N_21659);
or U21822 (N_21822,N_21676,N_21661);
nor U21823 (N_21823,N_21736,N_21665);
nor U21824 (N_21824,N_21600,N_21728);
nor U21825 (N_21825,N_21609,N_21686);
and U21826 (N_21826,N_21555,N_21700);
or U21827 (N_21827,N_21536,N_21578);
nor U21828 (N_21828,N_21718,N_21597);
and U21829 (N_21829,N_21640,N_21504);
or U21830 (N_21830,N_21544,N_21741);
or U21831 (N_21831,N_21611,N_21529);
or U21832 (N_21832,N_21744,N_21641);
nor U21833 (N_21833,N_21656,N_21639);
or U21834 (N_21834,N_21680,N_21635);
nor U21835 (N_21835,N_21574,N_21581);
nand U21836 (N_21836,N_21501,N_21523);
nand U21837 (N_21837,N_21694,N_21726);
or U21838 (N_21838,N_21669,N_21672);
or U21839 (N_21839,N_21559,N_21542);
xor U21840 (N_21840,N_21548,N_21602);
xor U21841 (N_21841,N_21634,N_21712);
or U21842 (N_21842,N_21642,N_21685);
and U21843 (N_21843,N_21537,N_21654);
nor U21844 (N_21844,N_21681,N_21593);
nor U21845 (N_21845,N_21552,N_21738);
xor U21846 (N_21846,N_21596,N_21500);
xnor U21847 (N_21847,N_21565,N_21506);
or U21848 (N_21848,N_21520,N_21748);
nor U21849 (N_21849,N_21533,N_21531);
or U21850 (N_21850,N_21604,N_21598);
and U21851 (N_21851,N_21535,N_21687);
and U21852 (N_21852,N_21660,N_21695);
or U21853 (N_21853,N_21704,N_21708);
and U21854 (N_21854,N_21614,N_21737);
and U21855 (N_21855,N_21652,N_21684);
nor U21856 (N_21856,N_21649,N_21690);
xor U21857 (N_21857,N_21505,N_21677);
nor U21858 (N_21858,N_21577,N_21557);
nand U21859 (N_21859,N_21585,N_21541);
nand U21860 (N_21860,N_21599,N_21746);
or U21861 (N_21861,N_21740,N_21551);
and U21862 (N_21862,N_21590,N_21517);
or U21863 (N_21863,N_21546,N_21723);
or U21864 (N_21864,N_21626,N_21576);
nor U21865 (N_21865,N_21528,N_21603);
nor U21866 (N_21866,N_21666,N_21663);
nor U21867 (N_21867,N_21539,N_21651);
nand U21868 (N_21868,N_21584,N_21696);
nand U21869 (N_21869,N_21735,N_21707);
or U21870 (N_21870,N_21745,N_21722);
xor U21871 (N_21871,N_21588,N_21518);
nor U21872 (N_21872,N_21547,N_21521);
nor U21873 (N_21873,N_21605,N_21579);
nand U21874 (N_21874,N_21706,N_21670);
nor U21875 (N_21875,N_21716,N_21568);
nand U21876 (N_21876,N_21639,N_21590);
and U21877 (N_21877,N_21660,N_21694);
or U21878 (N_21878,N_21632,N_21645);
nor U21879 (N_21879,N_21611,N_21574);
and U21880 (N_21880,N_21551,N_21602);
and U21881 (N_21881,N_21548,N_21735);
or U21882 (N_21882,N_21524,N_21570);
nand U21883 (N_21883,N_21509,N_21693);
nor U21884 (N_21884,N_21580,N_21600);
or U21885 (N_21885,N_21516,N_21625);
nand U21886 (N_21886,N_21529,N_21696);
nor U21887 (N_21887,N_21533,N_21667);
xnor U21888 (N_21888,N_21697,N_21748);
nand U21889 (N_21889,N_21503,N_21597);
or U21890 (N_21890,N_21533,N_21565);
and U21891 (N_21891,N_21642,N_21688);
or U21892 (N_21892,N_21500,N_21629);
and U21893 (N_21893,N_21619,N_21708);
xor U21894 (N_21894,N_21681,N_21736);
xnor U21895 (N_21895,N_21633,N_21740);
nand U21896 (N_21896,N_21689,N_21544);
nor U21897 (N_21897,N_21560,N_21603);
xor U21898 (N_21898,N_21665,N_21525);
or U21899 (N_21899,N_21701,N_21634);
and U21900 (N_21900,N_21526,N_21685);
and U21901 (N_21901,N_21579,N_21608);
nor U21902 (N_21902,N_21539,N_21727);
and U21903 (N_21903,N_21592,N_21686);
and U21904 (N_21904,N_21525,N_21567);
nor U21905 (N_21905,N_21553,N_21571);
nor U21906 (N_21906,N_21582,N_21745);
and U21907 (N_21907,N_21654,N_21747);
or U21908 (N_21908,N_21691,N_21500);
nor U21909 (N_21909,N_21591,N_21542);
nand U21910 (N_21910,N_21572,N_21504);
and U21911 (N_21911,N_21597,N_21724);
nand U21912 (N_21912,N_21715,N_21622);
nand U21913 (N_21913,N_21556,N_21583);
and U21914 (N_21914,N_21648,N_21623);
nor U21915 (N_21915,N_21606,N_21547);
or U21916 (N_21916,N_21559,N_21516);
or U21917 (N_21917,N_21610,N_21681);
or U21918 (N_21918,N_21508,N_21589);
and U21919 (N_21919,N_21506,N_21582);
or U21920 (N_21920,N_21666,N_21525);
or U21921 (N_21921,N_21672,N_21571);
or U21922 (N_21922,N_21567,N_21637);
and U21923 (N_21923,N_21591,N_21519);
nand U21924 (N_21924,N_21535,N_21639);
and U21925 (N_21925,N_21614,N_21585);
nand U21926 (N_21926,N_21682,N_21540);
nand U21927 (N_21927,N_21577,N_21546);
xor U21928 (N_21928,N_21516,N_21658);
nand U21929 (N_21929,N_21619,N_21703);
or U21930 (N_21930,N_21738,N_21537);
nor U21931 (N_21931,N_21744,N_21617);
nor U21932 (N_21932,N_21624,N_21562);
nor U21933 (N_21933,N_21744,N_21718);
nand U21934 (N_21934,N_21702,N_21662);
nand U21935 (N_21935,N_21584,N_21620);
and U21936 (N_21936,N_21571,N_21522);
nand U21937 (N_21937,N_21577,N_21537);
and U21938 (N_21938,N_21587,N_21589);
and U21939 (N_21939,N_21575,N_21505);
xnor U21940 (N_21940,N_21724,N_21646);
or U21941 (N_21941,N_21561,N_21730);
and U21942 (N_21942,N_21674,N_21645);
and U21943 (N_21943,N_21613,N_21513);
and U21944 (N_21944,N_21648,N_21748);
and U21945 (N_21945,N_21701,N_21648);
nor U21946 (N_21946,N_21733,N_21652);
xor U21947 (N_21947,N_21644,N_21581);
and U21948 (N_21948,N_21692,N_21529);
nand U21949 (N_21949,N_21707,N_21538);
nand U21950 (N_21950,N_21601,N_21605);
and U21951 (N_21951,N_21638,N_21581);
nand U21952 (N_21952,N_21591,N_21644);
or U21953 (N_21953,N_21510,N_21664);
or U21954 (N_21954,N_21634,N_21623);
xor U21955 (N_21955,N_21728,N_21637);
nor U21956 (N_21956,N_21534,N_21731);
nor U21957 (N_21957,N_21714,N_21643);
xnor U21958 (N_21958,N_21735,N_21629);
and U21959 (N_21959,N_21610,N_21684);
nor U21960 (N_21960,N_21616,N_21721);
nor U21961 (N_21961,N_21680,N_21638);
and U21962 (N_21962,N_21681,N_21660);
nor U21963 (N_21963,N_21723,N_21665);
and U21964 (N_21964,N_21578,N_21590);
and U21965 (N_21965,N_21727,N_21722);
and U21966 (N_21966,N_21733,N_21728);
nand U21967 (N_21967,N_21609,N_21646);
and U21968 (N_21968,N_21739,N_21724);
and U21969 (N_21969,N_21597,N_21734);
xnor U21970 (N_21970,N_21608,N_21611);
or U21971 (N_21971,N_21737,N_21665);
xnor U21972 (N_21972,N_21717,N_21589);
nand U21973 (N_21973,N_21624,N_21580);
nor U21974 (N_21974,N_21645,N_21627);
and U21975 (N_21975,N_21549,N_21601);
nor U21976 (N_21976,N_21742,N_21693);
nor U21977 (N_21977,N_21692,N_21516);
nand U21978 (N_21978,N_21741,N_21643);
or U21979 (N_21979,N_21716,N_21684);
or U21980 (N_21980,N_21504,N_21614);
or U21981 (N_21981,N_21729,N_21508);
xnor U21982 (N_21982,N_21572,N_21527);
and U21983 (N_21983,N_21520,N_21616);
or U21984 (N_21984,N_21643,N_21657);
nor U21985 (N_21985,N_21661,N_21553);
and U21986 (N_21986,N_21745,N_21690);
nor U21987 (N_21987,N_21588,N_21742);
nand U21988 (N_21988,N_21513,N_21628);
nor U21989 (N_21989,N_21602,N_21520);
or U21990 (N_21990,N_21616,N_21713);
nand U21991 (N_21991,N_21502,N_21662);
or U21992 (N_21992,N_21705,N_21588);
and U21993 (N_21993,N_21689,N_21537);
and U21994 (N_21994,N_21733,N_21515);
nand U21995 (N_21995,N_21676,N_21645);
or U21996 (N_21996,N_21655,N_21646);
nor U21997 (N_21997,N_21714,N_21560);
xnor U21998 (N_21998,N_21620,N_21721);
nand U21999 (N_21999,N_21673,N_21703);
or U22000 (N_22000,N_21812,N_21995);
or U22001 (N_22001,N_21755,N_21774);
and U22002 (N_22002,N_21970,N_21789);
nor U22003 (N_22003,N_21933,N_21968);
nor U22004 (N_22004,N_21967,N_21998);
or U22005 (N_22005,N_21751,N_21989);
or U22006 (N_22006,N_21969,N_21920);
or U22007 (N_22007,N_21916,N_21990);
nor U22008 (N_22008,N_21800,N_21884);
nand U22009 (N_22009,N_21823,N_21770);
and U22010 (N_22010,N_21963,N_21972);
and U22011 (N_22011,N_21831,N_21956);
or U22012 (N_22012,N_21799,N_21775);
nand U22013 (N_22013,N_21997,N_21937);
nor U22014 (N_22014,N_21826,N_21790);
xor U22015 (N_22015,N_21944,N_21830);
or U22016 (N_22016,N_21861,N_21858);
xnor U22017 (N_22017,N_21960,N_21795);
nor U22018 (N_22018,N_21763,N_21885);
and U22019 (N_22019,N_21759,N_21992);
or U22020 (N_22020,N_21864,N_21750);
nor U22021 (N_22021,N_21932,N_21982);
and U22022 (N_22022,N_21985,N_21808);
nand U22023 (N_22023,N_21881,N_21886);
nor U22024 (N_22024,N_21787,N_21895);
or U22025 (N_22025,N_21964,N_21948);
xnor U22026 (N_22026,N_21862,N_21913);
and U22027 (N_22027,N_21760,N_21804);
xor U22028 (N_22028,N_21966,N_21805);
nor U22029 (N_22029,N_21910,N_21957);
and U22030 (N_22030,N_21865,N_21902);
xor U22031 (N_22031,N_21827,N_21840);
nand U22032 (N_22032,N_21922,N_21797);
or U22033 (N_22033,N_21767,N_21941);
nand U22034 (N_22034,N_21839,N_21961);
nor U22035 (N_22035,N_21938,N_21834);
nor U22036 (N_22036,N_21946,N_21953);
nand U22037 (N_22037,N_21987,N_21842);
xnor U22038 (N_22038,N_21815,N_21757);
nand U22039 (N_22039,N_21809,N_21904);
nand U22040 (N_22040,N_21911,N_21894);
nor U22041 (N_22041,N_21859,N_21926);
nor U22042 (N_22042,N_21977,N_21768);
nand U22043 (N_22043,N_21818,N_21927);
or U22044 (N_22044,N_21955,N_21753);
and U22045 (N_22045,N_21792,N_21785);
and U22046 (N_22046,N_21841,N_21869);
and U22047 (N_22047,N_21801,N_21912);
and U22048 (N_22048,N_21848,N_21876);
nand U22049 (N_22049,N_21903,N_21929);
nor U22050 (N_22050,N_21798,N_21890);
xnor U22051 (N_22051,N_21892,N_21822);
and U22052 (N_22052,N_21984,N_21991);
or U22053 (N_22053,N_21843,N_21889);
and U22054 (N_22054,N_21762,N_21971);
nor U22055 (N_22055,N_21816,N_21891);
nand U22056 (N_22056,N_21959,N_21882);
xor U22057 (N_22057,N_21974,N_21777);
nand U22058 (N_22058,N_21878,N_21786);
or U22059 (N_22059,N_21952,N_21877);
nor U22060 (N_22060,N_21871,N_21875);
and U22061 (N_22061,N_21958,N_21752);
and U22062 (N_22062,N_21888,N_21975);
and U22063 (N_22063,N_21887,N_21907);
nand U22064 (N_22064,N_21851,N_21925);
or U22065 (N_22065,N_21979,N_21986);
nor U22066 (N_22066,N_21771,N_21921);
nor U22067 (N_22067,N_21880,N_21849);
or U22068 (N_22068,N_21973,N_21761);
and U22069 (N_22069,N_21931,N_21993);
nor U22070 (N_22070,N_21898,N_21817);
xor U22071 (N_22071,N_21819,N_21949);
or U22072 (N_22072,N_21951,N_21793);
xnor U22073 (N_22073,N_21821,N_21872);
and U22074 (N_22074,N_21778,N_21807);
nand U22075 (N_22075,N_21814,N_21847);
nand U22076 (N_22076,N_21780,N_21772);
or U22077 (N_22077,N_21838,N_21782);
nor U22078 (N_22078,N_21994,N_21873);
or U22079 (N_22079,N_21874,N_21999);
or U22080 (N_22080,N_21908,N_21914);
and U22081 (N_22081,N_21917,N_21844);
and U22082 (N_22082,N_21954,N_21923);
and U22083 (N_22083,N_21924,N_21883);
nor U22084 (N_22084,N_21835,N_21947);
or U22085 (N_22085,N_21853,N_21791);
nor U22086 (N_22086,N_21756,N_21776);
nor U22087 (N_22087,N_21996,N_21900);
and U22088 (N_22088,N_21909,N_21940);
nand U22089 (N_22089,N_21879,N_21779);
or U22090 (N_22090,N_21943,N_21802);
nor U22091 (N_22091,N_21936,N_21857);
or U22092 (N_22092,N_21813,N_21988);
nor U22093 (N_22093,N_21811,N_21983);
and U22094 (N_22094,N_21846,N_21837);
or U22095 (N_22095,N_21765,N_21784);
xnor U22096 (N_22096,N_21935,N_21764);
nor U22097 (N_22097,N_21928,N_21930);
xor U22098 (N_22098,N_21769,N_21897);
and U22099 (N_22099,N_21945,N_21773);
or U22100 (N_22100,N_21976,N_21950);
and U22101 (N_22101,N_21980,N_21833);
nor U22102 (N_22102,N_21828,N_21758);
and U22103 (N_22103,N_21829,N_21965);
or U22104 (N_22104,N_21836,N_21824);
nand U22105 (N_22105,N_21981,N_21868);
nor U22106 (N_22106,N_21810,N_21766);
nor U22107 (N_22107,N_21796,N_21934);
or U22108 (N_22108,N_21825,N_21896);
nor U22109 (N_22109,N_21942,N_21806);
and U22110 (N_22110,N_21850,N_21863);
or U22111 (N_22111,N_21905,N_21870);
and U22112 (N_22112,N_21783,N_21978);
or U22113 (N_22113,N_21860,N_21856);
nand U22114 (N_22114,N_21867,N_21919);
xor U22115 (N_22115,N_21918,N_21906);
nor U22116 (N_22116,N_21915,N_21866);
or U22117 (N_22117,N_21901,N_21832);
nor U22118 (N_22118,N_21754,N_21854);
and U22119 (N_22119,N_21852,N_21899);
nor U22120 (N_22120,N_21845,N_21820);
and U22121 (N_22121,N_21803,N_21939);
and U22122 (N_22122,N_21893,N_21794);
and U22123 (N_22123,N_21781,N_21962);
nor U22124 (N_22124,N_21788,N_21855);
or U22125 (N_22125,N_21789,N_21863);
and U22126 (N_22126,N_21867,N_21753);
nor U22127 (N_22127,N_21795,N_21782);
nor U22128 (N_22128,N_21836,N_21891);
and U22129 (N_22129,N_21921,N_21757);
nor U22130 (N_22130,N_21965,N_21844);
nor U22131 (N_22131,N_21880,N_21795);
nand U22132 (N_22132,N_21980,N_21970);
or U22133 (N_22133,N_21996,N_21990);
or U22134 (N_22134,N_21873,N_21923);
xor U22135 (N_22135,N_21758,N_21751);
or U22136 (N_22136,N_21800,N_21850);
nor U22137 (N_22137,N_21831,N_21799);
nor U22138 (N_22138,N_21999,N_21756);
and U22139 (N_22139,N_21950,N_21969);
and U22140 (N_22140,N_21871,N_21836);
or U22141 (N_22141,N_21758,N_21992);
nand U22142 (N_22142,N_21804,N_21847);
nand U22143 (N_22143,N_21917,N_21831);
and U22144 (N_22144,N_21803,N_21996);
and U22145 (N_22145,N_21836,N_21808);
nor U22146 (N_22146,N_21865,N_21864);
nand U22147 (N_22147,N_21901,N_21801);
xor U22148 (N_22148,N_21870,N_21789);
xnor U22149 (N_22149,N_21750,N_21865);
nand U22150 (N_22150,N_21807,N_21885);
nand U22151 (N_22151,N_21878,N_21935);
xor U22152 (N_22152,N_21959,N_21927);
nor U22153 (N_22153,N_21989,N_21852);
or U22154 (N_22154,N_21915,N_21827);
xnor U22155 (N_22155,N_21948,N_21917);
or U22156 (N_22156,N_21960,N_21790);
nor U22157 (N_22157,N_21914,N_21836);
or U22158 (N_22158,N_21827,N_21800);
or U22159 (N_22159,N_21760,N_21977);
nor U22160 (N_22160,N_21849,N_21989);
nor U22161 (N_22161,N_21985,N_21862);
nor U22162 (N_22162,N_21877,N_21833);
or U22163 (N_22163,N_21991,N_21924);
nand U22164 (N_22164,N_21790,N_21991);
xnor U22165 (N_22165,N_21754,N_21780);
nand U22166 (N_22166,N_21978,N_21928);
and U22167 (N_22167,N_21814,N_21934);
xor U22168 (N_22168,N_21753,N_21931);
or U22169 (N_22169,N_21961,N_21896);
and U22170 (N_22170,N_21866,N_21769);
and U22171 (N_22171,N_21865,N_21818);
xor U22172 (N_22172,N_21943,N_21797);
or U22173 (N_22173,N_21844,N_21846);
and U22174 (N_22174,N_21970,N_21895);
xor U22175 (N_22175,N_21811,N_21838);
and U22176 (N_22176,N_21823,N_21972);
and U22177 (N_22177,N_21818,N_21782);
or U22178 (N_22178,N_21939,N_21775);
nor U22179 (N_22179,N_21838,N_21757);
xor U22180 (N_22180,N_21991,N_21963);
nand U22181 (N_22181,N_21903,N_21963);
or U22182 (N_22182,N_21774,N_21949);
nand U22183 (N_22183,N_21897,N_21751);
nor U22184 (N_22184,N_21916,N_21895);
nand U22185 (N_22185,N_21840,N_21932);
or U22186 (N_22186,N_21995,N_21756);
nand U22187 (N_22187,N_21967,N_21836);
nor U22188 (N_22188,N_21787,N_21845);
and U22189 (N_22189,N_21948,N_21909);
or U22190 (N_22190,N_21777,N_21790);
or U22191 (N_22191,N_21819,N_21933);
and U22192 (N_22192,N_21794,N_21973);
and U22193 (N_22193,N_21902,N_21984);
or U22194 (N_22194,N_21954,N_21835);
and U22195 (N_22195,N_21982,N_21858);
nor U22196 (N_22196,N_21784,N_21993);
and U22197 (N_22197,N_21841,N_21911);
xnor U22198 (N_22198,N_21868,N_21781);
nand U22199 (N_22199,N_21841,N_21810);
xnor U22200 (N_22200,N_21825,N_21773);
nor U22201 (N_22201,N_21881,N_21866);
and U22202 (N_22202,N_21937,N_21811);
or U22203 (N_22203,N_21878,N_21899);
nand U22204 (N_22204,N_21803,N_21765);
or U22205 (N_22205,N_21883,N_21870);
xnor U22206 (N_22206,N_21796,N_21878);
nand U22207 (N_22207,N_21974,N_21799);
or U22208 (N_22208,N_21771,N_21935);
or U22209 (N_22209,N_21985,N_21860);
nor U22210 (N_22210,N_21988,N_21820);
nor U22211 (N_22211,N_21830,N_21951);
nor U22212 (N_22212,N_21886,N_21900);
and U22213 (N_22213,N_21828,N_21929);
or U22214 (N_22214,N_21905,N_21894);
or U22215 (N_22215,N_21976,N_21790);
nor U22216 (N_22216,N_21903,N_21827);
and U22217 (N_22217,N_21972,N_21785);
nor U22218 (N_22218,N_21845,N_21968);
and U22219 (N_22219,N_21985,N_21891);
or U22220 (N_22220,N_21906,N_21832);
nand U22221 (N_22221,N_21911,N_21851);
xor U22222 (N_22222,N_21898,N_21900);
and U22223 (N_22223,N_21947,N_21933);
and U22224 (N_22224,N_21820,N_21788);
or U22225 (N_22225,N_21922,N_21752);
or U22226 (N_22226,N_21920,N_21767);
or U22227 (N_22227,N_21761,N_21776);
nor U22228 (N_22228,N_21898,N_21848);
and U22229 (N_22229,N_21886,N_21925);
and U22230 (N_22230,N_21903,N_21818);
nor U22231 (N_22231,N_21829,N_21956);
xor U22232 (N_22232,N_21973,N_21830);
or U22233 (N_22233,N_21773,N_21906);
nor U22234 (N_22234,N_21780,N_21824);
nor U22235 (N_22235,N_21896,N_21758);
nand U22236 (N_22236,N_21903,N_21994);
and U22237 (N_22237,N_21828,N_21893);
or U22238 (N_22238,N_21892,N_21905);
nand U22239 (N_22239,N_21893,N_21829);
or U22240 (N_22240,N_21994,N_21769);
and U22241 (N_22241,N_21817,N_21838);
and U22242 (N_22242,N_21909,N_21770);
and U22243 (N_22243,N_21994,N_21939);
and U22244 (N_22244,N_21772,N_21868);
nand U22245 (N_22245,N_21920,N_21899);
nor U22246 (N_22246,N_21800,N_21910);
or U22247 (N_22247,N_21875,N_21892);
nor U22248 (N_22248,N_21973,N_21930);
xor U22249 (N_22249,N_21943,N_21785);
nor U22250 (N_22250,N_22160,N_22077);
and U22251 (N_22251,N_22125,N_22248);
or U22252 (N_22252,N_22226,N_22026);
or U22253 (N_22253,N_22153,N_22146);
nor U22254 (N_22254,N_22064,N_22011);
nor U22255 (N_22255,N_22196,N_22131);
nor U22256 (N_22256,N_22169,N_22166);
nand U22257 (N_22257,N_22022,N_22006);
and U22258 (N_22258,N_22200,N_22052);
nor U22259 (N_22259,N_22147,N_22163);
nand U22260 (N_22260,N_22055,N_22034);
or U22261 (N_22261,N_22050,N_22079);
or U22262 (N_22262,N_22193,N_22175);
nor U22263 (N_22263,N_22205,N_22121);
or U22264 (N_22264,N_22112,N_22132);
or U22265 (N_22265,N_22224,N_22211);
and U22266 (N_22266,N_22056,N_22015);
nor U22267 (N_22267,N_22029,N_22133);
nor U22268 (N_22268,N_22094,N_22066);
or U22269 (N_22269,N_22234,N_22012);
nor U22270 (N_22270,N_22092,N_22067);
nor U22271 (N_22271,N_22217,N_22018);
nor U22272 (N_22272,N_22148,N_22020);
nor U22273 (N_22273,N_22222,N_22192);
xnor U22274 (N_22274,N_22204,N_22157);
or U22275 (N_22275,N_22093,N_22209);
nand U22276 (N_22276,N_22127,N_22110);
or U22277 (N_22277,N_22071,N_22098);
nor U22278 (N_22278,N_22138,N_22244);
nor U22279 (N_22279,N_22025,N_22048);
or U22280 (N_22280,N_22164,N_22075);
and U22281 (N_22281,N_22197,N_22241);
xor U22282 (N_22282,N_22177,N_22059);
xnor U22283 (N_22283,N_22158,N_22060);
and U22284 (N_22284,N_22027,N_22028);
or U22285 (N_22285,N_22238,N_22199);
and U22286 (N_22286,N_22046,N_22171);
or U22287 (N_22287,N_22231,N_22080);
nand U22288 (N_22288,N_22201,N_22172);
nor U22289 (N_22289,N_22150,N_22096);
nor U22290 (N_22290,N_22030,N_22017);
nor U22291 (N_22291,N_22188,N_22249);
nor U22292 (N_22292,N_22154,N_22237);
nand U22293 (N_22293,N_22165,N_22085);
nor U22294 (N_22294,N_22207,N_22223);
nand U22295 (N_22295,N_22108,N_22101);
and U22296 (N_22296,N_22024,N_22074);
nand U22297 (N_22297,N_22116,N_22004);
and U22298 (N_22298,N_22083,N_22062);
nor U22299 (N_22299,N_22161,N_22078);
and U22300 (N_22300,N_22016,N_22123);
nor U22301 (N_22301,N_22183,N_22118);
or U22302 (N_22302,N_22076,N_22242);
nor U22303 (N_22303,N_22245,N_22122);
nand U22304 (N_22304,N_22103,N_22182);
nand U22305 (N_22305,N_22065,N_22220);
nor U22306 (N_22306,N_22229,N_22097);
and U22307 (N_22307,N_22106,N_22117);
and U22308 (N_22308,N_22187,N_22124);
and U22309 (N_22309,N_22084,N_22159);
nor U22310 (N_22310,N_22023,N_22049);
nand U22311 (N_22311,N_22168,N_22152);
nand U22312 (N_22312,N_22235,N_22202);
and U22313 (N_22313,N_22082,N_22212);
or U22314 (N_22314,N_22007,N_22215);
nor U22315 (N_22315,N_22019,N_22038);
and U22316 (N_22316,N_22173,N_22151);
nand U22317 (N_22317,N_22128,N_22099);
and U22318 (N_22318,N_22115,N_22195);
or U22319 (N_22319,N_22070,N_22189);
nor U22320 (N_22320,N_22013,N_22180);
nand U22321 (N_22321,N_22031,N_22185);
or U22322 (N_22322,N_22156,N_22134);
nor U22323 (N_22323,N_22051,N_22179);
and U22324 (N_22324,N_22032,N_22144);
and U22325 (N_22325,N_22073,N_22155);
and U22326 (N_22326,N_22184,N_22221);
and U22327 (N_22327,N_22087,N_22143);
nor U22328 (N_22328,N_22109,N_22044);
nor U22329 (N_22329,N_22176,N_22054);
nor U22330 (N_22330,N_22010,N_22061);
nor U22331 (N_22331,N_22174,N_22053);
or U22332 (N_22332,N_22203,N_22063);
or U22333 (N_22333,N_22130,N_22045);
nor U22334 (N_22334,N_22047,N_22145);
or U22335 (N_22335,N_22005,N_22002);
nand U22336 (N_22336,N_22039,N_22001);
or U22337 (N_22337,N_22190,N_22178);
or U22338 (N_22338,N_22068,N_22000);
or U22339 (N_22339,N_22072,N_22233);
nand U22340 (N_22340,N_22236,N_22230);
or U22341 (N_22341,N_22239,N_22043);
nand U22342 (N_22342,N_22009,N_22170);
or U22343 (N_22343,N_22058,N_22141);
and U22344 (N_22344,N_22186,N_22014);
nor U22345 (N_22345,N_22240,N_22140);
nor U22346 (N_22346,N_22088,N_22129);
or U22347 (N_22347,N_22191,N_22021);
or U22348 (N_22348,N_22081,N_22003);
and U22349 (N_22349,N_22210,N_22126);
and U22350 (N_22350,N_22162,N_22095);
nor U22351 (N_22351,N_22033,N_22206);
nor U22352 (N_22352,N_22246,N_22137);
or U22353 (N_22353,N_22213,N_22036);
or U22354 (N_22354,N_22090,N_22104);
nand U22355 (N_22355,N_22089,N_22119);
and U22356 (N_22356,N_22194,N_22136);
and U22357 (N_22357,N_22105,N_22069);
nand U22358 (N_22358,N_22139,N_22142);
nand U22359 (N_22359,N_22214,N_22113);
nor U22360 (N_22360,N_22167,N_22086);
nor U22361 (N_22361,N_22225,N_22218);
or U22362 (N_22362,N_22111,N_22042);
or U22363 (N_22363,N_22091,N_22107);
and U22364 (N_22364,N_22041,N_22040);
nand U22365 (N_22365,N_22114,N_22035);
or U22366 (N_22366,N_22198,N_22243);
and U22367 (N_22367,N_22181,N_22219);
and U22368 (N_22368,N_22135,N_22149);
and U22369 (N_22369,N_22120,N_22232);
and U22370 (N_22370,N_22037,N_22227);
or U22371 (N_22371,N_22057,N_22247);
nand U22372 (N_22372,N_22228,N_22102);
nor U22373 (N_22373,N_22100,N_22216);
xor U22374 (N_22374,N_22008,N_22208);
nand U22375 (N_22375,N_22081,N_22077);
nor U22376 (N_22376,N_22155,N_22093);
and U22377 (N_22377,N_22120,N_22002);
or U22378 (N_22378,N_22004,N_22050);
nand U22379 (N_22379,N_22016,N_22025);
nand U22380 (N_22380,N_22171,N_22081);
xnor U22381 (N_22381,N_22222,N_22070);
or U22382 (N_22382,N_22007,N_22145);
or U22383 (N_22383,N_22053,N_22038);
nor U22384 (N_22384,N_22164,N_22045);
nor U22385 (N_22385,N_22002,N_22129);
or U22386 (N_22386,N_22020,N_22092);
and U22387 (N_22387,N_22234,N_22122);
nand U22388 (N_22388,N_22093,N_22178);
nand U22389 (N_22389,N_22054,N_22239);
xnor U22390 (N_22390,N_22110,N_22139);
nand U22391 (N_22391,N_22152,N_22151);
or U22392 (N_22392,N_22080,N_22200);
nor U22393 (N_22393,N_22235,N_22142);
or U22394 (N_22394,N_22174,N_22181);
nor U22395 (N_22395,N_22052,N_22210);
and U22396 (N_22396,N_22107,N_22210);
nor U22397 (N_22397,N_22067,N_22179);
nand U22398 (N_22398,N_22023,N_22111);
nor U22399 (N_22399,N_22244,N_22021);
nor U22400 (N_22400,N_22098,N_22226);
xnor U22401 (N_22401,N_22207,N_22092);
nand U22402 (N_22402,N_22052,N_22211);
and U22403 (N_22403,N_22067,N_22055);
nor U22404 (N_22404,N_22057,N_22194);
and U22405 (N_22405,N_22187,N_22077);
or U22406 (N_22406,N_22024,N_22037);
xor U22407 (N_22407,N_22026,N_22175);
or U22408 (N_22408,N_22102,N_22148);
and U22409 (N_22409,N_22024,N_22144);
xor U22410 (N_22410,N_22104,N_22230);
nor U22411 (N_22411,N_22144,N_22033);
or U22412 (N_22412,N_22155,N_22238);
nand U22413 (N_22413,N_22192,N_22246);
xnor U22414 (N_22414,N_22034,N_22234);
nand U22415 (N_22415,N_22207,N_22104);
or U22416 (N_22416,N_22161,N_22006);
and U22417 (N_22417,N_22004,N_22052);
or U22418 (N_22418,N_22188,N_22027);
and U22419 (N_22419,N_22136,N_22144);
and U22420 (N_22420,N_22166,N_22192);
or U22421 (N_22421,N_22105,N_22073);
or U22422 (N_22422,N_22146,N_22073);
nand U22423 (N_22423,N_22154,N_22087);
or U22424 (N_22424,N_22078,N_22057);
nor U22425 (N_22425,N_22173,N_22116);
and U22426 (N_22426,N_22116,N_22193);
and U22427 (N_22427,N_22028,N_22227);
and U22428 (N_22428,N_22011,N_22102);
nor U22429 (N_22429,N_22191,N_22136);
or U22430 (N_22430,N_22178,N_22136);
and U22431 (N_22431,N_22006,N_22234);
or U22432 (N_22432,N_22206,N_22000);
nor U22433 (N_22433,N_22213,N_22165);
or U22434 (N_22434,N_22104,N_22084);
or U22435 (N_22435,N_22194,N_22107);
nor U22436 (N_22436,N_22063,N_22021);
nor U22437 (N_22437,N_22047,N_22008);
nand U22438 (N_22438,N_22025,N_22070);
xor U22439 (N_22439,N_22114,N_22170);
nand U22440 (N_22440,N_22110,N_22162);
xor U22441 (N_22441,N_22107,N_22049);
nand U22442 (N_22442,N_22067,N_22087);
or U22443 (N_22443,N_22162,N_22101);
or U22444 (N_22444,N_22078,N_22195);
nand U22445 (N_22445,N_22174,N_22113);
and U22446 (N_22446,N_22067,N_22029);
or U22447 (N_22447,N_22226,N_22021);
and U22448 (N_22448,N_22026,N_22091);
nand U22449 (N_22449,N_22093,N_22032);
nand U22450 (N_22450,N_22016,N_22026);
and U22451 (N_22451,N_22244,N_22049);
nand U22452 (N_22452,N_22183,N_22152);
nor U22453 (N_22453,N_22097,N_22140);
and U22454 (N_22454,N_22097,N_22238);
nor U22455 (N_22455,N_22024,N_22216);
or U22456 (N_22456,N_22099,N_22182);
nand U22457 (N_22457,N_22037,N_22172);
and U22458 (N_22458,N_22054,N_22211);
or U22459 (N_22459,N_22243,N_22082);
or U22460 (N_22460,N_22000,N_22053);
and U22461 (N_22461,N_22067,N_22020);
nand U22462 (N_22462,N_22016,N_22175);
nor U22463 (N_22463,N_22063,N_22243);
or U22464 (N_22464,N_22100,N_22171);
nand U22465 (N_22465,N_22060,N_22170);
nor U22466 (N_22466,N_22129,N_22132);
or U22467 (N_22467,N_22140,N_22098);
nand U22468 (N_22468,N_22234,N_22021);
and U22469 (N_22469,N_22228,N_22230);
or U22470 (N_22470,N_22187,N_22042);
or U22471 (N_22471,N_22235,N_22165);
or U22472 (N_22472,N_22105,N_22206);
and U22473 (N_22473,N_22095,N_22158);
or U22474 (N_22474,N_22189,N_22221);
and U22475 (N_22475,N_22125,N_22148);
and U22476 (N_22476,N_22234,N_22248);
nand U22477 (N_22477,N_22072,N_22079);
or U22478 (N_22478,N_22055,N_22181);
nor U22479 (N_22479,N_22062,N_22099);
and U22480 (N_22480,N_22238,N_22154);
nor U22481 (N_22481,N_22224,N_22200);
or U22482 (N_22482,N_22145,N_22159);
nor U22483 (N_22483,N_22203,N_22175);
xnor U22484 (N_22484,N_22137,N_22158);
xnor U22485 (N_22485,N_22231,N_22128);
nor U22486 (N_22486,N_22147,N_22198);
or U22487 (N_22487,N_22157,N_22216);
and U22488 (N_22488,N_22115,N_22008);
nand U22489 (N_22489,N_22061,N_22117);
and U22490 (N_22490,N_22112,N_22012);
xnor U22491 (N_22491,N_22208,N_22184);
or U22492 (N_22492,N_22093,N_22085);
xor U22493 (N_22493,N_22137,N_22047);
nor U22494 (N_22494,N_22055,N_22101);
nand U22495 (N_22495,N_22212,N_22073);
and U22496 (N_22496,N_22026,N_22217);
nor U22497 (N_22497,N_22023,N_22244);
nor U22498 (N_22498,N_22157,N_22123);
xnor U22499 (N_22499,N_22045,N_22034);
xnor U22500 (N_22500,N_22420,N_22259);
and U22501 (N_22501,N_22365,N_22432);
and U22502 (N_22502,N_22343,N_22421);
nor U22503 (N_22503,N_22426,N_22256);
or U22504 (N_22504,N_22311,N_22443);
nor U22505 (N_22505,N_22285,N_22358);
or U22506 (N_22506,N_22368,N_22482);
xor U22507 (N_22507,N_22377,N_22332);
xnor U22508 (N_22508,N_22264,N_22401);
or U22509 (N_22509,N_22307,N_22354);
nor U22510 (N_22510,N_22488,N_22429);
or U22511 (N_22511,N_22312,N_22396);
xor U22512 (N_22512,N_22331,N_22308);
nor U22513 (N_22513,N_22323,N_22367);
xnor U22514 (N_22514,N_22437,N_22398);
nor U22515 (N_22515,N_22340,N_22382);
and U22516 (N_22516,N_22250,N_22469);
and U22517 (N_22517,N_22444,N_22355);
and U22518 (N_22518,N_22471,N_22325);
nand U22519 (N_22519,N_22497,N_22288);
nand U22520 (N_22520,N_22484,N_22479);
nand U22521 (N_22521,N_22392,N_22274);
nand U22522 (N_22522,N_22269,N_22347);
nor U22523 (N_22523,N_22334,N_22427);
or U22524 (N_22524,N_22478,N_22456);
and U22525 (N_22525,N_22493,N_22295);
or U22526 (N_22526,N_22492,N_22321);
xnor U22527 (N_22527,N_22359,N_22489);
and U22528 (N_22528,N_22273,N_22362);
xnor U22529 (N_22529,N_22291,N_22394);
nand U22530 (N_22530,N_22294,N_22279);
and U22531 (N_22531,N_22281,N_22389);
nand U22532 (N_22532,N_22344,N_22267);
nor U22533 (N_22533,N_22298,N_22387);
and U22534 (N_22534,N_22391,N_22485);
and U22535 (N_22535,N_22254,N_22322);
or U22536 (N_22536,N_22345,N_22413);
nor U22537 (N_22537,N_22402,N_22495);
nand U22538 (N_22538,N_22341,N_22491);
nand U22539 (N_22539,N_22380,N_22449);
or U22540 (N_22540,N_22350,N_22370);
nand U22541 (N_22541,N_22318,N_22352);
nor U22542 (N_22542,N_22494,N_22351);
and U22543 (N_22543,N_22319,N_22463);
nand U22544 (N_22544,N_22460,N_22303);
nand U22545 (N_22545,N_22376,N_22328);
nand U22546 (N_22546,N_22446,N_22476);
xor U22547 (N_22547,N_22473,N_22409);
and U22548 (N_22548,N_22379,N_22299);
nor U22549 (N_22549,N_22272,N_22411);
and U22550 (N_22550,N_22356,N_22378);
nor U22551 (N_22551,N_22405,N_22470);
xnor U22552 (N_22552,N_22324,N_22410);
nor U22553 (N_22553,N_22252,N_22258);
or U22554 (N_22554,N_22422,N_22255);
nor U22555 (N_22555,N_22280,N_22305);
or U22556 (N_22556,N_22498,N_22459);
xnor U22557 (N_22557,N_22468,N_22373);
nand U22558 (N_22558,N_22477,N_22284);
nand U22559 (N_22559,N_22461,N_22474);
xor U22560 (N_22560,N_22266,N_22363);
and U22561 (N_22561,N_22458,N_22399);
nand U22562 (N_22562,N_22374,N_22412);
and U22563 (N_22563,N_22403,N_22466);
and U22564 (N_22564,N_22360,N_22270);
nand U22565 (N_22565,N_22440,N_22293);
nand U22566 (N_22566,N_22261,N_22447);
nor U22567 (N_22567,N_22297,N_22278);
nand U22568 (N_22568,N_22357,N_22407);
nor U22569 (N_22569,N_22381,N_22450);
nor U22570 (N_22570,N_22486,N_22283);
and U22571 (N_22571,N_22408,N_22275);
and U22572 (N_22572,N_22309,N_22304);
nand U22573 (N_22573,N_22435,N_22472);
nand U22574 (N_22574,N_22263,N_22465);
nor U22575 (N_22575,N_22251,N_22336);
xnor U22576 (N_22576,N_22260,N_22433);
xor U22577 (N_22577,N_22310,N_22454);
nor U22578 (N_22578,N_22296,N_22384);
or U22579 (N_22579,N_22430,N_22404);
nor U22580 (N_22580,N_22400,N_22349);
or U22581 (N_22581,N_22397,N_22306);
nor U22582 (N_22582,N_22483,N_22439);
nor U22583 (N_22583,N_22438,N_22496);
or U22584 (N_22584,N_22369,N_22346);
nand U22585 (N_22585,N_22320,N_22316);
nand U22586 (N_22586,N_22366,N_22480);
nor U22587 (N_22587,N_22462,N_22428);
nor U22588 (N_22588,N_22499,N_22395);
nor U22589 (N_22589,N_22327,N_22414);
nand U22590 (N_22590,N_22424,N_22431);
nand U22591 (N_22591,N_22330,N_22406);
xor U22592 (N_22592,N_22417,N_22451);
nor U22593 (N_22593,N_22385,N_22475);
nand U22594 (N_22594,N_22372,N_22300);
and U22595 (N_22595,N_22289,N_22353);
or U22596 (N_22596,N_22448,N_22388);
nor U22597 (N_22597,N_22423,N_22277);
nand U22598 (N_22598,N_22361,N_22425);
or U22599 (N_22599,N_22442,N_22271);
or U22600 (N_22600,N_22490,N_22386);
or U22601 (N_22601,N_22290,N_22419);
nor U22602 (N_22602,N_22457,N_22276);
nand U22603 (N_22603,N_22282,N_22464);
and U22604 (N_22604,N_22302,N_22467);
or U22605 (N_22605,N_22416,N_22329);
and U22606 (N_22606,N_22393,N_22415);
or U22607 (N_22607,N_22265,N_22326);
nand U22608 (N_22608,N_22418,N_22487);
nand U22609 (N_22609,N_22338,N_22434);
nand U22610 (N_22610,N_22436,N_22253);
nand U22611 (N_22611,N_22262,N_22453);
xor U22612 (N_22612,N_22301,N_22390);
or U22613 (N_22613,N_22371,N_22286);
and U22614 (N_22614,N_22348,N_22337);
and U22615 (N_22615,N_22339,N_22481);
and U22616 (N_22616,N_22452,N_22335);
or U22617 (N_22617,N_22314,N_22441);
or U22618 (N_22618,N_22383,N_22375);
nand U22619 (N_22619,N_22364,N_22292);
and U22620 (N_22620,N_22313,N_22333);
nand U22621 (N_22621,N_22315,N_22317);
nor U22622 (N_22622,N_22268,N_22257);
and U22623 (N_22623,N_22455,N_22342);
and U22624 (N_22624,N_22445,N_22287);
nand U22625 (N_22625,N_22436,N_22299);
nand U22626 (N_22626,N_22300,N_22448);
nor U22627 (N_22627,N_22411,N_22310);
or U22628 (N_22628,N_22499,N_22315);
nor U22629 (N_22629,N_22391,N_22358);
nor U22630 (N_22630,N_22260,N_22348);
and U22631 (N_22631,N_22438,N_22384);
and U22632 (N_22632,N_22263,N_22353);
nand U22633 (N_22633,N_22382,N_22361);
or U22634 (N_22634,N_22322,N_22403);
and U22635 (N_22635,N_22490,N_22285);
or U22636 (N_22636,N_22340,N_22264);
and U22637 (N_22637,N_22307,N_22318);
nand U22638 (N_22638,N_22460,N_22350);
and U22639 (N_22639,N_22445,N_22487);
and U22640 (N_22640,N_22263,N_22379);
nand U22641 (N_22641,N_22310,N_22267);
or U22642 (N_22642,N_22298,N_22486);
or U22643 (N_22643,N_22326,N_22472);
nor U22644 (N_22644,N_22429,N_22326);
and U22645 (N_22645,N_22273,N_22470);
nor U22646 (N_22646,N_22438,N_22352);
nor U22647 (N_22647,N_22443,N_22455);
or U22648 (N_22648,N_22375,N_22432);
or U22649 (N_22649,N_22454,N_22401);
nor U22650 (N_22650,N_22416,N_22402);
or U22651 (N_22651,N_22279,N_22429);
xnor U22652 (N_22652,N_22284,N_22285);
and U22653 (N_22653,N_22396,N_22304);
and U22654 (N_22654,N_22274,N_22393);
or U22655 (N_22655,N_22300,N_22286);
and U22656 (N_22656,N_22377,N_22474);
and U22657 (N_22657,N_22474,N_22447);
and U22658 (N_22658,N_22343,N_22493);
nor U22659 (N_22659,N_22332,N_22405);
nand U22660 (N_22660,N_22417,N_22407);
xor U22661 (N_22661,N_22409,N_22255);
nand U22662 (N_22662,N_22269,N_22349);
and U22663 (N_22663,N_22354,N_22403);
nand U22664 (N_22664,N_22316,N_22252);
and U22665 (N_22665,N_22476,N_22441);
or U22666 (N_22666,N_22493,N_22480);
or U22667 (N_22667,N_22426,N_22310);
nor U22668 (N_22668,N_22265,N_22485);
or U22669 (N_22669,N_22493,N_22252);
and U22670 (N_22670,N_22349,N_22263);
nand U22671 (N_22671,N_22267,N_22449);
or U22672 (N_22672,N_22480,N_22388);
and U22673 (N_22673,N_22469,N_22359);
nand U22674 (N_22674,N_22381,N_22271);
nand U22675 (N_22675,N_22276,N_22355);
or U22676 (N_22676,N_22346,N_22312);
nand U22677 (N_22677,N_22317,N_22418);
and U22678 (N_22678,N_22472,N_22459);
xor U22679 (N_22679,N_22278,N_22313);
and U22680 (N_22680,N_22306,N_22398);
nor U22681 (N_22681,N_22499,N_22455);
nor U22682 (N_22682,N_22445,N_22384);
xor U22683 (N_22683,N_22329,N_22458);
nor U22684 (N_22684,N_22380,N_22357);
nor U22685 (N_22685,N_22283,N_22360);
nand U22686 (N_22686,N_22253,N_22467);
and U22687 (N_22687,N_22303,N_22490);
and U22688 (N_22688,N_22269,N_22429);
and U22689 (N_22689,N_22292,N_22493);
or U22690 (N_22690,N_22251,N_22402);
nand U22691 (N_22691,N_22270,N_22292);
or U22692 (N_22692,N_22339,N_22334);
and U22693 (N_22693,N_22492,N_22411);
nand U22694 (N_22694,N_22379,N_22431);
and U22695 (N_22695,N_22333,N_22312);
nor U22696 (N_22696,N_22264,N_22465);
or U22697 (N_22697,N_22468,N_22270);
nand U22698 (N_22698,N_22409,N_22456);
or U22699 (N_22699,N_22468,N_22445);
and U22700 (N_22700,N_22347,N_22373);
and U22701 (N_22701,N_22321,N_22269);
and U22702 (N_22702,N_22269,N_22460);
and U22703 (N_22703,N_22484,N_22318);
nand U22704 (N_22704,N_22285,N_22292);
and U22705 (N_22705,N_22277,N_22304);
and U22706 (N_22706,N_22348,N_22476);
or U22707 (N_22707,N_22314,N_22358);
or U22708 (N_22708,N_22399,N_22331);
nor U22709 (N_22709,N_22435,N_22258);
nor U22710 (N_22710,N_22407,N_22268);
and U22711 (N_22711,N_22355,N_22489);
and U22712 (N_22712,N_22350,N_22462);
xor U22713 (N_22713,N_22352,N_22403);
xor U22714 (N_22714,N_22457,N_22266);
nand U22715 (N_22715,N_22427,N_22280);
or U22716 (N_22716,N_22446,N_22396);
or U22717 (N_22717,N_22453,N_22274);
or U22718 (N_22718,N_22349,N_22466);
xnor U22719 (N_22719,N_22263,N_22439);
or U22720 (N_22720,N_22379,N_22440);
nor U22721 (N_22721,N_22311,N_22418);
nor U22722 (N_22722,N_22314,N_22399);
nand U22723 (N_22723,N_22448,N_22433);
or U22724 (N_22724,N_22264,N_22289);
nand U22725 (N_22725,N_22371,N_22440);
or U22726 (N_22726,N_22281,N_22319);
and U22727 (N_22727,N_22399,N_22334);
and U22728 (N_22728,N_22284,N_22313);
and U22729 (N_22729,N_22456,N_22344);
or U22730 (N_22730,N_22463,N_22271);
and U22731 (N_22731,N_22467,N_22418);
nand U22732 (N_22732,N_22436,N_22347);
nor U22733 (N_22733,N_22369,N_22475);
xor U22734 (N_22734,N_22299,N_22471);
nand U22735 (N_22735,N_22374,N_22423);
and U22736 (N_22736,N_22271,N_22462);
or U22737 (N_22737,N_22496,N_22309);
or U22738 (N_22738,N_22375,N_22446);
or U22739 (N_22739,N_22283,N_22296);
or U22740 (N_22740,N_22424,N_22264);
or U22741 (N_22741,N_22369,N_22374);
or U22742 (N_22742,N_22310,N_22338);
or U22743 (N_22743,N_22317,N_22362);
nor U22744 (N_22744,N_22266,N_22418);
nor U22745 (N_22745,N_22413,N_22467);
nor U22746 (N_22746,N_22325,N_22350);
nor U22747 (N_22747,N_22362,N_22324);
or U22748 (N_22748,N_22348,N_22394);
nor U22749 (N_22749,N_22400,N_22297);
and U22750 (N_22750,N_22568,N_22586);
xor U22751 (N_22751,N_22621,N_22613);
or U22752 (N_22752,N_22683,N_22670);
and U22753 (N_22753,N_22561,N_22678);
and U22754 (N_22754,N_22713,N_22714);
and U22755 (N_22755,N_22723,N_22605);
nand U22756 (N_22756,N_22644,N_22533);
nand U22757 (N_22757,N_22588,N_22708);
and U22758 (N_22758,N_22570,N_22550);
nand U22759 (N_22759,N_22579,N_22505);
and U22760 (N_22760,N_22688,N_22659);
and U22761 (N_22761,N_22735,N_22686);
nor U22762 (N_22762,N_22571,N_22652);
nor U22763 (N_22763,N_22709,N_22639);
or U22764 (N_22764,N_22573,N_22749);
and U22765 (N_22765,N_22508,N_22632);
or U22766 (N_22766,N_22675,N_22507);
nor U22767 (N_22767,N_22737,N_22656);
xor U22768 (N_22768,N_22562,N_22720);
and U22769 (N_22769,N_22619,N_22515);
nor U22770 (N_22770,N_22549,N_22685);
and U22771 (N_22771,N_22544,N_22576);
xnor U22772 (N_22772,N_22698,N_22551);
nor U22773 (N_22773,N_22651,N_22597);
nand U22774 (N_22774,N_22658,N_22635);
or U22775 (N_22775,N_22691,N_22612);
and U22776 (N_22776,N_22682,N_22733);
or U22777 (N_22777,N_22643,N_22578);
nand U22778 (N_22778,N_22542,N_22598);
and U22779 (N_22779,N_22523,N_22673);
nand U22780 (N_22780,N_22717,N_22539);
nand U22781 (N_22781,N_22731,N_22648);
and U22782 (N_22782,N_22694,N_22501);
or U22783 (N_22783,N_22596,N_22581);
xor U22784 (N_22784,N_22564,N_22693);
and U22785 (N_22785,N_22603,N_22585);
nand U22786 (N_22786,N_22524,N_22679);
nor U22787 (N_22787,N_22608,N_22728);
and U22788 (N_22788,N_22663,N_22594);
nor U22789 (N_22789,N_22672,N_22531);
nand U22790 (N_22790,N_22512,N_22516);
and U22791 (N_22791,N_22620,N_22530);
and U22792 (N_22792,N_22525,N_22640);
and U22793 (N_22793,N_22615,N_22616);
nand U22794 (N_22794,N_22702,N_22521);
and U22795 (N_22795,N_22725,N_22610);
nor U22796 (N_22796,N_22569,N_22747);
nand U22797 (N_22797,N_22538,N_22669);
nor U22798 (N_22798,N_22695,N_22630);
and U22799 (N_22799,N_22722,N_22633);
xor U22800 (N_22800,N_22537,N_22556);
xnor U22801 (N_22801,N_22591,N_22730);
and U22802 (N_22802,N_22677,N_22684);
xor U22803 (N_22803,N_22736,N_22590);
nor U22804 (N_22804,N_22503,N_22528);
and U22805 (N_22805,N_22552,N_22706);
or U22806 (N_22806,N_22506,N_22710);
nand U22807 (N_22807,N_22554,N_22522);
or U22808 (N_22808,N_22606,N_22664);
xnor U22809 (N_22809,N_22583,N_22517);
nand U22810 (N_22810,N_22641,N_22607);
or U22811 (N_22811,N_22744,N_22726);
or U22812 (N_22812,N_22721,N_22614);
and U22813 (N_22813,N_22666,N_22631);
or U22814 (N_22814,N_22611,N_22657);
nor U22815 (N_22815,N_22662,N_22734);
nand U22816 (N_22816,N_22689,N_22577);
or U22817 (N_22817,N_22676,N_22638);
and U22818 (N_22818,N_22500,N_22526);
or U22819 (N_22819,N_22534,N_22604);
or U22820 (N_22820,N_22584,N_22547);
nor U22821 (N_22821,N_22599,N_22671);
and U22822 (N_22822,N_22540,N_22558);
and U22823 (N_22823,N_22582,N_22545);
or U22824 (N_22824,N_22541,N_22642);
or U22825 (N_22825,N_22668,N_22511);
or U22826 (N_22826,N_22575,N_22535);
nand U22827 (N_22827,N_22715,N_22626);
xor U22828 (N_22828,N_22567,N_22649);
or U22829 (N_22829,N_22628,N_22543);
or U22830 (N_22830,N_22574,N_22680);
or U22831 (N_22831,N_22687,N_22654);
and U22832 (N_22832,N_22636,N_22513);
nor U22833 (N_22833,N_22529,N_22559);
nand U22834 (N_22834,N_22510,N_22661);
nor U22835 (N_22835,N_22719,N_22690);
nor U22836 (N_22836,N_22716,N_22520);
and U22837 (N_22837,N_22646,N_22718);
nand U22838 (N_22838,N_22637,N_22699);
and U22839 (N_22839,N_22625,N_22692);
xnor U22840 (N_22840,N_22572,N_22509);
xnor U22841 (N_22841,N_22742,N_22667);
and U22842 (N_22842,N_22622,N_22623);
and U22843 (N_22843,N_22563,N_22727);
and U22844 (N_22844,N_22660,N_22624);
nand U22845 (N_22845,N_22743,N_22697);
and U22846 (N_22846,N_22645,N_22729);
nor U22847 (N_22847,N_22711,N_22674);
nand U22848 (N_22848,N_22592,N_22665);
nand U22849 (N_22849,N_22740,N_22724);
or U22850 (N_22850,N_22555,N_22518);
nand U22851 (N_22851,N_22600,N_22593);
nand U22852 (N_22852,N_22629,N_22560);
or U22853 (N_22853,N_22704,N_22601);
nand U22854 (N_22854,N_22748,N_22587);
nand U22855 (N_22855,N_22504,N_22746);
or U22856 (N_22856,N_22527,N_22536);
or U22857 (N_22857,N_22609,N_22566);
or U22858 (N_22858,N_22532,N_22738);
or U22859 (N_22859,N_22589,N_22627);
nor U22860 (N_22860,N_22565,N_22634);
nand U22861 (N_22861,N_22557,N_22701);
nand U22862 (N_22862,N_22705,N_22519);
nand U22863 (N_22863,N_22707,N_22739);
and U22864 (N_22864,N_22548,N_22732);
nor U22865 (N_22865,N_22602,N_22681);
nor U22866 (N_22866,N_22655,N_22502);
nand U22867 (N_22867,N_22514,N_22712);
xnor U22868 (N_22868,N_22580,N_22546);
xor U22869 (N_22869,N_22703,N_22650);
xor U22870 (N_22870,N_22618,N_22700);
nand U22871 (N_22871,N_22653,N_22745);
xor U22872 (N_22872,N_22595,N_22696);
or U22873 (N_22873,N_22617,N_22553);
nand U22874 (N_22874,N_22647,N_22741);
nand U22875 (N_22875,N_22561,N_22721);
nor U22876 (N_22876,N_22731,N_22627);
or U22877 (N_22877,N_22548,N_22505);
nor U22878 (N_22878,N_22701,N_22682);
or U22879 (N_22879,N_22686,N_22733);
and U22880 (N_22880,N_22723,N_22742);
and U22881 (N_22881,N_22531,N_22530);
nand U22882 (N_22882,N_22505,N_22704);
xor U22883 (N_22883,N_22536,N_22599);
and U22884 (N_22884,N_22651,N_22536);
nand U22885 (N_22885,N_22520,N_22631);
and U22886 (N_22886,N_22569,N_22702);
nand U22887 (N_22887,N_22692,N_22720);
nor U22888 (N_22888,N_22731,N_22532);
nand U22889 (N_22889,N_22564,N_22506);
and U22890 (N_22890,N_22632,N_22624);
xnor U22891 (N_22891,N_22602,N_22595);
nand U22892 (N_22892,N_22609,N_22730);
nor U22893 (N_22893,N_22573,N_22557);
or U22894 (N_22894,N_22711,N_22600);
nor U22895 (N_22895,N_22566,N_22706);
and U22896 (N_22896,N_22665,N_22650);
or U22897 (N_22897,N_22653,N_22706);
nand U22898 (N_22898,N_22724,N_22534);
nor U22899 (N_22899,N_22545,N_22645);
and U22900 (N_22900,N_22585,N_22541);
or U22901 (N_22901,N_22500,N_22675);
nor U22902 (N_22902,N_22617,N_22581);
and U22903 (N_22903,N_22707,N_22544);
nand U22904 (N_22904,N_22670,N_22523);
nor U22905 (N_22905,N_22537,N_22741);
nand U22906 (N_22906,N_22692,N_22605);
nor U22907 (N_22907,N_22501,N_22568);
nor U22908 (N_22908,N_22639,N_22680);
xor U22909 (N_22909,N_22670,N_22576);
nor U22910 (N_22910,N_22559,N_22609);
nor U22911 (N_22911,N_22567,N_22711);
nand U22912 (N_22912,N_22661,N_22550);
nor U22913 (N_22913,N_22586,N_22721);
nand U22914 (N_22914,N_22510,N_22576);
nand U22915 (N_22915,N_22550,N_22712);
and U22916 (N_22916,N_22563,N_22504);
and U22917 (N_22917,N_22563,N_22737);
or U22918 (N_22918,N_22646,N_22586);
or U22919 (N_22919,N_22544,N_22744);
and U22920 (N_22920,N_22535,N_22719);
nor U22921 (N_22921,N_22649,N_22576);
nand U22922 (N_22922,N_22556,N_22611);
and U22923 (N_22923,N_22699,N_22727);
nor U22924 (N_22924,N_22739,N_22709);
or U22925 (N_22925,N_22505,N_22553);
and U22926 (N_22926,N_22512,N_22723);
xnor U22927 (N_22927,N_22592,N_22601);
and U22928 (N_22928,N_22699,N_22747);
and U22929 (N_22929,N_22667,N_22568);
or U22930 (N_22930,N_22502,N_22728);
or U22931 (N_22931,N_22668,N_22665);
or U22932 (N_22932,N_22577,N_22612);
nor U22933 (N_22933,N_22613,N_22562);
nor U22934 (N_22934,N_22690,N_22546);
nand U22935 (N_22935,N_22734,N_22699);
xor U22936 (N_22936,N_22546,N_22532);
and U22937 (N_22937,N_22716,N_22652);
nand U22938 (N_22938,N_22639,N_22594);
nor U22939 (N_22939,N_22724,N_22718);
nor U22940 (N_22940,N_22634,N_22530);
or U22941 (N_22941,N_22706,N_22657);
or U22942 (N_22942,N_22541,N_22530);
nand U22943 (N_22943,N_22544,N_22547);
xor U22944 (N_22944,N_22506,N_22555);
nor U22945 (N_22945,N_22607,N_22541);
and U22946 (N_22946,N_22728,N_22534);
and U22947 (N_22947,N_22551,N_22685);
nor U22948 (N_22948,N_22744,N_22508);
and U22949 (N_22949,N_22596,N_22650);
and U22950 (N_22950,N_22529,N_22545);
nor U22951 (N_22951,N_22692,N_22740);
nor U22952 (N_22952,N_22515,N_22683);
or U22953 (N_22953,N_22632,N_22582);
or U22954 (N_22954,N_22690,N_22672);
nand U22955 (N_22955,N_22687,N_22544);
or U22956 (N_22956,N_22517,N_22707);
xor U22957 (N_22957,N_22678,N_22554);
nor U22958 (N_22958,N_22674,N_22582);
nor U22959 (N_22959,N_22632,N_22563);
and U22960 (N_22960,N_22687,N_22532);
or U22961 (N_22961,N_22560,N_22562);
and U22962 (N_22962,N_22649,N_22641);
and U22963 (N_22963,N_22621,N_22514);
xor U22964 (N_22964,N_22711,N_22725);
xnor U22965 (N_22965,N_22525,N_22564);
nand U22966 (N_22966,N_22640,N_22505);
or U22967 (N_22967,N_22569,N_22636);
nor U22968 (N_22968,N_22635,N_22516);
nand U22969 (N_22969,N_22687,N_22747);
and U22970 (N_22970,N_22679,N_22600);
and U22971 (N_22971,N_22582,N_22682);
nand U22972 (N_22972,N_22616,N_22699);
nand U22973 (N_22973,N_22689,N_22583);
nand U22974 (N_22974,N_22699,N_22556);
nor U22975 (N_22975,N_22645,N_22732);
nor U22976 (N_22976,N_22681,N_22520);
nand U22977 (N_22977,N_22718,N_22744);
and U22978 (N_22978,N_22635,N_22526);
or U22979 (N_22979,N_22746,N_22524);
and U22980 (N_22980,N_22555,N_22709);
or U22981 (N_22981,N_22711,N_22668);
and U22982 (N_22982,N_22716,N_22542);
nor U22983 (N_22983,N_22561,N_22650);
nand U22984 (N_22984,N_22619,N_22596);
or U22985 (N_22985,N_22541,N_22524);
nand U22986 (N_22986,N_22705,N_22605);
nand U22987 (N_22987,N_22639,N_22634);
nand U22988 (N_22988,N_22728,N_22705);
nand U22989 (N_22989,N_22625,N_22666);
and U22990 (N_22990,N_22717,N_22708);
xor U22991 (N_22991,N_22623,N_22675);
nor U22992 (N_22992,N_22610,N_22686);
or U22993 (N_22993,N_22510,N_22738);
nand U22994 (N_22994,N_22566,N_22699);
nor U22995 (N_22995,N_22683,N_22525);
or U22996 (N_22996,N_22520,N_22722);
or U22997 (N_22997,N_22646,N_22544);
nand U22998 (N_22998,N_22733,N_22617);
nor U22999 (N_22999,N_22646,N_22707);
nor U23000 (N_23000,N_22983,N_22857);
nand U23001 (N_23001,N_22979,N_22831);
or U23002 (N_23002,N_22957,N_22981);
or U23003 (N_23003,N_22952,N_22969);
nand U23004 (N_23004,N_22753,N_22951);
and U23005 (N_23005,N_22846,N_22794);
xor U23006 (N_23006,N_22885,N_22887);
nor U23007 (N_23007,N_22752,N_22907);
xnor U23008 (N_23008,N_22998,N_22903);
and U23009 (N_23009,N_22927,N_22793);
and U23010 (N_23010,N_22762,N_22980);
nor U23011 (N_23011,N_22865,N_22932);
xnor U23012 (N_23012,N_22913,N_22953);
and U23013 (N_23013,N_22766,N_22770);
nand U23014 (N_23014,N_22835,N_22959);
nand U23015 (N_23015,N_22909,N_22806);
nand U23016 (N_23016,N_22904,N_22947);
and U23017 (N_23017,N_22935,N_22996);
or U23018 (N_23018,N_22876,N_22811);
nand U23019 (N_23019,N_22815,N_22813);
or U23020 (N_23020,N_22999,N_22944);
or U23021 (N_23021,N_22829,N_22816);
xor U23022 (N_23022,N_22804,N_22869);
or U23023 (N_23023,N_22905,N_22978);
nand U23024 (N_23024,N_22933,N_22968);
or U23025 (N_23025,N_22859,N_22841);
xor U23026 (N_23026,N_22986,N_22915);
and U23027 (N_23027,N_22967,N_22833);
nand U23028 (N_23028,N_22757,N_22945);
nor U23029 (N_23029,N_22849,N_22760);
nor U23030 (N_23030,N_22761,N_22782);
nor U23031 (N_23031,N_22964,N_22858);
xor U23032 (N_23032,N_22823,N_22792);
xnor U23033 (N_23033,N_22779,N_22754);
and U23034 (N_23034,N_22960,N_22916);
and U23035 (N_23035,N_22897,N_22817);
or U23036 (N_23036,N_22778,N_22809);
nor U23037 (N_23037,N_22862,N_22898);
nor U23038 (N_23038,N_22772,N_22771);
nor U23039 (N_23039,N_22860,N_22901);
nand U23040 (N_23040,N_22873,N_22848);
nand U23041 (N_23041,N_22840,N_22917);
nor U23042 (N_23042,N_22845,N_22821);
nor U23043 (N_23043,N_22977,N_22870);
or U23044 (N_23044,N_22926,N_22796);
nor U23045 (N_23045,N_22874,N_22941);
or U23046 (N_23046,N_22852,N_22801);
nand U23047 (N_23047,N_22994,N_22883);
or U23048 (N_23048,N_22930,N_22958);
or U23049 (N_23049,N_22995,N_22975);
xor U23050 (N_23050,N_22972,N_22925);
or U23051 (N_23051,N_22825,N_22881);
xor U23052 (N_23052,N_22893,N_22919);
nor U23053 (N_23053,N_22934,N_22832);
xnor U23054 (N_23054,N_22877,N_22820);
nand U23055 (N_23055,N_22884,N_22861);
and U23056 (N_23056,N_22764,N_22847);
xnor U23057 (N_23057,N_22868,N_22851);
or U23058 (N_23058,N_22931,N_22973);
and U23059 (N_23059,N_22989,N_22795);
or U23060 (N_23060,N_22949,N_22818);
and U23061 (N_23061,N_22819,N_22908);
or U23062 (N_23062,N_22902,N_22988);
nor U23063 (N_23063,N_22939,N_22943);
or U23064 (N_23064,N_22954,N_22769);
nor U23065 (N_23065,N_22950,N_22910);
or U23066 (N_23066,N_22826,N_22997);
xnor U23067 (N_23067,N_22850,N_22987);
and U23068 (N_23068,N_22843,N_22781);
and U23069 (N_23069,N_22889,N_22777);
and U23070 (N_23070,N_22948,N_22937);
or U23071 (N_23071,N_22992,N_22856);
nand U23072 (N_23072,N_22786,N_22878);
nor U23073 (N_23073,N_22854,N_22991);
nor U23074 (N_23074,N_22837,N_22788);
and U23075 (N_23075,N_22803,N_22797);
or U23076 (N_23076,N_22808,N_22842);
nor U23077 (N_23077,N_22929,N_22767);
and U23078 (N_23078,N_22800,N_22871);
or U23079 (N_23079,N_22789,N_22955);
nor U23080 (N_23080,N_22836,N_22834);
xor U23081 (N_23081,N_22805,N_22890);
nor U23082 (N_23082,N_22882,N_22880);
and U23083 (N_23083,N_22758,N_22923);
nand U23084 (N_23084,N_22921,N_22918);
nand U23085 (N_23085,N_22828,N_22783);
or U23086 (N_23086,N_22751,N_22892);
or U23087 (N_23087,N_22791,N_22824);
or U23088 (N_23088,N_22928,N_22924);
nor U23089 (N_23089,N_22936,N_22961);
nand U23090 (N_23090,N_22785,N_22888);
nor U23091 (N_23091,N_22895,N_22750);
or U23092 (N_23092,N_22814,N_22894);
or U23093 (N_23093,N_22798,N_22938);
nand U23094 (N_23094,N_22993,N_22875);
or U23095 (N_23095,N_22775,N_22946);
or U23096 (N_23096,N_22864,N_22965);
xor U23097 (N_23097,N_22971,N_22812);
nand U23098 (N_23098,N_22914,N_22863);
or U23099 (N_23099,N_22906,N_22759);
nor U23100 (N_23100,N_22976,N_22962);
nand U23101 (N_23101,N_22787,N_22807);
xor U23102 (N_23102,N_22912,N_22956);
nand U23103 (N_23103,N_22940,N_22922);
and U23104 (N_23104,N_22810,N_22822);
or U23105 (N_23105,N_22830,N_22802);
nor U23106 (N_23106,N_22774,N_22867);
or U23107 (N_23107,N_22970,N_22886);
xnor U23108 (N_23108,N_22990,N_22879);
or U23109 (N_23109,N_22984,N_22911);
or U23110 (N_23110,N_22963,N_22966);
or U23111 (N_23111,N_22985,N_22896);
xnor U23112 (N_23112,N_22780,N_22899);
or U23113 (N_23113,N_22920,N_22755);
and U23114 (N_23114,N_22866,N_22900);
nor U23115 (N_23115,N_22891,N_22853);
or U23116 (N_23116,N_22844,N_22763);
nor U23117 (N_23117,N_22765,N_22942);
nand U23118 (N_23118,N_22784,N_22974);
and U23119 (N_23119,N_22790,N_22982);
and U23120 (N_23120,N_22799,N_22776);
and U23121 (N_23121,N_22827,N_22773);
nor U23122 (N_23122,N_22855,N_22838);
nand U23123 (N_23123,N_22768,N_22872);
xor U23124 (N_23124,N_22839,N_22756);
nor U23125 (N_23125,N_22764,N_22752);
nor U23126 (N_23126,N_22804,N_22826);
nor U23127 (N_23127,N_22895,N_22846);
or U23128 (N_23128,N_22785,N_22813);
and U23129 (N_23129,N_22764,N_22769);
or U23130 (N_23130,N_22970,N_22752);
nand U23131 (N_23131,N_22874,N_22814);
or U23132 (N_23132,N_22874,N_22858);
nand U23133 (N_23133,N_22774,N_22947);
nand U23134 (N_23134,N_22988,N_22898);
xnor U23135 (N_23135,N_22852,N_22908);
nor U23136 (N_23136,N_22951,N_22970);
nand U23137 (N_23137,N_22843,N_22916);
nor U23138 (N_23138,N_22876,N_22882);
and U23139 (N_23139,N_22838,N_22874);
xor U23140 (N_23140,N_22753,N_22882);
and U23141 (N_23141,N_22990,N_22937);
nand U23142 (N_23142,N_22784,N_22955);
or U23143 (N_23143,N_22974,N_22963);
nand U23144 (N_23144,N_22837,N_22844);
nand U23145 (N_23145,N_22941,N_22806);
xor U23146 (N_23146,N_22930,N_22994);
nor U23147 (N_23147,N_22911,N_22767);
or U23148 (N_23148,N_22836,N_22891);
and U23149 (N_23149,N_22986,N_22784);
xnor U23150 (N_23150,N_22782,N_22842);
or U23151 (N_23151,N_22947,N_22954);
and U23152 (N_23152,N_22926,N_22753);
nand U23153 (N_23153,N_22864,N_22942);
nor U23154 (N_23154,N_22911,N_22903);
nand U23155 (N_23155,N_22786,N_22765);
xnor U23156 (N_23156,N_22916,N_22958);
or U23157 (N_23157,N_22857,N_22757);
xnor U23158 (N_23158,N_22762,N_22815);
nand U23159 (N_23159,N_22917,N_22930);
and U23160 (N_23160,N_22897,N_22779);
nor U23161 (N_23161,N_22884,N_22818);
and U23162 (N_23162,N_22752,N_22873);
nand U23163 (N_23163,N_22826,N_22844);
or U23164 (N_23164,N_22878,N_22789);
nor U23165 (N_23165,N_22851,N_22903);
or U23166 (N_23166,N_22842,N_22978);
and U23167 (N_23167,N_22963,N_22935);
xnor U23168 (N_23168,N_22890,N_22811);
nor U23169 (N_23169,N_22858,N_22939);
and U23170 (N_23170,N_22775,N_22937);
or U23171 (N_23171,N_22889,N_22860);
nor U23172 (N_23172,N_22802,N_22908);
nand U23173 (N_23173,N_22859,N_22900);
nor U23174 (N_23174,N_22991,N_22966);
nor U23175 (N_23175,N_22782,N_22789);
and U23176 (N_23176,N_22866,N_22975);
xnor U23177 (N_23177,N_22842,N_22824);
nor U23178 (N_23178,N_22883,N_22885);
nand U23179 (N_23179,N_22878,N_22946);
nor U23180 (N_23180,N_22792,N_22958);
nand U23181 (N_23181,N_22813,N_22882);
xor U23182 (N_23182,N_22793,N_22766);
and U23183 (N_23183,N_22957,N_22975);
or U23184 (N_23184,N_22963,N_22759);
nand U23185 (N_23185,N_22824,N_22991);
or U23186 (N_23186,N_22787,N_22781);
nand U23187 (N_23187,N_22793,N_22835);
xnor U23188 (N_23188,N_22931,N_22857);
xor U23189 (N_23189,N_22877,N_22779);
or U23190 (N_23190,N_22996,N_22825);
nand U23191 (N_23191,N_22953,N_22911);
nor U23192 (N_23192,N_22770,N_22803);
nor U23193 (N_23193,N_22926,N_22846);
nand U23194 (N_23194,N_22910,N_22976);
and U23195 (N_23195,N_22886,N_22837);
xor U23196 (N_23196,N_22754,N_22935);
or U23197 (N_23197,N_22983,N_22831);
nand U23198 (N_23198,N_22990,N_22866);
xor U23199 (N_23199,N_22773,N_22768);
nor U23200 (N_23200,N_22772,N_22883);
and U23201 (N_23201,N_22825,N_22945);
and U23202 (N_23202,N_22881,N_22824);
nor U23203 (N_23203,N_22751,N_22932);
or U23204 (N_23204,N_22824,N_22993);
xnor U23205 (N_23205,N_22782,N_22893);
xnor U23206 (N_23206,N_22802,N_22845);
xor U23207 (N_23207,N_22793,N_22991);
nor U23208 (N_23208,N_22799,N_22837);
and U23209 (N_23209,N_22962,N_22830);
and U23210 (N_23210,N_22806,N_22984);
nand U23211 (N_23211,N_22930,N_22750);
nand U23212 (N_23212,N_22940,N_22841);
nor U23213 (N_23213,N_22795,N_22825);
nor U23214 (N_23214,N_22873,N_22766);
nor U23215 (N_23215,N_22954,N_22934);
nand U23216 (N_23216,N_22785,N_22763);
or U23217 (N_23217,N_22894,N_22797);
nand U23218 (N_23218,N_22924,N_22836);
nand U23219 (N_23219,N_22832,N_22801);
xnor U23220 (N_23220,N_22997,N_22892);
nor U23221 (N_23221,N_22810,N_22900);
nor U23222 (N_23222,N_22921,N_22929);
xnor U23223 (N_23223,N_22933,N_22764);
nor U23224 (N_23224,N_22977,N_22757);
xor U23225 (N_23225,N_22916,N_22800);
and U23226 (N_23226,N_22774,N_22994);
and U23227 (N_23227,N_22825,N_22933);
and U23228 (N_23228,N_22883,N_22960);
nand U23229 (N_23229,N_22858,N_22961);
and U23230 (N_23230,N_22828,N_22954);
nand U23231 (N_23231,N_22954,N_22810);
xor U23232 (N_23232,N_22942,N_22796);
and U23233 (N_23233,N_22937,N_22860);
or U23234 (N_23234,N_22892,N_22788);
and U23235 (N_23235,N_22958,N_22863);
nand U23236 (N_23236,N_22764,N_22949);
nor U23237 (N_23237,N_22820,N_22924);
xnor U23238 (N_23238,N_22969,N_22917);
and U23239 (N_23239,N_22905,N_22830);
nor U23240 (N_23240,N_22917,N_22947);
or U23241 (N_23241,N_22914,N_22838);
and U23242 (N_23242,N_22880,N_22845);
nand U23243 (N_23243,N_22941,N_22990);
nor U23244 (N_23244,N_22793,N_22816);
nor U23245 (N_23245,N_22989,N_22771);
nor U23246 (N_23246,N_22772,N_22918);
or U23247 (N_23247,N_22901,N_22962);
and U23248 (N_23248,N_22954,N_22868);
nor U23249 (N_23249,N_22879,N_22919);
and U23250 (N_23250,N_23188,N_23036);
nand U23251 (N_23251,N_23099,N_23000);
and U23252 (N_23252,N_23090,N_23059);
and U23253 (N_23253,N_23084,N_23212);
nand U23254 (N_23254,N_23048,N_23030);
and U23255 (N_23255,N_23160,N_23066);
or U23256 (N_23256,N_23051,N_23010);
or U23257 (N_23257,N_23168,N_23068);
nor U23258 (N_23258,N_23131,N_23045);
nand U23259 (N_23259,N_23189,N_23127);
xnor U23260 (N_23260,N_23028,N_23025);
nor U23261 (N_23261,N_23110,N_23038);
or U23262 (N_23262,N_23141,N_23146);
or U23263 (N_23263,N_23216,N_23184);
nor U23264 (N_23264,N_23083,N_23179);
nand U23265 (N_23265,N_23075,N_23171);
nand U23266 (N_23266,N_23107,N_23016);
and U23267 (N_23267,N_23227,N_23202);
nor U23268 (N_23268,N_23225,N_23012);
nand U23269 (N_23269,N_23133,N_23047);
or U23270 (N_23270,N_23150,N_23101);
or U23271 (N_23271,N_23204,N_23166);
nor U23272 (N_23272,N_23206,N_23040);
nor U23273 (N_23273,N_23191,N_23230);
nand U23274 (N_23274,N_23219,N_23123);
and U23275 (N_23275,N_23244,N_23240);
xor U23276 (N_23276,N_23019,N_23155);
or U23277 (N_23277,N_23170,N_23238);
xor U23278 (N_23278,N_23120,N_23174);
nor U23279 (N_23279,N_23163,N_23178);
or U23280 (N_23280,N_23065,N_23096);
nor U23281 (N_23281,N_23069,N_23079);
nor U23282 (N_23282,N_23094,N_23034);
nor U23283 (N_23283,N_23004,N_23176);
or U23284 (N_23284,N_23013,N_23035);
nand U23285 (N_23285,N_23195,N_23249);
and U23286 (N_23286,N_23237,N_23167);
and U23287 (N_23287,N_23067,N_23214);
nand U23288 (N_23288,N_23073,N_23064);
and U23289 (N_23289,N_23095,N_23236);
or U23290 (N_23290,N_23104,N_23109);
nand U23291 (N_23291,N_23217,N_23115);
nand U23292 (N_23292,N_23147,N_23097);
or U23293 (N_23293,N_23126,N_23011);
nand U23294 (N_23294,N_23226,N_23239);
or U23295 (N_23295,N_23041,N_23149);
nor U23296 (N_23296,N_23112,N_23006);
or U23297 (N_23297,N_23161,N_23005);
nand U23298 (N_23298,N_23098,N_23119);
xor U23299 (N_23299,N_23210,N_23007);
or U23300 (N_23300,N_23091,N_23208);
nor U23301 (N_23301,N_23049,N_23046);
or U23302 (N_23302,N_23029,N_23232);
or U23303 (N_23303,N_23039,N_23231);
and U23304 (N_23304,N_23224,N_23003);
and U23305 (N_23305,N_23196,N_23203);
nor U23306 (N_23306,N_23100,N_23173);
or U23307 (N_23307,N_23023,N_23218);
nor U23308 (N_23308,N_23116,N_23205);
or U23309 (N_23309,N_23086,N_23021);
nor U23310 (N_23310,N_23114,N_23072);
nand U23311 (N_23311,N_23229,N_23001);
nor U23312 (N_23312,N_23140,N_23220);
nor U23313 (N_23313,N_23103,N_23213);
and U23314 (N_23314,N_23077,N_23071);
and U23315 (N_23315,N_23130,N_23246);
or U23316 (N_23316,N_23145,N_23093);
or U23317 (N_23317,N_23061,N_23033);
nand U23318 (N_23318,N_23136,N_23024);
or U23319 (N_23319,N_23215,N_23043);
or U23320 (N_23320,N_23234,N_23143);
and U23321 (N_23321,N_23125,N_23128);
xor U23322 (N_23322,N_23026,N_23076);
nand U23323 (N_23323,N_23192,N_23135);
nand U23324 (N_23324,N_23017,N_23177);
or U23325 (N_23325,N_23020,N_23154);
or U23326 (N_23326,N_23018,N_23053);
xnor U23327 (N_23327,N_23037,N_23002);
and U23328 (N_23328,N_23193,N_23241);
and U23329 (N_23329,N_23102,N_23106);
and U23330 (N_23330,N_23118,N_23198);
nor U23331 (N_23331,N_23031,N_23222);
and U23332 (N_23332,N_23144,N_23008);
nor U23333 (N_23333,N_23138,N_23165);
nor U23334 (N_23334,N_23044,N_23129);
nand U23335 (N_23335,N_23242,N_23190);
and U23336 (N_23336,N_23207,N_23124);
or U23337 (N_23337,N_23159,N_23054);
nand U23338 (N_23338,N_23153,N_23183);
or U23339 (N_23339,N_23164,N_23182);
and U23340 (N_23340,N_23134,N_23108);
and U23341 (N_23341,N_23181,N_23089);
nor U23342 (N_23342,N_23172,N_23200);
xnor U23343 (N_23343,N_23022,N_23169);
nand U23344 (N_23344,N_23080,N_23209);
or U23345 (N_23345,N_23087,N_23032);
or U23346 (N_23346,N_23156,N_23199);
or U23347 (N_23347,N_23223,N_23132);
and U23348 (N_23348,N_23197,N_23070);
nor U23349 (N_23349,N_23148,N_23085);
nand U23350 (N_23350,N_23247,N_23063);
nand U23351 (N_23351,N_23186,N_23122);
and U23352 (N_23352,N_23175,N_23088);
nand U23353 (N_23353,N_23014,N_23078);
and U23354 (N_23354,N_23187,N_23092);
nand U23355 (N_23355,N_23152,N_23009);
and U23356 (N_23356,N_23180,N_23042);
nor U23357 (N_23357,N_23062,N_23248);
and U23358 (N_23358,N_23050,N_23060);
nor U23359 (N_23359,N_23105,N_23233);
and U23360 (N_23360,N_23058,N_23157);
and U23361 (N_23361,N_23211,N_23082);
xnor U23362 (N_23362,N_23245,N_23243);
and U23363 (N_23363,N_23057,N_23201);
and U23364 (N_23364,N_23228,N_23151);
or U23365 (N_23365,N_23185,N_23056);
nor U23366 (N_23366,N_23121,N_23158);
and U23367 (N_23367,N_23111,N_23055);
nand U23368 (N_23368,N_23074,N_23139);
and U23369 (N_23369,N_23015,N_23137);
or U23370 (N_23370,N_23027,N_23162);
nand U23371 (N_23371,N_23052,N_23142);
nand U23372 (N_23372,N_23081,N_23117);
nor U23373 (N_23373,N_23235,N_23113);
nand U23374 (N_23374,N_23221,N_23194);
nand U23375 (N_23375,N_23083,N_23226);
nor U23376 (N_23376,N_23087,N_23043);
nand U23377 (N_23377,N_23072,N_23101);
and U23378 (N_23378,N_23028,N_23160);
xnor U23379 (N_23379,N_23039,N_23042);
nand U23380 (N_23380,N_23012,N_23114);
xor U23381 (N_23381,N_23232,N_23044);
xnor U23382 (N_23382,N_23238,N_23171);
xnor U23383 (N_23383,N_23042,N_23068);
nand U23384 (N_23384,N_23106,N_23088);
and U23385 (N_23385,N_23245,N_23063);
nand U23386 (N_23386,N_23057,N_23078);
xor U23387 (N_23387,N_23011,N_23155);
nand U23388 (N_23388,N_23095,N_23223);
and U23389 (N_23389,N_23077,N_23156);
nand U23390 (N_23390,N_23139,N_23211);
and U23391 (N_23391,N_23220,N_23240);
nand U23392 (N_23392,N_23011,N_23081);
nand U23393 (N_23393,N_23203,N_23170);
nor U23394 (N_23394,N_23033,N_23050);
or U23395 (N_23395,N_23137,N_23126);
nand U23396 (N_23396,N_23116,N_23004);
nor U23397 (N_23397,N_23101,N_23130);
or U23398 (N_23398,N_23174,N_23215);
nand U23399 (N_23399,N_23182,N_23114);
nand U23400 (N_23400,N_23027,N_23024);
nand U23401 (N_23401,N_23185,N_23039);
nor U23402 (N_23402,N_23099,N_23123);
nand U23403 (N_23403,N_23088,N_23015);
and U23404 (N_23404,N_23142,N_23069);
and U23405 (N_23405,N_23205,N_23005);
or U23406 (N_23406,N_23071,N_23079);
nor U23407 (N_23407,N_23231,N_23113);
nor U23408 (N_23408,N_23122,N_23042);
nor U23409 (N_23409,N_23169,N_23171);
and U23410 (N_23410,N_23099,N_23183);
nand U23411 (N_23411,N_23149,N_23245);
nor U23412 (N_23412,N_23155,N_23013);
and U23413 (N_23413,N_23073,N_23213);
nand U23414 (N_23414,N_23079,N_23085);
xnor U23415 (N_23415,N_23249,N_23209);
xnor U23416 (N_23416,N_23014,N_23041);
and U23417 (N_23417,N_23066,N_23142);
xor U23418 (N_23418,N_23222,N_23242);
or U23419 (N_23419,N_23241,N_23115);
nand U23420 (N_23420,N_23166,N_23039);
nand U23421 (N_23421,N_23210,N_23102);
nor U23422 (N_23422,N_23139,N_23087);
or U23423 (N_23423,N_23140,N_23247);
nor U23424 (N_23424,N_23163,N_23093);
nand U23425 (N_23425,N_23178,N_23220);
nor U23426 (N_23426,N_23057,N_23218);
and U23427 (N_23427,N_23115,N_23100);
nand U23428 (N_23428,N_23156,N_23074);
nand U23429 (N_23429,N_23069,N_23201);
or U23430 (N_23430,N_23021,N_23046);
and U23431 (N_23431,N_23016,N_23138);
nand U23432 (N_23432,N_23018,N_23098);
nor U23433 (N_23433,N_23002,N_23022);
and U23434 (N_23434,N_23223,N_23183);
nand U23435 (N_23435,N_23114,N_23191);
nor U23436 (N_23436,N_23240,N_23241);
nor U23437 (N_23437,N_23216,N_23043);
nand U23438 (N_23438,N_23168,N_23127);
nor U23439 (N_23439,N_23239,N_23049);
or U23440 (N_23440,N_23157,N_23156);
nor U23441 (N_23441,N_23093,N_23026);
nor U23442 (N_23442,N_23208,N_23114);
or U23443 (N_23443,N_23137,N_23089);
or U23444 (N_23444,N_23012,N_23193);
nand U23445 (N_23445,N_23060,N_23059);
nand U23446 (N_23446,N_23238,N_23126);
xor U23447 (N_23447,N_23150,N_23160);
or U23448 (N_23448,N_23201,N_23033);
nor U23449 (N_23449,N_23021,N_23078);
or U23450 (N_23450,N_23116,N_23171);
or U23451 (N_23451,N_23223,N_23242);
or U23452 (N_23452,N_23159,N_23239);
nor U23453 (N_23453,N_23215,N_23145);
or U23454 (N_23454,N_23159,N_23198);
nor U23455 (N_23455,N_23190,N_23196);
and U23456 (N_23456,N_23103,N_23207);
and U23457 (N_23457,N_23224,N_23128);
and U23458 (N_23458,N_23059,N_23151);
nand U23459 (N_23459,N_23073,N_23241);
nor U23460 (N_23460,N_23092,N_23045);
nand U23461 (N_23461,N_23163,N_23046);
nand U23462 (N_23462,N_23100,N_23022);
nor U23463 (N_23463,N_23005,N_23054);
nand U23464 (N_23464,N_23023,N_23185);
nor U23465 (N_23465,N_23168,N_23138);
nand U23466 (N_23466,N_23239,N_23119);
or U23467 (N_23467,N_23077,N_23235);
xnor U23468 (N_23468,N_23078,N_23097);
xor U23469 (N_23469,N_23205,N_23057);
nor U23470 (N_23470,N_23221,N_23105);
nor U23471 (N_23471,N_23128,N_23065);
nor U23472 (N_23472,N_23002,N_23215);
and U23473 (N_23473,N_23143,N_23090);
or U23474 (N_23474,N_23187,N_23185);
or U23475 (N_23475,N_23005,N_23045);
nand U23476 (N_23476,N_23028,N_23049);
nand U23477 (N_23477,N_23091,N_23083);
xor U23478 (N_23478,N_23014,N_23209);
nor U23479 (N_23479,N_23189,N_23008);
nand U23480 (N_23480,N_23164,N_23065);
nand U23481 (N_23481,N_23007,N_23013);
nor U23482 (N_23482,N_23201,N_23090);
and U23483 (N_23483,N_23073,N_23174);
and U23484 (N_23484,N_23182,N_23107);
nor U23485 (N_23485,N_23229,N_23171);
nor U23486 (N_23486,N_23036,N_23100);
nand U23487 (N_23487,N_23079,N_23022);
and U23488 (N_23488,N_23145,N_23005);
nor U23489 (N_23489,N_23060,N_23171);
and U23490 (N_23490,N_23074,N_23173);
or U23491 (N_23491,N_23109,N_23169);
nor U23492 (N_23492,N_23019,N_23100);
nor U23493 (N_23493,N_23074,N_23123);
or U23494 (N_23494,N_23181,N_23073);
nand U23495 (N_23495,N_23201,N_23158);
nor U23496 (N_23496,N_23182,N_23040);
nand U23497 (N_23497,N_23224,N_23181);
xnor U23498 (N_23498,N_23127,N_23239);
nor U23499 (N_23499,N_23228,N_23013);
nor U23500 (N_23500,N_23305,N_23391);
and U23501 (N_23501,N_23415,N_23311);
nand U23502 (N_23502,N_23250,N_23326);
and U23503 (N_23503,N_23447,N_23404);
nand U23504 (N_23504,N_23303,N_23372);
nand U23505 (N_23505,N_23416,N_23364);
nand U23506 (N_23506,N_23429,N_23499);
nor U23507 (N_23507,N_23370,N_23251);
and U23508 (N_23508,N_23304,N_23266);
and U23509 (N_23509,N_23320,N_23402);
nand U23510 (N_23510,N_23354,N_23388);
or U23511 (N_23511,N_23452,N_23287);
xnor U23512 (N_23512,N_23394,N_23437);
and U23513 (N_23513,N_23414,N_23397);
xor U23514 (N_23514,N_23475,N_23264);
nor U23515 (N_23515,N_23374,N_23342);
and U23516 (N_23516,N_23408,N_23260);
and U23517 (N_23517,N_23435,N_23276);
nor U23518 (N_23518,N_23403,N_23459);
or U23519 (N_23519,N_23420,N_23498);
xnor U23520 (N_23520,N_23300,N_23446);
xnor U23521 (N_23521,N_23261,N_23466);
xor U23522 (N_23522,N_23375,N_23280);
nor U23523 (N_23523,N_23302,N_23453);
nand U23524 (N_23524,N_23484,N_23357);
xnor U23525 (N_23525,N_23497,N_23360);
and U23526 (N_23526,N_23263,N_23451);
xor U23527 (N_23527,N_23379,N_23477);
nand U23528 (N_23528,N_23438,N_23335);
and U23529 (N_23529,N_23361,N_23398);
or U23530 (N_23530,N_23426,N_23461);
nor U23531 (N_23531,N_23473,N_23355);
or U23532 (N_23532,N_23285,N_23295);
nand U23533 (N_23533,N_23373,N_23298);
and U23534 (N_23534,N_23389,N_23327);
and U23535 (N_23535,N_23490,N_23347);
or U23536 (N_23536,N_23259,N_23424);
or U23537 (N_23537,N_23339,N_23328);
nand U23538 (N_23538,N_23319,N_23277);
nand U23539 (N_23539,N_23377,N_23376);
nor U23540 (N_23540,N_23367,N_23419);
and U23541 (N_23541,N_23381,N_23468);
nor U23542 (N_23542,N_23455,N_23428);
or U23543 (N_23543,N_23333,N_23488);
and U23544 (N_23544,N_23380,N_23464);
and U23545 (N_23545,N_23341,N_23332);
and U23546 (N_23546,N_23393,N_23293);
and U23547 (N_23547,N_23431,N_23443);
and U23548 (N_23548,N_23353,N_23427);
nand U23549 (N_23549,N_23337,N_23485);
xor U23550 (N_23550,N_23494,N_23495);
or U23551 (N_23551,N_23396,N_23281);
or U23552 (N_23552,N_23423,N_23299);
nand U23553 (N_23553,N_23318,N_23313);
nand U23554 (N_23554,N_23352,N_23349);
nor U23555 (N_23555,N_23493,N_23297);
or U23556 (N_23556,N_23254,N_23314);
and U23557 (N_23557,N_23400,N_23253);
and U23558 (N_23558,N_23366,N_23385);
xor U23559 (N_23559,N_23257,N_23309);
and U23560 (N_23560,N_23476,N_23390);
nand U23561 (N_23561,N_23441,N_23343);
or U23562 (N_23562,N_23480,N_23255);
nor U23563 (N_23563,N_23483,N_23369);
xor U23564 (N_23564,N_23282,N_23418);
and U23565 (N_23565,N_23344,N_23417);
nor U23566 (N_23566,N_23334,N_23256);
nand U23567 (N_23567,N_23413,N_23262);
or U23568 (N_23568,N_23383,N_23442);
or U23569 (N_23569,N_23368,N_23445);
nor U23570 (N_23570,N_23481,N_23284);
xor U23571 (N_23571,N_23486,N_23283);
nand U23572 (N_23572,N_23350,N_23411);
and U23573 (N_23573,N_23382,N_23439);
nor U23574 (N_23574,N_23306,N_23492);
nor U23575 (N_23575,N_23315,N_23422);
nand U23576 (N_23576,N_23338,N_23340);
or U23577 (N_23577,N_23433,N_23288);
and U23578 (N_23578,N_23491,N_23478);
nor U23579 (N_23579,N_23440,N_23258);
and U23580 (N_23580,N_23265,N_23407);
nand U23581 (N_23581,N_23467,N_23378);
or U23582 (N_23582,N_23336,N_23412);
or U23583 (N_23583,N_23275,N_23454);
and U23584 (N_23584,N_23425,N_23365);
nand U23585 (N_23585,N_23312,N_23330);
and U23586 (N_23586,N_23474,N_23325);
and U23587 (N_23587,N_23324,N_23308);
and U23588 (N_23588,N_23270,N_23289);
and U23589 (N_23589,N_23321,N_23401);
xnor U23590 (N_23590,N_23363,N_23267);
and U23591 (N_23591,N_23462,N_23448);
or U23592 (N_23592,N_23430,N_23409);
nand U23593 (N_23593,N_23406,N_23436);
nor U23594 (N_23594,N_23371,N_23399);
or U23595 (N_23595,N_23449,N_23405);
nand U23596 (N_23596,N_23317,N_23358);
or U23597 (N_23597,N_23482,N_23450);
and U23598 (N_23598,N_23434,N_23487);
and U23599 (N_23599,N_23286,N_23322);
nor U23600 (N_23600,N_23463,N_23274);
and U23601 (N_23601,N_23296,N_23294);
nand U23602 (N_23602,N_23279,N_23331);
and U23603 (N_23603,N_23465,N_23395);
nand U23604 (N_23604,N_23301,N_23346);
nor U23605 (N_23605,N_23348,N_23291);
nor U23606 (N_23606,N_23307,N_23496);
xor U23607 (N_23607,N_23269,N_23460);
or U23608 (N_23608,N_23386,N_23356);
or U23609 (N_23609,N_23273,N_23469);
or U23610 (N_23610,N_23471,N_23479);
nand U23611 (N_23611,N_23456,N_23329);
and U23612 (N_23612,N_23410,N_23457);
or U23613 (N_23613,N_23271,N_23489);
nand U23614 (N_23614,N_23316,N_23387);
or U23615 (N_23615,N_23384,N_23323);
nand U23616 (N_23616,N_23392,N_23252);
nand U23617 (N_23617,N_23470,N_23421);
or U23618 (N_23618,N_23290,N_23359);
and U23619 (N_23619,N_23351,N_23310);
and U23620 (N_23620,N_23292,N_23345);
or U23621 (N_23621,N_23458,N_23472);
nor U23622 (N_23622,N_23268,N_23432);
and U23623 (N_23623,N_23278,N_23444);
nand U23624 (N_23624,N_23272,N_23362);
xnor U23625 (N_23625,N_23425,N_23399);
nand U23626 (N_23626,N_23425,N_23378);
xnor U23627 (N_23627,N_23363,N_23347);
xnor U23628 (N_23628,N_23333,N_23273);
or U23629 (N_23629,N_23496,N_23292);
and U23630 (N_23630,N_23488,N_23444);
and U23631 (N_23631,N_23340,N_23396);
nand U23632 (N_23632,N_23424,N_23342);
xor U23633 (N_23633,N_23372,N_23352);
or U23634 (N_23634,N_23493,N_23320);
nor U23635 (N_23635,N_23341,N_23306);
or U23636 (N_23636,N_23438,N_23420);
or U23637 (N_23637,N_23369,N_23432);
nand U23638 (N_23638,N_23388,N_23475);
xnor U23639 (N_23639,N_23379,N_23498);
nor U23640 (N_23640,N_23358,N_23472);
or U23641 (N_23641,N_23333,N_23316);
nand U23642 (N_23642,N_23263,N_23376);
nor U23643 (N_23643,N_23472,N_23478);
or U23644 (N_23644,N_23391,N_23279);
nor U23645 (N_23645,N_23354,N_23251);
nor U23646 (N_23646,N_23474,N_23400);
or U23647 (N_23647,N_23278,N_23422);
and U23648 (N_23648,N_23375,N_23483);
or U23649 (N_23649,N_23449,N_23387);
nand U23650 (N_23650,N_23261,N_23320);
nand U23651 (N_23651,N_23333,N_23321);
nor U23652 (N_23652,N_23324,N_23253);
or U23653 (N_23653,N_23456,N_23290);
or U23654 (N_23654,N_23457,N_23437);
and U23655 (N_23655,N_23366,N_23480);
nor U23656 (N_23656,N_23474,N_23314);
or U23657 (N_23657,N_23461,N_23470);
nand U23658 (N_23658,N_23413,N_23334);
or U23659 (N_23659,N_23366,N_23267);
or U23660 (N_23660,N_23274,N_23435);
nand U23661 (N_23661,N_23289,N_23351);
and U23662 (N_23662,N_23310,N_23291);
xor U23663 (N_23663,N_23415,N_23327);
xnor U23664 (N_23664,N_23404,N_23468);
and U23665 (N_23665,N_23387,N_23384);
xor U23666 (N_23666,N_23360,N_23375);
or U23667 (N_23667,N_23270,N_23262);
xnor U23668 (N_23668,N_23497,N_23452);
or U23669 (N_23669,N_23295,N_23424);
nand U23670 (N_23670,N_23384,N_23487);
and U23671 (N_23671,N_23403,N_23303);
nand U23672 (N_23672,N_23284,N_23409);
nand U23673 (N_23673,N_23421,N_23422);
and U23674 (N_23674,N_23466,N_23472);
xor U23675 (N_23675,N_23300,N_23438);
nor U23676 (N_23676,N_23263,N_23334);
or U23677 (N_23677,N_23420,N_23497);
and U23678 (N_23678,N_23279,N_23374);
or U23679 (N_23679,N_23365,N_23423);
and U23680 (N_23680,N_23492,N_23445);
nand U23681 (N_23681,N_23362,N_23397);
nor U23682 (N_23682,N_23434,N_23360);
or U23683 (N_23683,N_23401,N_23357);
or U23684 (N_23684,N_23483,N_23411);
xor U23685 (N_23685,N_23268,N_23446);
nor U23686 (N_23686,N_23393,N_23397);
and U23687 (N_23687,N_23262,N_23444);
and U23688 (N_23688,N_23293,N_23344);
or U23689 (N_23689,N_23326,N_23348);
or U23690 (N_23690,N_23309,N_23322);
nor U23691 (N_23691,N_23259,N_23375);
nand U23692 (N_23692,N_23372,N_23467);
and U23693 (N_23693,N_23311,N_23260);
nor U23694 (N_23694,N_23466,N_23339);
nor U23695 (N_23695,N_23457,N_23443);
nand U23696 (N_23696,N_23328,N_23268);
or U23697 (N_23697,N_23253,N_23317);
nand U23698 (N_23698,N_23470,N_23484);
or U23699 (N_23699,N_23261,N_23331);
nand U23700 (N_23700,N_23316,N_23262);
or U23701 (N_23701,N_23335,N_23303);
nand U23702 (N_23702,N_23497,N_23473);
nor U23703 (N_23703,N_23288,N_23303);
or U23704 (N_23704,N_23263,N_23495);
or U23705 (N_23705,N_23496,N_23321);
or U23706 (N_23706,N_23251,N_23294);
and U23707 (N_23707,N_23292,N_23434);
or U23708 (N_23708,N_23392,N_23402);
xor U23709 (N_23709,N_23300,N_23344);
xor U23710 (N_23710,N_23473,N_23377);
xor U23711 (N_23711,N_23260,N_23265);
nor U23712 (N_23712,N_23317,N_23271);
or U23713 (N_23713,N_23353,N_23417);
nand U23714 (N_23714,N_23283,N_23259);
nand U23715 (N_23715,N_23301,N_23484);
nor U23716 (N_23716,N_23473,N_23427);
or U23717 (N_23717,N_23316,N_23435);
nand U23718 (N_23718,N_23253,N_23345);
and U23719 (N_23719,N_23329,N_23280);
and U23720 (N_23720,N_23371,N_23372);
nor U23721 (N_23721,N_23336,N_23268);
xnor U23722 (N_23722,N_23319,N_23265);
xor U23723 (N_23723,N_23455,N_23361);
and U23724 (N_23724,N_23278,N_23399);
nor U23725 (N_23725,N_23487,N_23388);
and U23726 (N_23726,N_23458,N_23390);
or U23727 (N_23727,N_23279,N_23493);
and U23728 (N_23728,N_23484,N_23344);
or U23729 (N_23729,N_23441,N_23305);
or U23730 (N_23730,N_23446,N_23292);
or U23731 (N_23731,N_23318,N_23449);
nor U23732 (N_23732,N_23444,N_23371);
or U23733 (N_23733,N_23437,N_23290);
nor U23734 (N_23734,N_23315,N_23329);
nor U23735 (N_23735,N_23445,N_23365);
and U23736 (N_23736,N_23374,N_23459);
nand U23737 (N_23737,N_23279,N_23262);
xor U23738 (N_23738,N_23419,N_23449);
xor U23739 (N_23739,N_23457,N_23419);
and U23740 (N_23740,N_23347,N_23498);
nand U23741 (N_23741,N_23351,N_23265);
nand U23742 (N_23742,N_23321,N_23379);
nand U23743 (N_23743,N_23315,N_23452);
nand U23744 (N_23744,N_23326,N_23410);
nor U23745 (N_23745,N_23324,N_23264);
and U23746 (N_23746,N_23406,N_23407);
and U23747 (N_23747,N_23398,N_23444);
and U23748 (N_23748,N_23266,N_23404);
and U23749 (N_23749,N_23318,N_23421);
nor U23750 (N_23750,N_23680,N_23518);
nand U23751 (N_23751,N_23587,N_23524);
and U23752 (N_23752,N_23519,N_23503);
xor U23753 (N_23753,N_23728,N_23513);
nor U23754 (N_23754,N_23722,N_23535);
nand U23755 (N_23755,N_23664,N_23707);
or U23756 (N_23756,N_23739,N_23696);
nor U23757 (N_23757,N_23539,N_23555);
or U23758 (N_23758,N_23700,N_23536);
xnor U23759 (N_23759,N_23584,N_23640);
or U23760 (N_23760,N_23588,N_23529);
and U23761 (N_23761,N_23515,N_23599);
or U23762 (N_23762,N_23646,N_23512);
nand U23763 (N_23763,N_23718,N_23694);
and U23764 (N_23764,N_23733,N_23674);
xnor U23765 (N_23765,N_23604,N_23569);
nand U23766 (N_23766,N_23730,N_23721);
and U23767 (N_23767,N_23617,N_23670);
nor U23768 (N_23768,N_23608,N_23528);
xnor U23769 (N_23769,N_23594,N_23595);
nand U23770 (N_23770,N_23724,N_23574);
or U23771 (N_23771,N_23625,N_23601);
nand U23772 (N_23772,N_23687,N_23649);
nor U23773 (N_23773,N_23633,N_23705);
xor U23774 (N_23774,N_23671,N_23603);
nor U23775 (N_23775,N_23740,N_23581);
nand U23776 (N_23776,N_23702,N_23712);
nand U23777 (N_23777,N_23666,N_23634);
and U23778 (N_23778,N_23719,N_23637);
and U23779 (N_23779,N_23623,N_23660);
and U23780 (N_23780,N_23532,N_23662);
and U23781 (N_23781,N_23520,N_23709);
or U23782 (N_23782,N_23648,N_23554);
or U23783 (N_23783,N_23745,N_23641);
and U23784 (N_23784,N_23579,N_23575);
and U23785 (N_23785,N_23685,N_23639);
and U23786 (N_23786,N_23615,N_23585);
nand U23787 (N_23787,N_23635,N_23600);
nor U23788 (N_23788,N_23727,N_23668);
nand U23789 (N_23789,N_23573,N_23619);
and U23790 (N_23790,N_23563,N_23720);
or U23791 (N_23791,N_23507,N_23571);
and U23792 (N_23792,N_23557,N_23568);
or U23793 (N_23793,N_23653,N_23676);
nand U23794 (N_23794,N_23693,N_23586);
and U23795 (N_23795,N_23688,N_23683);
nor U23796 (N_23796,N_23741,N_23642);
and U23797 (N_23797,N_23697,N_23692);
and U23798 (N_23798,N_23606,N_23643);
or U23799 (N_23799,N_23716,N_23531);
and U23800 (N_23800,N_23734,N_23678);
and U23801 (N_23801,N_23597,N_23703);
xnor U23802 (N_23802,N_23592,N_23713);
nor U23803 (N_23803,N_23548,N_23723);
nor U23804 (N_23804,N_23704,N_23570);
nand U23805 (N_23805,N_23549,N_23744);
nor U23806 (N_23806,N_23542,N_23647);
xnor U23807 (N_23807,N_23673,N_23725);
nor U23808 (N_23808,N_23747,N_23508);
and U23809 (N_23809,N_23552,N_23657);
and U23810 (N_23810,N_23686,N_23636);
nand U23811 (N_23811,N_23627,N_23746);
nor U23812 (N_23812,N_23525,N_23620);
nand U23813 (N_23813,N_23501,N_23714);
nand U23814 (N_23814,N_23644,N_23630);
nor U23815 (N_23815,N_23749,N_23726);
and U23816 (N_23816,N_23511,N_23577);
nand U23817 (N_23817,N_23596,N_23613);
or U23818 (N_23818,N_23560,N_23624);
and U23819 (N_23819,N_23504,N_23576);
and U23820 (N_23820,N_23682,N_23706);
and U23821 (N_23821,N_23699,N_23609);
or U23822 (N_23822,N_23616,N_23559);
or U23823 (N_23823,N_23663,N_23654);
nand U23824 (N_23824,N_23530,N_23611);
nor U23825 (N_23825,N_23672,N_23534);
nor U23826 (N_23826,N_23506,N_23543);
and U23827 (N_23827,N_23517,N_23658);
xnor U23828 (N_23828,N_23545,N_23553);
xor U23829 (N_23829,N_23593,N_23677);
nor U23830 (N_23830,N_23684,N_23516);
and U23831 (N_23831,N_23665,N_23522);
nor U23832 (N_23832,N_23629,N_23566);
nand U23833 (N_23833,N_23655,N_23500);
xor U23834 (N_23834,N_23510,N_23731);
or U23835 (N_23835,N_23523,N_23729);
or U23836 (N_23836,N_23578,N_23590);
xor U23837 (N_23837,N_23614,N_23556);
nand U23838 (N_23838,N_23743,N_23715);
nand U23839 (N_23839,N_23567,N_23622);
nor U23840 (N_23840,N_23711,N_23689);
nor U23841 (N_23841,N_23580,N_23502);
nand U23842 (N_23842,N_23695,N_23652);
xor U23843 (N_23843,N_23610,N_23583);
nand U23844 (N_23844,N_23565,N_23618);
nor U23845 (N_23845,N_23607,N_23669);
and U23846 (N_23846,N_23572,N_23717);
xor U23847 (N_23847,N_23732,N_23667);
nand U23848 (N_23848,N_23538,N_23544);
nand U23849 (N_23849,N_23701,N_23748);
or U23850 (N_23850,N_23564,N_23736);
or U23851 (N_23851,N_23679,N_23632);
nor U23852 (N_23852,N_23675,N_23561);
nand U23853 (N_23853,N_23735,N_23650);
nand U23854 (N_23854,N_23537,N_23526);
nor U23855 (N_23855,N_23605,N_23690);
nand U23856 (N_23856,N_23742,N_23626);
and U23857 (N_23857,N_23708,N_23546);
or U23858 (N_23858,N_23638,N_23505);
or U23859 (N_23859,N_23551,N_23533);
nand U23860 (N_23860,N_23550,N_23541);
nor U23861 (N_23861,N_23656,N_23547);
and U23862 (N_23862,N_23602,N_23691);
and U23863 (N_23863,N_23589,N_23738);
and U23864 (N_23864,N_23591,N_23645);
or U23865 (N_23865,N_23540,N_23598);
nor U23866 (N_23866,N_23681,N_23582);
or U23867 (N_23867,N_23710,N_23621);
or U23868 (N_23868,N_23651,N_23527);
or U23869 (N_23869,N_23698,N_23562);
nor U23870 (N_23870,N_23514,N_23521);
or U23871 (N_23871,N_23659,N_23737);
nand U23872 (N_23872,N_23509,N_23631);
and U23873 (N_23873,N_23558,N_23628);
and U23874 (N_23874,N_23612,N_23661);
or U23875 (N_23875,N_23523,N_23580);
nor U23876 (N_23876,N_23552,N_23646);
or U23877 (N_23877,N_23680,N_23517);
nand U23878 (N_23878,N_23739,N_23737);
nor U23879 (N_23879,N_23618,N_23652);
xor U23880 (N_23880,N_23578,N_23559);
and U23881 (N_23881,N_23693,N_23712);
or U23882 (N_23882,N_23515,N_23695);
xnor U23883 (N_23883,N_23533,N_23549);
and U23884 (N_23884,N_23600,N_23602);
and U23885 (N_23885,N_23525,N_23611);
nor U23886 (N_23886,N_23519,N_23574);
nand U23887 (N_23887,N_23724,N_23697);
or U23888 (N_23888,N_23724,N_23735);
or U23889 (N_23889,N_23658,N_23531);
xor U23890 (N_23890,N_23589,N_23654);
nand U23891 (N_23891,N_23714,N_23741);
nand U23892 (N_23892,N_23706,N_23516);
nand U23893 (N_23893,N_23635,N_23748);
nor U23894 (N_23894,N_23589,N_23573);
nand U23895 (N_23895,N_23600,N_23611);
nor U23896 (N_23896,N_23627,N_23530);
nand U23897 (N_23897,N_23527,N_23621);
nand U23898 (N_23898,N_23546,N_23609);
or U23899 (N_23899,N_23516,N_23542);
nor U23900 (N_23900,N_23565,N_23634);
nor U23901 (N_23901,N_23526,N_23543);
nand U23902 (N_23902,N_23687,N_23721);
and U23903 (N_23903,N_23734,N_23629);
and U23904 (N_23904,N_23716,N_23602);
nand U23905 (N_23905,N_23722,N_23612);
or U23906 (N_23906,N_23710,N_23669);
nand U23907 (N_23907,N_23629,N_23720);
and U23908 (N_23908,N_23717,N_23716);
nand U23909 (N_23909,N_23549,N_23616);
nor U23910 (N_23910,N_23631,N_23681);
and U23911 (N_23911,N_23566,N_23721);
nor U23912 (N_23912,N_23682,N_23597);
and U23913 (N_23913,N_23622,N_23585);
and U23914 (N_23914,N_23669,N_23651);
nor U23915 (N_23915,N_23504,N_23546);
nor U23916 (N_23916,N_23545,N_23550);
and U23917 (N_23917,N_23678,N_23525);
and U23918 (N_23918,N_23688,N_23511);
and U23919 (N_23919,N_23665,N_23543);
and U23920 (N_23920,N_23695,N_23546);
nor U23921 (N_23921,N_23630,N_23578);
nand U23922 (N_23922,N_23648,N_23553);
xor U23923 (N_23923,N_23683,N_23505);
nand U23924 (N_23924,N_23722,N_23631);
xor U23925 (N_23925,N_23745,N_23554);
nand U23926 (N_23926,N_23589,N_23742);
or U23927 (N_23927,N_23502,N_23718);
or U23928 (N_23928,N_23622,N_23661);
and U23929 (N_23929,N_23546,N_23736);
nor U23930 (N_23930,N_23545,N_23514);
and U23931 (N_23931,N_23543,N_23640);
nor U23932 (N_23932,N_23583,N_23525);
xnor U23933 (N_23933,N_23518,N_23594);
and U23934 (N_23934,N_23748,N_23504);
nor U23935 (N_23935,N_23577,N_23659);
and U23936 (N_23936,N_23530,N_23683);
nand U23937 (N_23937,N_23686,N_23712);
xor U23938 (N_23938,N_23525,N_23659);
nor U23939 (N_23939,N_23608,N_23664);
nand U23940 (N_23940,N_23589,N_23585);
nor U23941 (N_23941,N_23560,N_23656);
and U23942 (N_23942,N_23633,N_23536);
and U23943 (N_23943,N_23657,N_23624);
nor U23944 (N_23944,N_23521,N_23619);
or U23945 (N_23945,N_23574,N_23509);
and U23946 (N_23946,N_23606,N_23610);
nor U23947 (N_23947,N_23707,N_23684);
nor U23948 (N_23948,N_23730,N_23509);
xor U23949 (N_23949,N_23529,N_23688);
nand U23950 (N_23950,N_23657,N_23655);
nand U23951 (N_23951,N_23510,N_23579);
nand U23952 (N_23952,N_23515,N_23551);
and U23953 (N_23953,N_23598,N_23525);
and U23954 (N_23954,N_23700,N_23535);
or U23955 (N_23955,N_23557,N_23646);
nand U23956 (N_23956,N_23622,N_23695);
or U23957 (N_23957,N_23694,N_23663);
nand U23958 (N_23958,N_23530,N_23518);
or U23959 (N_23959,N_23642,N_23669);
nand U23960 (N_23960,N_23590,N_23643);
nand U23961 (N_23961,N_23633,N_23569);
and U23962 (N_23962,N_23676,N_23701);
and U23963 (N_23963,N_23556,N_23666);
nand U23964 (N_23964,N_23659,N_23719);
and U23965 (N_23965,N_23729,N_23555);
nor U23966 (N_23966,N_23713,N_23549);
and U23967 (N_23967,N_23734,N_23613);
nand U23968 (N_23968,N_23654,N_23592);
nor U23969 (N_23969,N_23700,N_23614);
nand U23970 (N_23970,N_23505,N_23696);
nand U23971 (N_23971,N_23538,N_23593);
nor U23972 (N_23972,N_23716,N_23608);
or U23973 (N_23973,N_23646,N_23671);
and U23974 (N_23974,N_23654,N_23554);
or U23975 (N_23975,N_23534,N_23656);
nor U23976 (N_23976,N_23660,N_23544);
nand U23977 (N_23977,N_23588,N_23708);
nor U23978 (N_23978,N_23725,N_23609);
or U23979 (N_23979,N_23720,N_23590);
nand U23980 (N_23980,N_23509,N_23582);
nor U23981 (N_23981,N_23703,N_23508);
nor U23982 (N_23982,N_23734,N_23626);
nor U23983 (N_23983,N_23666,N_23714);
nand U23984 (N_23984,N_23553,N_23521);
nand U23985 (N_23985,N_23508,N_23718);
and U23986 (N_23986,N_23500,N_23521);
nand U23987 (N_23987,N_23555,N_23635);
nor U23988 (N_23988,N_23597,N_23509);
nor U23989 (N_23989,N_23745,N_23690);
nand U23990 (N_23990,N_23624,N_23541);
nor U23991 (N_23991,N_23682,N_23612);
or U23992 (N_23992,N_23614,N_23698);
or U23993 (N_23993,N_23599,N_23683);
nor U23994 (N_23994,N_23725,N_23672);
nand U23995 (N_23995,N_23720,N_23668);
and U23996 (N_23996,N_23716,N_23673);
or U23997 (N_23997,N_23660,N_23553);
xnor U23998 (N_23998,N_23546,N_23515);
and U23999 (N_23999,N_23680,N_23695);
nor U24000 (N_24000,N_23987,N_23811);
and U24001 (N_24001,N_23925,N_23947);
nor U24002 (N_24002,N_23978,N_23972);
nand U24003 (N_24003,N_23817,N_23999);
nand U24004 (N_24004,N_23906,N_23815);
or U24005 (N_24005,N_23968,N_23901);
nor U24006 (N_24006,N_23837,N_23903);
or U24007 (N_24007,N_23945,N_23919);
nor U24008 (N_24008,N_23851,N_23823);
or U24009 (N_24009,N_23878,N_23854);
and U24010 (N_24010,N_23967,N_23904);
nor U24011 (N_24011,N_23950,N_23994);
nor U24012 (N_24012,N_23835,N_23969);
nor U24013 (N_24013,N_23764,N_23866);
nor U24014 (N_24014,N_23850,N_23882);
and U24015 (N_24015,N_23941,N_23816);
and U24016 (N_24016,N_23852,N_23791);
and U24017 (N_24017,N_23812,N_23921);
or U24018 (N_24018,N_23979,N_23807);
or U24019 (N_24019,N_23920,N_23803);
and U24020 (N_24020,N_23965,N_23958);
xor U24021 (N_24021,N_23779,N_23960);
and U24022 (N_24022,N_23778,N_23966);
and U24023 (N_24023,N_23822,N_23896);
and U24024 (N_24024,N_23813,N_23897);
or U24025 (N_24025,N_23927,N_23917);
or U24026 (N_24026,N_23944,N_23908);
or U24027 (N_24027,N_23819,N_23998);
and U24028 (N_24028,N_23770,N_23842);
nand U24029 (N_24029,N_23772,N_23847);
or U24030 (N_24030,N_23980,N_23981);
and U24031 (N_24031,N_23789,N_23993);
and U24032 (N_24032,N_23776,N_23991);
or U24033 (N_24033,N_23804,N_23780);
nand U24034 (N_24034,N_23754,N_23957);
and U24035 (N_24035,N_23887,N_23801);
or U24036 (N_24036,N_23809,N_23894);
and U24037 (N_24037,N_23964,N_23939);
nor U24038 (N_24038,N_23821,N_23885);
and U24039 (N_24039,N_23975,N_23907);
nand U24040 (N_24040,N_23860,N_23955);
and U24041 (N_24041,N_23762,N_23900);
and U24042 (N_24042,N_23771,N_23932);
or U24043 (N_24043,N_23784,N_23948);
nand U24044 (N_24044,N_23783,N_23752);
nor U24045 (N_24045,N_23787,N_23858);
or U24046 (N_24046,N_23984,N_23832);
nand U24047 (N_24047,N_23983,N_23830);
and U24048 (N_24048,N_23889,N_23874);
or U24049 (N_24049,N_23761,N_23846);
nor U24050 (N_24050,N_23888,N_23956);
and U24051 (N_24051,N_23794,N_23872);
or U24052 (N_24052,N_23940,N_23934);
nand U24053 (N_24053,N_23829,N_23886);
xor U24054 (N_24054,N_23949,N_23954);
nor U24055 (N_24055,N_23997,N_23871);
or U24056 (N_24056,N_23833,N_23962);
nor U24057 (N_24057,N_23792,N_23861);
xor U24058 (N_24058,N_23953,N_23814);
nand U24059 (N_24059,N_23773,N_23827);
nor U24060 (N_24060,N_23961,N_23884);
nor U24061 (N_24061,N_23877,N_23828);
nand U24062 (N_24062,N_23938,N_23777);
nand U24063 (N_24063,N_23763,N_23862);
nand U24064 (N_24064,N_23793,N_23859);
or U24065 (N_24065,N_23899,N_23911);
and U24066 (N_24066,N_23766,N_23916);
or U24067 (N_24067,N_23869,N_23856);
xor U24068 (N_24068,N_23865,N_23922);
nor U24069 (N_24069,N_23826,N_23912);
or U24070 (N_24070,N_23843,N_23988);
nor U24071 (N_24071,N_23805,N_23818);
xnor U24072 (N_24072,N_23775,N_23937);
xor U24073 (N_24073,N_23910,N_23756);
or U24074 (N_24074,N_23790,N_23879);
nand U24075 (N_24075,N_23845,N_23942);
nor U24076 (N_24076,N_23923,N_23751);
and U24077 (N_24077,N_23909,N_23799);
and U24078 (N_24078,N_23838,N_23785);
nand U24079 (N_24079,N_23935,N_23782);
nand U24080 (N_24080,N_23902,N_23982);
nand U24081 (N_24081,N_23769,N_23929);
xor U24082 (N_24082,N_23825,N_23802);
nand U24083 (N_24083,N_23924,N_23952);
and U24084 (N_24084,N_23855,N_23795);
xor U24085 (N_24085,N_23959,N_23798);
xor U24086 (N_24086,N_23992,N_23824);
nand U24087 (N_24087,N_23977,N_23931);
and U24088 (N_24088,N_23863,N_23893);
xnor U24089 (N_24089,N_23974,N_23786);
or U24090 (N_24090,N_23881,N_23868);
or U24091 (N_24091,N_23928,N_23853);
xor U24092 (N_24092,N_23774,N_23839);
xnor U24093 (N_24093,N_23963,N_23831);
nand U24094 (N_24094,N_23848,N_23836);
xor U24095 (N_24095,N_23913,N_23759);
nand U24096 (N_24096,N_23951,N_23767);
xor U24097 (N_24097,N_23875,N_23765);
xor U24098 (N_24098,N_23989,N_23883);
or U24099 (N_24099,N_23758,N_23936);
and U24100 (N_24100,N_23797,N_23890);
nand U24101 (N_24101,N_23757,N_23844);
and U24102 (N_24102,N_23976,N_23808);
nand U24103 (N_24103,N_23985,N_23760);
nand U24104 (N_24104,N_23990,N_23841);
nand U24105 (N_24105,N_23898,N_23905);
xor U24106 (N_24106,N_23946,N_23820);
or U24107 (N_24107,N_23800,N_23870);
nand U24108 (N_24108,N_23788,N_23973);
nor U24109 (N_24109,N_23750,N_23810);
nand U24110 (N_24110,N_23995,N_23781);
or U24111 (N_24111,N_23864,N_23753);
or U24112 (N_24112,N_23996,N_23930);
nand U24113 (N_24113,N_23796,N_23915);
nor U24114 (N_24114,N_23768,N_23891);
and U24115 (N_24115,N_23943,N_23857);
or U24116 (N_24116,N_23867,N_23880);
nor U24117 (N_24117,N_23914,N_23986);
xor U24118 (N_24118,N_23971,N_23834);
and U24119 (N_24119,N_23895,N_23873);
nor U24120 (N_24120,N_23806,N_23918);
nor U24121 (N_24121,N_23926,N_23755);
and U24122 (N_24122,N_23933,N_23840);
and U24123 (N_24123,N_23970,N_23892);
nand U24124 (N_24124,N_23849,N_23876);
xnor U24125 (N_24125,N_23796,N_23845);
or U24126 (N_24126,N_23963,N_23954);
nor U24127 (N_24127,N_23955,N_23761);
or U24128 (N_24128,N_23890,N_23947);
xnor U24129 (N_24129,N_23780,N_23948);
nand U24130 (N_24130,N_23960,N_23800);
or U24131 (N_24131,N_23891,N_23982);
nand U24132 (N_24132,N_23752,N_23827);
nand U24133 (N_24133,N_23791,N_23869);
or U24134 (N_24134,N_23926,N_23960);
and U24135 (N_24135,N_23895,N_23887);
or U24136 (N_24136,N_23848,N_23979);
nor U24137 (N_24137,N_23938,N_23884);
nor U24138 (N_24138,N_23840,N_23901);
nand U24139 (N_24139,N_23798,N_23750);
xor U24140 (N_24140,N_23996,N_23904);
or U24141 (N_24141,N_23821,N_23751);
or U24142 (N_24142,N_23809,N_23859);
nor U24143 (N_24143,N_23788,N_23799);
nor U24144 (N_24144,N_23841,N_23910);
and U24145 (N_24145,N_23871,N_23985);
or U24146 (N_24146,N_23893,N_23959);
and U24147 (N_24147,N_23830,N_23887);
nand U24148 (N_24148,N_23916,N_23851);
or U24149 (N_24149,N_23760,N_23902);
nor U24150 (N_24150,N_23876,N_23886);
and U24151 (N_24151,N_23794,N_23767);
nand U24152 (N_24152,N_23857,N_23974);
and U24153 (N_24153,N_23875,N_23872);
nand U24154 (N_24154,N_23915,N_23926);
nor U24155 (N_24155,N_23794,N_23958);
nor U24156 (N_24156,N_23896,N_23887);
nor U24157 (N_24157,N_23810,N_23944);
nand U24158 (N_24158,N_23854,N_23903);
nand U24159 (N_24159,N_23933,N_23811);
xor U24160 (N_24160,N_23814,N_23876);
and U24161 (N_24161,N_23766,N_23971);
xnor U24162 (N_24162,N_23793,N_23813);
nor U24163 (N_24163,N_23950,N_23906);
and U24164 (N_24164,N_23785,N_23916);
or U24165 (N_24165,N_23857,N_23950);
nor U24166 (N_24166,N_23919,N_23898);
nor U24167 (N_24167,N_23775,N_23829);
nor U24168 (N_24168,N_23753,N_23929);
xor U24169 (N_24169,N_23776,N_23877);
or U24170 (N_24170,N_23777,N_23910);
or U24171 (N_24171,N_23759,N_23816);
xor U24172 (N_24172,N_23761,N_23962);
xor U24173 (N_24173,N_23854,N_23851);
nor U24174 (N_24174,N_23958,N_23778);
nor U24175 (N_24175,N_23904,N_23997);
and U24176 (N_24176,N_23894,N_23903);
xor U24177 (N_24177,N_23839,N_23808);
nor U24178 (N_24178,N_23757,N_23833);
and U24179 (N_24179,N_23751,N_23838);
nor U24180 (N_24180,N_23776,N_23995);
or U24181 (N_24181,N_23905,N_23891);
or U24182 (N_24182,N_23958,N_23891);
and U24183 (N_24183,N_23832,N_23928);
and U24184 (N_24184,N_23944,N_23913);
nor U24185 (N_24185,N_23762,N_23842);
and U24186 (N_24186,N_23775,N_23784);
or U24187 (N_24187,N_23841,N_23918);
nor U24188 (N_24188,N_23921,N_23953);
and U24189 (N_24189,N_23988,N_23944);
and U24190 (N_24190,N_23762,N_23795);
nand U24191 (N_24191,N_23869,N_23811);
or U24192 (N_24192,N_23936,N_23753);
or U24193 (N_24193,N_23818,N_23751);
nor U24194 (N_24194,N_23797,N_23919);
nor U24195 (N_24195,N_23879,N_23786);
or U24196 (N_24196,N_23992,N_23895);
xnor U24197 (N_24197,N_23960,N_23936);
nor U24198 (N_24198,N_23858,N_23832);
or U24199 (N_24199,N_23785,N_23835);
and U24200 (N_24200,N_23812,N_23774);
nor U24201 (N_24201,N_23957,N_23852);
or U24202 (N_24202,N_23756,N_23815);
nor U24203 (N_24203,N_23979,N_23952);
and U24204 (N_24204,N_23817,N_23772);
or U24205 (N_24205,N_23991,N_23926);
and U24206 (N_24206,N_23848,N_23846);
xor U24207 (N_24207,N_23886,N_23894);
or U24208 (N_24208,N_23872,N_23799);
nor U24209 (N_24209,N_23885,N_23819);
and U24210 (N_24210,N_23871,N_23827);
and U24211 (N_24211,N_23844,N_23805);
nand U24212 (N_24212,N_23977,N_23840);
and U24213 (N_24213,N_23924,N_23871);
and U24214 (N_24214,N_23952,N_23977);
nor U24215 (N_24215,N_23976,N_23967);
nand U24216 (N_24216,N_23897,N_23777);
and U24217 (N_24217,N_23813,N_23809);
and U24218 (N_24218,N_23934,N_23831);
and U24219 (N_24219,N_23784,N_23943);
nand U24220 (N_24220,N_23960,N_23796);
nor U24221 (N_24221,N_23823,N_23962);
and U24222 (N_24222,N_23851,N_23764);
or U24223 (N_24223,N_23932,N_23796);
or U24224 (N_24224,N_23976,N_23986);
or U24225 (N_24225,N_23894,N_23970);
or U24226 (N_24226,N_23934,N_23922);
and U24227 (N_24227,N_23796,N_23779);
and U24228 (N_24228,N_23961,N_23862);
nand U24229 (N_24229,N_23999,N_23938);
or U24230 (N_24230,N_23855,N_23771);
xor U24231 (N_24231,N_23948,N_23839);
nand U24232 (N_24232,N_23911,N_23815);
and U24233 (N_24233,N_23938,N_23869);
nand U24234 (N_24234,N_23910,N_23912);
and U24235 (N_24235,N_23827,N_23876);
nand U24236 (N_24236,N_23848,N_23817);
and U24237 (N_24237,N_23831,N_23777);
and U24238 (N_24238,N_23998,N_23883);
nand U24239 (N_24239,N_23884,N_23759);
nor U24240 (N_24240,N_23878,N_23922);
nor U24241 (N_24241,N_23778,N_23850);
nor U24242 (N_24242,N_23894,N_23817);
and U24243 (N_24243,N_23997,N_23929);
nor U24244 (N_24244,N_23839,N_23978);
nor U24245 (N_24245,N_23977,N_23788);
or U24246 (N_24246,N_23945,N_23846);
or U24247 (N_24247,N_23935,N_23812);
nand U24248 (N_24248,N_23984,N_23987);
nand U24249 (N_24249,N_23999,N_23852);
or U24250 (N_24250,N_24030,N_24236);
or U24251 (N_24251,N_24006,N_24108);
nor U24252 (N_24252,N_24079,N_24090);
xor U24253 (N_24253,N_24103,N_24166);
nor U24254 (N_24254,N_24092,N_24242);
nand U24255 (N_24255,N_24181,N_24057);
nor U24256 (N_24256,N_24104,N_24048);
nor U24257 (N_24257,N_24110,N_24188);
nand U24258 (N_24258,N_24225,N_24240);
and U24259 (N_24259,N_24034,N_24131);
and U24260 (N_24260,N_24222,N_24126);
nor U24261 (N_24261,N_24196,N_24217);
or U24262 (N_24262,N_24113,N_24117);
nand U24263 (N_24263,N_24195,N_24033);
xnor U24264 (N_24264,N_24139,N_24074);
nand U24265 (N_24265,N_24172,N_24244);
nor U24266 (N_24266,N_24043,N_24032);
or U24267 (N_24267,N_24071,N_24054);
and U24268 (N_24268,N_24206,N_24067);
or U24269 (N_24269,N_24098,N_24159);
xor U24270 (N_24270,N_24189,N_24066);
nor U24271 (N_24271,N_24199,N_24115);
nor U24272 (N_24272,N_24132,N_24152);
or U24273 (N_24273,N_24018,N_24137);
nor U24274 (N_24274,N_24101,N_24239);
nor U24275 (N_24275,N_24022,N_24216);
nor U24276 (N_24276,N_24121,N_24047);
or U24277 (N_24277,N_24096,N_24142);
and U24278 (N_24278,N_24220,N_24144);
or U24279 (N_24279,N_24102,N_24243);
and U24280 (N_24280,N_24192,N_24179);
nand U24281 (N_24281,N_24176,N_24028);
or U24282 (N_24282,N_24190,N_24191);
and U24283 (N_24283,N_24171,N_24045);
and U24284 (N_24284,N_24037,N_24138);
xor U24285 (N_24285,N_24241,N_24174);
nand U24286 (N_24286,N_24201,N_24182);
or U24287 (N_24287,N_24249,N_24170);
nand U24288 (N_24288,N_24025,N_24233);
and U24289 (N_24289,N_24133,N_24080);
or U24290 (N_24290,N_24061,N_24178);
and U24291 (N_24291,N_24013,N_24146);
and U24292 (N_24292,N_24085,N_24149);
and U24293 (N_24293,N_24135,N_24040);
xor U24294 (N_24294,N_24058,N_24050);
and U24295 (N_24295,N_24002,N_24091);
and U24296 (N_24296,N_24031,N_24122);
nand U24297 (N_24297,N_24016,N_24087);
and U24298 (N_24298,N_24237,N_24062);
nand U24299 (N_24299,N_24059,N_24235);
xnor U24300 (N_24300,N_24214,N_24036);
nor U24301 (N_24301,N_24218,N_24183);
nand U24302 (N_24302,N_24095,N_24046);
nor U24303 (N_24303,N_24082,N_24205);
and U24304 (N_24304,N_24068,N_24078);
and U24305 (N_24305,N_24223,N_24177);
and U24306 (N_24306,N_24084,N_24215);
nor U24307 (N_24307,N_24148,N_24111);
and U24308 (N_24308,N_24160,N_24020);
or U24309 (N_24309,N_24150,N_24136);
nor U24310 (N_24310,N_24155,N_24081);
and U24311 (N_24311,N_24075,N_24187);
nand U24312 (N_24312,N_24118,N_24209);
nand U24313 (N_24313,N_24051,N_24023);
or U24314 (N_24314,N_24093,N_24105);
or U24315 (N_24315,N_24055,N_24112);
nor U24316 (N_24316,N_24140,N_24197);
nand U24317 (N_24317,N_24017,N_24001);
and U24318 (N_24318,N_24041,N_24232);
nor U24319 (N_24319,N_24106,N_24130);
xnor U24320 (N_24320,N_24229,N_24119);
or U24321 (N_24321,N_24060,N_24029);
nand U24322 (N_24322,N_24238,N_24035);
or U24323 (N_24323,N_24077,N_24154);
xnor U24324 (N_24324,N_24076,N_24009);
nand U24325 (N_24325,N_24194,N_24210);
and U24326 (N_24326,N_24168,N_24014);
nand U24327 (N_24327,N_24158,N_24024);
xnor U24328 (N_24328,N_24072,N_24193);
or U24329 (N_24329,N_24147,N_24202);
xnor U24330 (N_24330,N_24019,N_24008);
and U24331 (N_24331,N_24246,N_24129);
or U24332 (N_24332,N_24185,N_24186);
or U24333 (N_24333,N_24162,N_24089);
nor U24334 (N_24334,N_24083,N_24004);
or U24335 (N_24335,N_24143,N_24044);
xor U24336 (N_24336,N_24107,N_24021);
xnor U24337 (N_24337,N_24027,N_24000);
nor U24338 (N_24338,N_24204,N_24100);
or U24339 (N_24339,N_24073,N_24151);
xor U24340 (N_24340,N_24169,N_24094);
nand U24341 (N_24341,N_24226,N_24065);
nand U24342 (N_24342,N_24114,N_24026);
nor U24343 (N_24343,N_24049,N_24015);
or U24344 (N_24344,N_24247,N_24120);
nor U24345 (N_24345,N_24056,N_24200);
xnor U24346 (N_24346,N_24231,N_24180);
nand U24347 (N_24347,N_24141,N_24003);
nand U24348 (N_24348,N_24039,N_24245);
nor U24349 (N_24349,N_24128,N_24153);
xnor U24350 (N_24350,N_24234,N_24156);
nor U24351 (N_24351,N_24012,N_24167);
nor U24352 (N_24352,N_24212,N_24184);
and U24353 (N_24353,N_24228,N_24207);
or U24354 (N_24354,N_24007,N_24099);
and U24355 (N_24355,N_24010,N_24097);
nor U24356 (N_24356,N_24164,N_24219);
nand U24357 (N_24357,N_24005,N_24213);
or U24358 (N_24358,N_24124,N_24063);
nand U24359 (N_24359,N_24165,N_24161);
or U24360 (N_24360,N_24042,N_24230);
nand U24361 (N_24361,N_24125,N_24163);
nand U24362 (N_24362,N_24064,N_24157);
and U24363 (N_24363,N_24134,N_24227);
nand U24364 (N_24364,N_24109,N_24069);
nand U24365 (N_24365,N_24123,N_24052);
or U24366 (N_24366,N_24175,N_24116);
xor U24367 (N_24367,N_24070,N_24203);
xor U24368 (N_24368,N_24088,N_24011);
or U24369 (N_24369,N_24145,N_24053);
xnor U24370 (N_24370,N_24127,N_24173);
nand U24371 (N_24371,N_24198,N_24208);
or U24372 (N_24372,N_24086,N_24038);
or U24373 (N_24373,N_24211,N_24224);
nor U24374 (N_24374,N_24221,N_24248);
nor U24375 (N_24375,N_24231,N_24002);
or U24376 (N_24376,N_24018,N_24164);
nand U24377 (N_24377,N_24038,N_24143);
nand U24378 (N_24378,N_24002,N_24201);
nor U24379 (N_24379,N_24231,N_24106);
nor U24380 (N_24380,N_24042,N_24232);
nand U24381 (N_24381,N_24228,N_24236);
and U24382 (N_24382,N_24124,N_24187);
nand U24383 (N_24383,N_24170,N_24164);
and U24384 (N_24384,N_24014,N_24185);
nand U24385 (N_24385,N_24234,N_24055);
nor U24386 (N_24386,N_24031,N_24224);
and U24387 (N_24387,N_24038,N_24032);
xor U24388 (N_24388,N_24123,N_24209);
nand U24389 (N_24389,N_24122,N_24103);
and U24390 (N_24390,N_24149,N_24018);
nand U24391 (N_24391,N_24020,N_24038);
or U24392 (N_24392,N_24032,N_24132);
nand U24393 (N_24393,N_24009,N_24221);
nand U24394 (N_24394,N_24225,N_24010);
or U24395 (N_24395,N_24129,N_24159);
nor U24396 (N_24396,N_24163,N_24061);
xor U24397 (N_24397,N_24166,N_24067);
and U24398 (N_24398,N_24118,N_24049);
or U24399 (N_24399,N_24035,N_24146);
nor U24400 (N_24400,N_24064,N_24072);
and U24401 (N_24401,N_24179,N_24237);
and U24402 (N_24402,N_24229,N_24200);
nor U24403 (N_24403,N_24172,N_24215);
nand U24404 (N_24404,N_24176,N_24217);
or U24405 (N_24405,N_24213,N_24107);
and U24406 (N_24406,N_24047,N_24157);
nor U24407 (N_24407,N_24185,N_24202);
nand U24408 (N_24408,N_24035,N_24055);
nor U24409 (N_24409,N_24012,N_24221);
and U24410 (N_24410,N_24002,N_24084);
xnor U24411 (N_24411,N_24065,N_24208);
and U24412 (N_24412,N_24003,N_24171);
nand U24413 (N_24413,N_24041,N_24133);
nand U24414 (N_24414,N_24060,N_24048);
and U24415 (N_24415,N_24013,N_24187);
nor U24416 (N_24416,N_24100,N_24047);
xor U24417 (N_24417,N_24205,N_24242);
or U24418 (N_24418,N_24238,N_24009);
nand U24419 (N_24419,N_24046,N_24182);
nor U24420 (N_24420,N_24214,N_24019);
nand U24421 (N_24421,N_24220,N_24060);
xnor U24422 (N_24422,N_24058,N_24113);
nor U24423 (N_24423,N_24078,N_24035);
or U24424 (N_24424,N_24026,N_24225);
and U24425 (N_24425,N_24034,N_24006);
xnor U24426 (N_24426,N_24240,N_24053);
nand U24427 (N_24427,N_24178,N_24183);
and U24428 (N_24428,N_24160,N_24120);
or U24429 (N_24429,N_24079,N_24145);
or U24430 (N_24430,N_24045,N_24248);
and U24431 (N_24431,N_24016,N_24219);
or U24432 (N_24432,N_24113,N_24162);
nor U24433 (N_24433,N_24030,N_24227);
nor U24434 (N_24434,N_24075,N_24005);
xnor U24435 (N_24435,N_24244,N_24226);
and U24436 (N_24436,N_24020,N_24060);
or U24437 (N_24437,N_24202,N_24084);
nand U24438 (N_24438,N_24010,N_24091);
or U24439 (N_24439,N_24094,N_24223);
nor U24440 (N_24440,N_24192,N_24045);
nand U24441 (N_24441,N_24211,N_24212);
and U24442 (N_24442,N_24084,N_24168);
or U24443 (N_24443,N_24181,N_24054);
nor U24444 (N_24444,N_24213,N_24025);
and U24445 (N_24445,N_24125,N_24195);
nor U24446 (N_24446,N_24111,N_24040);
nand U24447 (N_24447,N_24018,N_24168);
xor U24448 (N_24448,N_24093,N_24186);
or U24449 (N_24449,N_24104,N_24152);
nor U24450 (N_24450,N_24181,N_24110);
xor U24451 (N_24451,N_24161,N_24180);
and U24452 (N_24452,N_24146,N_24231);
or U24453 (N_24453,N_24218,N_24056);
nand U24454 (N_24454,N_24133,N_24113);
and U24455 (N_24455,N_24100,N_24151);
nor U24456 (N_24456,N_24224,N_24193);
xnor U24457 (N_24457,N_24120,N_24156);
xnor U24458 (N_24458,N_24112,N_24196);
nand U24459 (N_24459,N_24021,N_24045);
nor U24460 (N_24460,N_24046,N_24165);
xnor U24461 (N_24461,N_24048,N_24133);
nor U24462 (N_24462,N_24050,N_24212);
and U24463 (N_24463,N_24098,N_24132);
nand U24464 (N_24464,N_24173,N_24197);
xor U24465 (N_24465,N_24171,N_24021);
xnor U24466 (N_24466,N_24217,N_24087);
nand U24467 (N_24467,N_24048,N_24011);
or U24468 (N_24468,N_24231,N_24047);
nand U24469 (N_24469,N_24039,N_24071);
and U24470 (N_24470,N_24242,N_24047);
nor U24471 (N_24471,N_24008,N_24153);
and U24472 (N_24472,N_24052,N_24186);
xnor U24473 (N_24473,N_24011,N_24244);
or U24474 (N_24474,N_24201,N_24138);
or U24475 (N_24475,N_24138,N_24215);
and U24476 (N_24476,N_24176,N_24214);
nor U24477 (N_24477,N_24084,N_24140);
nor U24478 (N_24478,N_24172,N_24223);
or U24479 (N_24479,N_24014,N_24103);
or U24480 (N_24480,N_24031,N_24187);
or U24481 (N_24481,N_24089,N_24232);
and U24482 (N_24482,N_24076,N_24177);
nand U24483 (N_24483,N_24007,N_24029);
xor U24484 (N_24484,N_24040,N_24249);
nand U24485 (N_24485,N_24038,N_24016);
or U24486 (N_24486,N_24123,N_24183);
nand U24487 (N_24487,N_24118,N_24101);
xor U24488 (N_24488,N_24195,N_24243);
nor U24489 (N_24489,N_24116,N_24044);
nand U24490 (N_24490,N_24232,N_24088);
and U24491 (N_24491,N_24087,N_24092);
or U24492 (N_24492,N_24078,N_24190);
nand U24493 (N_24493,N_24143,N_24080);
nor U24494 (N_24494,N_24127,N_24163);
or U24495 (N_24495,N_24029,N_24045);
nor U24496 (N_24496,N_24054,N_24176);
and U24497 (N_24497,N_24130,N_24019);
nor U24498 (N_24498,N_24225,N_24152);
nor U24499 (N_24499,N_24071,N_24065);
nand U24500 (N_24500,N_24302,N_24442);
nor U24501 (N_24501,N_24493,N_24342);
xor U24502 (N_24502,N_24437,N_24388);
or U24503 (N_24503,N_24319,N_24262);
and U24504 (N_24504,N_24270,N_24325);
or U24505 (N_24505,N_24484,N_24488);
nor U24506 (N_24506,N_24457,N_24369);
xnor U24507 (N_24507,N_24382,N_24337);
nand U24508 (N_24508,N_24349,N_24474);
or U24509 (N_24509,N_24313,N_24362);
or U24510 (N_24510,N_24403,N_24404);
nand U24511 (N_24511,N_24451,N_24256);
nor U24512 (N_24512,N_24315,N_24425);
or U24513 (N_24513,N_24408,N_24334);
nand U24514 (N_24514,N_24459,N_24423);
and U24515 (N_24515,N_24291,N_24265);
or U24516 (N_24516,N_24267,N_24417);
nand U24517 (N_24517,N_24480,N_24399);
and U24518 (N_24518,N_24298,N_24483);
and U24519 (N_24519,N_24365,N_24301);
or U24520 (N_24520,N_24416,N_24329);
nand U24521 (N_24521,N_24448,N_24432);
nor U24522 (N_24522,N_24295,N_24309);
nor U24523 (N_24523,N_24438,N_24418);
nand U24524 (N_24524,N_24394,N_24429);
nor U24525 (N_24525,N_24494,N_24278);
or U24526 (N_24526,N_24328,N_24391);
and U24527 (N_24527,N_24443,N_24297);
nand U24528 (N_24528,N_24387,N_24456);
nor U24529 (N_24529,N_24414,N_24435);
or U24530 (N_24530,N_24348,N_24396);
or U24531 (N_24531,N_24286,N_24282);
or U24532 (N_24532,N_24486,N_24402);
nand U24533 (N_24533,N_24499,N_24462);
nor U24534 (N_24534,N_24268,N_24340);
and U24535 (N_24535,N_24312,N_24424);
or U24536 (N_24536,N_24250,N_24271);
nor U24537 (N_24537,N_24284,N_24273);
and U24538 (N_24538,N_24401,N_24446);
or U24539 (N_24539,N_24283,N_24374);
nor U24540 (N_24540,N_24279,N_24415);
xor U24541 (N_24541,N_24377,N_24386);
or U24542 (N_24542,N_24281,N_24287);
xor U24543 (N_24543,N_24489,N_24272);
xor U24544 (N_24544,N_24449,N_24350);
nand U24545 (N_24545,N_24398,N_24355);
nor U24546 (N_24546,N_24294,N_24371);
xor U24547 (N_24547,N_24364,N_24482);
and U24548 (N_24548,N_24370,N_24367);
and U24549 (N_24549,N_24338,N_24336);
nand U24550 (N_24550,N_24277,N_24257);
nand U24551 (N_24551,N_24352,N_24412);
and U24552 (N_24552,N_24356,N_24330);
and U24553 (N_24553,N_24254,N_24314);
and U24554 (N_24554,N_24373,N_24419);
nor U24555 (N_24555,N_24375,N_24263);
nand U24556 (N_24556,N_24380,N_24491);
or U24557 (N_24557,N_24469,N_24379);
nor U24558 (N_24558,N_24485,N_24339);
and U24559 (N_24559,N_24308,N_24310);
nand U24560 (N_24560,N_24467,N_24395);
nor U24561 (N_24561,N_24280,N_24397);
and U24562 (N_24562,N_24269,N_24468);
and U24563 (N_24563,N_24343,N_24274);
or U24564 (N_24564,N_24357,N_24420);
or U24565 (N_24565,N_24345,N_24458);
xor U24566 (N_24566,N_24441,N_24430);
or U24567 (N_24567,N_24450,N_24445);
or U24568 (N_24568,N_24498,N_24361);
nor U24569 (N_24569,N_24368,N_24487);
and U24570 (N_24570,N_24358,N_24320);
nand U24571 (N_24571,N_24427,N_24296);
or U24572 (N_24572,N_24477,N_24366);
nand U24573 (N_24573,N_24495,N_24479);
nor U24574 (N_24574,N_24376,N_24318);
nor U24575 (N_24575,N_24436,N_24347);
nor U24576 (N_24576,N_24390,N_24316);
nor U24577 (N_24577,N_24306,N_24255);
or U24578 (N_24578,N_24260,N_24351);
nand U24579 (N_24579,N_24431,N_24473);
and U24580 (N_24580,N_24292,N_24251);
and U24581 (N_24581,N_24496,N_24470);
nor U24582 (N_24582,N_24406,N_24407);
nor U24583 (N_24583,N_24475,N_24454);
xor U24584 (N_24584,N_24461,N_24490);
nand U24585 (N_24585,N_24497,N_24321);
or U24586 (N_24586,N_24428,N_24266);
and U24587 (N_24587,N_24264,N_24384);
nor U24588 (N_24588,N_24466,N_24317);
nand U24589 (N_24589,N_24422,N_24444);
or U24590 (N_24590,N_24307,N_24259);
xor U24591 (N_24591,N_24332,N_24465);
nor U24592 (N_24592,N_24289,N_24413);
nor U24593 (N_24593,N_24344,N_24288);
nand U24594 (N_24594,N_24372,N_24275);
or U24595 (N_24595,N_24359,N_24433);
nand U24596 (N_24596,N_24447,N_24324);
nor U24597 (N_24597,N_24405,N_24290);
nor U24598 (N_24598,N_24305,N_24327);
or U24599 (N_24599,N_24363,N_24392);
and U24600 (N_24600,N_24385,N_24426);
and U24601 (N_24601,N_24476,N_24421);
nand U24602 (N_24602,N_24460,N_24439);
and U24603 (N_24603,N_24393,N_24378);
or U24604 (N_24604,N_24455,N_24472);
nand U24605 (N_24605,N_24492,N_24303);
or U24606 (N_24606,N_24440,N_24410);
xor U24607 (N_24607,N_24354,N_24383);
and U24608 (N_24608,N_24253,N_24400);
nand U24609 (N_24609,N_24285,N_24331);
nor U24610 (N_24610,N_24335,N_24300);
xor U24611 (N_24611,N_24353,N_24299);
nor U24612 (N_24612,N_24326,N_24411);
and U24613 (N_24613,N_24463,N_24293);
xnor U24614 (N_24614,N_24478,N_24434);
nor U24615 (N_24615,N_24261,N_24471);
xnor U24616 (N_24616,N_24323,N_24409);
xor U24617 (N_24617,N_24464,N_24452);
xnor U24618 (N_24618,N_24481,N_24346);
nor U24619 (N_24619,N_24252,N_24322);
nor U24620 (N_24620,N_24304,N_24389);
and U24621 (N_24621,N_24311,N_24333);
nor U24622 (N_24622,N_24341,N_24381);
and U24623 (N_24623,N_24453,N_24360);
nor U24624 (N_24624,N_24258,N_24276);
or U24625 (N_24625,N_24490,N_24418);
or U24626 (N_24626,N_24406,N_24342);
or U24627 (N_24627,N_24470,N_24280);
nand U24628 (N_24628,N_24289,N_24291);
or U24629 (N_24629,N_24481,N_24482);
or U24630 (N_24630,N_24272,N_24497);
and U24631 (N_24631,N_24293,N_24308);
nand U24632 (N_24632,N_24272,N_24397);
nand U24633 (N_24633,N_24387,N_24360);
nand U24634 (N_24634,N_24292,N_24340);
nand U24635 (N_24635,N_24311,N_24413);
nor U24636 (N_24636,N_24295,N_24413);
nor U24637 (N_24637,N_24314,N_24286);
xnor U24638 (N_24638,N_24414,N_24369);
and U24639 (N_24639,N_24322,N_24492);
nand U24640 (N_24640,N_24289,N_24389);
and U24641 (N_24641,N_24465,N_24282);
nor U24642 (N_24642,N_24381,N_24331);
nand U24643 (N_24643,N_24318,N_24408);
and U24644 (N_24644,N_24486,N_24262);
or U24645 (N_24645,N_24418,N_24399);
nand U24646 (N_24646,N_24265,N_24375);
and U24647 (N_24647,N_24270,N_24445);
nand U24648 (N_24648,N_24264,N_24480);
nor U24649 (N_24649,N_24416,N_24273);
or U24650 (N_24650,N_24354,N_24336);
nand U24651 (N_24651,N_24414,N_24363);
or U24652 (N_24652,N_24305,N_24486);
nor U24653 (N_24653,N_24257,N_24293);
nand U24654 (N_24654,N_24393,N_24486);
nor U24655 (N_24655,N_24379,N_24334);
nor U24656 (N_24656,N_24289,N_24328);
and U24657 (N_24657,N_24296,N_24344);
nor U24658 (N_24658,N_24395,N_24278);
or U24659 (N_24659,N_24397,N_24401);
xor U24660 (N_24660,N_24407,N_24293);
and U24661 (N_24661,N_24359,N_24264);
and U24662 (N_24662,N_24411,N_24444);
and U24663 (N_24663,N_24498,N_24492);
nand U24664 (N_24664,N_24317,N_24345);
or U24665 (N_24665,N_24307,N_24329);
or U24666 (N_24666,N_24449,N_24303);
nand U24667 (N_24667,N_24365,N_24282);
and U24668 (N_24668,N_24451,N_24497);
or U24669 (N_24669,N_24336,N_24465);
nand U24670 (N_24670,N_24339,N_24422);
or U24671 (N_24671,N_24433,N_24311);
or U24672 (N_24672,N_24421,N_24409);
xnor U24673 (N_24673,N_24460,N_24391);
nand U24674 (N_24674,N_24458,N_24462);
nor U24675 (N_24675,N_24491,N_24433);
nand U24676 (N_24676,N_24393,N_24473);
nand U24677 (N_24677,N_24262,N_24452);
and U24678 (N_24678,N_24403,N_24317);
and U24679 (N_24679,N_24367,N_24305);
nor U24680 (N_24680,N_24493,N_24379);
or U24681 (N_24681,N_24415,N_24423);
or U24682 (N_24682,N_24325,N_24266);
or U24683 (N_24683,N_24368,N_24467);
xor U24684 (N_24684,N_24304,N_24375);
and U24685 (N_24685,N_24263,N_24422);
nand U24686 (N_24686,N_24269,N_24310);
nor U24687 (N_24687,N_24389,N_24498);
nor U24688 (N_24688,N_24411,N_24416);
or U24689 (N_24689,N_24445,N_24265);
nand U24690 (N_24690,N_24375,N_24416);
and U24691 (N_24691,N_24314,N_24262);
or U24692 (N_24692,N_24384,N_24328);
nand U24693 (N_24693,N_24327,N_24314);
or U24694 (N_24694,N_24494,N_24463);
xor U24695 (N_24695,N_24251,N_24349);
or U24696 (N_24696,N_24265,N_24491);
nor U24697 (N_24697,N_24312,N_24386);
nor U24698 (N_24698,N_24307,N_24475);
and U24699 (N_24699,N_24259,N_24326);
nand U24700 (N_24700,N_24371,N_24497);
xor U24701 (N_24701,N_24426,N_24369);
nand U24702 (N_24702,N_24284,N_24344);
nand U24703 (N_24703,N_24395,N_24309);
nor U24704 (N_24704,N_24325,N_24286);
and U24705 (N_24705,N_24431,N_24438);
or U24706 (N_24706,N_24412,N_24491);
nand U24707 (N_24707,N_24277,N_24481);
and U24708 (N_24708,N_24272,N_24364);
xor U24709 (N_24709,N_24413,N_24375);
nand U24710 (N_24710,N_24383,N_24309);
nor U24711 (N_24711,N_24444,N_24437);
xor U24712 (N_24712,N_24385,N_24254);
nand U24713 (N_24713,N_24413,N_24496);
or U24714 (N_24714,N_24282,N_24435);
nand U24715 (N_24715,N_24403,N_24472);
nor U24716 (N_24716,N_24395,N_24373);
nor U24717 (N_24717,N_24375,N_24362);
and U24718 (N_24718,N_24428,N_24449);
nor U24719 (N_24719,N_24344,N_24493);
xor U24720 (N_24720,N_24386,N_24316);
nand U24721 (N_24721,N_24259,N_24372);
nor U24722 (N_24722,N_24303,N_24495);
and U24723 (N_24723,N_24339,N_24477);
and U24724 (N_24724,N_24496,N_24351);
xnor U24725 (N_24725,N_24358,N_24352);
nor U24726 (N_24726,N_24436,N_24327);
and U24727 (N_24727,N_24379,N_24391);
nor U24728 (N_24728,N_24384,N_24485);
nor U24729 (N_24729,N_24372,N_24473);
and U24730 (N_24730,N_24422,N_24327);
or U24731 (N_24731,N_24313,N_24283);
or U24732 (N_24732,N_24382,N_24278);
or U24733 (N_24733,N_24402,N_24345);
or U24734 (N_24734,N_24353,N_24260);
nand U24735 (N_24735,N_24480,N_24404);
or U24736 (N_24736,N_24491,N_24498);
or U24737 (N_24737,N_24367,N_24412);
xnor U24738 (N_24738,N_24301,N_24394);
and U24739 (N_24739,N_24303,N_24454);
and U24740 (N_24740,N_24269,N_24358);
nand U24741 (N_24741,N_24425,N_24375);
nand U24742 (N_24742,N_24380,N_24472);
and U24743 (N_24743,N_24258,N_24420);
or U24744 (N_24744,N_24312,N_24331);
nand U24745 (N_24745,N_24311,N_24404);
or U24746 (N_24746,N_24422,N_24461);
xnor U24747 (N_24747,N_24402,N_24285);
nand U24748 (N_24748,N_24268,N_24380);
and U24749 (N_24749,N_24280,N_24456);
xor U24750 (N_24750,N_24693,N_24609);
nor U24751 (N_24751,N_24697,N_24724);
and U24752 (N_24752,N_24517,N_24510);
nand U24753 (N_24753,N_24643,N_24619);
or U24754 (N_24754,N_24637,N_24587);
and U24755 (N_24755,N_24727,N_24599);
nor U24756 (N_24756,N_24584,N_24733);
nand U24757 (N_24757,N_24570,N_24509);
xnor U24758 (N_24758,N_24628,N_24748);
xnor U24759 (N_24759,N_24592,N_24665);
and U24760 (N_24760,N_24514,N_24681);
xor U24761 (N_24761,N_24565,N_24554);
nand U24762 (N_24762,N_24660,N_24677);
nand U24763 (N_24763,N_24690,N_24647);
nand U24764 (N_24764,N_24729,N_24708);
or U24765 (N_24765,N_24664,N_24683);
nand U24766 (N_24766,N_24616,N_24745);
nor U24767 (N_24767,N_24659,N_24550);
or U24768 (N_24768,N_24582,N_24607);
and U24769 (N_24769,N_24601,N_24544);
nand U24770 (N_24770,N_24534,N_24716);
and U24771 (N_24771,N_24692,N_24728);
nor U24772 (N_24772,N_24702,N_24615);
xor U24773 (N_24773,N_24563,N_24541);
or U24774 (N_24774,N_24537,N_24680);
or U24775 (N_24775,N_24649,N_24545);
or U24776 (N_24776,N_24663,N_24633);
nor U24777 (N_24777,N_24654,N_24595);
or U24778 (N_24778,N_24551,N_24608);
and U24779 (N_24779,N_24524,N_24610);
or U24780 (N_24780,N_24548,N_24596);
xnor U24781 (N_24781,N_24536,N_24526);
nand U24782 (N_24782,N_24682,N_24604);
nor U24783 (N_24783,N_24679,N_24723);
and U24784 (N_24784,N_24673,N_24618);
or U24785 (N_24785,N_24585,N_24533);
nand U24786 (N_24786,N_24711,N_24624);
and U24787 (N_24787,N_24675,N_24655);
or U24788 (N_24788,N_24661,N_24560);
xnor U24789 (N_24789,N_24612,N_24549);
nor U24790 (N_24790,N_24606,N_24740);
or U24791 (N_24791,N_24735,N_24527);
and U24792 (N_24792,N_24694,N_24676);
or U24793 (N_24793,N_24742,N_24744);
nor U24794 (N_24794,N_24622,N_24629);
nor U24795 (N_24795,N_24505,N_24648);
and U24796 (N_24796,N_24642,N_24546);
and U24797 (N_24797,N_24695,N_24523);
and U24798 (N_24798,N_24645,N_24652);
and U24799 (N_24799,N_24686,N_24502);
xnor U24800 (N_24800,N_24623,N_24666);
or U24801 (N_24801,N_24580,N_24578);
nand U24802 (N_24802,N_24700,N_24688);
or U24803 (N_24803,N_24743,N_24719);
nand U24804 (N_24804,N_24540,N_24671);
xnor U24805 (N_24805,N_24529,N_24552);
nand U24806 (N_24806,N_24588,N_24626);
and U24807 (N_24807,N_24662,N_24500);
nor U24808 (N_24808,N_24709,N_24589);
nand U24809 (N_24809,N_24670,N_24739);
and U24810 (N_24810,N_24571,N_24625);
and U24811 (N_24811,N_24641,N_24577);
xor U24812 (N_24812,N_24558,N_24515);
nor U24813 (N_24813,N_24568,N_24520);
or U24814 (N_24814,N_24600,N_24583);
xor U24815 (N_24815,N_24525,N_24516);
nor U24816 (N_24816,N_24542,N_24547);
and U24817 (N_24817,N_24746,N_24653);
nand U24818 (N_24818,N_24712,N_24621);
nor U24819 (N_24819,N_24593,N_24614);
xnor U24820 (N_24820,N_24513,N_24731);
and U24821 (N_24821,N_24687,N_24557);
and U24822 (N_24822,N_24736,N_24564);
nor U24823 (N_24823,N_24539,N_24672);
nor U24824 (N_24824,N_24576,N_24506);
or U24825 (N_24825,N_24636,N_24574);
or U24826 (N_24826,N_24689,N_24705);
or U24827 (N_24827,N_24635,N_24566);
and U24828 (N_24828,N_24611,N_24669);
or U24829 (N_24829,N_24602,N_24646);
nor U24830 (N_24830,N_24696,N_24556);
or U24831 (N_24831,N_24530,N_24734);
nand U24832 (N_24832,N_24532,N_24749);
nand U24833 (N_24833,N_24598,N_24522);
and U24834 (N_24834,N_24722,N_24703);
and U24835 (N_24835,N_24569,N_24627);
nand U24836 (N_24836,N_24644,N_24685);
nand U24837 (N_24837,N_24507,N_24630);
nor U24838 (N_24838,N_24720,N_24535);
nor U24839 (N_24839,N_24543,N_24603);
nor U24840 (N_24840,N_24613,N_24737);
and U24841 (N_24841,N_24590,N_24741);
or U24842 (N_24842,N_24704,N_24504);
nor U24843 (N_24843,N_24718,N_24519);
or U24844 (N_24844,N_24573,N_24555);
nor U24845 (N_24845,N_24632,N_24650);
and U24846 (N_24846,N_24553,N_24725);
nand U24847 (N_24847,N_24691,N_24605);
and U24848 (N_24848,N_24710,N_24738);
or U24849 (N_24849,N_24620,N_24579);
nand U24850 (N_24850,N_24528,N_24698);
xnor U24851 (N_24851,N_24617,N_24674);
xnor U24852 (N_24852,N_24631,N_24699);
nor U24853 (N_24853,N_24684,N_24634);
xor U24854 (N_24854,N_24591,N_24581);
nor U24855 (N_24855,N_24658,N_24562);
and U24856 (N_24856,N_24713,N_24726);
nand U24857 (N_24857,N_24586,N_24521);
nor U24858 (N_24858,N_24730,N_24668);
nand U24859 (N_24859,N_24638,N_24657);
or U24860 (N_24860,N_24508,N_24512);
and U24861 (N_24861,N_24503,N_24561);
nand U24862 (N_24862,N_24732,N_24747);
and U24863 (N_24863,N_24594,N_24715);
xor U24864 (N_24864,N_24721,N_24651);
nor U24865 (N_24865,N_24667,N_24575);
nor U24866 (N_24866,N_24656,N_24678);
nor U24867 (N_24867,N_24518,N_24531);
xor U24868 (N_24868,N_24707,N_24567);
and U24869 (N_24869,N_24639,N_24640);
nand U24870 (N_24870,N_24701,N_24717);
or U24871 (N_24871,N_24706,N_24714);
and U24872 (N_24872,N_24572,N_24511);
nor U24873 (N_24873,N_24597,N_24538);
and U24874 (N_24874,N_24559,N_24501);
or U24875 (N_24875,N_24534,N_24736);
and U24876 (N_24876,N_24539,N_24670);
xnor U24877 (N_24877,N_24617,N_24530);
and U24878 (N_24878,N_24618,N_24613);
or U24879 (N_24879,N_24508,N_24666);
xor U24880 (N_24880,N_24573,N_24585);
nor U24881 (N_24881,N_24713,N_24720);
nand U24882 (N_24882,N_24675,N_24544);
xor U24883 (N_24883,N_24706,N_24663);
and U24884 (N_24884,N_24588,N_24614);
or U24885 (N_24885,N_24663,N_24694);
and U24886 (N_24886,N_24671,N_24703);
nor U24887 (N_24887,N_24637,N_24547);
nor U24888 (N_24888,N_24674,N_24582);
or U24889 (N_24889,N_24544,N_24566);
nor U24890 (N_24890,N_24664,N_24690);
and U24891 (N_24891,N_24548,N_24527);
nor U24892 (N_24892,N_24716,N_24565);
or U24893 (N_24893,N_24739,N_24602);
or U24894 (N_24894,N_24616,N_24713);
nor U24895 (N_24895,N_24585,N_24637);
nand U24896 (N_24896,N_24717,N_24592);
nand U24897 (N_24897,N_24586,N_24709);
or U24898 (N_24898,N_24741,N_24747);
nor U24899 (N_24899,N_24525,N_24692);
nor U24900 (N_24900,N_24587,N_24534);
nor U24901 (N_24901,N_24579,N_24712);
or U24902 (N_24902,N_24565,N_24661);
or U24903 (N_24903,N_24519,N_24728);
nor U24904 (N_24904,N_24741,N_24693);
nor U24905 (N_24905,N_24510,N_24529);
xor U24906 (N_24906,N_24516,N_24564);
and U24907 (N_24907,N_24543,N_24742);
or U24908 (N_24908,N_24740,N_24612);
nor U24909 (N_24909,N_24711,N_24561);
nor U24910 (N_24910,N_24572,N_24688);
or U24911 (N_24911,N_24748,N_24688);
xnor U24912 (N_24912,N_24727,N_24733);
and U24913 (N_24913,N_24557,N_24725);
nand U24914 (N_24914,N_24550,N_24679);
nand U24915 (N_24915,N_24720,N_24537);
nor U24916 (N_24916,N_24505,N_24560);
and U24917 (N_24917,N_24703,N_24514);
xnor U24918 (N_24918,N_24534,N_24559);
nor U24919 (N_24919,N_24631,N_24690);
and U24920 (N_24920,N_24670,N_24712);
nand U24921 (N_24921,N_24532,N_24704);
nand U24922 (N_24922,N_24580,N_24545);
nand U24923 (N_24923,N_24575,N_24719);
nor U24924 (N_24924,N_24705,N_24628);
and U24925 (N_24925,N_24580,N_24542);
or U24926 (N_24926,N_24590,N_24591);
nand U24927 (N_24927,N_24531,N_24502);
or U24928 (N_24928,N_24734,N_24658);
nor U24929 (N_24929,N_24746,N_24638);
and U24930 (N_24930,N_24690,N_24502);
xor U24931 (N_24931,N_24736,N_24543);
nand U24932 (N_24932,N_24514,N_24706);
and U24933 (N_24933,N_24681,N_24626);
and U24934 (N_24934,N_24588,N_24545);
nand U24935 (N_24935,N_24631,N_24632);
or U24936 (N_24936,N_24568,N_24715);
or U24937 (N_24937,N_24719,N_24589);
or U24938 (N_24938,N_24708,N_24749);
and U24939 (N_24939,N_24624,N_24731);
and U24940 (N_24940,N_24650,N_24619);
and U24941 (N_24941,N_24539,N_24637);
and U24942 (N_24942,N_24600,N_24616);
and U24943 (N_24943,N_24547,N_24503);
nand U24944 (N_24944,N_24528,N_24635);
nand U24945 (N_24945,N_24664,N_24723);
or U24946 (N_24946,N_24718,N_24553);
nand U24947 (N_24947,N_24581,N_24740);
and U24948 (N_24948,N_24561,N_24682);
nor U24949 (N_24949,N_24741,N_24551);
and U24950 (N_24950,N_24691,N_24731);
xnor U24951 (N_24951,N_24516,N_24530);
and U24952 (N_24952,N_24599,N_24633);
or U24953 (N_24953,N_24507,N_24626);
and U24954 (N_24954,N_24581,N_24736);
xnor U24955 (N_24955,N_24704,N_24538);
xor U24956 (N_24956,N_24563,N_24601);
and U24957 (N_24957,N_24513,N_24666);
nor U24958 (N_24958,N_24637,N_24569);
nand U24959 (N_24959,N_24654,N_24742);
and U24960 (N_24960,N_24580,N_24667);
nand U24961 (N_24961,N_24519,N_24604);
and U24962 (N_24962,N_24589,N_24636);
and U24963 (N_24963,N_24532,N_24625);
nand U24964 (N_24964,N_24535,N_24700);
nor U24965 (N_24965,N_24603,N_24641);
and U24966 (N_24966,N_24645,N_24622);
and U24967 (N_24967,N_24703,N_24700);
nand U24968 (N_24968,N_24522,N_24712);
or U24969 (N_24969,N_24620,N_24594);
nor U24970 (N_24970,N_24730,N_24527);
or U24971 (N_24971,N_24713,N_24627);
xor U24972 (N_24972,N_24653,N_24654);
xnor U24973 (N_24973,N_24635,N_24665);
xor U24974 (N_24974,N_24677,N_24549);
and U24975 (N_24975,N_24596,N_24521);
nor U24976 (N_24976,N_24678,N_24537);
nand U24977 (N_24977,N_24628,N_24548);
or U24978 (N_24978,N_24511,N_24741);
nand U24979 (N_24979,N_24568,N_24670);
nand U24980 (N_24980,N_24678,N_24558);
nor U24981 (N_24981,N_24528,N_24707);
or U24982 (N_24982,N_24739,N_24532);
nor U24983 (N_24983,N_24613,N_24521);
nor U24984 (N_24984,N_24687,N_24612);
and U24985 (N_24985,N_24585,N_24545);
or U24986 (N_24986,N_24539,N_24674);
and U24987 (N_24987,N_24655,N_24646);
and U24988 (N_24988,N_24680,N_24725);
nor U24989 (N_24989,N_24521,N_24571);
xnor U24990 (N_24990,N_24562,N_24519);
xnor U24991 (N_24991,N_24711,N_24669);
nor U24992 (N_24992,N_24638,N_24680);
or U24993 (N_24993,N_24607,N_24504);
and U24994 (N_24994,N_24540,N_24562);
and U24995 (N_24995,N_24711,N_24574);
and U24996 (N_24996,N_24639,N_24664);
or U24997 (N_24997,N_24673,N_24591);
or U24998 (N_24998,N_24663,N_24603);
nor U24999 (N_24999,N_24657,N_24653);
nor UO_0 (O_0,N_24910,N_24772);
and UO_1 (O_1,N_24903,N_24855);
nand UO_2 (O_2,N_24791,N_24988);
nor UO_3 (O_3,N_24845,N_24783);
nor UO_4 (O_4,N_24941,N_24752);
nor UO_5 (O_5,N_24937,N_24897);
and UO_6 (O_6,N_24890,N_24840);
nor UO_7 (O_7,N_24873,N_24756);
or UO_8 (O_8,N_24814,N_24971);
or UO_9 (O_9,N_24757,N_24964);
nor UO_10 (O_10,N_24750,N_24809);
nand UO_11 (O_11,N_24771,N_24758);
nor UO_12 (O_12,N_24872,N_24821);
and UO_13 (O_13,N_24792,N_24904);
nor UO_14 (O_14,N_24898,N_24906);
nand UO_15 (O_15,N_24879,N_24947);
and UO_16 (O_16,N_24887,N_24769);
or UO_17 (O_17,N_24826,N_24891);
nor UO_18 (O_18,N_24972,N_24975);
nand UO_19 (O_19,N_24944,N_24822);
nor UO_20 (O_20,N_24942,N_24781);
and UO_21 (O_21,N_24852,N_24779);
nor UO_22 (O_22,N_24962,N_24886);
or UO_23 (O_23,N_24768,N_24755);
and UO_24 (O_24,N_24784,N_24895);
or UO_25 (O_25,N_24961,N_24878);
xor UO_26 (O_26,N_24973,N_24935);
or UO_27 (O_27,N_24848,N_24837);
nor UO_28 (O_28,N_24950,N_24853);
and UO_29 (O_29,N_24869,N_24860);
and UO_30 (O_30,N_24923,N_24811);
nor UO_31 (O_31,N_24918,N_24862);
nor UO_32 (O_32,N_24829,N_24987);
nor UO_33 (O_33,N_24767,N_24877);
xnor UO_34 (O_34,N_24966,N_24785);
or UO_35 (O_35,N_24760,N_24948);
and UO_36 (O_36,N_24883,N_24881);
or UO_37 (O_37,N_24907,N_24958);
nand UO_38 (O_38,N_24924,N_24774);
nand UO_39 (O_39,N_24828,N_24936);
nor UO_40 (O_40,N_24765,N_24857);
or UO_41 (O_41,N_24911,N_24797);
or UO_42 (O_42,N_24876,N_24794);
nor UO_43 (O_43,N_24938,N_24925);
or UO_44 (O_44,N_24901,N_24919);
nor UO_45 (O_45,N_24915,N_24846);
or UO_46 (O_46,N_24759,N_24838);
and UO_47 (O_47,N_24946,N_24868);
nor UO_48 (O_48,N_24833,N_24775);
xnor UO_49 (O_49,N_24843,N_24920);
nor UO_50 (O_50,N_24778,N_24932);
nand UO_51 (O_51,N_24863,N_24815);
nand UO_52 (O_52,N_24956,N_24914);
nand UO_53 (O_53,N_24929,N_24803);
xor UO_54 (O_54,N_24945,N_24931);
nand UO_55 (O_55,N_24810,N_24882);
nor UO_56 (O_56,N_24866,N_24812);
or UO_57 (O_57,N_24844,N_24908);
and UO_58 (O_58,N_24871,N_24900);
nand UO_59 (O_59,N_24856,N_24796);
nor UO_60 (O_60,N_24993,N_24793);
xor UO_61 (O_61,N_24850,N_24786);
nand UO_62 (O_62,N_24770,N_24800);
and UO_63 (O_63,N_24957,N_24787);
or UO_64 (O_64,N_24762,N_24991);
and UO_65 (O_65,N_24992,N_24912);
nor UO_66 (O_66,N_24825,N_24806);
or UO_67 (O_67,N_24830,N_24959);
nand UO_68 (O_68,N_24969,N_24854);
nand UO_69 (O_69,N_24974,N_24953);
and UO_70 (O_70,N_24776,N_24965);
or UO_71 (O_71,N_24888,N_24817);
nor UO_72 (O_72,N_24978,N_24799);
nand UO_73 (O_73,N_24819,N_24847);
nor UO_74 (O_74,N_24870,N_24824);
nor UO_75 (O_75,N_24788,N_24808);
nor UO_76 (O_76,N_24789,N_24841);
nor UO_77 (O_77,N_24928,N_24864);
nor UO_78 (O_78,N_24996,N_24827);
nand UO_79 (O_79,N_24985,N_24754);
nor UO_80 (O_80,N_24939,N_24979);
and UO_81 (O_81,N_24943,N_24976);
nand UO_82 (O_82,N_24867,N_24885);
and UO_83 (O_83,N_24980,N_24970);
nor UO_84 (O_84,N_24861,N_24902);
nand UO_85 (O_85,N_24875,N_24832);
nand UO_86 (O_86,N_24795,N_24982);
xor UO_87 (O_87,N_24999,N_24751);
or UO_88 (O_88,N_24851,N_24802);
or UO_89 (O_89,N_24986,N_24820);
nor UO_90 (O_90,N_24884,N_24984);
or UO_91 (O_91,N_24955,N_24842);
nor UO_92 (O_92,N_24916,N_24753);
nand UO_93 (O_93,N_24927,N_24913);
or UO_94 (O_94,N_24761,N_24983);
nand UO_95 (O_95,N_24951,N_24835);
nor UO_96 (O_96,N_24990,N_24934);
or UO_97 (O_97,N_24880,N_24989);
xor UO_98 (O_98,N_24816,N_24773);
nand UO_99 (O_99,N_24926,N_24892);
and UO_100 (O_100,N_24813,N_24998);
and UO_101 (O_101,N_24899,N_24865);
nand UO_102 (O_102,N_24954,N_24798);
xnor UO_103 (O_103,N_24801,N_24968);
nor UO_104 (O_104,N_24849,N_24807);
or UO_105 (O_105,N_24922,N_24858);
xor UO_106 (O_106,N_24874,N_24930);
nor UO_107 (O_107,N_24764,N_24949);
and UO_108 (O_108,N_24896,N_24834);
and UO_109 (O_109,N_24952,N_24940);
or UO_110 (O_110,N_24766,N_24777);
or UO_111 (O_111,N_24818,N_24894);
and UO_112 (O_112,N_24823,N_24960);
nor UO_113 (O_113,N_24805,N_24994);
or UO_114 (O_114,N_24933,N_24790);
or UO_115 (O_115,N_24836,N_24977);
and UO_116 (O_116,N_24995,N_24997);
and UO_117 (O_117,N_24859,N_24780);
and UO_118 (O_118,N_24967,N_24782);
nand UO_119 (O_119,N_24831,N_24963);
xor UO_120 (O_120,N_24839,N_24763);
nand UO_121 (O_121,N_24889,N_24893);
nand UO_122 (O_122,N_24905,N_24921);
nand UO_123 (O_123,N_24909,N_24917);
nor UO_124 (O_124,N_24804,N_24981);
nand UO_125 (O_125,N_24962,N_24882);
nor UO_126 (O_126,N_24978,N_24951);
nand UO_127 (O_127,N_24943,N_24817);
or UO_128 (O_128,N_24755,N_24945);
nand UO_129 (O_129,N_24823,N_24761);
xnor UO_130 (O_130,N_24818,N_24991);
or UO_131 (O_131,N_24897,N_24977);
nand UO_132 (O_132,N_24762,N_24919);
nor UO_133 (O_133,N_24758,N_24972);
and UO_134 (O_134,N_24941,N_24871);
or UO_135 (O_135,N_24827,N_24969);
nor UO_136 (O_136,N_24816,N_24791);
nand UO_137 (O_137,N_24798,N_24828);
nor UO_138 (O_138,N_24957,N_24828);
or UO_139 (O_139,N_24803,N_24758);
nand UO_140 (O_140,N_24798,N_24857);
nand UO_141 (O_141,N_24923,N_24981);
xor UO_142 (O_142,N_24889,N_24776);
nand UO_143 (O_143,N_24797,N_24793);
or UO_144 (O_144,N_24827,N_24798);
nand UO_145 (O_145,N_24772,N_24791);
and UO_146 (O_146,N_24813,N_24770);
nand UO_147 (O_147,N_24762,N_24752);
nor UO_148 (O_148,N_24933,N_24777);
and UO_149 (O_149,N_24951,N_24875);
and UO_150 (O_150,N_24931,N_24822);
xnor UO_151 (O_151,N_24922,N_24917);
or UO_152 (O_152,N_24775,N_24902);
and UO_153 (O_153,N_24800,N_24850);
nor UO_154 (O_154,N_24894,N_24954);
or UO_155 (O_155,N_24790,N_24849);
or UO_156 (O_156,N_24896,N_24849);
nor UO_157 (O_157,N_24785,N_24933);
and UO_158 (O_158,N_24833,N_24996);
nand UO_159 (O_159,N_24996,N_24877);
and UO_160 (O_160,N_24963,N_24771);
and UO_161 (O_161,N_24947,N_24991);
xor UO_162 (O_162,N_24952,N_24876);
xnor UO_163 (O_163,N_24777,N_24830);
nand UO_164 (O_164,N_24757,N_24821);
xnor UO_165 (O_165,N_24815,N_24867);
xor UO_166 (O_166,N_24977,N_24841);
nand UO_167 (O_167,N_24891,N_24840);
and UO_168 (O_168,N_24833,N_24976);
or UO_169 (O_169,N_24845,N_24907);
or UO_170 (O_170,N_24998,N_24948);
nor UO_171 (O_171,N_24855,N_24770);
nor UO_172 (O_172,N_24850,N_24766);
nand UO_173 (O_173,N_24970,N_24773);
and UO_174 (O_174,N_24784,N_24967);
xnor UO_175 (O_175,N_24823,N_24804);
nor UO_176 (O_176,N_24890,N_24895);
nor UO_177 (O_177,N_24760,N_24946);
nor UO_178 (O_178,N_24908,N_24871);
or UO_179 (O_179,N_24843,N_24824);
nor UO_180 (O_180,N_24788,N_24864);
xor UO_181 (O_181,N_24986,N_24839);
nor UO_182 (O_182,N_24844,N_24839);
nor UO_183 (O_183,N_24845,N_24850);
or UO_184 (O_184,N_24812,N_24988);
nor UO_185 (O_185,N_24772,N_24888);
and UO_186 (O_186,N_24949,N_24752);
nand UO_187 (O_187,N_24956,N_24929);
and UO_188 (O_188,N_24930,N_24836);
nand UO_189 (O_189,N_24981,N_24934);
nor UO_190 (O_190,N_24981,N_24762);
and UO_191 (O_191,N_24868,N_24768);
nor UO_192 (O_192,N_24922,N_24999);
nor UO_193 (O_193,N_24884,N_24806);
xor UO_194 (O_194,N_24893,N_24946);
and UO_195 (O_195,N_24755,N_24918);
or UO_196 (O_196,N_24827,N_24929);
or UO_197 (O_197,N_24772,N_24783);
and UO_198 (O_198,N_24913,N_24836);
or UO_199 (O_199,N_24977,N_24786);
and UO_200 (O_200,N_24851,N_24911);
and UO_201 (O_201,N_24780,N_24799);
and UO_202 (O_202,N_24842,N_24992);
nor UO_203 (O_203,N_24753,N_24960);
nor UO_204 (O_204,N_24851,N_24817);
or UO_205 (O_205,N_24982,N_24827);
and UO_206 (O_206,N_24849,N_24990);
xnor UO_207 (O_207,N_24878,N_24913);
and UO_208 (O_208,N_24837,N_24992);
and UO_209 (O_209,N_24825,N_24983);
nor UO_210 (O_210,N_24859,N_24752);
nand UO_211 (O_211,N_24868,N_24851);
or UO_212 (O_212,N_24983,N_24997);
and UO_213 (O_213,N_24804,N_24881);
or UO_214 (O_214,N_24918,N_24905);
and UO_215 (O_215,N_24853,N_24945);
and UO_216 (O_216,N_24760,N_24878);
nand UO_217 (O_217,N_24878,N_24875);
xnor UO_218 (O_218,N_24927,N_24835);
and UO_219 (O_219,N_24973,N_24879);
and UO_220 (O_220,N_24968,N_24897);
or UO_221 (O_221,N_24833,N_24883);
nand UO_222 (O_222,N_24751,N_24882);
xnor UO_223 (O_223,N_24921,N_24801);
xnor UO_224 (O_224,N_24955,N_24908);
or UO_225 (O_225,N_24774,N_24841);
or UO_226 (O_226,N_24942,N_24981);
and UO_227 (O_227,N_24760,N_24817);
or UO_228 (O_228,N_24843,N_24801);
and UO_229 (O_229,N_24839,N_24971);
and UO_230 (O_230,N_24818,N_24911);
or UO_231 (O_231,N_24834,N_24949);
or UO_232 (O_232,N_24968,N_24799);
nor UO_233 (O_233,N_24758,N_24750);
or UO_234 (O_234,N_24985,N_24803);
nand UO_235 (O_235,N_24769,N_24964);
or UO_236 (O_236,N_24788,N_24754);
or UO_237 (O_237,N_24931,N_24943);
or UO_238 (O_238,N_24994,N_24853);
nor UO_239 (O_239,N_24863,N_24882);
xnor UO_240 (O_240,N_24886,N_24881);
and UO_241 (O_241,N_24867,N_24988);
xor UO_242 (O_242,N_24887,N_24822);
nor UO_243 (O_243,N_24789,N_24986);
and UO_244 (O_244,N_24981,N_24956);
and UO_245 (O_245,N_24957,N_24905);
nand UO_246 (O_246,N_24840,N_24937);
nand UO_247 (O_247,N_24942,N_24784);
and UO_248 (O_248,N_24906,N_24785);
nand UO_249 (O_249,N_24824,N_24982);
xnor UO_250 (O_250,N_24887,N_24804);
and UO_251 (O_251,N_24811,N_24982);
nor UO_252 (O_252,N_24895,N_24910);
or UO_253 (O_253,N_24906,N_24916);
nand UO_254 (O_254,N_24925,N_24838);
nand UO_255 (O_255,N_24921,N_24785);
or UO_256 (O_256,N_24902,N_24921);
nand UO_257 (O_257,N_24986,N_24879);
nor UO_258 (O_258,N_24797,N_24952);
nand UO_259 (O_259,N_24825,N_24878);
or UO_260 (O_260,N_24777,N_24888);
or UO_261 (O_261,N_24796,N_24870);
or UO_262 (O_262,N_24881,N_24778);
xor UO_263 (O_263,N_24954,N_24855);
nand UO_264 (O_264,N_24790,N_24929);
and UO_265 (O_265,N_24896,N_24932);
nand UO_266 (O_266,N_24895,N_24952);
and UO_267 (O_267,N_24950,N_24891);
nor UO_268 (O_268,N_24772,N_24867);
or UO_269 (O_269,N_24952,N_24824);
nor UO_270 (O_270,N_24855,N_24934);
nand UO_271 (O_271,N_24836,N_24831);
nor UO_272 (O_272,N_24799,N_24935);
nand UO_273 (O_273,N_24974,N_24924);
and UO_274 (O_274,N_24986,N_24817);
nand UO_275 (O_275,N_24996,N_24900);
or UO_276 (O_276,N_24949,N_24974);
nand UO_277 (O_277,N_24999,N_24987);
or UO_278 (O_278,N_24927,N_24977);
and UO_279 (O_279,N_24885,N_24945);
nor UO_280 (O_280,N_24982,N_24820);
nand UO_281 (O_281,N_24933,N_24750);
nand UO_282 (O_282,N_24834,N_24782);
nand UO_283 (O_283,N_24987,N_24942);
and UO_284 (O_284,N_24871,N_24828);
xor UO_285 (O_285,N_24792,N_24941);
or UO_286 (O_286,N_24835,N_24924);
xor UO_287 (O_287,N_24830,N_24891);
or UO_288 (O_288,N_24812,N_24979);
nand UO_289 (O_289,N_24794,N_24960);
nand UO_290 (O_290,N_24935,N_24824);
and UO_291 (O_291,N_24772,N_24828);
and UO_292 (O_292,N_24778,N_24860);
nand UO_293 (O_293,N_24765,N_24809);
nor UO_294 (O_294,N_24906,N_24753);
nand UO_295 (O_295,N_24877,N_24870);
or UO_296 (O_296,N_24950,N_24990);
nor UO_297 (O_297,N_24810,N_24796);
nand UO_298 (O_298,N_24927,N_24803);
and UO_299 (O_299,N_24948,N_24964);
or UO_300 (O_300,N_24867,N_24790);
nor UO_301 (O_301,N_24879,N_24821);
nand UO_302 (O_302,N_24980,N_24914);
or UO_303 (O_303,N_24851,N_24844);
nor UO_304 (O_304,N_24918,N_24903);
and UO_305 (O_305,N_24823,N_24810);
nor UO_306 (O_306,N_24907,N_24820);
xnor UO_307 (O_307,N_24902,N_24768);
nor UO_308 (O_308,N_24934,N_24800);
nand UO_309 (O_309,N_24902,N_24988);
xor UO_310 (O_310,N_24922,N_24981);
and UO_311 (O_311,N_24984,N_24898);
or UO_312 (O_312,N_24927,N_24992);
nand UO_313 (O_313,N_24914,N_24978);
or UO_314 (O_314,N_24964,N_24987);
nor UO_315 (O_315,N_24784,N_24999);
nand UO_316 (O_316,N_24961,N_24919);
nor UO_317 (O_317,N_24808,N_24854);
nor UO_318 (O_318,N_24985,N_24759);
nor UO_319 (O_319,N_24933,N_24900);
and UO_320 (O_320,N_24999,N_24973);
and UO_321 (O_321,N_24968,N_24843);
nor UO_322 (O_322,N_24778,N_24837);
and UO_323 (O_323,N_24780,N_24916);
nand UO_324 (O_324,N_24965,N_24826);
nor UO_325 (O_325,N_24802,N_24825);
nand UO_326 (O_326,N_24761,N_24758);
nor UO_327 (O_327,N_24798,N_24841);
and UO_328 (O_328,N_24998,N_24910);
nor UO_329 (O_329,N_24780,N_24912);
and UO_330 (O_330,N_24778,N_24993);
nand UO_331 (O_331,N_24993,N_24927);
and UO_332 (O_332,N_24856,N_24841);
or UO_333 (O_333,N_24806,N_24935);
or UO_334 (O_334,N_24844,N_24774);
or UO_335 (O_335,N_24882,N_24979);
nor UO_336 (O_336,N_24926,N_24805);
nor UO_337 (O_337,N_24850,N_24914);
or UO_338 (O_338,N_24789,N_24773);
or UO_339 (O_339,N_24814,N_24778);
xnor UO_340 (O_340,N_24961,N_24992);
and UO_341 (O_341,N_24824,N_24822);
and UO_342 (O_342,N_24920,N_24998);
or UO_343 (O_343,N_24956,N_24906);
nand UO_344 (O_344,N_24969,N_24852);
xnor UO_345 (O_345,N_24764,N_24852);
nand UO_346 (O_346,N_24802,N_24801);
nand UO_347 (O_347,N_24776,N_24924);
nand UO_348 (O_348,N_24886,N_24946);
or UO_349 (O_349,N_24814,N_24962);
nand UO_350 (O_350,N_24865,N_24819);
nand UO_351 (O_351,N_24823,N_24988);
xor UO_352 (O_352,N_24884,N_24809);
or UO_353 (O_353,N_24996,N_24848);
nor UO_354 (O_354,N_24789,N_24904);
nand UO_355 (O_355,N_24953,N_24763);
nor UO_356 (O_356,N_24787,N_24878);
or UO_357 (O_357,N_24775,N_24977);
nand UO_358 (O_358,N_24944,N_24953);
nor UO_359 (O_359,N_24840,N_24905);
nand UO_360 (O_360,N_24868,N_24923);
nand UO_361 (O_361,N_24893,N_24856);
nor UO_362 (O_362,N_24925,N_24774);
and UO_363 (O_363,N_24784,N_24896);
nand UO_364 (O_364,N_24940,N_24873);
or UO_365 (O_365,N_24999,N_24863);
nand UO_366 (O_366,N_24903,N_24819);
nor UO_367 (O_367,N_24794,N_24918);
or UO_368 (O_368,N_24958,N_24971);
nor UO_369 (O_369,N_24960,N_24925);
or UO_370 (O_370,N_24779,N_24966);
and UO_371 (O_371,N_24832,N_24886);
nand UO_372 (O_372,N_24945,N_24929);
nand UO_373 (O_373,N_24753,N_24975);
nand UO_374 (O_374,N_24797,N_24794);
nor UO_375 (O_375,N_24834,N_24859);
and UO_376 (O_376,N_24957,N_24813);
or UO_377 (O_377,N_24755,N_24881);
or UO_378 (O_378,N_24758,N_24935);
nand UO_379 (O_379,N_24930,N_24834);
nand UO_380 (O_380,N_24811,N_24855);
and UO_381 (O_381,N_24899,N_24971);
and UO_382 (O_382,N_24918,N_24753);
or UO_383 (O_383,N_24867,N_24886);
nor UO_384 (O_384,N_24998,N_24982);
or UO_385 (O_385,N_24988,N_24761);
or UO_386 (O_386,N_24802,N_24949);
nand UO_387 (O_387,N_24764,N_24930);
nor UO_388 (O_388,N_24819,N_24765);
xnor UO_389 (O_389,N_24752,N_24959);
nand UO_390 (O_390,N_24774,N_24897);
nor UO_391 (O_391,N_24780,N_24965);
nand UO_392 (O_392,N_24770,N_24939);
nor UO_393 (O_393,N_24954,N_24869);
nand UO_394 (O_394,N_24777,N_24882);
xor UO_395 (O_395,N_24840,N_24832);
or UO_396 (O_396,N_24774,N_24975);
nand UO_397 (O_397,N_24862,N_24750);
nand UO_398 (O_398,N_24908,N_24802);
nor UO_399 (O_399,N_24762,N_24852);
and UO_400 (O_400,N_24949,N_24890);
xnor UO_401 (O_401,N_24843,N_24859);
xor UO_402 (O_402,N_24806,N_24783);
nor UO_403 (O_403,N_24772,N_24864);
nor UO_404 (O_404,N_24911,N_24839);
and UO_405 (O_405,N_24829,N_24858);
nand UO_406 (O_406,N_24804,N_24839);
or UO_407 (O_407,N_24924,N_24936);
nor UO_408 (O_408,N_24987,N_24761);
nand UO_409 (O_409,N_24912,N_24963);
nand UO_410 (O_410,N_24860,N_24885);
xnor UO_411 (O_411,N_24912,N_24988);
nand UO_412 (O_412,N_24819,N_24894);
and UO_413 (O_413,N_24962,N_24911);
nor UO_414 (O_414,N_24976,N_24885);
and UO_415 (O_415,N_24993,N_24785);
and UO_416 (O_416,N_24918,N_24893);
and UO_417 (O_417,N_24781,N_24839);
and UO_418 (O_418,N_24755,N_24769);
and UO_419 (O_419,N_24892,N_24976);
nand UO_420 (O_420,N_24859,N_24903);
nand UO_421 (O_421,N_24770,N_24772);
or UO_422 (O_422,N_24848,N_24959);
and UO_423 (O_423,N_24799,N_24897);
xor UO_424 (O_424,N_24928,N_24839);
and UO_425 (O_425,N_24862,N_24967);
nor UO_426 (O_426,N_24958,N_24875);
nor UO_427 (O_427,N_24913,N_24767);
xnor UO_428 (O_428,N_24965,N_24854);
and UO_429 (O_429,N_24951,N_24853);
and UO_430 (O_430,N_24907,N_24763);
or UO_431 (O_431,N_24791,N_24811);
nor UO_432 (O_432,N_24994,N_24910);
nand UO_433 (O_433,N_24977,N_24826);
xnor UO_434 (O_434,N_24966,N_24983);
nor UO_435 (O_435,N_24953,N_24910);
or UO_436 (O_436,N_24776,N_24874);
or UO_437 (O_437,N_24940,N_24844);
nand UO_438 (O_438,N_24999,N_24986);
nor UO_439 (O_439,N_24896,N_24973);
nor UO_440 (O_440,N_24989,N_24915);
nor UO_441 (O_441,N_24773,N_24828);
nor UO_442 (O_442,N_24987,N_24904);
xor UO_443 (O_443,N_24916,N_24875);
xnor UO_444 (O_444,N_24824,N_24902);
nand UO_445 (O_445,N_24950,N_24803);
and UO_446 (O_446,N_24988,N_24783);
and UO_447 (O_447,N_24822,N_24961);
nand UO_448 (O_448,N_24839,N_24917);
nand UO_449 (O_449,N_24783,N_24902);
nor UO_450 (O_450,N_24938,N_24813);
or UO_451 (O_451,N_24936,N_24773);
nor UO_452 (O_452,N_24790,N_24783);
nor UO_453 (O_453,N_24825,N_24971);
and UO_454 (O_454,N_24912,N_24959);
xnor UO_455 (O_455,N_24835,N_24752);
and UO_456 (O_456,N_24929,N_24992);
xor UO_457 (O_457,N_24778,N_24826);
xor UO_458 (O_458,N_24863,N_24830);
and UO_459 (O_459,N_24961,N_24827);
and UO_460 (O_460,N_24814,N_24849);
or UO_461 (O_461,N_24972,N_24946);
or UO_462 (O_462,N_24916,N_24940);
or UO_463 (O_463,N_24903,N_24824);
nand UO_464 (O_464,N_24856,N_24770);
or UO_465 (O_465,N_24844,N_24953);
and UO_466 (O_466,N_24979,N_24854);
and UO_467 (O_467,N_24836,N_24957);
or UO_468 (O_468,N_24974,N_24945);
and UO_469 (O_469,N_24766,N_24803);
and UO_470 (O_470,N_24866,N_24992);
xor UO_471 (O_471,N_24755,N_24929);
and UO_472 (O_472,N_24776,N_24984);
nor UO_473 (O_473,N_24983,N_24869);
or UO_474 (O_474,N_24908,N_24879);
and UO_475 (O_475,N_24904,N_24963);
or UO_476 (O_476,N_24824,N_24752);
nand UO_477 (O_477,N_24802,N_24866);
and UO_478 (O_478,N_24759,N_24940);
and UO_479 (O_479,N_24759,N_24988);
nor UO_480 (O_480,N_24999,N_24982);
nor UO_481 (O_481,N_24862,N_24898);
nor UO_482 (O_482,N_24949,N_24793);
and UO_483 (O_483,N_24977,N_24929);
nand UO_484 (O_484,N_24993,N_24872);
nor UO_485 (O_485,N_24771,N_24986);
and UO_486 (O_486,N_24830,N_24857);
or UO_487 (O_487,N_24839,N_24955);
nand UO_488 (O_488,N_24901,N_24835);
xor UO_489 (O_489,N_24997,N_24791);
xnor UO_490 (O_490,N_24980,N_24986);
nand UO_491 (O_491,N_24843,N_24948);
nor UO_492 (O_492,N_24903,N_24897);
nand UO_493 (O_493,N_24825,N_24866);
or UO_494 (O_494,N_24929,N_24797);
and UO_495 (O_495,N_24876,N_24809);
or UO_496 (O_496,N_24830,N_24852);
and UO_497 (O_497,N_24991,N_24848);
nor UO_498 (O_498,N_24863,N_24906);
xnor UO_499 (O_499,N_24804,N_24816);
nand UO_500 (O_500,N_24785,N_24931);
or UO_501 (O_501,N_24769,N_24806);
and UO_502 (O_502,N_24975,N_24795);
or UO_503 (O_503,N_24750,N_24932);
nor UO_504 (O_504,N_24828,N_24946);
and UO_505 (O_505,N_24808,N_24772);
or UO_506 (O_506,N_24751,N_24750);
nand UO_507 (O_507,N_24754,N_24752);
xor UO_508 (O_508,N_24825,N_24831);
or UO_509 (O_509,N_24962,N_24957);
nand UO_510 (O_510,N_24957,N_24942);
or UO_511 (O_511,N_24986,N_24772);
or UO_512 (O_512,N_24877,N_24864);
or UO_513 (O_513,N_24931,N_24938);
nand UO_514 (O_514,N_24983,N_24828);
and UO_515 (O_515,N_24892,N_24854);
nand UO_516 (O_516,N_24891,N_24964);
or UO_517 (O_517,N_24779,N_24988);
nor UO_518 (O_518,N_24915,N_24890);
nor UO_519 (O_519,N_24971,N_24906);
or UO_520 (O_520,N_24926,N_24867);
nand UO_521 (O_521,N_24798,N_24790);
nand UO_522 (O_522,N_24978,N_24952);
nand UO_523 (O_523,N_24801,N_24764);
and UO_524 (O_524,N_24950,N_24954);
or UO_525 (O_525,N_24874,N_24918);
nor UO_526 (O_526,N_24779,N_24879);
and UO_527 (O_527,N_24969,N_24924);
or UO_528 (O_528,N_24835,N_24957);
or UO_529 (O_529,N_24938,N_24898);
nor UO_530 (O_530,N_24992,N_24770);
nand UO_531 (O_531,N_24985,N_24927);
nand UO_532 (O_532,N_24756,N_24814);
or UO_533 (O_533,N_24755,N_24927);
or UO_534 (O_534,N_24974,N_24842);
or UO_535 (O_535,N_24895,N_24861);
and UO_536 (O_536,N_24971,N_24781);
xnor UO_537 (O_537,N_24991,N_24892);
nor UO_538 (O_538,N_24959,N_24751);
nand UO_539 (O_539,N_24784,N_24880);
nor UO_540 (O_540,N_24949,N_24851);
or UO_541 (O_541,N_24851,N_24833);
and UO_542 (O_542,N_24957,N_24838);
nand UO_543 (O_543,N_24885,N_24880);
nor UO_544 (O_544,N_24793,N_24826);
or UO_545 (O_545,N_24991,N_24890);
and UO_546 (O_546,N_24817,N_24898);
nor UO_547 (O_547,N_24863,N_24778);
or UO_548 (O_548,N_24765,N_24878);
or UO_549 (O_549,N_24879,N_24859);
and UO_550 (O_550,N_24764,N_24980);
nand UO_551 (O_551,N_24897,N_24805);
nor UO_552 (O_552,N_24959,N_24923);
or UO_553 (O_553,N_24758,N_24782);
xor UO_554 (O_554,N_24775,N_24790);
or UO_555 (O_555,N_24980,N_24873);
nor UO_556 (O_556,N_24887,N_24798);
or UO_557 (O_557,N_24816,N_24886);
or UO_558 (O_558,N_24795,N_24787);
or UO_559 (O_559,N_24752,N_24944);
nor UO_560 (O_560,N_24766,N_24783);
nor UO_561 (O_561,N_24800,N_24977);
and UO_562 (O_562,N_24933,N_24854);
or UO_563 (O_563,N_24939,N_24763);
or UO_564 (O_564,N_24911,N_24885);
nand UO_565 (O_565,N_24791,N_24809);
or UO_566 (O_566,N_24925,N_24755);
nand UO_567 (O_567,N_24820,N_24873);
nor UO_568 (O_568,N_24836,N_24807);
nand UO_569 (O_569,N_24997,N_24902);
nand UO_570 (O_570,N_24874,N_24892);
nor UO_571 (O_571,N_24818,N_24773);
and UO_572 (O_572,N_24991,N_24978);
nand UO_573 (O_573,N_24977,N_24855);
nand UO_574 (O_574,N_24944,N_24928);
nand UO_575 (O_575,N_24946,N_24897);
nand UO_576 (O_576,N_24774,N_24796);
nor UO_577 (O_577,N_24834,N_24952);
and UO_578 (O_578,N_24803,N_24761);
or UO_579 (O_579,N_24878,N_24911);
nand UO_580 (O_580,N_24927,N_24953);
and UO_581 (O_581,N_24966,N_24783);
nand UO_582 (O_582,N_24799,N_24765);
and UO_583 (O_583,N_24802,N_24915);
nand UO_584 (O_584,N_24974,N_24844);
or UO_585 (O_585,N_24982,N_24976);
nand UO_586 (O_586,N_24779,N_24921);
or UO_587 (O_587,N_24930,N_24996);
or UO_588 (O_588,N_24892,N_24973);
and UO_589 (O_589,N_24843,N_24762);
nand UO_590 (O_590,N_24834,N_24923);
xnor UO_591 (O_591,N_24779,N_24915);
and UO_592 (O_592,N_24829,N_24911);
nor UO_593 (O_593,N_24969,N_24765);
or UO_594 (O_594,N_24886,N_24897);
nor UO_595 (O_595,N_24856,N_24948);
nand UO_596 (O_596,N_24850,N_24806);
and UO_597 (O_597,N_24874,N_24885);
nand UO_598 (O_598,N_24826,N_24970);
nand UO_599 (O_599,N_24811,N_24920);
nor UO_600 (O_600,N_24797,N_24906);
and UO_601 (O_601,N_24762,N_24833);
and UO_602 (O_602,N_24880,N_24994);
nand UO_603 (O_603,N_24759,N_24815);
nand UO_604 (O_604,N_24974,N_24992);
nand UO_605 (O_605,N_24952,N_24827);
xor UO_606 (O_606,N_24991,N_24846);
nor UO_607 (O_607,N_24995,N_24931);
xnor UO_608 (O_608,N_24767,N_24991);
nand UO_609 (O_609,N_24885,N_24952);
nand UO_610 (O_610,N_24982,N_24752);
and UO_611 (O_611,N_24826,N_24851);
nor UO_612 (O_612,N_24860,N_24976);
nor UO_613 (O_613,N_24912,N_24936);
nand UO_614 (O_614,N_24872,N_24836);
and UO_615 (O_615,N_24845,N_24809);
or UO_616 (O_616,N_24974,N_24896);
nand UO_617 (O_617,N_24939,N_24914);
nand UO_618 (O_618,N_24812,N_24874);
and UO_619 (O_619,N_24915,N_24835);
and UO_620 (O_620,N_24916,N_24800);
nor UO_621 (O_621,N_24906,N_24945);
or UO_622 (O_622,N_24850,N_24842);
nand UO_623 (O_623,N_24805,N_24780);
nor UO_624 (O_624,N_24840,N_24848);
nor UO_625 (O_625,N_24763,N_24913);
nand UO_626 (O_626,N_24920,N_24952);
nor UO_627 (O_627,N_24996,N_24898);
and UO_628 (O_628,N_24965,N_24814);
or UO_629 (O_629,N_24995,N_24973);
nor UO_630 (O_630,N_24908,N_24834);
nor UO_631 (O_631,N_24921,N_24792);
nand UO_632 (O_632,N_24881,N_24871);
or UO_633 (O_633,N_24990,N_24884);
nor UO_634 (O_634,N_24793,N_24866);
xnor UO_635 (O_635,N_24811,N_24974);
and UO_636 (O_636,N_24794,N_24945);
xor UO_637 (O_637,N_24939,N_24970);
nand UO_638 (O_638,N_24936,N_24767);
or UO_639 (O_639,N_24772,N_24769);
nand UO_640 (O_640,N_24901,N_24777);
nor UO_641 (O_641,N_24889,N_24935);
or UO_642 (O_642,N_24756,N_24882);
nor UO_643 (O_643,N_24911,N_24802);
or UO_644 (O_644,N_24881,N_24927);
and UO_645 (O_645,N_24903,N_24961);
nor UO_646 (O_646,N_24844,N_24983);
and UO_647 (O_647,N_24788,N_24914);
or UO_648 (O_648,N_24880,N_24865);
nor UO_649 (O_649,N_24959,N_24824);
and UO_650 (O_650,N_24904,N_24942);
and UO_651 (O_651,N_24816,N_24974);
or UO_652 (O_652,N_24835,N_24922);
or UO_653 (O_653,N_24991,N_24966);
nand UO_654 (O_654,N_24895,N_24915);
xor UO_655 (O_655,N_24960,N_24848);
nor UO_656 (O_656,N_24782,N_24801);
and UO_657 (O_657,N_24972,N_24887);
xnor UO_658 (O_658,N_24908,N_24827);
nand UO_659 (O_659,N_24999,N_24779);
nor UO_660 (O_660,N_24839,N_24871);
or UO_661 (O_661,N_24848,N_24835);
and UO_662 (O_662,N_24973,N_24838);
and UO_663 (O_663,N_24996,N_24835);
or UO_664 (O_664,N_24921,N_24989);
nand UO_665 (O_665,N_24769,N_24818);
xor UO_666 (O_666,N_24902,N_24779);
xor UO_667 (O_667,N_24853,N_24818);
or UO_668 (O_668,N_24915,N_24919);
or UO_669 (O_669,N_24879,N_24776);
nor UO_670 (O_670,N_24905,N_24963);
and UO_671 (O_671,N_24873,N_24917);
nor UO_672 (O_672,N_24936,N_24958);
and UO_673 (O_673,N_24899,N_24883);
or UO_674 (O_674,N_24884,N_24818);
nand UO_675 (O_675,N_24975,N_24948);
or UO_676 (O_676,N_24806,N_24764);
nand UO_677 (O_677,N_24884,N_24980);
nand UO_678 (O_678,N_24856,N_24855);
nand UO_679 (O_679,N_24992,N_24884);
nor UO_680 (O_680,N_24759,N_24904);
or UO_681 (O_681,N_24771,N_24778);
nand UO_682 (O_682,N_24836,N_24762);
nor UO_683 (O_683,N_24952,N_24753);
nor UO_684 (O_684,N_24947,N_24974);
and UO_685 (O_685,N_24778,N_24945);
nand UO_686 (O_686,N_24943,N_24929);
nand UO_687 (O_687,N_24782,N_24750);
and UO_688 (O_688,N_24957,N_24953);
and UO_689 (O_689,N_24988,N_24995);
nand UO_690 (O_690,N_24924,N_24754);
nand UO_691 (O_691,N_24775,N_24845);
nor UO_692 (O_692,N_24953,N_24773);
or UO_693 (O_693,N_24933,N_24973);
or UO_694 (O_694,N_24764,N_24866);
or UO_695 (O_695,N_24886,N_24871);
or UO_696 (O_696,N_24784,N_24865);
nand UO_697 (O_697,N_24834,N_24802);
nor UO_698 (O_698,N_24941,N_24894);
nor UO_699 (O_699,N_24883,N_24994);
nand UO_700 (O_700,N_24802,N_24870);
and UO_701 (O_701,N_24918,N_24987);
nand UO_702 (O_702,N_24827,N_24820);
and UO_703 (O_703,N_24828,N_24872);
nor UO_704 (O_704,N_24912,N_24923);
or UO_705 (O_705,N_24860,N_24982);
nor UO_706 (O_706,N_24757,N_24932);
nand UO_707 (O_707,N_24838,N_24862);
and UO_708 (O_708,N_24960,N_24890);
nor UO_709 (O_709,N_24773,N_24998);
or UO_710 (O_710,N_24962,N_24884);
nand UO_711 (O_711,N_24808,N_24886);
nand UO_712 (O_712,N_24981,N_24897);
and UO_713 (O_713,N_24977,N_24891);
xnor UO_714 (O_714,N_24770,N_24980);
and UO_715 (O_715,N_24788,N_24814);
and UO_716 (O_716,N_24771,N_24799);
nand UO_717 (O_717,N_24791,N_24755);
nor UO_718 (O_718,N_24818,N_24919);
or UO_719 (O_719,N_24846,N_24803);
and UO_720 (O_720,N_24827,N_24847);
nand UO_721 (O_721,N_24805,N_24800);
or UO_722 (O_722,N_24774,N_24846);
or UO_723 (O_723,N_24893,N_24759);
or UO_724 (O_724,N_24926,N_24782);
nor UO_725 (O_725,N_24867,N_24972);
nor UO_726 (O_726,N_24844,N_24990);
or UO_727 (O_727,N_24958,N_24887);
nand UO_728 (O_728,N_24813,N_24917);
nor UO_729 (O_729,N_24863,N_24847);
and UO_730 (O_730,N_24857,N_24913);
and UO_731 (O_731,N_24963,N_24779);
or UO_732 (O_732,N_24887,N_24977);
and UO_733 (O_733,N_24935,N_24922);
xnor UO_734 (O_734,N_24989,N_24869);
or UO_735 (O_735,N_24763,N_24835);
xor UO_736 (O_736,N_24883,N_24916);
xor UO_737 (O_737,N_24982,N_24840);
and UO_738 (O_738,N_24889,N_24833);
or UO_739 (O_739,N_24801,N_24856);
xor UO_740 (O_740,N_24990,N_24772);
xnor UO_741 (O_741,N_24775,N_24791);
nand UO_742 (O_742,N_24764,N_24904);
and UO_743 (O_743,N_24922,N_24852);
xnor UO_744 (O_744,N_24893,N_24798);
and UO_745 (O_745,N_24975,N_24982);
nand UO_746 (O_746,N_24812,N_24754);
nor UO_747 (O_747,N_24786,N_24956);
and UO_748 (O_748,N_24983,N_24808);
nand UO_749 (O_749,N_24969,N_24867);
nand UO_750 (O_750,N_24817,N_24891);
nor UO_751 (O_751,N_24975,N_24998);
or UO_752 (O_752,N_24902,N_24876);
and UO_753 (O_753,N_24792,N_24903);
nor UO_754 (O_754,N_24853,N_24829);
xor UO_755 (O_755,N_24938,N_24990);
and UO_756 (O_756,N_24801,N_24963);
nor UO_757 (O_757,N_24922,N_24842);
or UO_758 (O_758,N_24799,N_24793);
and UO_759 (O_759,N_24966,N_24871);
nand UO_760 (O_760,N_24961,N_24982);
nand UO_761 (O_761,N_24889,N_24969);
nor UO_762 (O_762,N_24968,N_24977);
nand UO_763 (O_763,N_24778,N_24750);
nor UO_764 (O_764,N_24850,N_24946);
nand UO_765 (O_765,N_24871,N_24752);
nand UO_766 (O_766,N_24790,N_24912);
nor UO_767 (O_767,N_24989,N_24761);
xor UO_768 (O_768,N_24977,N_24923);
and UO_769 (O_769,N_24923,N_24836);
nand UO_770 (O_770,N_24978,N_24811);
xor UO_771 (O_771,N_24916,N_24761);
or UO_772 (O_772,N_24919,N_24997);
and UO_773 (O_773,N_24817,N_24755);
nand UO_774 (O_774,N_24801,N_24837);
nand UO_775 (O_775,N_24954,N_24860);
nand UO_776 (O_776,N_24881,N_24964);
xor UO_777 (O_777,N_24796,N_24925);
and UO_778 (O_778,N_24752,N_24805);
nor UO_779 (O_779,N_24850,N_24982);
nor UO_780 (O_780,N_24932,N_24939);
and UO_781 (O_781,N_24893,N_24756);
nand UO_782 (O_782,N_24885,N_24918);
or UO_783 (O_783,N_24851,N_24846);
nor UO_784 (O_784,N_24885,N_24940);
nor UO_785 (O_785,N_24958,N_24869);
or UO_786 (O_786,N_24875,N_24818);
nand UO_787 (O_787,N_24837,N_24932);
nand UO_788 (O_788,N_24864,N_24758);
or UO_789 (O_789,N_24906,N_24966);
nor UO_790 (O_790,N_24931,N_24919);
and UO_791 (O_791,N_24761,N_24869);
xnor UO_792 (O_792,N_24933,N_24951);
nor UO_793 (O_793,N_24945,N_24951);
and UO_794 (O_794,N_24899,N_24930);
nor UO_795 (O_795,N_24996,N_24768);
xor UO_796 (O_796,N_24899,N_24945);
nor UO_797 (O_797,N_24845,N_24928);
xnor UO_798 (O_798,N_24953,N_24764);
nand UO_799 (O_799,N_24929,N_24780);
nor UO_800 (O_800,N_24914,N_24845);
nand UO_801 (O_801,N_24849,N_24784);
and UO_802 (O_802,N_24839,N_24877);
or UO_803 (O_803,N_24999,N_24839);
xnor UO_804 (O_804,N_24899,N_24803);
and UO_805 (O_805,N_24921,N_24811);
and UO_806 (O_806,N_24899,N_24752);
or UO_807 (O_807,N_24880,N_24943);
nor UO_808 (O_808,N_24848,N_24875);
or UO_809 (O_809,N_24945,N_24954);
or UO_810 (O_810,N_24953,N_24880);
nand UO_811 (O_811,N_24884,N_24897);
nand UO_812 (O_812,N_24859,N_24810);
or UO_813 (O_813,N_24767,N_24929);
or UO_814 (O_814,N_24821,N_24870);
nand UO_815 (O_815,N_24761,N_24867);
and UO_816 (O_816,N_24917,N_24916);
nand UO_817 (O_817,N_24852,N_24944);
and UO_818 (O_818,N_24969,N_24830);
nor UO_819 (O_819,N_24989,N_24801);
and UO_820 (O_820,N_24827,N_24850);
and UO_821 (O_821,N_24847,N_24933);
and UO_822 (O_822,N_24944,N_24850);
or UO_823 (O_823,N_24942,N_24802);
nand UO_824 (O_824,N_24925,N_24894);
nor UO_825 (O_825,N_24831,N_24851);
and UO_826 (O_826,N_24918,N_24989);
and UO_827 (O_827,N_24797,N_24835);
nand UO_828 (O_828,N_24846,N_24752);
nand UO_829 (O_829,N_24972,N_24808);
xor UO_830 (O_830,N_24801,N_24795);
nor UO_831 (O_831,N_24954,N_24842);
xnor UO_832 (O_832,N_24851,N_24867);
or UO_833 (O_833,N_24955,N_24780);
nand UO_834 (O_834,N_24861,N_24934);
and UO_835 (O_835,N_24923,N_24918);
nor UO_836 (O_836,N_24958,N_24931);
or UO_837 (O_837,N_24995,N_24920);
or UO_838 (O_838,N_24826,N_24998);
xnor UO_839 (O_839,N_24821,N_24909);
and UO_840 (O_840,N_24883,N_24776);
and UO_841 (O_841,N_24798,N_24797);
and UO_842 (O_842,N_24806,N_24925);
nand UO_843 (O_843,N_24814,N_24817);
nand UO_844 (O_844,N_24944,N_24835);
and UO_845 (O_845,N_24864,N_24824);
and UO_846 (O_846,N_24929,N_24942);
nor UO_847 (O_847,N_24889,N_24873);
or UO_848 (O_848,N_24775,N_24947);
xor UO_849 (O_849,N_24962,N_24989);
and UO_850 (O_850,N_24883,N_24751);
or UO_851 (O_851,N_24936,N_24858);
and UO_852 (O_852,N_24869,N_24764);
or UO_853 (O_853,N_24954,N_24837);
or UO_854 (O_854,N_24940,N_24843);
nand UO_855 (O_855,N_24754,N_24785);
or UO_856 (O_856,N_24871,N_24784);
or UO_857 (O_857,N_24785,N_24868);
and UO_858 (O_858,N_24964,N_24787);
and UO_859 (O_859,N_24942,N_24881);
nand UO_860 (O_860,N_24793,N_24818);
nor UO_861 (O_861,N_24815,N_24881);
and UO_862 (O_862,N_24906,N_24937);
xor UO_863 (O_863,N_24756,N_24800);
or UO_864 (O_864,N_24971,N_24826);
nor UO_865 (O_865,N_24975,N_24757);
and UO_866 (O_866,N_24862,N_24773);
or UO_867 (O_867,N_24776,N_24830);
nand UO_868 (O_868,N_24952,N_24836);
nand UO_869 (O_869,N_24823,N_24947);
and UO_870 (O_870,N_24926,N_24857);
xor UO_871 (O_871,N_24817,N_24960);
or UO_872 (O_872,N_24765,N_24839);
nand UO_873 (O_873,N_24955,N_24894);
or UO_874 (O_874,N_24885,N_24855);
nand UO_875 (O_875,N_24762,N_24834);
nor UO_876 (O_876,N_24782,N_24772);
and UO_877 (O_877,N_24800,N_24821);
nand UO_878 (O_878,N_24982,N_24927);
xor UO_879 (O_879,N_24841,N_24819);
or UO_880 (O_880,N_24990,N_24752);
nor UO_881 (O_881,N_24980,N_24781);
nor UO_882 (O_882,N_24951,N_24834);
or UO_883 (O_883,N_24969,N_24829);
or UO_884 (O_884,N_24883,N_24761);
or UO_885 (O_885,N_24790,N_24752);
nor UO_886 (O_886,N_24930,N_24965);
xor UO_887 (O_887,N_24849,N_24968);
nor UO_888 (O_888,N_24809,N_24928);
nor UO_889 (O_889,N_24851,N_24996);
nor UO_890 (O_890,N_24944,N_24894);
nor UO_891 (O_891,N_24784,N_24866);
nand UO_892 (O_892,N_24782,N_24756);
nor UO_893 (O_893,N_24859,N_24899);
nand UO_894 (O_894,N_24952,N_24926);
and UO_895 (O_895,N_24918,N_24847);
and UO_896 (O_896,N_24854,N_24793);
nand UO_897 (O_897,N_24959,N_24845);
and UO_898 (O_898,N_24918,N_24882);
nand UO_899 (O_899,N_24860,N_24798);
nor UO_900 (O_900,N_24921,N_24818);
and UO_901 (O_901,N_24840,N_24833);
and UO_902 (O_902,N_24857,N_24935);
nor UO_903 (O_903,N_24753,N_24930);
nor UO_904 (O_904,N_24772,N_24928);
nand UO_905 (O_905,N_24978,N_24797);
and UO_906 (O_906,N_24931,N_24991);
xnor UO_907 (O_907,N_24958,N_24799);
nor UO_908 (O_908,N_24923,N_24797);
or UO_909 (O_909,N_24793,N_24845);
nand UO_910 (O_910,N_24812,N_24791);
nand UO_911 (O_911,N_24825,N_24771);
and UO_912 (O_912,N_24781,N_24770);
nand UO_913 (O_913,N_24850,N_24992);
and UO_914 (O_914,N_24763,N_24997);
or UO_915 (O_915,N_24805,N_24758);
nor UO_916 (O_916,N_24868,N_24967);
or UO_917 (O_917,N_24832,N_24941);
and UO_918 (O_918,N_24989,N_24902);
nor UO_919 (O_919,N_24862,N_24830);
xnor UO_920 (O_920,N_24847,N_24824);
and UO_921 (O_921,N_24882,N_24899);
nor UO_922 (O_922,N_24883,N_24842);
nand UO_923 (O_923,N_24953,N_24937);
nor UO_924 (O_924,N_24983,N_24933);
or UO_925 (O_925,N_24823,N_24932);
or UO_926 (O_926,N_24807,N_24863);
nor UO_927 (O_927,N_24919,N_24801);
xor UO_928 (O_928,N_24981,N_24938);
nor UO_929 (O_929,N_24828,N_24970);
and UO_930 (O_930,N_24987,N_24864);
and UO_931 (O_931,N_24983,N_24753);
nor UO_932 (O_932,N_24918,N_24968);
nand UO_933 (O_933,N_24983,N_24879);
nor UO_934 (O_934,N_24766,N_24902);
nor UO_935 (O_935,N_24869,N_24775);
nor UO_936 (O_936,N_24971,N_24806);
or UO_937 (O_937,N_24938,N_24753);
and UO_938 (O_938,N_24984,N_24902);
or UO_939 (O_939,N_24931,N_24750);
and UO_940 (O_940,N_24784,N_24969);
or UO_941 (O_941,N_24995,N_24784);
nand UO_942 (O_942,N_24875,N_24901);
or UO_943 (O_943,N_24858,N_24854);
nand UO_944 (O_944,N_24880,N_24838);
nor UO_945 (O_945,N_24944,N_24808);
nand UO_946 (O_946,N_24788,N_24970);
and UO_947 (O_947,N_24859,N_24943);
or UO_948 (O_948,N_24921,N_24760);
and UO_949 (O_949,N_24930,N_24901);
xnor UO_950 (O_950,N_24832,N_24845);
nand UO_951 (O_951,N_24978,N_24755);
nor UO_952 (O_952,N_24922,N_24942);
or UO_953 (O_953,N_24753,N_24999);
nor UO_954 (O_954,N_24945,N_24859);
and UO_955 (O_955,N_24953,N_24932);
or UO_956 (O_956,N_24999,N_24844);
nand UO_957 (O_957,N_24939,N_24910);
nand UO_958 (O_958,N_24965,N_24844);
nor UO_959 (O_959,N_24933,N_24770);
nor UO_960 (O_960,N_24992,N_24799);
nand UO_961 (O_961,N_24940,N_24773);
nor UO_962 (O_962,N_24840,N_24794);
nor UO_963 (O_963,N_24998,N_24883);
nand UO_964 (O_964,N_24914,N_24787);
and UO_965 (O_965,N_24875,N_24931);
nor UO_966 (O_966,N_24990,N_24767);
xor UO_967 (O_967,N_24991,N_24823);
nand UO_968 (O_968,N_24864,N_24993);
nor UO_969 (O_969,N_24882,N_24994);
nand UO_970 (O_970,N_24769,N_24761);
and UO_971 (O_971,N_24933,N_24911);
or UO_972 (O_972,N_24787,N_24850);
nand UO_973 (O_973,N_24825,N_24842);
or UO_974 (O_974,N_24837,N_24814);
and UO_975 (O_975,N_24792,N_24901);
nor UO_976 (O_976,N_24769,N_24884);
nand UO_977 (O_977,N_24994,N_24890);
nand UO_978 (O_978,N_24951,N_24968);
nand UO_979 (O_979,N_24827,N_24869);
nand UO_980 (O_980,N_24887,N_24963);
or UO_981 (O_981,N_24899,N_24847);
nand UO_982 (O_982,N_24822,N_24883);
nor UO_983 (O_983,N_24962,N_24805);
nand UO_984 (O_984,N_24854,N_24855);
or UO_985 (O_985,N_24967,N_24821);
nor UO_986 (O_986,N_24987,N_24839);
or UO_987 (O_987,N_24835,N_24913);
nand UO_988 (O_988,N_24947,N_24834);
nor UO_989 (O_989,N_24869,N_24757);
nand UO_990 (O_990,N_24944,N_24917);
nor UO_991 (O_991,N_24878,N_24900);
or UO_992 (O_992,N_24864,N_24869);
and UO_993 (O_993,N_24800,N_24775);
or UO_994 (O_994,N_24956,N_24849);
or UO_995 (O_995,N_24831,N_24960);
nand UO_996 (O_996,N_24960,N_24801);
nand UO_997 (O_997,N_24913,N_24806);
or UO_998 (O_998,N_24973,N_24998);
or UO_999 (O_999,N_24877,N_24762);
nor UO_1000 (O_1000,N_24949,N_24909);
or UO_1001 (O_1001,N_24821,N_24858);
and UO_1002 (O_1002,N_24884,N_24976);
nor UO_1003 (O_1003,N_24939,N_24769);
or UO_1004 (O_1004,N_24794,N_24912);
nor UO_1005 (O_1005,N_24819,N_24767);
or UO_1006 (O_1006,N_24840,N_24800);
and UO_1007 (O_1007,N_24816,N_24836);
nand UO_1008 (O_1008,N_24850,N_24905);
or UO_1009 (O_1009,N_24926,N_24931);
or UO_1010 (O_1010,N_24876,N_24776);
or UO_1011 (O_1011,N_24936,N_24976);
nand UO_1012 (O_1012,N_24751,N_24814);
nor UO_1013 (O_1013,N_24832,N_24978);
and UO_1014 (O_1014,N_24987,N_24759);
or UO_1015 (O_1015,N_24991,N_24796);
nor UO_1016 (O_1016,N_24983,N_24799);
or UO_1017 (O_1017,N_24948,N_24956);
nor UO_1018 (O_1018,N_24866,N_24767);
xnor UO_1019 (O_1019,N_24767,N_24768);
or UO_1020 (O_1020,N_24941,N_24938);
or UO_1021 (O_1021,N_24857,N_24825);
and UO_1022 (O_1022,N_24892,N_24806);
or UO_1023 (O_1023,N_24955,N_24949);
and UO_1024 (O_1024,N_24789,N_24766);
or UO_1025 (O_1025,N_24874,N_24897);
and UO_1026 (O_1026,N_24940,N_24897);
nand UO_1027 (O_1027,N_24930,N_24823);
nor UO_1028 (O_1028,N_24915,N_24880);
and UO_1029 (O_1029,N_24775,N_24893);
or UO_1030 (O_1030,N_24847,N_24805);
nand UO_1031 (O_1031,N_24779,N_24959);
nor UO_1032 (O_1032,N_24963,N_24863);
xor UO_1033 (O_1033,N_24955,N_24887);
nand UO_1034 (O_1034,N_24775,N_24795);
nor UO_1035 (O_1035,N_24934,N_24804);
nor UO_1036 (O_1036,N_24967,N_24787);
or UO_1037 (O_1037,N_24812,N_24932);
and UO_1038 (O_1038,N_24833,N_24878);
nand UO_1039 (O_1039,N_24829,N_24826);
and UO_1040 (O_1040,N_24998,N_24872);
or UO_1041 (O_1041,N_24769,N_24947);
nor UO_1042 (O_1042,N_24784,N_24951);
and UO_1043 (O_1043,N_24897,N_24821);
or UO_1044 (O_1044,N_24809,N_24843);
or UO_1045 (O_1045,N_24808,N_24934);
or UO_1046 (O_1046,N_24845,N_24967);
and UO_1047 (O_1047,N_24814,N_24831);
nand UO_1048 (O_1048,N_24803,N_24845);
and UO_1049 (O_1049,N_24861,N_24775);
nor UO_1050 (O_1050,N_24821,N_24924);
and UO_1051 (O_1051,N_24840,N_24898);
and UO_1052 (O_1052,N_24853,N_24943);
and UO_1053 (O_1053,N_24848,N_24775);
or UO_1054 (O_1054,N_24936,N_24859);
and UO_1055 (O_1055,N_24750,N_24942);
and UO_1056 (O_1056,N_24899,N_24852);
nand UO_1057 (O_1057,N_24995,N_24987);
xnor UO_1058 (O_1058,N_24860,N_24973);
or UO_1059 (O_1059,N_24894,N_24857);
nand UO_1060 (O_1060,N_24994,N_24790);
nor UO_1061 (O_1061,N_24994,N_24894);
xnor UO_1062 (O_1062,N_24899,N_24891);
and UO_1063 (O_1063,N_24832,N_24763);
or UO_1064 (O_1064,N_24792,N_24834);
nand UO_1065 (O_1065,N_24781,N_24913);
nand UO_1066 (O_1066,N_24865,N_24972);
and UO_1067 (O_1067,N_24875,N_24950);
xor UO_1068 (O_1068,N_24788,N_24985);
nor UO_1069 (O_1069,N_24959,N_24873);
and UO_1070 (O_1070,N_24873,N_24893);
nand UO_1071 (O_1071,N_24840,N_24926);
or UO_1072 (O_1072,N_24803,N_24920);
or UO_1073 (O_1073,N_24764,N_24938);
or UO_1074 (O_1074,N_24901,N_24957);
and UO_1075 (O_1075,N_24827,N_24834);
and UO_1076 (O_1076,N_24835,N_24804);
and UO_1077 (O_1077,N_24965,N_24925);
nor UO_1078 (O_1078,N_24869,N_24811);
or UO_1079 (O_1079,N_24931,N_24975);
nor UO_1080 (O_1080,N_24929,N_24816);
or UO_1081 (O_1081,N_24782,N_24816);
and UO_1082 (O_1082,N_24979,N_24804);
xor UO_1083 (O_1083,N_24757,N_24762);
nor UO_1084 (O_1084,N_24825,N_24909);
nand UO_1085 (O_1085,N_24920,N_24950);
nor UO_1086 (O_1086,N_24997,N_24798);
nor UO_1087 (O_1087,N_24961,N_24933);
nand UO_1088 (O_1088,N_24838,N_24830);
and UO_1089 (O_1089,N_24790,N_24806);
or UO_1090 (O_1090,N_24811,N_24985);
nor UO_1091 (O_1091,N_24930,N_24779);
xor UO_1092 (O_1092,N_24886,N_24883);
or UO_1093 (O_1093,N_24767,N_24912);
nand UO_1094 (O_1094,N_24890,N_24973);
xor UO_1095 (O_1095,N_24861,N_24872);
and UO_1096 (O_1096,N_24820,N_24893);
nand UO_1097 (O_1097,N_24937,N_24831);
or UO_1098 (O_1098,N_24774,N_24825);
and UO_1099 (O_1099,N_24949,N_24882);
nand UO_1100 (O_1100,N_24805,N_24966);
and UO_1101 (O_1101,N_24786,N_24967);
nor UO_1102 (O_1102,N_24771,N_24783);
nor UO_1103 (O_1103,N_24988,N_24757);
nor UO_1104 (O_1104,N_24808,N_24790);
nor UO_1105 (O_1105,N_24783,N_24990);
or UO_1106 (O_1106,N_24900,N_24811);
nand UO_1107 (O_1107,N_24981,N_24994);
or UO_1108 (O_1108,N_24873,N_24994);
nand UO_1109 (O_1109,N_24969,N_24868);
or UO_1110 (O_1110,N_24950,N_24760);
nor UO_1111 (O_1111,N_24881,N_24836);
and UO_1112 (O_1112,N_24825,N_24785);
xor UO_1113 (O_1113,N_24900,N_24838);
nor UO_1114 (O_1114,N_24875,N_24961);
or UO_1115 (O_1115,N_24992,N_24858);
and UO_1116 (O_1116,N_24963,N_24753);
or UO_1117 (O_1117,N_24804,N_24844);
and UO_1118 (O_1118,N_24864,N_24751);
nand UO_1119 (O_1119,N_24936,N_24993);
or UO_1120 (O_1120,N_24811,N_24987);
and UO_1121 (O_1121,N_24761,N_24798);
xnor UO_1122 (O_1122,N_24772,N_24792);
and UO_1123 (O_1123,N_24807,N_24810);
nor UO_1124 (O_1124,N_24971,N_24854);
nor UO_1125 (O_1125,N_24976,N_24944);
nand UO_1126 (O_1126,N_24973,N_24757);
and UO_1127 (O_1127,N_24990,N_24754);
nand UO_1128 (O_1128,N_24837,N_24806);
nor UO_1129 (O_1129,N_24953,N_24836);
or UO_1130 (O_1130,N_24814,N_24879);
nand UO_1131 (O_1131,N_24768,N_24847);
nor UO_1132 (O_1132,N_24895,N_24781);
nor UO_1133 (O_1133,N_24892,N_24820);
nor UO_1134 (O_1134,N_24940,N_24919);
nand UO_1135 (O_1135,N_24790,N_24911);
nor UO_1136 (O_1136,N_24964,N_24975);
nor UO_1137 (O_1137,N_24864,N_24970);
and UO_1138 (O_1138,N_24922,N_24871);
nor UO_1139 (O_1139,N_24829,N_24887);
and UO_1140 (O_1140,N_24958,N_24830);
or UO_1141 (O_1141,N_24986,N_24899);
nand UO_1142 (O_1142,N_24836,N_24833);
and UO_1143 (O_1143,N_24959,N_24803);
xnor UO_1144 (O_1144,N_24755,N_24759);
or UO_1145 (O_1145,N_24904,N_24758);
nor UO_1146 (O_1146,N_24787,N_24821);
nand UO_1147 (O_1147,N_24795,N_24989);
xor UO_1148 (O_1148,N_24884,N_24900);
nand UO_1149 (O_1149,N_24998,N_24977);
and UO_1150 (O_1150,N_24786,N_24931);
or UO_1151 (O_1151,N_24823,N_24920);
xnor UO_1152 (O_1152,N_24860,N_24938);
nand UO_1153 (O_1153,N_24766,N_24840);
or UO_1154 (O_1154,N_24770,N_24990);
or UO_1155 (O_1155,N_24965,N_24756);
or UO_1156 (O_1156,N_24975,N_24781);
xor UO_1157 (O_1157,N_24792,N_24850);
xnor UO_1158 (O_1158,N_24830,N_24935);
or UO_1159 (O_1159,N_24998,N_24806);
nand UO_1160 (O_1160,N_24995,N_24787);
xor UO_1161 (O_1161,N_24803,N_24978);
or UO_1162 (O_1162,N_24956,N_24843);
xor UO_1163 (O_1163,N_24890,N_24912);
nand UO_1164 (O_1164,N_24850,N_24942);
nand UO_1165 (O_1165,N_24977,N_24805);
nand UO_1166 (O_1166,N_24783,N_24937);
nand UO_1167 (O_1167,N_24991,N_24782);
nor UO_1168 (O_1168,N_24965,N_24977);
nand UO_1169 (O_1169,N_24877,N_24995);
and UO_1170 (O_1170,N_24799,N_24820);
and UO_1171 (O_1171,N_24867,N_24974);
or UO_1172 (O_1172,N_24991,N_24768);
and UO_1173 (O_1173,N_24759,N_24927);
nor UO_1174 (O_1174,N_24924,N_24881);
or UO_1175 (O_1175,N_24756,N_24761);
nand UO_1176 (O_1176,N_24851,N_24898);
or UO_1177 (O_1177,N_24755,N_24770);
xnor UO_1178 (O_1178,N_24775,N_24770);
nand UO_1179 (O_1179,N_24766,N_24911);
nand UO_1180 (O_1180,N_24836,N_24752);
or UO_1181 (O_1181,N_24853,N_24845);
and UO_1182 (O_1182,N_24981,N_24912);
nand UO_1183 (O_1183,N_24758,N_24942);
and UO_1184 (O_1184,N_24912,N_24783);
or UO_1185 (O_1185,N_24996,N_24843);
or UO_1186 (O_1186,N_24853,N_24931);
nand UO_1187 (O_1187,N_24877,N_24794);
nor UO_1188 (O_1188,N_24801,N_24996);
nor UO_1189 (O_1189,N_24834,N_24962);
nor UO_1190 (O_1190,N_24869,N_24861);
or UO_1191 (O_1191,N_24851,N_24857);
nand UO_1192 (O_1192,N_24845,N_24940);
and UO_1193 (O_1193,N_24914,N_24964);
and UO_1194 (O_1194,N_24957,N_24753);
or UO_1195 (O_1195,N_24837,N_24951);
xnor UO_1196 (O_1196,N_24921,N_24799);
xnor UO_1197 (O_1197,N_24879,N_24991);
xnor UO_1198 (O_1198,N_24943,N_24836);
and UO_1199 (O_1199,N_24903,N_24760);
or UO_1200 (O_1200,N_24882,N_24902);
nor UO_1201 (O_1201,N_24823,N_24992);
or UO_1202 (O_1202,N_24960,N_24778);
nand UO_1203 (O_1203,N_24789,N_24861);
and UO_1204 (O_1204,N_24948,N_24918);
and UO_1205 (O_1205,N_24990,N_24982);
and UO_1206 (O_1206,N_24871,N_24903);
nor UO_1207 (O_1207,N_24889,N_24854);
nor UO_1208 (O_1208,N_24934,N_24891);
or UO_1209 (O_1209,N_24911,N_24956);
nand UO_1210 (O_1210,N_24913,N_24944);
and UO_1211 (O_1211,N_24874,N_24972);
nand UO_1212 (O_1212,N_24982,N_24877);
nand UO_1213 (O_1213,N_24812,N_24922);
or UO_1214 (O_1214,N_24901,N_24898);
nor UO_1215 (O_1215,N_24896,N_24999);
and UO_1216 (O_1216,N_24977,N_24842);
nor UO_1217 (O_1217,N_24881,N_24997);
or UO_1218 (O_1218,N_24842,N_24750);
nor UO_1219 (O_1219,N_24780,N_24811);
nor UO_1220 (O_1220,N_24945,N_24979);
and UO_1221 (O_1221,N_24792,N_24979);
and UO_1222 (O_1222,N_24848,N_24791);
nand UO_1223 (O_1223,N_24901,N_24794);
nand UO_1224 (O_1224,N_24891,N_24844);
xor UO_1225 (O_1225,N_24941,N_24758);
xnor UO_1226 (O_1226,N_24952,N_24904);
nand UO_1227 (O_1227,N_24810,N_24999);
nand UO_1228 (O_1228,N_24821,N_24795);
nand UO_1229 (O_1229,N_24879,N_24926);
and UO_1230 (O_1230,N_24969,N_24764);
nand UO_1231 (O_1231,N_24781,N_24784);
or UO_1232 (O_1232,N_24976,N_24776);
nor UO_1233 (O_1233,N_24758,N_24966);
nor UO_1234 (O_1234,N_24758,N_24794);
nand UO_1235 (O_1235,N_24937,N_24848);
and UO_1236 (O_1236,N_24803,N_24864);
and UO_1237 (O_1237,N_24939,N_24889);
xor UO_1238 (O_1238,N_24993,N_24923);
nor UO_1239 (O_1239,N_24913,N_24892);
and UO_1240 (O_1240,N_24908,N_24906);
xnor UO_1241 (O_1241,N_24793,N_24984);
and UO_1242 (O_1242,N_24895,N_24827);
and UO_1243 (O_1243,N_24881,N_24831);
nor UO_1244 (O_1244,N_24930,N_24876);
or UO_1245 (O_1245,N_24962,N_24912);
xor UO_1246 (O_1246,N_24988,N_24872);
or UO_1247 (O_1247,N_24848,N_24985);
or UO_1248 (O_1248,N_24918,N_24892);
or UO_1249 (O_1249,N_24809,N_24949);
nand UO_1250 (O_1250,N_24766,N_24945);
and UO_1251 (O_1251,N_24925,N_24920);
or UO_1252 (O_1252,N_24988,N_24960);
nand UO_1253 (O_1253,N_24993,N_24817);
xor UO_1254 (O_1254,N_24893,N_24902);
or UO_1255 (O_1255,N_24899,N_24977);
and UO_1256 (O_1256,N_24795,N_24784);
and UO_1257 (O_1257,N_24934,N_24865);
and UO_1258 (O_1258,N_24777,N_24836);
or UO_1259 (O_1259,N_24943,N_24900);
or UO_1260 (O_1260,N_24821,N_24794);
and UO_1261 (O_1261,N_24976,N_24841);
or UO_1262 (O_1262,N_24985,N_24791);
nor UO_1263 (O_1263,N_24802,N_24988);
nor UO_1264 (O_1264,N_24958,N_24842);
or UO_1265 (O_1265,N_24852,N_24813);
nand UO_1266 (O_1266,N_24828,N_24857);
nor UO_1267 (O_1267,N_24986,N_24767);
nand UO_1268 (O_1268,N_24832,N_24782);
nand UO_1269 (O_1269,N_24898,N_24960);
nor UO_1270 (O_1270,N_24890,N_24851);
xnor UO_1271 (O_1271,N_24816,N_24873);
xnor UO_1272 (O_1272,N_24971,N_24948);
nand UO_1273 (O_1273,N_24898,N_24909);
or UO_1274 (O_1274,N_24949,N_24958);
nor UO_1275 (O_1275,N_24887,N_24989);
nor UO_1276 (O_1276,N_24990,N_24932);
or UO_1277 (O_1277,N_24885,N_24752);
or UO_1278 (O_1278,N_24770,N_24829);
nor UO_1279 (O_1279,N_24812,N_24987);
nand UO_1280 (O_1280,N_24994,N_24977);
nor UO_1281 (O_1281,N_24758,N_24902);
nor UO_1282 (O_1282,N_24908,N_24848);
nand UO_1283 (O_1283,N_24809,N_24856);
or UO_1284 (O_1284,N_24966,N_24889);
or UO_1285 (O_1285,N_24863,N_24754);
or UO_1286 (O_1286,N_24887,N_24811);
nor UO_1287 (O_1287,N_24943,N_24822);
nand UO_1288 (O_1288,N_24878,N_24797);
xnor UO_1289 (O_1289,N_24860,N_24971);
or UO_1290 (O_1290,N_24993,N_24998);
nor UO_1291 (O_1291,N_24765,N_24926);
nor UO_1292 (O_1292,N_24971,N_24846);
nor UO_1293 (O_1293,N_24860,N_24801);
nor UO_1294 (O_1294,N_24909,N_24877);
nand UO_1295 (O_1295,N_24829,N_24907);
or UO_1296 (O_1296,N_24884,N_24889);
nand UO_1297 (O_1297,N_24889,N_24976);
and UO_1298 (O_1298,N_24827,N_24781);
and UO_1299 (O_1299,N_24781,N_24946);
nand UO_1300 (O_1300,N_24815,N_24933);
or UO_1301 (O_1301,N_24942,N_24755);
nand UO_1302 (O_1302,N_24796,N_24889);
or UO_1303 (O_1303,N_24873,N_24837);
nand UO_1304 (O_1304,N_24813,N_24873);
or UO_1305 (O_1305,N_24986,N_24919);
nor UO_1306 (O_1306,N_24786,N_24837);
or UO_1307 (O_1307,N_24791,N_24944);
nor UO_1308 (O_1308,N_24975,N_24791);
xnor UO_1309 (O_1309,N_24887,N_24781);
xnor UO_1310 (O_1310,N_24970,N_24819);
and UO_1311 (O_1311,N_24766,N_24943);
nor UO_1312 (O_1312,N_24857,N_24844);
nand UO_1313 (O_1313,N_24974,N_24775);
nand UO_1314 (O_1314,N_24959,N_24948);
xnor UO_1315 (O_1315,N_24849,N_24915);
and UO_1316 (O_1316,N_24835,N_24916);
xor UO_1317 (O_1317,N_24981,N_24884);
and UO_1318 (O_1318,N_24859,N_24852);
nor UO_1319 (O_1319,N_24971,N_24968);
or UO_1320 (O_1320,N_24919,N_24764);
and UO_1321 (O_1321,N_24956,N_24984);
and UO_1322 (O_1322,N_24920,N_24976);
or UO_1323 (O_1323,N_24770,N_24994);
nor UO_1324 (O_1324,N_24868,N_24953);
xor UO_1325 (O_1325,N_24860,N_24820);
and UO_1326 (O_1326,N_24779,N_24890);
or UO_1327 (O_1327,N_24853,N_24933);
and UO_1328 (O_1328,N_24802,N_24986);
nor UO_1329 (O_1329,N_24824,N_24764);
or UO_1330 (O_1330,N_24936,N_24760);
xnor UO_1331 (O_1331,N_24924,N_24919);
nor UO_1332 (O_1332,N_24959,N_24816);
nor UO_1333 (O_1333,N_24791,N_24864);
and UO_1334 (O_1334,N_24831,N_24891);
and UO_1335 (O_1335,N_24846,N_24892);
xnor UO_1336 (O_1336,N_24836,N_24813);
and UO_1337 (O_1337,N_24936,N_24888);
nand UO_1338 (O_1338,N_24992,N_24985);
nor UO_1339 (O_1339,N_24932,N_24922);
nor UO_1340 (O_1340,N_24824,N_24977);
or UO_1341 (O_1341,N_24997,N_24778);
nand UO_1342 (O_1342,N_24783,N_24882);
nand UO_1343 (O_1343,N_24987,N_24956);
and UO_1344 (O_1344,N_24762,N_24879);
and UO_1345 (O_1345,N_24868,N_24848);
nor UO_1346 (O_1346,N_24933,N_24956);
xnor UO_1347 (O_1347,N_24797,N_24868);
nand UO_1348 (O_1348,N_24865,N_24853);
and UO_1349 (O_1349,N_24974,N_24925);
nand UO_1350 (O_1350,N_24892,N_24855);
xnor UO_1351 (O_1351,N_24893,N_24777);
xnor UO_1352 (O_1352,N_24900,N_24899);
or UO_1353 (O_1353,N_24807,N_24806);
nor UO_1354 (O_1354,N_24765,N_24992);
and UO_1355 (O_1355,N_24896,N_24881);
nand UO_1356 (O_1356,N_24914,N_24755);
or UO_1357 (O_1357,N_24795,N_24793);
nor UO_1358 (O_1358,N_24761,N_24966);
or UO_1359 (O_1359,N_24773,N_24966);
or UO_1360 (O_1360,N_24933,N_24955);
nand UO_1361 (O_1361,N_24838,N_24960);
nor UO_1362 (O_1362,N_24860,N_24825);
nand UO_1363 (O_1363,N_24759,N_24812);
and UO_1364 (O_1364,N_24855,N_24781);
nand UO_1365 (O_1365,N_24912,N_24886);
or UO_1366 (O_1366,N_24993,N_24806);
nor UO_1367 (O_1367,N_24783,N_24999);
nand UO_1368 (O_1368,N_24914,N_24798);
and UO_1369 (O_1369,N_24905,N_24892);
nand UO_1370 (O_1370,N_24991,N_24861);
nand UO_1371 (O_1371,N_24756,N_24998);
or UO_1372 (O_1372,N_24912,N_24776);
nor UO_1373 (O_1373,N_24948,N_24821);
and UO_1374 (O_1374,N_24787,N_24901);
and UO_1375 (O_1375,N_24850,N_24967);
or UO_1376 (O_1376,N_24753,N_24902);
and UO_1377 (O_1377,N_24799,N_24760);
nor UO_1378 (O_1378,N_24985,N_24801);
or UO_1379 (O_1379,N_24818,N_24821);
xnor UO_1380 (O_1380,N_24803,N_24790);
nand UO_1381 (O_1381,N_24991,N_24908);
and UO_1382 (O_1382,N_24869,N_24910);
nor UO_1383 (O_1383,N_24857,N_24973);
nor UO_1384 (O_1384,N_24863,N_24760);
nand UO_1385 (O_1385,N_24835,N_24918);
or UO_1386 (O_1386,N_24924,N_24991);
nand UO_1387 (O_1387,N_24761,N_24998);
nand UO_1388 (O_1388,N_24865,N_24842);
nand UO_1389 (O_1389,N_24965,N_24888);
nand UO_1390 (O_1390,N_24830,N_24976);
and UO_1391 (O_1391,N_24811,N_24939);
xor UO_1392 (O_1392,N_24774,N_24966);
or UO_1393 (O_1393,N_24853,N_24906);
or UO_1394 (O_1394,N_24888,N_24791);
or UO_1395 (O_1395,N_24864,N_24764);
nand UO_1396 (O_1396,N_24903,N_24763);
nand UO_1397 (O_1397,N_24996,N_24974);
xor UO_1398 (O_1398,N_24759,N_24901);
nor UO_1399 (O_1399,N_24840,N_24854);
or UO_1400 (O_1400,N_24750,N_24858);
nand UO_1401 (O_1401,N_24758,N_24924);
nor UO_1402 (O_1402,N_24882,N_24897);
and UO_1403 (O_1403,N_24909,N_24968);
and UO_1404 (O_1404,N_24897,N_24825);
or UO_1405 (O_1405,N_24766,N_24859);
or UO_1406 (O_1406,N_24755,N_24905);
and UO_1407 (O_1407,N_24894,N_24947);
and UO_1408 (O_1408,N_24965,N_24981);
or UO_1409 (O_1409,N_24792,N_24929);
xor UO_1410 (O_1410,N_24866,N_24907);
and UO_1411 (O_1411,N_24896,N_24930);
xor UO_1412 (O_1412,N_24777,N_24796);
and UO_1413 (O_1413,N_24851,N_24913);
or UO_1414 (O_1414,N_24875,N_24847);
or UO_1415 (O_1415,N_24899,N_24964);
or UO_1416 (O_1416,N_24963,N_24896);
or UO_1417 (O_1417,N_24815,N_24847);
nor UO_1418 (O_1418,N_24995,N_24775);
nand UO_1419 (O_1419,N_24834,N_24984);
nand UO_1420 (O_1420,N_24880,N_24843);
and UO_1421 (O_1421,N_24945,N_24970);
nand UO_1422 (O_1422,N_24941,N_24995);
nor UO_1423 (O_1423,N_24848,N_24951);
nor UO_1424 (O_1424,N_24871,N_24991);
nand UO_1425 (O_1425,N_24801,N_24950);
or UO_1426 (O_1426,N_24957,N_24936);
xor UO_1427 (O_1427,N_24795,N_24885);
and UO_1428 (O_1428,N_24803,N_24885);
and UO_1429 (O_1429,N_24819,N_24873);
nor UO_1430 (O_1430,N_24921,N_24903);
and UO_1431 (O_1431,N_24983,N_24915);
nand UO_1432 (O_1432,N_24952,N_24799);
or UO_1433 (O_1433,N_24761,N_24843);
nor UO_1434 (O_1434,N_24788,N_24968);
or UO_1435 (O_1435,N_24908,N_24989);
nor UO_1436 (O_1436,N_24787,N_24871);
nor UO_1437 (O_1437,N_24797,N_24768);
nor UO_1438 (O_1438,N_24820,N_24968);
or UO_1439 (O_1439,N_24905,N_24751);
nand UO_1440 (O_1440,N_24819,N_24760);
and UO_1441 (O_1441,N_24893,N_24770);
or UO_1442 (O_1442,N_24933,N_24816);
nor UO_1443 (O_1443,N_24951,N_24952);
or UO_1444 (O_1444,N_24816,N_24934);
nand UO_1445 (O_1445,N_24750,N_24952);
and UO_1446 (O_1446,N_24777,N_24845);
xor UO_1447 (O_1447,N_24936,N_24929);
or UO_1448 (O_1448,N_24764,N_24757);
xnor UO_1449 (O_1449,N_24951,N_24764);
and UO_1450 (O_1450,N_24956,N_24989);
nor UO_1451 (O_1451,N_24900,N_24861);
xnor UO_1452 (O_1452,N_24871,N_24786);
and UO_1453 (O_1453,N_24789,N_24776);
nand UO_1454 (O_1454,N_24908,N_24860);
nand UO_1455 (O_1455,N_24857,N_24911);
nand UO_1456 (O_1456,N_24783,N_24804);
and UO_1457 (O_1457,N_24991,N_24960);
or UO_1458 (O_1458,N_24805,N_24918);
nor UO_1459 (O_1459,N_24859,N_24791);
xnor UO_1460 (O_1460,N_24909,N_24792);
xnor UO_1461 (O_1461,N_24834,N_24932);
and UO_1462 (O_1462,N_24872,N_24932);
or UO_1463 (O_1463,N_24825,N_24977);
nand UO_1464 (O_1464,N_24761,N_24750);
nor UO_1465 (O_1465,N_24894,N_24791);
or UO_1466 (O_1466,N_24885,N_24996);
or UO_1467 (O_1467,N_24792,N_24804);
nand UO_1468 (O_1468,N_24766,N_24947);
nor UO_1469 (O_1469,N_24999,N_24828);
and UO_1470 (O_1470,N_24992,N_24754);
or UO_1471 (O_1471,N_24858,N_24846);
xnor UO_1472 (O_1472,N_24774,N_24887);
and UO_1473 (O_1473,N_24809,N_24826);
or UO_1474 (O_1474,N_24998,N_24776);
nor UO_1475 (O_1475,N_24905,N_24820);
or UO_1476 (O_1476,N_24939,N_24755);
and UO_1477 (O_1477,N_24860,N_24928);
and UO_1478 (O_1478,N_24786,N_24826);
or UO_1479 (O_1479,N_24913,N_24867);
or UO_1480 (O_1480,N_24944,N_24837);
and UO_1481 (O_1481,N_24965,N_24809);
or UO_1482 (O_1482,N_24908,N_24973);
or UO_1483 (O_1483,N_24937,N_24862);
nand UO_1484 (O_1484,N_24896,N_24970);
nor UO_1485 (O_1485,N_24996,N_24774);
nand UO_1486 (O_1486,N_24830,N_24971);
or UO_1487 (O_1487,N_24945,N_24775);
or UO_1488 (O_1488,N_24789,N_24937);
or UO_1489 (O_1489,N_24932,N_24881);
or UO_1490 (O_1490,N_24952,N_24851);
or UO_1491 (O_1491,N_24958,N_24814);
or UO_1492 (O_1492,N_24827,N_24998);
nor UO_1493 (O_1493,N_24813,N_24951);
xnor UO_1494 (O_1494,N_24770,N_24991);
and UO_1495 (O_1495,N_24975,N_24983);
nor UO_1496 (O_1496,N_24836,N_24916);
and UO_1497 (O_1497,N_24919,N_24949);
and UO_1498 (O_1498,N_24751,N_24874);
nand UO_1499 (O_1499,N_24787,N_24909);
xnor UO_1500 (O_1500,N_24895,N_24866);
nand UO_1501 (O_1501,N_24785,N_24794);
or UO_1502 (O_1502,N_24929,N_24769);
or UO_1503 (O_1503,N_24937,N_24762);
and UO_1504 (O_1504,N_24775,N_24984);
nand UO_1505 (O_1505,N_24970,N_24823);
or UO_1506 (O_1506,N_24964,N_24870);
xor UO_1507 (O_1507,N_24948,N_24875);
or UO_1508 (O_1508,N_24974,N_24936);
or UO_1509 (O_1509,N_24944,N_24750);
nor UO_1510 (O_1510,N_24818,N_24756);
nor UO_1511 (O_1511,N_24976,N_24818);
nor UO_1512 (O_1512,N_24826,N_24920);
nor UO_1513 (O_1513,N_24907,N_24832);
xnor UO_1514 (O_1514,N_24850,N_24789);
xor UO_1515 (O_1515,N_24954,N_24789);
or UO_1516 (O_1516,N_24803,N_24777);
nand UO_1517 (O_1517,N_24934,N_24871);
nor UO_1518 (O_1518,N_24907,N_24968);
nor UO_1519 (O_1519,N_24764,N_24917);
or UO_1520 (O_1520,N_24842,N_24879);
or UO_1521 (O_1521,N_24792,N_24982);
or UO_1522 (O_1522,N_24988,N_24952);
nand UO_1523 (O_1523,N_24979,N_24922);
nand UO_1524 (O_1524,N_24794,N_24886);
or UO_1525 (O_1525,N_24825,N_24846);
or UO_1526 (O_1526,N_24767,N_24774);
xnor UO_1527 (O_1527,N_24921,N_24809);
nand UO_1528 (O_1528,N_24978,N_24787);
xnor UO_1529 (O_1529,N_24987,N_24835);
nor UO_1530 (O_1530,N_24812,N_24803);
nor UO_1531 (O_1531,N_24758,N_24879);
nand UO_1532 (O_1532,N_24813,N_24890);
or UO_1533 (O_1533,N_24937,N_24791);
or UO_1534 (O_1534,N_24876,N_24806);
nor UO_1535 (O_1535,N_24930,N_24804);
nand UO_1536 (O_1536,N_24956,N_24837);
or UO_1537 (O_1537,N_24760,N_24870);
nor UO_1538 (O_1538,N_24828,N_24889);
nor UO_1539 (O_1539,N_24866,N_24987);
and UO_1540 (O_1540,N_24815,N_24890);
or UO_1541 (O_1541,N_24894,N_24902);
xor UO_1542 (O_1542,N_24909,N_24888);
nor UO_1543 (O_1543,N_24865,N_24950);
xor UO_1544 (O_1544,N_24785,N_24924);
nand UO_1545 (O_1545,N_24979,N_24995);
nand UO_1546 (O_1546,N_24894,N_24827);
or UO_1547 (O_1547,N_24943,N_24919);
or UO_1548 (O_1548,N_24806,N_24818);
and UO_1549 (O_1549,N_24774,N_24952);
nor UO_1550 (O_1550,N_24977,N_24932);
nor UO_1551 (O_1551,N_24955,N_24835);
nor UO_1552 (O_1552,N_24969,N_24936);
and UO_1553 (O_1553,N_24913,N_24899);
and UO_1554 (O_1554,N_24792,N_24752);
and UO_1555 (O_1555,N_24817,N_24933);
xnor UO_1556 (O_1556,N_24990,N_24836);
or UO_1557 (O_1557,N_24873,N_24971);
nand UO_1558 (O_1558,N_24892,N_24950);
nor UO_1559 (O_1559,N_24951,N_24828);
nor UO_1560 (O_1560,N_24842,N_24863);
nand UO_1561 (O_1561,N_24788,N_24853);
and UO_1562 (O_1562,N_24787,N_24815);
and UO_1563 (O_1563,N_24842,N_24928);
or UO_1564 (O_1564,N_24831,N_24967);
or UO_1565 (O_1565,N_24819,N_24952);
nand UO_1566 (O_1566,N_24900,N_24795);
nand UO_1567 (O_1567,N_24755,N_24777);
nand UO_1568 (O_1568,N_24826,N_24838);
or UO_1569 (O_1569,N_24971,N_24782);
nor UO_1570 (O_1570,N_24797,N_24781);
or UO_1571 (O_1571,N_24953,N_24885);
nand UO_1572 (O_1572,N_24786,N_24881);
and UO_1573 (O_1573,N_24904,N_24920);
nor UO_1574 (O_1574,N_24835,N_24975);
nand UO_1575 (O_1575,N_24909,N_24959);
and UO_1576 (O_1576,N_24985,N_24853);
nand UO_1577 (O_1577,N_24951,N_24760);
nor UO_1578 (O_1578,N_24977,N_24946);
nor UO_1579 (O_1579,N_24807,N_24966);
nand UO_1580 (O_1580,N_24770,N_24985);
xnor UO_1581 (O_1581,N_24881,N_24987);
and UO_1582 (O_1582,N_24866,N_24860);
and UO_1583 (O_1583,N_24761,N_24934);
nor UO_1584 (O_1584,N_24788,N_24796);
nand UO_1585 (O_1585,N_24790,N_24842);
xnor UO_1586 (O_1586,N_24862,N_24871);
xor UO_1587 (O_1587,N_24886,N_24878);
or UO_1588 (O_1588,N_24894,N_24760);
and UO_1589 (O_1589,N_24773,N_24783);
xnor UO_1590 (O_1590,N_24860,N_24852);
or UO_1591 (O_1591,N_24818,N_24913);
and UO_1592 (O_1592,N_24847,N_24897);
and UO_1593 (O_1593,N_24838,N_24833);
nand UO_1594 (O_1594,N_24989,N_24936);
xnor UO_1595 (O_1595,N_24803,N_24842);
nor UO_1596 (O_1596,N_24939,N_24942);
nor UO_1597 (O_1597,N_24772,N_24887);
nor UO_1598 (O_1598,N_24813,N_24952);
nor UO_1599 (O_1599,N_24768,N_24834);
nor UO_1600 (O_1600,N_24944,N_24777);
xor UO_1601 (O_1601,N_24940,N_24879);
and UO_1602 (O_1602,N_24779,N_24980);
nor UO_1603 (O_1603,N_24917,N_24856);
nand UO_1604 (O_1604,N_24990,N_24815);
and UO_1605 (O_1605,N_24874,N_24777);
nor UO_1606 (O_1606,N_24811,N_24772);
nand UO_1607 (O_1607,N_24882,N_24916);
nand UO_1608 (O_1608,N_24910,N_24883);
or UO_1609 (O_1609,N_24858,N_24872);
xnor UO_1610 (O_1610,N_24762,N_24890);
and UO_1611 (O_1611,N_24833,N_24852);
or UO_1612 (O_1612,N_24933,N_24846);
or UO_1613 (O_1613,N_24903,N_24770);
nand UO_1614 (O_1614,N_24860,N_24859);
xor UO_1615 (O_1615,N_24990,N_24881);
nand UO_1616 (O_1616,N_24789,N_24935);
nor UO_1617 (O_1617,N_24952,N_24980);
or UO_1618 (O_1618,N_24781,N_24896);
nand UO_1619 (O_1619,N_24813,N_24906);
nand UO_1620 (O_1620,N_24800,N_24868);
or UO_1621 (O_1621,N_24793,N_24812);
nand UO_1622 (O_1622,N_24986,N_24844);
and UO_1623 (O_1623,N_24875,N_24993);
and UO_1624 (O_1624,N_24789,N_24792);
nand UO_1625 (O_1625,N_24895,N_24798);
or UO_1626 (O_1626,N_24994,N_24918);
or UO_1627 (O_1627,N_24817,N_24984);
nand UO_1628 (O_1628,N_24964,N_24970);
and UO_1629 (O_1629,N_24806,N_24770);
nand UO_1630 (O_1630,N_24876,N_24914);
nand UO_1631 (O_1631,N_24782,N_24863);
nand UO_1632 (O_1632,N_24855,N_24932);
nor UO_1633 (O_1633,N_24919,N_24968);
or UO_1634 (O_1634,N_24923,N_24949);
nand UO_1635 (O_1635,N_24944,N_24977);
xnor UO_1636 (O_1636,N_24936,N_24956);
and UO_1637 (O_1637,N_24790,N_24932);
nand UO_1638 (O_1638,N_24958,N_24845);
and UO_1639 (O_1639,N_24980,N_24816);
nor UO_1640 (O_1640,N_24817,N_24877);
nand UO_1641 (O_1641,N_24907,N_24900);
and UO_1642 (O_1642,N_24759,N_24970);
or UO_1643 (O_1643,N_24871,N_24847);
nor UO_1644 (O_1644,N_24937,N_24958);
and UO_1645 (O_1645,N_24950,N_24889);
nand UO_1646 (O_1646,N_24961,N_24764);
nor UO_1647 (O_1647,N_24808,N_24932);
xor UO_1648 (O_1648,N_24968,N_24764);
nor UO_1649 (O_1649,N_24772,N_24955);
or UO_1650 (O_1650,N_24881,N_24899);
and UO_1651 (O_1651,N_24790,N_24834);
xnor UO_1652 (O_1652,N_24960,N_24819);
or UO_1653 (O_1653,N_24751,N_24953);
or UO_1654 (O_1654,N_24960,N_24825);
or UO_1655 (O_1655,N_24974,N_24999);
or UO_1656 (O_1656,N_24891,N_24861);
and UO_1657 (O_1657,N_24964,N_24778);
xnor UO_1658 (O_1658,N_24778,N_24827);
xor UO_1659 (O_1659,N_24874,N_24788);
nand UO_1660 (O_1660,N_24798,N_24816);
nand UO_1661 (O_1661,N_24858,N_24782);
or UO_1662 (O_1662,N_24971,N_24987);
and UO_1663 (O_1663,N_24976,N_24910);
and UO_1664 (O_1664,N_24996,N_24787);
and UO_1665 (O_1665,N_24760,N_24751);
and UO_1666 (O_1666,N_24887,N_24795);
or UO_1667 (O_1667,N_24887,N_24790);
or UO_1668 (O_1668,N_24787,N_24801);
nand UO_1669 (O_1669,N_24770,N_24917);
or UO_1670 (O_1670,N_24916,N_24791);
and UO_1671 (O_1671,N_24781,N_24908);
and UO_1672 (O_1672,N_24870,N_24965);
nand UO_1673 (O_1673,N_24841,N_24892);
xnor UO_1674 (O_1674,N_24833,N_24985);
nand UO_1675 (O_1675,N_24751,N_24922);
xnor UO_1676 (O_1676,N_24783,N_24920);
or UO_1677 (O_1677,N_24944,N_24841);
nor UO_1678 (O_1678,N_24960,N_24947);
xnor UO_1679 (O_1679,N_24814,N_24904);
nor UO_1680 (O_1680,N_24773,N_24995);
or UO_1681 (O_1681,N_24757,N_24826);
and UO_1682 (O_1682,N_24786,N_24849);
or UO_1683 (O_1683,N_24890,N_24764);
and UO_1684 (O_1684,N_24915,N_24863);
nor UO_1685 (O_1685,N_24762,N_24826);
nor UO_1686 (O_1686,N_24998,N_24980);
nand UO_1687 (O_1687,N_24784,N_24928);
xor UO_1688 (O_1688,N_24789,N_24756);
and UO_1689 (O_1689,N_24945,N_24908);
nor UO_1690 (O_1690,N_24953,N_24802);
nand UO_1691 (O_1691,N_24913,N_24755);
nor UO_1692 (O_1692,N_24892,N_24898);
nor UO_1693 (O_1693,N_24761,N_24850);
and UO_1694 (O_1694,N_24998,N_24838);
nand UO_1695 (O_1695,N_24782,N_24852);
nand UO_1696 (O_1696,N_24753,N_24941);
or UO_1697 (O_1697,N_24843,N_24949);
nand UO_1698 (O_1698,N_24807,N_24790);
nand UO_1699 (O_1699,N_24982,N_24762);
nand UO_1700 (O_1700,N_24961,N_24828);
and UO_1701 (O_1701,N_24766,N_24858);
nand UO_1702 (O_1702,N_24871,N_24964);
or UO_1703 (O_1703,N_24899,N_24839);
nand UO_1704 (O_1704,N_24810,N_24920);
and UO_1705 (O_1705,N_24967,N_24863);
nand UO_1706 (O_1706,N_24756,N_24767);
or UO_1707 (O_1707,N_24993,N_24947);
and UO_1708 (O_1708,N_24834,N_24884);
nor UO_1709 (O_1709,N_24925,N_24763);
xor UO_1710 (O_1710,N_24975,N_24822);
and UO_1711 (O_1711,N_24781,N_24948);
nor UO_1712 (O_1712,N_24987,N_24867);
nor UO_1713 (O_1713,N_24891,N_24920);
nor UO_1714 (O_1714,N_24976,N_24764);
nand UO_1715 (O_1715,N_24759,N_24922);
or UO_1716 (O_1716,N_24781,N_24952);
nand UO_1717 (O_1717,N_24783,N_24916);
nor UO_1718 (O_1718,N_24906,N_24936);
xor UO_1719 (O_1719,N_24793,N_24898);
nand UO_1720 (O_1720,N_24798,N_24789);
nand UO_1721 (O_1721,N_24903,N_24889);
nand UO_1722 (O_1722,N_24814,N_24921);
nor UO_1723 (O_1723,N_24762,N_24946);
or UO_1724 (O_1724,N_24831,N_24793);
nor UO_1725 (O_1725,N_24936,N_24897);
nand UO_1726 (O_1726,N_24925,N_24881);
and UO_1727 (O_1727,N_24823,N_24906);
or UO_1728 (O_1728,N_24810,N_24784);
or UO_1729 (O_1729,N_24801,N_24828);
nor UO_1730 (O_1730,N_24752,N_24777);
nand UO_1731 (O_1731,N_24882,N_24957);
xnor UO_1732 (O_1732,N_24885,N_24844);
xor UO_1733 (O_1733,N_24969,N_24858);
and UO_1734 (O_1734,N_24858,N_24773);
and UO_1735 (O_1735,N_24762,N_24923);
nand UO_1736 (O_1736,N_24923,N_24931);
nand UO_1737 (O_1737,N_24908,N_24892);
and UO_1738 (O_1738,N_24924,N_24911);
or UO_1739 (O_1739,N_24950,N_24874);
nand UO_1740 (O_1740,N_24920,N_24800);
nor UO_1741 (O_1741,N_24821,N_24878);
nand UO_1742 (O_1742,N_24826,N_24843);
nand UO_1743 (O_1743,N_24938,N_24988);
nand UO_1744 (O_1744,N_24869,N_24773);
nor UO_1745 (O_1745,N_24753,N_24839);
nor UO_1746 (O_1746,N_24846,N_24807);
xor UO_1747 (O_1747,N_24896,N_24816);
nor UO_1748 (O_1748,N_24822,N_24985);
xnor UO_1749 (O_1749,N_24976,N_24955);
xnor UO_1750 (O_1750,N_24943,N_24868);
and UO_1751 (O_1751,N_24830,N_24900);
xnor UO_1752 (O_1752,N_24947,N_24785);
or UO_1753 (O_1753,N_24812,N_24881);
nand UO_1754 (O_1754,N_24768,N_24779);
and UO_1755 (O_1755,N_24985,N_24916);
xor UO_1756 (O_1756,N_24898,N_24750);
nand UO_1757 (O_1757,N_24896,N_24947);
nand UO_1758 (O_1758,N_24883,N_24935);
and UO_1759 (O_1759,N_24800,N_24906);
and UO_1760 (O_1760,N_24820,N_24999);
xor UO_1761 (O_1761,N_24907,N_24833);
nand UO_1762 (O_1762,N_24867,N_24767);
or UO_1763 (O_1763,N_24970,N_24865);
or UO_1764 (O_1764,N_24885,N_24845);
xor UO_1765 (O_1765,N_24828,N_24781);
xnor UO_1766 (O_1766,N_24772,N_24786);
or UO_1767 (O_1767,N_24762,N_24847);
nand UO_1768 (O_1768,N_24796,N_24772);
nand UO_1769 (O_1769,N_24892,N_24929);
nor UO_1770 (O_1770,N_24906,N_24804);
nor UO_1771 (O_1771,N_24775,N_24954);
xor UO_1772 (O_1772,N_24861,N_24807);
and UO_1773 (O_1773,N_24944,N_24921);
or UO_1774 (O_1774,N_24781,N_24788);
nand UO_1775 (O_1775,N_24814,N_24888);
or UO_1776 (O_1776,N_24970,N_24977);
nand UO_1777 (O_1777,N_24878,N_24793);
and UO_1778 (O_1778,N_24835,N_24836);
nor UO_1779 (O_1779,N_24903,N_24750);
or UO_1780 (O_1780,N_24830,N_24874);
and UO_1781 (O_1781,N_24875,N_24830);
or UO_1782 (O_1782,N_24935,N_24766);
nand UO_1783 (O_1783,N_24928,N_24921);
nand UO_1784 (O_1784,N_24830,N_24939);
nand UO_1785 (O_1785,N_24822,N_24802);
nand UO_1786 (O_1786,N_24917,N_24824);
or UO_1787 (O_1787,N_24779,N_24858);
xor UO_1788 (O_1788,N_24764,N_24811);
nand UO_1789 (O_1789,N_24811,N_24922);
or UO_1790 (O_1790,N_24945,N_24975);
and UO_1791 (O_1791,N_24803,N_24901);
and UO_1792 (O_1792,N_24902,N_24870);
and UO_1793 (O_1793,N_24913,N_24896);
nor UO_1794 (O_1794,N_24806,N_24952);
xor UO_1795 (O_1795,N_24853,N_24891);
nor UO_1796 (O_1796,N_24904,N_24865);
or UO_1797 (O_1797,N_24977,N_24785);
nor UO_1798 (O_1798,N_24854,N_24861);
nand UO_1799 (O_1799,N_24789,N_24796);
nand UO_1800 (O_1800,N_24945,N_24842);
or UO_1801 (O_1801,N_24803,N_24928);
and UO_1802 (O_1802,N_24972,N_24824);
nand UO_1803 (O_1803,N_24928,N_24844);
and UO_1804 (O_1804,N_24798,N_24848);
nor UO_1805 (O_1805,N_24989,N_24948);
nand UO_1806 (O_1806,N_24945,N_24893);
and UO_1807 (O_1807,N_24755,N_24926);
xnor UO_1808 (O_1808,N_24849,N_24853);
nor UO_1809 (O_1809,N_24971,N_24767);
nand UO_1810 (O_1810,N_24845,N_24796);
or UO_1811 (O_1811,N_24935,N_24767);
xnor UO_1812 (O_1812,N_24885,N_24960);
and UO_1813 (O_1813,N_24956,N_24852);
and UO_1814 (O_1814,N_24973,N_24902);
nand UO_1815 (O_1815,N_24771,N_24970);
or UO_1816 (O_1816,N_24925,N_24941);
or UO_1817 (O_1817,N_24940,N_24926);
or UO_1818 (O_1818,N_24802,N_24990);
xnor UO_1819 (O_1819,N_24975,N_24973);
or UO_1820 (O_1820,N_24765,N_24921);
xnor UO_1821 (O_1821,N_24996,N_24871);
nand UO_1822 (O_1822,N_24895,N_24754);
and UO_1823 (O_1823,N_24846,N_24936);
and UO_1824 (O_1824,N_24953,N_24765);
nor UO_1825 (O_1825,N_24852,N_24934);
or UO_1826 (O_1826,N_24925,N_24883);
and UO_1827 (O_1827,N_24802,N_24867);
nor UO_1828 (O_1828,N_24963,N_24842);
or UO_1829 (O_1829,N_24791,N_24890);
and UO_1830 (O_1830,N_24831,N_24849);
nand UO_1831 (O_1831,N_24977,N_24911);
xnor UO_1832 (O_1832,N_24979,N_24838);
or UO_1833 (O_1833,N_24841,N_24765);
and UO_1834 (O_1834,N_24807,N_24921);
xor UO_1835 (O_1835,N_24873,N_24918);
and UO_1836 (O_1836,N_24847,N_24825);
nor UO_1837 (O_1837,N_24899,N_24866);
and UO_1838 (O_1838,N_24772,N_24998);
nor UO_1839 (O_1839,N_24843,N_24868);
nor UO_1840 (O_1840,N_24767,N_24944);
nand UO_1841 (O_1841,N_24781,N_24983);
nand UO_1842 (O_1842,N_24947,N_24956);
nor UO_1843 (O_1843,N_24757,N_24933);
and UO_1844 (O_1844,N_24769,N_24877);
nand UO_1845 (O_1845,N_24895,N_24912);
and UO_1846 (O_1846,N_24851,N_24908);
or UO_1847 (O_1847,N_24893,N_24762);
and UO_1848 (O_1848,N_24918,N_24849);
or UO_1849 (O_1849,N_24886,N_24973);
nor UO_1850 (O_1850,N_24957,N_24997);
and UO_1851 (O_1851,N_24759,N_24802);
nor UO_1852 (O_1852,N_24945,N_24854);
nor UO_1853 (O_1853,N_24777,N_24758);
and UO_1854 (O_1854,N_24799,N_24856);
xor UO_1855 (O_1855,N_24801,N_24958);
xnor UO_1856 (O_1856,N_24967,N_24816);
nand UO_1857 (O_1857,N_24828,N_24873);
and UO_1858 (O_1858,N_24794,N_24995);
nand UO_1859 (O_1859,N_24771,N_24870);
nor UO_1860 (O_1860,N_24888,N_24874);
or UO_1861 (O_1861,N_24772,N_24891);
nor UO_1862 (O_1862,N_24915,N_24781);
nand UO_1863 (O_1863,N_24987,N_24861);
nor UO_1864 (O_1864,N_24994,N_24957);
and UO_1865 (O_1865,N_24850,N_24983);
and UO_1866 (O_1866,N_24978,N_24825);
or UO_1867 (O_1867,N_24968,N_24992);
and UO_1868 (O_1868,N_24888,N_24948);
nand UO_1869 (O_1869,N_24850,N_24962);
and UO_1870 (O_1870,N_24831,N_24903);
or UO_1871 (O_1871,N_24811,N_24841);
nor UO_1872 (O_1872,N_24811,N_24783);
or UO_1873 (O_1873,N_24998,N_24825);
nor UO_1874 (O_1874,N_24818,N_24808);
nor UO_1875 (O_1875,N_24864,N_24991);
or UO_1876 (O_1876,N_24869,N_24909);
nand UO_1877 (O_1877,N_24881,N_24959);
nor UO_1878 (O_1878,N_24824,N_24929);
and UO_1879 (O_1879,N_24801,N_24756);
and UO_1880 (O_1880,N_24792,N_24920);
or UO_1881 (O_1881,N_24791,N_24935);
nor UO_1882 (O_1882,N_24873,N_24863);
xor UO_1883 (O_1883,N_24816,N_24890);
xor UO_1884 (O_1884,N_24954,N_24815);
nor UO_1885 (O_1885,N_24750,N_24930);
and UO_1886 (O_1886,N_24948,N_24932);
nor UO_1887 (O_1887,N_24950,N_24982);
or UO_1888 (O_1888,N_24802,N_24973);
and UO_1889 (O_1889,N_24803,N_24820);
nor UO_1890 (O_1890,N_24846,N_24795);
nor UO_1891 (O_1891,N_24781,N_24837);
or UO_1892 (O_1892,N_24923,N_24786);
or UO_1893 (O_1893,N_24948,N_24928);
nor UO_1894 (O_1894,N_24987,N_24933);
or UO_1895 (O_1895,N_24811,N_24840);
nand UO_1896 (O_1896,N_24765,N_24891);
and UO_1897 (O_1897,N_24892,N_24891);
and UO_1898 (O_1898,N_24939,N_24948);
nor UO_1899 (O_1899,N_24865,N_24963);
or UO_1900 (O_1900,N_24846,N_24918);
or UO_1901 (O_1901,N_24878,N_24776);
nand UO_1902 (O_1902,N_24954,N_24816);
and UO_1903 (O_1903,N_24988,N_24763);
nand UO_1904 (O_1904,N_24971,N_24900);
and UO_1905 (O_1905,N_24778,N_24808);
nand UO_1906 (O_1906,N_24813,N_24855);
and UO_1907 (O_1907,N_24910,N_24950);
nand UO_1908 (O_1908,N_24907,N_24827);
nor UO_1909 (O_1909,N_24987,N_24909);
nor UO_1910 (O_1910,N_24832,N_24842);
nand UO_1911 (O_1911,N_24812,N_24944);
xnor UO_1912 (O_1912,N_24786,N_24998);
or UO_1913 (O_1913,N_24979,N_24953);
nor UO_1914 (O_1914,N_24950,N_24790);
or UO_1915 (O_1915,N_24935,N_24777);
nand UO_1916 (O_1916,N_24984,N_24918);
and UO_1917 (O_1917,N_24801,N_24935);
nor UO_1918 (O_1918,N_24784,N_24970);
or UO_1919 (O_1919,N_24932,N_24981);
nand UO_1920 (O_1920,N_24838,N_24964);
nand UO_1921 (O_1921,N_24800,N_24778);
or UO_1922 (O_1922,N_24998,N_24854);
and UO_1923 (O_1923,N_24894,N_24763);
or UO_1924 (O_1924,N_24923,N_24799);
nand UO_1925 (O_1925,N_24889,N_24958);
and UO_1926 (O_1926,N_24832,N_24795);
and UO_1927 (O_1927,N_24950,N_24948);
nor UO_1928 (O_1928,N_24951,N_24876);
or UO_1929 (O_1929,N_24782,N_24990);
nand UO_1930 (O_1930,N_24863,N_24948);
nand UO_1931 (O_1931,N_24781,N_24809);
nand UO_1932 (O_1932,N_24879,N_24787);
and UO_1933 (O_1933,N_24925,N_24798);
and UO_1934 (O_1934,N_24995,N_24918);
nor UO_1935 (O_1935,N_24996,N_24863);
nor UO_1936 (O_1936,N_24940,N_24776);
and UO_1937 (O_1937,N_24872,N_24916);
nand UO_1938 (O_1938,N_24891,N_24982);
and UO_1939 (O_1939,N_24753,N_24953);
or UO_1940 (O_1940,N_24796,N_24867);
nor UO_1941 (O_1941,N_24867,N_24907);
or UO_1942 (O_1942,N_24777,N_24926);
nand UO_1943 (O_1943,N_24774,N_24795);
nor UO_1944 (O_1944,N_24830,N_24928);
and UO_1945 (O_1945,N_24945,N_24982);
xnor UO_1946 (O_1946,N_24755,N_24983);
nand UO_1947 (O_1947,N_24855,N_24848);
and UO_1948 (O_1948,N_24944,N_24968);
or UO_1949 (O_1949,N_24969,N_24775);
or UO_1950 (O_1950,N_24853,N_24794);
or UO_1951 (O_1951,N_24920,N_24815);
and UO_1952 (O_1952,N_24949,N_24902);
nor UO_1953 (O_1953,N_24822,N_24855);
nor UO_1954 (O_1954,N_24912,N_24905);
nor UO_1955 (O_1955,N_24802,N_24936);
nor UO_1956 (O_1956,N_24893,N_24892);
nand UO_1957 (O_1957,N_24756,N_24784);
nor UO_1958 (O_1958,N_24769,N_24752);
nand UO_1959 (O_1959,N_24844,N_24852);
or UO_1960 (O_1960,N_24897,N_24956);
and UO_1961 (O_1961,N_24843,N_24812);
nor UO_1962 (O_1962,N_24916,N_24823);
or UO_1963 (O_1963,N_24870,N_24757);
xor UO_1964 (O_1964,N_24953,N_24750);
and UO_1965 (O_1965,N_24987,N_24826);
or UO_1966 (O_1966,N_24969,N_24932);
and UO_1967 (O_1967,N_24756,N_24936);
and UO_1968 (O_1968,N_24826,N_24847);
and UO_1969 (O_1969,N_24959,N_24927);
nand UO_1970 (O_1970,N_24870,N_24907);
or UO_1971 (O_1971,N_24788,N_24956);
nand UO_1972 (O_1972,N_24820,N_24856);
or UO_1973 (O_1973,N_24956,N_24866);
nand UO_1974 (O_1974,N_24943,N_24764);
nor UO_1975 (O_1975,N_24873,N_24975);
nor UO_1976 (O_1976,N_24961,N_24770);
nand UO_1977 (O_1977,N_24776,N_24985);
nand UO_1978 (O_1978,N_24783,N_24816);
and UO_1979 (O_1979,N_24901,N_24844);
nor UO_1980 (O_1980,N_24883,N_24895);
nand UO_1981 (O_1981,N_24895,N_24862);
or UO_1982 (O_1982,N_24955,N_24944);
nand UO_1983 (O_1983,N_24909,N_24757);
nor UO_1984 (O_1984,N_24920,N_24897);
nand UO_1985 (O_1985,N_24779,N_24841);
nand UO_1986 (O_1986,N_24908,N_24817);
and UO_1987 (O_1987,N_24926,N_24860);
nand UO_1988 (O_1988,N_24821,N_24949);
nand UO_1989 (O_1989,N_24801,N_24981);
and UO_1990 (O_1990,N_24896,N_24888);
and UO_1991 (O_1991,N_24916,N_24895);
or UO_1992 (O_1992,N_24822,N_24968);
or UO_1993 (O_1993,N_24855,N_24981);
nand UO_1994 (O_1994,N_24951,N_24750);
and UO_1995 (O_1995,N_24817,N_24923);
or UO_1996 (O_1996,N_24851,N_24883);
nor UO_1997 (O_1997,N_24979,N_24764);
or UO_1998 (O_1998,N_24853,N_24862);
nand UO_1999 (O_1999,N_24901,N_24761);
nand UO_2000 (O_2000,N_24919,N_24873);
and UO_2001 (O_2001,N_24818,N_24993);
and UO_2002 (O_2002,N_24840,N_24830);
and UO_2003 (O_2003,N_24917,N_24869);
nand UO_2004 (O_2004,N_24973,N_24834);
nand UO_2005 (O_2005,N_24887,N_24946);
and UO_2006 (O_2006,N_24958,N_24826);
nor UO_2007 (O_2007,N_24758,N_24907);
nor UO_2008 (O_2008,N_24798,N_24931);
and UO_2009 (O_2009,N_24953,N_24769);
nor UO_2010 (O_2010,N_24809,N_24895);
or UO_2011 (O_2011,N_24952,N_24933);
or UO_2012 (O_2012,N_24910,N_24909);
xnor UO_2013 (O_2013,N_24940,N_24810);
nor UO_2014 (O_2014,N_24960,N_24927);
nand UO_2015 (O_2015,N_24855,N_24902);
nand UO_2016 (O_2016,N_24948,N_24750);
nand UO_2017 (O_2017,N_24881,N_24784);
or UO_2018 (O_2018,N_24877,N_24756);
or UO_2019 (O_2019,N_24997,N_24861);
nor UO_2020 (O_2020,N_24860,N_24958);
nand UO_2021 (O_2021,N_24999,N_24831);
and UO_2022 (O_2022,N_24871,N_24895);
nor UO_2023 (O_2023,N_24772,N_24927);
and UO_2024 (O_2024,N_24950,N_24813);
and UO_2025 (O_2025,N_24832,N_24895);
or UO_2026 (O_2026,N_24904,N_24934);
nand UO_2027 (O_2027,N_24931,N_24889);
nand UO_2028 (O_2028,N_24805,N_24790);
or UO_2029 (O_2029,N_24958,N_24923);
or UO_2030 (O_2030,N_24962,N_24794);
xnor UO_2031 (O_2031,N_24801,N_24945);
and UO_2032 (O_2032,N_24789,N_24907);
or UO_2033 (O_2033,N_24896,N_24886);
nor UO_2034 (O_2034,N_24862,N_24865);
or UO_2035 (O_2035,N_24983,N_24818);
or UO_2036 (O_2036,N_24812,N_24989);
and UO_2037 (O_2037,N_24955,N_24799);
or UO_2038 (O_2038,N_24838,N_24914);
and UO_2039 (O_2039,N_24961,N_24995);
or UO_2040 (O_2040,N_24942,N_24770);
nor UO_2041 (O_2041,N_24939,N_24752);
nand UO_2042 (O_2042,N_24810,N_24856);
nor UO_2043 (O_2043,N_24925,N_24773);
nor UO_2044 (O_2044,N_24782,N_24968);
nand UO_2045 (O_2045,N_24931,N_24978);
nor UO_2046 (O_2046,N_24903,N_24807);
or UO_2047 (O_2047,N_24827,N_24886);
or UO_2048 (O_2048,N_24923,N_24753);
nand UO_2049 (O_2049,N_24978,N_24782);
or UO_2050 (O_2050,N_24786,N_24854);
xor UO_2051 (O_2051,N_24971,N_24962);
xor UO_2052 (O_2052,N_24824,N_24906);
xnor UO_2053 (O_2053,N_24927,N_24914);
nor UO_2054 (O_2054,N_24929,N_24863);
or UO_2055 (O_2055,N_24942,N_24828);
and UO_2056 (O_2056,N_24874,N_24864);
or UO_2057 (O_2057,N_24956,N_24785);
nand UO_2058 (O_2058,N_24822,N_24926);
nand UO_2059 (O_2059,N_24953,N_24840);
or UO_2060 (O_2060,N_24908,N_24846);
and UO_2061 (O_2061,N_24968,N_24814);
nor UO_2062 (O_2062,N_24755,N_24774);
nor UO_2063 (O_2063,N_24869,N_24987);
nor UO_2064 (O_2064,N_24753,N_24976);
and UO_2065 (O_2065,N_24982,N_24767);
nor UO_2066 (O_2066,N_24773,N_24968);
or UO_2067 (O_2067,N_24779,N_24871);
xnor UO_2068 (O_2068,N_24779,N_24909);
and UO_2069 (O_2069,N_24855,N_24880);
and UO_2070 (O_2070,N_24835,N_24756);
or UO_2071 (O_2071,N_24840,N_24858);
xor UO_2072 (O_2072,N_24854,N_24769);
nor UO_2073 (O_2073,N_24863,N_24940);
or UO_2074 (O_2074,N_24910,N_24885);
nand UO_2075 (O_2075,N_24910,N_24892);
or UO_2076 (O_2076,N_24938,N_24985);
nor UO_2077 (O_2077,N_24794,N_24930);
nor UO_2078 (O_2078,N_24764,N_24992);
or UO_2079 (O_2079,N_24786,N_24991);
xnor UO_2080 (O_2080,N_24753,N_24879);
nand UO_2081 (O_2081,N_24763,N_24985);
or UO_2082 (O_2082,N_24927,N_24843);
nand UO_2083 (O_2083,N_24852,N_24773);
nor UO_2084 (O_2084,N_24926,N_24964);
nand UO_2085 (O_2085,N_24866,N_24819);
or UO_2086 (O_2086,N_24751,N_24758);
xor UO_2087 (O_2087,N_24790,N_24787);
nand UO_2088 (O_2088,N_24936,N_24866);
nor UO_2089 (O_2089,N_24777,N_24909);
or UO_2090 (O_2090,N_24819,N_24761);
nor UO_2091 (O_2091,N_24868,N_24834);
nand UO_2092 (O_2092,N_24764,N_24983);
nand UO_2093 (O_2093,N_24751,N_24802);
and UO_2094 (O_2094,N_24788,N_24945);
nand UO_2095 (O_2095,N_24923,N_24889);
or UO_2096 (O_2096,N_24991,N_24865);
nor UO_2097 (O_2097,N_24917,N_24899);
nand UO_2098 (O_2098,N_24919,N_24952);
nor UO_2099 (O_2099,N_24836,N_24788);
nor UO_2100 (O_2100,N_24822,N_24974);
and UO_2101 (O_2101,N_24869,N_24879);
nand UO_2102 (O_2102,N_24943,N_24974);
and UO_2103 (O_2103,N_24865,N_24974);
or UO_2104 (O_2104,N_24787,N_24753);
nand UO_2105 (O_2105,N_24781,N_24899);
or UO_2106 (O_2106,N_24832,N_24912);
nand UO_2107 (O_2107,N_24752,N_24881);
nor UO_2108 (O_2108,N_24817,N_24784);
and UO_2109 (O_2109,N_24921,N_24974);
and UO_2110 (O_2110,N_24815,N_24828);
nand UO_2111 (O_2111,N_24868,N_24817);
and UO_2112 (O_2112,N_24777,N_24959);
xnor UO_2113 (O_2113,N_24903,N_24872);
or UO_2114 (O_2114,N_24884,N_24839);
or UO_2115 (O_2115,N_24790,N_24942);
and UO_2116 (O_2116,N_24907,N_24853);
nand UO_2117 (O_2117,N_24962,N_24769);
and UO_2118 (O_2118,N_24993,N_24957);
or UO_2119 (O_2119,N_24867,N_24786);
xor UO_2120 (O_2120,N_24847,N_24902);
nand UO_2121 (O_2121,N_24994,N_24999);
nor UO_2122 (O_2122,N_24889,N_24870);
and UO_2123 (O_2123,N_24832,N_24905);
nor UO_2124 (O_2124,N_24818,N_24912);
or UO_2125 (O_2125,N_24869,N_24839);
nand UO_2126 (O_2126,N_24951,N_24882);
or UO_2127 (O_2127,N_24774,N_24769);
nor UO_2128 (O_2128,N_24940,N_24819);
and UO_2129 (O_2129,N_24988,N_24914);
and UO_2130 (O_2130,N_24823,N_24826);
nand UO_2131 (O_2131,N_24813,N_24980);
or UO_2132 (O_2132,N_24868,N_24865);
or UO_2133 (O_2133,N_24874,N_24976);
nand UO_2134 (O_2134,N_24869,N_24966);
nor UO_2135 (O_2135,N_24971,N_24868);
or UO_2136 (O_2136,N_24993,N_24896);
nand UO_2137 (O_2137,N_24753,N_24850);
or UO_2138 (O_2138,N_24892,N_24779);
nor UO_2139 (O_2139,N_24917,N_24795);
or UO_2140 (O_2140,N_24940,N_24878);
xor UO_2141 (O_2141,N_24965,N_24817);
or UO_2142 (O_2142,N_24896,N_24783);
nand UO_2143 (O_2143,N_24785,N_24771);
nand UO_2144 (O_2144,N_24862,N_24971);
nor UO_2145 (O_2145,N_24814,N_24840);
xnor UO_2146 (O_2146,N_24995,N_24767);
nand UO_2147 (O_2147,N_24860,N_24821);
nand UO_2148 (O_2148,N_24872,N_24928);
nor UO_2149 (O_2149,N_24939,N_24756);
nor UO_2150 (O_2150,N_24851,N_24789);
nand UO_2151 (O_2151,N_24859,N_24967);
nor UO_2152 (O_2152,N_24985,N_24829);
xnor UO_2153 (O_2153,N_24893,N_24767);
nor UO_2154 (O_2154,N_24935,N_24772);
or UO_2155 (O_2155,N_24786,N_24953);
nor UO_2156 (O_2156,N_24784,N_24802);
nor UO_2157 (O_2157,N_24910,N_24971);
xor UO_2158 (O_2158,N_24781,N_24806);
or UO_2159 (O_2159,N_24886,N_24991);
xnor UO_2160 (O_2160,N_24896,N_24795);
xnor UO_2161 (O_2161,N_24924,N_24783);
xnor UO_2162 (O_2162,N_24885,N_24807);
and UO_2163 (O_2163,N_24776,N_24972);
nand UO_2164 (O_2164,N_24826,N_24927);
or UO_2165 (O_2165,N_24995,N_24888);
or UO_2166 (O_2166,N_24850,N_24949);
nor UO_2167 (O_2167,N_24757,N_24830);
or UO_2168 (O_2168,N_24903,N_24811);
nand UO_2169 (O_2169,N_24846,N_24848);
or UO_2170 (O_2170,N_24985,N_24879);
or UO_2171 (O_2171,N_24769,N_24758);
nor UO_2172 (O_2172,N_24869,N_24784);
or UO_2173 (O_2173,N_24884,N_24799);
and UO_2174 (O_2174,N_24973,N_24893);
or UO_2175 (O_2175,N_24854,N_24784);
and UO_2176 (O_2176,N_24964,N_24980);
nand UO_2177 (O_2177,N_24930,N_24765);
and UO_2178 (O_2178,N_24761,N_24865);
nor UO_2179 (O_2179,N_24966,N_24968);
nand UO_2180 (O_2180,N_24815,N_24806);
or UO_2181 (O_2181,N_24862,N_24965);
nand UO_2182 (O_2182,N_24912,N_24889);
nor UO_2183 (O_2183,N_24920,N_24927);
nand UO_2184 (O_2184,N_24942,N_24902);
nor UO_2185 (O_2185,N_24835,N_24845);
and UO_2186 (O_2186,N_24837,N_24937);
nor UO_2187 (O_2187,N_24892,N_24911);
or UO_2188 (O_2188,N_24982,N_24943);
and UO_2189 (O_2189,N_24984,N_24922);
nand UO_2190 (O_2190,N_24848,N_24830);
nand UO_2191 (O_2191,N_24888,N_24892);
or UO_2192 (O_2192,N_24875,N_24986);
and UO_2193 (O_2193,N_24955,N_24930);
nor UO_2194 (O_2194,N_24966,N_24777);
or UO_2195 (O_2195,N_24898,N_24994);
nor UO_2196 (O_2196,N_24768,N_24926);
nand UO_2197 (O_2197,N_24965,N_24770);
nand UO_2198 (O_2198,N_24963,N_24975);
and UO_2199 (O_2199,N_24829,N_24777);
and UO_2200 (O_2200,N_24949,N_24839);
and UO_2201 (O_2201,N_24919,N_24966);
or UO_2202 (O_2202,N_24886,N_24957);
or UO_2203 (O_2203,N_24964,N_24844);
and UO_2204 (O_2204,N_24790,N_24812);
xor UO_2205 (O_2205,N_24831,N_24930);
and UO_2206 (O_2206,N_24949,N_24948);
nand UO_2207 (O_2207,N_24891,N_24994);
or UO_2208 (O_2208,N_24884,N_24793);
xnor UO_2209 (O_2209,N_24753,N_24996);
or UO_2210 (O_2210,N_24806,N_24990);
nor UO_2211 (O_2211,N_24995,N_24906);
and UO_2212 (O_2212,N_24965,N_24942);
or UO_2213 (O_2213,N_24785,N_24789);
or UO_2214 (O_2214,N_24874,N_24894);
or UO_2215 (O_2215,N_24861,N_24791);
or UO_2216 (O_2216,N_24781,N_24787);
nor UO_2217 (O_2217,N_24915,N_24876);
or UO_2218 (O_2218,N_24793,N_24895);
nor UO_2219 (O_2219,N_24936,N_24838);
or UO_2220 (O_2220,N_24962,N_24933);
nand UO_2221 (O_2221,N_24876,N_24787);
nand UO_2222 (O_2222,N_24949,N_24776);
and UO_2223 (O_2223,N_24813,N_24968);
and UO_2224 (O_2224,N_24808,N_24897);
nand UO_2225 (O_2225,N_24772,N_24988);
nor UO_2226 (O_2226,N_24925,N_24814);
nand UO_2227 (O_2227,N_24961,N_24797);
nand UO_2228 (O_2228,N_24797,N_24937);
and UO_2229 (O_2229,N_24834,N_24924);
and UO_2230 (O_2230,N_24845,N_24791);
nor UO_2231 (O_2231,N_24928,N_24942);
and UO_2232 (O_2232,N_24773,N_24767);
nand UO_2233 (O_2233,N_24811,N_24877);
and UO_2234 (O_2234,N_24877,N_24840);
and UO_2235 (O_2235,N_24761,N_24951);
or UO_2236 (O_2236,N_24858,N_24836);
xor UO_2237 (O_2237,N_24800,N_24771);
nand UO_2238 (O_2238,N_24899,N_24827);
nand UO_2239 (O_2239,N_24933,N_24812);
or UO_2240 (O_2240,N_24813,N_24776);
or UO_2241 (O_2241,N_24867,N_24801);
and UO_2242 (O_2242,N_24954,N_24988);
xor UO_2243 (O_2243,N_24824,N_24910);
or UO_2244 (O_2244,N_24936,N_24886);
xnor UO_2245 (O_2245,N_24860,N_24823);
and UO_2246 (O_2246,N_24790,N_24762);
xnor UO_2247 (O_2247,N_24761,N_24896);
xor UO_2248 (O_2248,N_24978,N_24913);
or UO_2249 (O_2249,N_24886,N_24845);
xor UO_2250 (O_2250,N_24871,N_24857);
or UO_2251 (O_2251,N_24869,N_24895);
xnor UO_2252 (O_2252,N_24991,N_24809);
nor UO_2253 (O_2253,N_24993,N_24807);
and UO_2254 (O_2254,N_24815,N_24893);
nor UO_2255 (O_2255,N_24870,N_24930);
nor UO_2256 (O_2256,N_24886,N_24844);
or UO_2257 (O_2257,N_24921,N_24851);
nand UO_2258 (O_2258,N_24755,N_24947);
nor UO_2259 (O_2259,N_24945,N_24798);
and UO_2260 (O_2260,N_24999,N_24881);
xor UO_2261 (O_2261,N_24958,N_24793);
or UO_2262 (O_2262,N_24847,N_24813);
nand UO_2263 (O_2263,N_24927,N_24771);
nand UO_2264 (O_2264,N_24760,N_24775);
nand UO_2265 (O_2265,N_24916,N_24867);
xor UO_2266 (O_2266,N_24931,N_24990);
nor UO_2267 (O_2267,N_24869,N_24945);
nand UO_2268 (O_2268,N_24825,N_24911);
nand UO_2269 (O_2269,N_24941,N_24867);
xnor UO_2270 (O_2270,N_24855,N_24910);
or UO_2271 (O_2271,N_24913,N_24986);
or UO_2272 (O_2272,N_24922,N_24854);
or UO_2273 (O_2273,N_24817,N_24890);
nand UO_2274 (O_2274,N_24972,N_24949);
and UO_2275 (O_2275,N_24854,N_24963);
and UO_2276 (O_2276,N_24810,N_24894);
nor UO_2277 (O_2277,N_24810,N_24907);
or UO_2278 (O_2278,N_24886,N_24884);
nor UO_2279 (O_2279,N_24973,N_24867);
nor UO_2280 (O_2280,N_24808,N_24850);
nand UO_2281 (O_2281,N_24881,N_24961);
and UO_2282 (O_2282,N_24900,N_24805);
or UO_2283 (O_2283,N_24860,N_24984);
and UO_2284 (O_2284,N_24914,N_24868);
xor UO_2285 (O_2285,N_24828,N_24859);
nor UO_2286 (O_2286,N_24809,N_24786);
nor UO_2287 (O_2287,N_24892,N_24752);
nor UO_2288 (O_2288,N_24877,N_24787);
nor UO_2289 (O_2289,N_24982,N_24902);
or UO_2290 (O_2290,N_24977,N_24921);
xnor UO_2291 (O_2291,N_24966,N_24784);
nand UO_2292 (O_2292,N_24916,N_24925);
or UO_2293 (O_2293,N_24983,N_24917);
or UO_2294 (O_2294,N_24903,N_24958);
nor UO_2295 (O_2295,N_24955,N_24833);
nand UO_2296 (O_2296,N_24785,N_24997);
nor UO_2297 (O_2297,N_24760,N_24907);
or UO_2298 (O_2298,N_24980,N_24889);
or UO_2299 (O_2299,N_24889,N_24816);
xnor UO_2300 (O_2300,N_24753,N_24861);
or UO_2301 (O_2301,N_24962,N_24910);
nor UO_2302 (O_2302,N_24847,N_24892);
or UO_2303 (O_2303,N_24987,N_24799);
nand UO_2304 (O_2304,N_24942,N_24769);
nor UO_2305 (O_2305,N_24800,N_24797);
nand UO_2306 (O_2306,N_24977,N_24856);
and UO_2307 (O_2307,N_24783,N_24885);
or UO_2308 (O_2308,N_24984,N_24980);
nor UO_2309 (O_2309,N_24966,N_24810);
nand UO_2310 (O_2310,N_24903,N_24843);
xnor UO_2311 (O_2311,N_24937,N_24996);
nand UO_2312 (O_2312,N_24933,N_24833);
nor UO_2313 (O_2313,N_24833,N_24899);
xnor UO_2314 (O_2314,N_24792,N_24847);
nand UO_2315 (O_2315,N_24933,N_24804);
nand UO_2316 (O_2316,N_24983,N_24957);
xor UO_2317 (O_2317,N_24812,N_24773);
nor UO_2318 (O_2318,N_24967,N_24929);
nand UO_2319 (O_2319,N_24757,N_24913);
nor UO_2320 (O_2320,N_24819,N_24954);
or UO_2321 (O_2321,N_24925,N_24823);
nor UO_2322 (O_2322,N_24785,N_24851);
nand UO_2323 (O_2323,N_24798,N_24750);
and UO_2324 (O_2324,N_24942,N_24975);
or UO_2325 (O_2325,N_24853,N_24787);
and UO_2326 (O_2326,N_24828,N_24909);
xnor UO_2327 (O_2327,N_24951,N_24985);
nor UO_2328 (O_2328,N_24953,N_24902);
xor UO_2329 (O_2329,N_24982,N_24764);
nand UO_2330 (O_2330,N_24937,N_24926);
nor UO_2331 (O_2331,N_24900,N_24992);
or UO_2332 (O_2332,N_24928,N_24988);
or UO_2333 (O_2333,N_24773,N_24808);
and UO_2334 (O_2334,N_24858,N_24767);
nand UO_2335 (O_2335,N_24994,N_24909);
or UO_2336 (O_2336,N_24826,N_24966);
or UO_2337 (O_2337,N_24910,N_24757);
and UO_2338 (O_2338,N_24911,N_24792);
nand UO_2339 (O_2339,N_24798,N_24977);
and UO_2340 (O_2340,N_24946,N_24970);
nor UO_2341 (O_2341,N_24811,N_24753);
and UO_2342 (O_2342,N_24955,N_24889);
xor UO_2343 (O_2343,N_24831,N_24866);
nor UO_2344 (O_2344,N_24902,N_24991);
or UO_2345 (O_2345,N_24810,N_24778);
or UO_2346 (O_2346,N_24869,N_24968);
nor UO_2347 (O_2347,N_24907,N_24998);
nor UO_2348 (O_2348,N_24772,N_24899);
nor UO_2349 (O_2349,N_24753,N_24759);
and UO_2350 (O_2350,N_24896,N_24838);
and UO_2351 (O_2351,N_24752,N_24869);
and UO_2352 (O_2352,N_24950,N_24757);
nand UO_2353 (O_2353,N_24905,N_24891);
nor UO_2354 (O_2354,N_24765,N_24882);
or UO_2355 (O_2355,N_24770,N_24993);
and UO_2356 (O_2356,N_24991,N_24868);
or UO_2357 (O_2357,N_24900,N_24818);
nor UO_2358 (O_2358,N_24952,N_24917);
nor UO_2359 (O_2359,N_24961,N_24906);
nor UO_2360 (O_2360,N_24818,N_24958);
nand UO_2361 (O_2361,N_24892,N_24941);
and UO_2362 (O_2362,N_24919,N_24954);
nor UO_2363 (O_2363,N_24876,N_24796);
nand UO_2364 (O_2364,N_24878,N_24992);
or UO_2365 (O_2365,N_24860,N_24855);
nand UO_2366 (O_2366,N_24906,N_24895);
or UO_2367 (O_2367,N_24819,N_24906);
nor UO_2368 (O_2368,N_24829,N_24868);
and UO_2369 (O_2369,N_24936,N_24927);
and UO_2370 (O_2370,N_24796,N_24806);
nand UO_2371 (O_2371,N_24990,N_24863);
and UO_2372 (O_2372,N_24890,N_24863);
or UO_2373 (O_2373,N_24910,N_24754);
or UO_2374 (O_2374,N_24806,N_24870);
nor UO_2375 (O_2375,N_24825,N_24942);
xnor UO_2376 (O_2376,N_24855,N_24946);
xor UO_2377 (O_2377,N_24973,N_24859);
nor UO_2378 (O_2378,N_24916,N_24812);
nand UO_2379 (O_2379,N_24788,N_24997);
nor UO_2380 (O_2380,N_24862,N_24951);
and UO_2381 (O_2381,N_24789,N_24942);
and UO_2382 (O_2382,N_24985,N_24980);
nor UO_2383 (O_2383,N_24885,N_24846);
xnor UO_2384 (O_2384,N_24804,N_24909);
nand UO_2385 (O_2385,N_24762,N_24850);
or UO_2386 (O_2386,N_24753,N_24956);
nor UO_2387 (O_2387,N_24938,N_24793);
nor UO_2388 (O_2388,N_24971,N_24946);
and UO_2389 (O_2389,N_24884,N_24802);
and UO_2390 (O_2390,N_24968,N_24889);
and UO_2391 (O_2391,N_24759,N_24878);
nor UO_2392 (O_2392,N_24795,N_24806);
xnor UO_2393 (O_2393,N_24882,N_24817);
nand UO_2394 (O_2394,N_24950,N_24870);
or UO_2395 (O_2395,N_24909,N_24775);
nor UO_2396 (O_2396,N_24959,N_24759);
and UO_2397 (O_2397,N_24934,N_24988);
nand UO_2398 (O_2398,N_24814,N_24887);
nand UO_2399 (O_2399,N_24902,N_24937);
nand UO_2400 (O_2400,N_24857,N_24914);
or UO_2401 (O_2401,N_24951,N_24845);
nor UO_2402 (O_2402,N_24788,N_24873);
nor UO_2403 (O_2403,N_24783,N_24886);
xor UO_2404 (O_2404,N_24753,N_24925);
nor UO_2405 (O_2405,N_24818,N_24932);
and UO_2406 (O_2406,N_24977,N_24871);
or UO_2407 (O_2407,N_24851,N_24897);
or UO_2408 (O_2408,N_24856,N_24847);
nor UO_2409 (O_2409,N_24835,N_24888);
or UO_2410 (O_2410,N_24845,N_24837);
or UO_2411 (O_2411,N_24792,N_24985);
nand UO_2412 (O_2412,N_24920,N_24926);
nor UO_2413 (O_2413,N_24853,N_24908);
or UO_2414 (O_2414,N_24854,N_24886);
nor UO_2415 (O_2415,N_24760,N_24755);
nand UO_2416 (O_2416,N_24793,N_24765);
nor UO_2417 (O_2417,N_24908,N_24836);
and UO_2418 (O_2418,N_24754,N_24933);
and UO_2419 (O_2419,N_24891,N_24966);
or UO_2420 (O_2420,N_24903,N_24926);
nand UO_2421 (O_2421,N_24814,N_24907);
and UO_2422 (O_2422,N_24873,N_24848);
nor UO_2423 (O_2423,N_24889,N_24959);
nor UO_2424 (O_2424,N_24782,N_24918);
nand UO_2425 (O_2425,N_24783,N_24839);
nor UO_2426 (O_2426,N_24949,N_24931);
xnor UO_2427 (O_2427,N_24951,N_24956);
or UO_2428 (O_2428,N_24832,N_24812);
nand UO_2429 (O_2429,N_24905,N_24843);
nor UO_2430 (O_2430,N_24900,N_24785);
and UO_2431 (O_2431,N_24807,N_24754);
and UO_2432 (O_2432,N_24887,N_24933);
or UO_2433 (O_2433,N_24851,N_24891);
or UO_2434 (O_2434,N_24906,N_24924);
nor UO_2435 (O_2435,N_24945,N_24796);
and UO_2436 (O_2436,N_24823,N_24814);
or UO_2437 (O_2437,N_24887,N_24775);
nor UO_2438 (O_2438,N_24920,N_24866);
and UO_2439 (O_2439,N_24878,N_24995);
and UO_2440 (O_2440,N_24927,N_24846);
xnor UO_2441 (O_2441,N_24909,N_24957);
or UO_2442 (O_2442,N_24854,N_24817);
xor UO_2443 (O_2443,N_24835,N_24934);
or UO_2444 (O_2444,N_24957,N_24945);
and UO_2445 (O_2445,N_24894,N_24965);
and UO_2446 (O_2446,N_24838,N_24937);
and UO_2447 (O_2447,N_24870,N_24885);
nand UO_2448 (O_2448,N_24912,N_24917);
and UO_2449 (O_2449,N_24821,N_24845);
nand UO_2450 (O_2450,N_24914,N_24789);
nor UO_2451 (O_2451,N_24933,N_24997);
nand UO_2452 (O_2452,N_24921,N_24961);
nand UO_2453 (O_2453,N_24813,N_24841);
and UO_2454 (O_2454,N_24926,N_24863);
nand UO_2455 (O_2455,N_24797,N_24896);
or UO_2456 (O_2456,N_24928,N_24792);
nor UO_2457 (O_2457,N_24957,N_24877);
and UO_2458 (O_2458,N_24973,N_24852);
nor UO_2459 (O_2459,N_24893,N_24930);
xor UO_2460 (O_2460,N_24787,N_24889);
and UO_2461 (O_2461,N_24883,N_24790);
or UO_2462 (O_2462,N_24859,N_24815);
or UO_2463 (O_2463,N_24781,N_24813);
nor UO_2464 (O_2464,N_24827,N_24949);
nor UO_2465 (O_2465,N_24882,N_24778);
xor UO_2466 (O_2466,N_24805,N_24833);
nand UO_2467 (O_2467,N_24863,N_24934);
nand UO_2468 (O_2468,N_24813,N_24851);
or UO_2469 (O_2469,N_24777,N_24902);
and UO_2470 (O_2470,N_24767,N_24806);
and UO_2471 (O_2471,N_24992,N_24957);
xor UO_2472 (O_2472,N_24941,N_24954);
nor UO_2473 (O_2473,N_24866,N_24908);
or UO_2474 (O_2474,N_24863,N_24808);
nand UO_2475 (O_2475,N_24887,N_24755);
and UO_2476 (O_2476,N_24873,N_24849);
or UO_2477 (O_2477,N_24918,N_24823);
nand UO_2478 (O_2478,N_24922,N_24956);
nand UO_2479 (O_2479,N_24920,N_24968);
xor UO_2480 (O_2480,N_24806,N_24788);
nor UO_2481 (O_2481,N_24912,N_24831);
xor UO_2482 (O_2482,N_24880,N_24982);
nor UO_2483 (O_2483,N_24873,N_24796);
xor UO_2484 (O_2484,N_24962,N_24789);
xnor UO_2485 (O_2485,N_24861,N_24950);
and UO_2486 (O_2486,N_24909,N_24918);
and UO_2487 (O_2487,N_24986,N_24838);
and UO_2488 (O_2488,N_24862,N_24882);
or UO_2489 (O_2489,N_24871,N_24933);
and UO_2490 (O_2490,N_24966,N_24926);
nor UO_2491 (O_2491,N_24876,N_24755);
and UO_2492 (O_2492,N_24927,N_24947);
nand UO_2493 (O_2493,N_24954,N_24905);
nand UO_2494 (O_2494,N_24808,N_24898);
and UO_2495 (O_2495,N_24874,N_24896);
and UO_2496 (O_2496,N_24860,N_24796);
and UO_2497 (O_2497,N_24893,N_24874);
nand UO_2498 (O_2498,N_24980,N_24996);
and UO_2499 (O_2499,N_24946,N_24757);
nand UO_2500 (O_2500,N_24929,N_24768);
nor UO_2501 (O_2501,N_24837,N_24867);
nand UO_2502 (O_2502,N_24864,N_24823);
and UO_2503 (O_2503,N_24937,N_24938);
and UO_2504 (O_2504,N_24781,N_24963);
nor UO_2505 (O_2505,N_24850,N_24899);
nand UO_2506 (O_2506,N_24997,N_24822);
nor UO_2507 (O_2507,N_24895,N_24750);
and UO_2508 (O_2508,N_24781,N_24869);
or UO_2509 (O_2509,N_24773,N_24909);
nor UO_2510 (O_2510,N_24754,N_24784);
and UO_2511 (O_2511,N_24846,N_24906);
or UO_2512 (O_2512,N_24932,N_24777);
nand UO_2513 (O_2513,N_24773,N_24915);
xnor UO_2514 (O_2514,N_24984,N_24822);
nand UO_2515 (O_2515,N_24936,N_24881);
nor UO_2516 (O_2516,N_24896,N_24972);
and UO_2517 (O_2517,N_24962,N_24788);
nand UO_2518 (O_2518,N_24788,N_24966);
nand UO_2519 (O_2519,N_24900,N_24824);
or UO_2520 (O_2520,N_24984,N_24878);
or UO_2521 (O_2521,N_24998,N_24762);
and UO_2522 (O_2522,N_24810,N_24899);
and UO_2523 (O_2523,N_24777,N_24917);
or UO_2524 (O_2524,N_24864,N_24946);
nor UO_2525 (O_2525,N_24900,N_24978);
and UO_2526 (O_2526,N_24896,N_24813);
and UO_2527 (O_2527,N_24931,N_24856);
and UO_2528 (O_2528,N_24910,N_24825);
and UO_2529 (O_2529,N_24889,N_24874);
or UO_2530 (O_2530,N_24990,N_24826);
nor UO_2531 (O_2531,N_24810,N_24893);
and UO_2532 (O_2532,N_24802,N_24768);
nand UO_2533 (O_2533,N_24970,N_24938);
xnor UO_2534 (O_2534,N_24751,N_24913);
and UO_2535 (O_2535,N_24887,N_24925);
or UO_2536 (O_2536,N_24837,N_24835);
and UO_2537 (O_2537,N_24827,N_24902);
or UO_2538 (O_2538,N_24789,N_24974);
nor UO_2539 (O_2539,N_24984,N_24921);
nand UO_2540 (O_2540,N_24803,N_24850);
nand UO_2541 (O_2541,N_24952,N_24804);
or UO_2542 (O_2542,N_24951,N_24980);
and UO_2543 (O_2543,N_24979,N_24833);
xnor UO_2544 (O_2544,N_24910,N_24896);
nor UO_2545 (O_2545,N_24943,N_24947);
and UO_2546 (O_2546,N_24932,N_24971);
nand UO_2547 (O_2547,N_24918,N_24988);
or UO_2548 (O_2548,N_24975,N_24961);
nor UO_2549 (O_2549,N_24875,N_24980);
and UO_2550 (O_2550,N_24830,N_24811);
nand UO_2551 (O_2551,N_24995,N_24813);
nor UO_2552 (O_2552,N_24981,N_24940);
xor UO_2553 (O_2553,N_24832,N_24835);
nor UO_2554 (O_2554,N_24964,N_24960);
xnor UO_2555 (O_2555,N_24999,N_24956);
and UO_2556 (O_2556,N_24819,N_24809);
nand UO_2557 (O_2557,N_24949,N_24795);
nand UO_2558 (O_2558,N_24990,N_24976);
nand UO_2559 (O_2559,N_24771,N_24823);
nand UO_2560 (O_2560,N_24797,N_24779);
or UO_2561 (O_2561,N_24830,N_24906);
nor UO_2562 (O_2562,N_24850,N_24764);
nor UO_2563 (O_2563,N_24848,N_24820);
or UO_2564 (O_2564,N_24770,N_24847);
nand UO_2565 (O_2565,N_24930,N_24943);
or UO_2566 (O_2566,N_24958,N_24847);
and UO_2567 (O_2567,N_24931,N_24941);
and UO_2568 (O_2568,N_24957,N_24764);
nor UO_2569 (O_2569,N_24836,N_24844);
nor UO_2570 (O_2570,N_24847,N_24965);
xor UO_2571 (O_2571,N_24761,N_24773);
nand UO_2572 (O_2572,N_24814,N_24988);
xor UO_2573 (O_2573,N_24885,N_24908);
nand UO_2574 (O_2574,N_24858,N_24861);
and UO_2575 (O_2575,N_24848,N_24774);
or UO_2576 (O_2576,N_24821,N_24983);
nand UO_2577 (O_2577,N_24839,N_24912);
nand UO_2578 (O_2578,N_24867,N_24953);
or UO_2579 (O_2579,N_24993,N_24764);
or UO_2580 (O_2580,N_24906,N_24780);
nor UO_2581 (O_2581,N_24819,N_24976);
nand UO_2582 (O_2582,N_24800,N_24980);
nor UO_2583 (O_2583,N_24888,N_24942);
nor UO_2584 (O_2584,N_24883,N_24966);
or UO_2585 (O_2585,N_24860,N_24901);
or UO_2586 (O_2586,N_24911,N_24926);
nor UO_2587 (O_2587,N_24919,N_24758);
and UO_2588 (O_2588,N_24809,N_24948);
nand UO_2589 (O_2589,N_24953,N_24804);
nand UO_2590 (O_2590,N_24880,N_24798);
nor UO_2591 (O_2591,N_24870,N_24853);
or UO_2592 (O_2592,N_24873,N_24897);
nand UO_2593 (O_2593,N_24872,N_24970);
nand UO_2594 (O_2594,N_24812,N_24789);
nand UO_2595 (O_2595,N_24777,N_24838);
nor UO_2596 (O_2596,N_24934,N_24813);
xnor UO_2597 (O_2597,N_24995,N_24947);
nand UO_2598 (O_2598,N_24898,N_24885);
nand UO_2599 (O_2599,N_24836,N_24967);
nor UO_2600 (O_2600,N_24838,N_24761);
nor UO_2601 (O_2601,N_24904,N_24863);
nor UO_2602 (O_2602,N_24829,N_24806);
nor UO_2603 (O_2603,N_24877,N_24846);
and UO_2604 (O_2604,N_24979,N_24793);
nor UO_2605 (O_2605,N_24955,N_24919);
and UO_2606 (O_2606,N_24908,N_24889);
and UO_2607 (O_2607,N_24825,N_24800);
and UO_2608 (O_2608,N_24911,N_24783);
or UO_2609 (O_2609,N_24839,N_24890);
and UO_2610 (O_2610,N_24833,N_24980);
nor UO_2611 (O_2611,N_24872,N_24804);
or UO_2612 (O_2612,N_24896,N_24833);
or UO_2613 (O_2613,N_24878,N_24987);
and UO_2614 (O_2614,N_24942,N_24786);
nor UO_2615 (O_2615,N_24889,N_24888);
xor UO_2616 (O_2616,N_24938,N_24870);
or UO_2617 (O_2617,N_24989,N_24851);
nor UO_2618 (O_2618,N_24911,N_24887);
or UO_2619 (O_2619,N_24797,N_24959);
nand UO_2620 (O_2620,N_24968,N_24842);
nor UO_2621 (O_2621,N_24821,N_24782);
or UO_2622 (O_2622,N_24947,N_24904);
and UO_2623 (O_2623,N_24853,N_24885);
and UO_2624 (O_2624,N_24822,N_24823);
or UO_2625 (O_2625,N_24984,N_24988);
xnor UO_2626 (O_2626,N_24914,N_24963);
nand UO_2627 (O_2627,N_24856,N_24784);
nand UO_2628 (O_2628,N_24942,N_24852);
nor UO_2629 (O_2629,N_24850,N_24767);
and UO_2630 (O_2630,N_24870,N_24959);
nor UO_2631 (O_2631,N_24996,N_24861);
nand UO_2632 (O_2632,N_24988,N_24821);
or UO_2633 (O_2633,N_24789,N_24836);
xnor UO_2634 (O_2634,N_24992,N_24894);
or UO_2635 (O_2635,N_24979,N_24831);
nand UO_2636 (O_2636,N_24928,N_24756);
and UO_2637 (O_2637,N_24810,N_24967);
or UO_2638 (O_2638,N_24826,N_24856);
nand UO_2639 (O_2639,N_24830,N_24765);
nor UO_2640 (O_2640,N_24837,N_24927);
or UO_2641 (O_2641,N_24971,N_24980);
xnor UO_2642 (O_2642,N_24806,N_24997);
nor UO_2643 (O_2643,N_24966,N_24892);
xnor UO_2644 (O_2644,N_24819,N_24898);
nand UO_2645 (O_2645,N_24810,N_24750);
nand UO_2646 (O_2646,N_24924,N_24792);
nand UO_2647 (O_2647,N_24780,N_24989);
nor UO_2648 (O_2648,N_24773,N_24928);
or UO_2649 (O_2649,N_24789,N_24958);
or UO_2650 (O_2650,N_24900,N_24972);
nor UO_2651 (O_2651,N_24783,N_24831);
nor UO_2652 (O_2652,N_24924,N_24993);
and UO_2653 (O_2653,N_24954,N_24785);
nor UO_2654 (O_2654,N_24961,N_24753);
and UO_2655 (O_2655,N_24896,N_24765);
and UO_2656 (O_2656,N_24844,N_24753);
nand UO_2657 (O_2657,N_24766,N_24963);
nor UO_2658 (O_2658,N_24965,N_24971);
xor UO_2659 (O_2659,N_24868,N_24767);
nor UO_2660 (O_2660,N_24958,N_24941);
nor UO_2661 (O_2661,N_24782,N_24751);
and UO_2662 (O_2662,N_24903,N_24976);
nor UO_2663 (O_2663,N_24879,N_24883);
nor UO_2664 (O_2664,N_24961,N_24842);
or UO_2665 (O_2665,N_24906,N_24794);
nor UO_2666 (O_2666,N_24975,N_24895);
nor UO_2667 (O_2667,N_24934,N_24857);
nand UO_2668 (O_2668,N_24789,N_24934);
nand UO_2669 (O_2669,N_24754,N_24759);
nor UO_2670 (O_2670,N_24899,N_24873);
nand UO_2671 (O_2671,N_24858,N_24762);
xnor UO_2672 (O_2672,N_24795,N_24974);
and UO_2673 (O_2673,N_24791,N_24852);
nand UO_2674 (O_2674,N_24929,N_24919);
nor UO_2675 (O_2675,N_24958,N_24836);
nor UO_2676 (O_2676,N_24794,N_24900);
xnor UO_2677 (O_2677,N_24783,N_24900);
and UO_2678 (O_2678,N_24873,N_24898);
and UO_2679 (O_2679,N_24966,N_24768);
xnor UO_2680 (O_2680,N_24947,N_24923);
or UO_2681 (O_2681,N_24921,N_24906);
or UO_2682 (O_2682,N_24818,N_24795);
nand UO_2683 (O_2683,N_24942,N_24839);
nor UO_2684 (O_2684,N_24944,N_24836);
nor UO_2685 (O_2685,N_24813,N_24892);
nor UO_2686 (O_2686,N_24941,N_24991);
nor UO_2687 (O_2687,N_24859,N_24816);
nand UO_2688 (O_2688,N_24953,N_24851);
xnor UO_2689 (O_2689,N_24792,N_24803);
nor UO_2690 (O_2690,N_24836,N_24889);
xor UO_2691 (O_2691,N_24839,N_24797);
and UO_2692 (O_2692,N_24958,N_24878);
or UO_2693 (O_2693,N_24815,N_24884);
xnor UO_2694 (O_2694,N_24907,N_24805);
and UO_2695 (O_2695,N_24901,N_24890);
xor UO_2696 (O_2696,N_24813,N_24911);
or UO_2697 (O_2697,N_24855,N_24915);
or UO_2698 (O_2698,N_24961,N_24991);
xnor UO_2699 (O_2699,N_24941,N_24824);
xnor UO_2700 (O_2700,N_24877,N_24805);
and UO_2701 (O_2701,N_24777,N_24931);
nor UO_2702 (O_2702,N_24983,N_24866);
and UO_2703 (O_2703,N_24803,N_24811);
nor UO_2704 (O_2704,N_24995,N_24962);
nor UO_2705 (O_2705,N_24817,N_24930);
nand UO_2706 (O_2706,N_24919,N_24973);
nor UO_2707 (O_2707,N_24839,N_24944);
nand UO_2708 (O_2708,N_24833,N_24823);
and UO_2709 (O_2709,N_24855,N_24853);
or UO_2710 (O_2710,N_24942,N_24991);
nand UO_2711 (O_2711,N_24967,N_24981);
nor UO_2712 (O_2712,N_24936,N_24990);
nand UO_2713 (O_2713,N_24863,N_24911);
or UO_2714 (O_2714,N_24917,N_24930);
nand UO_2715 (O_2715,N_24763,N_24964);
nor UO_2716 (O_2716,N_24817,N_24833);
or UO_2717 (O_2717,N_24986,N_24997);
nand UO_2718 (O_2718,N_24847,N_24961);
xor UO_2719 (O_2719,N_24867,N_24877);
and UO_2720 (O_2720,N_24919,N_24811);
and UO_2721 (O_2721,N_24993,N_24915);
or UO_2722 (O_2722,N_24916,N_24865);
nor UO_2723 (O_2723,N_24830,N_24786);
xnor UO_2724 (O_2724,N_24991,N_24802);
nor UO_2725 (O_2725,N_24890,N_24891);
and UO_2726 (O_2726,N_24967,N_24817);
or UO_2727 (O_2727,N_24799,N_24834);
nor UO_2728 (O_2728,N_24901,N_24800);
nor UO_2729 (O_2729,N_24817,N_24940);
and UO_2730 (O_2730,N_24831,N_24846);
and UO_2731 (O_2731,N_24917,N_24943);
xor UO_2732 (O_2732,N_24934,N_24902);
nand UO_2733 (O_2733,N_24948,N_24899);
nand UO_2734 (O_2734,N_24917,N_24822);
nor UO_2735 (O_2735,N_24984,N_24925);
nor UO_2736 (O_2736,N_24979,N_24789);
nor UO_2737 (O_2737,N_24980,N_24937);
or UO_2738 (O_2738,N_24773,N_24959);
or UO_2739 (O_2739,N_24794,N_24767);
nand UO_2740 (O_2740,N_24888,N_24967);
nand UO_2741 (O_2741,N_24920,N_24837);
nor UO_2742 (O_2742,N_24819,N_24843);
and UO_2743 (O_2743,N_24969,N_24832);
or UO_2744 (O_2744,N_24885,N_24957);
nor UO_2745 (O_2745,N_24835,N_24854);
nor UO_2746 (O_2746,N_24994,N_24809);
or UO_2747 (O_2747,N_24998,N_24771);
or UO_2748 (O_2748,N_24795,N_24812);
or UO_2749 (O_2749,N_24948,N_24895);
or UO_2750 (O_2750,N_24825,N_24890);
nor UO_2751 (O_2751,N_24931,N_24857);
or UO_2752 (O_2752,N_24903,N_24943);
nand UO_2753 (O_2753,N_24769,N_24798);
nor UO_2754 (O_2754,N_24899,N_24862);
nor UO_2755 (O_2755,N_24869,N_24800);
xor UO_2756 (O_2756,N_24819,N_24875);
and UO_2757 (O_2757,N_24933,N_24836);
nand UO_2758 (O_2758,N_24809,N_24831);
or UO_2759 (O_2759,N_24992,N_24948);
or UO_2760 (O_2760,N_24982,N_24979);
nand UO_2761 (O_2761,N_24844,N_24878);
or UO_2762 (O_2762,N_24901,N_24921);
or UO_2763 (O_2763,N_24770,N_24973);
nand UO_2764 (O_2764,N_24782,N_24965);
and UO_2765 (O_2765,N_24850,N_24852);
nor UO_2766 (O_2766,N_24960,N_24847);
nand UO_2767 (O_2767,N_24896,N_24933);
nand UO_2768 (O_2768,N_24997,N_24809);
or UO_2769 (O_2769,N_24812,N_24940);
or UO_2770 (O_2770,N_24773,N_24753);
nand UO_2771 (O_2771,N_24780,N_24986);
nor UO_2772 (O_2772,N_24795,N_24997);
or UO_2773 (O_2773,N_24814,N_24994);
nor UO_2774 (O_2774,N_24838,N_24850);
nand UO_2775 (O_2775,N_24938,N_24953);
nand UO_2776 (O_2776,N_24919,N_24906);
nand UO_2777 (O_2777,N_24755,N_24842);
nand UO_2778 (O_2778,N_24845,N_24798);
nand UO_2779 (O_2779,N_24947,N_24832);
nand UO_2780 (O_2780,N_24856,N_24882);
and UO_2781 (O_2781,N_24975,N_24968);
nand UO_2782 (O_2782,N_24813,N_24886);
nor UO_2783 (O_2783,N_24847,N_24781);
nand UO_2784 (O_2784,N_24811,N_24964);
nor UO_2785 (O_2785,N_24777,N_24751);
xnor UO_2786 (O_2786,N_24851,N_24865);
and UO_2787 (O_2787,N_24763,N_24875);
or UO_2788 (O_2788,N_24903,N_24971);
nand UO_2789 (O_2789,N_24752,N_24855);
xor UO_2790 (O_2790,N_24805,N_24769);
nor UO_2791 (O_2791,N_24834,N_24850);
and UO_2792 (O_2792,N_24922,N_24841);
xnor UO_2793 (O_2793,N_24800,N_24976);
xnor UO_2794 (O_2794,N_24895,N_24870);
nand UO_2795 (O_2795,N_24853,N_24932);
and UO_2796 (O_2796,N_24836,N_24963);
nand UO_2797 (O_2797,N_24789,N_24849);
xor UO_2798 (O_2798,N_24783,N_24904);
nand UO_2799 (O_2799,N_24940,N_24802);
nand UO_2800 (O_2800,N_24918,N_24972);
nor UO_2801 (O_2801,N_24890,N_24954);
nor UO_2802 (O_2802,N_24788,N_24803);
or UO_2803 (O_2803,N_24982,N_24934);
nor UO_2804 (O_2804,N_24864,N_24965);
or UO_2805 (O_2805,N_24982,N_24863);
xor UO_2806 (O_2806,N_24983,N_24893);
or UO_2807 (O_2807,N_24865,N_24778);
nor UO_2808 (O_2808,N_24942,N_24787);
nor UO_2809 (O_2809,N_24871,N_24803);
nand UO_2810 (O_2810,N_24882,N_24876);
nand UO_2811 (O_2811,N_24886,N_24796);
nand UO_2812 (O_2812,N_24825,N_24982);
and UO_2813 (O_2813,N_24847,N_24806);
nor UO_2814 (O_2814,N_24780,N_24862);
nand UO_2815 (O_2815,N_24812,N_24868);
or UO_2816 (O_2816,N_24810,N_24854);
nand UO_2817 (O_2817,N_24995,N_24998);
nor UO_2818 (O_2818,N_24808,N_24891);
nor UO_2819 (O_2819,N_24866,N_24988);
and UO_2820 (O_2820,N_24887,N_24892);
and UO_2821 (O_2821,N_24763,N_24991);
or UO_2822 (O_2822,N_24902,N_24979);
nor UO_2823 (O_2823,N_24992,N_24825);
xor UO_2824 (O_2824,N_24787,N_24904);
or UO_2825 (O_2825,N_24911,N_24902);
nand UO_2826 (O_2826,N_24903,N_24898);
nor UO_2827 (O_2827,N_24925,N_24846);
xor UO_2828 (O_2828,N_24872,N_24889);
nand UO_2829 (O_2829,N_24791,N_24903);
and UO_2830 (O_2830,N_24887,N_24821);
or UO_2831 (O_2831,N_24768,N_24983);
or UO_2832 (O_2832,N_24860,N_24770);
nand UO_2833 (O_2833,N_24825,N_24881);
and UO_2834 (O_2834,N_24768,N_24766);
xnor UO_2835 (O_2835,N_24901,N_24868);
nand UO_2836 (O_2836,N_24908,N_24804);
nand UO_2837 (O_2837,N_24799,N_24966);
xnor UO_2838 (O_2838,N_24776,N_24772);
nor UO_2839 (O_2839,N_24773,N_24937);
xor UO_2840 (O_2840,N_24902,N_24987);
and UO_2841 (O_2841,N_24961,N_24830);
and UO_2842 (O_2842,N_24938,N_24883);
and UO_2843 (O_2843,N_24899,N_24906);
and UO_2844 (O_2844,N_24904,N_24875);
nor UO_2845 (O_2845,N_24853,N_24807);
xor UO_2846 (O_2846,N_24941,N_24920);
xor UO_2847 (O_2847,N_24921,N_24841);
and UO_2848 (O_2848,N_24860,N_24751);
nor UO_2849 (O_2849,N_24961,N_24775);
nand UO_2850 (O_2850,N_24992,N_24845);
xnor UO_2851 (O_2851,N_24819,N_24997);
nor UO_2852 (O_2852,N_24913,N_24979);
or UO_2853 (O_2853,N_24952,N_24801);
and UO_2854 (O_2854,N_24916,N_24855);
nand UO_2855 (O_2855,N_24847,N_24834);
nand UO_2856 (O_2856,N_24767,N_24978);
nand UO_2857 (O_2857,N_24801,N_24940);
and UO_2858 (O_2858,N_24751,N_24863);
xnor UO_2859 (O_2859,N_24757,N_24851);
and UO_2860 (O_2860,N_24879,N_24782);
and UO_2861 (O_2861,N_24873,N_24847);
and UO_2862 (O_2862,N_24950,N_24966);
nor UO_2863 (O_2863,N_24782,N_24952);
nor UO_2864 (O_2864,N_24923,N_24835);
xnor UO_2865 (O_2865,N_24965,N_24976);
and UO_2866 (O_2866,N_24815,N_24882);
nand UO_2867 (O_2867,N_24805,N_24979);
xnor UO_2868 (O_2868,N_24765,N_24939);
and UO_2869 (O_2869,N_24774,N_24880);
and UO_2870 (O_2870,N_24896,N_24801);
and UO_2871 (O_2871,N_24818,N_24848);
and UO_2872 (O_2872,N_24866,N_24927);
and UO_2873 (O_2873,N_24990,N_24898);
or UO_2874 (O_2874,N_24838,N_24767);
nor UO_2875 (O_2875,N_24904,N_24884);
nand UO_2876 (O_2876,N_24935,N_24751);
nand UO_2877 (O_2877,N_24754,N_24835);
nor UO_2878 (O_2878,N_24846,N_24957);
or UO_2879 (O_2879,N_24904,N_24948);
or UO_2880 (O_2880,N_24923,N_24828);
nor UO_2881 (O_2881,N_24913,N_24774);
nor UO_2882 (O_2882,N_24990,N_24956);
nor UO_2883 (O_2883,N_24907,N_24764);
nand UO_2884 (O_2884,N_24905,N_24824);
nor UO_2885 (O_2885,N_24871,N_24816);
nor UO_2886 (O_2886,N_24833,N_24947);
and UO_2887 (O_2887,N_24872,N_24800);
xor UO_2888 (O_2888,N_24856,N_24839);
nor UO_2889 (O_2889,N_24822,N_24941);
nand UO_2890 (O_2890,N_24856,N_24940);
nand UO_2891 (O_2891,N_24796,N_24966);
and UO_2892 (O_2892,N_24862,N_24783);
xor UO_2893 (O_2893,N_24941,N_24878);
nand UO_2894 (O_2894,N_24772,N_24894);
or UO_2895 (O_2895,N_24935,N_24938);
nor UO_2896 (O_2896,N_24882,N_24859);
nand UO_2897 (O_2897,N_24875,N_24921);
nor UO_2898 (O_2898,N_24967,N_24799);
or UO_2899 (O_2899,N_24838,N_24883);
or UO_2900 (O_2900,N_24803,N_24752);
nand UO_2901 (O_2901,N_24786,N_24801);
xor UO_2902 (O_2902,N_24875,N_24936);
and UO_2903 (O_2903,N_24779,N_24880);
nor UO_2904 (O_2904,N_24866,N_24990);
nand UO_2905 (O_2905,N_24995,N_24819);
or UO_2906 (O_2906,N_24951,N_24803);
nand UO_2907 (O_2907,N_24894,N_24751);
and UO_2908 (O_2908,N_24850,N_24849);
and UO_2909 (O_2909,N_24803,N_24921);
nand UO_2910 (O_2910,N_24856,N_24798);
or UO_2911 (O_2911,N_24950,N_24848);
and UO_2912 (O_2912,N_24917,N_24994);
or UO_2913 (O_2913,N_24760,N_24993);
nor UO_2914 (O_2914,N_24833,N_24975);
or UO_2915 (O_2915,N_24793,N_24952);
nor UO_2916 (O_2916,N_24888,N_24769);
xor UO_2917 (O_2917,N_24837,N_24908);
nand UO_2918 (O_2918,N_24774,N_24988);
xnor UO_2919 (O_2919,N_24897,N_24850);
nand UO_2920 (O_2920,N_24946,N_24816);
and UO_2921 (O_2921,N_24850,N_24943);
xnor UO_2922 (O_2922,N_24950,N_24930);
or UO_2923 (O_2923,N_24839,N_24761);
or UO_2924 (O_2924,N_24809,N_24868);
nand UO_2925 (O_2925,N_24790,N_24888);
nor UO_2926 (O_2926,N_24754,N_24959);
and UO_2927 (O_2927,N_24810,N_24956);
and UO_2928 (O_2928,N_24844,N_24754);
or UO_2929 (O_2929,N_24868,N_24847);
nor UO_2930 (O_2930,N_24891,N_24921);
and UO_2931 (O_2931,N_24763,N_24879);
and UO_2932 (O_2932,N_24948,N_24913);
nor UO_2933 (O_2933,N_24994,N_24825);
nand UO_2934 (O_2934,N_24892,N_24903);
nor UO_2935 (O_2935,N_24868,N_24879);
nand UO_2936 (O_2936,N_24837,N_24893);
nor UO_2937 (O_2937,N_24904,N_24911);
or UO_2938 (O_2938,N_24978,N_24817);
nor UO_2939 (O_2939,N_24755,N_24754);
and UO_2940 (O_2940,N_24869,N_24890);
nor UO_2941 (O_2941,N_24939,N_24794);
xor UO_2942 (O_2942,N_24886,N_24865);
nor UO_2943 (O_2943,N_24914,N_24752);
xor UO_2944 (O_2944,N_24930,N_24987);
and UO_2945 (O_2945,N_24853,N_24841);
or UO_2946 (O_2946,N_24848,N_24829);
nand UO_2947 (O_2947,N_24790,N_24856);
or UO_2948 (O_2948,N_24988,N_24969);
and UO_2949 (O_2949,N_24872,N_24780);
or UO_2950 (O_2950,N_24901,N_24785);
nor UO_2951 (O_2951,N_24808,N_24801);
nand UO_2952 (O_2952,N_24904,N_24958);
or UO_2953 (O_2953,N_24888,N_24902);
and UO_2954 (O_2954,N_24865,N_24810);
and UO_2955 (O_2955,N_24900,N_24797);
or UO_2956 (O_2956,N_24883,N_24873);
or UO_2957 (O_2957,N_24811,N_24792);
and UO_2958 (O_2958,N_24897,N_24914);
nand UO_2959 (O_2959,N_24863,N_24777);
or UO_2960 (O_2960,N_24970,N_24963);
nor UO_2961 (O_2961,N_24862,N_24789);
nor UO_2962 (O_2962,N_24906,N_24996);
and UO_2963 (O_2963,N_24841,N_24836);
nand UO_2964 (O_2964,N_24804,N_24838);
and UO_2965 (O_2965,N_24948,N_24880);
xor UO_2966 (O_2966,N_24783,N_24873);
nor UO_2967 (O_2967,N_24859,N_24775);
and UO_2968 (O_2968,N_24860,N_24881);
or UO_2969 (O_2969,N_24861,N_24859);
and UO_2970 (O_2970,N_24805,N_24815);
xnor UO_2971 (O_2971,N_24958,N_24975);
nor UO_2972 (O_2972,N_24921,N_24894);
and UO_2973 (O_2973,N_24949,N_24816);
or UO_2974 (O_2974,N_24823,N_24799);
xor UO_2975 (O_2975,N_24813,N_24978);
or UO_2976 (O_2976,N_24954,N_24821);
xnor UO_2977 (O_2977,N_24751,N_24806);
and UO_2978 (O_2978,N_24904,N_24974);
nand UO_2979 (O_2979,N_24772,N_24936);
or UO_2980 (O_2980,N_24818,N_24943);
nor UO_2981 (O_2981,N_24756,N_24880);
nor UO_2982 (O_2982,N_24786,N_24756);
nand UO_2983 (O_2983,N_24863,N_24764);
or UO_2984 (O_2984,N_24858,N_24945);
nor UO_2985 (O_2985,N_24922,N_24969);
or UO_2986 (O_2986,N_24868,N_24950);
nor UO_2987 (O_2987,N_24842,N_24791);
nor UO_2988 (O_2988,N_24896,N_24758);
nor UO_2989 (O_2989,N_24936,N_24939);
nand UO_2990 (O_2990,N_24891,N_24768);
or UO_2991 (O_2991,N_24772,N_24847);
nand UO_2992 (O_2992,N_24949,N_24970);
and UO_2993 (O_2993,N_24927,N_24773);
or UO_2994 (O_2994,N_24903,N_24852);
and UO_2995 (O_2995,N_24855,N_24872);
or UO_2996 (O_2996,N_24974,N_24770);
and UO_2997 (O_2997,N_24960,N_24761);
nor UO_2998 (O_2998,N_24789,N_24994);
xor UO_2999 (O_2999,N_24935,N_24859);
endmodule