module basic_2500_25000_3000_50_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_885,In_1944);
or U1 (N_1,In_1545,In_1660);
xor U2 (N_2,In_2478,In_1299);
or U3 (N_3,In_1678,In_1136);
or U4 (N_4,In_792,In_567);
nor U5 (N_5,In_149,In_1684);
nand U6 (N_6,In_2017,In_535);
and U7 (N_7,In_1329,In_2000);
nand U8 (N_8,In_112,In_846);
or U9 (N_9,In_1594,In_732);
or U10 (N_10,In_2497,In_600);
and U11 (N_11,In_1906,In_2084);
nand U12 (N_12,In_1346,In_801);
or U13 (N_13,In_1544,In_1367);
or U14 (N_14,In_887,In_1952);
and U15 (N_15,In_1252,In_849);
or U16 (N_16,In_890,In_1664);
or U17 (N_17,In_1873,In_1498);
xor U18 (N_18,In_2149,In_2254);
xnor U19 (N_19,In_652,In_314);
xnor U20 (N_20,In_2318,In_1358);
or U21 (N_21,In_1776,In_1300);
nor U22 (N_22,In_2447,In_568);
or U23 (N_23,In_1059,In_627);
nor U24 (N_24,In_2082,In_2422);
nor U25 (N_25,In_28,In_2044);
nand U26 (N_26,In_857,In_1224);
nand U27 (N_27,In_827,In_2411);
and U28 (N_28,In_1649,In_2224);
nand U29 (N_29,In_1117,In_2288);
and U30 (N_30,In_2294,In_1128);
or U31 (N_31,In_223,In_1953);
and U32 (N_32,In_2233,In_1641);
and U33 (N_33,In_2413,In_2186);
xor U34 (N_34,In_823,In_1663);
nand U35 (N_35,In_1854,In_984);
nor U36 (N_36,In_166,In_2326);
or U37 (N_37,In_1580,In_1824);
nor U38 (N_38,In_1942,In_411);
or U39 (N_39,In_144,In_1523);
xnor U40 (N_40,In_1303,In_327);
nor U41 (N_41,In_863,In_2457);
and U42 (N_42,In_2299,In_1880);
or U43 (N_43,In_2496,In_1898);
or U44 (N_44,In_444,In_2048);
or U45 (N_45,In_249,In_706);
and U46 (N_46,In_2490,In_2062);
nor U47 (N_47,In_501,In_1782);
or U48 (N_48,In_2032,In_1085);
or U49 (N_49,In_992,In_1381);
nand U50 (N_50,In_80,In_2260);
xnor U51 (N_51,In_796,In_1807);
nand U52 (N_52,In_2386,In_991);
or U53 (N_53,In_1628,In_879);
and U54 (N_54,In_313,In_2414);
xor U55 (N_55,In_1899,In_243);
xnor U56 (N_56,In_531,In_2453);
nand U57 (N_57,In_898,In_919);
or U58 (N_58,In_613,In_458);
nand U59 (N_59,In_945,In_23);
and U60 (N_60,In_2025,In_1861);
xor U61 (N_61,In_596,In_1020);
nor U62 (N_62,In_953,In_1486);
nor U63 (N_63,In_145,In_227);
nand U64 (N_64,In_1493,In_921);
nor U65 (N_65,In_2402,In_477);
nand U66 (N_66,In_1240,In_549);
nor U67 (N_67,In_1796,In_304);
xnor U68 (N_68,In_384,In_321);
and U69 (N_69,In_1399,In_33);
xnor U70 (N_70,In_32,In_641);
nand U71 (N_71,In_1140,In_2416);
or U72 (N_72,In_1410,In_1394);
nor U73 (N_73,In_2070,In_968);
nand U74 (N_74,In_1420,In_632);
nor U75 (N_75,In_1264,In_1558);
nand U76 (N_76,In_2107,In_1222);
and U77 (N_77,In_680,In_675);
nand U78 (N_78,In_1078,In_1166);
xor U79 (N_79,In_1500,In_664);
and U80 (N_80,In_2470,In_462);
nand U81 (N_81,In_1855,In_540);
nand U82 (N_82,In_1791,In_2383);
and U83 (N_83,In_1368,In_258);
xor U84 (N_84,In_2367,In_744);
or U85 (N_85,In_1588,In_1835);
xnor U86 (N_86,In_1050,In_2006);
or U87 (N_87,In_579,In_1075);
nor U88 (N_88,In_2214,In_2273);
xor U89 (N_89,In_2344,In_2170);
and U90 (N_90,In_790,In_1276);
nor U91 (N_91,In_193,In_1245);
or U92 (N_92,In_2406,In_181);
xor U93 (N_93,In_563,In_560);
nand U94 (N_94,In_785,In_2353);
and U95 (N_95,In_1654,In_688);
or U96 (N_96,In_2218,In_939);
nand U97 (N_97,In_2251,In_1675);
or U98 (N_98,In_1168,In_1055);
xor U99 (N_99,In_1056,In_2161);
nand U100 (N_100,In_1863,In_301);
nor U101 (N_101,In_2494,In_1416);
xor U102 (N_102,In_50,In_1097);
and U103 (N_103,In_1562,In_246);
and U104 (N_104,In_491,In_781);
nand U105 (N_105,In_1135,In_377);
xnor U106 (N_106,In_189,In_917);
nand U107 (N_107,In_1821,In_693);
nor U108 (N_108,In_427,In_753);
xor U109 (N_109,In_331,In_1503);
and U110 (N_110,In_1271,In_2271);
and U111 (N_111,In_1865,In_502);
and U112 (N_112,In_2142,In_867);
and U113 (N_113,In_1816,In_1029);
nand U114 (N_114,In_2210,In_1054);
nor U115 (N_115,In_1871,In_928);
and U116 (N_116,In_2162,In_194);
and U117 (N_117,In_1449,In_2136);
xnor U118 (N_118,In_1572,In_714);
and U119 (N_119,In_1391,In_2340);
and U120 (N_120,In_668,In_1279);
xnor U121 (N_121,In_281,In_683);
xor U122 (N_122,In_1062,In_2369);
nand U123 (N_123,In_320,In_87);
or U124 (N_124,In_1469,In_387);
and U125 (N_125,In_816,In_264);
nand U126 (N_126,In_1255,In_15);
or U127 (N_127,In_2141,In_1908);
nor U128 (N_128,In_1687,In_2331);
or U129 (N_129,In_982,In_230);
nor U130 (N_130,In_1784,In_2325);
or U131 (N_131,In_2019,In_2235);
and U132 (N_132,In_1987,In_2349);
and U133 (N_133,In_1444,In_1378);
or U134 (N_134,In_1762,In_963);
nor U135 (N_135,In_1602,In_908);
and U136 (N_136,In_2272,In_682);
nor U137 (N_137,In_2315,In_1370);
xnor U138 (N_138,In_432,In_68);
xor U139 (N_139,In_94,In_2259);
nor U140 (N_140,In_2289,In_1016);
and U141 (N_141,In_359,In_83);
nor U142 (N_142,In_390,In_1120);
xor U143 (N_143,In_186,In_2421);
nand U144 (N_144,In_1830,In_2092);
and U145 (N_145,In_1984,In_2011);
nand U146 (N_146,In_481,In_455);
or U147 (N_147,In_97,In_1977);
and U148 (N_148,In_2089,In_1696);
nor U149 (N_149,In_161,In_190);
xnor U150 (N_150,In_978,In_875);
nor U151 (N_151,In_2439,In_2454);
nand U152 (N_152,In_1199,In_860);
or U153 (N_153,In_242,In_1635);
nor U154 (N_154,In_1215,In_370);
nor U155 (N_155,In_392,In_39);
xnor U156 (N_156,In_1212,In_1905);
xor U157 (N_157,In_2231,In_1439);
and U158 (N_158,In_2042,In_957);
nand U159 (N_159,In_2074,In_736);
and U160 (N_160,In_1430,In_2035);
and U161 (N_161,In_1917,In_1126);
xnor U162 (N_162,In_226,In_2018);
xnor U163 (N_163,In_1686,In_1210);
and U164 (N_164,In_1341,In_1526);
and U165 (N_165,In_1886,In_1488);
xor U166 (N_166,In_891,In_2459);
nor U167 (N_167,In_2373,In_1448);
nand U168 (N_168,In_2007,In_920);
and U169 (N_169,In_1291,In_1679);
xnor U170 (N_170,In_904,In_374);
xnor U171 (N_171,In_1682,In_834);
or U172 (N_172,In_2088,In_2250);
or U173 (N_173,In_804,In_1094);
nand U174 (N_174,In_1067,In_1384);
or U175 (N_175,In_914,In_2319);
and U176 (N_176,In_1071,In_947);
and U177 (N_177,In_2311,In_1661);
xnor U178 (N_178,In_625,In_2185);
nand U179 (N_179,In_1313,In_1936);
or U180 (N_180,In_1389,In_578);
and U181 (N_181,In_752,In_2352);
xnor U182 (N_182,In_1709,In_1304);
xor U183 (N_183,In_1284,In_154);
and U184 (N_184,In_1758,In_1318);
or U185 (N_185,In_188,In_1233);
xnor U186 (N_186,In_1667,In_1322);
or U187 (N_187,In_260,In_2203);
and U188 (N_188,In_218,In_1465);
nor U189 (N_189,In_40,In_2304);
or U190 (N_190,In_332,In_1744);
and U191 (N_191,In_2206,In_2366);
nand U192 (N_192,In_761,In_287);
and U193 (N_193,In_2041,In_813);
nand U194 (N_194,In_585,In_107);
xnor U195 (N_195,In_141,In_1433);
xor U196 (N_196,In_1194,In_415);
nand U197 (N_197,In_1676,In_2105);
nand U198 (N_198,In_1819,In_1750);
and U199 (N_199,In_487,In_912);
nand U200 (N_200,In_1283,In_1575);
nand U201 (N_201,In_2390,In_1520);
nand U202 (N_202,In_1539,In_1866);
or U203 (N_203,In_1999,In_2342);
xnor U204 (N_204,In_1721,In_588);
xnor U205 (N_205,In_453,In_129);
or U206 (N_206,In_2111,In_811);
nor U207 (N_207,In_256,In_2365);
and U208 (N_208,In_967,In_1958);
nand U209 (N_209,In_835,In_864);
nor U210 (N_210,In_2110,In_2266);
or U211 (N_211,In_508,In_2347);
nor U212 (N_212,In_2096,In_105);
nand U213 (N_213,In_1738,In_770);
or U214 (N_214,In_2443,In_419);
nand U215 (N_215,In_1096,In_1243);
and U216 (N_216,In_1200,In_1447);
nand U217 (N_217,In_1306,In_2090);
nor U218 (N_218,In_2119,In_1841);
xnor U219 (N_219,In_1557,In_674);
nor U220 (N_220,In_323,In_1805);
or U221 (N_221,In_1175,In_412);
nor U222 (N_222,In_1177,In_608);
nand U223 (N_223,In_335,In_1388);
xnor U224 (N_224,In_1730,In_883);
or U225 (N_225,In_56,In_751);
or U226 (N_226,In_704,In_1357);
and U227 (N_227,In_1044,In_1251);
or U228 (N_228,In_1955,In_2465);
nor U229 (N_229,In_1006,In_1728);
nor U230 (N_230,In_926,In_1141);
or U231 (N_231,In_820,In_768);
and U232 (N_232,In_1543,In_728);
and U233 (N_233,In_2431,In_213);
or U234 (N_234,In_1561,In_818);
xor U235 (N_235,In_1962,In_956);
or U236 (N_236,In_584,In_372);
nor U237 (N_237,In_1147,In_470);
xor U238 (N_238,In_1483,In_1292);
xnor U239 (N_239,In_2243,In_303);
and U240 (N_240,In_1169,In_1626);
nor U241 (N_241,In_1497,In_2472);
nand U242 (N_242,In_29,In_1481);
nand U243 (N_243,In_143,In_70);
or U244 (N_244,In_1307,In_1302);
nor U245 (N_245,In_689,In_9);
and U246 (N_246,In_1531,In_155);
and U247 (N_247,In_559,In_1174);
xor U248 (N_248,In_763,In_1751);
nand U249 (N_249,In_2063,In_649);
xor U250 (N_250,In_999,In_643);
xnor U251 (N_251,In_20,In_2069);
or U252 (N_252,In_289,In_398);
nor U253 (N_253,In_1845,In_697);
and U254 (N_254,In_2002,In_1301);
and U255 (N_255,In_833,In_1473);
and U256 (N_256,In_1574,In_429);
nor U257 (N_257,In_2473,In_1643);
and U258 (N_258,In_1797,In_1564);
xnor U259 (N_259,In_1928,In_1004);
xnor U260 (N_260,In_1220,In_483);
xnor U261 (N_261,In_1515,In_1765);
nand U262 (N_262,In_1030,In_1221);
or U263 (N_263,In_2312,In_2479);
nand U264 (N_264,In_21,In_134);
nand U265 (N_265,In_1009,In_1812);
nor U266 (N_266,In_1691,In_1773);
xor U267 (N_267,In_1184,In_1074);
or U268 (N_268,In_285,In_117);
and U269 (N_269,In_77,In_2179);
nor U270 (N_270,In_1804,In_1436);
nor U271 (N_271,In_2424,In_205);
nand U272 (N_272,In_2392,In_2085);
xor U273 (N_273,In_1487,In_871);
and U274 (N_274,In_1429,In_308);
nand U275 (N_275,In_402,In_182);
nor U276 (N_276,In_2056,In_1069);
and U277 (N_277,In_355,In_1450);
and U278 (N_278,In_1619,In_2121);
or U279 (N_279,In_1235,In_1522);
nor U280 (N_280,In_1423,In_164);
or U281 (N_281,In_1530,In_36);
nand U282 (N_282,In_1369,In_1193);
and U283 (N_283,In_1008,In_617);
nand U284 (N_284,In_479,In_422);
nand U285 (N_285,In_1441,In_1716);
and U286 (N_286,In_2471,In_2122);
or U287 (N_287,In_2464,In_1890);
and U288 (N_288,In_646,In_615);
or U289 (N_289,In_1435,In_1412);
nor U290 (N_290,In_1883,In_1201);
and U291 (N_291,In_272,In_1548);
nand U292 (N_292,In_1010,In_581);
nor U293 (N_293,In_634,In_841);
nand U294 (N_294,In_2396,In_2034);
nand U295 (N_295,In_8,In_99);
xor U296 (N_296,In_1364,In_2348);
and U297 (N_297,In_2225,In_2204);
xnor U298 (N_298,In_1294,In_2112);
and U299 (N_299,In_520,In_1926);
and U300 (N_300,In_2128,In_2008);
xnor U301 (N_301,In_1070,In_1457);
or U302 (N_302,In_2076,In_137);
xor U303 (N_303,In_44,In_1502);
nand U304 (N_304,In_106,In_306);
xnor U305 (N_305,In_1261,In_2219);
and U306 (N_306,In_676,In_1516);
nor U307 (N_307,In_716,In_529);
nor U308 (N_308,In_1223,In_2200);
nand U309 (N_309,In_2387,In_1556);
nand U310 (N_310,In_211,In_1767);
and U311 (N_311,In_2426,In_448);
nand U312 (N_312,In_2481,In_1099);
nor U313 (N_313,In_4,In_525);
or U314 (N_314,In_337,In_2238);
nor U315 (N_315,In_2135,In_2);
xor U316 (N_316,In_397,In_1553);
and U317 (N_317,In_2058,In_1338);
or U318 (N_318,In_428,In_1312);
nor U319 (N_319,In_1589,In_1823);
nor U320 (N_320,In_27,In_1756);
nor U321 (N_321,In_973,In_1287);
xnor U322 (N_322,In_1850,In_530);
xor U323 (N_323,In_981,In_1569);
xor U324 (N_324,In_976,In_2079);
nor U325 (N_325,In_234,In_959);
nor U326 (N_326,In_1024,In_812);
or U327 (N_327,In_565,In_2316);
nand U328 (N_328,In_2242,In_1012);
nand U329 (N_329,In_271,In_1528);
xnor U330 (N_330,In_52,In_612);
or U331 (N_331,In_71,In_279);
nor U332 (N_332,In_899,In_558);
and U333 (N_333,In_1134,In_2480);
nor U334 (N_334,In_1615,In_1525);
xor U335 (N_335,In_1783,In_78);
nor U336 (N_336,In_366,In_1419);
or U337 (N_337,In_730,In_644);
nand U338 (N_338,In_1249,In_1072);
or U339 (N_339,In_780,In_1968);
xnor U340 (N_340,In_880,In_747);
or U341 (N_341,In_620,In_430);
and U342 (N_342,In_7,In_2484);
nand U343 (N_343,In_268,In_1809);
xnor U344 (N_344,In_1554,In_2038);
nor U345 (N_345,In_1409,In_1081);
or U346 (N_346,In_2449,In_1670);
and U347 (N_347,In_170,In_865);
or U348 (N_348,In_894,In_651);
nor U349 (N_349,In_1646,In_1013);
nor U350 (N_350,In_2292,In_2160);
or U351 (N_351,In_1327,In_1757);
nand U352 (N_352,In_379,In_1725);
nand U353 (N_353,In_1598,In_1295);
nor U354 (N_354,In_1417,In_1965);
xnor U355 (N_355,In_687,In_711);
nand U356 (N_356,In_1701,In_2418);
nand U357 (N_357,In_1887,In_2381);
or U358 (N_358,In_409,In_310);
or U359 (N_359,In_431,In_124);
xnor U360 (N_360,In_489,In_292);
nor U361 (N_361,In_2337,In_1242);
and U362 (N_362,In_616,In_1837);
nand U363 (N_363,In_179,In_37);
nor U364 (N_364,In_439,In_977);
and U365 (N_365,In_156,In_1902);
or U366 (N_366,In_1014,In_1188);
xnor U367 (N_367,In_1191,In_929);
and U368 (N_368,In_1155,In_576);
nand U369 (N_369,In_881,In_1);
or U370 (N_370,In_802,In_1546);
nor U371 (N_371,In_1133,In_807);
xor U372 (N_372,In_2169,In_1624);
nand U373 (N_373,In_2430,In_2498);
nand U374 (N_374,In_1142,In_72);
or U375 (N_375,In_1238,In_2216);
or U376 (N_376,In_2215,In_1610);
and U377 (N_377,In_266,In_510);
nand U378 (N_378,In_1086,In_1510);
nand U379 (N_379,In_2223,In_2336);
nand U380 (N_380,In_425,In_1495);
nor U381 (N_381,In_2379,In_1157);
xnor U382 (N_382,In_533,In_1180);
nor U383 (N_383,In_449,In_1179);
nor U384 (N_384,In_421,In_416);
xor U385 (N_385,In_361,In_1404);
nor U386 (N_386,In_941,In_2274);
nor U387 (N_387,In_1335,In_269);
and U388 (N_388,In_356,In_426);
or U389 (N_389,In_1743,In_1467);
nand U390 (N_390,In_325,In_1559);
xnor U391 (N_391,In_1266,In_1914);
nor U392 (N_392,In_657,In_441);
xnor U393 (N_393,In_1951,In_614);
nor U394 (N_394,In_760,In_1361);
or U395 (N_395,In_666,In_2207);
nor U396 (N_396,In_2239,In_2059);
or U397 (N_397,In_2358,In_532);
or U398 (N_398,In_451,In_1098);
xnor U399 (N_399,In_1470,In_962);
nor U400 (N_400,In_2033,In_798);
nand U401 (N_401,In_89,In_2094);
or U402 (N_402,In_707,In_2346);
nor U403 (N_403,In_1337,In_2176);
xnor U404 (N_404,In_197,In_14);
or U405 (N_405,In_1428,In_2361);
or U406 (N_406,In_2248,In_1395);
xor U407 (N_407,In_1285,In_1342);
or U408 (N_408,In_645,In_1456);
nor U409 (N_409,In_2165,In_284);
nor U410 (N_410,In_1480,In_836);
and U411 (N_411,In_1036,In_1981);
or U412 (N_412,In_1183,In_1611);
or U413 (N_413,In_173,In_2098);
or U414 (N_414,In_1267,In_1256);
and U415 (N_415,In_870,In_862);
nand U416 (N_416,In_153,In_2435);
nor U417 (N_417,In_2244,In_577);
nor U418 (N_418,In_438,In_2351);
and U419 (N_419,In_2305,In_858);
nand U420 (N_420,In_74,In_1627);
xnor U421 (N_421,In_2404,In_199);
nor U422 (N_422,In_2345,In_2043);
and U423 (N_423,In_690,In_1724);
xor U424 (N_424,In_949,In_1132);
nand U425 (N_425,In_1407,In_1365);
and U426 (N_426,In_618,In_930);
or U427 (N_427,In_866,In_878);
and U428 (N_428,In_2287,In_2436);
nor U429 (N_429,In_1351,In_964);
nor U430 (N_430,In_1974,In_1786);
nand U431 (N_431,In_1262,In_1669);
nand U432 (N_432,In_60,In_1032);
nor U433 (N_433,In_2317,In_2129);
nor U434 (N_434,In_1088,In_2145);
or U435 (N_435,In_1277,In_1241);
nor U436 (N_436,In_1232,In_1954);
nor U437 (N_437,In_1512,In_731);
or U438 (N_438,In_2495,In_1167);
or U439 (N_439,In_1801,In_2320);
nor U440 (N_440,In_1061,In_1550);
or U441 (N_441,In_2014,In_906);
xnor U442 (N_442,In_2055,In_1258);
and U443 (N_443,In_130,In_1702);
xnor U444 (N_444,In_2157,In_1431);
nand U445 (N_445,In_2073,In_622);
xnor U446 (N_446,In_1889,In_1021);
nand U447 (N_447,In_1053,In_1655);
or U448 (N_448,In_270,In_47);
nand U449 (N_449,In_1315,In_737);
or U450 (N_450,In_126,In_373);
xnor U451 (N_451,In_2211,In_1959);
nor U452 (N_452,In_1826,In_1604);
or U453 (N_453,In_1403,In_1349);
nand U454 (N_454,In_1163,In_1496);
xnor U455 (N_455,In_1025,In_286);
or U456 (N_456,In_461,In_1460);
or U457 (N_457,In_975,In_2020);
nor U458 (N_458,In_1991,In_1218);
nand U459 (N_459,In_670,In_1415);
and U460 (N_460,In_831,In_165);
nand U461 (N_461,In_342,In_989);
xor U462 (N_462,In_1396,In_282);
and U463 (N_463,In_2068,In_1386);
and U464 (N_464,In_66,In_278);
or U465 (N_465,In_980,In_609);
nor U466 (N_466,In_1585,In_803);
or U467 (N_467,In_1379,In_913);
or U468 (N_468,In_903,In_376);
or U469 (N_469,In_2280,In_1688);
or U470 (N_470,In_2137,In_2049);
nand U471 (N_471,In_1446,In_1633);
and U472 (N_472,In_273,In_556);
xnor U473 (N_473,In_897,In_2016);
and U474 (N_474,In_1583,In_1001);
xnor U475 (N_475,In_1461,In_1706);
nand U476 (N_476,In_809,In_248);
and U477 (N_477,In_2201,In_2183);
nand U478 (N_478,In_2477,In_659);
or U479 (N_479,In_54,In_315);
or U480 (N_480,In_678,In_2362);
nor U481 (N_481,In_497,In_316);
and U482 (N_482,In_1930,In_1031);
xor U483 (N_483,In_1995,In_2419);
or U484 (N_484,In_966,In_944);
nor U485 (N_485,In_1197,In_102);
nand U486 (N_486,In_1631,In_696);
xor U487 (N_487,In_2037,In_1625);
or U488 (N_488,In_515,In_892);
nor U489 (N_489,In_168,In_2232);
and U490 (N_490,In_405,In_985);
or U491 (N_491,In_10,In_1411);
or U492 (N_492,In_420,In_2103);
or U493 (N_493,In_305,In_460);
nor U494 (N_494,In_1376,In_597);
or U495 (N_495,In_1216,In_538);
nor U496 (N_496,In_326,In_786);
or U497 (N_497,In_553,In_2022);
nand U498 (N_498,In_773,In_2117);
nand U499 (N_499,In_2448,In_853);
or U500 (N_500,N_402,In_1173);
xor U501 (N_501,In_2188,In_1362);
and U502 (N_502,In_950,In_1116);
or U503 (N_503,In_67,In_2338);
and U504 (N_504,N_233,In_1219);
or U505 (N_505,In_772,In_200);
nand U506 (N_506,In_395,In_2335);
xor U507 (N_507,N_330,N_77);
nor U508 (N_508,In_2212,In_485);
or U509 (N_509,In_1940,In_2164);
or U510 (N_510,In_2226,N_196);
or U511 (N_511,In_2261,N_444);
and U512 (N_512,N_211,In_237);
or U513 (N_513,In_1761,N_11);
nor U514 (N_514,In_1996,In_1060);
or U515 (N_515,In_127,In_661);
nor U516 (N_516,In_1290,In_1760);
and U517 (N_517,In_1822,In_1039);
or U518 (N_518,In_1372,N_260);
nor U519 (N_519,In_31,In_1969);
nand U520 (N_520,In_723,In_583);
and U521 (N_521,In_1190,In_572);
nand U522 (N_522,In_2168,N_394);
or U523 (N_523,In_2343,In_61);
xnor U524 (N_524,In_136,N_419);
or U525 (N_525,In_1907,In_1288);
and U526 (N_526,In_1002,In_1217);
nand U527 (N_527,N_345,In_1192);
and U528 (N_528,In_1595,In_1492);
or U529 (N_529,In_699,In_109);
nand U530 (N_530,In_2474,In_232);
or U531 (N_531,N_484,N_351);
nor U532 (N_532,N_396,In_598);
xor U533 (N_533,N_372,In_1397);
or U534 (N_534,In_1455,In_217);
nor U535 (N_535,In_1127,N_168);
nand U536 (N_536,In_1269,In_523);
nor U537 (N_537,N_28,N_476);
xor U538 (N_538,N_276,In_1041);
nand U539 (N_539,In_1080,N_89);
nor U540 (N_540,N_438,In_2208);
or U541 (N_541,In_1922,In_1766);
xor U542 (N_542,In_909,In_294);
xor U543 (N_543,In_55,In_1451);
nor U544 (N_544,N_280,N_297);
nor U545 (N_545,In_1236,In_2191);
and U546 (N_546,In_2277,In_17);
nand U547 (N_547,N_442,In_994);
or U548 (N_548,N_127,N_35);
nand U549 (N_549,In_152,In_2228);
and U550 (N_550,In_2067,In_739);
xnor U551 (N_551,In_0,In_2444);
or U552 (N_552,In_745,In_2150);
or U553 (N_553,In_1937,In_1208);
and U554 (N_554,In_2227,In_2040);
nor U555 (N_555,In_825,N_178);
xnor U556 (N_556,N_273,In_222);
or U557 (N_557,In_1947,In_1323);
nor U558 (N_558,N_384,In_1617);
xnor U559 (N_559,In_2125,In_1356);
and U560 (N_560,In_507,In_1375);
nor U561 (N_561,In_1918,In_1909);
xor U562 (N_562,In_1815,In_1110);
nor U563 (N_563,In_1196,In_247);
nor U564 (N_564,N_190,In_2258);
or U565 (N_565,In_764,In_2463);
nand U566 (N_566,In_2154,In_360);
and U567 (N_567,In_2060,In_108);
nand U568 (N_568,In_907,N_482);
xnor U569 (N_569,In_51,In_2407);
nor U570 (N_570,In_1466,In_2360);
nand U571 (N_571,In_115,N_63);
xor U572 (N_572,In_1934,In_73);
nor U573 (N_573,In_1842,N_105);
nor U574 (N_574,In_2051,In_265);
nand U575 (N_575,In_1045,In_424);
nor U576 (N_576,In_1584,In_2302);
nand U577 (N_577,N_201,N_348);
or U578 (N_578,N_392,In_2144);
nand U579 (N_579,N_208,N_468);
and U580 (N_580,In_88,In_79);
xnor U581 (N_581,N_9,In_1103);
and U582 (N_582,In_1405,In_196);
and U583 (N_583,N_346,In_2451);
or U584 (N_584,In_57,In_1714);
nand U585 (N_585,In_1980,In_983);
xnor U586 (N_586,In_1779,In_718);
or U587 (N_587,N_478,In_621);
or U588 (N_588,N_164,In_488);
nand U589 (N_589,In_1671,In_1519);
and U590 (N_590,In_81,In_499);
or U591 (N_591,In_1418,In_974);
or U592 (N_592,In_1875,N_143);
xor U593 (N_593,N_325,N_187);
nand U594 (N_594,In_1272,In_555);
or U595 (N_595,In_844,In_450);
nor U596 (N_596,In_663,In_1745);
xor U597 (N_597,In_1772,N_203);
nand U598 (N_598,N_377,In_1148);
or U599 (N_599,In_219,In_1623);
xnor U600 (N_600,In_2004,In_90);
or U601 (N_601,In_603,In_1317);
or U602 (N_602,In_1535,In_1172);
or U603 (N_603,In_2202,N_207);
nand U604 (N_604,In_362,In_938);
or U605 (N_605,In_1770,In_93);
and U606 (N_606,In_1753,N_184);
nor U607 (N_607,N_61,In_472);
nor U608 (N_608,N_126,N_155);
and U609 (N_609,In_48,N_106);
nor U610 (N_610,In_1113,In_1401);
nor U611 (N_611,In_1434,N_269);
nand U612 (N_612,In_2087,In_1777);
and U613 (N_613,N_461,N_296);
and U614 (N_614,In_1383,N_455);
nand U615 (N_615,In_2275,In_1640);
nand U616 (N_616,In_1281,In_1852);
xor U617 (N_617,In_2264,In_1334);
xor U618 (N_618,N_284,In_2491);
nor U619 (N_619,N_238,In_2120);
xor U620 (N_620,In_2045,In_2341);
or U621 (N_621,In_1160,In_2469);
xor U622 (N_622,In_702,In_2359);
and U623 (N_623,In_2488,In_1833);
or U624 (N_624,In_1393,In_1634);
or U625 (N_625,In_2023,In_1382);
nand U626 (N_626,N_194,N_41);
nand U627 (N_627,In_685,N_191);
nor U628 (N_628,In_2140,In_2339);
nand U629 (N_629,N_424,In_1400);
nand U630 (N_630,N_379,In_936);
nand U631 (N_631,In_979,In_1813);
or U632 (N_632,In_1310,In_1596);
or U633 (N_633,In_469,In_340);
and U634 (N_634,In_2027,In_2247);
xnor U635 (N_635,In_590,In_1653);
or U636 (N_636,In_371,In_5);
xnor U637 (N_637,In_1093,In_175);
and U638 (N_638,N_475,In_1278);
and U639 (N_639,In_1587,In_410);
nor U640 (N_640,In_2196,In_2081);
and U641 (N_641,In_498,In_791);
nor U642 (N_642,In_257,In_1209);
nor U643 (N_643,In_2072,In_1632);
nand U644 (N_644,N_342,N_460);
and U645 (N_645,N_304,N_405);
nand U646 (N_646,In_1567,N_354);
nor U647 (N_647,In_1049,In_684);
nand U648 (N_648,N_339,In_1736);
nand U649 (N_649,In_1943,In_1979);
and U650 (N_650,In_1392,In_1234);
and U651 (N_651,In_2452,In_334);
and U652 (N_652,In_1897,In_1471);
xor U653 (N_653,In_724,In_1884);
xor U654 (N_654,N_366,N_452);
nand U655 (N_655,In_2438,N_485);
nor U656 (N_656,In_1214,In_905);
and U657 (N_657,In_1629,In_1818);
nand U658 (N_658,In_1225,In_1956);
nor U659 (N_659,N_286,In_467);
xnor U660 (N_660,In_26,In_954);
nor U661 (N_661,In_1607,In_838);
xor U662 (N_662,In_970,In_2252);
and U663 (N_663,N_430,In_872);
or U664 (N_664,In_2410,In_1458);
xnor U665 (N_665,In_1058,In_2066);
and U666 (N_666,N_398,In_1836);
nor U667 (N_667,In_354,N_439);
nand U668 (N_668,In_2279,In_214);
xor U669 (N_669,In_307,In_2323);
xnor U670 (N_670,In_2442,N_256);
and U671 (N_671,In_1158,In_2234);
or U672 (N_672,In_2171,N_65);
and U673 (N_673,In_1390,In_1452);
nand U674 (N_674,In_636,N_160);
and U675 (N_675,In_2409,In_333);
nand U676 (N_676,N_270,In_1911);
or U677 (N_677,In_1007,In_463);
or U678 (N_678,In_725,In_1674);
nand U679 (N_679,In_2009,In_43);
nand U680 (N_680,In_1119,In_582);
or U681 (N_681,N_193,In_698);
and U682 (N_682,N_8,In_1923);
xnor U683 (N_683,In_1079,In_1656);
nor U684 (N_684,In_1501,In_746);
or U685 (N_685,In_743,N_267);
nor U686 (N_686,In_45,In_1165);
xor U687 (N_687,N_236,In_2293);
nand U688 (N_688,In_1137,In_2230);
nand U689 (N_689,In_758,In_2205);
and U690 (N_690,In_1939,In_1901);
nand U691 (N_691,N_343,N_363);
or U692 (N_692,In_1989,N_180);
or U693 (N_693,N_380,In_695);
xor U694 (N_694,In_822,In_1414);
and U695 (N_695,In_569,N_298);
and U696 (N_696,In_1933,In_1373);
or U697 (N_697,In_2155,In_1690);
xor U698 (N_698,In_1286,In_1858);
and U699 (N_699,N_282,N_54);
xnor U700 (N_700,In_1839,In_210);
nand U701 (N_701,In_512,In_951);
or U702 (N_702,In_1570,In_662);
xnor U703 (N_703,In_1402,In_404);
xnor U704 (N_704,In_142,In_2077);
nor U705 (N_705,In_1957,In_1340);
xnor U706 (N_706,In_1946,N_213);
or U707 (N_707,N_224,In_1422);
nor U708 (N_708,In_309,In_1432);
and U709 (N_709,In_1665,In_2354);
and U710 (N_710,In_1521,In_208);
and U711 (N_711,N_100,N_358);
or U712 (N_712,N_26,In_1993);
and U713 (N_713,In_2100,In_1354);
xnor U714 (N_714,N_76,In_1637);
or U715 (N_715,In_592,In_1616);
and U716 (N_716,In_277,In_797);
xor U717 (N_717,In_509,In_987);
xor U718 (N_718,In_787,N_432);
nor U719 (N_719,In_1896,N_237);
nand U720 (N_720,In_1840,N_138);
nor U721 (N_721,In_1592,N_150);
or U722 (N_722,N_447,In_2291);
and U723 (N_723,In_1636,In_619);
nand U724 (N_724,In_1159,In_2476);
xor U725 (N_725,In_1028,In_1185);
and U726 (N_726,In_756,N_131);
and U727 (N_727,In_2329,In_1970);
nor U728 (N_728,In_1246,In_861);
and U729 (N_729,In_2330,N_158);
and U730 (N_730,In_1697,In_261);
nand U731 (N_731,In_757,In_806);
nor U732 (N_732,In_64,In_274);
and U733 (N_733,N_285,In_1311);
and U734 (N_734,In_319,N_82);
nor U735 (N_735,In_788,In_1489);
xor U736 (N_736,In_514,In_1352);
or U737 (N_737,In_2286,In_2256);
nand U738 (N_738,In_874,In_1213);
nor U739 (N_739,N_404,In_1095);
xnor U740 (N_740,N_449,In_1967);
nand U741 (N_741,N_483,In_2217);
or U742 (N_742,In_1413,In_774);
and U743 (N_743,In_564,In_1723);
nor U744 (N_744,N_383,In_842);
and U745 (N_745,In_1778,In_2321);
nand U746 (N_746,N_332,In_672);
or U747 (N_747,In_527,In_2499);
xnor U748 (N_748,N_52,In_993);
and U749 (N_749,In_640,In_1862);
and U750 (N_750,In_1344,In_121);
xnor U751 (N_751,In_341,In_925);
nand U752 (N_752,N_313,N_317);
nor U753 (N_753,In_403,N_5);
nand U754 (N_754,In_1527,In_547);
or U755 (N_755,In_2328,In_2270);
and U756 (N_756,In_911,N_374);
and U757 (N_757,In_900,In_562);
nor U758 (N_758,In_13,N_245);
xor U759 (N_759,In_2432,In_1296);
and U760 (N_760,In_1864,In_198);
and U761 (N_761,N_264,In_719);
and U762 (N_762,N_445,N_94);
and U763 (N_763,N_87,In_1207);
nand U764 (N_764,N_251,N_497);
nor U765 (N_765,In_873,In_2123);
xor U766 (N_766,In_96,In_220);
nand U767 (N_767,In_1695,N_353);
or U768 (N_768,In_2395,In_1244);
or U769 (N_769,In_703,N_227);
or U770 (N_770,In_177,In_721);
and U771 (N_771,In_1505,In_1612);
and U772 (N_772,In_2156,In_916);
xor U773 (N_773,N_307,In_2376);
nor U774 (N_774,In_2131,In_1749);
nand U775 (N_775,N_471,In_1844);
or U776 (N_776,In_575,In_1330);
and U777 (N_777,In_2450,In_942);
or U778 (N_778,In_255,N_136);
xnor U779 (N_779,In_1084,In_280);
or U780 (N_780,In_283,In_729);
xnor U781 (N_781,In_1538,In_1620);
nor U782 (N_782,In_1838,In_2308);
or U783 (N_783,N_375,N_426);
or U784 (N_784,In_2268,In_2108);
nand U785 (N_785,In_369,In_2193);
and U786 (N_786,In_1438,In_611);
nor U787 (N_787,In_2467,In_350);
and U788 (N_788,In_1718,In_2039);
xor U789 (N_789,In_2197,In_2475);
xnor U790 (N_790,N_170,N_253);
and U791 (N_791,N_71,In_296);
and U792 (N_792,N_327,In_236);
nand U793 (N_793,N_119,In_92);
or U794 (N_794,In_561,In_16);
or U795 (N_795,N_255,In_2093);
or U796 (N_796,In_1963,In_1717);
nor U797 (N_797,N_235,N_489);
xnor U798 (N_798,In_1692,In_471);
nand U799 (N_799,In_1945,N_200);
nor U800 (N_800,N_58,In_263);
nand U801 (N_801,In_1231,In_631);
nor U802 (N_802,In_1363,In_1941);
nor U803 (N_803,N_456,In_1518);
xnor U804 (N_804,N_23,In_1499);
nor U805 (N_805,In_1566,In_2408);
xnor U806 (N_806,N_453,N_294);
nor U807 (N_807,N_448,In_1618);
and U808 (N_808,In_146,N_31);
and U809 (N_809,In_399,In_1722);
nand U810 (N_810,In_537,In_1895);
nor U811 (N_811,In_1121,In_1517);
or U812 (N_812,In_35,N_29);
nor U813 (N_813,In_380,In_1156);
nand U814 (N_814,In_623,In_1090);
nor U815 (N_815,In_2364,In_734);
xor U816 (N_816,In_378,In_267);
xnor U817 (N_817,In_396,In_591);
nor U818 (N_818,In_1490,N_169);
or U819 (N_819,In_1710,In_1677);
nand U820 (N_820,In_539,In_225);
nor U821 (N_821,N_98,In_1398);
nor U822 (N_822,N_102,In_2133);
and U823 (N_823,In_2389,In_2099);
or U824 (N_824,N_42,In_457);
nand U825 (N_825,In_1022,In_738);
nor U826 (N_826,In_1638,In_2382);
or U827 (N_827,In_1555,In_1308);
nand U828 (N_828,N_333,In_1768);
or U829 (N_829,In_167,In_888);
xor U830 (N_830,In_769,In_1921);
and U831 (N_831,In_1748,In_345);
nand U832 (N_832,N_198,In_401);
or U833 (N_833,In_1982,In_375);
and U834 (N_834,In_650,N_334);
nand U835 (N_835,In_2461,In_2434);
or U836 (N_836,In_1077,In_969);
nand U837 (N_837,In_1426,In_1849);
or U838 (N_838,In_1793,In_2455);
or U839 (N_839,In_601,In_1339);
and U840 (N_840,N_412,In_740);
nor U841 (N_841,N_271,In_852);
nor U842 (N_842,In_224,In_231);
xnor U843 (N_843,In_2134,N_132);
or U844 (N_844,In_1542,In_1925);
and U845 (N_845,In_1533,In_1673);
nor U846 (N_846,N_171,In_2173);
nor U847 (N_847,In_1792,In_352);
or U848 (N_848,N_368,In_1949);
nor U849 (N_849,N_446,In_1443);
xnor U850 (N_850,In_2440,In_2064);
or U851 (N_851,In_2374,In_1347);
nand U852 (N_852,In_955,In_1440);
nor U853 (N_853,N_122,In_1018);
and U854 (N_854,In_1704,In_322);
nor U855 (N_855,In_135,N_303);
xor U856 (N_856,N_324,In_869);
and U857 (N_857,In_1983,In_1774);
and U858 (N_858,In_2332,In_1988);
and U859 (N_859,N_498,In_513);
or U860 (N_860,In_1794,N_275);
and U861 (N_861,N_157,In_239);
xor U862 (N_862,In_1827,N_192);
nand U863 (N_863,In_895,In_293);
or U864 (N_864,In_2429,N_145);
xor U865 (N_865,N_60,N_97);
and U866 (N_866,In_658,In_948);
nand U867 (N_867,In_830,N_263);
xor U868 (N_868,In_1164,N_49);
or U869 (N_869,N_311,In_34);
and U870 (N_870,In_116,In_2198);
or U871 (N_871,In_2118,In_1442);
nor U872 (N_872,In_18,In_593);
nor U873 (N_873,In_1763,In_58);
and U874 (N_874,In_383,In_1082);
nand U875 (N_875,N_335,In_1552);
and U876 (N_876,In_1986,In_705);
nand U877 (N_877,N_341,In_1817);
xnor U878 (N_878,N_434,In_766);
xnor U879 (N_879,In_607,In_782);
or U880 (N_880,N_162,In_542);
nor U881 (N_881,N_104,In_1648);
and U882 (N_882,In_1600,In_2026);
xor U883 (N_883,In_2182,In_2139);
xnor U884 (N_884,In_2333,N_146);
nand U885 (N_885,N_463,In_715);
xor U886 (N_886,In_1139,In_1810);
nand U887 (N_887,N_388,N_492);
xor U888 (N_888,In_1421,N_45);
or U889 (N_889,N_413,In_1549);
or U890 (N_890,N_50,N_16);
nand U891 (N_891,In_1033,In_2437);
nor U892 (N_892,In_111,N_79);
nor U893 (N_893,In_2267,In_1916);
and U894 (N_894,In_2028,In_990);
and U895 (N_895,In_2132,In_2172);
nand U896 (N_896,In_1424,In_435);
xor U897 (N_897,N_385,In_1445);
nand U898 (N_898,In_2412,N_141);
nand U899 (N_899,In_571,In_1003);
and U900 (N_900,In_1950,In_701);
nor U901 (N_901,In_1257,N_4);
nor U902 (N_902,In_1834,In_2061);
nor U903 (N_903,In_694,N_43);
nor U904 (N_904,In_1853,In_1966);
xor U905 (N_905,N_85,In_750);
nor U906 (N_906,N_74,In_655);
and U907 (N_907,In_915,In_859);
nand U908 (N_908,N_120,N_239);
xor U909 (N_909,In_160,N_174);
nor U910 (N_910,In_195,In_2036);
nand U911 (N_911,In_1975,In_876);
or U912 (N_912,In_784,N_397);
xnor U913 (N_913,N_6,In_389);
xnor U914 (N_914,In_275,In_1178);
and U915 (N_915,In_1608,In_599);
nand U916 (N_916,In_1913,N_209);
or U917 (N_917,N_369,In_1694);
or U918 (N_918,In_2046,In_2152);
and U919 (N_919,In_2050,In_1297);
nor U920 (N_920,In_829,In_817);
or U921 (N_921,In_1507,In_789);
xnor U922 (N_922,In_654,In_1681);
or U923 (N_923,In_1752,N_48);
nand U924 (N_924,In_171,In_1333);
or U925 (N_925,In_1891,In_163);
nor U926 (N_926,N_210,In_552);
and U927 (N_927,In_839,In_215);
nor U928 (N_928,In_1265,In_2355);
nor U929 (N_929,In_1230,N_166);
or U930 (N_930,In_465,In_1644);
nand U931 (N_931,In_290,In_918);
and U932 (N_932,N_212,In_1806);
nand U933 (N_933,In_492,In_1076);
nor U934 (N_934,N_159,In_1705);
and U935 (N_935,In_1874,In_1203);
nor U936 (N_936,In_1581,In_692);
nor U937 (N_937,In_775,In_1582);
xnor U938 (N_938,In_298,N_230);
nor U939 (N_939,In_351,In_1336);
nor U940 (N_940,N_490,N_205);
nand U941 (N_941,In_2415,In_1204);
or U942 (N_942,In_2114,In_1149);
nor U943 (N_943,In_59,N_78);
xnor U944 (N_944,N_128,In_2370);
and U945 (N_945,In_1109,In_1973);
nor U946 (N_946,In_318,N_378);
nor U947 (N_947,In_854,In_544);
xor U948 (N_948,In_192,In_1961);
or U949 (N_949,In_98,N_124);
nand U950 (N_950,In_1052,In_317);
or U951 (N_951,N_349,In_1829);
nor U952 (N_952,In_1726,In_2163);
nor U953 (N_953,N_243,In_1739);
and U954 (N_954,In_2313,In_679);
xnor U955 (N_955,In_291,In_1101);
nand U956 (N_956,In_2394,N_411);
or U957 (N_957,N_421,In_1248);
nand U958 (N_958,In_437,In_1043);
xnor U959 (N_959,N_319,In_1658);
and U960 (N_960,N_39,N_254);
xnor U961 (N_961,In_1034,In_1254);
and U962 (N_962,N_56,In_2368);
or U963 (N_963,In_519,In_276);
nand U964 (N_964,N_10,In_660);
and U965 (N_965,N_149,In_550);
nand U966 (N_966,N_75,In_847);
and U967 (N_967,N_22,In_49);
nand U968 (N_968,N_408,In_604);
nand U969 (N_969,In_1609,In_447);
and U970 (N_970,In_882,In_506);
nor U971 (N_971,In_1698,In_868);
or U972 (N_972,In_95,N_70);
nand U973 (N_973,In_545,In_1227);
nand U974 (N_974,In_1237,In_1847);
xor U975 (N_975,In_2184,In_671);
nand U976 (N_976,In_1972,In_1425);
nand U977 (N_977,N_152,In_125);
nand U978 (N_978,In_1803,N_95);
xor U979 (N_979,In_1878,In_808);
xor U980 (N_980,In_1540,In_511);
or U981 (N_981,In_169,In_1105);
nor U982 (N_982,In_1508,In_628);
and U983 (N_983,In_810,In_754);
nand U984 (N_984,N_231,In_1591);
xor U985 (N_985,In_2003,N_295);
xnor U986 (N_986,In_837,In_2104);
nand U987 (N_987,N_373,In_748);
nor U988 (N_988,N_409,In_1590);
nor U989 (N_989,In_635,N_258);
nor U990 (N_990,N_135,In_667);
and U991 (N_991,N_214,In_2240);
and U992 (N_992,In_2005,In_475);
nor U993 (N_993,In_120,In_1289);
nor U994 (N_994,In_2296,In_148);
xnor U995 (N_995,In_1437,In_2174);
or U996 (N_996,In_122,In_1998);
or U997 (N_997,N_247,In_1282);
nor U998 (N_998,In_1484,N_175);
nor U999 (N_999,N_88,N_462);
or U1000 (N_1000,In_2021,N_684);
nand U1001 (N_1001,In_1065,N_225);
nor U1002 (N_1002,In_1771,N_964);
xnor U1003 (N_1003,In_1073,N_165);
nand U1004 (N_1004,In_1532,N_173);
nand U1005 (N_1005,In_312,In_1647);
or U1006 (N_1006,N_51,In_901);
nor U1007 (N_1007,N_911,In_815);
and U1008 (N_1008,In_1759,In_1181);
nand U1009 (N_1009,N_667,In_2187);
and U1010 (N_1010,In_1274,In_494);
and U1011 (N_1011,N_878,N_885);
nand U1012 (N_1012,N_604,N_888);
xnor U1013 (N_1013,In_1463,In_1593);
nand U1014 (N_1014,N_429,In_1366);
nor U1015 (N_1015,N_927,In_1107);
nand U1016 (N_1016,In_2300,In_943);
nand U1017 (N_1017,In_201,In_2420);
nor U1018 (N_1018,N_437,N_504);
nand U1019 (N_1019,N_579,N_365);
nor U1020 (N_1020,In_495,In_19);
nor U1021 (N_1021,N_985,In_1689);
or U1022 (N_1022,N_537,N_129);
nand U1023 (N_1023,N_7,N_221);
nor U1024 (N_1024,In_1319,In_2221);
xor U1025 (N_1025,N_692,In_288);
nor U1026 (N_1026,N_548,In_856);
nor U1027 (N_1027,In_505,In_832);
or U1028 (N_1028,In_233,In_151);
nand U1029 (N_1029,N_112,In_1000);
xor U1030 (N_1030,N_0,In_299);
and U1031 (N_1031,In_1976,N_861);
or U1032 (N_1032,In_518,N_781);
or U1033 (N_1033,In_1769,N_808);
nand U1034 (N_1034,In_1831,N_918);
or U1035 (N_1035,N_519,N_843);
nand U1036 (N_1036,N_675,N_590);
nor U1037 (N_1037,N_794,In_187);
nand U1038 (N_1038,In_720,N_558);
nand U1039 (N_1039,In_1005,In_1800);
nor U1040 (N_1040,In_2126,In_1162);
xor U1041 (N_1041,In_2263,In_209);
and U1042 (N_1042,N_854,N_502);
nand U1043 (N_1043,N_841,N_668);
or U1044 (N_1044,In_1326,N_435);
xor U1045 (N_1045,In_2158,In_2080);
and U1046 (N_1046,In_2236,N_315);
and U1047 (N_1047,In_1707,In_1764);
xor U1048 (N_1048,N_839,In_339);
xor U1049 (N_1049,N_646,N_573);
nand U1050 (N_1050,N_735,In_2428);
or U1051 (N_1051,In_259,In_1063);
nand U1052 (N_1052,N_526,N_600);
xnor U1053 (N_1053,N_229,In_516);
nor U1054 (N_1054,In_1894,N_33);
and U1055 (N_1055,N_818,N_910);
nor U1056 (N_1056,In_1275,N_559);
nand U1057 (N_1057,N_228,N_578);
nand U1058 (N_1058,In_1733,In_1477);
xnor U1059 (N_1059,N_91,In_586);
and U1060 (N_1060,In_1035,In_2175);
nor U1061 (N_1061,N_391,N_356);
or U1062 (N_1062,N_586,In_1788);
nor U1063 (N_1063,N_110,N_977);
nor U1064 (N_1064,In_38,N_980);
nor U1065 (N_1065,In_1729,N_59);
nor U1066 (N_1066,In_665,N_287);
and U1067 (N_1067,N_115,In_1092);
nor U1068 (N_1068,In_602,In_347);
xor U1069 (N_1069,N_274,N_681);
nand U1070 (N_1070,In_119,N_522);
nor U1071 (N_1071,In_1563,N_840);
nand U1072 (N_1072,In_2377,In_185);
or U1073 (N_1073,N_147,N_218);
or U1074 (N_1074,N_176,In_1703);
nor U1075 (N_1075,In_2385,N_819);
nor U1076 (N_1076,In_1478,N_480);
nand U1077 (N_1077,In_336,N_851);
nor U1078 (N_1078,N_393,N_720);
or U1079 (N_1079,N_825,N_25);
nor U1080 (N_1080,N_967,In_726);
nor U1081 (N_1081,In_1789,N_433);
or U1082 (N_1082,N_134,N_499);
and U1083 (N_1083,In_1931,In_1494);
or U1084 (N_1084,N_40,In_2445);
or U1085 (N_1085,N_418,N_949);
nor U1086 (N_1086,N_727,N_19);
nor U1087 (N_1087,N_524,In_1273);
nor U1088 (N_1088,N_761,N_935);
nand U1089 (N_1089,In_191,In_923);
nand U1090 (N_1090,In_2327,N_625);
xor U1091 (N_1091,N_216,N_204);
or U1092 (N_1092,N_362,N_926);
nand U1093 (N_1093,In_998,In_2398);
nor U1094 (N_1094,N_717,N_680);
or U1095 (N_1095,N_778,In_1124);
and U1096 (N_1096,In_961,N_912);
nor U1097 (N_1097,N_706,In_2285);
nand U1098 (N_1098,N_493,N_399);
nor U1099 (N_1099,N_847,N_938);
or U1100 (N_1100,N_427,N_167);
nor U1101 (N_1101,N_756,N_922);
nand U1102 (N_1102,N_970,In_1129);
nand U1103 (N_1103,N_958,In_767);
xor U1104 (N_1104,N_1,In_1708);
or U1105 (N_1105,In_630,N_108);
or U1106 (N_1106,In_393,In_253);
and U1107 (N_1107,N_410,N_933);
nand U1108 (N_1108,In_1712,In_1305);
nor U1109 (N_1109,In_2115,In_522);
nand U1110 (N_1110,In_1026,In_486);
or U1111 (N_1111,N_865,N_487);
nor U1112 (N_1112,N_547,In_118);
and U1113 (N_1113,N_479,In_24);
and U1114 (N_1114,N_942,In_30);
nand U1115 (N_1115,In_624,In_765);
xor U1116 (N_1116,N_509,N_639);
nor U1117 (N_1117,In_1978,In_997);
nor U1118 (N_1118,In_2124,In_2116);
and U1119 (N_1119,In_1211,N_740);
nand U1120 (N_1120,N_921,N_266);
and U1121 (N_1121,In_2301,In_1859);
nor U1122 (N_1122,N_814,N_111);
nor U1123 (N_1123,In_1820,N_773);
nor U1124 (N_1124,In_1727,N_650);
xor U1125 (N_1125,N_308,In_2151);
xor U1126 (N_1126,In_1746,N_477);
and U1127 (N_1127,In_2417,N_826);
and U1128 (N_1128,N_81,N_571);
or U1129 (N_1129,In_965,N_505);
xor U1130 (N_1130,N_441,N_550);
and U1131 (N_1131,In_1314,N_989);
xnor U1132 (N_1132,N_64,N_821);
nor U1133 (N_1133,N_510,In_543);
nor U1134 (N_1134,N_987,In_82);
nor U1135 (N_1135,N_506,In_2024);
xnor U1136 (N_1136,In_1802,In_1171);
xor U1137 (N_1137,In_150,N_503);
or U1138 (N_1138,N_904,N_943);
nand U1139 (N_1139,In_1685,N_161);
nor U1140 (N_1140,N_440,N_853);
and U1141 (N_1141,N_466,N_265);
nand U1142 (N_1142,In_22,In_741);
nor U1143 (N_1143,N_486,N_541);
nor U1144 (N_1144,N_62,N_875);
nor U1145 (N_1145,N_884,In_1904);
or U1146 (N_1146,N_952,N_743);
or U1147 (N_1147,N_994,N_2);
or U1148 (N_1148,N_730,N_901);
nor U1149 (N_1149,N_978,N_734);
xnor U1150 (N_1150,In_2148,In_128);
xor U1151 (N_1151,N_609,N_154);
xnor U1152 (N_1152,N_139,In_1560);
nand U1153 (N_1153,In_1790,N_549);
xor U1154 (N_1154,N_199,In_1268);
xnor U1155 (N_1155,In_708,In_2199);
and U1156 (N_1156,In_2282,N_595);
and U1157 (N_1157,In_452,N_465);
xnor U1158 (N_1158,N_722,N_473);
or U1159 (N_1159,N_842,N_916);
xor U1160 (N_1160,N_118,In_311);
xor U1161 (N_1161,N_467,In_2143);
nor U1162 (N_1162,In_1881,In_686);
or U1163 (N_1163,N_713,N_770);
xnor U1164 (N_1164,In_42,In_1534);
and U1165 (N_1165,N_835,N_329);
xor U1166 (N_1166,N_371,N_494);
and U1167 (N_1167,N_67,In_1785);
nand U1168 (N_1168,N_917,N_774);
or U1169 (N_1169,In_391,N_953);
and U1170 (N_1170,In_1353,N_331);
nor U1171 (N_1171,In_594,In_2209);
or U1172 (N_1172,N_142,N_241);
nor U1173 (N_1173,In_566,In_2309);
or U1174 (N_1174,In_1485,In_1699);
and U1175 (N_1175,N_603,In_2130);
and U1176 (N_1176,In_2446,In_800);
nor U1177 (N_1177,N_937,N_696);
nor U1178 (N_1178,N_529,N_934);
or U1179 (N_1179,N_805,In_749);
or U1180 (N_1180,N_882,In_1742);
xnor U1181 (N_1181,N_662,In_845);
nor U1182 (N_1182,N_593,N_99);
and U1183 (N_1183,N_950,In_1048);
and U1184 (N_1184,In_2423,In_250);
or U1185 (N_1185,N_732,N_936);
or U1186 (N_1186,N_407,In_1316);
nor U1187 (N_1187,N_278,N_464);
xnor U1188 (N_1188,N_598,In_1144);
or U1189 (N_1189,N_742,In_1605);
nand U1190 (N_1190,N_903,In_1229);
nand U1191 (N_1191,In_1270,N_148);
or U1192 (N_1192,N_886,In_1613);
xnor U1193 (N_1193,In_394,In_1775);
or U1194 (N_1194,In_2356,N_830);
and U1195 (N_1195,In_2255,N_496);
xnor U1196 (N_1196,In_2334,N_21);
nand U1197 (N_1197,N_423,In_478);
and U1198 (N_1198,In_76,In_300);
nand U1199 (N_1199,In_476,In_254);
xnor U1200 (N_1200,In_1747,In_2054);
and U1201 (N_1201,N_828,In_653);
nor U1202 (N_1202,In_1606,N_133);
nand U1203 (N_1203,N_862,N_86);
nor U1204 (N_1204,N_807,N_849);
xnor U1205 (N_1205,N_645,N_915);
and U1206 (N_1206,In_2399,In_709);
xor U1207 (N_1207,In_1017,N_923);
xnor U1208 (N_1208,In_1651,In_454);
or U1209 (N_1209,N_871,In_2159);
nand U1210 (N_1210,In_147,N_272);
nand U1211 (N_1211,In_673,In_958);
nand U1212 (N_1212,N_992,In_2487);
and U1213 (N_1213,In_2262,N_749);
nand U1214 (N_1214,N_226,N_669);
or U1215 (N_1215,In_1038,N_364);
nand U1216 (N_1216,In_251,N_563);
and U1217 (N_1217,In_2095,In_1903);
and U1218 (N_1218,N_109,N_309);
and U1219 (N_1219,N_867,N_686);
nand U1220 (N_1220,N_451,In_436);
xor U1221 (N_1221,In_228,In_589);
nand U1222 (N_1222,In_1360,N_659);
and U1223 (N_1223,N_974,N_83);
and U1224 (N_1224,N_567,In_157);
and U1225 (N_1225,N_673,In_1672);
or U1226 (N_1226,N_795,N_786);
or U1227 (N_1227,N_850,In_2147);
nor U1228 (N_1228,N_976,In_41);
nor U1229 (N_1229,In_2493,In_2307);
nor U1230 (N_1230,N_664,N_540);
xor U1231 (N_1231,N_531,In_2371);
nand U1232 (N_1232,In_1719,In_1202);
nor U1233 (N_1233,N_188,In_1715);
or U1234 (N_1234,In_2378,In_1577);
xnor U1235 (N_1235,In_484,N_704);
xnor U1236 (N_1236,In_1586,In_433);
nand U1237 (N_1237,N_340,In_139);
xnor U1238 (N_1238,N_299,In_2485);
nor U1239 (N_1239,In_2403,In_826);
and U1240 (N_1240,In_381,N_940);
or U1241 (N_1241,In_1321,N_234);
xnor U1242 (N_1242,In_2283,In_1371);
and U1243 (N_1243,In_1332,N_852);
or U1244 (N_1244,N_249,In_2314);
xnor U1245 (N_1245,N_712,In_480);
nor U1246 (N_1246,N_705,N_597);
xnor U1247 (N_1247,N_769,In_1867);
xnor U1248 (N_1248,N_337,In_503);
nor U1249 (N_1249,N_417,In_2166);
nor U1250 (N_1250,N_602,In_2057);
xnor U1251 (N_1251,In_1350,In_713);
nand U1252 (N_1252,N_898,N_244);
nor U1253 (N_1253,In_1068,N_594);
xnor U1254 (N_1254,N_626,N_836);
nand U1255 (N_1255,In_2138,N_820);
and U1256 (N_1256,In_1639,In_159);
xnor U1257 (N_1257,In_65,In_986);
nand U1258 (N_1258,N_195,N_553);
and U1259 (N_1259,In_1464,In_2106);
and U1260 (N_1260,In_1123,In_794);
and U1261 (N_1261,In_1331,N_753);
nor U1262 (N_1262,In_1138,N_401);
and U1263 (N_1263,N_458,N_283);
xor U1264 (N_1264,N_80,N_389);
or U1265 (N_1265,N_719,N_638);
nand U1266 (N_1266,In_1992,N_996);
and U1267 (N_1267,N_988,In_302);
nand U1268 (N_1268,In_2384,N_568);
nand U1269 (N_1269,In_2281,N_376);
xnor U1270 (N_1270,N_738,N_491);
xnor U1271 (N_1271,N_792,In_368);
or U1272 (N_1272,In_443,In_1131);
nor U1273 (N_1273,N_762,N_472);
nand U1274 (N_1274,In_1828,N_708);
or U1275 (N_1275,In_184,In_434);
or U1276 (N_1276,N_975,In_53);
nand U1277 (N_1277,In_459,In_1454);
nor U1278 (N_1278,In_221,In_1799);
nand U1279 (N_1279,In_1622,N_585);
nor U1280 (N_1280,N_766,In_1506);
xnor U1281 (N_1281,In_2001,N_584);
or U1282 (N_1282,N_846,N_232);
and U1283 (N_1283,N_801,N_811);
xnor U1284 (N_1284,N_606,N_824);
xor U1285 (N_1285,In_1960,In_2486);
nand U1286 (N_1286,In_245,N_859);
nand U1287 (N_1287,N_474,In_1046);
or U1288 (N_1288,In_886,N_737);
and U1289 (N_1289,In_2482,In_482);
nand U1290 (N_1290,In_776,N_605);
and U1291 (N_1291,In_238,In_1057);
and U1292 (N_1292,N_893,In_937);
or U1293 (N_1293,In_1948,N_13);
nand U1294 (N_1294,N_37,N_587);
or U1295 (N_1295,N_156,In_1568);
and U1296 (N_1296,In_1731,In_1877);
and U1297 (N_1297,N_944,In_1741);
nand U1298 (N_1298,N_301,N_312);
nor U1299 (N_1299,N_666,N_791);
xor U1300 (N_1300,In_848,In_1253);
nor U1301 (N_1301,In_330,N_344);
xor U1302 (N_1302,N_941,N_665);
and U1303 (N_1303,N_137,In_1355);
or U1304 (N_1304,In_63,N_36);
nor U1305 (N_1305,In_1614,In_1228);
xnor U1306 (N_1306,In_1657,N_640);
xor U1307 (N_1307,In_417,N_711);
nor U1308 (N_1308,In_114,In_445);
xnor U1309 (N_1309,N_582,N_823);
and U1310 (N_1310,In_2278,In_91);
and U1311 (N_1311,In_1971,N_92);
and U1312 (N_1312,N_802,In_722);
nor U1313 (N_1313,N_125,In_656);
nor U1314 (N_1314,N_679,In_1579);
xnor U1315 (N_1315,In_1293,N_929);
nand U1316 (N_1316,N_355,In_2290);
or U1317 (N_1317,In_2015,N_561);
and U1318 (N_1318,N_386,In_357);
xor U1319 (N_1319,In_1047,In_587);
xnor U1320 (N_1320,N_222,In_2010);
nor U1321 (N_1321,In_1754,In_252);
nor U1322 (N_1322,In_988,In_1309);
xnor U1323 (N_1323,In_2065,In_2177);
or U1324 (N_1324,In_824,N_747);
xor U1325 (N_1325,In_133,N_876);
xnor U1326 (N_1326,In_1037,N_951);
and U1327 (N_1327,In_884,N_532);
or U1328 (N_1328,In_474,In_2405);
nand U1329 (N_1329,In_324,In_2253);
xnor U1330 (N_1330,N_18,N_784);
and U1331 (N_1331,N_252,In_414);
nand U1332 (N_1332,In_1102,In_1879);
nor U1333 (N_1333,In_1787,In_922);
nor U1334 (N_1334,N_390,In_1599);
xnor U1335 (N_1335,N_909,N_288);
nand U1336 (N_1336,N_863,N_671);
xnor U1337 (N_1337,In_1740,In_1359);
or U1338 (N_1338,In_889,N_624);
and U1339 (N_1339,In_534,N_153);
or U1340 (N_1340,In_212,In_364);
or U1341 (N_1341,In_2397,N_381);
xnor U1342 (N_1342,In_735,In_1459);
nor U1343 (N_1343,N_963,In_2167);
xor U1344 (N_1344,N_183,In_605);
nor U1345 (N_1345,N_443,In_338);
nor U1346 (N_1346,In_2350,N_694);
nor U1347 (N_1347,N_748,In_1734);
or U1348 (N_1348,In_960,N_848);
or U1349 (N_1349,N_858,N_990);
and U1350 (N_1350,N_751,N_972);
or U1351 (N_1351,In_1087,In_2298);
nor U1352 (N_1352,In_2109,N_661);
nand U1353 (N_1353,In_2322,In_1475);
xor U1354 (N_1354,In_382,N_518);
nand U1355 (N_1355,In_2401,In_365);
and U1356 (N_1356,In_2460,In_241);
nor U1357 (N_1357,N_632,N_688);
or U1358 (N_1358,In_1150,In_639);
xnor U1359 (N_1359,In_633,N_46);
xnor U1360 (N_1360,In_1662,N_599);
nand U1361 (N_1361,In_1468,N_262);
xnor U1362 (N_1362,N_971,In_329);
nand U1363 (N_1363,N_930,N_806);
or U1364 (N_1364,N_27,In_388);
nand U1365 (N_1365,In_1462,N_642);
nand U1366 (N_1366,In_971,In_1919);
and U1367 (N_1367,In_710,In_1176);
nand U1368 (N_1368,N_880,N_764);
nand U1369 (N_1369,In_1932,In_11);
nand U1370 (N_1370,N_767,N_577);
xnor U1371 (N_1371,In_712,N_631);
nand U1372 (N_1372,N_752,In_1693);
nor U1373 (N_1373,In_1182,In_353);
or U1374 (N_1374,N_869,N_306);
nor U1375 (N_1375,In_1320,In_132);
and U1376 (N_1376,In_202,N_797);
nand U1377 (N_1377,In_113,N_860);
and U1378 (N_1378,In_541,N_530);
nor U1379 (N_1379,In_1900,N_701);
xor U1380 (N_1380,In_1537,N_523);
and U1381 (N_1381,N_960,N_768);
xor U1382 (N_1382,N_783,In_1345);
nand U1383 (N_1383,N_24,N_457);
or U1384 (N_1384,In_2458,N_197);
and U1385 (N_1385,In_595,N_576);
and U1386 (N_1386,In_216,N_956);
nor U1387 (N_1387,N_635,In_2249);
and U1388 (N_1388,In_69,In_140);
or U1389 (N_1389,N_651,N_114);
or U1390 (N_1390,In_423,N_360);
nor U1391 (N_1391,N_887,In_1125);
nand U1392 (N_1392,In_1205,In_1189);
and U1393 (N_1393,N_47,N_630);
and U1394 (N_1394,N_614,N_202);
or U1395 (N_1395,In_1851,N_322);
nor U1396 (N_1396,In_172,In_1857);
nor U1397 (N_1397,In_408,N_517);
or U1398 (N_1398,N_592,In_1888);
or U1399 (N_1399,In_1737,N_20);
nor U1400 (N_1400,N_765,In_348);
or U1401 (N_1401,N_450,In_1151);
xnor U1402 (N_1402,In_946,N_261);
and U1403 (N_1403,In_1645,In_1511);
xor U1404 (N_1404,N_321,N_866);
nand U1405 (N_1405,N_731,In_343);
xor U1406 (N_1406,N_703,In_934);
nor U1407 (N_1407,N_803,N_812);
nor U1408 (N_1408,In_110,In_1260);
xor U1409 (N_1409,N_892,In_62);
xor U1410 (N_1410,N_914,N_900);
or U1411 (N_1411,N_182,N_924);
nor U1412 (N_1412,In_1935,In_1924);
or U1413 (N_1413,In_1482,In_1387);
nor U1414 (N_1414,N_347,N_527);
xor U1415 (N_1415,In_1659,In_84);
nand U1416 (N_1416,In_101,N_618);
and U1417 (N_1417,In_727,In_386);
xor U1418 (N_1418,In_2189,N_121);
nor U1419 (N_1419,N_415,In_104);
nor U1420 (N_1420,In_1187,N_682);
nor U1421 (N_1421,N_838,N_920);
nand U1422 (N_1422,N_760,In_828);
nand U1423 (N_1423,N_436,N_982);
nand U1424 (N_1424,N_588,N_895);
nor U1425 (N_1425,In_162,In_1154);
nand U1426 (N_1426,In_1652,N_248);
nand U1427 (N_1427,N_583,In_2097);
xnor U1428 (N_1428,In_1226,N_403);
and U1429 (N_1429,N_220,In_548);
xnor U1430 (N_1430,N_520,In_2372);
xor U1431 (N_1431,N_789,N_481);
nand U1432 (N_1432,N_350,N_804);
or U1433 (N_1433,N_961,In_1011);
and U1434 (N_1434,In_1541,In_1720);
or U1435 (N_1435,In_778,N_469);
nor U1436 (N_1436,N_107,In_2246);
xnor U1437 (N_1437,In_1406,In_1377);
nand U1438 (N_1438,N_965,N_181);
xnor U1439 (N_1439,N_833,N_627);
nor U1440 (N_1440,N_931,In_733);
nor U1441 (N_1441,N_314,In_1551);
nand U1442 (N_1442,In_2400,N_44);
nor U1443 (N_1443,In_1843,N_945);
and U1444 (N_1444,In_1920,In_677);
and U1445 (N_1445,N_906,N_674);
and U1446 (N_1446,N_744,N_361);
and U1447 (N_1447,N_454,In_2127);
and U1448 (N_1448,In_2146,N_739);
or U1449 (N_1449,In_606,In_1051);
or U1450 (N_1450,In_521,In_1474);
xnor U1451 (N_1451,In_2375,In_1700);
and U1452 (N_1452,N_827,In_1027);
and U1453 (N_1453,N_581,In_206);
and U1454 (N_1454,In_1910,N_370);
or U1455 (N_1455,N_103,In_464);
xnor U1456 (N_1456,N_683,In_3);
nand U1457 (N_1457,In_1603,In_2241);
and U1458 (N_1458,In_1206,In_1324);
and U1459 (N_1459,N_172,N_889);
and U1460 (N_1460,In_2101,N_796);
xor U1461 (N_1461,In_1536,N_151);
nor U1462 (N_1462,N_721,N_637);
and U1463 (N_1463,In_1732,In_235);
xnor U1464 (N_1464,In_466,In_496);
and U1465 (N_1465,N_318,N_293);
nor U1466 (N_1466,In_2102,N_723);
and U1467 (N_1467,N_733,In_2012);
or U1468 (N_1468,In_2483,In_2052);
nor U1469 (N_1469,In_638,N_163);
or U1470 (N_1470,N_395,In_406);
xor U1471 (N_1471,In_490,In_850);
and U1472 (N_1472,N_623,N_829);
or U1473 (N_1473,In_1152,N_785);
nor U1474 (N_1474,N_725,N_580);
or U1475 (N_1475,N_832,In_2462);
nand U1476 (N_1476,In_1912,In_2190);
and U1477 (N_1477,In_940,In_1513);
or U1478 (N_1478,In_1642,In_1735);
nor U1479 (N_1479,In_363,N_905);
nand U1480 (N_1480,N_268,N_844);
nand U1481 (N_1481,In_493,N_556);
or U1482 (N_1482,N_822,In_2295);
nor U1483 (N_1483,In_805,N_621);
nand U1484 (N_1484,N_709,In_504);
nand U1485 (N_1485,N_691,N_955);
nor U1486 (N_1486,In_207,N_873);
or U1487 (N_1487,In_204,N_554);
nand U1488 (N_1488,In_456,N_336);
xnor U1489 (N_1489,In_642,In_526);
nor U1490 (N_1490,In_2297,In_2029);
or U1491 (N_1491,N_995,N_755);
xnor U1492 (N_1492,N_570,N_856);
and U1493 (N_1493,N_714,In_2492);
nor U1494 (N_1494,In_2324,In_1870);
xnor U1495 (N_1495,In_1882,N_658);
or U1496 (N_1496,N_72,N_816);
xor U1497 (N_1497,N_695,In_1111);
and U1498 (N_1498,In_1106,In_12);
and U1499 (N_1499,N_908,In_2192);
or U1500 (N_1500,N_1094,N_1317);
xnor U1501 (N_1501,N_1438,N_1058);
or U1502 (N_1502,In_1997,N_1430);
or U1503 (N_1503,N_1279,N_1377);
or U1504 (N_1504,N_1161,N_928);
xnor U1505 (N_1505,In_771,In_2276);
xor U1506 (N_1506,N_1335,N_831);
nor U1507 (N_1507,N_729,N_754);
or U1508 (N_1508,N_962,N_1310);
and U1509 (N_1509,N_566,N_3);
or U1510 (N_1510,N_1088,N_1056);
or U1511 (N_1511,In_2031,N_1307);
or U1512 (N_1512,In_1153,N_1116);
or U1513 (N_1513,N_242,N_736);
nor U1514 (N_1514,N_1378,N_622);
and U1515 (N_1515,In_2306,N_993);
or U1516 (N_1516,N_1270,N_1469);
nor U1517 (N_1517,N_678,N_1403);
and U1518 (N_1518,In_1161,In_1814);
nand U1519 (N_1519,N_1142,N_1224);
nand U1520 (N_1520,In_626,In_1597);
and U1521 (N_1521,N_1240,N_1391);
nor U1522 (N_1522,N_1290,N_1209);
and U1523 (N_1523,In_1091,N_534);
nand U1524 (N_1524,N_793,N_113);
and U1525 (N_1525,N_1259,N_302);
nand U1526 (N_1526,In_932,N_607);
nor U1527 (N_1527,In_2489,N_1212);
and U1528 (N_1528,In_25,N_1086);
or U1529 (N_1529,N_1480,In_1239);
nor U1530 (N_1530,N_1376,N_1481);
nor U1531 (N_1531,N_1364,N_428);
nor U1532 (N_1532,N_1028,N_1351);
and U1533 (N_1533,N_919,N_1268);
or U1534 (N_1534,In_262,N_1462);
and U1535 (N_1535,N_1045,N_1172);
nor U1536 (N_1536,N_1258,In_418);
or U1537 (N_1537,N_305,N_574);
nor U1538 (N_1538,In_349,In_893);
or U1539 (N_1539,N_1429,N_946);
nor U1540 (N_1540,N_1341,N_1052);
nand U1541 (N_1541,N_1302,N_1138);
xor U1542 (N_1542,In_473,N_1402);
nor U1543 (N_1543,N_710,In_2357);
or U1544 (N_1544,N_1195,N_117);
xor U1545 (N_1545,N_1032,In_1892);
xor U1546 (N_1546,N_1387,N_34);
and U1547 (N_1547,N_1472,In_2030);
and U1548 (N_1548,In_2245,N_1320);
and U1549 (N_1549,In_1811,N_1063);
xnor U1550 (N_1550,N_1074,N_219);
or U1551 (N_1551,In_178,N_1308);
nand U1552 (N_1552,N_1175,In_647);
nand U1553 (N_1553,N_984,In_1408);
or U1554 (N_1554,N_758,N_1038);
nand U1555 (N_1555,In_1170,In_1145);
nor U1556 (N_1556,N_1078,N_677);
nor U1557 (N_1557,N_1339,N_968);
and U1558 (N_1558,N_179,N_1476);
xnor U1559 (N_1559,In_681,N_1273);
xnor U1560 (N_1560,N_707,N_1368);
nand U1561 (N_1561,N_1414,N_240);
nor U1562 (N_1562,N_1228,N_1083);
and U1563 (N_1563,In_570,N_777);
nor U1564 (N_1564,N_1277,N_1183);
nor U1565 (N_1565,N_1379,N_1437);
and U1566 (N_1566,N_1098,N_1075);
nor U1567 (N_1567,N_1122,N_1408);
and U1568 (N_1568,In_877,N_1455);
or U1569 (N_1569,N_1295,N_1050);
nor U1570 (N_1570,N_1162,N_1047);
nor U1571 (N_1571,N_1392,N_907);
nand U1572 (N_1572,In_446,N_420);
nor U1573 (N_1573,N_1176,N_1332);
nor U1574 (N_1574,In_407,N_431);
or U1575 (N_1575,N_533,In_1994);
nor U1576 (N_1576,N_672,N_1151);
xor U1577 (N_1577,N_1108,N_986);
nand U1578 (N_1578,N_1360,N_636);
xnor U1579 (N_1579,N_1060,In_524);
xor U1580 (N_1580,N_1386,N_1309);
nor U1581 (N_1581,N_1238,In_896);
nand U1582 (N_1582,N_655,In_843);
and U1583 (N_1583,In_2388,N_1323);
nand U1584 (N_1584,N_817,In_762);
nor U1585 (N_1585,N_1054,N_1287);
nand U1586 (N_1586,In_1795,N_1447);
nand U1587 (N_1587,N_1338,In_779);
xor U1588 (N_1588,In_755,N_1282);
nand U1589 (N_1589,N_775,N_470);
nor U1590 (N_1590,N_1483,N_641);
or U1591 (N_1591,N_562,N_1485);
nand U1592 (N_1592,N_1325,N_1255);
and U1593 (N_1593,N_277,N_1367);
and U1594 (N_1594,N_591,N_511);
or U1595 (N_1595,In_358,N_779);
nor U1596 (N_1596,N_1226,N_1460);
xor U1597 (N_1597,N_872,In_400);
or U1598 (N_1598,N_1157,In_851);
nand U1599 (N_1599,N_619,N_12);
nand U1600 (N_1600,N_913,In_2053);
nand U1601 (N_1601,N_1201,N_1445);
nor U1602 (N_1602,N_1107,N_1486);
or U1603 (N_1603,In_1066,N_1187);
xnor U1604 (N_1604,N_1291,N_617);
nor U1605 (N_1605,N_790,In_2427);
and U1606 (N_1606,N_1092,In_1524);
xnor U1607 (N_1607,N_1372,N_1019);
xor U1608 (N_1608,In_468,N_90);
and U1609 (N_1609,N_1362,N_1284);
or U1610 (N_1610,N_1231,N_782);
xor U1611 (N_1611,N_93,In_1680);
nand U1612 (N_1612,In_295,N_544);
xnor U1613 (N_1613,In_1915,N_1200);
xnor U1614 (N_1614,In_2222,N_1340);
xnor U1615 (N_1615,N_1356,N_698);
nor U1616 (N_1616,N_894,In_902);
or U1617 (N_1617,N_1070,N_1105);
nor U1618 (N_1618,N_414,N_1329);
and U1619 (N_1619,N_628,N_1036);
nor U1620 (N_1620,N_1464,N_1085);
and U1621 (N_1621,N_1327,N_1271);
or U1622 (N_1622,N_1363,N_1384);
nor U1623 (N_1623,In_2425,N_1194);
and U1624 (N_1624,N_250,N_1444);
or U1625 (N_1625,N_1048,N_991);
and U1626 (N_1626,N_676,N_983);
or U1627 (N_1627,N_1192,N_1448);
and U1628 (N_1628,N_1266,In_528);
nand U1629 (N_1629,In_1195,N_1010);
or U1630 (N_1630,In_821,N_959);
and U1631 (N_1631,N_1191,N_1352);
nor U1632 (N_1632,N_601,In_413);
and U1633 (N_1633,N_1267,N_1269);
or U1634 (N_1634,N_1081,In_1927);
and U1635 (N_1635,In_580,N_1043);
and U1636 (N_1636,N_615,N_1189);
and U1637 (N_1637,N_1446,In_1112);
and U1638 (N_1638,N_1229,N_246);
or U1639 (N_1639,In_637,In_840);
nor U1640 (N_1640,N_1237,N_352);
and U1641 (N_1641,N_1262,N_536);
nand U1642 (N_1642,N_1319,In_1755);
nand U1643 (N_1643,N_1416,N_1102);
xor U1644 (N_1644,In_1856,N_1206);
nand U1645 (N_1645,N_1205,N_1350);
nor U1646 (N_1646,N_1230,N_1173);
or U1647 (N_1647,N_1002,N_687);
xor U1648 (N_1648,N_1426,N_73);
xor U1649 (N_1649,N_1440,N_1158);
nor U1650 (N_1650,In_691,In_1298);
nor U1651 (N_1651,N_1202,N_647);
nor U1652 (N_1652,N_1423,N_1245);
nand U1653 (N_1653,In_1780,In_1186);
nand U1654 (N_1654,In_2433,N_1133);
nand U1655 (N_1655,N_981,N_870);
or U1656 (N_1656,N_1140,N_699);
nand U1657 (N_1657,N_1396,In_385);
or U1658 (N_1658,N_1400,N_14);
and U1659 (N_1659,N_38,N_1153);
nor U1660 (N_1660,N_69,N_1404);
and U1661 (N_1661,N_1280,N_1039);
xnor U1662 (N_1662,N_750,N_1257);
xnor U1663 (N_1663,N_279,N_1049);
xor U1664 (N_1664,N_1385,In_996);
xor U1665 (N_1665,N_1111,N_1288);
nand U1666 (N_1666,N_763,N_1236);
nor U1667 (N_1667,N_1170,N_1457);
or U1668 (N_1668,N_1190,N_874);
nor U1669 (N_1669,In_1848,In_297);
nand U1670 (N_1670,N_1064,N_1196);
and U1671 (N_1671,N_834,In_573);
xor U1672 (N_1672,N_663,N_1355);
xnor U1673 (N_1673,N_1215,N_1473);
xor U1674 (N_1674,N_1470,N_1082);
nand U1675 (N_1675,N_1233,N_1024);
nor U1676 (N_1676,N_1040,N_1235);
nand U1677 (N_1677,N_186,N_514);
nand U1678 (N_1678,N_660,In_2265);
or U1679 (N_1679,N_1421,N_1496);
xnor U1680 (N_1680,N_400,N_1097);
nor U1681 (N_1681,N_1459,N_634);
xnor U1682 (N_1682,N_1366,In_1650);
nor U1683 (N_1683,N_1110,In_1547);
xor U1684 (N_1684,N_1346,In_1385);
or U1685 (N_1685,In_2180,In_2456);
nor U1686 (N_1686,In_1514,In_2013);
nor U1687 (N_1687,N_130,N_1297);
xor U1688 (N_1688,N_1337,N_932);
and U1689 (N_1689,N_746,N_1020);
nor U1690 (N_1690,N_406,In_1578);
nand U1691 (N_1691,N_1358,N_759);
or U1692 (N_1692,In_1108,N_1390);
and U1693 (N_1693,N_1180,In_1504);
nor U1694 (N_1694,N_101,N_575);
or U1695 (N_1695,In_131,N_1080);
nand U1696 (N_1696,N_1204,In_1876);
nor U1697 (N_1697,N_1300,In_2083);
or U1698 (N_1698,N_1482,N_259);
nand U1699 (N_1699,N_320,In_1781);
nor U1700 (N_1700,N_1061,N_300);
nor U1701 (N_1701,N_1033,N_1221);
nor U1702 (N_1702,In_1565,N_1005);
xor U1703 (N_1703,N_620,N_1285);
xnor U1704 (N_1704,N_1458,In_795);
or U1705 (N_1705,In_1328,N_1071);
nor U1706 (N_1706,N_1318,N_1411);
and U1707 (N_1707,In_6,N_189);
nor U1708 (N_1708,N_656,In_1479);
xnor U1709 (N_1709,In_1666,N_359);
or U1710 (N_1710,N_1023,In_517);
nor U1711 (N_1711,N_1292,N_1431);
nand U1712 (N_1712,In_103,N_1463);
xor U1713 (N_1713,In_1114,N_416);
xor U1714 (N_1714,N_652,N_1330);
nor U1715 (N_1715,N_223,N_1304);
nand U1716 (N_1716,N_741,N_1249);
nor U1717 (N_1717,N_689,N_1027);
xnor U1718 (N_1718,N_326,N_697);
and U1719 (N_1719,N_1399,In_536);
and U1720 (N_1720,N_1106,N_864);
xnor U1721 (N_1721,N_1001,N_542);
xnor U1722 (N_1722,N_515,N_1178);
nand U1723 (N_1723,N_1349,N_68);
nand U1724 (N_1724,N_724,In_1040);
nor U1725 (N_1725,In_240,In_1143);
xnor U1726 (N_1726,N_979,N_1479);
xor U1727 (N_1727,In_1104,In_176);
or U1728 (N_1728,N_1492,N_459);
nor U1729 (N_1729,N_1119,N_1344);
or U1730 (N_1730,N_1099,N_1156);
nand U1731 (N_1731,In_1325,N_1003);
or U1732 (N_1732,In_931,N_969);
nor U1733 (N_1733,N_1150,N_799);
and U1734 (N_1734,N_500,N_815);
xnor U1735 (N_1735,N_1053,N_1418);
nand U1736 (N_1736,In_777,N_1031);
or U1737 (N_1737,N_1381,N_1343);
or U1738 (N_1738,N_1326,N_144);
nor U1739 (N_1739,N_1076,N_1345);
nand U1740 (N_1740,N_948,In_328);
and U1741 (N_1741,N_1454,In_717);
and U1742 (N_1742,N_1306,N_1383);
nor U1743 (N_1743,N_328,N_693);
or U1744 (N_1744,N_1186,N_1051);
or U1745 (N_1745,In_1601,N_1293);
or U1746 (N_1746,In_1985,N_954);
or U1747 (N_1747,N_1316,N_1419);
nor U1748 (N_1748,N_1129,N_1025);
xnor U1749 (N_1749,In_1832,In_669);
xnor U1750 (N_1750,In_1122,N_1424);
or U1751 (N_1751,N_30,N_1298);
and U1752 (N_1752,N_788,N_546);
xor U1753 (N_1753,In_910,In_244);
xnor U1754 (N_1754,In_2178,N_1167);
nand U1755 (N_1755,In_2393,N_1322);
or U1756 (N_1756,N_1365,In_935);
or U1757 (N_1757,N_643,N_1289);
nand U1758 (N_1758,In_2310,N_1185);
or U1759 (N_1759,N_1132,N_1008);
or U1760 (N_1760,In_1846,In_1860);
nand U1761 (N_1761,N_1114,In_554);
xor U1762 (N_1762,N_1207,In_1868);
nand U1763 (N_1763,In_1630,N_1118);
nand U1764 (N_1764,N_387,N_1435);
nor U1765 (N_1765,N_1220,N_96);
nor U1766 (N_1766,N_1250,N_702);
nor U1767 (N_1767,N_896,N_1135);
nand U1768 (N_1768,In_574,In_1869);
and U1769 (N_1769,In_1374,In_1263);
and U1770 (N_1770,N_1227,N_508);
or U1771 (N_1771,N_425,N_1466);
or U1772 (N_1772,N_1046,In_2380);
xor U1773 (N_1773,In_158,N_1370);
nor U1774 (N_1774,N_1272,In_629);
or U1775 (N_1775,N_1296,In_2153);
nand U1776 (N_1776,N_555,N_1144);
and U1777 (N_1777,N_1371,In_1042);
nand U1778 (N_1778,In_440,N_1188);
and U1779 (N_1779,N_1498,In_924);
or U1780 (N_1780,N_564,N_897);
xor U1781 (N_1781,N_1016,N_507);
or U1782 (N_1782,N_1354,N_1055);
xor U1783 (N_1783,N_1000,In_1259);
and U1784 (N_1784,N_1145,In_1621);
nand U1785 (N_1785,In_1083,N_1013);
nand U1786 (N_1786,N_1405,N_1096);
nor U1787 (N_1787,N_1251,N_1217);
and U1788 (N_1788,N_1148,In_85);
nor U1789 (N_1789,N_66,N_1398);
nand U1790 (N_1790,In_742,In_174);
or U1791 (N_1791,N_1265,N_1422);
xor U1792 (N_1792,N_966,N_1120);
nand U1793 (N_1793,N_545,N_1127);
xor U1794 (N_1794,In_1198,N_612);
or U1795 (N_1795,N_1283,N_1100);
nor U1796 (N_1796,In_1250,In_1019);
or U1797 (N_1797,N_780,N_868);
and U1798 (N_1798,N_367,N_1274);
and U1799 (N_1799,In_1576,In_2363);
xnor U1800 (N_1800,N_998,N_1213);
and U1801 (N_1801,N_1174,N_1253);
and U1802 (N_1802,N_1037,In_972);
nand U1803 (N_1803,N_1168,N_1147);
xnor U1804 (N_1804,N_495,N_1260);
xor U1805 (N_1805,N_1305,N_1434);
or U1806 (N_1806,N_1465,N_685);
xnor U1807 (N_1807,N_1152,N_997);
and U1808 (N_1808,N_1079,N_837);
and U1809 (N_1809,In_346,In_819);
nand U1810 (N_1810,N_1324,In_1893);
and U1811 (N_1811,N_1246,In_1453);
or U1812 (N_1812,In_1476,N_1263);
and U1813 (N_1813,N_1030,In_1100);
nand U1814 (N_1814,N_1276,N_543);
nor U1815 (N_1815,N_891,N_257);
nor U1816 (N_1816,N_1208,N_648);
or U1817 (N_1817,N_1136,N_1369);
xnor U1818 (N_1818,N_1439,In_1808);
or U1819 (N_1819,In_2220,N_316);
nand U1820 (N_1820,N_1427,In_1280);
nand U1821 (N_1821,N_957,N_1184);
xor U1822 (N_1822,N_1415,In_610);
and U1823 (N_1823,N_1128,N_291);
xor U1824 (N_1824,N_1433,N_1216);
nor U1825 (N_1825,N_1166,N_1035);
nand U1826 (N_1826,N_84,N_1456);
xnor U1827 (N_1827,N_1177,In_2237);
xor U1828 (N_1828,N_1059,In_551);
and U1829 (N_1829,N_1139,N_1089);
and U1830 (N_1830,N_1225,N_1382);
or U1831 (N_1831,In_2213,N_611);
nor U1832 (N_1832,In_1990,N_521);
nand U1833 (N_1833,N_1453,In_546);
xnor U1834 (N_1834,In_814,N_1171);
xor U1835 (N_1835,In_855,N_57);
or U1836 (N_1836,N_1163,N_1478);
xor U1837 (N_1837,In_1348,N_1353);
xnor U1838 (N_1838,N_1395,N_1256);
xor U1839 (N_1839,N_557,N_1181);
xnor U1840 (N_1840,In_2441,N_608);
or U1841 (N_1841,In_2468,N_1471);
or U1842 (N_1842,In_2047,N_1487);
xnor U1843 (N_1843,In_1130,N_899);
and U1844 (N_1844,N_535,N_718);
nor U1845 (N_1845,N_1091,N_1252);
xnor U1846 (N_1846,N_1328,N_1160);
nand U1847 (N_1847,N_1203,N_1103);
and U1848 (N_1848,N_716,N_947);
and U1849 (N_1849,N_516,N_1169);
or U1850 (N_1850,In_75,N_513);
nor U1851 (N_1851,N_1413,N_1067);
nor U1852 (N_1852,N_1467,N_116);
or U1853 (N_1853,N_610,In_700);
and U1854 (N_1854,N_1477,N_1125);
nand U1855 (N_1855,N_1068,N_1495);
and U1856 (N_1856,In_46,In_2466);
xor U1857 (N_1857,N_1179,In_1683);
xor U1858 (N_1858,In_2181,N_1104);
xnor U1859 (N_1859,N_338,In_2078);
or U1860 (N_1860,In_783,N_613);
or U1861 (N_1861,N_1388,N_1211);
nor U1862 (N_1862,In_2086,N_1159);
nor U1863 (N_1863,N_1347,N_629);
nor U1864 (N_1864,N_798,N_1087);
nand U1865 (N_1865,N_1137,N_1057);
or U1866 (N_1866,N_1123,N_1021);
nand U1867 (N_1867,N_1155,N_881);
nand U1868 (N_1868,N_1018,N_1334);
or U1869 (N_1869,N_1109,N_289);
or U1870 (N_1870,N_1389,N_1248);
or U1871 (N_1871,N_1361,N_1130);
and U1872 (N_1872,N_1149,In_799);
or U1873 (N_1873,N_1494,N_1484);
nand U1874 (N_1874,N_1012,In_1872);
xnor U1875 (N_1875,N_1301,N_488);
nand U1876 (N_1876,N_177,In_442);
xor U1877 (N_1877,In_1089,N_539);
or U1878 (N_1878,N_292,In_1023);
nand U1879 (N_1879,In_1115,N_382);
and U1880 (N_1880,N_1449,N_1131);
nand U1881 (N_1881,N_654,N_1084);
nor U1882 (N_1882,N_1443,N_1214);
and U1883 (N_1883,N_1393,N_1493);
xnor U1884 (N_1884,N_809,N_1475);
and U1885 (N_1885,N_1281,In_367);
xnor U1886 (N_1886,N_1342,In_1247);
or U1887 (N_1887,N_1218,In_759);
xor U1888 (N_1888,N_1294,N_1006);
nand U1889 (N_1889,N_1165,N_1333);
or U1890 (N_1890,N_1314,N_1017);
xor U1891 (N_1891,N_1243,N_1101);
xor U1892 (N_1892,N_596,N_1254);
and U1893 (N_1893,In_183,N_1041);
or U1894 (N_1894,N_1072,N_1499);
nand U1895 (N_1895,N_1275,N_1374);
nand U1896 (N_1896,N_215,N_1394);
xor U1897 (N_1897,N_925,N_1113);
or U1898 (N_1898,In_1491,N_290);
nor U1899 (N_1899,N_1321,N_565);
or U1900 (N_1900,In_138,N_1117);
nand U1901 (N_1901,N_1199,In_2269);
and U1902 (N_1902,N_1313,N_776);
nand U1903 (N_1903,N_810,N_1124);
or U1904 (N_1904,N_1336,N_1234);
xor U1905 (N_1905,N_1331,In_1668);
and U1906 (N_1906,In_1064,In_1529);
and U1907 (N_1907,N_123,N_1141);
nand U1908 (N_1908,N_1044,N_939);
xnor U1909 (N_1909,N_700,N_1451);
and U1910 (N_1910,N_1222,In_1929);
xor U1911 (N_1911,N_1164,N_633);
and U1912 (N_1912,In_2113,In_793);
nand U1913 (N_1913,N_726,N_1450);
or U1914 (N_1914,In_1427,N_1042);
nor U1915 (N_1915,In_123,N_17);
xnor U1916 (N_1916,N_877,N_1066);
nand U1917 (N_1917,N_653,N_1441);
nand U1918 (N_1918,In_995,N_1380);
or U1919 (N_1919,N_1242,N_771);
nand U1920 (N_1920,N_1143,N_1417);
nor U1921 (N_1921,In_1938,N_206);
nand U1922 (N_1922,In_648,N_1121);
and U1923 (N_1923,N_1412,N_32);
or U1924 (N_1924,N_1489,N_1115);
xor U1925 (N_1925,N_616,N_1011);
or U1926 (N_1926,In_2229,N_1442);
xnor U1927 (N_1927,N_745,N_501);
or U1928 (N_1928,N_1126,N_1095);
nand U1929 (N_1929,N_1425,N_310);
and U1930 (N_1930,N_1312,N_1303);
xnor U1931 (N_1931,In_1713,N_855);
or U1932 (N_1932,N_281,N_538);
nand U1933 (N_1933,N_1026,N_1198);
xor U1934 (N_1934,N_422,N_1134);
and U1935 (N_1935,N_1022,In_1343);
nand U1936 (N_1936,N_1436,In_100);
nand U1937 (N_1937,In_952,N_1488);
and U1938 (N_1938,N_1014,In_1964);
nor U1939 (N_1939,N_1375,In_1825);
or U1940 (N_1940,N_1286,In_1571);
and U1941 (N_1941,N_1420,N_1359);
nand U1942 (N_1942,In_2391,N_1077);
nor U1943 (N_1943,N_1239,N_1491);
or U1944 (N_1944,N_1034,N_879);
nor U1945 (N_1945,In_1015,N_185);
or U1946 (N_1946,N_1029,In_1509);
or U1947 (N_1947,N_1073,In_933);
xnor U1948 (N_1948,N_1407,N_1278);
xor U1949 (N_1949,N_715,N_1357);
and U1950 (N_1950,In_1711,N_528);
nand U1951 (N_1951,N_883,In_1885);
nand U1952 (N_1952,N_973,In_2075);
xnor U1953 (N_1953,In_2195,N_551);
nor U1954 (N_1954,In_86,N_902);
or U1955 (N_1955,In_2071,N_1299);
nor U1956 (N_1956,N_1015,N_787);
nor U1957 (N_1957,N_525,N_1461);
or U1958 (N_1958,N_1112,N_1004);
nor U1959 (N_1959,N_217,N_572);
or U1960 (N_1960,N_1241,N_569);
xor U1961 (N_1961,N_845,N_1232);
nand U1962 (N_1962,N_15,N_1219);
and U1963 (N_1963,N_1474,N_1223);
and U1964 (N_1964,N_644,N_1373);
nor U1965 (N_1965,N_772,N_1348);
xor U1966 (N_1966,N_1154,N_690);
nand U1967 (N_1967,In_1146,In_1380);
nor U1968 (N_1968,N_800,N_1264);
nand U1969 (N_1969,N_1261,N_1311);
and U1970 (N_1970,N_813,N_1432);
or U1971 (N_1971,N_1007,N_890);
xor U1972 (N_1972,In_1472,N_1182);
or U1973 (N_1973,N_1197,N_1193);
or U1974 (N_1974,In_2194,In_229);
and U1975 (N_1975,N_857,N_1409);
nand U1976 (N_1976,In_1573,In_180);
and U1977 (N_1977,N_1452,N_53);
or U1978 (N_1978,N_1397,N_552);
nor U1979 (N_1979,N_1244,N_1247);
or U1980 (N_1980,N_1069,N_657);
nor U1981 (N_1981,N_55,N_1410);
nand U1982 (N_1982,N_1210,N_1406);
or U1983 (N_1983,N_323,N_1401);
nand U1984 (N_1984,N_1062,In_2257);
xor U1985 (N_1985,N_757,In_2091);
xnor U1986 (N_1986,N_728,N_1428);
xnor U1987 (N_1987,In_203,N_1315);
or U1988 (N_1988,In_1118,N_357);
nand U1989 (N_1989,N_560,N_1009);
xor U1990 (N_1990,N_140,In_344);
nor U1991 (N_1991,N_1093,N_1468);
or U1992 (N_1992,In_2303,N_1490);
or U1993 (N_1993,In_927,N_649);
nand U1994 (N_1994,N_1146,N_1090);
xnor U1995 (N_1995,N_1065,N_1497);
nand U1996 (N_1996,N_999,In_2284);
xor U1997 (N_1997,N_589,N_670);
xnor U1998 (N_1998,N_512,In_1798);
nor U1999 (N_1999,In_500,In_557);
nor U2000 (N_2000,N_1564,N_1651);
or U2001 (N_2001,N_1875,N_1613);
nor U2002 (N_2002,N_1593,N_1544);
or U2003 (N_2003,N_1937,N_1604);
nand U2004 (N_2004,N_1511,N_1567);
xnor U2005 (N_2005,N_1541,N_1524);
xnor U2006 (N_2006,N_1594,N_1628);
and U2007 (N_2007,N_1566,N_1685);
or U2008 (N_2008,N_1974,N_1636);
nand U2009 (N_2009,N_1716,N_1958);
nor U2010 (N_2010,N_1939,N_1905);
nor U2011 (N_2011,N_1765,N_1982);
and U2012 (N_2012,N_1851,N_1833);
nand U2013 (N_2013,N_1728,N_1714);
or U2014 (N_2014,N_1616,N_1673);
or U2015 (N_2015,N_1839,N_1523);
xor U2016 (N_2016,N_1510,N_1725);
nor U2017 (N_2017,N_1907,N_1549);
nor U2018 (N_2018,N_1602,N_1805);
xor U2019 (N_2019,N_1630,N_1644);
xnor U2020 (N_2020,N_1737,N_1852);
nor U2021 (N_2021,N_1731,N_1516);
and U2022 (N_2022,N_1595,N_1850);
or U2023 (N_2023,N_1619,N_1965);
nand U2024 (N_2024,N_1788,N_1626);
and U2025 (N_2025,N_1978,N_1950);
nand U2026 (N_2026,N_1704,N_1976);
or U2027 (N_2027,N_1821,N_1669);
xnor U2028 (N_2028,N_1944,N_1543);
nand U2029 (N_2029,N_1649,N_1586);
nor U2030 (N_2030,N_1598,N_1954);
and U2031 (N_2031,N_1755,N_1932);
and U2032 (N_2032,N_1941,N_1994);
nand U2033 (N_2033,N_1947,N_1710);
nor U2034 (N_2034,N_1911,N_1966);
or U2035 (N_2035,N_1512,N_1934);
or U2036 (N_2036,N_1938,N_1583);
xnor U2037 (N_2037,N_1534,N_1980);
and U2038 (N_2038,N_1676,N_1836);
nand U2039 (N_2039,N_1995,N_1760);
nor U2040 (N_2040,N_1761,N_1736);
or U2041 (N_2041,N_1824,N_1927);
nor U2042 (N_2042,N_1780,N_1580);
nor U2043 (N_2043,N_1642,N_1589);
or U2044 (N_2044,N_1531,N_1828);
and U2045 (N_2045,N_1521,N_1734);
nor U2046 (N_2046,N_1538,N_1525);
and U2047 (N_2047,N_1945,N_1967);
or U2048 (N_2048,N_1518,N_1658);
nand U2049 (N_2049,N_1827,N_1720);
xor U2050 (N_2050,N_1849,N_1989);
nand U2051 (N_2051,N_1554,N_1930);
xor U2052 (N_2052,N_1777,N_1822);
and U2053 (N_2053,N_1575,N_1551);
and U2054 (N_2054,N_1587,N_1555);
or U2055 (N_2055,N_1897,N_1910);
and U2056 (N_2056,N_1817,N_1743);
nor U2057 (N_2057,N_1870,N_1834);
xor U2058 (N_2058,N_1763,N_1860);
or U2059 (N_2059,N_1574,N_1527);
and U2060 (N_2060,N_1672,N_1674);
or U2061 (N_2061,N_1882,N_1610);
nand U2062 (N_2062,N_1773,N_1590);
and U2063 (N_2063,N_1906,N_1768);
nor U2064 (N_2064,N_1711,N_1520);
and U2065 (N_2065,N_1991,N_1659);
xor U2066 (N_2066,N_1621,N_1996);
and U2067 (N_2067,N_1802,N_1746);
and U2068 (N_2068,N_1745,N_1990);
and U2069 (N_2069,N_1916,N_1874);
and U2070 (N_2070,N_1796,N_1936);
xor U2071 (N_2071,N_1638,N_1603);
xor U2072 (N_2072,N_1691,N_1885);
or U2073 (N_2073,N_1748,N_1539);
xor U2074 (N_2074,N_1793,N_1565);
nand U2075 (N_2075,N_1559,N_1979);
and U2076 (N_2076,N_1584,N_1942);
xnor U2077 (N_2077,N_1912,N_1892);
nor U2078 (N_2078,N_1902,N_1623);
nor U2079 (N_2079,N_1957,N_1532);
xnor U2080 (N_2080,N_1506,N_1722);
nor U2081 (N_2081,N_1650,N_1992);
nor U2082 (N_2082,N_1858,N_1770);
nor U2083 (N_2083,N_1960,N_1984);
or U2084 (N_2084,N_1964,N_1914);
and U2085 (N_2085,N_1867,N_1571);
or U2086 (N_2086,N_1985,N_1764);
xor U2087 (N_2087,N_1835,N_1872);
nand U2088 (N_2088,N_1536,N_1702);
nand U2089 (N_2089,N_1504,N_1781);
or U2090 (N_2090,N_1733,N_1522);
nand U2091 (N_2091,N_1550,N_1920);
and U2092 (N_2092,N_1675,N_1678);
nor U2093 (N_2093,N_1782,N_1861);
or U2094 (N_2094,N_1883,N_1791);
nand U2095 (N_2095,N_1726,N_1847);
and U2096 (N_2096,N_1500,N_1749);
nand U2097 (N_2097,N_1776,N_1918);
xor U2098 (N_2098,N_1792,N_1772);
nand U2099 (N_2099,N_1513,N_1816);
or U2100 (N_2100,N_1668,N_1663);
nand U2101 (N_2101,N_1854,N_1786);
nor U2102 (N_2102,N_1712,N_1609);
nor U2103 (N_2103,N_1687,N_1935);
nand U2104 (N_2104,N_1730,N_1643);
or U2105 (N_2105,N_1767,N_1751);
and U2106 (N_2106,N_1607,N_1963);
nor U2107 (N_2107,N_1693,N_1876);
nand U2108 (N_2108,N_1640,N_1614);
nand U2109 (N_2109,N_1624,N_1620);
nor U2110 (N_2110,N_1837,N_1840);
xor U2111 (N_2111,N_1787,N_1740);
nor U2112 (N_2112,N_1878,N_1661);
and U2113 (N_2113,N_1929,N_1856);
or U2114 (N_2114,N_1970,N_1646);
nor U2115 (N_2115,N_1535,N_1709);
and U2116 (N_2116,N_1913,N_1825);
or U2117 (N_2117,N_1832,N_1666);
and U2118 (N_2118,N_1533,N_1601);
and U2119 (N_2119,N_1799,N_1877);
nor U2120 (N_2120,N_1826,N_1612);
xnor U2121 (N_2121,N_1625,N_1810);
and U2122 (N_2122,N_1997,N_1697);
or U2123 (N_2123,N_1706,N_1975);
nand U2124 (N_2124,N_1775,N_1808);
nand U2125 (N_2125,N_1893,N_1784);
or U2126 (N_2126,N_1739,N_1841);
and U2127 (N_2127,N_1507,N_1648);
xnor U2128 (N_2128,N_1540,N_1868);
nor U2129 (N_2129,N_1968,N_1701);
xor U2130 (N_2130,N_1798,N_1732);
nor U2131 (N_2131,N_1946,N_1896);
nand U2132 (N_2132,N_1573,N_1608);
xor U2133 (N_2133,N_1591,N_1909);
nor U2134 (N_2134,N_1656,N_1599);
or U2135 (N_2135,N_1560,N_1880);
xor U2136 (N_2136,N_1509,N_1542);
and U2137 (N_2137,N_1569,N_1812);
xnor U2138 (N_2138,N_1708,N_1694);
xor U2139 (N_2139,N_1677,N_1572);
nor U2140 (N_2140,N_1742,N_1700);
nor U2141 (N_2141,N_1953,N_1806);
xnor U2142 (N_2142,N_1752,N_1629);
and U2143 (N_2143,N_1959,N_1688);
nor U2144 (N_2144,N_1890,N_1895);
nand U2145 (N_2145,N_1662,N_1859);
nor U2146 (N_2146,N_1718,N_1999);
and U2147 (N_2147,N_1756,N_1577);
or U2148 (N_2148,N_1923,N_1771);
and U2149 (N_2149,N_1652,N_1615);
or U2150 (N_2150,N_1800,N_1705);
and U2151 (N_2151,N_1690,N_1757);
xnor U2152 (N_2152,N_1981,N_1886);
or U2153 (N_2153,N_1972,N_1961);
and U2154 (N_2154,N_1528,N_1622);
and U2155 (N_2155,N_1881,N_1738);
nand U2156 (N_2156,N_1552,N_1795);
nand U2157 (N_2157,N_1790,N_1797);
and U2158 (N_2158,N_1545,N_1631);
and U2159 (N_2159,N_1955,N_1557);
nand U2160 (N_2160,N_1900,N_1818);
or U2161 (N_2161,N_1919,N_1655);
or U2162 (N_2162,N_1843,N_1888);
xor U2163 (N_2163,N_1546,N_1759);
xnor U2164 (N_2164,N_1887,N_1653);
or U2165 (N_2165,N_1721,N_1848);
xor U2166 (N_2166,N_1943,N_1667);
xor U2167 (N_2167,N_1921,N_1830);
xnor U2168 (N_2168,N_1588,N_1986);
nand U2169 (N_2169,N_1993,N_1926);
xnor U2170 (N_2170,N_1689,N_1820);
and U2171 (N_2171,N_1505,N_1562);
nand U2172 (N_2172,N_1842,N_1682);
nor U2173 (N_2173,N_1845,N_1962);
nand U2174 (N_2174,N_1719,N_1903);
and U2175 (N_2175,N_1537,N_1794);
nand U2176 (N_2176,N_1563,N_1568);
and U2177 (N_2177,N_1951,N_1683);
or U2178 (N_2178,N_1600,N_1846);
nor U2179 (N_2179,N_1547,N_1724);
or U2180 (N_2180,N_1741,N_1684);
nor U2181 (N_2181,N_1679,N_1898);
nand U2182 (N_2182,N_1618,N_1908);
or U2183 (N_2183,N_1879,N_1634);
or U2184 (N_2184,N_1699,N_1635);
or U2185 (N_2185,N_1713,N_1924);
or U2186 (N_2186,N_1815,N_1519);
and U2187 (N_2187,N_1804,N_1809);
and U2188 (N_2188,N_1639,N_1735);
nand U2189 (N_2189,N_1977,N_1948);
nor U2190 (N_2190,N_1758,N_1811);
nor U2191 (N_2191,N_1660,N_1855);
xor U2192 (N_2192,N_1863,N_1889);
nand U2193 (N_2193,N_1707,N_1973);
nand U2194 (N_2194,N_1823,N_1696);
xor U2195 (N_2195,N_1891,N_1779);
and U2196 (N_2196,N_1884,N_1515);
and U2197 (N_2197,N_1917,N_1664);
nor U2198 (N_2198,N_1969,N_1899);
xor U2199 (N_2199,N_1671,N_1592);
or U2200 (N_2200,N_1931,N_1581);
xnor U2201 (N_2201,N_1762,N_1647);
and U2202 (N_2202,N_1915,N_1692);
and U2203 (N_2203,N_1556,N_1750);
and U2204 (N_2204,N_1998,N_1933);
nand U2205 (N_2205,N_1727,N_1952);
and U2206 (N_2206,N_1596,N_1717);
nor U2207 (N_2207,N_1831,N_1838);
nand U2208 (N_2208,N_1789,N_1949);
nand U2209 (N_2209,N_1627,N_1695);
and U2210 (N_2210,N_1747,N_1853);
or U2211 (N_2211,N_1925,N_1502);
or U2212 (N_2212,N_1654,N_1829);
or U2213 (N_2213,N_1922,N_1753);
xnor U2214 (N_2214,N_1778,N_1570);
or U2215 (N_2215,N_1501,N_1605);
nand U2216 (N_2216,N_1987,N_1637);
nand U2217 (N_2217,N_1928,N_1611);
or U2218 (N_2218,N_1579,N_1814);
nor U2219 (N_2219,N_1582,N_1813);
and U2220 (N_2220,N_1641,N_1801);
nor U2221 (N_2221,N_1723,N_1866);
nand U2222 (N_2222,N_1657,N_1783);
nor U2223 (N_2223,N_1988,N_1526);
xor U2224 (N_2224,N_1803,N_1894);
xor U2225 (N_2225,N_1632,N_1971);
nand U2226 (N_2226,N_1904,N_1869);
nor U2227 (N_2227,N_1617,N_1585);
xor U2228 (N_2228,N_1956,N_1807);
or U2229 (N_2229,N_1871,N_1940);
xor U2230 (N_2230,N_1503,N_1715);
nand U2231 (N_2231,N_1785,N_1744);
or U2232 (N_2232,N_1901,N_1983);
nand U2233 (N_2233,N_1864,N_1681);
nor U2234 (N_2234,N_1517,N_1548);
nor U2235 (N_2235,N_1606,N_1754);
nand U2236 (N_2236,N_1865,N_1769);
and U2237 (N_2237,N_1508,N_1576);
xor U2238 (N_2238,N_1862,N_1703);
xor U2239 (N_2239,N_1680,N_1857);
and U2240 (N_2240,N_1670,N_1645);
nor U2241 (N_2241,N_1873,N_1558);
nor U2242 (N_2242,N_1729,N_1597);
and U2243 (N_2243,N_1561,N_1774);
xnor U2244 (N_2244,N_1553,N_1665);
nand U2245 (N_2245,N_1698,N_1578);
or U2246 (N_2246,N_1686,N_1530);
xnor U2247 (N_2247,N_1766,N_1514);
xor U2248 (N_2248,N_1844,N_1633);
nor U2249 (N_2249,N_1529,N_1819);
nor U2250 (N_2250,N_1790,N_1838);
nor U2251 (N_2251,N_1582,N_1796);
or U2252 (N_2252,N_1563,N_1633);
nand U2253 (N_2253,N_1672,N_1616);
and U2254 (N_2254,N_1675,N_1564);
or U2255 (N_2255,N_1867,N_1612);
nand U2256 (N_2256,N_1776,N_1934);
nor U2257 (N_2257,N_1555,N_1837);
nand U2258 (N_2258,N_1675,N_1813);
nor U2259 (N_2259,N_1850,N_1503);
nand U2260 (N_2260,N_1819,N_1869);
nor U2261 (N_2261,N_1826,N_1689);
nand U2262 (N_2262,N_1800,N_1995);
or U2263 (N_2263,N_1520,N_1635);
or U2264 (N_2264,N_1978,N_1765);
nand U2265 (N_2265,N_1956,N_1603);
xor U2266 (N_2266,N_1804,N_1709);
nand U2267 (N_2267,N_1776,N_1842);
or U2268 (N_2268,N_1924,N_1754);
xor U2269 (N_2269,N_1956,N_1986);
xnor U2270 (N_2270,N_1569,N_1874);
and U2271 (N_2271,N_1862,N_1992);
or U2272 (N_2272,N_1744,N_1865);
xnor U2273 (N_2273,N_1754,N_1851);
nor U2274 (N_2274,N_1940,N_1727);
nor U2275 (N_2275,N_1572,N_1590);
nand U2276 (N_2276,N_1524,N_1880);
nor U2277 (N_2277,N_1952,N_1666);
and U2278 (N_2278,N_1855,N_1815);
xor U2279 (N_2279,N_1852,N_1772);
nor U2280 (N_2280,N_1717,N_1811);
nand U2281 (N_2281,N_1549,N_1894);
and U2282 (N_2282,N_1905,N_1790);
nand U2283 (N_2283,N_1839,N_1991);
nand U2284 (N_2284,N_1765,N_1535);
nand U2285 (N_2285,N_1647,N_1751);
or U2286 (N_2286,N_1624,N_1879);
nor U2287 (N_2287,N_1841,N_1505);
xor U2288 (N_2288,N_1953,N_1816);
or U2289 (N_2289,N_1714,N_1875);
nand U2290 (N_2290,N_1857,N_1662);
nor U2291 (N_2291,N_1564,N_1782);
xnor U2292 (N_2292,N_1838,N_1507);
nor U2293 (N_2293,N_1889,N_1959);
nor U2294 (N_2294,N_1611,N_1544);
nor U2295 (N_2295,N_1826,N_1667);
and U2296 (N_2296,N_1614,N_1652);
nor U2297 (N_2297,N_1889,N_1607);
and U2298 (N_2298,N_1781,N_1819);
nand U2299 (N_2299,N_1895,N_1727);
nor U2300 (N_2300,N_1848,N_1958);
xnor U2301 (N_2301,N_1588,N_1691);
or U2302 (N_2302,N_1557,N_1996);
xnor U2303 (N_2303,N_1929,N_1667);
or U2304 (N_2304,N_1886,N_1906);
nor U2305 (N_2305,N_1529,N_1905);
nand U2306 (N_2306,N_1981,N_1943);
and U2307 (N_2307,N_1982,N_1550);
nor U2308 (N_2308,N_1962,N_1990);
and U2309 (N_2309,N_1877,N_1673);
nor U2310 (N_2310,N_1768,N_1938);
xor U2311 (N_2311,N_1879,N_1543);
nor U2312 (N_2312,N_1542,N_1927);
or U2313 (N_2313,N_1776,N_1979);
and U2314 (N_2314,N_1964,N_1542);
nand U2315 (N_2315,N_1557,N_1645);
xor U2316 (N_2316,N_1520,N_1961);
or U2317 (N_2317,N_1830,N_1607);
nand U2318 (N_2318,N_1930,N_1538);
nor U2319 (N_2319,N_1840,N_1902);
nor U2320 (N_2320,N_1626,N_1808);
xnor U2321 (N_2321,N_1743,N_1752);
nand U2322 (N_2322,N_1767,N_1539);
xor U2323 (N_2323,N_1557,N_1897);
nor U2324 (N_2324,N_1862,N_1902);
nand U2325 (N_2325,N_1796,N_1650);
nor U2326 (N_2326,N_1619,N_1954);
nand U2327 (N_2327,N_1661,N_1561);
nand U2328 (N_2328,N_1975,N_1851);
xnor U2329 (N_2329,N_1602,N_1674);
xor U2330 (N_2330,N_1882,N_1725);
nor U2331 (N_2331,N_1590,N_1698);
xor U2332 (N_2332,N_1658,N_1558);
and U2333 (N_2333,N_1913,N_1887);
nor U2334 (N_2334,N_1563,N_1674);
or U2335 (N_2335,N_1660,N_1830);
nand U2336 (N_2336,N_1578,N_1994);
nor U2337 (N_2337,N_1529,N_1976);
nand U2338 (N_2338,N_1905,N_1770);
nor U2339 (N_2339,N_1519,N_1809);
xnor U2340 (N_2340,N_1957,N_1689);
nand U2341 (N_2341,N_1590,N_1501);
xor U2342 (N_2342,N_1774,N_1576);
xor U2343 (N_2343,N_1673,N_1955);
nor U2344 (N_2344,N_1943,N_1552);
nand U2345 (N_2345,N_1758,N_1575);
nand U2346 (N_2346,N_1944,N_1617);
nor U2347 (N_2347,N_1702,N_1592);
xor U2348 (N_2348,N_1622,N_1579);
nand U2349 (N_2349,N_1986,N_1763);
or U2350 (N_2350,N_1784,N_1708);
nor U2351 (N_2351,N_1613,N_1645);
or U2352 (N_2352,N_1546,N_1677);
xor U2353 (N_2353,N_1933,N_1728);
nand U2354 (N_2354,N_1681,N_1691);
and U2355 (N_2355,N_1612,N_1534);
or U2356 (N_2356,N_1737,N_1583);
and U2357 (N_2357,N_1909,N_1805);
and U2358 (N_2358,N_1906,N_1850);
or U2359 (N_2359,N_1864,N_1991);
or U2360 (N_2360,N_1833,N_1654);
and U2361 (N_2361,N_1961,N_1870);
and U2362 (N_2362,N_1845,N_1661);
and U2363 (N_2363,N_1921,N_1704);
xor U2364 (N_2364,N_1528,N_1520);
xnor U2365 (N_2365,N_1772,N_1932);
and U2366 (N_2366,N_1975,N_1858);
or U2367 (N_2367,N_1610,N_1550);
nand U2368 (N_2368,N_1826,N_1961);
or U2369 (N_2369,N_1901,N_1631);
and U2370 (N_2370,N_1695,N_1704);
nand U2371 (N_2371,N_1636,N_1743);
or U2372 (N_2372,N_1731,N_1740);
or U2373 (N_2373,N_1660,N_1842);
and U2374 (N_2374,N_1667,N_1891);
nand U2375 (N_2375,N_1773,N_1694);
and U2376 (N_2376,N_1671,N_1998);
or U2377 (N_2377,N_1815,N_1646);
and U2378 (N_2378,N_1946,N_1670);
and U2379 (N_2379,N_1662,N_1955);
or U2380 (N_2380,N_1996,N_1693);
nand U2381 (N_2381,N_1935,N_1642);
or U2382 (N_2382,N_1700,N_1699);
or U2383 (N_2383,N_1511,N_1916);
and U2384 (N_2384,N_1533,N_1998);
nand U2385 (N_2385,N_1926,N_1637);
xor U2386 (N_2386,N_1873,N_1553);
and U2387 (N_2387,N_1887,N_1762);
xor U2388 (N_2388,N_1893,N_1559);
and U2389 (N_2389,N_1860,N_1778);
or U2390 (N_2390,N_1521,N_1917);
nand U2391 (N_2391,N_1805,N_1655);
and U2392 (N_2392,N_1976,N_1663);
nor U2393 (N_2393,N_1662,N_1711);
nor U2394 (N_2394,N_1653,N_1776);
and U2395 (N_2395,N_1868,N_1587);
nor U2396 (N_2396,N_1912,N_1858);
nor U2397 (N_2397,N_1612,N_1842);
xor U2398 (N_2398,N_1666,N_1589);
nand U2399 (N_2399,N_1802,N_1837);
xor U2400 (N_2400,N_1556,N_1595);
xor U2401 (N_2401,N_1975,N_1549);
nand U2402 (N_2402,N_1850,N_1902);
xor U2403 (N_2403,N_1653,N_1782);
or U2404 (N_2404,N_1759,N_1988);
and U2405 (N_2405,N_1922,N_1854);
nor U2406 (N_2406,N_1841,N_1690);
or U2407 (N_2407,N_1589,N_1754);
nor U2408 (N_2408,N_1964,N_1801);
and U2409 (N_2409,N_1883,N_1667);
nand U2410 (N_2410,N_1911,N_1624);
and U2411 (N_2411,N_1835,N_1777);
and U2412 (N_2412,N_1716,N_1783);
and U2413 (N_2413,N_1637,N_1809);
nor U2414 (N_2414,N_1651,N_1734);
or U2415 (N_2415,N_1880,N_1700);
or U2416 (N_2416,N_1874,N_1900);
or U2417 (N_2417,N_1883,N_1733);
and U2418 (N_2418,N_1647,N_1543);
and U2419 (N_2419,N_1778,N_1992);
nand U2420 (N_2420,N_1631,N_1982);
nand U2421 (N_2421,N_1808,N_1805);
and U2422 (N_2422,N_1840,N_1836);
and U2423 (N_2423,N_1838,N_1916);
nor U2424 (N_2424,N_1878,N_1572);
nand U2425 (N_2425,N_1694,N_1963);
and U2426 (N_2426,N_1868,N_1624);
and U2427 (N_2427,N_1739,N_1530);
xor U2428 (N_2428,N_1654,N_1527);
or U2429 (N_2429,N_1684,N_1657);
and U2430 (N_2430,N_1594,N_1677);
nand U2431 (N_2431,N_1674,N_1653);
nor U2432 (N_2432,N_1514,N_1829);
nand U2433 (N_2433,N_1692,N_1732);
and U2434 (N_2434,N_1857,N_1843);
xnor U2435 (N_2435,N_1745,N_1600);
nand U2436 (N_2436,N_1978,N_1882);
and U2437 (N_2437,N_1906,N_1774);
and U2438 (N_2438,N_1866,N_1855);
or U2439 (N_2439,N_1816,N_1870);
nor U2440 (N_2440,N_1773,N_1627);
nand U2441 (N_2441,N_1502,N_1979);
nand U2442 (N_2442,N_1734,N_1913);
or U2443 (N_2443,N_1567,N_1978);
nand U2444 (N_2444,N_1816,N_1823);
and U2445 (N_2445,N_1811,N_1618);
xnor U2446 (N_2446,N_1851,N_1840);
or U2447 (N_2447,N_1982,N_1770);
and U2448 (N_2448,N_1972,N_1923);
nor U2449 (N_2449,N_1506,N_1910);
xor U2450 (N_2450,N_1552,N_1543);
xor U2451 (N_2451,N_1644,N_1915);
and U2452 (N_2452,N_1565,N_1639);
xor U2453 (N_2453,N_1544,N_1562);
and U2454 (N_2454,N_1556,N_1672);
nor U2455 (N_2455,N_1860,N_1672);
or U2456 (N_2456,N_1715,N_1641);
nand U2457 (N_2457,N_1919,N_1977);
nor U2458 (N_2458,N_1970,N_1791);
nor U2459 (N_2459,N_1535,N_1879);
and U2460 (N_2460,N_1666,N_1513);
nor U2461 (N_2461,N_1665,N_1567);
xnor U2462 (N_2462,N_1818,N_1959);
nand U2463 (N_2463,N_1660,N_1773);
xor U2464 (N_2464,N_1753,N_1556);
xor U2465 (N_2465,N_1751,N_1858);
xor U2466 (N_2466,N_1553,N_1558);
xor U2467 (N_2467,N_1900,N_1843);
and U2468 (N_2468,N_1675,N_1521);
nor U2469 (N_2469,N_1535,N_1526);
xnor U2470 (N_2470,N_1968,N_1575);
nor U2471 (N_2471,N_1986,N_1526);
xor U2472 (N_2472,N_1877,N_1935);
nor U2473 (N_2473,N_1555,N_1951);
or U2474 (N_2474,N_1960,N_1831);
or U2475 (N_2475,N_1647,N_1788);
nor U2476 (N_2476,N_1965,N_1523);
xor U2477 (N_2477,N_1779,N_1967);
nand U2478 (N_2478,N_1665,N_1934);
nor U2479 (N_2479,N_1953,N_1950);
nand U2480 (N_2480,N_1566,N_1832);
or U2481 (N_2481,N_1513,N_1687);
nor U2482 (N_2482,N_1660,N_1813);
and U2483 (N_2483,N_1925,N_1671);
xor U2484 (N_2484,N_1823,N_1907);
and U2485 (N_2485,N_1956,N_1650);
xor U2486 (N_2486,N_1676,N_1554);
nor U2487 (N_2487,N_1756,N_1516);
and U2488 (N_2488,N_1666,N_1578);
nor U2489 (N_2489,N_1684,N_1692);
or U2490 (N_2490,N_1764,N_1581);
and U2491 (N_2491,N_1845,N_1581);
nand U2492 (N_2492,N_1628,N_1707);
xor U2493 (N_2493,N_1846,N_1704);
or U2494 (N_2494,N_1777,N_1600);
and U2495 (N_2495,N_1643,N_1848);
and U2496 (N_2496,N_1954,N_1543);
or U2497 (N_2497,N_1819,N_1608);
nor U2498 (N_2498,N_1937,N_1508);
and U2499 (N_2499,N_1830,N_1579);
or U2500 (N_2500,N_2387,N_2246);
or U2501 (N_2501,N_2239,N_2057);
or U2502 (N_2502,N_2376,N_2398);
or U2503 (N_2503,N_2178,N_2261);
or U2504 (N_2504,N_2386,N_2306);
xor U2505 (N_2505,N_2450,N_2379);
or U2506 (N_2506,N_2277,N_2392);
or U2507 (N_2507,N_2226,N_2099);
xnor U2508 (N_2508,N_2391,N_2173);
and U2509 (N_2509,N_2230,N_2124);
xnor U2510 (N_2510,N_2498,N_2161);
nor U2511 (N_2511,N_2445,N_2499);
xor U2512 (N_2512,N_2107,N_2443);
xnor U2513 (N_2513,N_2065,N_2263);
xnor U2514 (N_2514,N_2265,N_2411);
nor U2515 (N_2515,N_2211,N_2412);
xor U2516 (N_2516,N_2356,N_2399);
nand U2517 (N_2517,N_2217,N_2334);
and U2518 (N_2518,N_2479,N_2336);
nor U2519 (N_2519,N_2153,N_2472);
or U2520 (N_2520,N_2458,N_2191);
xor U2521 (N_2521,N_2313,N_2342);
or U2522 (N_2522,N_2011,N_2007);
nor U2523 (N_2523,N_2468,N_2378);
xnor U2524 (N_2524,N_2419,N_2372);
and U2525 (N_2525,N_2351,N_2492);
nand U2526 (N_2526,N_2421,N_2118);
xor U2527 (N_2527,N_2081,N_2369);
xnor U2528 (N_2528,N_2119,N_2070);
and U2529 (N_2529,N_2112,N_2269);
xor U2530 (N_2530,N_2426,N_2255);
xnor U2531 (N_2531,N_2290,N_2035);
xor U2532 (N_2532,N_2475,N_2234);
nand U2533 (N_2533,N_2013,N_2402);
and U2534 (N_2534,N_2061,N_2141);
nor U2535 (N_2535,N_2100,N_2190);
xnor U2536 (N_2536,N_2159,N_2497);
and U2537 (N_2537,N_2270,N_2338);
xnor U2538 (N_2538,N_2415,N_2477);
xnor U2539 (N_2539,N_2375,N_2194);
nor U2540 (N_2540,N_2340,N_2483);
nand U2541 (N_2541,N_2046,N_2276);
xor U2542 (N_2542,N_2327,N_2051);
or U2543 (N_2543,N_2082,N_2127);
and U2544 (N_2544,N_2158,N_2353);
nand U2545 (N_2545,N_2203,N_2397);
or U2546 (N_2546,N_2320,N_2478);
xnor U2547 (N_2547,N_2089,N_2489);
nor U2548 (N_2548,N_2060,N_2400);
xnor U2549 (N_2549,N_2037,N_2389);
and U2550 (N_2550,N_2009,N_2097);
and U2551 (N_2551,N_2449,N_2147);
xor U2552 (N_2552,N_2283,N_2052);
and U2553 (N_2553,N_2197,N_2288);
and U2554 (N_2554,N_2145,N_2018);
nand U2555 (N_2555,N_2362,N_2106);
nand U2556 (N_2556,N_2414,N_2062);
nand U2557 (N_2557,N_2413,N_2245);
and U2558 (N_2558,N_2078,N_2408);
and U2559 (N_2559,N_2388,N_2136);
or U2560 (N_2560,N_2019,N_2028);
nand U2561 (N_2561,N_2222,N_2115);
nand U2562 (N_2562,N_2359,N_2325);
xnor U2563 (N_2563,N_2303,N_2022);
xor U2564 (N_2564,N_2451,N_2132);
nor U2565 (N_2565,N_2485,N_2014);
and U2566 (N_2566,N_2300,N_2355);
or U2567 (N_2567,N_2491,N_2071);
nand U2568 (N_2568,N_2495,N_2461);
xnor U2569 (N_2569,N_2224,N_2252);
or U2570 (N_2570,N_2405,N_2015);
or U2571 (N_2571,N_2010,N_2347);
nor U2572 (N_2572,N_2103,N_2020);
or U2573 (N_2573,N_2464,N_2282);
and U2574 (N_2574,N_2429,N_2123);
or U2575 (N_2575,N_2098,N_2446);
xor U2576 (N_2576,N_2248,N_2243);
and U2577 (N_2577,N_2104,N_2213);
xnor U2578 (N_2578,N_2436,N_2095);
and U2579 (N_2579,N_2278,N_2292);
or U2580 (N_2580,N_2091,N_2208);
xor U2581 (N_2581,N_2148,N_2382);
nor U2582 (N_2582,N_2108,N_2349);
or U2583 (N_2583,N_2048,N_2033);
nor U2584 (N_2584,N_2202,N_2316);
nand U2585 (N_2585,N_2326,N_2096);
xor U2586 (N_2586,N_2371,N_2343);
nand U2587 (N_2587,N_2184,N_2357);
or U2588 (N_2588,N_2437,N_2006);
and U2589 (N_2589,N_2040,N_2434);
nand U2590 (N_2590,N_2162,N_2044);
and U2591 (N_2591,N_2187,N_2249);
or U2592 (N_2592,N_2486,N_2182);
nor U2593 (N_2593,N_2469,N_2189);
nor U2594 (N_2594,N_2286,N_2215);
and U2595 (N_2595,N_2370,N_2385);
xnor U2596 (N_2596,N_2487,N_2134);
or U2597 (N_2597,N_2396,N_2142);
or U2598 (N_2598,N_2474,N_2031);
nor U2599 (N_2599,N_2420,N_2348);
and U2600 (N_2600,N_2305,N_2237);
and U2601 (N_2601,N_2333,N_2253);
or U2602 (N_2602,N_2465,N_2418);
or U2603 (N_2603,N_2125,N_2318);
or U2604 (N_2604,N_2409,N_2235);
nor U2605 (N_2605,N_2068,N_2242);
xor U2606 (N_2606,N_2144,N_2149);
nor U2607 (N_2607,N_2001,N_2043);
and U2608 (N_2608,N_2428,N_2012);
or U2609 (N_2609,N_2188,N_2133);
nor U2610 (N_2610,N_2105,N_2076);
xnor U2611 (N_2611,N_2319,N_2023);
nand U2612 (N_2612,N_2181,N_2274);
nor U2613 (N_2613,N_2488,N_2185);
nor U2614 (N_2614,N_2030,N_2176);
nand U2615 (N_2615,N_2111,N_2496);
nand U2616 (N_2616,N_2467,N_2287);
xor U2617 (N_2617,N_2170,N_2207);
xnor U2618 (N_2618,N_2317,N_2410);
nor U2619 (N_2619,N_2077,N_2271);
and U2620 (N_2620,N_2135,N_2085);
nand U2621 (N_2621,N_2452,N_2383);
xnor U2622 (N_2622,N_2481,N_2175);
xnor U2623 (N_2623,N_2093,N_2140);
nand U2624 (N_2624,N_2435,N_2150);
nand U2625 (N_2625,N_2427,N_2312);
nand U2626 (N_2626,N_2262,N_2110);
nor U2627 (N_2627,N_2291,N_2193);
nand U2628 (N_2628,N_2373,N_2216);
or U2629 (N_2629,N_2328,N_2214);
nor U2630 (N_2630,N_2027,N_2000);
xor U2631 (N_2631,N_2201,N_2024);
and U2632 (N_2632,N_2247,N_2352);
nor U2633 (N_2633,N_2032,N_2180);
xnor U2634 (N_2634,N_2354,N_2120);
xnor U2635 (N_2635,N_2459,N_2160);
xnor U2636 (N_2636,N_2155,N_2460);
or U2637 (N_2637,N_2425,N_2301);
and U2638 (N_2638,N_2102,N_2494);
and U2639 (N_2639,N_2116,N_2337);
or U2640 (N_2640,N_2374,N_2165);
xnor U2641 (N_2641,N_2361,N_2063);
and U2642 (N_2642,N_2439,N_2285);
and U2643 (N_2643,N_2205,N_2039);
nor U2644 (N_2644,N_2322,N_2315);
or U2645 (N_2645,N_2447,N_2209);
and U2646 (N_2646,N_2232,N_2090);
or U2647 (N_2647,N_2130,N_2302);
nand U2648 (N_2648,N_2101,N_2395);
nor U2649 (N_2649,N_2053,N_2131);
xnor U2650 (N_2650,N_2422,N_2471);
or U2651 (N_2651,N_2438,N_2067);
or U2652 (N_2652,N_2219,N_2368);
or U2653 (N_2653,N_2143,N_2050);
and U2654 (N_2654,N_2284,N_2117);
xnor U2655 (N_2655,N_2056,N_2365);
and U2656 (N_2656,N_2138,N_2266);
or U2657 (N_2657,N_2025,N_2304);
and U2658 (N_2658,N_2059,N_2168);
or U2659 (N_2659,N_2146,N_2186);
and U2660 (N_2660,N_2254,N_2042);
or U2661 (N_2661,N_2114,N_2324);
xor U2662 (N_2662,N_2416,N_2021);
or U2663 (N_2663,N_2323,N_2473);
nor U2664 (N_2664,N_2250,N_2331);
and U2665 (N_2665,N_2058,N_2272);
and U2666 (N_2666,N_2454,N_2074);
or U2667 (N_2667,N_2453,N_2199);
and U2668 (N_2668,N_2212,N_2003);
nand U2669 (N_2669,N_2448,N_2251);
or U2670 (N_2670,N_2360,N_2164);
and U2671 (N_2671,N_2423,N_2220);
nand U2672 (N_2672,N_2268,N_2179);
nand U2673 (N_2673,N_2086,N_2256);
and U2674 (N_2674,N_2345,N_2047);
nand U2675 (N_2675,N_2476,N_2433);
nor U2676 (N_2676,N_2005,N_2083);
and U2677 (N_2677,N_2281,N_2380);
or U2678 (N_2678,N_2238,N_2137);
nand U2679 (N_2679,N_2169,N_2192);
and U2680 (N_2680,N_2075,N_2299);
nor U2681 (N_2681,N_2417,N_2484);
nand U2682 (N_2682,N_2126,N_2297);
nand U2683 (N_2683,N_2321,N_2157);
or U2684 (N_2684,N_2258,N_2041);
nand U2685 (N_2685,N_2094,N_2339);
nand U2686 (N_2686,N_2172,N_2384);
or U2687 (N_2687,N_2335,N_2390);
or U2688 (N_2688,N_2279,N_2457);
xnor U2689 (N_2689,N_2004,N_2069);
and U2690 (N_2690,N_2377,N_2204);
xor U2691 (N_2691,N_2171,N_2314);
and U2692 (N_2692,N_2480,N_2442);
nor U2693 (N_2693,N_2330,N_2311);
nand U2694 (N_2694,N_2294,N_2257);
nand U2695 (N_2695,N_2231,N_2432);
or U2696 (N_2696,N_2295,N_2198);
xnor U2697 (N_2697,N_2393,N_2072);
and U2698 (N_2698,N_2309,N_2228);
xor U2699 (N_2699,N_2407,N_2151);
nor U2700 (N_2700,N_2403,N_2308);
nor U2701 (N_2701,N_2275,N_2195);
or U2702 (N_2702,N_2406,N_2087);
nor U2703 (N_2703,N_2455,N_2394);
nand U2704 (N_2704,N_2128,N_2260);
nand U2705 (N_2705,N_2367,N_2092);
or U2706 (N_2706,N_2240,N_2358);
and U2707 (N_2707,N_2241,N_2167);
xnor U2708 (N_2708,N_2259,N_2152);
nand U2709 (N_2709,N_2470,N_2364);
nor U2710 (N_2710,N_2200,N_2493);
nor U2711 (N_2711,N_2049,N_2332);
xor U2712 (N_2712,N_2344,N_2002);
or U2713 (N_2713,N_2462,N_2034);
and U2714 (N_2714,N_2431,N_2066);
and U2715 (N_2715,N_2366,N_2036);
nand U2716 (N_2716,N_2139,N_2008);
and U2717 (N_2717,N_2298,N_2223);
and U2718 (N_2718,N_2440,N_2154);
nand U2719 (N_2719,N_2401,N_2026);
xor U2720 (N_2720,N_2221,N_2054);
and U2721 (N_2721,N_2045,N_2490);
and U2722 (N_2722,N_2079,N_2463);
or U2723 (N_2723,N_2381,N_2177);
and U2724 (N_2724,N_2273,N_2233);
nor U2725 (N_2725,N_2163,N_2196);
nor U2726 (N_2726,N_2113,N_2329);
or U2727 (N_2727,N_2227,N_2236);
nand U2728 (N_2728,N_2307,N_2156);
nand U2729 (N_2729,N_2441,N_2080);
and U2730 (N_2730,N_2404,N_2064);
and U2731 (N_2731,N_2363,N_2029);
nor U2732 (N_2732,N_2430,N_2341);
and U2733 (N_2733,N_2183,N_2073);
or U2734 (N_2734,N_2084,N_2296);
and U2735 (N_2735,N_2244,N_2218);
and U2736 (N_2736,N_2129,N_2289);
nand U2737 (N_2737,N_2310,N_2121);
or U2738 (N_2738,N_2122,N_2038);
nor U2739 (N_2739,N_2424,N_2206);
and U2740 (N_2740,N_2280,N_2055);
xor U2741 (N_2741,N_2210,N_2350);
nand U2742 (N_2742,N_2088,N_2166);
and U2743 (N_2743,N_2466,N_2444);
and U2744 (N_2744,N_2225,N_2267);
nand U2745 (N_2745,N_2017,N_2264);
or U2746 (N_2746,N_2482,N_2456);
xnor U2747 (N_2747,N_2016,N_2174);
or U2748 (N_2748,N_2346,N_2293);
or U2749 (N_2749,N_2229,N_2109);
nor U2750 (N_2750,N_2166,N_2050);
nand U2751 (N_2751,N_2305,N_2352);
nor U2752 (N_2752,N_2036,N_2168);
nand U2753 (N_2753,N_2267,N_2104);
or U2754 (N_2754,N_2003,N_2172);
or U2755 (N_2755,N_2236,N_2437);
nor U2756 (N_2756,N_2490,N_2442);
xnor U2757 (N_2757,N_2214,N_2050);
nor U2758 (N_2758,N_2056,N_2126);
nor U2759 (N_2759,N_2418,N_2498);
nand U2760 (N_2760,N_2101,N_2441);
nor U2761 (N_2761,N_2390,N_2325);
nand U2762 (N_2762,N_2399,N_2186);
nand U2763 (N_2763,N_2385,N_2322);
nand U2764 (N_2764,N_2224,N_2147);
or U2765 (N_2765,N_2150,N_2131);
nand U2766 (N_2766,N_2143,N_2450);
nand U2767 (N_2767,N_2345,N_2098);
and U2768 (N_2768,N_2060,N_2486);
nor U2769 (N_2769,N_2191,N_2374);
nand U2770 (N_2770,N_2017,N_2040);
xor U2771 (N_2771,N_2331,N_2030);
nor U2772 (N_2772,N_2436,N_2328);
nor U2773 (N_2773,N_2294,N_2185);
and U2774 (N_2774,N_2260,N_2044);
nor U2775 (N_2775,N_2005,N_2222);
or U2776 (N_2776,N_2067,N_2064);
and U2777 (N_2777,N_2039,N_2248);
nor U2778 (N_2778,N_2281,N_2497);
or U2779 (N_2779,N_2495,N_2250);
or U2780 (N_2780,N_2038,N_2480);
or U2781 (N_2781,N_2155,N_2203);
and U2782 (N_2782,N_2105,N_2069);
xnor U2783 (N_2783,N_2110,N_2215);
nor U2784 (N_2784,N_2135,N_2351);
nor U2785 (N_2785,N_2382,N_2496);
and U2786 (N_2786,N_2422,N_2343);
xnor U2787 (N_2787,N_2356,N_2205);
nand U2788 (N_2788,N_2186,N_2488);
xnor U2789 (N_2789,N_2425,N_2232);
nor U2790 (N_2790,N_2220,N_2449);
and U2791 (N_2791,N_2453,N_2051);
nand U2792 (N_2792,N_2076,N_2448);
nand U2793 (N_2793,N_2068,N_2085);
nor U2794 (N_2794,N_2455,N_2201);
and U2795 (N_2795,N_2150,N_2367);
nor U2796 (N_2796,N_2463,N_2173);
nor U2797 (N_2797,N_2369,N_2030);
xnor U2798 (N_2798,N_2372,N_2168);
nand U2799 (N_2799,N_2484,N_2261);
nand U2800 (N_2800,N_2414,N_2327);
and U2801 (N_2801,N_2329,N_2206);
and U2802 (N_2802,N_2464,N_2243);
and U2803 (N_2803,N_2126,N_2332);
nor U2804 (N_2804,N_2081,N_2258);
xnor U2805 (N_2805,N_2444,N_2041);
nand U2806 (N_2806,N_2032,N_2165);
nand U2807 (N_2807,N_2161,N_2112);
nor U2808 (N_2808,N_2039,N_2075);
nor U2809 (N_2809,N_2331,N_2378);
or U2810 (N_2810,N_2178,N_2365);
or U2811 (N_2811,N_2486,N_2484);
nand U2812 (N_2812,N_2177,N_2374);
or U2813 (N_2813,N_2016,N_2401);
or U2814 (N_2814,N_2179,N_2081);
or U2815 (N_2815,N_2353,N_2309);
or U2816 (N_2816,N_2139,N_2115);
xor U2817 (N_2817,N_2484,N_2282);
nand U2818 (N_2818,N_2463,N_2200);
nand U2819 (N_2819,N_2051,N_2472);
nand U2820 (N_2820,N_2041,N_2285);
and U2821 (N_2821,N_2191,N_2248);
nor U2822 (N_2822,N_2369,N_2160);
nand U2823 (N_2823,N_2361,N_2149);
and U2824 (N_2824,N_2138,N_2276);
xnor U2825 (N_2825,N_2156,N_2018);
nand U2826 (N_2826,N_2277,N_2349);
xor U2827 (N_2827,N_2487,N_2145);
nand U2828 (N_2828,N_2367,N_2316);
xor U2829 (N_2829,N_2444,N_2072);
nor U2830 (N_2830,N_2282,N_2144);
nor U2831 (N_2831,N_2317,N_2451);
or U2832 (N_2832,N_2430,N_2426);
nand U2833 (N_2833,N_2346,N_2284);
nor U2834 (N_2834,N_2466,N_2315);
xnor U2835 (N_2835,N_2108,N_2424);
and U2836 (N_2836,N_2042,N_2212);
and U2837 (N_2837,N_2426,N_2110);
nor U2838 (N_2838,N_2096,N_2447);
xor U2839 (N_2839,N_2058,N_2218);
xnor U2840 (N_2840,N_2035,N_2049);
nand U2841 (N_2841,N_2494,N_2465);
nand U2842 (N_2842,N_2219,N_2184);
or U2843 (N_2843,N_2185,N_2012);
or U2844 (N_2844,N_2053,N_2251);
or U2845 (N_2845,N_2103,N_2027);
xor U2846 (N_2846,N_2240,N_2283);
or U2847 (N_2847,N_2051,N_2336);
or U2848 (N_2848,N_2379,N_2010);
xor U2849 (N_2849,N_2094,N_2120);
xnor U2850 (N_2850,N_2388,N_2477);
nand U2851 (N_2851,N_2160,N_2096);
or U2852 (N_2852,N_2352,N_2023);
or U2853 (N_2853,N_2403,N_2048);
or U2854 (N_2854,N_2116,N_2102);
xor U2855 (N_2855,N_2496,N_2309);
xor U2856 (N_2856,N_2488,N_2187);
nor U2857 (N_2857,N_2440,N_2173);
nor U2858 (N_2858,N_2342,N_2424);
or U2859 (N_2859,N_2315,N_2233);
and U2860 (N_2860,N_2130,N_2323);
and U2861 (N_2861,N_2281,N_2235);
xnor U2862 (N_2862,N_2469,N_2395);
and U2863 (N_2863,N_2196,N_2424);
and U2864 (N_2864,N_2347,N_2035);
xor U2865 (N_2865,N_2386,N_2129);
and U2866 (N_2866,N_2082,N_2117);
nor U2867 (N_2867,N_2241,N_2223);
nand U2868 (N_2868,N_2383,N_2234);
or U2869 (N_2869,N_2319,N_2048);
and U2870 (N_2870,N_2491,N_2449);
and U2871 (N_2871,N_2187,N_2408);
and U2872 (N_2872,N_2392,N_2139);
or U2873 (N_2873,N_2333,N_2435);
xnor U2874 (N_2874,N_2340,N_2276);
nand U2875 (N_2875,N_2294,N_2467);
nor U2876 (N_2876,N_2436,N_2455);
or U2877 (N_2877,N_2470,N_2300);
or U2878 (N_2878,N_2098,N_2234);
nor U2879 (N_2879,N_2031,N_2479);
xnor U2880 (N_2880,N_2308,N_2203);
and U2881 (N_2881,N_2253,N_2062);
nand U2882 (N_2882,N_2217,N_2054);
and U2883 (N_2883,N_2013,N_2078);
or U2884 (N_2884,N_2202,N_2149);
or U2885 (N_2885,N_2084,N_2150);
or U2886 (N_2886,N_2194,N_2356);
nor U2887 (N_2887,N_2455,N_2271);
and U2888 (N_2888,N_2172,N_2392);
nor U2889 (N_2889,N_2410,N_2440);
xor U2890 (N_2890,N_2161,N_2438);
or U2891 (N_2891,N_2293,N_2207);
nor U2892 (N_2892,N_2094,N_2208);
and U2893 (N_2893,N_2330,N_2177);
nor U2894 (N_2894,N_2373,N_2469);
or U2895 (N_2895,N_2462,N_2168);
and U2896 (N_2896,N_2020,N_2472);
xor U2897 (N_2897,N_2162,N_2449);
and U2898 (N_2898,N_2375,N_2352);
and U2899 (N_2899,N_2129,N_2293);
nand U2900 (N_2900,N_2361,N_2498);
or U2901 (N_2901,N_2498,N_2175);
nor U2902 (N_2902,N_2450,N_2087);
and U2903 (N_2903,N_2045,N_2246);
xnor U2904 (N_2904,N_2362,N_2063);
or U2905 (N_2905,N_2027,N_2390);
nor U2906 (N_2906,N_2273,N_2096);
nor U2907 (N_2907,N_2281,N_2093);
xor U2908 (N_2908,N_2148,N_2414);
nand U2909 (N_2909,N_2388,N_2413);
nand U2910 (N_2910,N_2090,N_2123);
nor U2911 (N_2911,N_2101,N_2489);
and U2912 (N_2912,N_2154,N_2202);
nor U2913 (N_2913,N_2095,N_2068);
or U2914 (N_2914,N_2485,N_2273);
xor U2915 (N_2915,N_2407,N_2470);
and U2916 (N_2916,N_2288,N_2200);
nor U2917 (N_2917,N_2121,N_2076);
nor U2918 (N_2918,N_2126,N_2128);
xor U2919 (N_2919,N_2270,N_2389);
nand U2920 (N_2920,N_2125,N_2276);
xnor U2921 (N_2921,N_2037,N_2330);
nand U2922 (N_2922,N_2184,N_2028);
and U2923 (N_2923,N_2354,N_2299);
and U2924 (N_2924,N_2020,N_2299);
nand U2925 (N_2925,N_2220,N_2450);
nand U2926 (N_2926,N_2467,N_2244);
xor U2927 (N_2927,N_2160,N_2436);
xnor U2928 (N_2928,N_2135,N_2231);
and U2929 (N_2929,N_2107,N_2440);
nor U2930 (N_2930,N_2279,N_2200);
xnor U2931 (N_2931,N_2491,N_2421);
or U2932 (N_2932,N_2272,N_2226);
nor U2933 (N_2933,N_2365,N_2043);
and U2934 (N_2934,N_2105,N_2171);
or U2935 (N_2935,N_2122,N_2493);
and U2936 (N_2936,N_2069,N_2236);
nand U2937 (N_2937,N_2120,N_2358);
and U2938 (N_2938,N_2316,N_2427);
xnor U2939 (N_2939,N_2218,N_2412);
and U2940 (N_2940,N_2141,N_2418);
xnor U2941 (N_2941,N_2239,N_2182);
or U2942 (N_2942,N_2461,N_2315);
nor U2943 (N_2943,N_2000,N_2320);
and U2944 (N_2944,N_2224,N_2413);
or U2945 (N_2945,N_2243,N_2303);
and U2946 (N_2946,N_2314,N_2352);
xnor U2947 (N_2947,N_2122,N_2466);
nand U2948 (N_2948,N_2071,N_2145);
nand U2949 (N_2949,N_2084,N_2129);
or U2950 (N_2950,N_2141,N_2001);
xnor U2951 (N_2951,N_2032,N_2040);
nor U2952 (N_2952,N_2396,N_2469);
or U2953 (N_2953,N_2379,N_2482);
and U2954 (N_2954,N_2473,N_2200);
or U2955 (N_2955,N_2041,N_2050);
nor U2956 (N_2956,N_2087,N_2157);
and U2957 (N_2957,N_2000,N_2067);
and U2958 (N_2958,N_2366,N_2495);
or U2959 (N_2959,N_2009,N_2017);
and U2960 (N_2960,N_2308,N_2372);
xnor U2961 (N_2961,N_2489,N_2243);
and U2962 (N_2962,N_2029,N_2275);
xnor U2963 (N_2963,N_2046,N_2017);
nand U2964 (N_2964,N_2291,N_2416);
and U2965 (N_2965,N_2301,N_2283);
xor U2966 (N_2966,N_2068,N_2267);
and U2967 (N_2967,N_2320,N_2449);
nand U2968 (N_2968,N_2258,N_2328);
and U2969 (N_2969,N_2281,N_2498);
and U2970 (N_2970,N_2000,N_2066);
xnor U2971 (N_2971,N_2175,N_2013);
nand U2972 (N_2972,N_2172,N_2150);
xor U2973 (N_2973,N_2193,N_2153);
or U2974 (N_2974,N_2409,N_2394);
and U2975 (N_2975,N_2495,N_2044);
nand U2976 (N_2976,N_2291,N_2324);
xnor U2977 (N_2977,N_2220,N_2455);
and U2978 (N_2978,N_2423,N_2477);
and U2979 (N_2979,N_2182,N_2240);
nor U2980 (N_2980,N_2083,N_2065);
or U2981 (N_2981,N_2118,N_2251);
nor U2982 (N_2982,N_2217,N_2246);
and U2983 (N_2983,N_2485,N_2193);
or U2984 (N_2984,N_2375,N_2378);
nor U2985 (N_2985,N_2026,N_2233);
xnor U2986 (N_2986,N_2264,N_2195);
xnor U2987 (N_2987,N_2282,N_2020);
or U2988 (N_2988,N_2066,N_2154);
nand U2989 (N_2989,N_2192,N_2031);
or U2990 (N_2990,N_2312,N_2072);
xor U2991 (N_2991,N_2094,N_2336);
and U2992 (N_2992,N_2116,N_2363);
and U2993 (N_2993,N_2065,N_2361);
xnor U2994 (N_2994,N_2490,N_2127);
or U2995 (N_2995,N_2073,N_2306);
xor U2996 (N_2996,N_2104,N_2220);
xor U2997 (N_2997,N_2028,N_2358);
and U2998 (N_2998,N_2214,N_2413);
nor U2999 (N_2999,N_2065,N_2304);
and U3000 (N_3000,N_2971,N_2874);
or U3001 (N_3001,N_2606,N_2886);
nand U3002 (N_3002,N_2529,N_2657);
and U3003 (N_3003,N_2982,N_2940);
and U3004 (N_3004,N_2770,N_2921);
and U3005 (N_3005,N_2740,N_2787);
nor U3006 (N_3006,N_2765,N_2648);
nor U3007 (N_3007,N_2711,N_2880);
and U3008 (N_3008,N_2684,N_2892);
xnor U3009 (N_3009,N_2650,N_2885);
nor U3010 (N_3010,N_2973,N_2852);
nor U3011 (N_3011,N_2777,N_2965);
nor U3012 (N_3012,N_2534,N_2881);
nand U3013 (N_3013,N_2978,N_2997);
xor U3014 (N_3014,N_2564,N_2794);
nor U3015 (N_3015,N_2535,N_2966);
and U3016 (N_3016,N_2867,N_2736);
and U3017 (N_3017,N_2757,N_2840);
and U3018 (N_3018,N_2907,N_2876);
xor U3019 (N_3019,N_2789,N_2592);
xnor U3020 (N_3020,N_2687,N_2561);
xnor U3021 (N_3021,N_2796,N_2584);
nand U3022 (N_3022,N_2912,N_2824);
xnor U3023 (N_3023,N_2663,N_2572);
xnor U3024 (N_3024,N_2926,N_2775);
nand U3025 (N_3025,N_2848,N_2567);
nand U3026 (N_3026,N_2888,N_2842);
or U3027 (N_3027,N_2990,N_2678);
nor U3028 (N_3028,N_2550,N_2516);
or U3029 (N_3029,N_2785,N_2944);
nor U3030 (N_3030,N_2506,N_2565);
xor U3031 (N_3031,N_2636,N_2836);
nor U3032 (N_3032,N_2622,N_2788);
nand U3033 (N_3033,N_2941,N_2672);
and U3034 (N_3034,N_2810,N_2715);
nand U3035 (N_3035,N_2823,N_2862);
xor U3036 (N_3036,N_2820,N_2799);
nor U3037 (N_3037,N_2590,N_2625);
and U3038 (N_3038,N_2955,N_2919);
xnor U3039 (N_3039,N_2679,N_2859);
or U3040 (N_3040,N_2682,N_2968);
xnor U3041 (N_3041,N_2598,N_2922);
or U3042 (N_3042,N_2509,N_2538);
and U3043 (N_3043,N_2868,N_2675);
and U3044 (N_3044,N_2952,N_2722);
or U3045 (N_3045,N_2994,N_2716);
or U3046 (N_3046,N_2644,N_2605);
nand U3047 (N_3047,N_2897,N_2658);
nand U3048 (N_3048,N_2557,N_2809);
xor U3049 (N_3049,N_2714,N_2577);
xor U3050 (N_3050,N_2913,N_2642);
or U3051 (N_3051,N_2596,N_2668);
nor U3052 (N_3052,N_2967,N_2523);
xor U3053 (N_3053,N_2974,N_2957);
xor U3054 (N_3054,N_2582,N_2615);
nand U3055 (N_3055,N_2815,N_2917);
xor U3056 (N_3056,N_2635,N_2960);
or U3057 (N_3057,N_2838,N_2681);
nor U3058 (N_3058,N_2540,N_2560);
nand U3059 (N_3059,N_2725,N_2959);
or U3060 (N_3060,N_2520,N_2686);
xor U3061 (N_3061,N_2786,N_2549);
xor U3062 (N_3062,N_2833,N_2539);
nand U3063 (N_3063,N_2846,N_2805);
nor U3064 (N_3064,N_2694,N_2619);
nor U3065 (N_3065,N_2710,N_2993);
nor U3066 (N_3066,N_2507,N_2871);
nand U3067 (N_3067,N_2814,N_2578);
and U3068 (N_3068,N_2847,N_2901);
nand U3069 (N_3069,N_2975,N_2697);
nor U3070 (N_3070,N_2843,N_2515);
xnor U3071 (N_3071,N_2562,N_2500);
nand U3072 (N_3072,N_2626,N_2837);
nor U3073 (N_3073,N_2870,N_2734);
or U3074 (N_3074,N_2612,N_2904);
nor U3075 (N_3075,N_2841,N_2728);
nand U3076 (N_3076,N_2915,N_2695);
and U3077 (N_3077,N_2743,N_2653);
nor U3078 (N_3078,N_2513,N_2646);
or U3079 (N_3079,N_2649,N_2522);
or U3080 (N_3080,N_2989,N_2717);
xor U3081 (N_3081,N_2637,N_2568);
or U3082 (N_3082,N_2772,N_2898);
xor U3083 (N_3083,N_2700,N_2832);
xnor U3084 (N_3084,N_2835,N_2660);
nor U3085 (N_3085,N_2609,N_2571);
xor U3086 (N_3086,N_2961,N_2517);
and U3087 (N_3087,N_2603,N_2748);
or U3088 (N_3088,N_2807,N_2712);
xor U3089 (N_3089,N_2827,N_2858);
and U3090 (N_3090,N_2632,N_2692);
nor U3091 (N_3091,N_2614,N_2911);
or U3092 (N_3092,N_2895,N_2667);
nor U3093 (N_3093,N_2942,N_2768);
xnor U3094 (N_3094,N_2766,N_2864);
xor U3095 (N_3095,N_2747,N_2671);
xor U3096 (N_3096,N_2834,N_2970);
xor U3097 (N_3097,N_2628,N_2875);
and U3098 (N_3098,N_2845,N_2738);
and U3099 (N_3099,N_2878,N_2854);
nor U3100 (N_3100,N_2666,N_2899);
and U3101 (N_3101,N_2776,N_2623);
xor U3102 (N_3102,N_2928,N_2977);
xor U3103 (N_3103,N_2593,N_2599);
nand U3104 (N_3104,N_2633,N_2784);
nand U3105 (N_3105,N_2797,N_2631);
and U3106 (N_3106,N_2643,N_2532);
nand U3107 (N_3107,N_2719,N_2869);
xnor U3108 (N_3108,N_2691,N_2662);
nand U3109 (N_3109,N_2951,N_2709);
xnor U3110 (N_3110,N_2983,N_2801);
and U3111 (N_3111,N_2587,N_2718);
nor U3112 (N_3112,N_2872,N_2791);
nand U3113 (N_3113,N_2894,N_2808);
or U3114 (N_3114,N_2893,N_2616);
or U3115 (N_3115,N_2783,N_2986);
xnor U3116 (N_3116,N_2943,N_2987);
or U3117 (N_3117,N_2689,N_2769);
xor U3118 (N_3118,N_2927,N_2849);
and U3119 (N_3119,N_2802,N_2767);
xor U3120 (N_3120,N_2621,N_2936);
nand U3121 (N_3121,N_2591,N_2905);
nand U3122 (N_3122,N_2713,N_2638);
xnor U3123 (N_3123,N_2884,N_2857);
and U3124 (N_3124,N_2762,N_2937);
xor U3125 (N_3125,N_2699,N_2601);
and U3126 (N_3126,N_2861,N_2580);
nand U3127 (N_3127,N_2761,N_2627);
and U3128 (N_3128,N_2879,N_2720);
and U3129 (N_3129,N_2558,N_2798);
xor U3130 (N_3130,N_2831,N_2505);
nand U3131 (N_3131,N_2597,N_2524);
nand U3132 (N_3132,N_2737,N_2556);
nand U3133 (N_3133,N_2702,N_2931);
nor U3134 (N_3134,N_2502,N_2803);
and U3135 (N_3135,N_2563,N_2526);
and U3136 (N_3136,N_2726,N_2521);
nor U3137 (N_3137,N_2826,N_2611);
nand U3138 (N_3138,N_2948,N_2533);
nand U3139 (N_3139,N_2721,N_2552);
nand U3140 (N_3140,N_2906,N_2882);
nand U3141 (N_3141,N_2669,N_2602);
nand U3142 (N_3142,N_2963,N_2690);
nor U3143 (N_3143,N_2503,N_2555);
xor U3144 (N_3144,N_2839,N_2877);
xnor U3145 (N_3145,N_2610,N_2519);
xnor U3146 (N_3146,N_2673,N_2964);
nand U3147 (N_3147,N_2929,N_2760);
or U3148 (N_3148,N_2908,N_2569);
or U3149 (N_3149,N_2751,N_2756);
nand U3150 (N_3150,N_2918,N_2741);
nor U3151 (N_3151,N_2570,N_2817);
or U3152 (N_3152,N_2950,N_2510);
nor U3153 (N_3153,N_2991,N_2607);
nor U3154 (N_3154,N_2508,N_2739);
xnor U3155 (N_3155,N_2780,N_2903);
nor U3156 (N_3156,N_2980,N_2851);
and U3157 (N_3157,N_2932,N_2822);
or U3158 (N_3158,N_2956,N_2630);
nor U3159 (N_3159,N_2850,N_2958);
nand U3160 (N_3160,N_2579,N_2863);
nor U3161 (N_3161,N_2909,N_2828);
nand U3162 (N_3162,N_2693,N_2812);
nor U3163 (N_3163,N_2962,N_2703);
and U3164 (N_3164,N_2543,N_2585);
nand U3165 (N_3165,N_2853,N_2883);
xor U3166 (N_3166,N_2742,N_2652);
nand U3167 (N_3167,N_2920,N_2573);
or U3168 (N_3168,N_2856,N_2764);
xnor U3169 (N_3169,N_2589,N_2800);
nand U3170 (N_3170,N_2542,N_2536);
or U3171 (N_3171,N_2661,N_2685);
and U3172 (N_3172,N_2745,N_2530);
or U3173 (N_3173,N_2654,N_2746);
and U3174 (N_3174,N_2995,N_2758);
and U3175 (N_3175,N_2581,N_2825);
and U3176 (N_3176,N_2954,N_2829);
nand U3177 (N_3177,N_2795,N_2647);
or U3178 (N_3178,N_2566,N_2525);
xnor U3179 (N_3179,N_2866,N_2934);
xnor U3180 (N_3180,N_2900,N_2511);
nand U3181 (N_3181,N_2945,N_2811);
and U3182 (N_3182,N_2890,N_2860);
xor U3183 (N_3183,N_2735,N_2501);
or U3184 (N_3184,N_2541,N_2939);
nand U3185 (N_3185,N_2670,N_2781);
or U3186 (N_3186,N_2586,N_2916);
and U3187 (N_3187,N_2792,N_2553);
or U3188 (N_3188,N_2656,N_2819);
nand U3189 (N_3189,N_2608,N_2664);
or U3190 (N_3190,N_2773,N_2655);
xor U3191 (N_3191,N_2724,N_2574);
or U3192 (N_3192,N_2680,N_2696);
or U3193 (N_3193,N_2755,N_2708);
and U3194 (N_3194,N_2759,N_2730);
and U3195 (N_3195,N_2969,N_2984);
nor U3196 (N_3196,N_2545,N_2996);
and U3197 (N_3197,N_2749,N_2999);
or U3198 (N_3198,N_2620,N_2544);
nor U3199 (N_3199,N_2947,N_2548);
xor U3200 (N_3200,N_2729,N_2816);
and U3201 (N_3201,N_2546,N_2683);
and U3202 (N_3202,N_2813,N_2972);
nor U3203 (N_3203,N_2778,N_2732);
nand U3204 (N_3204,N_2651,N_2504);
xor U3205 (N_3205,N_2583,N_2855);
or U3206 (N_3206,N_2528,N_2576);
or U3207 (N_3207,N_2537,N_2613);
xnor U3208 (N_3208,N_2518,N_2998);
nand U3209 (N_3209,N_2705,N_2896);
nor U3210 (N_3210,N_2688,N_2806);
xnor U3211 (N_3211,N_2992,N_2873);
nor U3212 (N_3212,N_2559,N_2804);
or U3213 (N_3213,N_2514,N_2731);
xor U3214 (N_3214,N_2782,N_2793);
xor U3215 (N_3215,N_2698,N_2930);
nor U3216 (N_3216,N_2641,N_2531);
nand U3217 (N_3217,N_2645,N_2551);
and U3218 (N_3218,N_2985,N_2924);
nor U3219 (N_3219,N_2818,N_2910);
and U3220 (N_3220,N_2923,N_2704);
nand U3221 (N_3221,N_2887,N_2865);
nand U3222 (N_3222,N_2595,N_2844);
xnor U3223 (N_3223,N_2723,N_2588);
nand U3224 (N_3224,N_2981,N_2727);
and U3225 (N_3225,N_2665,N_2953);
and U3226 (N_3226,N_2790,N_2659);
or U3227 (N_3227,N_2639,N_2754);
and U3228 (N_3228,N_2527,N_2779);
xnor U3229 (N_3229,N_2594,N_2706);
or U3230 (N_3230,N_2547,N_2676);
nand U3231 (N_3231,N_2707,N_2830);
nand U3232 (N_3232,N_2624,N_2925);
nand U3233 (N_3233,N_2617,N_2750);
or U3234 (N_3234,N_2938,N_2744);
and U3235 (N_3235,N_2677,N_2774);
xnor U3236 (N_3236,N_2701,N_2604);
nor U3237 (N_3237,N_2575,N_2600);
and U3238 (N_3238,N_2988,N_2821);
and U3239 (N_3239,N_2902,N_2634);
and U3240 (N_3240,N_2771,N_2891);
nand U3241 (N_3241,N_2976,N_2512);
and U3242 (N_3242,N_2554,N_2763);
xnor U3243 (N_3243,N_2752,N_2733);
nor U3244 (N_3244,N_2935,N_2753);
nor U3245 (N_3245,N_2640,N_2946);
or U3246 (N_3246,N_2674,N_2914);
nand U3247 (N_3247,N_2949,N_2979);
nand U3248 (N_3248,N_2629,N_2889);
xnor U3249 (N_3249,N_2933,N_2618);
nor U3250 (N_3250,N_2723,N_2863);
nand U3251 (N_3251,N_2724,N_2810);
and U3252 (N_3252,N_2827,N_2739);
nand U3253 (N_3253,N_2961,N_2625);
xnor U3254 (N_3254,N_2745,N_2901);
nor U3255 (N_3255,N_2651,N_2801);
nor U3256 (N_3256,N_2579,N_2613);
xor U3257 (N_3257,N_2926,N_2618);
xor U3258 (N_3258,N_2983,N_2941);
xnor U3259 (N_3259,N_2867,N_2684);
and U3260 (N_3260,N_2604,N_2613);
nor U3261 (N_3261,N_2938,N_2917);
nor U3262 (N_3262,N_2702,N_2863);
xnor U3263 (N_3263,N_2893,N_2888);
nor U3264 (N_3264,N_2804,N_2898);
xnor U3265 (N_3265,N_2608,N_2920);
and U3266 (N_3266,N_2783,N_2887);
nor U3267 (N_3267,N_2656,N_2519);
or U3268 (N_3268,N_2735,N_2708);
nand U3269 (N_3269,N_2880,N_2888);
or U3270 (N_3270,N_2897,N_2885);
and U3271 (N_3271,N_2863,N_2714);
and U3272 (N_3272,N_2588,N_2911);
or U3273 (N_3273,N_2533,N_2933);
nand U3274 (N_3274,N_2919,N_2806);
nand U3275 (N_3275,N_2537,N_2705);
or U3276 (N_3276,N_2683,N_2742);
and U3277 (N_3277,N_2711,N_2773);
and U3278 (N_3278,N_2544,N_2974);
xnor U3279 (N_3279,N_2629,N_2639);
nor U3280 (N_3280,N_2923,N_2588);
xor U3281 (N_3281,N_2969,N_2595);
nand U3282 (N_3282,N_2648,N_2581);
and U3283 (N_3283,N_2873,N_2887);
and U3284 (N_3284,N_2579,N_2966);
xnor U3285 (N_3285,N_2749,N_2701);
xnor U3286 (N_3286,N_2964,N_2728);
and U3287 (N_3287,N_2511,N_2623);
and U3288 (N_3288,N_2646,N_2742);
xnor U3289 (N_3289,N_2746,N_2954);
nand U3290 (N_3290,N_2604,N_2562);
nor U3291 (N_3291,N_2837,N_2972);
nand U3292 (N_3292,N_2752,N_2940);
and U3293 (N_3293,N_2829,N_2939);
and U3294 (N_3294,N_2574,N_2762);
and U3295 (N_3295,N_2715,N_2603);
nand U3296 (N_3296,N_2523,N_2621);
nand U3297 (N_3297,N_2890,N_2768);
or U3298 (N_3298,N_2608,N_2590);
or U3299 (N_3299,N_2724,N_2576);
xnor U3300 (N_3300,N_2834,N_2909);
and U3301 (N_3301,N_2657,N_2938);
and U3302 (N_3302,N_2594,N_2891);
nor U3303 (N_3303,N_2762,N_2585);
nor U3304 (N_3304,N_2750,N_2889);
or U3305 (N_3305,N_2928,N_2597);
and U3306 (N_3306,N_2889,N_2524);
nand U3307 (N_3307,N_2612,N_2950);
xor U3308 (N_3308,N_2980,N_2753);
or U3309 (N_3309,N_2628,N_2594);
xor U3310 (N_3310,N_2817,N_2811);
or U3311 (N_3311,N_2952,N_2592);
and U3312 (N_3312,N_2569,N_2983);
nand U3313 (N_3313,N_2826,N_2659);
and U3314 (N_3314,N_2551,N_2859);
nor U3315 (N_3315,N_2662,N_2539);
nor U3316 (N_3316,N_2760,N_2774);
xnor U3317 (N_3317,N_2868,N_2567);
or U3318 (N_3318,N_2565,N_2664);
nand U3319 (N_3319,N_2559,N_2516);
nand U3320 (N_3320,N_2673,N_2597);
xor U3321 (N_3321,N_2636,N_2592);
nand U3322 (N_3322,N_2687,N_2511);
nor U3323 (N_3323,N_2532,N_2522);
xor U3324 (N_3324,N_2634,N_2751);
or U3325 (N_3325,N_2930,N_2573);
nand U3326 (N_3326,N_2844,N_2539);
and U3327 (N_3327,N_2637,N_2611);
nor U3328 (N_3328,N_2526,N_2737);
nand U3329 (N_3329,N_2568,N_2583);
or U3330 (N_3330,N_2747,N_2716);
xor U3331 (N_3331,N_2522,N_2755);
or U3332 (N_3332,N_2732,N_2631);
xor U3333 (N_3333,N_2844,N_2559);
or U3334 (N_3334,N_2550,N_2895);
or U3335 (N_3335,N_2927,N_2741);
xor U3336 (N_3336,N_2698,N_2685);
xnor U3337 (N_3337,N_2660,N_2554);
xor U3338 (N_3338,N_2894,N_2500);
nand U3339 (N_3339,N_2890,N_2553);
xnor U3340 (N_3340,N_2602,N_2659);
or U3341 (N_3341,N_2713,N_2512);
nand U3342 (N_3342,N_2739,N_2690);
nor U3343 (N_3343,N_2889,N_2936);
nand U3344 (N_3344,N_2617,N_2598);
and U3345 (N_3345,N_2823,N_2608);
and U3346 (N_3346,N_2680,N_2646);
or U3347 (N_3347,N_2691,N_2868);
and U3348 (N_3348,N_2931,N_2893);
xor U3349 (N_3349,N_2653,N_2654);
xor U3350 (N_3350,N_2559,N_2619);
and U3351 (N_3351,N_2911,N_2730);
or U3352 (N_3352,N_2982,N_2528);
nand U3353 (N_3353,N_2990,N_2701);
or U3354 (N_3354,N_2535,N_2510);
nor U3355 (N_3355,N_2543,N_2643);
nor U3356 (N_3356,N_2933,N_2834);
nor U3357 (N_3357,N_2543,N_2619);
and U3358 (N_3358,N_2797,N_2520);
nand U3359 (N_3359,N_2958,N_2928);
and U3360 (N_3360,N_2664,N_2680);
and U3361 (N_3361,N_2584,N_2576);
or U3362 (N_3362,N_2857,N_2905);
and U3363 (N_3363,N_2920,N_2646);
or U3364 (N_3364,N_2504,N_2623);
nand U3365 (N_3365,N_2505,N_2752);
nand U3366 (N_3366,N_2743,N_2635);
nor U3367 (N_3367,N_2987,N_2728);
nand U3368 (N_3368,N_2742,N_2559);
xor U3369 (N_3369,N_2661,N_2779);
or U3370 (N_3370,N_2882,N_2978);
nand U3371 (N_3371,N_2844,N_2561);
or U3372 (N_3372,N_2846,N_2706);
nor U3373 (N_3373,N_2700,N_2648);
and U3374 (N_3374,N_2558,N_2761);
and U3375 (N_3375,N_2828,N_2984);
or U3376 (N_3376,N_2736,N_2957);
and U3377 (N_3377,N_2937,N_2638);
and U3378 (N_3378,N_2708,N_2505);
and U3379 (N_3379,N_2704,N_2872);
or U3380 (N_3380,N_2896,N_2683);
nor U3381 (N_3381,N_2883,N_2620);
nor U3382 (N_3382,N_2868,N_2805);
or U3383 (N_3383,N_2689,N_2852);
nand U3384 (N_3384,N_2843,N_2757);
nor U3385 (N_3385,N_2932,N_2754);
nand U3386 (N_3386,N_2752,N_2802);
xnor U3387 (N_3387,N_2512,N_2525);
or U3388 (N_3388,N_2922,N_2835);
nand U3389 (N_3389,N_2775,N_2690);
or U3390 (N_3390,N_2999,N_2539);
nand U3391 (N_3391,N_2685,N_2824);
or U3392 (N_3392,N_2687,N_2951);
and U3393 (N_3393,N_2886,N_2723);
and U3394 (N_3394,N_2853,N_2994);
xnor U3395 (N_3395,N_2837,N_2720);
xnor U3396 (N_3396,N_2814,N_2673);
nor U3397 (N_3397,N_2633,N_2928);
or U3398 (N_3398,N_2919,N_2634);
nor U3399 (N_3399,N_2849,N_2635);
nor U3400 (N_3400,N_2826,N_2873);
and U3401 (N_3401,N_2515,N_2542);
and U3402 (N_3402,N_2589,N_2622);
nand U3403 (N_3403,N_2732,N_2877);
or U3404 (N_3404,N_2669,N_2972);
or U3405 (N_3405,N_2696,N_2532);
xnor U3406 (N_3406,N_2642,N_2688);
xnor U3407 (N_3407,N_2647,N_2540);
nand U3408 (N_3408,N_2975,N_2873);
nor U3409 (N_3409,N_2647,N_2544);
xnor U3410 (N_3410,N_2802,N_2760);
nand U3411 (N_3411,N_2528,N_2580);
xor U3412 (N_3412,N_2771,N_2797);
nand U3413 (N_3413,N_2969,N_2806);
and U3414 (N_3414,N_2588,N_2522);
or U3415 (N_3415,N_2591,N_2703);
nor U3416 (N_3416,N_2869,N_2990);
nand U3417 (N_3417,N_2835,N_2808);
or U3418 (N_3418,N_2924,N_2977);
or U3419 (N_3419,N_2545,N_2700);
or U3420 (N_3420,N_2767,N_2523);
and U3421 (N_3421,N_2913,N_2676);
xor U3422 (N_3422,N_2935,N_2963);
and U3423 (N_3423,N_2825,N_2679);
nor U3424 (N_3424,N_2747,N_2885);
xor U3425 (N_3425,N_2932,N_2555);
xor U3426 (N_3426,N_2968,N_2969);
or U3427 (N_3427,N_2882,N_2792);
and U3428 (N_3428,N_2739,N_2560);
and U3429 (N_3429,N_2633,N_2996);
nand U3430 (N_3430,N_2822,N_2769);
xor U3431 (N_3431,N_2626,N_2594);
and U3432 (N_3432,N_2874,N_2598);
or U3433 (N_3433,N_2781,N_2696);
xor U3434 (N_3434,N_2953,N_2961);
nand U3435 (N_3435,N_2914,N_2677);
nand U3436 (N_3436,N_2762,N_2809);
and U3437 (N_3437,N_2517,N_2644);
nand U3438 (N_3438,N_2551,N_2526);
nor U3439 (N_3439,N_2893,N_2973);
nor U3440 (N_3440,N_2517,N_2525);
nor U3441 (N_3441,N_2509,N_2950);
and U3442 (N_3442,N_2623,N_2676);
xnor U3443 (N_3443,N_2799,N_2667);
and U3444 (N_3444,N_2596,N_2557);
xor U3445 (N_3445,N_2618,N_2617);
nor U3446 (N_3446,N_2854,N_2764);
or U3447 (N_3447,N_2761,N_2805);
nand U3448 (N_3448,N_2951,N_2506);
or U3449 (N_3449,N_2695,N_2899);
or U3450 (N_3450,N_2740,N_2691);
nand U3451 (N_3451,N_2596,N_2904);
nor U3452 (N_3452,N_2561,N_2821);
xnor U3453 (N_3453,N_2597,N_2969);
or U3454 (N_3454,N_2641,N_2571);
xor U3455 (N_3455,N_2742,N_2772);
or U3456 (N_3456,N_2940,N_2634);
nor U3457 (N_3457,N_2977,N_2966);
xor U3458 (N_3458,N_2701,N_2774);
and U3459 (N_3459,N_2766,N_2820);
nor U3460 (N_3460,N_2650,N_2605);
and U3461 (N_3461,N_2550,N_2648);
or U3462 (N_3462,N_2777,N_2500);
nand U3463 (N_3463,N_2609,N_2826);
nor U3464 (N_3464,N_2507,N_2670);
nor U3465 (N_3465,N_2592,N_2860);
nand U3466 (N_3466,N_2601,N_2514);
or U3467 (N_3467,N_2911,N_2668);
nand U3468 (N_3468,N_2800,N_2543);
or U3469 (N_3469,N_2682,N_2846);
nor U3470 (N_3470,N_2607,N_2926);
and U3471 (N_3471,N_2886,N_2724);
nor U3472 (N_3472,N_2759,N_2645);
xor U3473 (N_3473,N_2657,N_2507);
nor U3474 (N_3474,N_2974,N_2712);
nand U3475 (N_3475,N_2573,N_2751);
xnor U3476 (N_3476,N_2630,N_2880);
or U3477 (N_3477,N_2962,N_2723);
nand U3478 (N_3478,N_2935,N_2508);
and U3479 (N_3479,N_2566,N_2540);
nor U3480 (N_3480,N_2891,N_2719);
nor U3481 (N_3481,N_2860,N_2889);
and U3482 (N_3482,N_2848,N_2898);
or U3483 (N_3483,N_2713,N_2966);
xor U3484 (N_3484,N_2514,N_2827);
nor U3485 (N_3485,N_2527,N_2847);
or U3486 (N_3486,N_2796,N_2985);
or U3487 (N_3487,N_2637,N_2955);
nand U3488 (N_3488,N_2765,N_2558);
xnor U3489 (N_3489,N_2968,N_2828);
and U3490 (N_3490,N_2812,N_2888);
or U3491 (N_3491,N_2911,N_2754);
nand U3492 (N_3492,N_2622,N_2590);
and U3493 (N_3493,N_2556,N_2791);
nand U3494 (N_3494,N_2670,N_2934);
nand U3495 (N_3495,N_2773,N_2630);
xor U3496 (N_3496,N_2802,N_2669);
nor U3497 (N_3497,N_2689,N_2911);
nor U3498 (N_3498,N_2785,N_2778);
or U3499 (N_3499,N_2968,N_2854);
and U3500 (N_3500,N_3159,N_3233);
and U3501 (N_3501,N_3196,N_3395);
nor U3502 (N_3502,N_3062,N_3108);
nand U3503 (N_3503,N_3273,N_3322);
and U3504 (N_3504,N_3317,N_3275);
and U3505 (N_3505,N_3231,N_3292);
or U3506 (N_3506,N_3099,N_3149);
nor U3507 (N_3507,N_3369,N_3312);
nor U3508 (N_3508,N_3213,N_3324);
nor U3509 (N_3509,N_3125,N_3359);
and U3510 (N_3510,N_3335,N_3470);
and U3511 (N_3511,N_3022,N_3490);
nand U3512 (N_3512,N_3461,N_3462);
or U3513 (N_3513,N_3091,N_3449);
and U3514 (N_3514,N_3259,N_3001);
xor U3515 (N_3515,N_3241,N_3323);
or U3516 (N_3516,N_3178,N_3267);
nand U3517 (N_3517,N_3129,N_3372);
xor U3518 (N_3518,N_3043,N_3058);
xnor U3519 (N_3519,N_3230,N_3309);
and U3520 (N_3520,N_3409,N_3176);
nand U3521 (N_3521,N_3009,N_3417);
or U3522 (N_3522,N_3356,N_3250);
nand U3523 (N_3523,N_3036,N_3383);
nor U3524 (N_3524,N_3332,N_3475);
nand U3525 (N_3525,N_3430,N_3158);
or U3526 (N_3526,N_3450,N_3177);
xnor U3527 (N_3527,N_3445,N_3459);
xor U3528 (N_3528,N_3366,N_3494);
nand U3529 (N_3529,N_3018,N_3133);
or U3530 (N_3530,N_3113,N_3377);
or U3531 (N_3531,N_3346,N_3368);
or U3532 (N_3532,N_3466,N_3394);
or U3533 (N_3533,N_3270,N_3287);
nand U3534 (N_3534,N_3402,N_3049);
and U3535 (N_3535,N_3362,N_3135);
or U3536 (N_3536,N_3358,N_3418);
xnor U3537 (N_3537,N_3334,N_3225);
and U3538 (N_3538,N_3126,N_3115);
nand U3539 (N_3539,N_3077,N_3281);
xor U3540 (N_3540,N_3298,N_3145);
or U3541 (N_3541,N_3151,N_3226);
and U3542 (N_3542,N_3097,N_3232);
nor U3543 (N_3543,N_3416,N_3160);
nand U3544 (N_3544,N_3191,N_3382);
nor U3545 (N_3545,N_3146,N_3215);
and U3546 (N_3546,N_3085,N_3199);
xor U3547 (N_3547,N_3396,N_3123);
nor U3548 (N_3548,N_3350,N_3139);
nor U3549 (N_3549,N_3076,N_3200);
nor U3550 (N_3550,N_3423,N_3235);
or U3551 (N_3551,N_3119,N_3031);
nand U3552 (N_3552,N_3472,N_3051);
and U3553 (N_3553,N_3063,N_3242);
nand U3554 (N_3554,N_3238,N_3035);
nand U3555 (N_3555,N_3040,N_3329);
xnor U3556 (N_3556,N_3157,N_3258);
nor U3557 (N_3557,N_3069,N_3061);
nor U3558 (N_3558,N_3384,N_3353);
nand U3559 (N_3559,N_3081,N_3072);
nor U3560 (N_3560,N_3143,N_3240);
or U3561 (N_3561,N_3337,N_3015);
and U3562 (N_3562,N_3385,N_3060);
and U3563 (N_3563,N_3348,N_3279);
xor U3564 (N_3564,N_3357,N_3165);
xnor U3565 (N_3565,N_3310,N_3419);
and U3566 (N_3566,N_3024,N_3016);
or U3567 (N_3567,N_3155,N_3308);
or U3568 (N_3568,N_3217,N_3412);
nand U3569 (N_3569,N_3020,N_3276);
and U3570 (N_3570,N_3255,N_3150);
or U3571 (N_3571,N_3488,N_3278);
nand U3572 (N_3572,N_3048,N_3340);
or U3573 (N_3573,N_3437,N_3166);
or U3574 (N_3574,N_3065,N_3447);
nand U3575 (N_3575,N_3074,N_3026);
nor U3576 (N_3576,N_3127,N_3376);
or U3577 (N_3577,N_3465,N_3037);
nand U3578 (N_3578,N_3254,N_3451);
nand U3579 (N_3579,N_3138,N_3087);
and U3580 (N_3580,N_3304,N_3364);
or U3581 (N_3581,N_3011,N_3136);
nand U3582 (N_3582,N_3397,N_3390);
xnor U3583 (N_3583,N_3244,N_3468);
xor U3584 (N_3584,N_3429,N_3311);
nand U3585 (N_3585,N_3030,N_3482);
or U3586 (N_3586,N_3454,N_3438);
nand U3587 (N_3587,N_3425,N_3131);
xor U3588 (N_3588,N_3361,N_3209);
and U3589 (N_3589,N_3453,N_3455);
xnor U3590 (N_3590,N_3010,N_3476);
nor U3591 (N_3591,N_3406,N_3251);
and U3592 (N_3592,N_3027,N_3245);
nand U3593 (N_3593,N_3321,N_3021);
nand U3594 (N_3594,N_3497,N_3189);
or U3595 (N_3595,N_3260,N_3073);
xnor U3596 (N_3596,N_3354,N_3435);
or U3597 (N_3597,N_3486,N_3389);
nand U3598 (N_3598,N_3089,N_3103);
nand U3599 (N_3599,N_3094,N_3263);
or U3600 (N_3600,N_3173,N_3481);
xor U3601 (N_3601,N_3344,N_3285);
and U3602 (N_3602,N_3100,N_3485);
nor U3603 (N_3603,N_3047,N_3201);
nand U3604 (N_3604,N_3112,N_3056);
nor U3605 (N_3605,N_3380,N_3493);
xor U3606 (N_3606,N_3474,N_3274);
and U3607 (N_3607,N_3243,N_3228);
or U3608 (N_3608,N_3296,N_3197);
xor U3609 (N_3609,N_3104,N_3339);
xnor U3610 (N_3610,N_3118,N_3148);
nand U3611 (N_3611,N_3247,N_3294);
nor U3612 (N_3612,N_3156,N_3163);
nand U3613 (N_3613,N_3443,N_3489);
nor U3614 (N_3614,N_3144,N_3008);
or U3615 (N_3615,N_3052,N_3257);
nand U3616 (N_3616,N_3034,N_3130);
xnor U3617 (N_3617,N_3019,N_3479);
or U3618 (N_3618,N_3162,N_3224);
xor U3619 (N_3619,N_3044,N_3183);
or U3620 (N_3620,N_3401,N_3253);
nand U3621 (N_3621,N_3057,N_3439);
nand U3622 (N_3622,N_3208,N_3411);
or U3623 (N_3623,N_3404,N_3261);
xnor U3624 (N_3624,N_3068,N_3315);
and U3625 (N_3625,N_3038,N_3484);
or U3626 (N_3626,N_3137,N_3473);
or U3627 (N_3627,N_3387,N_3110);
nand U3628 (N_3628,N_3098,N_3088);
nor U3629 (N_3629,N_3050,N_3070);
nor U3630 (N_3630,N_3202,N_3181);
and U3631 (N_3631,N_3326,N_3117);
or U3632 (N_3632,N_3028,N_3206);
and U3633 (N_3633,N_3442,N_3054);
xor U3634 (N_3634,N_3420,N_3071);
nand U3635 (N_3635,N_3268,N_3182);
xnor U3636 (N_3636,N_3121,N_3288);
nor U3637 (N_3637,N_3345,N_3082);
and U3638 (N_3638,N_3154,N_3105);
nor U3639 (N_3639,N_3301,N_3469);
and U3640 (N_3640,N_3046,N_3114);
nand U3641 (N_3641,N_3053,N_3391);
and U3642 (N_3642,N_3214,N_3014);
nand U3643 (N_3643,N_3471,N_3079);
nor U3644 (N_3644,N_3033,N_3271);
nand U3645 (N_3645,N_3295,N_3341);
xnor U3646 (N_3646,N_3055,N_3107);
and U3647 (N_3647,N_3192,N_3167);
and U3648 (N_3648,N_3306,N_3371);
and U3649 (N_3649,N_3221,N_3421);
and U3650 (N_3650,N_3313,N_3205);
nor U3651 (N_3651,N_3381,N_3092);
or U3652 (N_3652,N_3239,N_3360);
and U3653 (N_3653,N_3378,N_3218);
or U3654 (N_3654,N_3483,N_3161);
and U3655 (N_3655,N_3075,N_3370);
nor U3656 (N_3656,N_3272,N_3477);
or U3657 (N_3657,N_3175,N_3349);
or U3658 (N_3658,N_3480,N_3499);
xor U3659 (N_3659,N_3080,N_3227);
and U3660 (N_3660,N_3399,N_3492);
nand U3661 (N_3661,N_3219,N_3203);
or U3662 (N_3662,N_3180,N_3194);
xor U3663 (N_3663,N_3106,N_3434);
or U3664 (N_3664,N_3210,N_3000);
and U3665 (N_3665,N_3463,N_3005);
nand U3666 (N_3666,N_3122,N_3365);
and U3667 (N_3667,N_3414,N_3086);
and U3668 (N_3668,N_3456,N_3211);
nor U3669 (N_3669,N_3032,N_3336);
nand U3670 (N_3670,N_3084,N_3460);
nor U3671 (N_3671,N_3169,N_3207);
xor U3672 (N_3672,N_3045,N_3286);
nand U3673 (N_3673,N_3327,N_3299);
or U3674 (N_3674,N_3029,N_3140);
nor U3675 (N_3675,N_3120,N_3374);
or U3676 (N_3676,N_3342,N_3023);
and U3677 (N_3677,N_3152,N_3393);
nand U3678 (N_3678,N_3164,N_3495);
nor U3679 (N_3679,N_3293,N_3059);
nor U3680 (N_3680,N_3006,N_3067);
nand U3681 (N_3681,N_3392,N_3428);
nand U3682 (N_3682,N_3190,N_3109);
xnor U3683 (N_3683,N_3187,N_3237);
and U3684 (N_3684,N_3212,N_3330);
and U3685 (N_3685,N_3170,N_3351);
xor U3686 (N_3686,N_3093,N_3320);
nor U3687 (N_3687,N_3407,N_3436);
and U3688 (N_3688,N_3179,N_3262);
nor U3689 (N_3689,N_3432,N_3496);
or U3690 (N_3690,N_3386,N_3193);
nor U3691 (N_3691,N_3444,N_3427);
and U3692 (N_3692,N_3252,N_3379);
and U3693 (N_3693,N_3352,N_3116);
xor U3694 (N_3694,N_3440,N_3266);
nor U3695 (N_3695,N_3355,N_3012);
nor U3696 (N_3696,N_3498,N_3216);
nand U3697 (N_3697,N_3171,N_3464);
and U3698 (N_3698,N_3403,N_3467);
nor U3699 (N_3699,N_3318,N_3373);
nor U3700 (N_3700,N_3367,N_3039);
xor U3701 (N_3701,N_3277,N_3302);
nor U3702 (N_3702,N_3290,N_3111);
nand U3703 (N_3703,N_3487,N_3446);
and U3704 (N_3704,N_3064,N_3338);
and U3705 (N_3705,N_3017,N_3248);
and U3706 (N_3706,N_3234,N_3134);
nand U3707 (N_3707,N_3007,N_3422);
xnor U3708 (N_3708,N_3185,N_3002);
nor U3709 (N_3709,N_3375,N_3025);
nand U3710 (N_3710,N_3147,N_3303);
nor U3711 (N_3711,N_3066,N_3413);
nor U3712 (N_3712,N_3405,N_3013);
nor U3713 (N_3713,N_3433,N_3452);
nor U3714 (N_3714,N_3282,N_3083);
xor U3715 (N_3715,N_3003,N_3153);
and U3716 (N_3716,N_3325,N_3101);
nor U3717 (N_3717,N_3408,N_3004);
or U3718 (N_3718,N_3289,N_3090);
or U3719 (N_3719,N_3305,N_3280);
nor U3720 (N_3720,N_3491,N_3431);
nand U3721 (N_3721,N_3041,N_3195);
or U3722 (N_3722,N_3236,N_3174);
nand U3723 (N_3723,N_3220,N_3400);
and U3724 (N_3724,N_3347,N_3300);
nor U3725 (N_3725,N_3102,N_3314);
and U3726 (N_3726,N_3283,N_3222);
nor U3727 (N_3727,N_3410,N_3095);
xor U3728 (N_3728,N_3457,N_3398);
and U3729 (N_3729,N_3042,N_3168);
or U3730 (N_3730,N_3096,N_3388);
or U3731 (N_3731,N_3172,N_3331);
nand U3732 (N_3732,N_3297,N_3333);
and U3733 (N_3733,N_3188,N_3284);
and U3734 (N_3734,N_3204,N_3256);
nand U3735 (N_3735,N_3426,N_3223);
nor U3736 (N_3736,N_3441,N_3246);
and U3737 (N_3737,N_3316,N_3229);
nor U3738 (N_3738,N_3249,N_3269);
and U3739 (N_3739,N_3184,N_3128);
and U3740 (N_3740,N_3186,N_3458);
or U3741 (N_3741,N_3291,N_3448);
xor U3742 (N_3742,N_3124,N_3198);
nor U3743 (N_3743,N_3132,N_3078);
nor U3744 (N_3744,N_3307,N_3142);
and U3745 (N_3745,N_3424,N_3363);
nand U3746 (N_3746,N_3319,N_3265);
and U3747 (N_3747,N_3141,N_3478);
and U3748 (N_3748,N_3343,N_3415);
nand U3749 (N_3749,N_3264,N_3328);
or U3750 (N_3750,N_3442,N_3051);
and U3751 (N_3751,N_3259,N_3010);
and U3752 (N_3752,N_3127,N_3486);
nand U3753 (N_3753,N_3005,N_3177);
nor U3754 (N_3754,N_3439,N_3008);
xnor U3755 (N_3755,N_3446,N_3357);
and U3756 (N_3756,N_3459,N_3426);
and U3757 (N_3757,N_3498,N_3197);
xor U3758 (N_3758,N_3004,N_3296);
xnor U3759 (N_3759,N_3123,N_3156);
and U3760 (N_3760,N_3255,N_3212);
nor U3761 (N_3761,N_3107,N_3276);
and U3762 (N_3762,N_3094,N_3424);
nand U3763 (N_3763,N_3333,N_3165);
nand U3764 (N_3764,N_3093,N_3468);
and U3765 (N_3765,N_3142,N_3178);
and U3766 (N_3766,N_3264,N_3274);
nand U3767 (N_3767,N_3222,N_3225);
or U3768 (N_3768,N_3370,N_3160);
or U3769 (N_3769,N_3245,N_3390);
nand U3770 (N_3770,N_3068,N_3319);
or U3771 (N_3771,N_3175,N_3067);
nand U3772 (N_3772,N_3186,N_3097);
nor U3773 (N_3773,N_3095,N_3272);
xor U3774 (N_3774,N_3218,N_3282);
and U3775 (N_3775,N_3143,N_3221);
or U3776 (N_3776,N_3431,N_3468);
nor U3777 (N_3777,N_3269,N_3116);
xnor U3778 (N_3778,N_3254,N_3331);
nor U3779 (N_3779,N_3469,N_3494);
nor U3780 (N_3780,N_3113,N_3101);
xor U3781 (N_3781,N_3203,N_3459);
or U3782 (N_3782,N_3378,N_3101);
and U3783 (N_3783,N_3025,N_3282);
nor U3784 (N_3784,N_3079,N_3111);
nand U3785 (N_3785,N_3493,N_3218);
xnor U3786 (N_3786,N_3108,N_3059);
nor U3787 (N_3787,N_3126,N_3257);
xnor U3788 (N_3788,N_3159,N_3021);
nand U3789 (N_3789,N_3402,N_3302);
and U3790 (N_3790,N_3471,N_3414);
nand U3791 (N_3791,N_3036,N_3022);
nand U3792 (N_3792,N_3241,N_3182);
and U3793 (N_3793,N_3122,N_3112);
nand U3794 (N_3794,N_3445,N_3235);
nand U3795 (N_3795,N_3382,N_3391);
nand U3796 (N_3796,N_3351,N_3423);
nand U3797 (N_3797,N_3314,N_3284);
and U3798 (N_3798,N_3316,N_3438);
nor U3799 (N_3799,N_3126,N_3455);
and U3800 (N_3800,N_3201,N_3146);
or U3801 (N_3801,N_3082,N_3016);
nor U3802 (N_3802,N_3349,N_3294);
and U3803 (N_3803,N_3003,N_3108);
nor U3804 (N_3804,N_3266,N_3103);
or U3805 (N_3805,N_3460,N_3244);
and U3806 (N_3806,N_3120,N_3136);
nor U3807 (N_3807,N_3035,N_3069);
xnor U3808 (N_3808,N_3096,N_3446);
nor U3809 (N_3809,N_3263,N_3213);
nand U3810 (N_3810,N_3248,N_3476);
or U3811 (N_3811,N_3281,N_3045);
and U3812 (N_3812,N_3457,N_3397);
or U3813 (N_3813,N_3324,N_3452);
nor U3814 (N_3814,N_3067,N_3277);
and U3815 (N_3815,N_3466,N_3072);
nand U3816 (N_3816,N_3101,N_3055);
nor U3817 (N_3817,N_3173,N_3064);
or U3818 (N_3818,N_3155,N_3242);
xor U3819 (N_3819,N_3307,N_3092);
or U3820 (N_3820,N_3306,N_3292);
xor U3821 (N_3821,N_3069,N_3173);
xor U3822 (N_3822,N_3298,N_3311);
xnor U3823 (N_3823,N_3388,N_3310);
xor U3824 (N_3824,N_3131,N_3454);
xor U3825 (N_3825,N_3449,N_3082);
xnor U3826 (N_3826,N_3056,N_3139);
or U3827 (N_3827,N_3216,N_3080);
xnor U3828 (N_3828,N_3262,N_3150);
nand U3829 (N_3829,N_3430,N_3116);
and U3830 (N_3830,N_3492,N_3401);
nor U3831 (N_3831,N_3152,N_3355);
xnor U3832 (N_3832,N_3449,N_3206);
nand U3833 (N_3833,N_3018,N_3309);
and U3834 (N_3834,N_3256,N_3159);
or U3835 (N_3835,N_3048,N_3397);
and U3836 (N_3836,N_3465,N_3304);
and U3837 (N_3837,N_3008,N_3099);
nand U3838 (N_3838,N_3465,N_3233);
nor U3839 (N_3839,N_3452,N_3104);
nor U3840 (N_3840,N_3471,N_3245);
nor U3841 (N_3841,N_3417,N_3412);
nand U3842 (N_3842,N_3027,N_3091);
and U3843 (N_3843,N_3339,N_3205);
and U3844 (N_3844,N_3168,N_3214);
nor U3845 (N_3845,N_3417,N_3160);
and U3846 (N_3846,N_3160,N_3356);
nand U3847 (N_3847,N_3055,N_3452);
xnor U3848 (N_3848,N_3134,N_3091);
xor U3849 (N_3849,N_3025,N_3136);
nor U3850 (N_3850,N_3488,N_3082);
nand U3851 (N_3851,N_3011,N_3267);
nand U3852 (N_3852,N_3389,N_3146);
nor U3853 (N_3853,N_3362,N_3087);
nor U3854 (N_3854,N_3164,N_3478);
nand U3855 (N_3855,N_3077,N_3107);
and U3856 (N_3856,N_3293,N_3241);
nand U3857 (N_3857,N_3130,N_3410);
and U3858 (N_3858,N_3138,N_3476);
xnor U3859 (N_3859,N_3218,N_3437);
xnor U3860 (N_3860,N_3057,N_3088);
and U3861 (N_3861,N_3477,N_3254);
nand U3862 (N_3862,N_3316,N_3094);
nand U3863 (N_3863,N_3467,N_3487);
and U3864 (N_3864,N_3328,N_3350);
xor U3865 (N_3865,N_3308,N_3396);
and U3866 (N_3866,N_3327,N_3281);
nand U3867 (N_3867,N_3048,N_3449);
or U3868 (N_3868,N_3183,N_3450);
or U3869 (N_3869,N_3035,N_3121);
and U3870 (N_3870,N_3148,N_3139);
nand U3871 (N_3871,N_3206,N_3469);
and U3872 (N_3872,N_3066,N_3498);
xnor U3873 (N_3873,N_3026,N_3082);
or U3874 (N_3874,N_3445,N_3049);
nand U3875 (N_3875,N_3258,N_3163);
nor U3876 (N_3876,N_3288,N_3406);
and U3877 (N_3877,N_3144,N_3123);
nand U3878 (N_3878,N_3044,N_3280);
xor U3879 (N_3879,N_3304,N_3195);
and U3880 (N_3880,N_3000,N_3085);
nor U3881 (N_3881,N_3277,N_3091);
nand U3882 (N_3882,N_3265,N_3059);
nor U3883 (N_3883,N_3425,N_3162);
nor U3884 (N_3884,N_3181,N_3127);
nand U3885 (N_3885,N_3002,N_3176);
and U3886 (N_3886,N_3460,N_3044);
xor U3887 (N_3887,N_3431,N_3147);
or U3888 (N_3888,N_3463,N_3209);
nand U3889 (N_3889,N_3160,N_3382);
xor U3890 (N_3890,N_3171,N_3261);
nor U3891 (N_3891,N_3220,N_3136);
nor U3892 (N_3892,N_3352,N_3322);
xnor U3893 (N_3893,N_3166,N_3471);
xnor U3894 (N_3894,N_3090,N_3292);
xnor U3895 (N_3895,N_3163,N_3132);
or U3896 (N_3896,N_3172,N_3092);
nor U3897 (N_3897,N_3104,N_3430);
nand U3898 (N_3898,N_3078,N_3115);
xnor U3899 (N_3899,N_3398,N_3342);
and U3900 (N_3900,N_3332,N_3066);
or U3901 (N_3901,N_3403,N_3249);
nand U3902 (N_3902,N_3082,N_3124);
or U3903 (N_3903,N_3187,N_3423);
or U3904 (N_3904,N_3324,N_3447);
and U3905 (N_3905,N_3493,N_3115);
or U3906 (N_3906,N_3271,N_3290);
nand U3907 (N_3907,N_3005,N_3255);
and U3908 (N_3908,N_3301,N_3461);
and U3909 (N_3909,N_3101,N_3025);
and U3910 (N_3910,N_3466,N_3279);
xor U3911 (N_3911,N_3023,N_3230);
xor U3912 (N_3912,N_3395,N_3199);
nor U3913 (N_3913,N_3236,N_3395);
and U3914 (N_3914,N_3304,N_3414);
xnor U3915 (N_3915,N_3025,N_3298);
nor U3916 (N_3916,N_3259,N_3402);
or U3917 (N_3917,N_3306,N_3017);
or U3918 (N_3918,N_3401,N_3052);
or U3919 (N_3919,N_3191,N_3395);
or U3920 (N_3920,N_3191,N_3276);
and U3921 (N_3921,N_3360,N_3029);
nor U3922 (N_3922,N_3104,N_3072);
xor U3923 (N_3923,N_3343,N_3414);
xor U3924 (N_3924,N_3475,N_3293);
nor U3925 (N_3925,N_3174,N_3392);
and U3926 (N_3926,N_3361,N_3356);
and U3927 (N_3927,N_3186,N_3298);
xnor U3928 (N_3928,N_3056,N_3116);
nand U3929 (N_3929,N_3353,N_3387);
or U3930 (N_3930,N_3421,N_3085);
nand U3931 (N_3931,N_3014,N_3413);
nor U3932 (N_3932,N_3455,N_3009);
and U3933 (N_3933,N_3242,N_3100);
nand U3934 (N_3934,N_3312,N_3498);
nand U3935 (N_3935,N_3377,N_3408);
and U3936 (N_3936,N_3016,N_3154);
nor U3937 (N_3937,N_3393,N_3165);
nor U3938 (N_3938,N_3043,N_3482);
nor U3939 (N_3939,N_3258,N_3221);
xor U3940 (N_3940,N_3115,N_3268);
xor U3941 (N_3941,N_3008,N_3120);
or U3942 (N_3942,N_3045,N_3051);
nand U3943 (N_3943,N_3477,N_3308);
nor U3944 (N_3944,N_3375,N_3345);
and U3945 (N_3945,N_3070,N_3089);
nor U3946 (N_3946,N_3066,N_3436);
nor U3947 (N_3947,N_3421,N_3201);
nand U3948 (N_3948,N_3279,N_3110);
and U3949 (N_3949,N_3343,N_3309);
nand U3950 (N_3950,N_3184,N_3467);
nand U3951 (N_3951,N_3462,N_3150);
nor U3952 (N_3952,N_3038,N_3428);
xor U3953 (N_3953,N_3221,N_3347);
nor U3954 (N_3954,N_3407,N_3155);
or U3955 (N_3955,N_3331,N_3146);
nand U3956 (N_3956,N_3482,N_3097);
nand U3957 (N_3957,N_3067,N_3343);
or U3958 (N_3958,N_3298,N_3129);
nor U3959 (N_3959,N_3484,N_3058);
nor U3960 (N_3960,N_3113,N_3303);
nor U3961 (N_3961,N_3366,N_3079);
nor U3962 (N_3962,N_3310,N_3434);
xor U3963 (N_3963,N_3278,N_3155);
nand U3964 (N_3964,N_3375,N_3190);
nor U3965 (N_3965,N_3252,N_3341);
xnor U3966 (N_3966,N_3092,N_3423);
nand U3967 (N_3967,N_3149,N_3395);
xor U3968 (N_3968,N_3085,N_3353);
and U3969 (N_3969,N_3382,N_3062);
or U3970 (N_3970,N_3481,N_3195);
or U3971 (N_3971,N_3184,N_3428);
xor U3972 (N_3972,N_3388,N_3222);
nand U3973 (N_3973,N_3472,N_3079);
or U3974 (N_3974,N_3337,N_3412);
nor U3975 (N_3975,N_3013,N_3488);
and U3976 (N_3976,N_3332,N_3495);
xor U3977 (N_3977,N_3273,N_3205);
nand U3978 (N_3978,N_3021,N_3423);
or U3979 (N_3979,N_3099,N_3220);
or U3980 (N_3980,N_3467,N_3245);
or U3981 (N_3981,N_3107,N_3378);
and U3982 (N_3982,N_3146,N_3167);
or U3983 (N_3983,N_3159,N_3124);
or U3984 (N_3984,N_3475,N_3310);
xnor U3985 (N_3985,N_3333,N_3466);
or U3986 (N_3986,N_3237,N_3001);
or U3987 (N_3987,N_3285,N_3035);
or U3988 (N_3988,N_3495,N_3161);
and U3989 (N_3989,N_3414,N_3131);
nand U3990 (N_3990,N_3487,N_3308);
or U3991 (N_3991,N_3198,N_3345);
xnor U3992 (N_3992,N_3032,N_3190);
and U3993 (N_3993,N_3337,N_3438);
and U3994 (N_3994,N_3332,N_3478);
xor U3995 (N_3995,N_3116,N_3101);
nand U3996 (N_3996,N_3097,N_3084);
xor U3997 (N_3997,N_3113,N_3085);
and U3998 (N_3998,N_3265,N_3022);
nor U3999 (N_3999,N_3167,N_3115);
or U4000 (N_4000,N_3630,N_3643);
or U4001 (N_4001,N_3507,N_3709);
and U4002 (N_4002,N_3846,N_3549);
or U4003 (N_4003,N_3972,N_3789);
nor U4004 (N_4004,N_3819,N_3690);
nor U4005 (N_4005,N_3601,N_3682);
xnor U4006 (N_4006,N_3925,N_3628);
nand U4007 (N_4007,N_3978,N_3573);
nand U4008 (N_4008,N_3835,N_3769);
xor U4009 (N_4009,N_3512,N_3553);
xor U4010 (N_4010,N_3710,N_3716);
nor U4011 (N_4011,N_3566,N_3941);
or U4012 (N_4012,N_3797,N_3656);
or U4013 (N_4013,N_3645,N_3613);
and U4014 (N_4014,N_3733,N_3689);
and U4015 (N_4015,N_3794,N_3693);
and U4016 (N_4016,N_3775,N_3675);
nand U4017 (N_4017,N_3815,N_3806);
nor U4018 (N_4018,N_3639,N_3829);
and U4019 (N_4019,N_3917,N_3950);
and U4020 (N_4020,N_3793,N_3580);
nor U4021 (N_4021,N_3855,N_3625);
xnor U4022 (N_4022,N_3953,N_3878);
xnor U4023 (N_4023,N_3896,N_3697);
nand U4024 (N_4024,N_3754,N_3776);
and U4025 (N_4025,N_3755,N_3871);
or U4026 (N_4026,N_3823,N_3581);
xor U4027 (N_4027,N_3844,N_3652);
xor U4028 (N_4028,N_3686,N_3773);
nor U4029 (N_4029,N_3929,N_3830);
xnor U4030 (N_4030,N_3809,N_3884);
nor U4031 (N_4031,N_3914,N_3559);
nand U4032 (N_4032,N_3770,N_3713);
nor U4033 (N_4033,N_3670,N_3927);
nand U4034 (N_4034,N_3564,N_3665);
and U4035 (N_4035,N_3662,N_3707);
and U4036 (N_4036,N_3746,N_3872);
nand U4037 (N_4037,N_3781,N_3801);
xnor U4038 (N_4038,N_3936,N_3839);
and U4039 (N_4039,N_3785,N_3873);
nand U4040 (N_4040,N_3816,N_3623);
xnor U4041 (N_4041,N_3533,N_3582);
nand U4042 (N_4042,N_3536,N_3821);
or U4043 (N_4043,N_3931,N_3547);
xor U4044 (N_4044,N_3605,N_3525);
nor U4045 (N_4045,N_3933,N_3901);
nor U4046 (N_4046,N_3937,N_3699);
nor U4047 (N_4047,N_3779,N_3894);
and U4048 (N_4048,N_3555,N_3758);
nor U4049 (N_4049,N_3622,N_3934);
or U4050 (N_4050,N_3864,N_3597);
xnor U4051 (N_4051,N_3657,N_3585);
nand U4052 (N_4052,N_3834,N_3869);
xnor U4053 (N_4053,N_3938,N_3500);
and U4054 (N_4054,N_3552,N_3556);
xnor U4055 (N_4055,N_3868,N_3765);
nand U4056 (N_4056,N_3791,N_3833);
nor U4057 (N_4057,N_3870,N_3768);
nand U4058 (N_4058,N_3711,N_3596);
nand U4059 (N_4059,N_3983,N_3749);
xor U4060 (N_4060,N_3528,N_3703);
nor U4061 (N_4061,N_3893,N_3683);
and U4062 (N_4062,N_3503,N_3606);
nor U4063 (N_4063,N_3919,N_3629);
nor U4064 (N_4064,N_3837,N_3600);
and U4065 (N_4065,N_3522,N_3957);
xor U4066 (N_4066,N_3910,N_3620);
and U4067 (N_4067,N_3804,N_3539);
xor U4068 (N_4068,N_3644,N_3838);
nor U4069 (N_4069,N_3958,N_3861);
or U4070 (N_4070,N_3646,N_3718);
nor U4071 (N_4071,N_3965,N_3537);
xnor U4072 (N_4072,N_3681,N_3874);
nand U4073 (N_4073,N_3908,N_3915);
and U4074 (N_4074,N_3952,N_3742);
xnor U4075 (N_4075,N_3905,N_3848);
or U4076 (N_4076,N_3860,N_3722);
nor U4077 (N_4077,N_3603,N_3799);
nand U4078 (N_4078,N_3611,N_3966);
or U4079 (N_4079,N_3663,N_3532);
nand U4080 (N_4080,N_3863,N_3787);
or U4081 (N_4081,N_3761,N_3569);
nor U4082 (N_4082,N_3780,N_3955);
xnor U4083 (N_4083,N_3612,N_3543);
or U4084 (N_4084,N_3803,N_3760);
and U4085 (N_4085,N_3747,N_3947);
or U4086 (N_4086,N_3579,N_3546);
nor U4087 (N_4087,N_3825,N_3667);
xor U4088 (N_4088,N_3633,N_3880);
and U4089 (N_4089,N_3968,N_3999);
or U4090 (N_4090,N_3715,N_3504);
and U4091 (N_4091,N_3526,N_3614);
or U4092 (N_4092,N_3827,N_3788);
nand U4093 (N_4093,N_3949,N_3859);
and U4094 (N_4094,N_3772,N_3554);
nand U4095 (N_4095,N_3923,N_3777);
and U4096 (N_4096,N_3882,N_3990);
and U4097 (N_4097,N_3598,N_3700);
nor U4098 (N_4098,N_3530,N_3920);
nor U4099 (N_4099,N_3756,N_3515);
nor U4100 (N_4100,N_3624,N_3531);
nor U4101 (N_4101,N_3994,N_3694);
nand U4102 (N_4102,N_3841,N_3857);
xnor U4103 (N_4103,N_3850,N_3545);
nor U4104 (N_4104,N_3684,N_3971);
xor U4105 (N_4105,N_3640,N_3964);
and U4106 (N_4106,N_3724,N_3508);
and U4107 (N_4107,N_3664,N_3890);
nor U4108 (N_4108,N_3842,N_3895);
or U4109 (N_4109,N_3560,N_3784);
or U4110 (N_4110,N_3510,N_3858);
nor U4111 (N_4111,N_3669,N_3988);
nor U4112 (N_4112,N_3790,N_3509);
xnor U4113 (N_4113,N_3570,N_3744);
nand U4114 (N_4114,N_3759,N_3969);
nand U4115 (N_4115,N_3558,N_3604);
nor U4116 (N_4116,N_3691,N_3951);
nand U4117 (N_4117,N_3728,N_3668);
and U4118 (N_4118,N_3659,N_3617);
xnor U4119 (N_4119,N_3698,N_3942);
nand U4120 (N_4120,N_3609,N_3902);
nor U4121 (N_4121,N_3702,N_3960);
or U4122 (N_4122,N_3666,N_3680);
nor U4123 (N_4123,N_3701,N_3602);
or U4124 (N_4124,N_3762,N_3692);
and U4125 (N_4125,N_3538,N_3996);
or U4126 (N_4126,N_3725,N_3774);
nor U4127 (N_4127,N_3677,N_3524);
or U4128 (N_4128,N_3592,N_3610);
nor U4129 (N_4129,N_3995,N_3648);
and U4130 (N_4130,N_3527,N_3847);
xnor U4131 (N_4131,N_3735,N_3913);
xor U4132 (N_4132,N_3757,N_3717);
xnor U4133 (N_4133,N_3575,N_3740);
or U4134 (N_4134,N_3736,N_3578);
or U4135 (N_4135,N_3589,N_3705);
and U4136 (N_4136,N_3911,N_3587);
xor U4137 (N_4137,N_3907,N_3608);
or U4138 (N_4138,N_3909,N_3977);
xor U4139 (N_4139,N_3635,N_3976);
or U4140 (N_4140,N_3607,N_3655);
and U4141 (N_4141,N_3695,N_3822);
nor U4142 (N_4142,N_3583,N_3906);
or U4143 (N_4143,N_3814,N_3514);
or U4144 (N_4144,N_3866,N_3594);
or U4145 (N_4145,N_3731,N_3828);
and U4146 (N_4146,N_3678,N_3888);
nand U4147 (N_4147,N_3948,N_3634);
or U4148 (N_4148,N_3922,N_3892);
and U4149 (N_4149,N_3631,N_3981);
nand U4150 (N_4150,N_3732,N_3885);
nor U4151 (N_4151,N_3738,N_3904);
and U4152 (N_4152,N_3616,N_3889);
nand U4153 (N_4153,N_3807,N_3748);
nor U4154 (N_4154,N_3567,N_3752);
nor U4155 (N_4155,N_3518,N_3641);
nand U4156 (N_4156,N_3921,N_3877);
and U4157 (N_4157,N_3708,N_3562);
nor U4158 (N_4158,N_3540,N_3986);
and U4159 (N_4159,N_3824,N_3865);
and U4160 (N_4160,N_3796,N_3912);
nand U4161 (N_4161,N_3544,N_3820);
or U4162 (N_4162,N_3661,N_3529);
nor U4163 (N_4163,N_3706,N_3817);
and U4164 (N_4164,N_3939,N_3930);
xnor U4165 (N_4165,N_3924,N_3903);
xor U4166 (N_4166,N_3897,N_3517);
xor U4167 (N_4167,N_3973,N_3811);
xor U4168 (N_4168,N_3520,N_3654);
xor U4169 (N_4169,N_3626,N_3926);
and U4170 (N_4170,N_3980,N_3993);
xnor U4171 (N_4171,N_3962,N_3967);
and U4172 (N_4172,N_3808,N_3511);
or U4173 (N_4173,N_3795,N_3739);
and U4174 (N_4174,N_3997,N_3805);
and U4175 (N_4175,N_3741,N_3851);
or U4176 (N_4176,N_3568,N_3506);
nor U4177 (N_4177,N_3852,N_3551);
or U4178 (N_4178,N_3685,N_3541);
xnor U4179 (N_4179,N_3813,N_3723);
xor U4180 (N_4180,N_3638,N_3764);
or U4181 (N_4181,N_3737,N_3845);
nor U4182 (N_4182,N_3688,N_3672);
and U4183 (N_4183,N_3862,N_3619);
nor U4184 (N_4184,N_3875,N_3876);
and U4185 (N_4185,N_3812,N_3674);
nor U4186 (N_4186,N_3632,N_3800);
nand U4187 (N_4187,N_3928,N_3954);
or U4188 (N_4188,N_3687,N_3879);
xor U4189 (N_4189,N_3783,N_3900);
nor U4190 (N_4190,N_3577,N_3548);
nor U4191 (N_4191,N_3647,N_3658);
and U4192 (N_4192,N_3513,N_3588);
nand U4193 (N_4193,N_3721,N_3726);
or U4194 (N_4194,N_3572,N_3679);
and U4195 (N_4195,N_3563,N_3730);
nand U4196 (N_4196,N_3676,N_3763);
xor U4197 (N_4197,N_3959,N_3883);
nand U4198 (N_4198,N_3898,N_3649);
nor U4199 (N_4199,N_3970,N_3586);
or U4200 (N_4200,N_3849,N_3867);
or U4201 (N_4201,N_3918,N_3615);
or U4202 (N_4202,N_3734,N_3557);
xor U4203 (N_4203,N_3502,N_3987);
nand U4204 (N_4204,N_3714,N_3712);
and U4205 (N_4205,N_3992,N_3627);
nor U4206 (N_4206,N_3576,N_3571);
or U4207 (N_4207,N_3961,N_3565);
and U4208 (N_4208,N_3767,N_3982);
nand U4209 (N_4209,N_3956,N_3642);
xnor U4210 (N_4210,N_3963,N_3534);
or U4211 (N_4211,N_3940,N_3831);
nand U4212 (N_4212,N_3836,N_3745);
nand U4213 (N_4213,N_3561,N_3653);
xnor U4214 (N_4214,N_3550,N_3886);
nand U4215 (N_4215,N_3943,N_3771);
and U4216 (N_4216,N_3542,N_3535);
nand U4217 (N_4217,N_3998,N_3974);
or U4218 (N_4218,N_3854,N_3818);
or U4219 (N_4219,N_3719,N_3750);
nor U4220 (N_4220,N_3887,N_3671);
xnor U4221 (N_4221,N_3891,N_3810);
nor U4222 (N_4222,N_3636,N_3826);
nand U4223 (N_4223,N_3519,N_3899);
nor U4224 (N_4224,N_3975,N_3932);
xnor U4225 (N_4225,N_3651,N_3621);
xor U4226 (N_4226,N_3945,N_3786);
or U4227 (N_4227,N_3673,N_3985);
xor U4228 (N_4228,N_3751,N_3618);
nand U4229 (N_4229,N_3729,N_3798);
and U4230 (N_4230,N_3916,N_3782);
xor U4231 (N_4231,N_3505,N_3720);
nand U4232 (N_4232,N_3660,N_3853);
or U4233 (N_4233,N_3591,N_3935);
or U4234 (N_4234,N_3856,N_3727);
and U4235 (N_4235,N_3593,N_3574);
nand U4236 (N_4236,N_3802,N_3704);
or U4237 (N_4237,N_3637,N_3979);
nor U4238 (N_4238,N_3595,N_3843);
xor U4239 (N_4239,N_3501,N_3944);
or U4240 (N_4240,N_3521,N_3584);
nor U4241 (N_4241,N_3792,N_3989);
or U4242 (N_4242,N_3832,N_3516);
and U4243 (N_4243,N_3946,N_3743);
nand U4244 (N_4244,N_3523,N_3650);
nand U4245 (N_4245,N_3881,N_3991);
nor U4246 (N_4246,N_3778,N_3766);
nor U4247 (N_4247,N_3590,N_3599);
nand U4248 (N_4248,N_3984,N_3696);
xor U4249 (N_4249,N_3753,N_3840);
xnor U4250 (N_4250,N_3990,N_3750);
nor U4251 (N_4251,N_3983,N_3905);
xor U4252 (N_4252,N_3517,N_3649);
nor U4253 (N_4253,N_3758,N_3816);
nor U4254 (N_4254,N_3832,N_3500);
nand U4255 (N_4255,N_3952,N_3819);
nor U4256 (N_4256,N_3671,N_3520);
nor U4257 (N_4257,N_3577,N_3809);
nor U4258 (N_4258,N_3710,N_3888);
nand U4259 (N_4259,N_3784,N_3981);
nand U4260 (N_4260,N_3738,N_3552);
or U4261 (N_4261,N_3744,N_3717);
xor U4262 (N_4262,N_3712,N_3626);
nand U4263 (N_4263,N_3979,N_3774);
or U4264 (N_4264,N_3674,N_3876);
or U4265 (N_4265,N_3885,N_3580);
and U4266 (N_4266,N_3940,N_3603);
nand U4267 (N_4267,N_3696,N_3774);
or U4268 (N_4268,N_3814,N_3599);
xnor U4269 (N_4269,N_3820,N_3793);
nor U4270 (N_4270,N_3669,N_3782);
nand U4271 (N_4271,N_3770,N_3763);
nand U4272 (N_4272,N_3541,N_3861);
nand U4273 (N_4273,N_3895,N_3538);
or U4274 (N_4274,N_3864,N_3740);
xnor U4275 (N_4275,N_3732,N_3568);
xnor U4276 (N_4276,N_3909,N_3504);
xnor U4277 (N_4277,N_3970,N_3837);
or U4278 (N_4278,N_3726,N_3781);
xnor U4279 (N_4279,N_3553,N_3565);
xnor U4280 (N_4280,N_3614,N_3520);
nand U4281 (N_4281,N_3787,N_3728);
nand U4282 (N_4282,N_3878,N_3806);
and U4283 (N_4283,N_3698,N_3682);
nor U4284 (N_4284,N_3708,N_3566);
nor U4285 (N_4285,N_3755,N_3912);
xnor U4286 (N_4286,N_3654,N_3743);
nor U4287 (N_4287,N_3736,N_3514);
nand U4288 (N_4288,N_3961,N_3952);
nand U4289 (N_4289,N_3565,N_3710);
nor U4290 (N_4290,N_3689,N_3766);
or U4291 (N_4291,N_3560,N_3908);
xor U4292 (N_4292,N_3864,N_3775);
nand U4293 (N_4293,N_3599,N_3630);
nand U4294 (N_4294,N_3752,N_3974);
nand U4295 (N_4295,N_3980,N_3516);
nor U4296 (N_4296,N_3617,N_3516);
xor U4297 (N_4297,N_3737,N_3510);
nor U4298 (N_4298,N_3845,N_3656);
xor U4299 (N_4299,N_3869,N_3986);
or U4300 (N_4300,N_3690,N_3806);
or U4301 (N_4301,N_3530,N_3871);
nand U4302 (N_4302,N_3520,N_3537);
nor U4303 (N_4303,N_3900,N_3815);
nor U4304 (N_4304,N_3916,N_3581);
or U4305 (N_4305,N_3967,N_3849);
and U4306 (N_4306,N_3973,N_3619);
and U4307 (N_4307,N_3679,N_3847);
nand U4308 (N_4308,N_3781,N_3584);
xor U4309 (N_4309,N_3811,N_3859);
nor U4310 (N_4310,N_3940,N_3513);
and U4311 (N_4311,N_3600,N_3580);
and U4312 (N_4312,N_3595,N_3758);
xnor U4313 (N_4313,N_3764,N_3553);
nand U4314 (N_4314,N_3694,N_3533);
or U4315 (N_4315,N_3689,N_3527);
xor U4316 (N_4316,N_3562,N_3966);
xnor U4317 (N_4317,N_3570,N_3627);
or U4318 (N_4318,N_3568,N_3758);
and U4319 (N_4319,N_3656,N_3798);
or U4320 (N_4320,N_3904,N_3799);
and U4321 (N_4321,N_3986,N_3929);
or U4322 (N_4322,N_3774,N_3989);
nor U4323 (N_4323,N_3908,N_3581);
xor U4324 (N_4324,N_3609,N_3822);
nand U4325 (N_4325,N_3750,N_3541);
nand U4326 (N_4326,N_3948,N_3513);
and U4327 (N_4327,N_3902,N_3577);
nand U4328 (N_4328,N_3706,N_3589);
or U4329 (N_4329,N_3519,N_3598);
nand U4330 (N_4330,N_3855,N_3856);
or U4331 (N_4331,N_3592,N_3588);
or U4332 (N_4332,N_3811,N_3976);
and U4333 (N_4333,N_3638,N_3851);
or U4334 (N_4334,N_3770,N_3859);
nor U4335 (N_4335,N_3557,N_3761);
or U4336 (N_4336,N_3510,N_3716);
nor U4337 (N_4337,N_3616,N_3960);
and U4338 (N_4338,N_3931,N_3649);
nor U4339 (N_4339,N_3624,N_3610);
nand U4340 (N_4340,N_3620,N_3979);
or U4341 (N_4341,N_3849,N_3579);
or U4342 (N_4342,N_3953,N_3675);
nand U4343 (N_4343,N_3847,N_3909);
nand U4344 (N_4344,N_3971,N_3950);
or U4345 (N_4345,N_3866,N_3841);
or U4346 (N_4346,N_3596,N_3787);
nor U4347 (N_4347,N_3506,N_3914);
xnor U4348 (N_4348,N_3852,N_3529);
xnor U4349 (N_4349,N_3940,N_3808);
or U4350 (N_4350,N_3723,N_3697);
xnor U4351 (N_4351,N_3860,N_3918);
or U4352 (N_4352,N_3655,N_3823);
or U4353 (N_4353,N_3581,N_3866);
nor U4354 (N_4354,N_3645,N_3779);
xnor U4355 (N_4355,N_3955,N_3814);
or U4356 (N_4356,N_3635,N_3657);
nor U4357 (N_4357,N_3992,N_3655);
xor U4358 (N_4358,N_3715,N_3711);
xnor U4359 (N_4359,N_3562,N_3945);
xnor U4360 (N_4360,N_3599,N_3916);
nand U4361 (N_4361,N_3591,N_3705);
xnor U4362 (N_4362,N_3547,N_3927);
nand U4363 (N_4363,N_3849,N_3898);
and U4364 (N_4364,N_3980,N_3660);
nor U4365 (N_4365,N_3765,N_3948);
xnor U4366 (N_4366,N_3623,N_3919);
nor U4367 (N_4367,N_3569,N_3853);
nand U4368 (N_4368,N_3824,N_3931);
and U4369 (N_4369,N_3519,N_3542);
xnor U4370 (N_4370,N_3605,N_3823);
xnor U4371 (N_4371,N_3903,N_3627);
xor U4372 (N_4372,N_3948,N_3734);
and U4373 (N_4373,N_3914,N_3659);
nor U4374 (N_4374,N_3554,N_3622);
nand U4375 (N_4375,N_3837,N_3730);
xor U4376 (N_4376,N_3807,N_3855);
and U4377 (N_4377,N_3876,N_3732);
nand U4378 (N_4378,N_3818,N_3723);
or U4379 (N_4379,N_3635,N_3915);
nand U4380 (N_4380,N_3603,N_3861);
nand U4381 (N_4381,N_3907,N_3706);
nor U4382 (N_4382,N_3900,N_3734);
and U4383 (N_4383,N_3990,N_3810);
or U4384 (N_4384,N_3936,N_3763);
nand U4385 (N_4385,N_3556,N_3568);
nand U4386 (N_4386,N_3932,N_3944);
and U4387 (N_4387,N_3912,N_3580);
and U4388 (N_4388,N_3685,N_3893);
nor U4389 (N_4389,N_3539,N_3814);
nor U4390 (N_4390,N_3558,N_3862);
nand U4391 (N_4391,N_3954,N_3609);
xnor U4392 (N_4392,N_3937,N_3822);
nand U4393 (N_4393,N_3770,N_3789);
xor U4394 (N_4394,N_3651,N_3895);
nor U4395 (N_4395,N_3872,N_3724);
nor U4396 (N_4396,N_3634,N_3923);
nor U4397 (N_4397,N_3524,N_3573);
xnor U4398 (N_4398,N_3785,N_3540);
nand U4399 (N_4399,N_3648,N_3530);
nand U4400 (N_4400,N_3692,N_3913);
xor U4401 (N_4401,N_3506,N_3772);
or U4402 (N_4402,N_3740,N_3642);
xnor U4403 (N_4403,N_3737,N_3789);
and U4404 (N_4404,N_3663,N_3884);
or U4405 (N_4405,N_3590,N_3889);
and U4406 (N_4406,N_3857,N_3974);
and U4407 (N_4407,N_3996,N_3523);
or U4408 (N_4408,N_3526,N_3945);
and U4409 (N_4409,N_3703,N_3594);
xnor U4410 (N_4410,N_3922,N_3839);
and U4411 (N_4411,N_3964,N_3563);
nor U4412 (N_4412,N_3865,N_3698);
nor U4413 (N_4413,N_3537,N_3745);
nor U4414 (N_4414,N_3889,N_3887);
nor U4415 (N_4415,N_3959,N_3733);
nand U4416 (N_4416,N_3666,N_3603);
nor U4417 (N_4417,N_3707,N_3865);
nand U4418 (N_4418,N_3650,N_3794);
nand U4419 (N_4419,N_3879,N_3887);
xor U4420 (N_4420,N_3675,N_3533);
or U4421 (N_4421,N_3966,N_3738);
nor U4422 (N_4422,N_3909,N_3943);
or U4423 (N_4423,N_3638,N_3687);
and U4424 (N_4424,N_3906,N_3737);
nand U4425 (N_4425,N_3738,N_3729);
and U4426 (N_4426,N_3821,N_3991);
nand U4427 (N_4427,N_3989,N_3936);
nor U4428 (N_4428,N_3656,N_3857);
xor U4429 (N_4429,N_3757,N_3715);
nor U4430 (N_4430,N_3595,N_3905);
or U4431 (N_4431,N_3562,N_3925);
xnor U4432 (N_4432,N_3871,N_3808);
nand U4433 (N_4433,N_3614,N_3735);
nand U4434 (N_4434,N_3509,N_3942);
or U4435 (N_4435,N_3590,N_3940);
xnor U4436 (N_4436,N_3569,N_3735);
and U4437 (N_4437,N_3983,N_3583);
nand U4438 (N_4438,N_3954,N_3965);
or U4439 (N_4439,N_3753,N_3628);
and U4440 (N_4440,N_3917,N_3919);
xnor U4441 (N_4441,N_3507,N_3687);
xnor U4442 (N_4442,N_3782,N_3968);
and U4443 (N_4443,N_3509,N_3622);
or U4444 (N_4444,N_3693,N_3584);
nand U4445 (N_4445,N_3848,N_3774);
or U4446 (N_4446,N_3697,N_3903);
or U4447 (N_4447,N_3887,N_3683);
nor U4448 (N_4448,N_3845,N_3549);
and U4449 (N_4449,N_3874,N_3818);
or U4450 (N_4450,N_3819,N_3510);
xnor U4451 (N_4451,N_3759,N_3613);
or U4452 (N_4452,N_3520,N_3594);
and U4453 (N_4453,N_3985,N_3689);
and U4454 (N_4454,N_3956,N_3923);
or U4455 (N_4455,N_3647,N_3765);
xnor U4456 (N_4456,N_3662,N_3520);
or U4457 (N_4457,N_3930,N_3594);
or U4458 (N_4458,N_3527,N_3546);
or U4459 (N_4459,N_3666,N_3809);
and U4460 (N_4460,N_3993,N_3663);
nand U4461 (N_4461,N_3608,N_3692);
or U4462 (N_4462,N_3854,N_3667);
xnor U4463 (N_4463,N_3515,N_3532);
and U4464 (N_4464,N_3674,N_3989);
nand U4465 (N_4465,N_3746,N_3581);
and U4466 (N_4466,N_3667,N_3801);
or U4467 (N_4467,N_3637,N_3636);
and U4468 (N_4468,N_3803,N_3893);
nor U4469 (N_4469,N_3636,N_3550);
or U4470 (N_4470,N_3656,N_3957);
or U4471 (N_4471,N_3903,N_3822);
xnor U4472 (N_4472,N_3779,N_3821);
nand U4473 (N_4473,N_3570,N_3581);
nand U4474 (N_4474,N_3695,N_3954);
nor U4475 (N_4475,N_3963,N_3957);
nand U4476 (N_4476,N_3712,N_3596);
or U4477 (N_4477,N_3788,N_3976);
xnor U4478 (N_4478,N_3621,N_3700);
nand U4479 (N_4479,N_3613,N_3888);
xor U4480 (N_4480,N_3741,N_3953);
nor U4481 (N_4481,N_3958,N_3635);
nor U4482 (N_4482,N_3784,N_3537);
nor U4483 (N_4483,N_3567,N_3537);
or U4484 (N_4484,N_3705,N_3948);
xor U4485 (N_4485,N_3852,N_3579);
and U4486 (N_4486,N_3642,N_3639);
nand U4487 (N_4487,N_3542,N_3872);
or U4488 (N_4488,N_3934,N_3665);
xor U4489 (N_4489,N_3611,N_3959);
nand U4490 (N_4490,N_3579,N_3663);
nor U4491 (N_4491,N_3992,N_3841);
nand U4492 (N_4492,N_3722,N_3798);
or U4493 (N_4493,N_3976,N_3562);
and U4494 (N_4494,N_3718,N_3621);
nand U4495 (N_4495,N_3736,N_3596);
and U4496 (N_4496,N_3939,N_3740);
and U4497 (N_4497,N_3792,N_3775);
and U4498 (N_4498,N_3697,N_3802);
xnor U4499 (N_4499,N_3694,N_3663);
or U4500 (N_4500,N_4186,N_4461);
xor U4501 (N_4501,N_4226,N_4297);
nor U4502 (N_4502,N_4205,N_4006);
and U4503 (N_4503,N_4056,N_4265);
and U4504 (N_4504,N_4247,N_4048);
nor U4505 (N_4505,N_4143,N_4123);
nor U4506 (N_4506,N_4302,N_4422);
and U4507 (N_4507,N_4151,N_4380);
nor U4508 (N_4508,N_4209,N_4419);
and U4509 (N_4509,N_4045,N_4451);
xnor U4510 (N_4510,N_4442,N_4409);
nor U4511 (N_4511,N_4458,N_4218);
nand U4512 (N_4512,N_4373,N_4393);
nand U4513 (N_4513,N_4341,N_4215);
nand U4514 (N_4514,N_4402,N_4464);
and U4515 (N_4515,N_4032,N_4348);
and U4516 (N_4516,N_4110,N_4483);
nand U4517 (N_4517,N_4054,N_4162);
and U4518 (N_4518,N_4147,N_4026);
and U4519 (N_4519,N_4079,N_4099);
or U4520 (N_4520,N_4087,N_4234);
xnor U4521 (N_4521,N_4498,N_4421);
nor U4522 (N_4522,N_4038,N_4342);
nand U4523 (N_4523,N_4133,N_4331);
xnor U4524 (N_4524,N_4330,N_4183);
nor U4525 (N_4525,N_4303,N_4130);
and U4526 (N_4526,N_4202,N_4431);
and U4527 (N_4527,N_4138,N_4379);
or U4528 (N_4528,N_4263,N_4077);
nand U4529 (N_4529,N_4013,N_4453);
xnor U4530 (N_4530,N_4018,N_4352);
nor U4531 (N_4531,N_4141,N_4166);
xor U4532 (N_4532,N_4259,N_4069);
xnor U4533 (N_4533,N_4168,N_4043);
or U4534 (N_4534,N_4028,N_4105);
and U4535 (N_4535,N_4065,N_4493);
nand U4536 (N_4536,N_4125,N_4411);
nor U4537 (N_4537,N_4232,N_4437);
nor U4538 (N_4538,N_4358,N_4078);
xnor U4539 (N_4539,N_4176,N_4314);
and U4540 (N_4540,N_4128,N_4208);
nand U4541 (N_4541,N_4024,N_4333);
xor U4542 (N_4542,N_4478,N_4086);
nand U4543 (N_4543,N_4154,N_4093);
xnor U4544 (N_4544,N_4334,N_4175);
nor U4545 (N_4545,N_4378,N_4426);
nor U4546 (N_4546,N_4061,N_4363);
and U4547 (N_4547,N_4152,N_4413);
and U4548 (N_4548,N_4111,N_4137);
and U4549 (N_4549,N_4395,N_4047);
or U4550 (N_4550,N_4499,N_4441);
nor U4551 (N_4551,N_4295,N_4120);
xor U4552 (N_4552,N_4062,N_4200);
and U4553 (N_4553,N_4073,N_4354);
xor U4554 (N_4554,N_4273,N_4389);
and U4555 (N_4555,N_4067,N_4323);
xor U4556 (N_4556,N_4280,N_4156);
nor U4557 (N_4557,N_4456,N_4287);
nand U4558 (N_4558,N_4398,N_4148);
and U4559 (N_4559,N_4015,N_4091);
or U4560 (N_4560,N_4284,N_4479);
or U4561 (N_4561,N_4094,N_4212);
nand U4562 (N_4562,N_4353,N_4064);
and U4563 (N_4563,N_4374,N_4220);
and U4564 (N_4564,N_4468,N_4113);
or U4565 (N_4565,N_4324,N_4471);
and U4566 (N_4566,N_4249,N_4058);
nand U4567 (N_4567,N_4188,N_4177);
nor U4568 (N_4568,N_4288,N_4052);
nand U4569 (N_4569,N_4372,N_4443);
and U4570 (N_4570,N_4115,N_4486);
nand U4571 (N_4571,N_4294,N_4401);
or U4572 (N_4572,N_4410,N_4368);
or U4573 (N_4573,N_4037,N_4490);
nor U4574 (N_4574,N_4108,N_4083);
and U4575 (N_4575,N_4020,N_4440);
and U4576 (N_4576,N_4262,N_4469);
nand U4577 (N_4577,N_4167,N_4072);
or U4578 (N_4578,N_4060,N_4124);
nor U4579 (N_4579,N_4217,N_4362);
xnor U4580 (N_4580,N_4198,N_4477);
and U4581 (N_4581,N_4206,N_4261);
and U4582 (N_4582,N_4452,N_4325);
nor U4583 (N_4583,N_4191,N_4213);
or U4584 (N_4584,N_4116,N_4428);
nand U4585 (N_4585,N_4196,N_4491);
nor U4586 (N_4586,N_4278,N_4350);
or U4587 (N_4587,N_4383,N_4436);
nand U4588 (N_4588,N_4150,N_4327);
xor U4589 (N_4589,N_4246,N_4408);
or U4590 (N_4590,N_4290,N_4369);
xnor U4591 (N_4591,N_4158,N_4476);
nand U4592 (N_4592,N_4257,N_4255);
or U4593 (N_4593,N_4169,N_4454);
xnor U4594 (N_4594,N_4121,N_4224);
or U4595 (N_4595,N_4328,N_4082);
nand U4596 (N_4596,N_4267,N_4204);
or U4597 (N_4597,N_4495,N_4240);
xor U4598 (N_4598,N_4460,N_4256);
nor U4599 (N_4599,N_4384,N_4173);
nor U4600 (N_4600,N_4207,N_4236);
nor U4601 (N_4601,N_4397,N_4201);
and U4602 (N_4602,N_4134,N_4185);
and U4603 (N_4603,N_4466,N_4070);
and U4604 (N_4604,N_4429,N_4400);
and U4605 (N_4605,N_4475,N_4057);
xnor U4606 (N_4606,N_4161,N_4068);
or U4607 (N_4607,N_4049,N_4066);
and U4608 (N_4608,N_4434,N_4274);
xor U4609 (N_4609,N_4438,N_4301);
nand U4610 (N_4610,N_4364,N_4392);
and U4611 (N_4611,N_4322,N_4455);
nand U4612 (N_4612,N_4450,N_4423);
nor U4613 (N_4613,N_4055,N_4310);
or U4614 (N_4614,N_4473,N_4085);
xor U4615 (N_4615,N_4031,N_4326);
nor U4616 (N_4616,N_4140,N_4007);
nor U4617 (N_4617,N_4357,N_4251);
nor U4618 (N_4618,N_4386,N_4272);
and U4619 (N_4619,N_4193,N_4285);
nor U4620 (N_4620,N_4371,N_4223);
or U4621 (N_4621,N_4035,N_4109);
or U4622 (N_4622,N_4306,N_4157);
or U4623 (N_4623,N_4399,N_4027);
and U4624 (N_4624,N_4396,N_4404);
nor U4625 (N_4625,N_4470,N_4416);
nor U4626 (N_4626,N_4343,N_4114);
nor U4627 (N_4627,N_4139,N_4427);
nand U4628 (N_4628,N_4254,N_4155);
and U4629 (N_4629,N_4430,N_4317);
xor U4630 (N_4630,N_4203,N_4266);
or U4631 (N_4631,N_4283,N_4112);
nand U4632 (N_4632,N_4277,N_4033);
and U4633 (N_4633,N_4172,N_4019);
or U4634 (N_4634,N_4126,N_4300);
xnor U4635 (N_4635,N_4012,N_4252);
nor U4636 (N_4636,N_4009,N_4448);
nor U4637 (N_4637,N_4039,N_4349);
nor U4638 (N_4638,N_4275,N_4046);
or U4639 (N_4639,N_4394,N_4420);
nand U4640 (N_4640,N_4474,N_4102);
nor U4641 (N_4641,N_4377,N_4316);
or U4642 (N_4642,N_4041,N_4345);
xnor U4643 (N_4643,N_4304,N_4281);
nor U4644 (N_4644,N_4279,N_4403);
nand U4645 (N_4645,N_4210,N_4312);
xor U4646 (N_4646,N_4346,N_4367);
nand U4647 (N_4647,N_4117,N_4268);
and U4648 (N_4648,N_4230,N_4182);
xor U4649 (N_4649,N_4164,N_4090);
nand U4650 (N_4650,N_4309,N_4003);
nor U4651 (N_4651,N_4320,N_4189);
or U4652 (N_4652,N_4307,N_4004);
xnor U4653 (N_4653,N_4299,N_4017);
xor U4654 (N_4654,N_4487,N_4233);
nand U4655 (N_4655,N_4344,N_4445);
nor U4656 (N_4656,N_4036,N_4365);
and U4657 (N_4657,N_4488,N_4005);
nor U4658 (N_4658,N_4329,N_4075);
xor U4659 (N_4659,N_4135,N_4418);
nor U4660 (N_4660,N_4104,N_4253);
nor U4661 (N_4661,N_4076,N_4412);
nor U4662 (N_4662,N_4339,N_4286);
nand U4663 (N_4663,N_4485,N_4228);
nand U4664 (N_4664,N_4472,N_4489);
xor U4665 (N_4665,N_4163,N_4089);
xor U4666 (N_4666,N_4180,N_4034);
or U4667 (N_4667,N_4237,N_4029);
nor U4668 (N_4668,N_4264,N_4282);
nand U4669 (N_4669,N_4424,N_4332);
or U4670 (N_4670,N_4023,N_4337);
xnor U4671 (N_4671,N_4214,N_4435);
or U4672 (N_4672,N_4092,N_4366);
or U4673 (N_4673,N_4336,N_4227);
and U4674 (N_4674,N_4225,N_4293);
xnor U4675 (N_4675,N_4291,N_4088);
nand U4676 (N_4676,N_4145,N_4390);
and U4677 (N_4677,N_4480,N_4107);
and U4678 (N_4678,N_4002,N_4462);
xor U4679 (N_4679,N_4229,N_4417);
or U4680 (N_4680,N_4439,N_4181);
or U4681 (N_4681,N_4482,N_4248);
nor U4682 (N_4682,N_4053,N_4360);
and U4683 (N_4683,N_4381,N_4496);
and U4684 (N_4684,N_4391,N_4465);
or U4685 (N_4685,N_4347,N_4221);
nor U4686 (N_4686,N_4165,N_4425);
xnor U4687 (N_4687,N_4197,N_4071);
or U4688 (N_4688,N_4179,N_4101);
and U4689 (N_4689,N_4359,N_4433);
xor U4690 (N_4690,N_4040,N_4042);
xor U4691 (N_4691,N_4447,N_4340);
nand U4692 (N_4692,N_4497,N_4244);
xnor U4693 (N_4693,N_4296,N_4415);
or U4694 (N_4694,N_4119,N_4080);
nor U4695 (N_4695,N_4335,N_4387);
and U4696 (N_4696,N_4298,N_4001);
and U4697 (N_4697,N_4351,N_4376);
and U4698 (N_4698,N_4484,N_4097);
or U4699 (N_4699,N_4492,N_4219);
nor U4700 (N_4700,N_4239,N_4190);
nand U4701 (N_4701,N_4096,N_4030);
or U4702 (N_4702,N_4014,N_4449);
nor U4703 (N_4703,N_4074,N_4270);
nand U4704 (N_4704,N_4481,N_4370);
nand U4705 (N_4705,N_4171,N_4463);
or U4706 (N_4706,N_4315,N_4242);
or U4707 (N_4707,N_4355,N_4414);
nand U4708 (N_4708,N_4245,N_4318);
xnor U4709 (N_4709,N_4269,N_4241);
or U4710 (N_4710,N_4051,N_4127);
nand U4711 (N_4711,N_4160,N_4149);
nor U4712 (N_4712,N_4385,N_4235);
xnor U4713 (N_4713,N_4081,N_4243);
and U4714 (N_4714,N_4199,N_4016);
and U4715 (N_4715,N_4432,N_4192);
xor U4716 (N_4716,N_4338,N_4407);
nand U4717 (N_4717,N_4044,N_4025);
nor U4718 (N_4718,N_4178,N_4313);
or U4719 (N_4719,N_4382,N_4406);
xnor U4720 (N_4720,N_4021,N_4142);
or U4721 (N_4721,N_4184,N_4457);
nand U4722 (N_4722,N_4100,N_4146);
nand U4723 (N_4723,N_4276,N_4098);
nand U4724 (N_4724,N_4136,N_4194);
or U4725 (N_4725,N_4132,N_4319);
xor U4726 (N_4726,N_4170,N_4010);
nor U4727 (N_4727,N_4159,N_4063);
and U4728 (N_4728,N_4467,N_4059);
nor U4729 (N_4729,N_4305,N_4405);
nor U4730 (N_4730,N_4289,N_4388);
nand U4731 (N_4731,N_4011,N_4271);
xor U4732 (N_4732,N_4308,N_4459);
or U4733 (N_4733,N_4250,N_4311);
nor U4734 (N_4734,N_4144,N_4195);
or U4735 (N_4735,N_4231,N_4375);
xor U4736 (N_4736,N_4103,N_4494);
and U4737 (N_4737,N_4084,N_4211);
xor U4738 (N_4738,N_4118,N_4444);
and U4739 (N_4739,N_4008,N_4187);
or U4740 (N_4740,N_4153,N_4260);
or U4741 (N_4741,N_4000,N_4129);
or U4742 (N_4742,N_4131,N_4238);
nor U4743 (N_4743,N_4446,N_4216);
nand U4744 (N_4744,N_4258,N_4174);
xor U4745 (N_4745,N_4321,N_4356);
nand U4746 (N_4746,N_4050,N_4022);
nor U4747 (N_4747,N_4222,N_4361);
or U4748 (N_4748,N_4106,N_4095);
and U4749 (N_4749,N_4292,N_4122);
nand U4750 (N_4750,N_4119,N_4168);
or U4751 (N_4751,N_4204,N_4207);
or U4752 (N_4752,N_4033,N_4174);
nor U4753 (N_4753,N_4222,N_4266);
nor U4754 (N_4754,N_4470,N_4257);
xnor U4755 (N_4755,N_4161,N_4039);
nand U4756 (N_4756,N_4339,N_4412);
nor U4757 (N_4757,N_4496,N_4054);
nor U4758 (N_4758,N_4243,N_4252);
nand U4759 (N_4759,N_4096,N_4330);
xor U4760 (N_4760,N_4116,N_4406);
nand U4761 (N_4761,N_4155,N_4061);
and U4762 (N_4762,N_4122,N_4346);
and U4763 (N_4763,N_4099,N_4222);
nor U4764 (N_4764,N_4209,N_4131);
and U4765 (N_4765,N_4289,N_4355);
or U4766 (N_4766,N_4260,N_4137);
and U4767 (N_4767,N_4152,N_4019);
nor U4768 (N_4768,N_4416,N_4078);
nor U4769 (N_4769,N_4129,N_4329);
nand U4770 (N_4770,N_4068,N_4078);
nand U4771 (N_4771,N_4292,N_4421);
or U4772 (N_4772,N_4032,N_4109);
nor U4773 (N_4773,N_4260,N_4236);
xor U4774 (N_4774,N_4358,N_4235);
or U4775 (N_4775,N_4367,N_4272);
xor U4776 (N_4776,N_4437,N_4211);
xor U4777 (N_4777,N_4234,N_4424);
nand U4778 (N_4778,N_4267,N_4459);
and U4779 (N_4779,N_4367,N_4412);
or U4780 (N_4780,N_4337,N_4309);
xnor U4781 (N_4781,N_4455,N_4084);
xor U4782 (N_4782,N_4031,N_4470);
nand U4783 (N_4783,N_4195,N_4310);
or U4784 (N_4784,N_4253,N_4049);
nand U4785 (N_4785,N_4368,N_4417);
or U4786 (N_4786,N_4431,N_4273);
nor U4787 (N_4787,N_4306,N_4332);
nand U4788 (N_4788,N_4426,N_4482);
nand U4789 (N_4789,N_4281,N_4386);
nor U4790 (N_4790,N_4318,N_4322);
nand U4791 (N_4791,N_4368,N_4380);
xnor U4792 (N_4792,N_4176,N_4275);
and U4793 (N_4793,N_4337,N_4169);
or U4794 (N_4794,N_4096,N_4014);
nor U4795 (N_4795,N_4352,N_4104);
nor U4796 (N_4796,N_4066,N_4341);
nor U4797 (N_4797,N_4335,N_4400);
xor U4798 (N_4798,N_4312,N_4207);
and U4799 (N_4799,N_4459,N_4021);
or U4800 (N_4800,N_4284,N_4356);
and U4801 (N_4801,N_4346,N_4301);
or U4802 (N_4802,N_4281,N_4163);
nand U4803 (N_4803,N_4131,N_4139);
and U4804 (N_4804,N_4277,N_4040);
xnor U4805 (N_4805,N_4111,N_4148);
and U4806 (N_4806,N_4220,N_4249);
xor U4807 (N_4807,N_4171,N_4465);
and U4808 (N_4808,N_4163,N_4327);
xor U4809 (N_4809,N_4070,N_4416);
and U4810 (N_4810,N_4191,N_4272);
nor U4811 (N_4811,N_4153,N_4217);
or U4812 (N_4812,N_4454,N_4154);
and U4813 (N_4813,N_4315,N_4328);
xnor U4814 (N_4814,N_4224,N_4471);
nand U4815 (N_4815,N_4329,N_4223);
nand U4816 (N_4816,N_4320,N_4094);
xor U4817 (N_4817,N_4414,N_4166);
xor U4818 (N_4818,N_4202,N_4263);
nand U4819 (N_4819,N_4046,N_4350);
xnor U4820 (N_4820,N_4119,N_4318);
nor U4821 (N_4821,N_4155,N_4035);
xor U4822 (N_4822,N_4201,N_4207);
nand U4823 (N_4823,N_4009,N_4393);
or U4824 (N_4824,N_4499,N_4266);
or U4825 (N_4825,N_4378,N_4389);
nor U4826 (N_4826,N_4491,N_4473);
or U4827 (N_4827,N_4194,N_4196);
nand U4828 (N_4828,N_4086,N_4197);
xnor U4829 (N_4829,N_4438,N_4218);
xor U4830 (N_4830,N_4273,N_4429);
or U4831 (N_4831,N_4460,N_4437);
nor U4832 (N_4832,N_4114,N_4184);
nand U4833 (N_4833,N_4404,N_4080);
xnor U4834 (N_4834,N_4387,N_4434);
nand U4835 (N_4835,N_4344,N_4309);
xor U4836 (N_4836,N_4426,N_4382);
nand U4837 (N_4837,N_4312,N_4163);
or U4838 (N_4838,N_4423,N_4131);
and U4839 (N_4839,N_4248,N_4211);
nand U4840 (N_4840,N_4099,N_4448);
and U4841 (N_4841,N_4152,N_4200);
and U4842 (N_4842,N_4473,N_4267);
xnor U4843 (N_4843,N_4165,N_4364);
xnor U4844 (N_4844,N_4135,N_4267);
and U4845 (N_4845,N_4384,N_4101);
nand U4846 (N_4846,N_4326,N_4335);
nor U4847 (N_4847,N_4239,N_4475);
and U4848 (N_4848,N_4016,N_4441);
and U4849 (N_4849,N_4476,N_4219);
or U4850 (N_4850,N_4357,N_4078);
nand U4851 (N_4851,N_4268,N_4299);
nand U4852 (N_4852,N_4397,N_4005);
and U4853 (N_4853,N_4267,N_4152);
and U4854 (N_4854,N_4229,N_4224);
nor U4855 (N_4855,N_4426,N_4411);
xor U4856 (N_4856,N_4457,N_4138);
nand U4857 (N_4857,N_4237,N_4491);
or U4858 (N_4858,N_4423,N_4362);
nor U4859 (N_4859,N_4009,N_4201);
nand U4860 (N_4860,N_4407,N_4438);
and U4861 (N_4861,N_4015,N_4362);
nand U4862 (N_4862,N_4072,N_4423);
nor U4863 (N_4863,N_4124,N_4441);
and U4864 (N_4864,N_4352,N_4006);
nor U4865 (N_4865,N_4320,N_4125);
nand U4866 (N_4866,N_4294,N_4217);
xor U4867 (N_4867,N_4300,N_4381);
nor U4868 (N_4868,N_4329,N_4258);
or U4869 (N_4869,N_4047,N_4415);
nor U4870 (N_4870,N_4495,N_4355);
or U4871 (N_4871,N_4302,N_4215);
nand U4872 (N_4872,N_4384,N_4457);
xor U4873 (N_4873,N_4270,N_4238);
nand U4874 (N_4874,N_4055,N_4269);
or U4875 (N_4875,N_4391,N_4268);
nor U4876 (N_4876,N_4016,N_4419);
xor U4877 (N_4877,N_4252,N_4003);
nor U4878 (N_4878,N_4101,N_4158);
nor U4879 (N_4879,N_4423,N_4344);
nor U4880 (N_4880,N_4033,N_4342);
nor U4881 (N_4881,N_4332,N_4151);
and U4882 (N_4882,N_4008,N_4222);
nand U4883 (N_4883,N_4039,N_4422);
nor U4884 (N_4884,N_4090,N_4401);
nor U4885 (N_4885,N_4119,N_4287);
or U4886 (N_4886,N_4311,N_4173);
nor U4887 (N_4887,N_4266,N_4106);
and U4888 (N_4888,N_4367,N_4381);
or U4889 (N_4889,N_4463,N_4335);
nand U4890 (N_4890,N_4450,N_4173);
or U4891 (N_4891,N_4035,N_4167);
and U4892 (N_4892,N_4034,N_4032);
nand U4893 (N_4893,N_4406,N_4332);
or U4894 (N_4894,N_4001,N_4103);
and U4895 (N_4895,N_4282,N_4470);
and U4896 (N_4896,N_4384,N_4058);
xnor U4897 (N_4897,N_4110,N_4130);
nand U4898 (N_4898,N_4100,N_4383);
xnor U4899 (N_4899,N_4479,N_4107);
nand U4900 (N_4900,N_4027,N_4462);
and U4901 (N_4901,N_4451,N_4421);
or U4902 (N_4902,N_4226,N_4210);
nand U4903 (N_4903,N_4421,N_4004);
or U4904 (N_4904,N_4417,N_4113);
xnor U4905 (N_4905,N_4297,N_4196);
and U4906 (N_4906,N_4102,N_4381);
or U4907 (N_4907,N_4430,N_4274);
nand U4908 (N_4908,N_4077,N_4367);
xor U4909 (N_4909,N_4302,N_4049);
and U4910 (N_4910,N_4395,N_4158);
xnor U4911 (N_4911,N_4450,N_4244);
nand U4912 (N_4912,N_4422,N_4092);
nand U4913 (N_4913,N_4337,N_4197);
and U4914 (N_4914,N_4118,N_4395);
xor U4915 (N_4915,N_4178,N_4411);
nor U4916 (N_4916,N_4045,N_4286);
nor U4917 (N_4917,N_4322,N_4040);
nand U4918 (N_4918,N_4117,N_4403);
nand U4919 (N_4919,N_4361,N_4450);
xnor U4920 (N_4920,N_4176,N_4135);
or U4921 (N_4921,N_4335,N_4389);
nor U4922 (N_4922,N_4120,N_4304);
nand U4923 (N_4923,N_4079,N_4028);
nand U4924 (N_4924,N_4224,N_4298);
or U4925 (N_4925,N_4259,N_4200);
xor U4926 (N_4926,N_4130,N_4439);
nor U4927 (N_4927,N_4185,N_4346);
or U4928 (N_4928,N_4305,N_4172);
and U4929 (N_4929,N_4061,N_4293);
or U4930 (N_4930,N_4459,N_4257);
nor U4931 (N_4931,N_4478,N_4105);
or U4932 (N_4932,N_4434,N_4297);
and U4933 (N_4933,N_4411,N_4166);
and U4934 (N_4934,N_4089,N_4069);
or U4935 (N_4935,N_4309,N_4200);
and U4936 (N_4936,N_4279,N_4273);
xnor U4937 (N_4937,N_4135,N_4238);
nand U4938 (N_4938,N_4278,N_4394);
and U4939 (N_4939,N_4342,N_4315);
or U4940 (N_4940,N_4412,N_4158);
and U4941 (N_4941,N_4072,N_4074);
and U4942 (N_4942,N_4422,N_4234);
and U4943 (N_4943,N_4245,N_4117);
xor U4944 (N_4944,N_4149,N_4151);
nor U4945 (N_4945,N_4027,N_4107);
xnor U4946 (N_4946,N_4028,N_4011);
nand U4947 (N_4947,N_4067,N_4358);
nor U4948 (N_4948,N_4047,N_4203);
and U4949 (N_4949,N_4467,N_4185);
xor U4950 (N_4950,N_4006,N_4151);
xor U4951 (N_4951,N_4388,N_4157);
nand U4952 (N_4952,N_4025,N_4216);
nand U4953 (N_4953,N_4078,N_4425);
and U4954 (N_4954,N_4456,N_4250);
or U4955 (N_4955,N_4231,N_4408);
and U4956 (N_4956,N_4331,N_4051);
xnor U4957 (N_4957,N_4154,N_4029);
or U4958 (N_4958,N_4211,N_4190);
nand U4959 (N_4959,N_4063,N_4001);
nand U4960 (N_4960,N_4340,N_4149);
and U4961 (N_4961,N_4185,N_4433);
nand U4962 (N_4962,N_4177,N_4397);
nand U4963 (N_4963,N_4482,N_4346);
nand U4964 (N_4964,N_4058,N_4342);
xnor U4965 (N_4965,N_4053,N_4218);
or U4966 (N_4966,N_4302,N_4016);
nand U4967 (N_4967,N_4201,N_4430);
nor U4968 (N_4968,N_4049,N_4070);
nor U4969 (N_4969,N_4097,N_4064);
nand U4970 (N_4970,N_4302,N_4243);
and U4971 (N_4971,N_4388,N_4360);
and U4972 (N_4972,N_4050,N_4074);
nand U4973 (N_4973,N_4393,N_4069);
and U4974 (N_4974,N_4387,N_4357);
nor U4975 (N_4975,N_4426,N_4338);
xnor U4976 (N_4976,N_4369,N_4106);
or U4977 (N_4977,N_4432,N_4310);
nor U4978 (N_4978,N_4306,N_4265);
and U4979 (N_4979,N_4370,N_4149);
xnor U4980 (N_4980,N_4248,N_4489);
or U4981 (N_4981,N_4100,N_4455);
and U4982 (N_4982,N_4303,N_4286);
xor U4983 (N_4983,N_4455,N_4067);
and U4984 (N_4984,N_4328,N_4011);
nor U4985 (N_4985,N_4004,N_4017);
or U4986 (N_4986,N_4417,N_4388);
and U4987 (N_4987,N_4126,N_4401);
xnor U4988 (N_4988,N_4450,N_4122);
or U4989 (N_4989,N_4359,N_4423);
xnor U4990 (N_4990,N_4220,N_4144);
or U4991 (N_4991,N_4265,N_4196);
nor U4992 (N_4992,N_4202,N_4495);
and U4993 (N_4993,N_4318,N_4103);
nor U4994 (N_4994,N_4151,N_4124);
xor U4995 (N_4995,N_4280,N_4386);
nor U4996 (N_4996,N_4488,N_4343);
or U4997 (N_4997,N_4464,N_4409);
or U4998 (N_4998,N_4155,N_4206);
or U4999 (N_4999,N_4395,N_4497);
nor U5000 (N_5000,N_4848,N_4877);
nand U5001 (N_5001,N_4713,N_4680);
nor U5002 (N_5002,N_4801,N_4997);
nand U5003 (N_5003,N_4571,N_4780);
nand U5004 (N_5004,N_4628,N_4561);
nor U5005 (N_5005,N_4541,N_4810);
and U5006 (N_5006,N_4649,N_4808);
xnor U5007 (N_5007,N_4904,N_4932);
xor U5008 (N_5008,N_4839,N_4703);
nor U5009 (N_5009,N_4934,N_4684);
xnor U5010 (N_5010,N_4554,N_4662);
xnor U5011 (N_5011,N_4724,N_4720);
or U5012 (N_5012,N_4874,N_4772);
and U5013 (N_5013,N_4778,N_4697);
nor U5014 (N_5014,N_4719,N_4721);
nand U5015 (N_5015,N_4855,N_4610);
or U5016 (N_5016,N_4613,N_4798);
or U5017 (N_5017,N_4601,N_4756);
xor U5018 (N_5018,N_4592,N_4923);
nor U5019 (N_5019,N_4889,N_4815);
nor U5020 (N_5020,N_4735,N_4811);
or U5021 (N_5021,N_4971,N_4841);
nor U5022 (N_5022,N_4599,N_4786);
nor U5023 (N_5023,N_4701,N_4645);
nand U5024 (N_5024,N_4709,N_4749);
xor U5025 (N_5025,N_4885,N_4830);
or U5026 (N_5026,N_4819,N_4531);
xnor U5027 (N_5027,N_4942,N_4573);
nor U5028 (N_5028,N_4667,N_4868);
nand U5029 (N_5029,N_4569,N_4818);
nor U5030 (N_5030,N_4898,N_4725);
nor U5031 (N_5031,N_4681,N_4560);
xnor U5032 (N_5032,N_4948,N_4553);
xnor U5033 (N_5033,N_4957,N_4859);
or U5034 (N_5034,N_4979,N_4500);
or U5035 (N_5035,N_4551,N_4552);
nand U5036 (N_5036,N_4911,N_4805);
xor U5037 (N_5037,N_4717,N_4529);
nor U5038 (N_5038,N_4807,N_4890);
xor U5039 (N_5039,N_4823,N_4856);
xnor U5040 (N_5040,N_4776,N_4799);
nor U5041 (N_5041,N_4639,N_4520);
nor U5042 (N_5042,N_4521,N_4764);
xor U5043 (N_5043,N_4590,N_4967);
nand U5044 (N_5044,N_4501,N_4995);
or U5045 (N_5045,N_4666,N_4692);
and U5046 (N_5046,N_4733,N_4643);
nor U5047 (N_5047,N_4753,N_4982);
and U5048 (N_5048,N_4837,N_4872);
nor U5049 (N_5049,N_4887,N_4793);
nor U5050 (N_5050,N_4984,N_4705);
and U5051 (N_5051,N_4609,N_4527);
xor U5052 (N_5052,N_4858,N_4828);
nand U5053 (N_5053,N_4739,N_4802);
xnor U5054 (N_5054,N_4936,N_4897);
xnor U5055 (N_5055,N_4655,N_4933);
nand U5056 (N_5056,N_4876,N_4760);
nor U5057 (N_5057,N_4998,N_4675);
nand U5058 (N_5058,N_4768,N_4952);
or U5059 (N_5059,N_4714,N_4690);
nor U5060 (N_5060,N_4706,N_4635);
nor U5061 (N_5061,N_4921,N_4939);
nand U5062 (N_5062,N_4908,N_4530);
and U5063 (N_5063,N_4992,N_4761);
nor U5064 (N_5064,N_4730,N_4814);
xor U5065 (N_5065,N_4652,N_4928);
nand U5066 (N_5066,N_4833,N_4914);
xor U5067 (N_5067,N_4661,N_4836);
and U5068 (N_5068,N_4976,N_4895);
or U5069 (N_5069,N_4926,N_4779);
and U5070 (N_5070,N_4827,N_4822);
nand U5071 (N_5071,N_4596,N_4674);
xor U5072 (N_5072,N_4647,N_4862);
nand U5073 (N_5073,N_4960,N_4962);
and U5074 (N_5074,N_4737,N_4965);
nor U5075 (N_5075,N_4850,N_4712);
nor U5076 (N_5076,N_4611,N_4945);
nand U5077 (N_5077,N_4742,N_4708);
or U5078 (N_5078,N_4977,N_4624);
and U5079 (N_5079,N_4563,N_4526);
or U5080 (N_5080,N_4784,N_4988);
or U5081 (N_5081,N_4843,N_4758);
or U5082 (N_5082,N_4627,N_4658);
nand U5083 (N_5083,N_4838,N_4671);
and U5084 (N_5084,N_4679,N_4585);
nand U5085 (N_5085,N_4752,N_4966);
or U5086 (N_5086,N_4791,N_4702);
xnor U5087 (N_5087,N_4864,N_4806);
nor U5088 (N_5088,N_4794,N_4961);
xor U5089 (N_5089,N_4564,N_4881);
nand U5090 (N_5090,N_4700,N_4729);
and U5091 (N_5091,N_4555,N_4594);
xor U5092 (N_5092,N_4673,N_4688);
and U5093 (N_5093,N_4536,N_4935);
nand U5094 (N_5094,N_4931,N_4999);
or U5095 (N_5095,N_4882,N_4623);
xnor U5096 (N_5096,N_4920,N_4654);
or U5097 (N_5097,N_4912,N_4574);
nand U5098 (N_5098,N_4835,N_4734);
nand U5099 (N_5099,N_4570,N_4777);
xnor U5100 (N_5100,N_4583,N_4980);
or U5101 (N_5101,N_4567,N_4532);
nand U5102 (N_5102,N_4608,N_4746);
nand U5103 (N_5103,N_4634,N_4901);
nand U5104 (N_5104,N_4670,N_4875);
and U5105 (N_5105,N_4891,N_4580);
nand U5106 (N_5106,N_4540,N_4750);
xnor U5107 (N_5107,N_4506,N_4595);
nor U5108 (N_5108,N_4907,N_4754);
and U5109 (N_5109,N_4860,N_4696);
nand U5110 (N_5110,N_4845,N_4925);
xor U5111 (N_5111,N_4727,N_4863);
xor U5112 (N_5112,N_4755,N_4512);
and U5113 (N_5113,N_4584,N_4759);
and U5114 (N_5114,N_4668,N_4677);
and U5115 (N_5115,N_4869,N_4549);
nor U5116 (N_5116,N_4964,N_4958);
xor U5117 (N_5117,N_4657,N_4972);
nand U5118 (N_5118,N_4622,N_4689);
nand U5119 (N_5119,N_4517,N_4723);
or U5120 (N_5120,N_4782,N_4975);
or U5121 (N_5121,N_4896,N_4844);
nor U5122 (N_5122,N_4743,N_4947);
xnor U5123 (N_5123,N_4938,N_4909);
or U5124 (N_5124,N_4796,N_4842);
nor U5125 (N_5125,N_4870,N_4765);
nand U5126 (N_5126,N_4762,N_4691);
nand U5127 (N_5127,N_4974,N_4534);
and U5128 (N_5128,N_4543,N_4582);
nand U5129 (N_5129,N_4899,N_4538);
xor U5130 (N_5130,N_4698,N_4820);
or U5131 (N_5131,N_4824,N_4978);
and U5132 (N_5132,N_4736,N_4804);
or U5133 (N_5133,N_4883,N_4941);
nand U5134 (N_5134,N_4731,N_4663);
or U5135 (N_5135,N_4878,N_4886);
nand U5136 (N_5136,N_4726,N_4771);
and U5137 (N_5137,N_4616,N_4812);
and U5138 (N_5138,N_4959,N_4792);
or U5139 (N_5139,N_4787,N_4809);
nand U5140 (N_5140,N_4800,N_4644);
or U5141 (N_5141,N_4572,N_4528);
nor U5142 (N_5142,N_4544,N_4910);
nand U5143 (N_5143,N_4789,N_4873);
nand U5144 (N_5144,N_4950,N_4954);
and U5145 (N_5145,N_4699,N_4871);
xnor U5146 (N_5146,N_4607,N_4525);
nor U5147 (N_5147,N_4790,N_4600);
or U5148 (N_5148,N_4550,N_4865);
xnor U5149 (N_5149,N_4857,N_4515);
nor U5150 (N_5150,N_4744,N_4615);
and U5151 (N_5151,N_4880,N_4919);
or U5152 (N_5152,N_4846,N_4519);
xnor U5153 (N_5153,N_4922,N_4718);
nor U5154 (N_5154,N_4946,N_4523);
nor U5155 (N_5155,N_4953,N_4900);
nor U5156 (N_5156,N_4606,N_4940);
and U5157 (N_5157,N_4638,N_4659);
and U5158 (N_5158,N_4686,N_4695);
or U5159 (N_5159,N_4867,N_4617);
nor U5160 (N_5160,N_4591,N_4505);
xor U5161 (N_5161,N_4587,N_4566);
nor U5162 (N_5162,N_4711,N_4763);
nor U5163 (N_5163,N_4769,N_4956);
nand U5164 (N_5164,N_4785,N_4803);
or U5165 (N_5165,N_4944,N_4969);
or U5166 (N_5166,N_4559,N_4510);
xnor U5167 (N_5167,N_4605,N_4851);
or U5168 (N_5168,N_4770,N_4775);
nor U5169 (N_5169,N_4545,N_4852);
xor U5170 (N_5170,N_4631,N_4604);
and U5171 (N_5171,N_4704,N_4716);
or U5172 (N_5172,N_4577,N_4766);
xor U5173 (N_5173,N_4546,N_4568);
or U5174 (N_5174,N_4665,N_4913);
nor U5175 (N_5175,N_4949,N_4993);
nor U5176 (N_5176,N_4522,N_4924);
nand U5177 (N_5177,N_4906,N_4508);
and U5178 (N_5178,N_4651,N_4916);
and U5179 (N_5179,N_4715,N_4829);
xor U5180 (N_5180,N_4660,N_4575);
or U5181 (N_5181,N_4586,N_4621);
or U5182 (N_5182,N_4581,N_4648);
and U5183 (N_5183,N_4745,N_4630);
and U5184 (N_5184,N_4576,N_4633);
nor U5185 (N_5185,N_4637,N_4682);
and U5186 (N_5186,N_4902,N_4866);
or U5187 (N_5187,N_4884,N_4894);
nand U5188 (N_5188,N_4504,N_4915);
xor U5189 (N_5189,N_4847,N_4767);
or U5190 (N_5190,N_4646,N_4507);
nand U5191 (N_5191,N_4539,N_4970);
nand U5192 (N_5192,N_4535,N_4558);
and U5193 (N_5193,N_4813,N_4991);
or U5194 (N_5194,N_4831,N_4636);
nor U5195 (N_5195,N_4816,N_4748);
or U5196 (N_5196,N_4641,N_4879);
or U5197 (N_5197,N_4732,N_4516);
nor U5198 (N_5198,N_4840,N_4518);
nor U5199 (N_5199,N_4687,N_4951);
or U5200 (N_5200,N_4537,N_4513);
and U5201 (N_5201,N_4524,N_4547);
nor U5202 (N_5202,N_4968,N_4849);
nor U5203 (N_5203,N_4985,N_4728);
nor U5204 (N_5204,N_4625,N_4511);
xor U5205 (N_5205,N_4937,N_4738);
nor U5206 (N_5206,N_4579,N_4987);
xor U5207 (N_5207,N_4888,N_4741);
xnor U5208 (N_5208,N_4996,N_4614);
nor U5209 (N_5209,N_4757,N_4853);
and U5210 (N_5210,N_4640,N_4905);
and U5211 (N_5211,N_4892,N_4593);
xor U5212 (N_5212,N_4672,N_4983);
xnor U5213 (N_5213,N_4986,N_4854);
nor U5214 (N_5214,N_4557,N_4795);
nor U5215 (N_5215,N_4740,N_4990);
xor U5216 (N_5216,N_4797,N_4642);
or U5217 (N_5217,N_4955,N_4917);
xnor U5218 (N_5218,N_4783,N_4722);
xnor U5219 (N_5219,N_4533,N_4626);
and U5220 (N_5220,N_4825,N_4502);
xnor U5221 (N_5221,N_4685,N_4562);
or U5222 (N_5222,N_4602,N_4612);
nand U5223 (N_5223,N_4994,N_4632);
nand U5224 (N_5224,N_4650,N_4514);
nand U5225 (N_5225,N_4751,N_4683);
nand U5226 (N_5226,N_4973,N_4509);
nor U5227 (N_5227,N_4918,N_4588);
or U5228 (N_5228,N_4597,N_4963);
xnor U5229 (N_5229,N_4618,N_4893);
nor U5230 (N_5230,N_4619,N_4694);
nand U5231 (N_5231,N_4565,N_4503);
xnor U5232 (N_5232,N_4821,N_4603);
xor U5233 (N_5233,N_4861,N_4927);
nor U5234 (N_5234,N_4556,N_4817);
nor U5235 (N_5235,N_4930,N_4656);
xor U5236 (N_5236,N_4781,N_4664);
xor U5237 (N_5237,N_4678,N_4747);
or U5238 (N_5238,N_4707,N_4548);
nor U5239 (N_5239,N_4989,N_4629);
or U5240 (N_5240,N_4929,N_4669);
nand U5241 (N_5241,N_4826,N_4693);
xor U5242 (N_5242,N_4578,N_4788);
xor U5243 (N_5243,N_4676,N_4773);
nor U5244 (N_5244,N_4710,N_4943);
nand U5245 (N_5245,N_4653,N_4589);
and U5246 (N_5246,N_4832,N_4903);
and U5247 (N_5247,N_4542,N_4834);
nand U5248 (N_5248,N_4774,N_4598);
xor U5249 (N_5249,N_4981,N_4620);
and U5250 (N_5250,N_4971,N_4586);
and U5251 (N_5251,N_4969,N_4546);
or U5252 (N_5252,N_4626,N_4897);
nor U5253 (N_5253,N_4958,N_4733);
xnor U5254 (N_5254,N_4879,N_4529);
or U5255 (N_5255,N_4526,N_4578);
xnor U5256 (N_5256,N_4770,N_4709);
nand U5257 (N_5257,N_4915,N_4862);
xnor U5258 (N_5258,N_4727,N_4818);
nand U5259 (N_5259,N_4765,N_4947);
xnor U5260 (N_5260,N_4726,N_4625);
nand U5261 (N_5261,N_4912,N_4559);
nor U5262 (N_5262,N_4570,N_4697);
nor U5263 (N_5263,N_4857,N_4972);
nand U5264 (N_5264,N_4914,N_4556);
nor U5265 (N_5265,N_4677,N_4763);
xor U5266 (N_5266,N_4512,N_4542);
nand U5267 (N_5267,N_4714,N_4853);
xnor U5268 (N_5268,N_4774,N_4757);
and U5269 (N_5269,N_4674,N_4864);
nand U5270 (N_5270,N_4711,N_4629);
or U5271 (N_5271,N_4512,N_4607);
or U5272 (N_5272,N_4704,N_4665);
xor U5273 (N_5273,N_4534,N_4978);
or U5274 (N_5274,N_4973,N_4682);
xor U5275 (N_5275,N_4539,N_4929);
nor U5276 (N_5276,N_4686,N_4711);
nand U5277 (N_5277,N_4844,N_4855);
xor U5278 (N_5278,N_4537,N_4931);
nor U5279 (N_5279,N_4903,N_4555);
nor U5280 (N_5280,N_4524,N_4551);
or U5281 (N_5281,N_4740,N_4604);
nor U5282 (N_5282,N_4875,N_4609);
xnor U5283 (N_5283,N_4522,N_4877);
xor U5284 (N_5284,N_4522,N_4965);
nand U5285 (N_5285,N_4881,N_4917);
and U5286 (N_5286,N_4746,N_4520);
nand U5287 (N_5287,N_4713,N_4837);
and U5288 (N_5288,N_4622,N_4939);
nor U5289 (N_5289,N_4513,N_4659);
or U5290 (N_5290,N_4786,N_4541);
or U5291 (N_5291,N_4539,N_4861);
nor U5292 (N_5292,N_4978,N_4868);
and U5293 (N_5293,N_4969,N_4773);
xor U5294 (N_5294,N_4893,N_4850);
or U5295 (N_5295,N_4573,N_4727);
xor U5296 (N_5296,N_4779,N_4937);
or U5297 (N_5297,N_4887,N_4574);
xor U5298 (N_5298,N_4713,N_4666);
or U5299 (N_5299,N_4720,N_4705);
xnor U5300 (N_5300,N_4617,N_4994);
and U5301 (N_5301,N_4935,N_4867);
and U5302 (N_5302,N_4877,N_4680);
xor U5303 (N_5303,N_4717,N_4552);
nand U5304 (N_5304,N_4534,N_4940);
and U5305 (N_5305,N_4608,N_4752);
nand U5306 (N_5306,N_4947,N_4615);
nand U5307 (N_5307,N_4937,N_4853);
nand U5308 (N_5308,N_4793,N_4946);
xor U5309 (N_5309,N_4566,N_4871);
and U5310 (N_5310,N_4743,N_4944);
nand U5311 (N_5311,N_4519,N_4722);
and U5312 (N_5312,N_4931,N_4937);
or U5313 (N_5313,N_4896,N_4923);
nand U5314 (N_5314,N_4926,N_4915);
nand U5315 (N_5315,N_4758,N_4542);
nor U5316 (N_5316,N_4802,N_4938);
and U5317 (N_5317,N_4548,N_4642);
and U5318 (N_5318,N_4542,N_4725);
or U5319 (N_5319,N_4597,N_4919);
nor U5320 (N_5320,N_4595,N_4957);
and U5321 (N_5321,N_4992,N_4529);
or U5322 (N_5322,N_4550,N_4721);
and U5323 (N_5323,N_4778,N_4687);
nor U5324 (N_5324,N_4773,N_4991);
and U5325 (N_5325,N_4703,N_4998);
nand U5326 (N_5326,N_4828,N_4678);
nor U5327 (N_5327,N_4829,N_4810);
nor U5328 (N_5328,N_4608,N_4969);
or U5329 (N_5329,N_4564,N_4704);
xnor U5330 (N_5330,N_4711,N_4513);
xor U5331 (N_5331,N_4897,N_4542);
or U5332 (N_5332,N_4619,N_4775);
nor U5333 (N_5333,N_4648,N_4568);
nand U5334 (N_5334,N_4625,N_4633);
xor U5335 (N_5335,N_4679,N_4617);
or U5336 (N_5336,N_4854,N_4849);
xnor U5337 (N_5337,N_4765,N_4666);
and U5338 (N_5338,N_4673,N_4775);
nor U5339 (N_5339,N_4789,N_4857);
xor U5340 (N_5340,N_4927,N_4694);
or U5341 (N_5341,N_4790,N_4989);
nor U5342 (N_5342,N_4562,N_4721);
and U5343 (N_5343,N_4938,N_4554);
and U5344 (N_5344,N_4743,N_4750);
or U5345 (N_5345,N_4905,N_4509);
xor U5346 (N_5346,N_4587,N_4542);
xor U5347 (N_5347,N_4976,N_4516);
nand U5348 (N_5348,N_4795,N_4909);
or U5349 (N_5349,N_4505,N_4841);
nand U5350 (N_5350,N_4723,N_4671);
nand U5351 (N_5351,N_4548,N_4522);
and U5352 (N_5352,N_4673,N_4653);
nor U5353 (N_5353,N_4970,N_4860);
and U5354 (N_5354,N_4590,N_4638);
and U5355 (N_5355,N_4870,N_4590);
nand U5356 (N_5356,N_4711,N_4823);
nor U5357 (N_5357,N_4848,N_4940);
nand U5358 (N_5358,N_4985,N_4665);
nor U5359 (N_5359,N_4640,N_4926);
xnor U5360 (N_5360,N_4742,N_4925);
nand U5361 (N_5361,N_4547,N_4666);
xnor U5362 (N_5362,N_4656,N_4727);
xor U5363 (N_5363,N_4575,N_4795);
xnor U5364 (N_5364,N_4754,N_4782);
xor U5365 (N_5365,N_4585,N_4826);
nor U5366 (N_5366,N_4771,N_4791);
nor U5367 (N_5367,N_4527,N_4865);
and U5368 (N_5368,N_4638,N_4885);
xnor U5369 (N_5369,N_4821,N_4549);
nor U5370 (N_5370,N_4838,N_4943);
xor U5371 (N_5371,N_4660,N_4598);
xor U5372 (N_5372,N_4587,N_4947);
nor U5373 (N_5373,N_4922,N_4845);
and U5374 (N_5374,N_4863,N_4685);
or U5375 (N_5375,N_4797,N_4548);
or U5376 (N_5376,N_4688,N_4992);
and U5377 (N_5377,N_4521,N_4586);
nand U5378 (N_5378,N_4541,N_4771);
or U5379 (N_5379,N_4719,N_4522);
and U5380 (N_5380,N_4799,N_4547);
and U5381 (N_5381,N_4588,N_4561);
xnor U5382 (N_5382,N_4912,N_4682);
nor U5383 (N_5383,N_4742,N_4662);
and U5384 (N_5384,N_4985,N_4850);
and U5385 (N_5385,N_4920,N_4839);
xor U5386 (N_5386,N_4996,N_4795);
nor U5387 (N_5387,N_4667,N_4810);
xor U5388 (N_5388,N_4801,N_4912);
nor U5389 (N_5389,N_4683,N_4846);
xor U5390 (N_5390,N_4630,N_4907);
nor U5391 (N_5391,N_4736,N_4655);
and U5392 (N_5392,N_4798,N_4915);
nand U5393 (N_5393,N_4741,N_4966);
or U5394 (N_5394,N_4780,N_4834);
nor U5395 (N_5395,N_4733,N_4604);
nor U5396 (N_5396,N_4795,N_4876);
or U5397 (N_5397,N_4727,N_4699);
nand U5398 (N_5398,N_4878,N_4725);
and U5399 (N_5399,N_4890,N_4634);
xnor U5400 (N_5400,N_4554,N_4668);
nand U5401 (N_5401,N_4681,N_4558);
nor U5402 (N_5402,N_4763,N_4846);
or U5403 (N_5403,N_4760,N_4741);
xnor U5404 (N_5404,N_4565,N_4659);
and U5405 (N_5405,N_4748,N_4940);
nor U5406 (N_5406,N_4549,N_4591);
nand U5407 (N_5407,N_4550,N_4989);
nor U5408 (N_5408,N_4781,N_4842);
and U5409 (N_5409,N_4939,N_4637);
and U5410 (N_5410,N_4506,N_4608);
nand U5411 (N_5411,N_4767,N_4875);
nor U5412 (N_5412,N_4948,N_4616);
nand U5413 (N_5413,N_4869,N_4833);
and U5414 (N_5414,N_4502,N_4522);
xor U5415 (N_5415,N_4884,N_4897);
or U5416 (N_5416,N_4845,N_4755);
nor U5417 (N_5417,N_4896,N_4736);
nor U5418 (N_5418,N_4939,N_4549);
nor U5419 (N_5419,N_4702,N_4642);
nor U5420 (N_5420,N_4875,N_4898);
nand U5421 (N_5421,N_4803,N_4840);
nand U5422 (N_5422,N_4686,N_4698);
or U5423 (N_5423,N_4766,N_4758);
nor U5424 (N_5424,N_4940,N_4942);
and U5425 (N_5425,N_4910,N_4707);
or U5426 (N_5426,N_4763,N_4506);
and U5427 (N_5427,N_4999,N_4850);
nor U5428 (N_5428,N_4598,N_4667);
nand U5429 (N_5429,N_4820,N_4552);
or U5430 (N_5430,N_4684,N_4946);
xnor U5431 (N_5431,N_4663,N_4544);
nand U5432 (N_5432,N_4905,N_4802);
nand U5433 (N_5433,N_4545,N_4645);
xnor U5434 (N_5434,N_4537,N_4573);
nor U5435 (N_5435,N_4852,N_4854);
and U5436 (N_5436,N_4514,N_4798);
nand U5437 (N_5437,N_4697,N_4716);
or U5438 (N_5438,N_4809,N_4924);
nand U5439 (N_5439,N_4956,N_4610);
nand U5440 (N_5440,N_4761,N_4552);
and U5441 (N_5441,N_4947,N_4734);
xor U5442 (N_5442,N_4514,N_4925);
nand U5443 (N_5443,N_4937,N_4818);
or U5444 (N_5444,N_4540,N_4906);
xnor U5445 (N_5445,N_4899,N_4512);
xor U5446 (N_5446,N_4619,N_4998);
xnor U5447 (N_5447,N_4761,N_4553);
nor U5448 (N_5448,N_4869,N_4779);
xnor U5449 (N_5449,N_4655,N_4913);
nand U5450 (N_5450,N_4704,N_4785);
xor U5451 (N_5451,N_4561,N_4587);
xor U5452 (N_5452,N_4733,N_4672);
nand U5453 (N_5453,N_4828,N_4622);
xor U5454 (N_5454,N_4576,N_4614);
nor U5455 (N_5455,N_4737,N_4867);
nor U5456 (N_5456,N_4887,N_4946);
or U5457 (N_5457,N_4517,N_4870);
nand U5458 (N_5458,N_4595,N_4623);
nand U5459 (N_5459,N_4902,N_4862);
nor U5460 (N_5460,N_4844,N_4547);
xnor U5461 (N_5461,N_4937,N_4500);
xor U5462 (N_5462,N_4780,N_4618);
xnor U5463 (N_5463,N_4842,N_4728);
and U5464 (N_5464,N_4945,N_4800);
xnor U5465 (N_5465,N_4980,N_4687);
and U5466 (N_5466,N_4705,N_4972);
and U5467 (N_5467,N_4659,N_4954);
nor U5468 (N_5468,N_4675,N_4662);
and U5469 (N_5469,N_4501,N_4922);
xnor U5470 (N_5470,N_4883,N_4971);
nor U5471 (N_5471,N_4733,N_4803);
xor U5472 (N_5472,N_4908,N_4569);
and U5473 (N_5473,N_4923,N_4869);
nor U5474 (N_5474,N_4720,N_4781);
xnor U5475 (N_5475,N_4618,N_4678);
and U5476 (N_5476,N_4877,N_4972);
and U5477 (N_5477,N_4691,N_4954);
and U5478 (N_5478,N_4638,N_4923);
and U5479 (N_5479,N_4943,N_4777);
nor U5480 (N_5480,N_4635,N_4945);
nand U5481 (N_5481,N_4714,N_4583);
or U5482 (N_5482,N_4890,N_4707);
nor U5483 (N_5483,N_4728,N_4598);
or U5484 (N_5484,N_4644,N_4919);
or U5485 (N_5485,N_4582,N_4951);
nor U5486 (N_5486,N_4975,N_4991);
nor U5487 (N_5487,N_4893,N_4667);
or U5488 (N_5488,N_4839,N_4902);
or U5489 (N_5489,N_4914,N_4639);
nor U5490 (N_5490,N_4646,N_4891);
nand U5491 (N_5491,N_4523,N_4824);
and U5492 (N_5492,N_4929,N_4553);
and U5493 (N_5493,N_4718,N_4940);
and U5494 (N_5494,N_4930,N_4781);
or U5495 (N_5495,N_4747,N_4832);
and U5496 (N_5496,N_4760,N_4703);
xor U5497 (N_5497,N_4983,N_4836);
xor U5498 (N_5498,N_4500,N_4680);
and U5499 (N_5499,N_4693,N_4989);
xnor U5500 (N_5500,N_5090,N_5250);
nand U5501 (N_5501,N_5007,N_5378);
or U5502 (N_5502,N_5211,N_5222);
nor U5503 (N_5503,N_5472,N_5372);
or U5504 (N_5504,N_5315,N_5075);
and U5505 (N_5505,N_5328,N_5413);
nor U5506 (N_5506,N_5411,N_5246);
or U5507 (N_5507,N_5135,N_5052);
and U5508 (N_5508,N_5420,N_5095);
or U5509 (N_5509,N_5055,N_5051);
or U5510 (N_5510,N_5048,N_5039);
xor U5511 (N_5511,N_5253,N_5321);
and U5512 (N_5512,N_5174,N_5395);
nand U5513 (N_5513,N_5412,N_5102);
nand U5514 (N_5514,N_5429,N_5162);
and U5515 (N_5515,N_5088,N_5049);
xor U5516 (N_5516,N_5282,N_5063);
and U5517 (N_5517,N_5004,N_5151);
or U5518 (N_5518,N_5340,N_5020);
or U5519 (N_5519,N_5379,N_5115);
xnor U5520 (N_5520,N_5225,N_5233);
nand U5521 (N_5521,N_5193,N_5139);
nor U5522 (N_5522,N_5251,N_5281);
or U5523 (N_5523,N_5147,N_5261);
nand U5524 (N_5524,N_5138,N_5334);
or U5525 (N_5525,N_5118,N_5122);
and U5526 (N_5526,N_5214,N_5346);
nor U5527 (N_5527,N_5305,N_5414);
xor U5528 (N_5528,N_5476,N_5309);
nand U5529 (N_5529,N_5169,N_5084);
xor U5530 (N_5530,N_5178,N_5053);
or U5531 (N_5531,N_5080,N_5215);
nand U5532 (N_5532,N_5175,N_5109);
nor U5533 (N_5533,N_5184,N_5245);
nand U5534 (N_5534,N_5078,N_5360);
xor U5535 (N_5535,N_5207,N_5304);
nand U5536 (N_5536,N_5392,N_5074);
nor U5537 (N_5537,N_5449,N_5436);
or U5538 (N_5538,N_5066,N_5212);
nor U5539 (N_5539,N_5432,N_5000);
nor U5540 (N_5540,N_5418,N_5177);
or U5541 (N_5541,N_5168,N_5110);
xor U5542 (N_5542,N_5355,N_5032);
or U5543 (N_5543,N_5114,N_5462);
nand U5544 (N_5544,N_5031,N_5489);
xnor U5545 (N_5545,N_5479,N_5111);
and U5546 (N_5546,N_5023,N_5042);
nand U5547 (N_5547,N_5314,N_5240);
nor U5548 (N_5548,N_5347,N_5339);
xor U5549 (N_5549,N_5009,N_5033);
or U5550 (N_5550,N_5142,N_5167);
or U5551 (N_5551,N_5450,N_5461);
nand U5552 (N_5552,N_5201,N_5179);
nand U5553 (N_5553,N_5335,N_5438);
and U5554 (N_5554,N_5493,N_5308);
xor U5555 (N_5555,N_5025,N_5386);
and U5556 (N_5556,N_5083,N_5017);
xor U5557 (N_5557,N_5137,N_5202);
and U5558 (N_5558,N_5027,N_5481);
or U5559 (N_5559,N_5243,N_5124);
xnor U5560 (N_5560,N_5037,N_5041);
nor U5561 (N_5561,N_5230,N_5359);
xor U5562 (N_5562,N_5036,N_5463);
nand U5563 (N_5563,N_5047,N_5297);
nand U5564 (N_5564,N_5043,N_5464);
and U5565 (N_5565,N_5030,N_5403);
and U5566 (N_5566,N_5430,N_5157);
nor U5567 (N_5567,N_5192,N_5389);
nand U5568 (N_5568,N_5387,N_5331);
xor U5569 (N_5569,N_5302,N_5380);
and U5570 (N_5570,N_5097,N_5272);
or U5571 (N_5571,N_5426,N_5185);
or U5572 (N_5572,N_5236,N_5100);
or U5573 (N_5573,N_5393,N_5356);
nor U5574 (N_5574,N_5105,N_5241);
and U5575 (N_5575,N_5363,N_5330);
and U5576 (N_5576,N_5350,N_5265);
and U5577 (N_5577,N_5087,N_5498);
nand U5578 (N_5578,N_5399,N_5307);
or U5579 (N_5579,N_5401,N_5150);
xor U5580 (N_5580,N_5348,N_5040);
nor U5581 (N_5581,N_5451,N_5434);
or U5582 (N_5582,N_5235,N_5373);
nor U5583 (N_5583,N_5466,N_5285);
and U5584 (N_5584,N_5491,N_5024);
xnor U5585 (N_5585,N_5271,N_5322);
and U5586 (N_5586,N_5164,N_5216);
nand U5587 (N_5587,N_5034,N_5270);
and U5588 (N_5588,N_5086,N_5312);
nor U5589 (N_5589,N_5146,N_5370);
nor U5590 (N_5590,N_5351,N_5259);
or U5591 (N_5591,N_5148,N_5054);
nor U5592 (N_5592,N_5345,N_5364);
xor U5593 (N_5593,N_5467,N_5155);
xnor U5594 (N_5594,N_5226,N_5209);
xnor U5595 (N_5595,N_5064,N_5490);
xor U5596 (N_5596,N_5289,N_5311);
or U5597 (N_5597,N_5070,N_5424);
or U5598 (N_5598,N_5077,N_5447);
and U5599 (N_5599,N_5495,N_5190);
nor U5600 (N_5600,N_5059,N_5362);
nand U5601 (N_5601,N_5484,N_5208);
or U5602 (N_5602,N_5385,N_5093);
and U5603 (N_5603,N_5057,N_5357);
or U5604 (N_5604,N_5197,N_5329);
and U5605 (N_5605,N_5455,N_5152);
xor U5606 (N_5606,N_5213,N_5191);
and U5607 (N_5607,N_5431,N_5267);
nand U5608 (N_5608,N_5354,N_5407);
or U5609 (N_5609,N_5323,N_5170);
xor U5610 (N_5610,N_5256,N_5288);
or U5611 (N_5611,N_5003,N_5200);
and U5612 (N_5612,N_5283,N_5195);
and U5613 (N_5613,N_5268,N_5465);
xnor U5614 (N_5614,N_5013,N_5113);
nor U5615 (N_5615,N_5158,N_5428);
and U5616 (N_5616,N_5448,N_5296);
or U5617 (N_5617,N_5341,N_5486);
and U5618 (N_5618,N_5189,N_5306);
xnor U5619 (N_5619,N_5327,N_5408);
or U5620 (N_5620,N_5249,N_5182);
nand U5621 (N_5621,N_5478,N_5210);
nor U5622 (N_5622,N_5018,N_5482);
or U5623 (N_5623,N_5145,N_5494);
xnor U5624 (N_5624,N_5497,N_5483);
nand U5625 (N_5625,N_5369,N_5130);
nor U5626 (N_5626,N_5276,N_5287);
and U5627 (N_5627,N_5273,N_5459);
nor U5628 (N_5628,N_5358,N_5325);
and U5629 (N_5629,N_5284,N_5433);
nand U5630 (N_5630,N_5224,N_5120);
xor U5631 (N_5631,N_5166,N_5026);
nor U5632 (N_5632,N_5223,N_5444);
and U5633 (N_5633,N_5487,N_5353);
nor U5634 (N_5634,N_5133,N_5238);
or U5635 (N_5635,N_5390,N_5143);
nand U5636 (N_5636,N_5458,N_5320);
nand U5637 (N_5637,N_5313,N_5452);
and U5638 (N_5638,N_5473,N_5128);
or U5639 (N_5639,N_5028,N_5468);
or U5640 (N_5640,N_5252,N_5469);
and U5641 (N_5641,N_5263,N_5257);
or U5642 (N_5642,N_5376,N_5293);
xor U5643 (N_5643,N_5094,N_5286);
nor U5644 (N_5644,N_5422,N_5069);
nand U5645 (N_5645,N_5262,N_5480);
nand U5646 (N_5646,N_5199,N_5269);
nor U5647 (N_5647,N_5406,N_5391);
or U5648 (N_5648,N_5485,N_5300);
nand U5649 (N_5649,N_5035,N_5014);
or U5650 (N_5650,N_5384,N_5126);
or U5651 (N_5651,N_5132,N_5475);
or U5652 (N_5652,N_5220,N_5474);
nor U5653 (N_5653,N_5344,N_5388);
and U5654 (N_5654,N_5471,N_5046);
or U5655 (N_5655,N_5136,N_5439);
and U5656 (N_5656,N_5073,N_5010);
and U5657 (N_5657,N_5092,N_5125);
xor U5658 (N_5658,N_5409,N_5274);
and U5659 (N_5659,N_5044,N_5006);
nand U5660 (N_5660,N_5237,N_5375);
or U5661 (N_5661,N_5280,N_5361);
and U5662 (N_5662,N_5317,N_5396);
nand U5663 (N_5663,N_5368,N_5012);
nor U5664 (N_5664,N_5154,N_5050);
nor U5665 (N_5665,N_5333,N_5324);
nor U5666 (N_5666,N_5453,N_5203);
xor U5667 (N_5667,N_5338,N_5415);
xnor U5668 (N_5668,N_5127,N_5398);
or U5669 (N_5669,N_5319,N_5255);
or U5670 (N_5670,N_5460,N_5076);
nand U5671 (N_5671,N_5266,N_5183);
and U5672 (N_5672,N_5492,N_5163);
or U5673 (N_5673,N_5247,N_5374);
or U5674 (N_5674,N_5310,N_5254);
and U5675 (N_5675,N_5228,N_5291);
or U5676 (N_5676,N_5275,N_5103);
and U5677 (N_5677,N_5081,N_5499);
nor U5678 (N_5678,N_5290,N_5316);
or U5679 (N_5679,N_5365,N_5058);
and U5680 (N_5680,N_5352,N_5045);
xnor U5681 (N_5681,N_5336,N_5419);
and U5682 (N_5682,N_5221,N_5104);
nor U5683 (N_5683,N_5258,N_5421);
nand U5684 (N_5684,N_5021,N_5425);
or U5685 (N_5685,N_5457,N_5488);
nand U5686 (N_5686,N_5101,N_5377);
nand U5687 (N_5687,N_5405,N_5106);
nand U5688 (N_5688,N_5496,N_5180);
and U5689 (N_5689,N_5065,N_5382);
nand U5690 (N_5690,N_5061,N_5068);
nor U5691 (N_5691,N_5016,N_5298);
or U5692 (N_5692,N_5062,N_5441);
nand U5693 (N_5693,N_5292,N_5349);
nand U5694 (N_5694,N_5056,N_5244);
nor U5695 (N_5695,N_5091,N_5402);
or U5696 (N_5696,N_5108,N_5446);
nand U5697 (N_5697,N_5187,N_5165);
nor U5698 (N_5698,N_5144,N_5117);
nand U5699 (N_5699,N_5089,N_5008);
nand U5700 (N_5700,N_5219,N_5015);
xor U5701 (N_5701,N_5326,N_5159);
nor U5702 (N_5702,N_5248,N_5440);
nor U5703 (N_5703,N_5022,N_5129);
and U5704 (N_5704,N_5002,N_5301);
xnor U5705 (N_5705,N_5227,N_5140);
nand U5706 (N_5706,N_5295,N_5299);
xnor U5707 (N_5707,N_5218,N_5205);
and U5708 (N_5708,N_5367,N_5071);
and U5709 (N_5709,N_5161,N_5067);
and U5710 (N_5710,N_5204,N_5029);
or U5711 (N_5711,N_5303,N_5371);
or U5712 (N_5712,N_5239,N_5383);
xnor U5713 (N_5713,N_5435,N_5096);
and U5714 (N_5714,N_5477,N_5232);
and U5715 (N_5715,N_5381,N_5242);
xnor U5716 (N_5716,N_5149,N_5141);
xnor U5717 (N_5717,N_5264,N_5160);
or U5718 (N_5718,N_5427,N_5131);
and U5719 (N_5719,N_5229,N_5337);
or U5720 (N_5720,N_5005,N_5366);
or U5721 (N_5721,N_5343,N_5456);
nand U5722 (N_5722,N_5417,N_5176);
or U5723 (N_5723,N_5318,N_5279);
and U5724 (N_5724,N_5134,N_5198);
or U5725 (N_5725,N_5196,N_5173);
xor U5726 (N_5726,N_5085,N_5112);
or U5727 (N_5727,N_5231,N_5019);
and U5728 (N_5728,N_5001,N_5437);
xor U5729 (N_5729,N_5206,N_5107);
nand U5730 (N_5730,N_5172,N_5153);
xnor U5731 (N_5731,N_5397,N_5400);
xor U5732 (N_5732,N_5294,N_5260);
nor U5733 (N_5733,N_5443,N_5060);
or U5734 (N_5734,N_5416,N_5194);
nand U5735 (N_5735,N_5011,N_5186);
and U5736 (N_5736,N_5470,N_5079);
or U5737 (N_5737,N_5454,N_5082);
xor U5738 (N_5738,N_5171,N_5072);
nand U5739 (N_5739,N_5119,N_5278);
nand U5740 (N_5740,N_5217,N_5277);
and U5741 (N_5741,N_5121,N_5342);
nand U5742 (N_5742,N_5445,N_5123);
nand U5743 (N_5743,N_5181,N_5234);
and U5744 (N_5744,N_5332,N_5156);
or U5745 (N_5745,N_5410,N_5098);
xnor U5746 (N_5746,N_5423,N_5442);
xor U5747 (N_5747,N_5404,N_5099);
and U5748 (N_5748,N_5116,N_5188);
xnor U5749 (N_5749,N_5394,N_5038);
and U5750 (N_5750,N_5107,N_5175);
nand U5751 (N_5751,N_5070,N_5165);
or U5752 (N_5752,N_5425,N_5432);
or U5753 (N_5753,N_5185,N_5334);
nand U5754 (N_5754,N_5234,N_5136);
and U5755 (N_5755,N_5055,N_5366);
xnor U5756 (N_5756,N_5050,N_5131);
xor U5757 (N_5757,N_5387,N_5016);
or U5758 (N_5758,N_5439,N_5455);
nand U5759 (N_5759,N_5313,N_5426);
nand U5760 (N_5760,N_5208,N_5350);
or U5761 (N_5761,N_5098,N_5356);
and U5762 (N_5762,N_5153,N_5035);
or U5763 (N_5763,N_5149,N_5409);
xor U5764 (N_5764,N_5346,N_5370);
nor U5765 (N_5765,N_5016,N_5166);
and U5766 (N_5766,N_5075,N_5461);
and U5767 (N_5767,N_5488,N_5472);
xnor U5768 (N_5768,N_5005,N_5441);
nand U5769 (N_5769,N_5168,N_5488);
nor U5770 (N_5770,N_5404,N_5085);
or U5771 (N_5771,N_5325,N_5330);
and U5772 (N_5772,N_5207,N_5365);
and U5773 (N_5773,N_5397,N_5280);
nor U5774 (N_5774,N_5258,N_5206);
and U5775 (N_5775,N_5287,N_5213);
and U5776 (N_5776,N_5438,N_5307);
xor U5777 (N_5777,N_5468,N_5247);
nor U5778 (N_5778,N_5252,N_5345);
nand U5779 (N_5779,N_5275,N_5296);
and U5780 (N_5780,N_5199,N_5419);
xor U5781 (N_5781,N_5285,N_5362);
and U5782 (N_5782,N_5272,N_5011);
or U5783 (N_5783,N_5313,N_5036);
nor U5784 (N_5784,N_5316,N_5312);
nor U5785 (N_5785,N_5139,N_5486);
nor U5786 (N_5786,N_5198,N_5210);
and U5787 (N_5787,N_5001,N_5285);
nand U5788 (N_5788,N_5404,N_5241);
nand U5789 (N_5789,N_5306,N_5330);
and U5790 (N_5790,N_5468,N_5332);
xor U5791 (N_5791,N_5017,N_5253);
or U5792 (N_5792,N_5000,N_5256);
and U5793 (N_5793,N_5095,N_5388);
and U5794 (N_5794,N_5034,N_5085);
nand U5795 (N_5795,N_5374,N_5194);
xor U5796 (N_5796,N_5157,N_5079);
xnor U5797 (N_5797,N_5492,N_5369);
nor U5798 (N_5798,N_5256,N_5272);
xnor U5799 (N_5799,N_5384,N_5460);
and U5800 (N_5800,N_5185,N_5320);
and U5801 (N_5801,N_5291,N_5369);
xor U5802 (N_5802,N_5071,N_5371);
xnor U5803 (N_5803,N_5348,N_5067);
xor U5804 (N_5804,N_5257,N_5455);
or U5805 (N_5805,N_5128,N_5241);
xor U5806 (N_5806,N_5232,N_5378);
or U5807 (N_5807,N_5483,N_5097);
nor U5808 (N_5808,N_5355,N_5004);
nor U5809 (N_5809,N_5104,N_5396);
nor U5810 (N_5810,N_5097,N_5284);
xnor U5811 (N_5811,N_5108,N_5279);
nor U5812 (N_5812,N_5439,N_5085);
nor U5813 (N_5813,N_5209,N_5150);
or U5814 (N_5814,N_5433,N_5277);
xnor U5815 (N_5815,N_5401,N_5078);
or U5816 (N_5816,N_5145,N_5370);
or U5817 (N_5817,N_5448,N_5459);
and U5818 (N_5818,N_5138,N_5352);
and U5819 (N_5819,N_5174,N_5089);
xnor U5820 (N_5820,N_5447,N_5067);
xnor U5821 (N_5821,N_5085,N_5001);
nand U5822 (N_5822,N_5248,N_5048);
and U5823 (N_5823,N_5202,N_5181);
and U5824 (N_5824,N_5204,N_5372);
nor U5825 (N_5825,N_5197,N_5279);
or U5826 (N_5826,N_5072,N_5259);
xor U5827 (N_5827,N_5336,N_5084);
or U5828 (N_5828,N_5313,N_5101);
nor U5829 (N_5829,N_5014,N_5394);
and U5830 (N_5830,N_5216,N_5306);
xor U5831 (N_5831,N_5260,N_5416);
nor U5832 (N_5832,N_5127,N_5333);
or U5833 (N_5833,N_5253,N_5004);
and U5834 (N_5834,N_5245,N_5281);
nand U5835 (N_5835,N_5248,N_5123);
or U5836 (N_5836,N_5422,N_5482);
xor U5837 (N_5837,N_5093,N_5021);
or U5838 (N_5838,N_5275,N_5151);
nor U5839 (N_5839,N_5292,N_5044);
nor U5840 (N_5840,N_5053,N_5349);
xor U5841 (N_5841,N_5097,N_5273);
nor U5842 (N_5842,N_5288,N_5390);
xor U5843 (N_5843,N_5179,N_5349);
nand U5844 (N_5844,N_5101,N_5128);
nor U5845 (N_5845,N_5477,N_5448);
and U5846 (N_5846,N_5199,N_5040);
and U5847 (N_5847,N_5390,N_5057);
nand U5848 (N_5848,N_5414,N_5306);
nor U5849 (N_5849,N_5241,N_5061);
xor U5850 (N_5850,N_5475,N_5244);
nor U5851 (N_5851,N_5426,N_5187);
or U5852 (N_5852,N_5335,N_5217);
nand U5853 (N_5853,N_5034,N_5431);
xnor U5854 (N_5854,N_5476,N_5152);
nor U5855 (N_5855,N_5263,N_5044);
nand U5856 (N_5856,N_5192,N_5230);
xor U5857 (N_5857,N_5213,N_5137);
nor U5858 (N_5858,N_5491,N_5144);
or U5859 (N_5859,N_5467,N_5204);
nor U5860 (N_5860,N_5152,N_5005);
nand U5861 (N_5861,N_5201,N_5307);
nor U5862 (N_5862,N_5123,N_5351);
nand U5863 (N_5863,N_5209,N_5398);
and U5864 (N_5864,N_5152,N_5285);
or U5865 (N_5865,N_5181,N_5424);
xnor U5866 (N_5866,N_5235,N_5499);
or U5867 (N_5867,N_5472,N_5465);
or U5868 (N_5868,N_5302,N_5331);
nand U5869 (N_5869,N_5402,N_5217);
nor U5870 (N_5870,N_5112,N_5190);
and U5871 (N_5871,N_5324,N_5289);
and U5872 (N_5872,N_5319,N_5346);
nor U5873 (N_5873,N_5418,N_5488);
nand U5874 (N_5874,N_5384,N_5417);
nor U5875 (N_5875,N_5009,N_5459);
and U5876 (N_5876,N_5487,N_5435);
nor U5877 (N_5877,N_5205,N_5326);
and U5878 (N_5878,N_5106,N_5490);
and U5879 (N_5879,N_5316,N_5315);
nor U5880 (N_5880,N_5299,N_5306);
nor U5881 (N_5881,N_5445,N_5471);
xnor U5882 (N_5882,N_5114,N_5421);
nor U5883 (N_5883,N_5142,N_5434);
xor U5884 (N_5884,N_5345,N_5457);
nand U5885 (N_5885,N_5129,N_5114);
or U5886 (N_5886,N_5256,N_5157);
and U5887 (N_5887,N_5451,N_5104);
nand U5888 (N_5888,N_5230,N_5476);
nor U5889 (N_5889,N_5094,N_5059);
and U5890 (N_5890,N_5064,N_5494);
nor U5891 (N_5891,N_5241,N_5096);
or U5892 (N_5892,N_5021,N_5205);
xnor U5893 (N_5893,N_5254,N_5370);
xnor U5894 (N_5894,N_5191,N_5166);
and U5895 (N_5895,N_5352,N_5407);
nand U5896 (N_5896,N_5030,N_5322);
and U5897 (N_5897,N_5173,N_5296);
nand U5898 (N_5898,N_5170,N_5402);
nor U5899 (N_5899,N_5375,N_5179);
xor U5900 (N_5900,N_5256,N_5423);
and U5901 (N_5901,N_5093,N_5427);
xnor U5902 (N_5902,N_5404,N_5494);
nor U5903 (N_5903,N_5441,N_5032);
nand U5904 (N_5904,N_5147,N_5454);
xnor U5905 (N_5905,N_5400,N_5086);
xor U5906 (N_5906,N_5313,N_5163);
nor U5907 (N_5907,N_5272,N_5398);
nor U5908 (N_5908,N_5293,N_5010);
or U5909 (N_5909,N_5499,N_5273);
xnor U5910 (N_5910,N_5240,N_5109);
nand U5911 (N_5911,N_5139,N_5239);
nand U5912 (N_5912,N_5454,N_5195);
nor U5913 (N_5913,N_5032,N_5051);
xor U5914 (N_5914,N_5338,N_5201);
nand U5915 (N_5915,N_5240,N_5495);
nor U5916 (N_5916,N_5076,N_5060);
and U5917 (N_5917,N_5079,N_5124);
nor U5918 (N_5918,N_5124,N_5372);
xor U5919 (N_5919,N_5489,N_5231);
or U5920 (N_5920,N_5097,N_5383);
nor U5921 (N_5921,N_5428,N_5172);
nand U5922 (N_5922,N_5437,N_5261);
and U5923 (N_5923,N_5421,N_5443);
nand U5924 (N_5924,N_5486,N_5300);
nor U5925 (N_5925,N_5086,N_5084);
xor U5926 (N_5926,N_5436,N_5359);
and U5927 (N_5927,N_5017,N_5163);
and U5928 (N_5928,N_5463,N_5085);
and U5929 (N_5929,N_5244,N_5094);
xor U5930 (N_5930,N_5222,N_5085);
and U5931 (N_5931,N_5192,N_5472);
nand U5932 (N_5932,N_5257,N_5073);
or U5933 (N_5933,N_5291,N_5060);
xnor U5934 (N_5934,N_5477,N_5122);
and U5935 (N_5935,N_5365,N_5438);
or U5936 (N_5936,N_5270,N_5264);
xnor U5937 (N_5937,N_5425,N_5447);
nand U5938 (N_5938,N_5438,N_5237);
or U5939 (N_5939,N_5139,N_5326);
and U5940 (N_5940,N_5078,N_5284);
or U5941 (N_5941,N_5421,N_5169);
nand U5942 (N_5942,N_5166,N_5380);
nand U5943 (N_5943,N_5027,N_5455);
or U5944 (N_5944,N_5409,N_5437);
and U5945 (N_5945,N_5241,N_5485);
or U5946 (N_5946,N_5202,N_5313);
nand U5947 (N_5947,N_5189,N_5087);
nor U5948 (N_5948,N_5185,N_5109);
and U5949 (N_5949,N_5183,N_5068);
nor U5950 (N_5950,N_5308,N_5045);
and U5951 (N_5951,N_5063,N_5297);
or U5952 (N_5952,N_5323,N_5036);
and U5953 (N_5953,N_5220,N_5072);
nand U5954 (N_5954,N_5164,N_5369);
or U5955 (N_5955,N_5081,N_5050);
nor U5956 (N_5956,N_5001,N_5461);
nor U5957 (N_5957,N_5162,N_5361);
and U5958 (N_5958,N_5212,N_5409);
xnor U5959 (N_5959,N_5487,N_5032);
or U5960 (N_5960,N_5360,N_5119);
xor U5961 (N_5961,N_5089,N_5310);
xor U5962 (N_5962,N_5276,N_5069);
or U5963 (N_5963,N_5492,N_5371);
and U5964 (N_5964,N_5278,N_5099);
xnor U5965 (N_5965,N_5214,N_5033);
nand U5966 (N_5966,N_5356,N_5154);
xnor U5967 (N_5967,N_5374,N_5461);
nand U5968 (N_5968,N_5479,N_5304);
and U5969 (N_5969,N_5415,N_5149);
and U5970 (N_5970,N_5250,N_5445);
nand U5971 (N_5971,N_5168,N_5471);
xnor U5972 (N_5972,N_5466,N_5380);
nor U5973 (N_5973,N_5124,N_5047);
nand U5974 (N_5974,N_5480,N_5275);
and U5975 (N_5975,N_5051,N_5085);
and U5976 (N_5976,N_5206,N_5417);
and U5977 (N_5977,N_5150,N_5218);
nor U5978 (N_5978,N_5358,N_5333);
or U5979 (N_5979,N_5119,N_5330);
and U5980 (N_5980,N_5345,N_5486);
and U5981 (N_5981,N_5492,N_5218);
nand U5982 (N_5982,N_5328,N_5019);
nor U5983 (N_5983,N_5291,N_5110);
or U5984 (N_5984,N_5064,N_5354);
and U5985 (N_5985,N_5335,N_5094);
xnor U5986 (N_5986,N_5258,N_5059);
nor U5987 (N_5987,N_5304,N_5182);
xnor U5988 (N_5988,N_5467,N_5227);
nand U5989 (N_5989,N_5354,N_5166);
nand U5990 (N_5990,N_5082,N_5110);
and U5991 (N_5991,N_5014,N_5392);
nand U5992 (N_5992,N_5281,N_5435);
and U5993 (N_5993,N_5347,N_5415);
nor U5994 (N_5994,N_5319,N_5149);
and U5995 (N_5995,N_5215,N_5469);
nand U5996 (N_5996,N_5438,N_5376);
xnor U5997 (N_5997,N_5469,N_5132);
nor U5998 (N_5998,N_5036,N_5406);
nand U5999 (N_5999,N_5235,N_5433);
xnor U6000 (N_6000,N_5737,N_5640);
nand U6001 (N_6001,N_5528,N_5571);
nor U6002 (N_6002,N_5855,N_5920);
or U6003 (N_6003,N_5516,N_5746);
nor U6004 (N_6004,N_5934,N_5545);
xor U6005 (N_6005,N_5685,N_5797);
nand U6006 (N_6006,N_5661,N_5727);
or U6007 (N_6007,N_5662,N_5874);
nor U6008 (N_6008,N_5778,N_5579);
and U6009 (N_6009,N_5651,N_5834);
or U6010 (N_6010,N_5719,N_5506);
nand U6011 (N_6011,N_5782,N_5846);
nand U6012 (N_6012,N_5523,N_5677);
nand U6013 (N_6013,N_5619,N_5665);
nand U6014 (N_6014,N_5938,N_5533);
and U6015 (N_6015,N_5713,N_5577);
nor U6016 (N_6016,N_5763,N_5900);
xor U6017 (N_6017,N_5546,N_5784);
or U6018 (N_6018,N_5927,N_5954);
nor U6019 (N_6019,N_5936,N_5884);
and U6020 (N_6020,N_5872,N_5957);
xnor U6021 (N_6021,N_5978,N_5827);
nor U6022 (N_6022,N_5632,N_5606);
and U6023 (N_6023,N_5725,N_5531);
nor U6024 (N_6024,N_5948,N_5892);
nand U6025 (N_6025,N_5572,N_5880);
xor U6026 (N_6026,N_5617,N_5734);
nor U6027 (N_6027,N_5692,N_5802);
or U6028 (N_6028,N_5966,N_5578);
or U6029 (N_6029,N_5645,N_5564);
nand U6030 (N_6030,N_5736,N_5553);
nand U6031 (N_6031,N_5696,N_5870);
nand U6032 (N_6032,N_5952,N_5684);
and U6033 (N_6033,N_5994,N_5702);
xnor U6034 (N_6034,N_5964,N_5961);
xnor U6035 (N_6035,N_5507,N_5897);
nor U6036 (N_6036,N_5607,N_5730);
and U6037 (N_6037,N_5574,N_5982);
nand U6038 (N_6038,N_5840,N_5621);
and U6039 (N_6039,N_5896,N_5613);
and U6040 (N_6040,N_5803,N_5799);
or U6041 (N_6041,N_5521,N_5551);
xor U6042 (N_6042,N_5882,N_5538);
xnor U6043 (N_6043,N_5996,N_5805);
nand U6044 (N_6044,N_5536,N_5723);
and U6045 (N_6045,N_5541,N_5556);
and U6046 (N_6046,N_5804,N_5829);
or U6047 (N_6047,N_5659,N_5945);
nand U6048 (N_6048,N_5749,N_5599);
nor U6049 (N_6049,N_5597,N_5608);
xor U6050 (N_6050,N_5540,N_5776);
or U6051 (N_6051,N_5976,N_5745);
nor U6052 (N_6052,N_5625,N_5604);
and U6053 (N_6053,N_5601,N_5844);
or U6054 (N_6054,N_5832,N_5637);
nor U6055 (N_6055,N_5714,N_5841);
or U6056 (N_6056,N_5825,N_5594);
nand U6057 (N_6057,N_5974,N_5548);
xnor U6058 (N_6058,N_5807,N_5850);
nand U6059 (N_6059,N_5911,N_5694);
xnor U6060 (N_6060,N_5849,N_5647);
nor U6061 (N_6061,N_5678,N_5753);
nand U6062 (N_6062,N_5770,N_5583);
or U6063 (N_6063,N_5916,N_5837);
or U6064 (N_6064,N_5886,N_5748);
nand U6065 (N_6065,N_5854,N_5923);
nor U6066 (N_6066,N_5666,N_5906);
and U6067 (N_6067,N_5699,N_5649);
or U6068 (N_6068,N_5963,N_5510);
and U6069 (N_6069,N_5986,N_5774);
or U6070 (N_6070,N_5527,N_5971);
nand U6071 (N_6071,N_5672,N_5819);
nand U6072 (N_6072,N_5838,N_5915);
nand U6073 (N_6073,N_5650,N_5783);
nand U6074 (N_6074,N_5806,N_5925);
nor U6075 (N_6075,N_5522,N_5544);
and U6076 (N_6076,N_5997,N_5519);
and U6077 (N_6077,N_5969,N_5983);
nor U6078 (N_6078,N_5566,N_5673);
xor U6079 (N_6079,N_5740,N_5861);
nor U6080 (N_6080,N_5656,N_5798);
xnor U6081 (N_6081,N_5909,N_5683);
nand U6082 (N_6082,N_5929,N_5575);
or U6083 (N_6083,N_5639,N_5705);
nand U6084 (N_6084,N_5524,N_5990);
and U6085 (N_6085,N_5977,N_5959);
nand U6086 (N_6086,N_5750,N_5771);
xor U6087 (N_6087,N_5813,N_5901);
or U6088 (N_6088,N_5542,N_5612);
nand U6089 (N_6089,N_5823,N_5967);
or U6090 (N_6090,N_5590,N_5922);
or U6091 (N_6091,N_5693,N_5554);
nor U6092 (N_6092,N_5570,N_5998);
nand U6093 (N_6093,N_5831,N_5532);
or U6094 (N_6094,N_5576,N_5586);
xnor U6095 (N_6095,N_5615,N_5931);
nand U6096 (N_6096,N_5557,N_5535);
xor U6097 (N_6097,N_5739,N_5968);
xor U6098 (N_6098,N_5944,N_5883);
and U6099 (N_6099,N_5985,N_5518);
nand U6100 (N_6100,N_5869,N_5603);
nor U6101 (N_6101,N_5709,N_5843);
and U6102 (N_6102,N_5525,N_5933);
nor U6103 (N_6103,N_5867,N_5851);
nand U6104 (N_6104,N_5853,N_5898);
and U6105 (N_6105,N_5756,N_5708);
and U6106 (N_6106,N_5835,N_5779);
nand U6107 (N_6107,N_5686,N_5690);
or U6108 (N_6108,N_5777,N_5676);
xor U6109 (N_6109,N_5620,N_5790);
and U6110 (N_6110,N_5689,N_5633);
nor U6111 (N_6111,N_5947,N_5810);
nand U6112 (N_6112,N_5537,N_5657);
nor U6113 (N_6113,N_5800,N_5818);
xnor U6114 (N_6114,N_5664,N_5926);
and U6115 (N_6115,N_5724,N_5588);
and U6116 (N_6116,N_5644,N_5887);
xor U6117 (N_6117,N_5668,N_5716);
nor U6118 (N_6118,N_5755,N_5768);
nor U6119 (N_6119,N_5559,N_5914);
nand U6120 (N_6120,N_5932,N_5503);
or U6121 (N_6121,N_5866,N_5589);
xnor U6122 (N_6122,N_5711,N_5600);
and U6123 (N_6123,N_5616,N_5773);
and U6124 (N_6124,N_5529,N_5757);
nand U6125 (N_6125,N_5842,N_5654);
or U6126 (N_6126,N_5808,N_5965);
and U6127 (N_6127,N_5951,N_5735);
nor U6128 (N_6128,N_5940,N_5772);
nor U6129 (N_6129,N_5609,N_5707);
nand U6130 (N_6130,N_5681,N_5949);
or U6131 (N_6131,N_5717,N_5895);
nor U6132 (N_6132,N_5928,N_5581);
nor U6133 (N_6133,N_5863,N_5520);
xnor U6134 (N_6134,N_5549,N_5624);
and U6135 (N_6135,N_5824,N_5862);
or U6136 (N_6136,N_5917,N_5913);
nand U6137 (N_6137,N_5688,N_5958);
or U6138 (N_6138,N_5631,N_5674);
nor U6139 (N_6139,N_5787,N_5858);
nor U6140 (N_6140,N_5747,N_5742);
and U6141 (N_6141,N_5955,N_5698);
xor U6142 (N_6142,N_5643,N_5703);
xnor U6143 (N_6143,N_5560,N_5663);
nor U6144 (N_6144,N_5960,N_5878);
and U6145 (N_6145,N_5598,N_5762);
or U6146 (N_6146,N_5511,N_5973);
nor U6147 (N_6147,N_5513,N_5732);
xnor U6148 (N_6148,N_5836,N_5890);
or U6149 (N_6149,N_5902,N_5515);
nor U6150 (N_6150,N_5764,N_5567);
and U6151 (N_6151,N_5828,N_5852);
nor U6152 (N_6152,N_5543,N_5585);
xnor U6153 (N_6153,N_5814,N_5864);
or U6154 (N_6154,N_5697,N_5539);
nor U6155 (N_6155,N_5670,N_5738);
nand U6156 (N_6156,N_5918,N_5587);
nand U6157 (N_6157,N_5565,N_5817);
nor U6158 (N_6158,N_5675,N_5962);
nor U6159 (N_6159,N_5526,N_5839);
and U6160 (N_6160,N_5642,N_5593);
and U6161 (N_6161,N_5903,N_5975);
nand U6162 (N_6162,N_5752,N_5530);
or U6163 (N_6163,N_5634,N_5879);
or U6164 (N_6164,N_5584,N_5569);
xnor U6165 (N_6165,N_5627,N_5641);
xor U6166 (N_6166,N_5899,N_5726);
nand U6167 (N_6167,N_5626,N_5534);
nand U6168 (N_6168,N_5793,N_5759);
or U6169 (N_6169,N_5781,N_5956);
nand U6170 (N_6170,N_5706,N_5871);
xor U6171 (N_6171,N_5780,N_5943);
and U6172 (N_6172,N_5789,N_5667);
and U6173 (N_6173,N_5991,N_5580);
or U6174 (N_6174,N_5988,N_5939);
or U6175 (N_6175,N_5905,N_5636);
xor U6176 (N_6176,N_5505,N_5652);
and U6177 (N_6177,N_5733,N_5595);
or U6178 (N_6178,N_5791,N_5721);
and U6179 (N_6179,N_5761,N_5989);
and U6180 (N_6180,N_5875,N_5618);
nand U6181 (N_6181,N_5517,N_5891);
nand U6182 (N_6182,N_5816,N_5833);
nand U6183 (N_6183,N_5728,N_5942);
and U6184 (N_6184,N_5704,N_5876);
or U6185 (N_6185,N_5582,N_5889);
nand U6186 (N_6186,N_5552,N_5741);
xor U6187 (N_6187,N_5970,N_5504);
nand U6188 (N_6188,N_5687,N_5812);
nand U6189 (N_6189,N_5826,N_5710);
or U6190 (N_6190,N_5563,N_5547);
and U6191 (N_6191,N_5775,N_5946);
and U6192 (N_6192,N_5981,N_5561);
or U6193 (N_6193,N_5910,N_5655);
or U6194 (N_6194,N_5795,N_5820);
xor U6195 (N_6195,N_5701,N_5907);
nand U6196 (N_6196,N_5682,N_5822);
or U6197 (N_6197,N_5646,N_5873);
nor U6198 (N_6198,N_5999,N_5658);
or U6199 (N_6199,N_5785,N_5865);
nor U6200 (N_6200,N_5950,N_5514);
nand U6201 (N_6201,N_5502,N_5729);
xnor U6202 (N_6202,N_5629,N_5767);
nor U6203 (N_6203,N_5691,N_5671);
xnor U6204 (N_6204,N_5630,N_5592);
nor U6205 (N_6205,N_5648,N_5792);
or U6206 (N_6206,N_5635,N_5765);
or U6207 (N_6207,N_5602,N_5758);
nand U6208 (N_6208,N_5788,N_5937);
or U6209 (N_6209,N_5857,N_5794);
nor U6210 (N_6210,N_5848,N_5766);
and U6211 (N_6211,N_5550,N_5801);
xnor U6212 (N_6212,N_5953,N_5611);
or U6213 (N_6213,N_5786,N_5980);
nor U6214 (N_6214,N_5845,N_5509);
xor U6215 (N_6215,N_5501,N_5679);
and U6216 (N_6216,N_5568,N_5894);
or U6217 (N_6217,N_5815,N_5984);
or U6218 (N_6218,N_5860,N_5500);
xnor U6219 (N_6219,N_5993,N_5904);
xnor U6220 (N_6220,N_5888,N_5660);
nand U6221 (N_6221,N_5508,N_5605);
or U6222 (N_6222,N_5893,N_5614);
xor U6223 (N_6223,N_5669,N_5722);
nand U6224 (N_6224,N_5856,N_5638);
xor U6225 (N_6225,N_5847,N_5811);
nand U6226 (N_6226,N_5596,N_5715);
xnor U6227 (N_6227,N_5720,N_5751);
nor U6228 (N_6228,N_5718,N_5743);
and U6229 (N_6229,N_5995,N_5695);
or U6230 (N_6230,N_5912,N_5591);
nand U6231 (N_6231,N_5744,N_5859);
or U6232 (N_6232,N_5908,N_5628);
xor U6233 (N_6233,N_5809,N_5979);
and U6234 (N_6234,N_5760,N_5653);
nand U6235 (N_6235,N_5558,N_5921);
or U6236 (N_6236,N_5712,N_5992);
nand U6237 (N_6237,N_5935,N_5868);
nand U6238 (N_6238,N_5877,N_5796);
nor U6239 (N_6239,N_5830,N_5680);
or U6240 (N_6240,N_5573,N_5512);
and U6241 (N_6241,N_5622,N_5623);
xor U6242 (N_6242,N_5881,N_5972);
or U6243 (N_6243,N_5941,N_5731);
nor U6244 (N_6244,N_5555,N_5700);
nor U6245 (N_6245,N_5610,N_5919);
or U6246 (N_6246,N_5924,N_5754);
or U6247 (N_6247,N_5930,N_5769);
xor U6248 (N_6248,N_5987,N_5562);
xor U6249 (N_6249,N_5821,N_5885);
or U6250 (N_6250,N_5674,N_5754);
nand U6251 (N_6251,N_5653,N_5713);
and U6252 (N_6252,N_5603,N_5952);
or U6253 (N_6253,N_5621,N_5594);
nand U6254 (N_6254,N_5837,N_5759);
xor U6255 (N_6255,N_5985,N_5824);
nor U6256 (N_6256,N_5773,N_5528);
or U6257 (N_6257,N_5638,N_5912);
xor U6258 (N_6258,N_5896,N_5827);
or U6259 (N_6259,N_5884,N_5800);
or U6260 (N_6260,N_5571,N_5855);
nand U6261 (N_6261,N_5624,N_5524);
or U6262 (N_6262,N_5719,N_5818);
and U6263 (N_6263,N_5608,N_5783);
or U6264 (N_6264,N_5765,N_5676);
or U6265 (N_6265,N_5854,N_5628);
nor U6266 (N_6266,N_5528,N_5976);
or U6267 (N_6267,N_5914,N_5785);
nand U6268 (N_6268,N_5973,N_5521);
nand U6269 (N_6269,N_5676,N_5709);
xnor U6270 (N_6270,N_5908,N_5916);
xor U6271 (N_6271,N_5951,N_5500);
xnor U6272 (N_6272,N_5689,N_5573);
and U6273 (N_6273,N_5881,N_5736);
nor U6274 (N_6274,N_5834,N_5817);
xor U6275 (N_6275,N_5831,N_5633);
and U6276 (N_6276,N_5788,N_5841);
or U6277 (N_6277,N_5892,N_5945);
nand U6278 (N_6278,N_5763,N_5643);
and U6279 (N_6279,N_5616,N_5834);
or U6280 (N_6280,N_5732,N_5706);
nor U6281 (N_6281,N_5975,N_5653);
xnor U6282 (N_6282,N_5597,N_5995);
xor U6283 (N_6283,N_5568,N_5663);
or U6284 (N_6284,N_5506,N_5671);
nand U6285 (N_6285,N_5737,N_5945);
xnor U6286 (N_6286,N_5904,N_5585);
xnor U6287 (N_6287,N_5528,N_5513);
or U6288 (N_6288,N_5811,N_5628);
and U6289 (N_6289,N_5733,N_5830);
and U6290 (N_6290,N_5888,N_5985);
or U6291 (N_6291,N_5716,N_5973);
or U6292 (N_6292,N_5738,N_5906);
xor U6293 (N_6293,N_5877,N_5542);
nand U6294 (N_6294,N_5991,N_5951);
nor U6295 (N_6295,N_5729,N_5763);
and U6296 (N_6296,N_5588,N_5729);
and U6297 (N_6297,N_5614,N_5892);
xor U6298 (N_6298,N_5538,N_5766);
and U6299 (N_6299,N_5681,N_5684);
nor U6300 (N_6300,N_5772,N_5801);
nand U6301 (N_6301,N_5836,N_5891);
xnor U6302 (N_6302,N_5803,N_5671);
xnor U6303 (N_6303,N_5637,N_5682);
or U6304 (N_6304,N_5989,N_5921);
and U6305 (N_6305,N_5608,N_5940);
or U6306 (N_6306,N_5692,N_5576);
and U6307 (N_6307,N_5962,N_5999);
xor U6308 (N_6308,N_5647,N_5881);
or U6309 (N_6309,N_5808,N_5825);
nand U6310 (N_6310,N_5954,N_5743);
or U6311 (N_6311,N_5640,N_5827);
xor U6312 (N_6312,N_5832,N_5646);
and U6313 (N_6313,N_5610,N_5804);
and U6314 (N_6314,N_5500,N_5515);
nand U6315 (N_6315,N_5898,N_5887);
or U6316 (N_6316,N_5847,N_5643);
nor U6317 (N_6317,N_5546,N_5683);
or U6318 (N_6318,N_5712,N_5943);
nor U6319 (N_6319,N_5672,N_5871);
and U6320 (N_6320,N_5786,N_5948);
nand U6321 (N_6321,N_5745,N_5921);
nor U6322 (N_6322,N_5513,N_5634);
nor U6323 (N_6323,N_5749,N_5854);
nand U6324 (N_6324,N_5641,N_5745);
and U6325 (N_6325,N_5938,N_5651);
nand U6326 (N_6326,N_5865,N_5706);
or U6327 (N_6327,N_5933,N_5957);
and U6328 (N_6328,N_5653,N_5614);
or U6329 (N_6329,N_5939,N_5736);
and U6330 (N_6330,N_5568,N_5702);
nand U6331 (N_6331,N_5753,N_5623);
nor U6332 (N_6332,N_5876,N_5868);
nand U6333 (N_6333,N_5632,N_5993);
xnor U6334 (N_6334,N_5800,N_5663);
and U6335 (N_6335,N_5949,N_5736);
xor U6336 (N_6336,N_5559,N_5727);
xor U6337 (N_6337,N_5768,N_5756);
nand U6338 (N_6338,N_5973,N_5532);
and U6339 (N_6339,N_5578,N_5577);
nand U6340 (N_6340,N_5907,N_5717);
xnor U6341 (N_6341,N_5911,N_5936);
nand U6342 (N_6342,N_5707,N_5829);
nor U6343 (N_6343,N_5964,N_5547);
nand U6344 (N_6344,N_5701,N_5860);
or U6345 (N_6345,N_5521,N_5947);
and U6346 (N_6346,N_5526,N_5851);
and U6347 (N_6347,N_5768,N_5598);
nor U6348 (N_6348,N_5713,N_5884);
nor U6349 (N_6349,N_5972,N_5550);
and U6350 (N_6350,N_5564,N_5607);
xnor U6351 (N_6351,N_5905,N_5913);
or U6352 (N_6352,N_5797,N_5849);
and U6353 (N_6353,N_5516,N_5648);
nor U6354 (N_6354,N_5877,N_5747);
nor U6355 (N_6355,N_5995,N_5742);
nor U6356 (N_6356,N_5710,N_5937);
or U6357 (N_6357,N_5719,N_5702);
nor U6358 (N_6358,N_5533,N_5865);
and U6359 (N_6359,N_5529,N_5992);
and U6360 (N_6360,N_5759,N_5689);
nand U6361 (N_6361,N_5885,N_5718);
nor U6362 (N_6362,N_5565,N_5959);
and U6363 (N_6363,N_5880,N_5700);
or U6364 (N_6364,N_5977,N_5552);
and U6365 (N_6365,N_5946,N_5898);
nand U6366 (N_6366,N_5883,N_5659);
nand U6367 (N_6367,N_5730,N_5915);
or U6368 (N_6368,N_5537,N_5746);
or U6369 (N_6369,N_5962,N_5529);
nand U6370 (N_6370,N_5600,N_5578);
nor U6371 (N_6371,N_5757,N_5921);
xnor U6372 (N_6372,N_5684,N_5602);
or U6373 (N_6373,N_5927,N_5804);
nor U6374 (N_6374,N_5750,N_5766);
nor U6375 (N_6375,N_5780,N_5997);
nand U6376 (N_6376,N_5794,N_5697);
or U6377 (N_6377,N_5778,N_5646);
nand U6378 (N_6378,N_5979,N_5812);
and U6379 (N_6379,N_5624,N_5925);
xnor U6380 (N_6380,N_5520,N_5952);
nor U6381 (N_6381,N_5549,N_5871);
or U6382 (N_6382,N_5900,N_5759);
nand U6383 (N_6383,N_5560,N_5687);
or U6384 (N_6384,N_5988,N_5670);
or U6385 (N_6385,N_5667,N_5543);
and U6386 (N_6386,N_5715,N_5878);
xnor U6387 (N_6387,N_5713,N_5790);
or U6388 (N_6388,N_5510,N_5707);
or U6389 (N_6389,N_5815,N_5587);
nand U6390 (N_6390,N_5608,N_5721);
or U6391 (N_6391,N_5976,N_5599);
and U6392 (N_6392,N_5668,N_5984);
nor U6393 (N_6393,N_5832,N_5530);
xnor U6394 (N_6394,N_5749,N_5670);
nor U6395 (N_6395,N_5880,N_5655);
and U6396 (N_6396,N_5610,N_5531);
or U6397 (N_6397,N_5514,N_5941);
xor U6398 (N_6398,N_5855,N_5629);
nand U6399 (N_6399,N_5625,N_5526);
nand U6400 (N_6400,N_5692,N_5598);
xnor U6401 (N_6401,N_5978,N_5860);
and U6402 (N_6402,N_5688,N_5979);
and U6403 (N_6403,N_5932,N_5510);
and U6404 (N_6404,N_5712,N_5556);
nor U6405 (N_6405,N_5669,N_5829);
xnor U6406 (N_6406,N_5544,N_5916);
and U6407 (N_6407,N_5956,N_5535);
and U6408 (N_6408,N_5811,N_5917);
or U6409 (N_6409,N_5652,N_5720);
and U6410 (N_6410,N_5916,N_5993);
or U6411 (N_6411,N_5816,N_5960);
nand U6412 (N_6412,N_5933,N_5713);
xor U6413 (N_6413,N_5606,N_5654);
nor U6414 (N_6414,N_5608,N_5808);
and U6415 (N_6415,N_5881,N_5729);
nor U6416 (N_6416,N_5800,N_5886);
nor U6417 (N_6417,N_5776,N_5911);
or U6418 (N_6418,N_5589,N_5801);
and U6419 (N_6419,N_5875,N_5566);
nor U6420 (N_6420,N_5893,N_5692);
nand U6421 (N_6421,N_5622,N_5841);
xnor U6422 (N_6422,N_5968,N_5660);
and U6423 (N_6423,N_5838,N_5926);
and U6424 (N_6424,N_5942,N_5965);
nor U6425 (N_6425,N_5566,N_5956);
nor U6426 (N_6426,N_5637,N_5915);
nor U6427 (N_6427,N_5552,N_5731);
and U6428 (N_6428,N_5625,N_5885);
or U6429 (N_6429,N_5801,N_5982);
xnor U6430 (N_6430,N_5952,N_5640);
nor U6431 (N_6431,N_5723,N_5626);
or U6432 (N_6432,N_5705,N_5856);
xnor U6433 (N_6433,N_5576,N_5605);
nand U6434 (N_6434,N_5868,N_5519);
and U6435 (N_6435,N_5869,N_5952);
nor U6436 (N_6436,N_5677,N_5563);
nor U6437 (N_6437,N_5820,N_5528);
or U6438 (N_6438,N_5604,N_5871);
xor U6439 (N_6439,N_5845,N_5506);
nand U6440 (N_6440,N_5677,N_5559);
nor U6441 (N_6441,N_5504,N_5840);
nor U6442 (N_6442,N_5643,N_5765);
xnor U6443 (N_6443,N_5648,N_5786);
and U6444 (N_6444,N_5503,N_5778);
nand U6445 (N_6445,N_5673,N_5770);
and U6446 (N_6446,N_5588,N_5559);
xnor U6447 (N_6447,N_5772,N_5763);
or U6448 (N_6448,N_5886,N_5993);
nand U6449 (N_6449,N_5686,N_5542);
and U6450 (N_6450,N_5619,N_5577);
and U6451 (N_6451,N_5583,N_5756);
nand U6452 (N_6452,N_5975,N_5671);
nand U6453 (N_6453,N_5994,N_5922);
or U6454 (N_6454,N_5584,N_5627);
xor U6455 (N_6455,N_5844,N_5655);
nand U6456 (N_6456,N_5863,N_5963);
and U6457 (N_6457,N_5931,N_5691);
nor U6458 (N_6458,N_5729,N_5718);
xnor U6459 (N_6459,N_5893,N_5947);
or U6460 (N_6460,N_5725,N_5813);
and U6461 (N_6461,N_5781,N_5627);
and U6462 (N_6462,N_5912,N_5863);
or U6463 (N_6463,N_5815,N_5961);
nor U6464 (N_6464,N_5647,N_5517);
and U6465 (N_6465,N_5690,N_5664);
and U6466 (N_6466,N_5718,N_5600);
nor U6467 (N_6467,N_5864,N_5879);
or U6468 (N_6468,N_5931,N_5679);
xnor U6469 (N_6469,N_5591,N_5639);
xnor U6470 (N_6470,N_5953,N_5903);
or U6471 (N_6471,N_5860,N_5790);
and U6472 (N_6472,N_5739,N_5963);
nor U6473 (N_6473,N_5809,N_5646);
and U6474 (N_6474,N_5589,N_5973);
or U6475 (N_6475,N_5707,N_5775);
nor U6476 (N_6476,N_5646,N_5754);
nor U6477 (N_6477,N_5836,N_5646);
or U6478 (N_6478,N_5960,N_5956);
nand U6479 (N_6479,N_5557,N_5692);
and U6480 (N_6480,N_5957,N_5689);
nand U6481 (N_6481,N_5800,N_5759);
or U6482 (N_6482,N_5673,N_5680);
nor U6483 (N_6483,N_5771,N_5557);
or U6484 (N_6484,N_5676,N_5657);
nor U6485 (N_6485,N_5675,N_5623);
or U6486 (N_6486,N_5518,N_5637);
nand U6487 (N_6487,N_5901,N_5938);
nand U6488 (N_6488,N_5715,N_5636);
and U6489 (N_6489,N_5754,N_5619);
xnor U6490 (N_6490,N_5534,N_5655);
xnor U6491 (N_6491,N_5615,N_5843);
nand U6492 (N_6492,N_5687,N_5562);
and U6493 (N_6493,N_5594,N_5751);
nor U6494 (N_6494,N_5576,N_5941);
and U6495 (N_6495,N_5666,N_5687);
nor U6496 (N_6496,N_5736,N_5929);
nand U6497 (N_6497,N_5766,N_5881);
or U6498 (N_6498,N_5934,N_5758);
nor U6499 (N_6499,N_5500,N_5861);
xor U6500 (N_6500,N_6164,N_6078);
xnor U6501 (N_6501,N_6006,N_6094);
or U6502 (N_6502,N_6466,N_6000);
nand U6503 (N_6503,N_6417,N_6082);
or U6504 (N_6504,N_6367,N_6349);
xor U6505 (N_6505,N_6056,N_6184);
nand U6506 (N_6506,N_6409,N_6015);
nor U6507 (N_6507,N_6479,N_6033);
or U6508 (N_6508,N_6263,N_6259);
nor U6509 (N_6509,N_6273,N_6356);
and U6510 (N_6510,N_6211,N_6122);
or U6511 (N_6511,N_6221,N_6197);
nor U6512 (N_6512,N_6494,N_6061);
and U6513 (N_6513,N_6213,N_6181);
or U6514 (N_6514,N_6168,N_6342);
or U6515 (N_6515,N_6465,N_6423);
nor U6516 (N_6516,N_6125,N_6130);
xnor U6517 (N_6517,N_6176,N_6257);
and U6518 (N_6518,N_6270,N_6171);
nand U6519 (N_6519,N_6162,N_6388);
xnor U6520 (N_6520,N_6419,N_6426);
and U6521 (N_6521,N_6458,N_6253);
or U6522 (N_6522,N_6261,N_6452);
xnor U6523 (N_6523,N_6454,N_6413);
and U6524 (N_6524,N_6063,N_6072);
or U6525 (N_6525,N_6234,N_6028);
nand U6526 (N_6526,N_6475,N_6214);
nor U6527 (N_6527,N_6037,N_6498);
nand U6528 (N_6528,N_6442,N_6060);
or U6529 (N_6529,N_6222,N_6397);
xnor U6530 (N_6530,N_6414,N_6274);
nand U6531 (N_6531,N_6084,N_6205);
or U6532 (N_6532,N_6382,N_6100);
nand U6533 (N_6533,N_6371,N_6308);
xor U6534 (N_6534,N_6411,N_6251);
or U6535 (N_6535,N_6146,N_6359);
or U6536 (N_6536,N_6416,N_6286);
and U6537 (N_6537,N_6380,N_6188);
or U6538 (N_6538,N_6361,N_6480);
nand U6539 (N_6539,N_6165,N_6314);
xor U6540 (N_6540,N_6040,N_6212);
xor U6541 (N_6541,N_6249,N_6027);
or U6542 (N_6542,N_6155,N_6310);
nor U6543 (N_6543,N_6365,N_6473);
nor U6544 (N_6544,N_6300,N_6394);
nand U6545 (N_6545,N_6119,N_6085);
and U6546 (N_6546,N_6076,N_6333);
nand U6547 (N_6547,N_6192,N_6347);
nor U6548 (N_6548,N_6112,N_6116);
xor U6549 (N_6549,N_6421,N_6256);
nor U6550 (N_6550,N_6150,N_6358);
nand U6551 (N_6551,N_6364,N_6145);
or U6552 (N_6552,N_6489,N_6204);
nor U6553 (N_6553,N_6373,N_6231);
or U6554 (N_6554,N_6460,N_6478);
and U6555 (N_6555,N_6362,N_6280);
and U6556 (N_6556,N_6190,N_6011);
or U6557 (N_6557,N_6046,N_6449);
nor U6558 (N_6558,N_6317,N_6220);
or U6559 (N_6559,N_6346,N_6096);
nand U6560 (N_6560,N_6104,N_6341);
xor U6561 (N_6561,N_6081,N_6147);
nand U6562 (N_6562,N_6402,N_6293);
xnor U6563 (N_6563,N_6157,N_6114);
xnor U6564 (N_6564,N_6276,N_6319);
nand U6565 (N_6565,N_6003,N_6495);
nor U6566 (N_6566,N_6309,N_6343);
xnor U6567 (N_6567,N_6004,N_6327);
or U6568 (N_6568,N_6187,N_6185);
nand U6569 (N_6569,N_6170,N_6024);
nor U6570 (N_6570,N_6332,N_6196);
xor U6571 (N_6571,N_6316,N_6127);
nand U6572 (N_6572,N_6227,N_6313);
nor U6573 (N_6573,N_6101,N_6330);
nand U6574 (N_6574,N_6048,N_6376);
nor U6575 (N_6575,N_6285,N_6065);
or U6576 (N_6576,N_6203,N_6095);
and U6577 (N_6577,N_6363,N_6216);
xor U6578 (N_6578,N_6070,N_6225);
xor U6579 (N_6579,N_6183,N_6210);
or U6580 (N_6580,N_6055,N_6338);
xnor U6581 (N_6581,N_6329,N_6236);
nand U6582 (N_6582,N_6025,N_6389);
nand U6583 (N_6583,N_6215,N_6246);
or U6584 (N_6584,N_6008,N_6488);
nand U6585 (N_6585,N_6339,N_6174);
xnor U6586 (N_6586,N_6415,N_6194);
or U6587 (N_6587,N_6075,N_6272);
and U6588 (N_6588,N_6237,N_6120);
xnor U6589 (N_6589,N_6115,N_6090);
nor U6590 (N_6590,N_6296,N_6436);
and U6591 (N_6591,N_6400,N_6303);
or U6592 (N_6592,N_6250,N_6492);
nor U6593 (N_6593,N_6306,N_6066);
nor U6594 (N_6594,N_6158,N_6392);
xnor U6595 (N_6595,N_6219,N_6391);
xnor U6596 (N_6596,N_6351,N_6337);
nand U6597 (N_6597,N_6305,N_6186);
or U6598 (N_6598,N_6057,N_6434);
nor U6599 (N_6599,N_6019,N_6079);
xnor U6600 (N_6600,N_6062,N_6163);
nand U6601 (N_6601,N_6177,N_6258);
nor U6602 (N_6602,N_6029,N_6229);
xnor U6603 (N_6603,N_6036,N_6136);
nand U6604 (N_6604,N_6232,N_6375);
nor U6605 (N_6605,N_6265,N_6427);
nor U6606 (N_6606,N_6068,N_6050);
nand U6607 (N_6607,N_6422,N_6357);
or U6608 (N_6608,N_6175,N_6111);
nand U6609 (N_6609,N_6279,N_6401);
or U6610 (N_6610,N_6113,N_6148);
nor U6611 (N_6611,N_6200,N_6487);
nand U6612 (N_6612,N_6195,N_6178);
and U6613 (N_6613,N_6044,N_6097);
nor U6614 (N_6614,N_6016,N_6462);
xor U6615 (N_6615,N_6073,N_6277);
xnor U6616 (N_6616,N_6233,N_6052);
and U6617 (N_6617,N_6430,N_6266);
and U6618 (N_6618,N_6135,N_6297);
xor U6619 (N_6619,N_6433,N_6443);
and U6620 (N_6620,N_6385,N_6355);
nand U6621 (N_6621,N_6173,N_6269);
nor U6622 (N_6622,N_6344,N_6252);
or U6623 (N_6623,N_6091,N_6153);
nor U6624 (N_6624,N_6399,N_6491);
or U6625 (N_6625,N_6340,N_6047);
and U6626 (N_6626,N_6322,N_6275);
or U6627 (N_6627,N_6404,N_6141);
and U6628 (N_6628,N_6242,N_6374);
xor U6629 (N_6629,N_6467,N_6009);
and U6630 (N_6630,N_6331,N_6372);
or U6631 (N_6631,N_6217,N_6154);
nand U6632 (N_6632,N_6228,N_6323);
xnor U6633 (N_6633,N_6335,N_6034);
and U6634 (N_6634,N_6395,N_6282);
xnor U6635 (N_6635,N_6247,N_6124);
nor U6636 (N_6636,N_6243,N_6106);
nor U6637 (N_6637,N_6051,N_6360);
and U6638 (N_6638,N_6386,N_6069);
nand U6639 (N_6639,N_6118,N_6291);
xnor U6640 (N_6640,N_6302,N_6167);
xnor U6641 (N_6641,N_6117,N_6131);
or U6642 (N_6642,N_6030,N_6484);
or U6643 (N_6643,N_6447,N_6172);
and U6644 (N_6644,N_6469,N_6288);
or U6645 (N_6645,N_6295,N_6020);
xnor U6646 (N_6646,N_6089,N_6224);
nand U6647 (N_6647,N_6226,N_6180);
nand U6648 (N_6648,N_6022,N_6405);
xnor U6649 (N_6649,N_6451,N_6348);
nand U6650 (N_6650,N_6189,N_6059);
nor U6651 (N_6651,N_6099,N_6312);
nor U6652 (N_6652,N_6023,N_6448);
nor U6653 (N_6653,N_6207,N_6005);
nand U6654 (N_6654,N_6352,N_6370);
nand U6655 (N_6655,N_6139,N_6407);
nand U6656 (N_6656,N_6420,N_6456);
xor U6657 (N_6657,N_6126,N_6369);
nand U6658 (N_6658,N_6102,N_6377);
xor U6659 (N_6659,N_6138,N_6396);
and U6660 (N_6660,N_6461,N_6301);
nor U6661 (N_6661,N_6235,N_6384);
nand U6662 (N_6662,N_6408,N_6074);
nand U6663 (N_6663,N_6425,N_6080);
xor U6664 (N_6664,N_6156,N_6424);
xnor U6665 (N_6665,N_6109,N_6497);
nor U6666 (N_6666,N_6381,N_6268);
and U6667 (N_6667,N_6486,N_6318);
nor U6668 (N_6668,N_6262,N_6445);
and U6669 (N_6669,N_6209,N_6092);
xnor U6670 (N_6670,N_6083,N_6134);
xnor U6671 (N_6671,N_6483,N_6298);
xor U6672 (N_6672,N_6107,N_6328);
or U6673 (N_6673,N_6311,N_6455);
nand U6674 (N_6674,N_6453,N_6431);
nand U6675 (N_6675,N_6087,N_6432);
nand U6676 (N_6676,N_6325,N_6206);
xor U6677 (N_6677,N_6468,N_6035);
or U6678 (N_6678,N_6041,N_6179);
and U6679 (N_6679,N_6260,N_6238);
or U6680 (N_6680,N_6437,N_6086);
nor U6681 (N_6681,N_6129,N_6284);
nand U6682 (N_6682,N_6151,N_6105);
nor U6683 (N_6683,N_6198,N_6496);
nand U6684 (N_6684,N_6410,N_6470);
xnor U6685 (N_6685,N_6320,N_6240);
nand U6686 (N_6686,N_6199,N_6045);
and U6687 (N_6687,N_6223,N_6441);
and U6688 (N_6688,N_6039,N_6121);
nand U6689 (N_6689,N_6239,N_6058);
xnor U6690 (N_6690,N_6393,N_6354);
xor U6691 (N_6691,N_6038,N_6053);
and U6692 (N_6692,N_6334,N_6439);
nand U6693 (N_6693,N_6166,N_6387);
nor U6694 (N_6694,N_6191,N_6324);
and U6695 (N_6695,N_6123,N_6294);
xor U6696 (N_6696,N_6103,N_6007);
nand U6697 (N_6697,N_6481,N_6290);
and U6698 (N_6698,N_6013,N_6292);
and U6699 (N_6699,N_6304,N_6281);
and U6700 (N_6700,N_6042,N_6368);
nor U6701 (N_6701,N_6093,N_6098);
nand U6702 (N_6702,N_6110,N_6152);
xor U6703 (N_6703,N_6383,N_6321);
nand U6704 (N_6704,N_6471,N_6485);
nor U6705 (N_6705,N_6472,N_6245);
xor U6706 (N_6706,N_6350,N_6278);
or U6707 (N_6707,N_6026,N_6476);
and U6708 (N_6708,N_6149,N_6255);
and U6709 (N_6709,N_6429,N_6271);
nor U6710 (N_6710,N_6017,N_6398);
nand U6711 (N_6711,N_6128,N_6390);
nor U6712 (N_6712,N_6144,N_6012);
nand U6713 (N_6713,N_6244,N_6071);
or U6714 (N_6714,N_6435,N_6446);
xnor U6715 (N_6715,N_6326,N_6459);
and U6716 (N_6716,N_6193,N_6001);
xor U6717 (N_6717,N_6160,N_6307);
xor U6718 (N_6718,N_6406,N_6132);
and U6719 (N_6719,N_6287,N_6182);
nor U6720 (N_6720,N_6440,N_6201);
xor U6721 (N_6721,N_6267,N_6378);
nand U6722 (N_6722,N_6088,N_6379);
nor U6723 (N_6723,N_6064,N_6450);
nand U6724 (N_6724,N_6018,N_6049);
and U6725 (N_6725,N_6457,N_6463);
nand U6726 (N_6726,N_6067,N_6254);
nand U6727 (N_6727,N_6464,N_6031);
nor U6728 (N_6728,N_6299,N_6161);
nand U6729 (N_6729,N_6428,N_6202);
xnor U6730 (N_6730,N_6032,N_6002);
xor U6731 (N_6731,N_6137,N_6169);
or U6732 (N_6732,N_6021,N_6366);
nand U6733 (N_6733,N_6248,N_6283);
or U6734 (N_6734,N_6108,N_6499);
and U6735 (N_6735,N_6403,N_6159);
or U6736 (N_6736,N_6077,N_6444);
xor U6737 (N_6737,N_6482,N_6353);
and U6738 (N_6738,N_6140,N_6289);
or U6739 (N_6739,N_6241,N_6208);
and U6740 (N_6740,N_6315,N_6230);
or U6741 (N_6741,N_6477,N_6490);
xnor U6742 (N_6742,N_6218,N_6438);
xor U6743 (N_6743,N_6493,N_6142);
xnor U6744 (N_6744,N_6014,N_6010);
nand U6745 (N_6745,N_6143,N_6412);
nand U6746 (N_6746,N_6474,N_6336);
or U6747 (N_6747,N_6264,N_6418);
nand U6748 (N_6748,N_6133,N_6054);
or U6749 (N_6749,N_6043,N_6345);
nor U6750 (N_6750,N_6315,N_6166);
nor U6751 (N_6751,N_6254,N_6288);
nor U6752 (N_6752,N_6371,N_6404);
and U6753 (N_6753,N_6036,N_6302);
xor U6754 (N_6754,N_6207,N_6331);
xor U6755 (N_6755,N_6479,N_6371);
nor U6756 (N_6756,N_6168,N_6426);
nand U6757 (N_6757,N_6118,N_6180);
nand U6758 (N_6758,N_6065,N_6308);
nor U6759 (N_6759,N_6314,N_6370);
and U6760 (N_6760,N_6393,N_6300);
nor U6761 (N_6761,N_6303,N_6321);
nand U6762 (N_6762,N_6282,N_6343);
nor U6763 (N_6763,N_6305,N_6054);
nand U6764 (N_6764,N_6025,N_6426);
xor U6765 (N_6765,N_6071,N_6252);
nand U6766 (N_6766,N_6041,N_6461);
xor U6767 (N_6767,N_6046,N_6258);
and U6768 (N_6768,N_6389,N_6431);
xor U6769 (N_6769,N_6035,N_6414);
nor U6770 (N_6770,N_6197,N_6029);
nand U6771 (N_6771,N_6253,N_6272);
xnor U6772 (N_6772,N_6008,N_6280);
or U6773 (N_6773,N_6026,N_6376);
and U6774 (N_6774,N_6133,N_6038);
nand U6775 (N_6775,N_6203,N_6052);
and U6776 (N_6776,N_6212,N_6376);
xor U6777 (N_6777,N_6144,N_6056);
or U6778 (N_6778,N_6327,N_6367);
nor U6779 (N_6779,N_6447,N_6009);
nor U6780 (N_6780,N_6347,N_6313);
nor U6781 (N_6781,N_6169,N_6092);
nor U6782 (N_6782,N_6410,N_6383);
or U6783 (N_6783,N_6271,N_6479);
xor U6784 (N_6784,N_6359,N_6443);
nand U6785 (N_6785,N_6448,N_6018);
nor U6786 (N_6786,N_6376,N_6448);
and U6787 (N_6787,N_6412,N_6010);
and U6788 (N_6788,N_6292,N_6207);
and U6789 (N_6789,N_6322,N_6085);
and U6790 (N_6790,N_6315,N_6203);
nand U6791 (N_6791,N_6302,N_6237);
xor U6792 (N_6792,N_6048,N_6195);
or U6793 (N_6793,N_6129,N_6191);
and U6794 (N_6794,N_6417,N_6413);
xnor U6795 (N_6795,N_6432,N_6120);
xor U6796 (N_6796,N_6026,N_6044);
and U6797 (N_6797,N_6445,N_6134);
nor U6798 (N_6798,N_6492,N_6038);
nand U6799 (N_6799,N_6061,N_6427);
xnor U6800 (N_6800,N_6148,N_6064);
xnor U6801 (N_6801,N_6043,N_6152);
and U6802 (N_6802,N_6282,N_6406);
and U6803 (N_6803,N_6095,N_6075);
nor U6804 (N_6804,N_6136,N_6311);
nor U6805 (N_6805,N_6400,N_6323);
nand U6806 (N_6806,N_6318,N_6406);
nand U6807 (N_6807,N_6486,N_6370);
and U6808 (N_6808,N_6477,N_6133);
and U6809 (N_6809,N_6254,N_6444);
xnor U6810 (N_6810,N_6088,N_6078);
nor U6811 (N_6811,N_6272,N_6312);
xnor U6812 (N_6812,N_6249,N_6000);
or U6813 (N_6813,N_6093,N_6294);
or U6814 (N_6814,N_6154,N_6261);
xor U6815 (N_6815,N_6113,N_6007);
nand U6816 (N_6816,N_6391,N_6446);
nand U6817 (N_6817,N_6388,N_6238);
nor U6818 (N_6818,N_6053,N_6027);
nor U6819 (N_6819,N_6153,N_6303);
nand U6820 (N_6820,N_6265,N_6287);
xnor U6821 (N_6821,N_6140,N_6480);
or U6822 (N_6822,N_6237,N_6377);
or U6823 (N_6823,N_6445,N_6192);
and U6824 (N_6824,N_6437,N_6369);
xor U6825 (N_6825,N_6234,N_6455);
nor U6826 (N_6826,N_6490,N_6248);
xnor U6827 (N_6827,N_6049,N_6417);
nand U6828 (N_6828,N_6328,N_6260);
nor U6829 (N_6829,N_6252,N_6065);
nand U6830 (N_6830,N_6035,N_6363);
nand U6831 (N_6831,N_6254,N_6268);
nor U6832 (N_6832,N_6124,N_6480);
and U6833 (N_6833,N_6343,N_6268);
xor U6834 (N_6834,N_6300,N_6456);
nor U6835 (N_6835,N_6357,N_6379);
nand U6836 (N_6836,N_6178,N_6323);
xor U6837 (N_6837,N_6478,N_6137);
xor U6838 (N_6838,N_6197,N_6446);
or U6839 (N_6839,N_6405,N_6297);
nand U6840 (N_6840,N_6299,N_6109);
and U6841 (N_6841,N_6076,N_6395);
nand U6842 (N_6842,N_6333,N_6212);
nor U6843 (N_6843,N_6015,N_6050);
or U6844 (N_6844,N_6482,N_6494);
and U6845 (N_6845,N_6216,N_6475);
nand U6846 (N_6846,N_6004,N_6273);
or U6847 (N_6847,N_6070,N_6085);
nor U6848 (N_6848,N_6316,N_6416);
nor U6849 (N_6849,N_6250,N_6477);
and U6850 (N_6850,N_6051,N_6251);
nand U6851 (N_6851,N_6008,N_6331);
and U6852 (N_6852,N_6064,N_6213);
and U6853 (N_6853,N_6152,N_6273);
nor U6854 (N_6854,N_6341,N_6201);
nor U6855 (N_6855,N_6255,N_6039);
and U6856 (N_6856,N_6222,N_6124);
nand U6857 (N_6857,N_6395,N_6473);
nor U6858 (N_6858,N_6252,N_6383);
or U6859 (N_6859,N_6012,N_6013);
nand U6860 (N_6860,N_6094,N_6072);
nor U6861 (N_6861,N_6304,N_6052);
or U6862 (N_6862,N_6483,N_6251);
nand U6863 (N_6863,N_6395,N_6413);
and U6864 (N_6864,N_6038,N_6300);
nor U6865 (N_6865,N_6440,N_6332);
or U6866 (N_6866,N_6333,N_6073);
xor U6867 (N_6867,N_6297,N_6045);
or U6868 (N_6868,N_6273,N_6412);
and U6869 (N_6869,N_6359,N_6019);
or U6870 (N_6870,N_6043,N_6034);
or U6871 (N_6871,N_6153,N_6269);
nor U6872 (N_6872,N_6499,N_6068);
and U6873 (N_6873,N_6117,N_6498);
xor U6874 (N_6874,N_6322,N_6434);
and U6875 (N_6875,N_6092,N_6286);
and U6876 (N_6876,N_6053,N_6485);
nor U6877 (N_6877,N_6010,N_6099);
nand U6878 (N_6878,N_6111,N_6245);
nand U6879 (N_6879,N_6230,N_6289);
nor U6880 (N_6880,N_6083,N_6058);
nand U6881 (N_6881,N_6202,N_6271);
nor U6882 (N_6882,N_6395,N_6280);
nand U6883 (N_6883,N_6224,N_6276);
or U6884 (N_6884,N_6367,N_6341);
and U6885 (N_6885,N_6173,N_6032);
or U6886 (N_6886,N_6080,N_6148);
nor U6887 (N_6887,N_6313,N_6325);
or U6888 (N_6888,N_6394,N_6271);
xnor U6889 (N_6889,N_6364,N_6316);
nor U6890 (N_6890,N_6054,N_6107);
nor U6891 (N_6891,N_6081,N_6265);
or U6892 (N_6892,N_6408,N_6076);
nor U6893 (N_6893,N_6475,N_6258);
xnor U6894 (N_6894,N_6069,N_6209);
or U6895 (N_6895,N_6174,N_6394);
nor U6896 (N_6896,N_6394,N_6426);
nor U6897 (N_6897,N_6157,N_6458);
nand U6898 (N_6898,N_6017,N_6139);
or U6899 (N_6899,N_6485,N_6214);
nand U6900 (N_6900,N_6369,N_6395);
and U6901 (N_6901,N_6384,N_6088);
nand U6902 (N_6902,N_6345,N_6458);
or U6903 (N_6903,N_6438,N_6170);
or U6904 (N_6904,N_6007,N_6305);
or U6905 (N_6905,N_6186,N_6112);
or U6906 (N_6906,N_6124,N_6437);
xnor U6907 (N_6907,N_6066,N_6394);
nor U6908 (N_6908,N_6090,N_6327);
nand U6909 (N_6909,N_6011,N_6441);
nand U6910 (N_6910,N_6341,N_6387);
or U6911 (N_6911,N_6276,N_6457);
nand U6912 (N_6912,N_6300,N_6112);
or U6913 (N_6913,N_6169,N_6422);
nand U6914 (N_6914,N_6416,N_6296);
xor U6915 (N_6915,N_6278,N_6406);
nor U6916 (N_6916,N_6288,N_6357);
and U6917 (N_6917,N_6120,N_6020);
xnor U6918 (N_6918,N_6011,N_6436);
or U6919 (N_6919,N_6097,N_6321);
xor U6920 (N_6920,N_6424,N_6418);
and U6921 (N_6921,N_6350,N_6307);
or U6922 (N_6922,N_6198,N_6374);
or U6923 (N_6923,N_6178,N_6183);
nor U6924 (N_6924,N_6123,N_6411);
xor U6925 (N_6925,N_6103,N_6031);
and U6926 (N_6926,N_6275,N_6193);
xor U6927 (N_6927,N_6113,N_6066);
nor U6928 (N_6928,N_6044,N_6299);
and U6929 (N_6929,N_6413,N_6378);
and U6930 (N_6930,N_6283,N_6372);
nand U6931 (N_6931,N_6357,N_6361);
nor U6932 (N_6932,N_6257,N_6349);
xor U6933 (N_6933,N_6032,N_6285);
and U6934 (N_6934,N_6050,N_6172);
xnor U6935 (N_6935,N_6141,N_6121);
xor U6936 (N_6936,N_6142,N_6283);
nor U6937 (N_6937,N_6372,N_6067);
and U6938 (N_6938,N_6184,N_6251);
xnor U6939 (N_6939,N_6414,N_6402);
or U6940 (N_6940,N_6065,N_6086);
and U6941 (N_6941,N_6261,N_6015);
or U6942 (N_6942,N_6222,N_6033);
or U6943 (N_6943,N_6416,N_6357);
nand U6944 (N_6944,N_6028,N_6298);
nor U6945 (N_6945,N_6162,N_6200);
nand U6946 (N_6946,N_6370,N_6281);
nor U6947 (N_6947,N_6237,N_6423);
nand U6948 (N_6948,N_6334,N_6373);
nor U6949 (N_6949,N_6085,N_6170);
and U6950 (N_6950,N_6035,N_6229);
nor U6951 (N_6951,N_6187,N_6048);
xnor U6952 (N_6952,N_6126,N_6291);
xor U6953 (N_6953,N_6386,N_6417);
xnor U6954 (N_6954,N_6376,N_6130);
and U6955 (N_6955,N_6276,N_6211);
nand U6956 (N_6956,N_6397,N_6081);
nor U6957 (N_6957,N_6151,N_6213);
xor U6958 (N_6958,N_6106,N_6486);
and U6959 (N_6959,N_6001,N_6316);
or U6960 (N_6960,N_6067,N_6270);
and U6961 (N_6961,N_6052,N_6183);
nand U6962 (N_6962,N_6194,N_6474);
nor U6963 (N_6963,N_6483,N_6122);
xor U6964 (N_6964,N_6422,N_6377);
and U6965 (N_6965,N_6467,N_6244);
or U6966 (N_6966,N_6337,N_6184);
xnor U6967 (N_6967,N_6280,N_6137);
and U6968 (N_6968,N_6096,N_6221);
nor U6969 (N_6969,N_6362,N_6088);
and U6970 (N_6970,N_6250,N_6022);
or U6971 (N_6971,N_6137,N_6364);
nor U6972 (N_6972,N_6158,N_6050);
xor U6973 (N_6973,N_6107,N_6315);
nor U6974 (N_6974,N_6035,N_6289);
nor U6975 (N_6975,N_6223,N_6209);
or U6976 (N_6976,N_6169,N_6070);
xor U6977 (N_6977,N_6057,N_6364);
or U6978 (N_6978,N_6264,N_6238);
and U6979 (N_6979,N_6148,N_6107);
nor U6980 (N_6980,N_6168,N_6048);
and U6981 (N_6981,N_6488,N_6169);
or U6982 (N_6982,N_6291,N_6010);
nand U6983 (N_6983,N_6050,N_6180);
nand U6984 (N_6984,N_6474,N_6299);
and U6985 (N_6985,N_6112,N_6416);
nor U6986 (N_6986,N_6414,N_6374);
nand U6987 (N_6987,N_6040,N_6256);
or U6988 (N_6988,N_6388,N_6114);
nor U6989 (N_6989,N_6499,N_6347);
or U6990 (N_6990,N_6388,N_6205);
xor U6991 (N_6991,N_6080,N_6232);
xnor U6992 (N_6992,N_6190,N_6205);
and U6993 (N_6993,N_6379,N_6285);
and U6994 (N_6994,N_6047,N_6458);
nand U6995 (N_6995,N_6275,N_6098);
nor U6996 (N_6996,N_6034,N_6051);
nor U6997 (N_6997,N_6246,N_6457);
nand U6998 (N_6998,N_6259,N_6106);
nand U6999 (N_6999,N_6160,N_6356);
nor U7000 (N_7000,N_6687,N_6764);
or U7001 (N_7001,N_6632,N_6866);
nand U7002 (N_7002,N_6539,N_6574);
nand U7003 (N_7003,N_6993,N_6942);
nor U7004 (N_7004,N_6703,N_6535);
xor U7005 (N_7005,N_6858,N_6540);
and U7006 (N_7006,N_6718,N_6874);
xnor U7007 (N_7007,N_6810,N_6926);
and U7008 (N_7008,N_6900,N_6946);
nor U7009 (N_7009,N_6629,N_6607);
and U7010 (N_7010,N_6784,N_6705);
or U7011 (N_7011,N_6627,N_6508);
and U7012 (N_7012,N_6511,N_6735);
and U7013 (N_7013,N_6948,N_6725);
xor U7014 (N_7014,N_6967,N_6904);
or U7015 (N_7015,N_6702,N_6956);
nand U7016 (N_7016,N_6851,N_6815);
or U7017 (N_7017,N_6595,N_6700);
xnor U7018 (N_7018,N_6988,N_6786);
nand U7019 (N_7019,N_6545,N_6501);
nor U7020 (N_7020,N_6892,N_6800);
or U7021 (N_7021,N_6562,N_6543);
xor U7022 (N_7022,N_6576,N_6751);
or U7023 (N_7023,N_6662,N_6594);
or U7024 (N_7024,N_6925,N_6955);
and U7025 (N_7025,N_6997,N_6531);
and U7026 (N_7026,N_6612,N_6526);
nand U7027 (N_7027,N_6914,N_6623);
nand U7028 (N_7028,N_6585,N_6773);
and U7029 (N_7029,N_6869,N_6610);
nor U7030 (N_7030,N_6709,N_6748);
xnor U7031 (N_7031,N_6514,N_6555);
nand U7032 (N_7032,N_6845,N_6846);
or U7033 (N_7033,N_6990,N_6986);
or U7034 (N_7034,N_6583,N_6536);
nor U7035 (N_7035,N_6631,N_6852);
nand U7036 (N_7036,N_6947,N_6621);
or U7037 (N_7037,N_6935,N_6516);
xor U7038 (N_7038,N_6762,N_6877);
or U7039 (N_7039,N_6575,N_6927);
nor U7040 (N_7040,N_6564,N_6818);
xor U7041 (N_7041,N_6635,N_6593);
nor U7042 (N_7042,N_6847,N_6739);
nor U7043 (N_7043,N_6596,N_6519);
or U7044 (N_7044,N_6711,N_6777);
or U7045 (N_7045,N_6512,N_6968);
nor U7046 (N_7046,N_6868,N_6862);
xor U7047 (N_7047,N_6626,N_6738);
nor U7048 (N_7048,N_6654,N_6671);
xor U7049 (N_7049,N_6857,N_6999);
xor U7050 (N_7050,N_6683,N_6776);
and U7051 (N_7051,N_6833,N_6680);
nand U7052 (N_7052,N_6779,N_6672);
or U7053 (N_7053,N_6691,N_6812);
and U7054 (N_7054,N_6592,N_6550);
and U7055 (N_7055,N_6951,N_6697);
xor U7056 (N_7056,N_6600,N_6970);
xor U7057 (N_7057,N_6732,N_6809);
or U7058 (N_7058,N_6641,N_6775);
or U7059 (N_7059,N_6766,N_6532);
xor U7060 (N_7060,N_6880,N_6832);
nand U7061 (N_7061,N_6974,N_6601);
nor U7062 (N_7062,N_6538,N_6878);
and U7063 (N_7063,N_6996,N_6941);
or U7064 (N_7064,N_6888,N_6876);
nand U7065 (N_7065,N_6677,N_6843);
or U7066 (N_7066,N_6782,N_6588);
nand U7067 (N_7067,N_6799,N_6960);
and U7068 (N_7068,N_6571,N_6890);
nand U7069 (N_7069,N_6681,N_6811);
and U7070 (N_7070,N_6903,N_6840);
or U7071 (N_7071,N_6989,N_6765);
xnor U7072 (N_7072,N_6597,N_6917);
and U7073 (N_7073,N_6673,N_6885);
nor U7074 (N_7074,N_6790,N_6801);
nor U7075 (N_7075,N_6909,N_6906);
and U7076 (N_7076,N_6805,N_6905);
and U7077 (N_7077,N_6769,N_6894);
or U7078 (N_7078,N_6870,N_6728);
xnor U7079 (N_7079,N_6643,N_6613);
and U7080 (N_7080,N_6850,N_6838);
nand U7081 (N_7081,N_6922,N_6618);
and U7082 (N_7082,N_6675,N_6882);
or U7083 (N_7083,N_6648,N_6723);
xor U7084 (N_7084,N_6579,N_6754);
nor U7085 (N_7085,N_6736,N_6706);
nand U7086 (N_7086,N_6837,N_6695);
nand U7087 (N_7087,N_6761,N_6789);
nor U7088 (N_7088,N_6568,N_6507);
xnor U7089 (N_7089,N_6994,N_6864);
xnor U7090 (N_7090,N_6759,N_6740);
and U7091 (N_7091,N_6821,N_6528);
nor U7092 (N_7092,N_6551,N_6676);
nand U7093 (N_7093,N_6795,N_6983);
xor U7094 (N_7094,N_6721,N_6717);
xnor U7095 (N_7095,N_6642,N_6719);
or U7096 (N_7096,N_6533,N_6685);
and U7097 (N_7097,N_6756,N_6659);
xnor U7098 (N_7098,N_6856,N_6558);
and U7099 (N_7099,N_6586,N_6502);
nand U7100 (N_7100,N_6932,N_6791);
nor U7101 (N_7101,N_6940,N_6962);
xor U7102 (N_7102,N_6710,N_6669);
xor U7103 (N_7103,N_6745,N_6911);
nand U7104 (N_7104,N_6844,N_6954);
nand U7105 (N_7105,N_6933,N_6901);
and U7106 (N_7106,N_6908,N_6729);
nand U7107 (N_7107,N_6806,N_6943);
nand U7108 (N_7108,N_6660,N_6871);
or U7109 (N_7109,N_6663,N_6981);
nor U7110 (N_7110,N_6615,N_6645);
and U7111 (N_7111,N_6887,N_6608);
nor U7112 (N_7112,N_6820,N_6853);
nand U7113 (N_7113,N_6835,N_6547);
xnor U7114 (N_7114,N_6658,N_6804);
and U7115 (N_7115,N_6860,N_6918);
and U7116 (N_7116,N_6763,N_6966);
and U7117 (N_7117,N_6733,N_6572);
or U7118 (N_7118,N_6639,N_6848);
nor U7119 (N_7119,N_6854,N_6530);
and U7120 (N_7120,N_6792,N_6771);
nand U7121 (N_7121,N_6505,N_6823);
xnor U7122 (N_7122,N_6578,N_6861);
or U7123 (N_7123,N_6923,N_6529);
xor U7124 (N_7124,N_6737,N_6628);
or U7125 (N_7125,N_6549,N_6573);
nor U7126 (N_7126,N_6541,N_6670);
nor U7127 (N_7127,N_6873,N_6916);
nor U7128 (N_7128,N_6743,N_6715);
or U7129 (N_7129,N_6624,N_6666);
nor U7130 (N_7130,N_6965,N_6783);
nor U7131 (N_7131,N_6686,N_6750);
nand U7132 (N_7132,N_6749,N_6696);
nand U7133 (N_7133,N_6652,N_6712);
nand U7134 (N_7134,N_6824,N_6977);
nand U7135 (N_7135,N_6650,N_6826);
nor U7136 (N_7136,N_6734,N_6865);
and U7137 (N_7137,N_6938,N_6972);
or U7138 (N_7138,N_6638,N_6598);
nor U7139 (N_7139,N_6544,N_6552);
xnor U7140 (N_7140,N_6995,N_6836);
xor U7141 (N_7141,N_6537,N_6839);
nand U7142 (N_7142,N_6611,N_6982);
nand U7143 (N_7143,N_6500,N_6570);
or U7144 (N_7144,N_6655,N_6971);
or U7145 (N_7145,N_6863,N_6707);
or U7146 (N_7146,N_6580,N_6620);
and U7147 (N_7147,N_6699,N_6602);
or U7148 (N_7148,N_6859,N_6684);
nand U7149 (N_7149,N_6559,N_6726);
xnor U7150 (N_7150,N_6931,N_6920);
nand U7151 (N_7151,N_6637,N_6730);
or U7152 (N_7152,N_6523,N_6930);
xor U7153 (N_7153,N_6589,N_6958);
nor U7154 (N_7154,N_6963,N_6757);
nand U7155 (N_7155,N_6944,N_6849);
nand U7156 (N_7156,N_6649,N_6599);
nor U7157 (N_7157,N_6991,N_6979);
nand U7158 (N_7158,N_6661,N_6886);
or U7159 (N_7159,N_6924,N_6636);
and U7160 (N_7160,N_6975,N_6959);
nand U7161 (N_7161,N_6557,N_6945);
nor U7162 (N_7162,N_6778,N_6912);
and U7163 (N_7163,N_6692,N_6964);
nor U7164 (N_7164,N_6919,N_6875);
or U7165 (N_7165,N_6881,N_6542);
and U7166 (N_7166,N_6617,N_6554);
or U7167 (N_7167,N_6814,N_6741);
nor U7168 (N_7168,N_6679,N_6828);
nand U7169 (N_7169,N_6755,N_6622);
xnor U7170 (N_7170,N_6998,N_6504);
nand U7171 (N_7171,N_6668,N_6774);
xor U7172 (N_7172,N_6934,N_6582);
nor U7173 (N_7173,N_6802,N_6907);
nand U7174 (N_7174,N_6605,N_6506);
or U7175 (N_7175,N_6758,N_6803);
and U7176 (N_7176,N_6902,N_6665);
or U7177 (N_7177,N_6704,N_6604);
and U7178 (N_7178,N_6744,N_6794);
xnor U7179 (N_7179,N_6560,N_6656);
or U7180 (N_7180,N_6807,N_6829);
nor U7181 (N_7181,N_6816,N_6587);
nand U7182 (N_7182,N_6952,N_6522);
or U7183 (N_7183,N_6788,N_6752);
xnor U7184 (N_7184,N_6682,N_6567);
and U7185 (N_7185,N_6978,N_6513);
nor U7186 (N_7186,N_6898,N_6614);
or U7187 (N_7187,N_6831,N_6722);
nand U7188 (N_7188,N_6842,N_6834);
or U7189 (N_7189,N_6561,N_6796);
nand U7190 (N_7190,N_6770,N_6524);
nor U7191 (N_7191,N_6724,N_6563);
and U7192 (N_7192,N_6780,N_6969);
nor U7193 (N_7193,N_6813,N_6891);
and U7194 (N_7194,N_6961,N_6694);
xnor U7195 (N_7195,N_6644,N_6581);
and U7196 (N_7196,N_6984,N_6667);
and U7197 (N_7197,N_6872,N_6760);
and U7198 (N_7198,N_6584,N_6577);
xnor U7199 (N_7199,N_6785,N_6553);
xnor U7200 (N_7200,N_6515,N_6913);
nor U7201 (N_7201,N_6619,N_6548);
and U7202 (N_7202,N_6787,N_6950);
and U7203 (N_7203,N_6767,N_6727);
nor U7204 (N_7204,N_6630,N_6742);
or U7205 (N_7205,N_6503,N_6896);
nor U7206 (N_7206,N_6937,N_6753);
and U7207 (N_7207,N_6616,N_6693);
nand U7208 (N_7208,N_6713,N_6746);
or U7209 (N_7209,N_6698,N_6899);
or U7210 (N_7210,N_6651,N_6509);
nand U7211 (N_7211,N_6939,N_6985);
nand U7212 (N_7212,N_6520,N_6678);
or U7213 (N_7213,N_6867,N_6830);
nand U7214 (N_7214,N_6714,N_6591);
xor U7215 (N_7215,N_6731,N_6772);
nor U7216 (N_7216,N_6657,N_6664);
nand U7217 (N_7217,N_6716,N_6590);
xor U7218 (N_7218,N_6521,N_6747);
nor U7219 (N_7219,N_6897,N_6936);
or U7220 (N_7220,N_6976,N_6688);
nand U7221 (N_7221,N_6546,N_6781);
nand U7222 (N_7222,N_6603,N_6634);
or U7223 (N_7223,N_6708,N_6825);
xor U7224 (N_7224,N_6953,N_6609);
or U7225 (N_7225,N_6987,N_6768);
xor U7226 (N_7226,N_6566,N_6674);
or U7227 (N_7227,N_6841,N_6633);
nor U7228 (N_7228,N_6690,N_6653);
nor U7229 (N_7229,N_6879,N_6973);
xor U7230 (N_7230,N_6895,N_6793);
nand U7231 (N_7231,N_6525,N_6915);
or U7232 (N_7232,N_6949,N_6646);
nor U7233 (N_7233,N_6534,N_6817);
and U7234 (N_7234,N_6510,N_6910);
and U7235 (N_7235,N_6798,N_6893);
or U7236 (N_7236,N_6928,N_6647);
nand U7237 (N_7237,N_6855,N_6797);
and U7238 (N_7238,N_6889,N_6689);
nor U7239 (N_7239,N_6720,N_6921);
and U7240 (N_7240,N_6929,N_6819);
or U7241 (N_7241,N_6517,N_6518);
nor U7242 (N_7242,N_6701,N_6992);
nand U7243 (N_7243,N_6827,N_6957);
nand U7244 (N_7244,N_6569,N_6822);
xor U7245 (N_7245,N_6640,N_6565);
nor U7246 (N_7246,N_6980,N_6556);
and U7247 (N_7247,N_6884,N_6527);
xor U7248 (N_7248,N_6606,N_6883);
xnor U7249 (N_7249,N_6808,N_6625);
nor U7250 (N_7250,N_6918,N_6914);
or U7251 (N_7251,N_6948,N_6781);
or U7252 (N_7252,N_6950,N_6561);
xor U7253 (N_7253,N_6996,N_6500);
nor U7254 (N_7254,N_6588,N_6713);
and U7255 (N_7255,N_6644,N_6584);
nor U7256 (N_7256,N_6752,N_6803);
xnor U7257 (N_7257,N_6901,N_6980);
or U7258 (N_7258,N_6982,N_6906);
nand U7259 (N_7259,N_6987,N_6549);
nand U7260 (N_7260,N_6748,N_6809);
and U7261 (N_7261,N_6859,N_6959);
xnor U7262 (N_7262,N_6981,N_6936);
or U7263 (N_7263,N_6796,N_6530);
xor U7264 (N_7264,N_6675,N_6749);
xor U7265 (N_7265,N_6821,N_6558);
xnor U7266 (N_7266,N_6924,N_6756);
or U7267 (N_7267,N_6505,N_6971);
nand U7268 (N_7268,N_6602,N_6598);
xor U7269 (N_7269,N_6856,N_6850);
and U7270 (N_7270,N_6920,N_6749);
and U7271 (N_7271,N_6966,N_6768);
and U7272 (N_7272,N_6684,N_6784);
and U7273 (N_7273,N_6697,N_6536);
and U7274 (N_7274,N_6533,N_6850);
xnor U7275 (N_7275,N_6695,N_6613);
nand U7276 (N_7276,N_6726,N_6703);
xor U7277 (N_7277,N_6988,N_6602);
and U7278 (N_7278,N_6859,N_6553);
or U7279 (N_7279,N_6776,N_6989);
or U7280 (N_7280,N_6525,N_6946);
and U7281 (N_7281,N_6722,N_6661);
nand U7282 (N_7282,N_6935,N_6839);
and U7283 (N_7283,N_6761,N_6525);
xnor U7284 (N_7284,N_6632,N_6672);
or U7285 (N_7285,N_6871,N_6625);
or U7286 (N_7286,N_6793,N_6911);
nor U7287 (N_7287,N_6620,N_6730);
and U7288 (N_7288,N_6626,N_6784);
and U7289 (N_7289,N_6948,N_6754);
nor U7290 (N_7290,N_6672,N_6520);
xnor U7291 (N_7291,N_6524,N_6768);
and U7292 (N_7292,N_6983,N_6740);
xnor U7293 (N_7293,N_6973,N_6730);
and U7294 (N_7294,N_6717,N_6742);
and U7295 (N_7295,N_6632,N_6681);
xnor U7296 (N_7296,N_6604,N_6685);
or U7297 (N_7297,N_6838,N_6504);
and U7298 (N_7298,N_6659,N_6963);
nor U7299 (N_7299,N_6851,N_6962);
xnor U7300 (N_7300,N_6821,N_6515);
and U7301 (N_7301,N_6760,N_6904);
or U7302 (N_7302,N_6533,N_6979);
xnor U7303 (N_7303,N_6574,N_6933);
or U7304 (N_7304,N_6586,N_6572);
nor U7305 (N_7305,N_6801,N_6973);
nand U7306 (N_7306,N_6863,N_6924);
nor U7307 (N_7307,N_6759,N_6529);
nor U7308 (N_7308,N_6648,N_6877);
or U7309 (N_7309,N_6820,N_6935);
nand U7310 (N_7310,N_6533,N_6501);
nand U7311 (N_7311,N_6643,N_6795);
and U7312 (N_7312,N_6735,N_6948);
nand U7313 (N_7313,N_6591,N_6764);
nor U7314 (N_7314,N_6642,N_6875);
and U7315 (N_7315,N_6606,N_6634);
and U7316 (N_7316,N_6915,N_6904);
xnor U7317 (N_7317,N_6880,N_6905);
xnor U7318 (N_7318,N_6858,N_6628);
and U7319 (N_7319,N_6982,N_6525);
and U7320 (N_7320,N_6543,N_6510);
and U7321 (N_7321,N_6796,N_6533);
or U7322 (N_7322,N_6843,N_6513);
nand U7323 (N_7323,N_6641,N_6908);
xor U7324 (N_7324,N_6627,N_6726);
nand U7325 (N_7325,N_6646,N_6690);
nand U7326 (N_7326,N_6943,N_6634);
nor U7327 (N_7327,N_6751,N_6589);
nand U7328 (N_7328,N_6659,N_6880);
xor U7329 (N_7329,N_6544,N_6857);
nor U7330 (N_7330,N_6740,N_6814);
or U7331 (N_7331,N_6678,N_6884);
xor U7332 (N_7332,N_6757,N_6986);
and U7333 (N_7333,N_6626,N_6692);
xnor U7334 (N_7334,N_6795,N_6511);
nor U7335 (N_7335,N_6581,N_6796);
or U7336 (N_7336,N_6750,N_6949);
or U7337 (N_7337,N_6608,N_6598);
nor U7338 (N_7338,N_6514,N_6885);
or U7339 (N_7339,N_6597,N_6721);
nand U7340 (N_7340,N_6697,N_6637);
nand U7341 (N_7341,N_6539,N_6997);
and U7342 (N_7342,N_6715,N_6920);
xor U7343 (N_7343,N_6999,N_6726);
nor U7344 (N_7344,N_6854,N_6921);
xor U7345 (N_7345,N_6669,N_6570);
or U7346 (N_7346,N_6525,N_6564);
nor U7347 (N_7347,N_6740,N_6571);
xor U7348 (N_7348,N_6588,N_6798);
xor U7349 (N_7349,N_6954,N_6969);
or U7350 (N_7350,N_6918,N_6569);
nor U7351 (N_7351,N_6775,N_6672);
and U7352 (N_7352,N_6969,N_6635);
or U7353 (N_7353,N_6566,N_6801);
nand U7354 (N_7354,N_6757,N_6896);
and U7355 (N_7355,N_6890,N_6954);
xnor U7356 (N_7356,N_6970,N_6815);
or U7357 (N_7357,N_6834,N_6799);
and U7358 (N_7358,N_6573,N_6806);
or U7359 (N_7359,N_6680,N_6939);
nand U7360 (N_7360,N_6786,N_6617);
xnor U7361 (N_7361,N_6906,N_6788);
or U7362 (N_7362,N_6512,N_6770);
xor U7363 (N_7363,N_6841,N_6664);
xor U7364 (N_7364,N_6577,N_6803);
nand U7365 (N_7365,N_6944,N_6660);
nand U7366 (N_7366,N_6722,N_6909);
and U7367 (N_7367,N_6967,N_6702);
or U7368 (N_7368,N_6652,N_6867);
xnor U7369 (N_7369,N_6647,N_6757);
or U7370 (N_7370,N_6891,N_6642);
nand U7371 (N_7371,N_6734,N_6855);
nand U7372 (N_7372,N_6532,N_6510);
nor U7373 (N_7373,N_6934,N_6997);
nand U7374 (N_7374,N_6775,N_6676);
nor U7375 (N_7375,N_6866,N_6761);
xor U7376 (N_7376,N_6744,N_6534);
or U7377 (N_7377,N_6805,N_6628);
nor U7378 (N_7378,N_6987,N_6592);
xnor U7379 (N_7379,N_6886,N_6729);
and U7380 (N_7380,N_6507,N_6692);
nand U7381 (N_7381,N_6714,N_6845);
xor U7382 (N_7382,N_6841,N_6933);
xnor U7383 (N_7383,N_6883,N_6727);
and U7384 (N_7384,N_6581,N_6719);
and U7385 (N_7385,N_6770,N_6901);
nand U7386 (N_7386,N_6577,N_6749);
xnor U7387 (N_7387,N_6869,N_6618);
xor U7388 (N_7388,N_6528,N_6937);
xor U7389 (N_7389,N_6659,N_6692);
and U7390 (N_7390,N_6505,N_6789);
or U7391 (N_7391,N_6549,N_6749);
nor U7392 (N_7392,N_6571,N_6522);
xnor U7393 (N_7393,N_6561,N_6761);
and U7394 (N_7394,N_6734,N_6693);
nand U7395 (N_7395,N_6602,N_6654);
nand U7396 (N_7396,N_6875,N_6910);
and U7397 (N_7397,N_6980,N_6914);
or U7398 (N_7398,N_6698,N_6516);
nand U7399 (N_7399,N_6863,N_6626);
and U7400 (N_7400,N_6889,N_6937);
nand U7401 (N_7401,N_6826,N_6854);
and U7402 (N_7402,N_6942,N_6715);
and U7403 (N_7403,N_6764,N_6816);
xor U7404 (N_7404,N_6834,N_6685);
and U7405 (N_7405,N_6795,N_6670);
xnor U7406 (N_7406,N_6882,N_6783);
nand U7407 (N_7407,N_6588,N_6987);
nand U7408 (N_7408,N_6638,N_6810);
nand U7409 (N_7409,N_6539,N_6534);
nor U7410 (N_7410,N_6922,N_6578);
xor U7411 (N_7411,N_6812,N_6845);
or U7412 (N_7412,N_6526,N_6932);
or U7413 (N_7413,N_6863,N_6860);
or U7414 (N_7414,N_6513,N_6800);
nor U7415 (N_7415,N_6865,N_6910);
xnor U7416 (N_7416,N_6676,N_6559);
and U7417 (N_7417,N_6833,N_6540);
xor U7418 (N_7418,N_6936,N_6788);
xor U7419 (N_7419,N_6579,N_6516);
xor U7420 (N_7420,N_6902,N_6931);
nand U7421 (N_7421,N_6880,N_6791);
nor U7422 (N_7422,N_6606,N_6948);
xnor U7423 (N_7423,N_6859,N_6528);
nand U7424 (N_7424,N_6846,N_6983);
xnor U7425 (N_7425,N_6882,N_6824);
xnor U7426 (N_7426,N_6751,N_6667);
nand U7427 (N_7427,N_6740,N_6833);
xor U7428 (N_7428,N_6659,N_6944);
nand U7429 (N_7429,N_6760,N_6700);
xnor U7430 (N_7430,N_6680,N_6933);
or U7431 (N_7431,N_6554,N_6569);
nand U7432 (N_7432,N_6620,N_6741);
xor U7433 (N_7433,N_6706,N_6829);
xnor U7434 (N_7434,N_6598,N_6763);
xnor U7435 (N_7435,N_6743,N_6934);
and U7436 (N_7436,N_6992,N_6998);
xor U7437 (N_7437,N_6518,N_6966);
and U7438 (N_7438,N_6696,N_6873);
xnor U7439 (N_7439,N_6699,N_6889);
nand U7440 (N_7440,N_6978,N_6627);
or U7441 (N_7441,N_6530,N_6532);
and U7442 (N_7442,N_6601,N_6578);
or U7443 (N_7443,N_6964,N_6742);
xor U7444 (N_7444,N_6723,N_6605);
or U7445 (N_7445,N_6632,N_6933);
nor U7446 (N_7446,N_6735,N_6730);
xnor U7447 (N_7447,N_6742,N_6697);
and U7448 (N_7448,N_6594,N_6575);
nand U7449 (N_7449,N_6518,N_6863);
and U7450 (N_7450,N_6577,N_6581);
and U7451 (N_7451,N_6693,N_6566);
or U7452 (N_7452,N_6822,N_6591);
nor U7453 (N_7453,N_6772,N_6671);
nand U7454 (N_7454,N_6910,N_6712);
nor U7455 (N_7455,N_6821,N_6789);
nor U7456 (N_7456,N_6943,N_6694);
nand U7457 (N_7457,N_6990,N_6810);
nor U7458 (N_7458,N_6835,N_6598);
nand U7459 (N_7459,N_6904,N_6894);
and U7460 (N_7460,N_6983,N_6746);
nand U7461 (N_7461,N_6586,N_6870);
and U7462 (N_7462,N_6568,N_6542);
and U7463 (N_7463,N_6614,N_6948);
nor U7464 (N_7464,N_6559,N_6563);
nor U7465 (N_7465,N_6699,N_6949);
nand U7466 (N_7466,N_6774,N_6824);
xnor U7467 (N_7467,N_6914,N_6839);
nand U7468 (N_7468,N_6755,N_6981);
and U7469 (N_7469,N_6886,N_6639);
nand U7470 (N_7470,N_6667,N_6825);
and U7471 (N_7471,N_6568,N_6526);
xor U7472 (N_7472,N_6845,N_6559);
nor U7473 (N_7473,N_6511,N_6724);
or U7474 (N_7474,N_6625,N_6663);
and U7475 (N_7475,N_6575,N_6611);
nor U7476 (N_7476,N_6620,N_6793);
nor U7477 (N_7477,N_6860,N_6853);
nand U7478 (N_7478,N_6855,N_6857);
or U7479 (N_7479,N_6605,N_6695);
and U7480 (N_7480,N_6949,N_6633);
nor U7481 (N_7481,N_6574,N_6601);
or U7482 (N_7482,N_6500,N_6791);
nor U7483 (N_7483,N_6933,N_6554);
nor U7484 (N_7484,N_6980,N_6557);
xnor U7485 (N_7485,N_6757,N_6705);
xor U7486 (N_7486,N_6916,N_6983);
xor U7487 (N_7487,N_6526,N_6965);
nor U7488 (N_7488,N_6677,N_6987);
xnor U7489 (N_7489,N_6561,N_6584);
or U7490 (N_7490,N_6862,N_6619);
and U7491 (N_7491,N_6759,N_6845);
xnor U7492 (N_7492,N_6925,N_6890);
xnor U7493 (N_7493,N_6590,N_6601);
nor U7494 (N_7494,N_6767,N_6992);
nand U7495 (N_7495,N_6842,N_6679);
nand U7496 (N_7496,N_6843,N_6516);
nand U7497 (N_7497,N_6994,N_6948);
nor U7498 (N_7498,N_6558,N_6742);
nor U7499 (N_7499,N_6996,N_6900);
nor U7500 (N_7500,N_7057,N_7477);
xnor U7501 (N_7501,N_7064,N_7379);
nand U7502 (N_7502,N_7149,N_7200);
or U7503 (N_7503,N_7278,N_7122);
and U7504 (N_7504,N_7013,N_7193);
xnor U7505 (N_7505,N_7382,N_7042);
nor U7506 (N_7506,N_7053,N_7160);
and U7507 (N_7507,N_7267,N_7047);
xor U7508 (N_7508,N_7484,N_7299);
xor U7509 (N_7509,N_7380,N_7217);
nand U7510 (N_7510,N_7405,N_7227);
nand U7511 (N_7511,N_7207,N_7082);
nand U7512 (N_7512,N_7445,N_7449);
and U7513 (N_7513,N_7376,N_7220);
and U7514 (N_7514,N_7451,N_7408);
nor U7515 (N_7515,N_7367,N_7325);
nand U7516 (N_7516,N_7173,N_7269);
or U7517 (N_7517,N_7184,N_7462);
and U7518 (N_7518,N_7113,N_7457);
nand U7519 (N_7519,N_7355,N_7192);
or U7520 (N_7520,N_7322,N_7313);
nand U7521 (N_7521,N_7212,N_7010);
nand U7522 (N_7522,N_7273,N_7389);
nand U7523 (N_7523,N_7438,N_7170);
nand U7524 (N_7524,N_7168,N_7241);
xnor U7525 (N_7525,N_7097,N_7260);
nor U7526 (N_7526,N_7134,N_7485);
or U7527 (N_7527,N_7056,N_7252);
nand U7528 (N_7528,N_7225,N_7307);
nor U7529 (N_7529,N_7391,N_7132);
or U7530 (N_7530,N_7282,N_7338);
xnor U7531 (N_7531,N_7377,N_7371);
and U7532 (N_7532,N_7480,N_7343);
and U7533 (N_7533,N_7366,N_7312);
nand U7534 (N_7534,N_7300,N_7060);
xnor U7535 (N_7535,N_7345,N_7319);
and U7536 (N_7536,N_7027,N_7100);
or U7537 (N_7537,N_7142,N_7265);
xnor U7538 (N_7538,N_7394,N_7250);
and U7539 (N_7539,N_7178,N_7197);
or U7540 (N_7540,N_7246,N_7350);
xnor U7541 (N_7541,N_7206,N_7049);
and U7542 (N_7542,N_7404,N_7364);
nor U7543 (N_7543,N_7009,N_7413);
or U7544 (N_7544,N_7439,N_7453);
nor U7545 (N_7545,N_7198,N_7456);
and U7546 (N_7546,N_7141,N_7043);
nand U7547 (N_7547,N_7335,N_7234);
xor U7548 (N_7548,N_7428,N_7257);
nand U7549 (N_7549,N_7023,N_7357);
xnor U7550 (N_7550,N_7336,N_7317);
nor U7551 (N_7551,N_7432,N_7497);
and U7552 (N_7552,N_7481,N_7196);
nor U7553 (N_7553,N_7446,N_7492);
nor U7554 (N_7554,N_7420,N_7264);
nand U7555 (N_7555,N_7067,N_7085);
nand U7556 (N_7556,N_7116,N_7020);
xnor U7557 (N_7557,N_7486,N_7240);
xor U7558 (N_7558,N_7354,N_7008);
nor U7559 (N_7559,N_7424,N_7383);
and U7560 (N_7560,N_7172,N_7219);
nand U7561 (N_7561,N_7393,N_7466);
nand U7562 (N_7562,N_7223,N_7140);
and U7563 (N_7563,N_7344,N_7414);
or U7564 (N_7564,N_7275,N_7150);
nor U7565 (N_7565,N_7059,N_7187);
nand U7566 (N_7566,N_7084,N_7174);
xor U7567 (N_7567,N_7330,N_7123);
and U7568 (N_7568,N_7270,N_7297);
and U7569 (N_7569,N_7306,N_7255);
xnor U7570 (N_7570,N_7320,N_7417);
nor U7571 (N_7571,N_7179,N_7156);
and U7572 (N_7572,N_7163,N_7069);
and U7573 (N_7573,N_7055,N_7472);
or U7574 (N_7574,N_7024,N_7396);
nor U7575 (N_7575,N_7347,N_7327);
xor U7576 (N_7576,N_7155,N_7012);
xor U7577 (N_7577,N_7274,N_7211);
or U7578 (N_7578,N_7426,N_7044);
and U7579 (N_7579,N_7189,N_7128);
nand U7580 (N_7580,N_7136,N_7215);
nand U7581 (N_7581,N_7133,N_7406);
and U7582 (N_7582,N_7348,N_7321);
nor U7583 (N_7583,N_7054,N_7353);
and U7584 (N_7584,N_7291,N_7425);
nor U7585 (N_7585,N_7440,N_7034);
xor U7586 (N_7586,N_7068,N_7016);
xor U7587 (N_7587,N_7304,N_7106);
and U7588 (N_7588,N_7203,N_7071);
nand U7589 (N_7589,N_7434,N_7450);
nand U7590 (N_7590,N_7375,N_7052);
and U7591 (N_7591,N_7369,N_7103);
or U7592 (N_7592,N_7385,N_7118);
nand U7593 (N_7593,N_7421,N_7422);
xnor U7594 (N_7594,N_7473,N_7022);
and U7595 (N_7595,N_7259,N_7311);
nand U7596 (N_7596,N_7239,N_7237);
or U7597 (N_7597,N_7469,N_7062);
nor U7598 (N_7598,N_7229,N_7114);
nor U7599 (N_7599,N_7111,N_7018);
nand U7600 (N_7600,N_7152,N_7230);
and U7601 (N_7601,N_7104,N_7416);
nor U7602 (N_7602,N_7323,N_7045);
nand U7603 (N_7603,N_7251,N_7436);
nor U7604 (N_7604,N_7400,N_7146);
xnor U7605 (N_7605,N_7268,N_7315);
and U7606 (N_7606,N_7046,N_7188);
or U7607 (N_7607,N_7444,N_7475);
nor U7608 (N_7608,N_7295,N_7249);
xnor U7609 (N_7609,N_7094,N_7078);
nand U7610 (N_7610,N_7096,N_7226);
xor U7611 (N_7611,N_7148,N_7166);
xor U7612 (N_7612,N_7063,N_7147);
xnor U7613 (N_7613,N_7429,N_7002);
xnor U7614 (N_7614,N_7177,N_7041);
xor U7615 (N_7615,N_7289,N_7489);
xor U7616 (N_7616,N_7075,N_7356);
nand U7617 (N_7617,N_7331,N_7247);
xor U7618 (N_7618,N_7037,N_7143);
xnor U7619 (N_7619,N_7244,N_7138);
nand U7620 (N_7620,N_7387,N_7081);
or U7621 (N_7621,N_7105,N_7488);
nand U7622 (N_7622,N_7032,N_7388);
or U7623 (N_7623,N_7093,N_7216);
nor U7624 (N_7624,N_7459,N_7378);
nand U7625 (N_7625,N_7029,N_7190);
and U7626 (N_7626,N_7410,N_7452);
nor U7627 (N_7627,N_7169,N_7314);
nand U7628 (N_7628,N_7340,N_7460);
xnor U7629 (N_7629,N_7030,N_7126);
xnor U7630 (N_7630,N_7154,N_7242);
or U7631 (N_7631,N_7231,N_7474);
or U7632 (N_7632,N_7341,N_7271);
and U7633 (N_7633,N_7194,N_7339);
and U7634 (N_7634,N_7007,N_7415);
xnor U7635 (N_7635,N_7115,N_7205);
xnor U7636 (N_7636,N_7175,N_7125);
xnor U7637 (N_7637,N_7153,N_7080);
or U7638 (N_7638,N_7083,N_7272);
and U7639 (N_7639,N_7427,N_7235);
or U7640 (N_7640,N_7491,N_7158);
nand U7641 (N_7641,N_7442,N_7435);
nor U7642 (N_7642,N_7066,N_7487);
nand U7643 (N_7643,N_7108,N_7232);
nor U7644 (N_7644,N_7465,N_7296);
xor U7645 (N_7645,N_7015,N_7333);
and U7646 (N_7646,N_7281,N_7411);
or U7647 (N_7647,N_7092,N_7395);
or U7648 (N_7648,N_7003,N_7361);
and U7649 (N_7649,N_7162,N_7471);
nor U7650 (N_7650,N_7039,N_7076);
nor U7651 (N_7651,N_7233,N_7329);
nor U7652 (N_7652,N_7455,N_7352);
nand U7653 (N_7653,N_7004,N_7384);
xor U7654 (N_7654,N_7180,N_7431);
nor U7655 (N_7655,N_7334,N_7412);
and U7656 (N_7656,N_7458,N_7483);
xor U7657 (N_7657,N_7266,N_7099);
xnor U7658 (N_7658,N_7280,N_7470);
nand U7659 (N_7659,N_7326,N_7072);
nand U7660 (N_7660,N_7409,N_7145);
and U7661 (N_7661,N_7351,N_7031);
nor U7662 (N_7662,N_7171,N_7358);
nor U7663 (N_7663,N_7495,N_7493);
and U7664 (N_7664,N_7496,N_7129);
or U7665 (N_7665,N_7107,N_7224);
xor U7666 (N_7666,N_7137,N_7028);
nand U7667 (N_7667,N_7077,N_7363);
or U7668 (N_7668,N_7119,N_7074);
nor U7669 (N_7669,N_7437,N_7310);
or U7670 (N_7670,N_7176,N_7430);
xnor U7671 (N_7671,N_7308,N_7290);
nor U7672 (N_7672,N_7288,N_7324);
or U7673 (N_7673,N_7183,N_7318);
xor U7674 (N_7674,N_7468,N_7478);
and U7675 (N_7675,N_7245,N_7098);
and U7676 (N_7676,N_7276,N_7441);
and U7677 (N_7677,N_7127,N_7418);
xnor U7678 (N_7678,N_7464,N_7112);
nor U7679 (N_7679,N_7087,N_7258);
nor U7680 (N_7680,N_7204,N_7403);
nor U7681 (N_7681,N_7236,N_7397);
xnor U7682 (N_7682,N_7359,N_7337);
nor U7683 (N_7683,N_7228,N_7167);
or U7684 (N_7684,N_7135,N_7293);
xnor U7685 (N_7685,N_7316,N_7292);
nor U7686 (N_7686,N_7482,N_7342);
and U7687 (N_7687,N_7349,N_7017);
or U7688 (N_7688,N_7121,N_7368);
xnor U7689 (N_7689,N_7284,N_7243);
xor U7690 (N_7690,N_7365,N_7201);
and U7691 (N_7691,N_7101,N_7423);
nor U7692 (N_7692,N_7181,N_7286);
and U7693 (N_7693,N_7253,N_7301);
and U7694 (N_7694,N_7210,N_7399);
nand U7695 (N_7695,N_7443,N_7185);
xnor U7696 (N_7696,N_7089,N_7157);
nand U7697 (N_7697,N_7014,N_7130);
and U7698 (N_7698,N_7195,N_7011);
or U7699 (N_7699,N_7191,N_7360);
or U7700 (N_7700,N_7209,N_7305);
nor U7701 (N_7701,N_7025,N_7079);
and U7702 (N_7702,N_7499,N_7479);
nor U7703 (N_7703,N_7287,N_7033);
and U7704 (N_7704,N_7373,N_7117);
xnor U7705 (N_7705,N_7221,N_7498);
and U7706 (N_7706,N_7494,N_7139);
xnor U7707 (N_7707,N_7222,N_7238);
and U7708 (N_7708,N_7454,N_7102);
nand U7709 (N_7709,N_7065,N_7303);
and U7710 (N_7710,N_7256,N_7447);
nor U7711 (N_7711,N_7309,N_7254);
or U7712 (N_7712,N_7298,N_7277);
and U7713 (N_7713,N_7261,N_7159);
or U7714 (N_7714,N_7164,N_7285);
xnor U7715 (N_7715,N_7419,N_7021);
and U7716 (N_7716,N_7073,N_7109);
xnor U7717 (N_7717,N_7263,N_7402);
and U7718 (N_7718,N_7302,N_7058);
nand U7719 (N_7719,N_7213,N_7202);
nor U7720 (N_7720,N_7248,N_7433);
nand U7721 (N_7721,N_7398,N_7199);
nor U7722 (N_7722,N_7131,N_7332);
or U7723 (N_7723,N_7461,N_7000);
nand U7724 (N_7724,N_7144,N_7086);
xor U7725 (N_7725,N_7294,N_7040);
nor U7726 (N_7726,N_7088,N_7005);
nor U7727 (N_7727,N_7182,N_7390);
nand U7728 (N_7728,N_7038,N_7048);
nor U7729 (N_7729,N_7346,N_7476);
or U7730 (N_7730,N_7463,N_7124);
nand U7731 (N_7731,N_7467,N_7186);
xor U7732 (N_7732,N_7448,N_7161);
nand U7733 (N_7733,N_7151,N_7401);
and U7734 (N_7734,N_7362,N_7392);
xor U7735 (N_7735,N_7374,N_7050);
and U7736 (N_7736,N_7407,N_7001);
nor U7737 (N_7737,N_7208,N_7091);
nor U7738 (N_7738,N_7214,N_7283);
or U7739 (N_7739,N_7051,N_7386);
or U7740 (N_7740,N_7370,N_7218);
and U7741 (N_7741,N_7006,N_7036);
nor U7742 (N_7742,N_7019,N_7165);
xor U7743 (N_7743,N_7279,N_7490);
xor U7744 (N_7744,N_7095,N_7090);
xor U7745 (N_7745,N_7035,N_7381);
and U7746 (N_7746,N_7110,N_7026);
nor U7747 (N_7747,N_7372,N_7070);
nor U7748 (N_7748,N_7120,N_7262);
xnor U7749 (N_7749,N_7061,N_7328);
xnor U7750 (N_7750,N_7295,N_7346);
and U7751 (N_7751,N_7433,N_7083);
xnor U7752 (N_7752,N_7049,N_7327);
xnor U7753 (N_7753,N_7415,N_7476);
xor U7754 (N_7754,N_7324,N_7046);
and U7755 (N_7755,N_7228,N_7218);
and U7756 (N_7756,N_7237,N_7304);
nor U7757 (N_7757,N_7349,N_7019);
or U7758 (N_7758,N_7426,N_7292);
and U7759 (N_7759,N_7471,N_7098);
and U7760 (N_7760,N_7287,N_7303);
nor U7761 (N_7761,N_7242,N_7089);
nor U7762 (N_7762,N_7160,N_7168);
or U7763 (N_7763,N_7317,N_7055);
and U7764 (N_7764,N_7482,N_7043);
nor U7765 (N_7765,N_7101,N_7191);
or U7766 (N_7766,N_7324,N_7028);
nor U7767 (N_7767,N_7295,N_7314);
xnor U7768 (N_7768,N_7288,N_7259);
or U7769 (N_7769,N_7064,N_7060);
or U7770 (N_7770,N_7485,N_7098);
or U7771 (N_7771,N_7460,N_7293);
and U7772 (N_7772,N_7123,N_7378);
and U7773 (N_7773,N_7195,N_7330);
or U7774 (N_7774,N_7484,N_7201);
or U7775 (N_7775,N_7442,N_7376);
nand U7776 (N_7776,N_7067,N_7209);
xor U7777 (N_7777,N_7482,N_7022);
and U7778 (N_7778,N_7170,N_7155);
xnor U7779 (N_7779,N_7453,N_7008);
nor U7780 (N_7780,N_7270,N_7080);
nor U7781 (N_7781,N_7140,N_7118);
nand U7782 (N_7782,N_7037,N_7460);
nor U7783 (N_7783,N_7489,N_7442);
xor U7784 (N_7784,N_7114,N_7149);
nor U7785 (N_7785,N_7381,N_7084);
or U7786 (N_7786,N_7391,N_7490);
and U7787 (N_7787,N_7412,N_7268);
and U7788 (N_7788,N_7262,N_7027);
and U7789 (N_7789,N_7118,N_7164);
nor U7790 (N_7790,N_7270,N_7301);
nor U7791 (N_7791,N_7452,N_7362);
or U7792 (N_7792,N_7047,N_7017);
and U7793 (N_7793,N_7324,N_7417);
xor U7794 (N_7794,N_7403,N_7438);
xnor U7795 (N_7795,N_7485,N_7138);
or U7796 (N_7796,N_7409,N_7174);
xnor U7797 (N_7797,N_7265,N_7209);
or U7798 (N_7798,N_7209,N_7327);
nor U7799 (N_7799,N_7200,N_7009);
and U7800 (N_7800,N_7270,N_7268);
nand U7801 (N_7801,N_7086,N_7366);
or U7802 (N_7802,N_7112,N_7398);
or U7803 (N_7803,N_7181,N_7000);
or U7804 (N_7804,N_7170,N_7369);
xor U7805 (N_7805,N_7478,N_7201);
or U7806 (N_7806,N_7201,N_7273);
nand U7807 (N_7807,N_7114,N_7401);
and U7808 (N_7808,N_7253,N_7071);
nor U7809 (N_7809,N_7351,N_7181);
and U7810 (N_7810,N_7259,N_7364);
xnor U7811 (N_7811,N_7003,N_7307);
xnor U7812 (N_7812,N_7303,N_7041);
xnor U7813 (N_7813,N_7274,N_7234);
or U7814 (N_7814,N_7467,N_7063);
or U7815 (N_7815,N_7378,N_7365);
or U7816 (N_7816,N_7423,N_7230);
and U7817 (N_7817,N_7173,N_7381);
nand U7818 (N_7818,N_7249,N_7138);
xor U7819 (N_7819,N_7432,N_7495);
and U7820 (N_7820,N_7392,N_7087);
nand U7821 (N_7821,N_7253,N_7157);
xor U7822 (N_7822,N_7351,N_7024);
nand U7823 (N_7823,N_7159,N_7233);
nor U7824 (N_7824,N_7426,N_7269);
nor U7825 (N_7825,N_7164,N_7186);
and U7826 (N_7826,N_7466,N_7185);
nor U7827 (N_7827,N_7003,N_7188);
nor U7828 (N_7828,N_7306,N_7302);
or U7829 (N_7829,N_7344,N_7443);
or U7830 (N_7830,N_7139,N_7142);
xnor U7831 (N_7831,N_7307,N_7354);
nor U7832 (N_7832,N_7077,N_7464);
xor U7833 (N_7833,N_7405,N_7341);
and U7834 (N_7834,N_7300,N_7125);
xor U7835 (N_7835,N_7078,N_7019);
nand U7836 (N_7836,N_7327,N_7296);
nand U7837 (N_7837,N_7408,N_7268);
or U7838 (N_7838,N_7174,N_7269);
and U7839 (N_7839,N_7110,N_7249);
nor U7840 (N_7840,N_7301,N_7408);
nand U7841 (N_7841,N_7138,N_7368);
and U7842 (N_7842,N_7031,N_7409);
or U7843 (N_7843,N_7402,N_7126);
and U7844 (N_7844,N_7328,N_7311);
nand U7845 (N_7845,N_7367,N_7390);
nor U7846 (N_7846,N_7336,N_7377);
xnor U7847 (N_7847,N_7487,N_7416);
nor U7848 (N_7848,N_7394,N_7213);
nand U7849 (N_7849,N_7183,N_7249);
or U7850 (N_7850,N_7444,N_7397);
and U7851 (N_7851,N_7148,N_7214);
xor U7852 (N_7852,N_7496,N_7274);
nor U7853 (N_7853,N_7393,N_7054);
and U7854 (N_7854,N_7028,N_7372);
or U7855 (N_7855,N_7024,N_7248);
and U7856 (N_7856,N_7172,N_7036);
nand U7857 (N_7857,N_7174,N_7320);
nand U7858 (N_7858,N_7060,N_7183);
nand U7859 (N_7859,N_7499,N_7485);
or U7860 (N_7860,N_7230,N_7209);
nor U7861 (N_7861,N_7246,N_7303);
nand U7862 (N_7862,N_7418,N_7115);
nor U7863 (N_7863,N_7331,N_7304);
and U7864 (N_7864,N_7009,N_7375);
xnor U7865 (N_7865,N_7142,N_7324);
nand U7866 (N_7866,N_7178,N_7074);
xor U7867 (N_7867,N_7321,N_7436);
nor U7868 (N_7868,N_7403,N_7120);
and U7869 (N_7869,N_7083,N_7469);
nand U7870 (N_7870,N_7264,N_7419);
or U7871 (N_7871,N_7016,N_7345);
nor U7872 (N_7872,N_7181,N_7337);
or U7873 (N_7873,N_7213,N_7280);
and U7874 (N_7874,N_7485,N_7089);
nor U7875 (N_7875,N_7141,N_7437);
xnor U7876 (N_7876,N_7470,N_7328);
and U7877 (N_7877,N_7257,N_7165);
nor U7878 (N_7878,N_7123,N_7246);
xnor U7879 (N_7879,N_7019,N_7296);
or U7880 (N_7880,N_7120,N_7269);
or U7881 (N_7881,N_7017,N_7079);
nand U7882 (N_7882,N_7285,N_7392);
nand U7883 (N_7883,N_7302,N_7101);
and U7884 (N_7884,N_7337,N_7434);
nor U7885 (N_7885,N_7277,N_7306);
nand U7886 (N_7886,N_7090,N_7094);
and U7887 (N_7887,N_7011,N_7417);
and U7888 (N_7888,N_7088,N_7036);
xor U7889 (N_7889,N_7041,N_7015);
or U7890 (N_7890,N_7196,N_7150);
xnor U7891 (N_7891,N_7393,N_7375);
or U7892 (N_7892,N_7171,N_7343);
and U7893 (N_7893,N_7164,N_7064);
xor U7894 (N_7894,N_7087,N_7319);
or U7895 (N_7895,N_7372,N_7495);
nor U7896 (N_7896,N_7041,N_7014);
xor U7897 (N_7897,N_7286,N_7137);
nor U7898 (N_7898,N_7082,N_7395);
xor U7899 (N_7899,N_7037,N_7016);
nand U7900 (N_7900,N_7387,N_7184);
nor U7901 (N_7901,N_7410,N_7132);
and U7902 (N_7902,N_7017,N_7248);
nor U7903 (N_7903,N_7080,N_7330);
nand U7904 (N_7904,N_7274,N_7127);
nor U7905 (N_7905,N_7386,N_7125);
xnor U7906 (N_7906,N_7225,N_7260);
or U7907 (N_7907,N_7082,N_7038);
nand U7908 (N_7908,N_7002,N_7124);
and U7909 (N_7909,N_7278,N_7491);
or U7910 (N_7910,N_7035,N_7162);
or U7911 (N_7911,N_7104,N_7216);
or U7912 (N_7912,N_7465,N_7284);
and U7913 (N_7913,N_7008,N_7040);
nor U7914 (N_7914,N_7475,N_7478);
nand U7915 (N_7915,N_7456,N_7053);
nand U7916 (N_7916,N_7199,N_7242);
xor U7917 (N_7917,N_7129,N_7205);
nand U7918 (N_7918,N_7152,N_7089);
or U7919 (N_7919,N_7034,N_7480);
and U7920 (N_7920,N_7088,N_7238);
or U7921 (N_7921,N_7105,N_7454);
nor U7922 (N_7922,N_7423,N_7445);
xor U7923 (N_7923,N_7008,N_7361);
xnor U7924 (N_7924,N_7215,N_7380);
nor U7925 (N_7925,N_7125,N_7161);
nor U7926 (N_7926,N_7094,N_7342);
or U7927 (N_7927,N_7376,N_7247);
nand U7928 (N_7928,N_7451,N_7092);
nor U7929 (N_7929,N_7346,N_7157);
nor U7930 (N_7930,N_7130,N_7400);
xnor U7931 (N_7931,N_7253,N_7199);
and U7932 (N_7932,N_7142,N_7052);
or U7933 (N_7933,N_7152,N_7318);
xor U7934 (N_7934,N_7485,N_7157);
nand U7935 (N_7935,N_7291,N_7097);
or U7936 (N_7936,N_7292,N_7207);
nand U7937 (N_7937,N_7205,N_7223);
xnor U7938 (N_7938,N_7458,N_7474);
xor U7939 (N_7939,N_7168,N_7055);
nor U7940 (N_7940,N_7090,N_7450);
and U7941 (N_7941,N_7168,N_7376);
nand U7942 (N_7942,N_7328,N_7462);
nand U7943 (N_7943,N_7213,N_7045);
or U7944 (N_7944,N_7069,N_7436);
nand U7945 (N_7945,N_7230,N_7268);
nor U7946 (N_7946,N_7206,N_7041);
or U7947 (N_7947,N_7179,N_7132);
and U7948 (N_7948,N_7277,N_7194);
and U7949 (N_7949,N_7089,N_7052);
or U7950 (N_7950,N_7360,N_7012);
or U7951 (N_7951,N_7144,N_7271);
nand U7952 (N_7952,N_7234,N_7210);
nand U7953 (N_7953,N_7184,N_7149);
nor U7954 (N_7954,N_7063,N_7342);
nand U7955 (N_7955,N_7471,N_7220);
xnor U7956 (N_7956,N_7381,N_7174);
nand U7957 (N_7957,N_7149,N_7407);
and U7958 (N_7958,N_7065,N_7391);
or U7959 (N_7959,N_7435,N_7307);
nor U7960 (N_7960,N_7432,N_7421);
nand U7961 (N_7961,N_7161,N_7383);
or U7962 (N_7962,N_7335,N_7071);
or U7963 (N_7963,N_7120,N_7418);
nand U7964 (N_7964,N_7161,N_7366);
xor U7965 (N_7965,N_7045,N_7170);
and U7966 (N_7966,N_7068,N_7370);
or U7967 (N_7967,N_7229,N_7275);
and U7968 (N_7968,N_7029,N_7495);
xor U7969 (N_7969,N_7258,N_7379);
and U7970 (N_7970,N_7083,N_7419);
xnor U7971 (N_7971,N_7285,N_7238);
xor U7972 (N_7972,N_7017,N_7444);
nor U7973 (N_7973,N_7340,N_7344);
nor U7974 (N_7974,N_7488,N_7168);
and U7975 (N_7975,N_7069,N_7455);
or U7976 (N_7976,N_7487,N_7208);
and U7977 (N_7977,N_7251,N_7148);
nor U7978 (N_7978,N_7464,N_7427);
nand U7979 (N_7979,N_7460,N_7493);
xor U7980 (N_7980,N_7083,N_7263);
nand U7981 (N_7981,N_7217,N_7479);
or U7982 (N_7982,N_7044,N_7137);
xor U7983 (N_7983,N_7047,N_7145);
xnor U7984 (N_7984,N_7448,N_7085);
nor U7985 (N_7985,N_7389,N_7371);
nand U7986 (N_7986,N_7231,N_7371);
and U7987 (N_7987,N_7359,N_7101);
or U7988 (N_7988,N_7376,N_7311);
xor U7989 (N_7989,N_7494,N_7492);
and U7990 (N_7990,N_7054,N_7099);
and U7991 (N_7991,N_7090,N_7240);
or U7992 (N_7992,N_7310,N_7435);
nor U7993 (N_7993,N_7207,N_7276);
or U7994 (N_7994,N_7446,N_7491);
or U7995 (N_7995,N_7497,N_7361);
and U7996 (N_7996,N_7402,N_7376);
nand U7997 (N_7997,N_7257,N_7158);
nor U7998 (N_7998,N_7165,N_7321);
nand U7999 (N_7999,N_7368,N_7456);
nand U8000 (N_8000,N_7948,N_7986);
and U8001 (N_8001,N_7654,N_7985);
nor U8002 (N_8002,N_7576,N_7844);
xor U8003 (N_8003,N_7624,N_7561);
xor U8004 (N_8004,N_7510,N_7688);
nor U8005 (N_8005,N_7863,N_7501);
nand U8006 (N_8006,N_7993,N_7586);
nand U8007 (N_8007,N_7583,N_7822);
or U8008 (N_8008,N_7771,N_7996);
or U8009 (N_8009,N_7836,N_7689);
or U8010 (N_8010,N_7871,N_7710);
or U8011 (N_8011,N_7641,N_7912);
and U8012 (N_8012,N_7678,N_7803);
and U8013 (N_8013,N_7589,N_7626);
and U8014 (N_8014,N_7747,N_7782);
nor U8015 (N_8015,N_7659,N_7954);
nand U8016 (N_8016,N_7698,N_7828);
nor U8017 (N_8017,N_7770,N_7581);
xor U8018 (N_8018,N_7570,N_7804);
or U8019 (N_8019,N_7805,N_7965);
and U8020 (N_8020,N_7646,N_7702);
xor U8021 (N_8021,N_7753,N_7612);
and U8022 (N_8022,N_7566,N_7787);
or U8023 (N_8023,N_7604,N_7521);
xor U8024 (N_8024,N_7642,N_7931);
xor U8025 (N_8025,N_7914,N_7731);
and U8026 (N_8026,N_7904,N_7736);
or U8027 (N_8027,N_7503,N_7826);
or U8028 (N_8028,N_7667,N_7808);
xnor U8029 (N_8029,N_7830,N_7937);
nand U8030 (N_8030,N_7725,N_7979);
nor U8031 (N_8031,N_7956,N_7973);
xor U8032 (N_8032,N_7567,N_7728);
xor U8033 (N_8033,N_7673,N_7706);
xnor U8034 (N_8034,N_7898,N_7674);
xnor U8035 (N_8035,N_7866,N_7927);
nor U8036 (N_8036,N_7950,N_7640);
xor U8037 (N_8037,N_7661,N_7941);
xor U8038 (N_8038,N_7902,N_7969);
and U8039 (N_8039,N_7686,N_7707);
nor U8040 (N_8040,N_7764,N_7504);
nand U8041 (N_8041,N_7621,N_7655);
nor U8042 (N_8042,N_7798,N_7638);
nor U8043 (N_8043,N_7629,N_7718);
xnor U8044 (N_8044,N_7639,N_7681);
nand U8045 (N_8045,N_7568,N_7806);
and U8046 (N_8046,N_7799,N_7729);
and U8047 (N_8047,N_7645,N_7522);
and U8048 (N_8048,N_7683,N_7978);
nor U8049 (N_8049,N_7769,N_7574);
nand U8050 (N_8050,N_7597,N_7989);
or U8051 (N_8051,N_7716,N_7607);
and U8052 (N_8052,N_7824,N_7974);
nor U8053 (N_8053,N_7953,N_7915);
xnor U8054 (N_8054,N_7745,N_7852);
nand U8055 (N_8055,N_7881,N_7890);
or U8056 (N_8056,N_7858,N_7791);
nand U8057 (N_8057,N_7773,N_7947);
and U8058 (N_8058,N_7529,N_7619);
or U8059 (N_8059,N_7699,N_7991);
xnor U8060 (N_8060,N_7899,N_7610);
xnor U8061 (N_8061,N_7740,N_7651);
and U8062 (N_8062,N_7869,N_7872);
xnor U8063 (N_8063,N_7853,N_7943);
xor U8064 (N_8064,N_7841,N_7783);
and U8065 (N_8065,N_7860,N_7809);
xnor U8066 (N_8066,N_7896,N_7967);
nand U8067 (N_8067,N_7755,N_7992);
nand U8068 (N_8068,N_7870,N_7751);
nor U8069 (N_8069,N_7560,N_7559);
xor U8070 (N_8070,N_7682,N_7821);
xor U8071 (N_8071,N_7971,N_7823);
or U8072 (N_8072,N_7905,N_7526);
or U8073 (N_8073,N_7994,N_7593);
nor U8074 (N_8074,N_7935,N_7636);
nor U8075 (N_8075,N_7724,N_7648);
nor U8076 (N_8076,N_7932,N_7502);
nor U8077 (N_8077,N_7835,N_7656);
nand U8078 (N_8078,N_7889,N_7572);
nor U8079 (N_8079,N_7776,N_7837);
and U8080 (N_8080,N_7917,N_7720);
and U8081 (N_8081,N_7714,N_7712);
nor U8082 (N_8082,N_7670,N_7966);
and U8083 (N_8083,N_7876,N_7602);
nor U8084 (N_8084,N_7553,N_7977);
nand U8085 (N_8085,N_7664,N_7634);
and U8086 (N_8086,N_7558,N_7882);
and U8087 (N_8087,N_7705,N_7756);
and U8088 (N_8088,N_7925,N_7878);
nor U8089 (N_8089,N_7868,N_7691);
and U8090 (N_8090,N_7669,N_7605);
nor U8091 (N_8091,N_7980,N_7732);
and U8092 (N_8092,N_7894,N_7792);
nand U8093 (N_8093,N_7573,N_7883);
nor U8094 (N_8094,N_7891,N_7599);
nor U8095 (N_8095,N_7800,N_7834);
and U8096 (N_8096,N_7831,N_7535);
and U8097 (N_8097,N_7666,N_7509);
nand U8098 (N_8098,N_7617,N_7812);
or U8099 (N_8099,N_7672,N_7671);
nor U8100 (N_8100,N_7608,N_7532);
xor U8101 (N_8101,N_7508,N_7960);
or U8102 (N_8102,N_7820,N_7727);
nand U8103 (N_8103,N_7913,N_7713);
or U8104 (N_8104,N_7926,N_7500);
xnor U8105 (N_8105,N_7680,N_7909);
nor U8106 (N_8106,N_7539,N_7722);
and U8107 (N_8107,N_7518,N_7923);
and U8108 (N_8108,N_7520,N_7797);
and U8109 (N_8109,N_7892,N_7613);
nor U8110 (N_8110,N_7657,N_7995);
or U8111 (N_8111,N_7571,N_7693);
or U8112 (N_8112,N_7949,N_7877);
and U8113 (N_8113,N_7616,N_7611);
nand U8114 (N_8114,N_7957,N_7708);
xor U8115 (N_8115,N_7647,N_7848);
or U8116 (N_8116,N_7507,N_7939);
nor U8117 (N_8117,N_7684,N_7748);
xnor U8118 (N_8118,N_7859,N_7794);
nor U8119 (N_8119,N_7580,N_7793);
xnor U8120 (N_8120,N_7813,N_7506);
xnor U8121 (N_8121,N_7660,N_7744);
xnor U8122 (N_8122,N_7505,N_7554);
nand U8123 (N_8123,N_7903,N_7885);
and U8124 (N_8124,N_7735,N_7919);
nor U8125 (N_8125,N_7618,N_7582);
or U8126 (N_8126,N_7615,N_7845);
and U8127 (N_8127,N_7763,N_7785);
or U8128 (N_8128,N_7998,N_7513);
nor U8129 (N_8129,N_7726,N_7528);
nor U8130 (N_8130,N_7862,N_7677);
or U8131 (N_8131,N_7694,N_7697);
or U8132 (N_8132,N_7757,N_7850);
nor U8133 (N_8133,N_7746,N_7623);
nand U8134 (N_8134,N_7983,N_7741);
nor U8135 (N_8135,N_7940,N_7700);
nand U8136 (N_8136,N_7537,N_7635);
nor U8137 (N_8137,N_7517,N_7833);
or U8138 (N_8138,N_7864,N_7933);
nor U8139 (N_8139,N_7564,N_7955);
and U8140 (N_8140,N_7970,N_7814);
nand U8141 (N_8141,N_7603,N_7695);
or U8142 (N_8142,N_7542,N_7591);
or U8143 (N_8143,N_7665,N_7963);
nor U8144 (N_8144,N_7644,N_7901);
xnor U8145 (N_8145,N_7704,N_7622);
nand U8146 (N_8146,N_7873,N_7549);
and U8147 (N_8147,N_7779,N_7551);
and U8148 (N_8148,N_7911,N_7907);
or U8149 (N_8149,N_7649,N_7762);
or U8150 (N_8150,N_7690,N_7525);
nor U8151 (N_8151,N_7592,N_7816);
and U8152 (N_8152,N_7633,N_7918);
or U8153 (N_8153,N_7723,N_7847);
nor U8154 (N_8154,N_7897,N_7719);
or U8155 (N_8155,N_7675,N_7575);
or U8156 (N_8156,N_7938,N_7679);
and U8157 (N_8157,N_7880,N_7772);
xnor U8158 (N_8158,N_7990,N_7865);
xnor U8159 (N_8159,N_7587,N_7766);
xor U8160 (N_8160,N_7565,N_7817);
xnor U8161 (N_8161,N_7851,N_7668);
and U8162 (N_8162,N_7606,N_7921);
nand U8163 (N_8163,N_7854,N_7519);
or U8164 (N_8164,N_7879,N_7934);
nand U8165 (N_8165,N_7534,N_7999);
nand U8166 (N_8166,N_7839,N_7569);
nor U8167 (N_8167,N_7768,N_7936);
nor U8168 (N_8168,N_7964,N_7596);
and U8169 (N_8169,N_7924,N_7540);
or U8170 (N_8170,N_7961,N_7663);
and U8171 (N_8171,N_7631,N_7951);
or U8172 (N_8172,N_7795,N_7846);
or U8173 (N_8173,N_7658,N_7536);
nand U8174 (N_8174,N_7562,N_7818);
nand U8175 (N_8175,N_7516,N_7584);
nand U8176 (N_8176,N_7550,N_7546);
nand U8177 (N_8177,N_7662,N_7538);
nand U8178 (N_8178,N_7984,N_7777);
or U8179 (N_8179,N_7531,N_7895);
xnor U8180 (N_8180,N_7888,N_7588);
xor U8181 (N_8181,N_7737,N_7721);
nand U8182 (N_8182,N_7887,N_7547);
and U8183 (N_8183,N_7595,N_7832);
xnor U8184 (N_8184,N_7807,N_7555);
nor U8185 (N_8185,N_7819,N_7856);
or U8186 (N_8186,N_7650,N_7838);
nor U8187 (N_8187,N_7515,N_7563);
nand U8188 (N_8188,N_7544,N_7743);
xor U8189 (N_8189,N_7976,N_7527);
nand U8190 (N_8190,N_7778,N_7717);
or U8191 (N_8191,N_7545,N_7676);
and U8192 (N_8192,N_7930,N_7796);
and U8193 (N_8193,N_7598,N_7780);
xnor U8194 (N_8194,N_7692,N_7715);
nand U8195 (N_8195,N_7758,N_7774);
nor U8196 (N_8196,N_7908,N_7946);
nand U8197 (N_8197,N_7750,N_7742);
xor U8198 (N_8198,N_7761,N_7942);
and U8199 (N_8199,N_7801,N_7514);
nand U8200 (N_8200,N_7653,N_7579);
or U8201 (N_8201,N_7524,N_7637);
xor U8202 (N_8202,N_7600,N_7767);
nor U8203 (N_8203,N_7533,N_7614);
nor U8204 (N_8204,N_7685,N_7512);
xnor U8205 (N_8205,N_7701,N_7988);
xnor U8206 (N_8206,N_7781,N_7875);
or U8207 (N_8207,N_7944,N_7749);
and U8208 (N_8208,N_7825,N_7906);
xor U8209 (N_8209,N_7541,N_7815);
and U8210 (N_8210,N_7530,N_7959);
and U8211 (N_8211,N_7789,N_7916);
and U8212 (N_8212,N_7703,N_7929);
or U8213 (N_8213,N_7855,N_7975);
or U8214 (N_8214,N_7543,N_7687);
nand U8215 (N_8215,N_7696,N_7958);
xnor U8216 (N_8216,N_7552,N_7628);
nand U8217 (N_8217,N_7594,N_7557);
xor U8218 (N_8218,N_7620,N_7754);
or U8219 (N_8219,N_7952,N_7920);
nor U8220 (N_8220,N_7861,N_7738);
nand U8221 (N_8221,N_7752,N_7625);
nand U8222 (N_8222,N_7627,N_7968);
or U8223 (N_8223,N_7730,N_7811);
and U8224 (N_8224,N_7786,N_7802);
nor U8225 (N_8225,N_7733,N_7827);
nand U8226 (N_8226,N_7981,N_7577);
or U8227 (N_8227,N_7857,N_7945);
nand U8228 (N_8228,N_7711,N_7849);
xnor U8229 (N_8229,N_7893,N_7734);
nor U8230 (N_8230,N_7982,N_7632);
and U8231 (N_8231,N_7829,N_7760);
nand U8232 (N_8232,N_7788,N_7765);
xnor U8233 (N_8233,N_7843,N_7630);
nor U8234 (N_8234,N_7585,N_7874);
xor U8235 (N_8235,N_7867,N_7884);
nand U8236 (N_8236,N_7652,N_7972);
nand U8237 (N_8237,N_7790,N_7928);
or U8238 (N_8238,N_7910,N_7590);
nand U8239 (N_8239,N_7922,N_7643);
nor U8240 (N_8240,N_7609,N_7548);
nand U8241 (N_8241,N_7784,N_7556);
nand U8242 (N_8242,N_7900,N_7997);
and U8243 (N_8243,N_7840,N_7987);
and U8244 (N_8244,N_7511,N_7775);
xnor U8245 (N_8245,N_7601,N_7842);
xnor U8246 (N_8246,N_7962,N_7739);
and U8247 (N_8247,N_7886,N_7523);
or U8248 (N_8248,N_7709,N_7759);
nor U8249 (N_8249,N_7810,N_7578);
and U8250 (N_8250,N_7873,N_7988);
nand U8251 (N_8251,N_7832,N_7596);
and U8252 (N_8252,N_7954,N_7695);
nor U8253 (N_8253,N_7764,N_7849);
xor U8254 (N_8254,N_7808,N_7841);
or U8255 (N_8255,N_7782,N_7519);
nor U8256 (N_8256,N_7834,N_7761);
xor U8257 (N_8257,N_7537,N_7853);
or U8258 (N_8258,N_7624,N_7515);
or U8259 (N_8259,N_7833,N_7870);
or U8260 (N_8260,N_7978,N_7530);
or U8261 (N_8261,N_7735,N_7738);
nand U8262 (N_8262,N_7948,N_7517);
nor U8263 (N_8263,N_7599,N_7951);
or U8264 (N_8264,N_7652,N_7716);
nor U8265 (N_8265,N_7546,N_7674);
or U8266 (N_8266,N_7923,N_7742);
nand U8267 (N_8267,N_7589,N_7938);
or U8268 (N_8268,N_7887,N_7751);
nand U8269 (N_8269,N_7623,N_7949);
or U8270 (N_8270,N_7674,N_7967);
xnor U8271 (N_8271,N_7868,N_7898);
xor U8272 (N_8272,N_7720,N_7941);
nand U8273 (N_8273,N_7849,N_7804);
nor U8274 (N_8274,N_7627,N_7840);
xnor U8275 (N_8275,N_7838,N_7611);
nor U8276 (N_8276,N_7946,N_7938);
or U8277 (N_8277,N_7542,N_7787);
nand U8278 (N_8278,N_7588,N_7536);
nor U8279 (N_8279,N_7990,N_7854);
and U8280 (N_8280,N_7870,N_7505);
and U8281 (N_8281,N_7549,N_7867);
nand U8282 (N_8282,N_7694,N_7875);
nor U8283 (N_8283,N_7567,N_7804);
nand U8284 (N_8284,N_7951,N_7593);
nor U8285 (N_8285,N_7848,N_7843);
nand U8286 (N_8286,N_7934,N_7799);
and U8287 (N_8287,N_7981,N_7738);
nor U8288 (N_8288,N_7933,N_7507);
nand U8289 (N_8289,N_7504,N_7500);
and U8290 (N_8290,N_7853,N_7596);
nor U8291 (N_8291,N_7609,N_7668);
nand U8292 (N_8292,N_7824,N_7777);
and U8293 (N_8293,N_7544,N_7714);
and U8294 (N_8294,N_7972,N_7813);
or U8295 (N_8295,N_7657,N_7634);
xor U8296 (N_8296,N_7760,N_7948);
and U8297 (N_8297,N_7772,N_7534);
nand U8298 (N_8298,N_7562,N_7904);
nand U8299 (N_8299,N_7615,N_7513);
and U8300 (N_8300,N_7703,N_7612);
and U8301 (N_8301,N_7867,N_7605);
nor U8302 (N_8302,N_7540,N_7818);
or U8303 (N_8303,N_7976,N_7928);
xnor U8304 (N_8304,N_7994,N_7922);
and U8305 (N_8305,N_7543,N_7943);
xnor U8306 (N_8306,N_7810,N_7889);
nor U8307 (N_8307,N_7835,N_7662);
or U8308 (N_8308,N_7648,N_7617);
and U8309 (N_8309,N_7693,N_7843);
nand U8310 (N_8310,N_7675,N_7994);
and U8311 (N_8311,N_7929,N_7791);
nand U8312 (N_8312,N_7726,N_7827);
or U8313 (N_8313,N_7703,N_7993);
and U8314 (N_8314,N_7758,N_7616);
nor U8315 (N_8315,N_7557,N_7848);
xnor U8316 (N_8316,N_7698,N_7603);
and U8317 (N_8317,N_7664,N_7817);
xnor U8318 (N_8318,N_7691,N_7538);
nand U8319 (N_8319,N_7989,N_7531);
nor U8320 (N_8320,N_7691,N_7618);
nand U8321 (N_8321,N_7554,N_7852);
nand U8322 (N_8322,N_7669,N_7784);
xor U8323 (N_8323,N_7640,N_7968);
xor U8324 (N_8324,N_7787,N_7633);
xor U8325 (N_8325,N_7797,N_7717);
nor U8326 (N_8326,N_7834,N_7714);
nand U8327 (N_8327,N_7896,N_7701);
or U8328 (N_8328,N_7956,N_7837);
nor U8329 (N_8329,N_7542,N_7634);
xnor U8330 (N_8330,N_7711,N_7926);
nand U8331 (N_8331,N_7582,N_7817);
or U8332 (N_8332,N_7723,N_7591);
nor U8333 (N_8333,N_7815,N_7566);
xor U8334 (N_8334,N_7679,N_7876);
nor U8335 (N_8335,N_7838,N_7919);
and U8336 (N_8336,N_7555,N_7627);
xor U8337 (N_8337,N_7932,N_7855);
or U8338 (N_8338,N_7960,N_7575);
xor U8339 (N_8339,N_7592,N_7661);
xor U8340 (N_8340,N_7730,N_7757);
nor U8341 (N_8341,N_7646,N_7577);
and U8342 (N_8342,N_7853,N_7561);
nand U8343 (N_8343,N_7959,N_7743);
xor U8344 (N_8344,N_7979,N_7659);
xor U8345 (N_8345,N_7693,N_7797);
and U8346 (N_8346,N_7705,N_7762);
nand U8347 (N_8347,N_7742,N_7707);
nand U8348 (N_8348,N_7553,N_7639);
or U8349 (N_8349,N_7966,N_7869);
or U8350 (N_8350,N_7784,N_7874);
xor U8351 (N_8351,N_7838,N_7797);
nand U8352 (N_8352,N_7718,N_7635);
nand U8353 (N_8353,N_7891,N_7852);
or U8354 (N_8354,N_7723,N_7511);
or U8355 (N_8355,N_7614,N_7824);
nor U8356 (N_8356,N_7753,N_7764);
nor U8357 (N_8357,N_7613,N_7548);
and U8358 (N_8358,N_7681,N_7710);
nor U8359 (N_8359,N_7603,N_7686);
and U8360 (N_8360,N_7775,N_7555);
xor U8361 (N_8361,N_7706,N_7850);
and U8362 (N_8362,N_7957,N_7980);
xor U8363 (N_8363,N_7955,N_7531);
or U8364 (N_8364,N_7636,N_7684);
nand U8365 (N_8365,N_7970,N_7523);
xnor U8366 (N_8366,N_7792,N_7988);
nor U8367 (N_8367,N_7597,N_7832);
xor U8368 (N_8368,N_7891,N_7596);
and U8369 (N_8369,N_7738,N_7691);
or U8370 (N_8370,N_7541,N_7996);
or U8371 (N_8371,N_7710,N_7848);
or U8372 (N_8372,N_7603,N_7567);
and U8373 (N_8373,N_7902,N_7755);
nand U8374 (N_8374,N_7606,N_7538);
and U8375 (N_8375,N_7624,N_7748);
or U8376 (N_8376,N_7536,N_7761);
nand U8377 (N_8377,N_7744,N_7813);
or U8378 (N_8378,N_7703,N_7978);
or U8379 (N_8379,N_7686,N_7849);
nor U8380 (N_8380,N_7696,N_7664);
or U8381 (N_8381,N_7510,N_7678);
xor U8382 (N_8382,N_7787,N_7928);
and U8383 (N_8383,N_7724,N_7555);
xnor U8384 (N_8384,N_7916,N_7774);
nor U8385 (N_8385,N_7534,N_7714);
nor U8386 (N_8386,N_7926,N_7957);
or U8387 (N_8387,N_7856,N_7748);
and U8388 (N_8388,N_7944,N_7908);
or U8389 (N_8389,N_7827,N_7615);
or U8390 (N_8390,N_7519,N_7542);
or U8391 (N_8391,N_7633,N_7590);
and U8392 (N_8392,N_7691,N_7684);
nand U8393 (N_8393,N_7707,N_7692);
and U8394 (N_8394,N_7561,N_7918);
nand U8395 (N_8395,N_7915,N_7925);
nand U8396 (N_8396,N_7697,N_7800);
xor U8397 (N_8397,N_7627,N_7611);
nor U8398 (N_8398,N_7522,N_7946);
or U8399 (N_8399,N_7964,N_7657);
nor U8400 (N_8400,N_7716,N_7827);
nor U8401 (N_8401,N_7933,N_7894);
and U8402 (N_8402,N_7818,N_7503);
nor U8403 (N_8403,N_7832,N_7757);
or U8404 (N_8404,N_7740,N_7941);
and U8405 (N_8405,N_7884,N_7782);
and U8406 (N_8406,N_7535,N_7835);
xnor U8407 (N_8407,N_7978,N_7901);
xor U8408 (N_8408,N_7975,N_7633);
nand U8409 (N_8409,N_7534,N_7823);
nand U8410 (N_8410,N_7987,N_7854);
or U8411 (N_8411,N_7758,N_7767);
nand U8412 (N_8412,N_7522,N_7910);
nor U8413 (N_8413,N_7836,N_7976);
xnor U8414 (N_8414,N_7636,N_7946);
xnor U8415 (N_8415,N_7987,N_7828);
and U8416 (N_8416,N_7668,N_7724);
and U8417 (N_8417,N_7891,N_7770);
nand U8418 (N_8418,N_7623,N_7761);
or U8419 (N_8419,N_7902,N_7927);
xor U8420 (N_8420,N_7671,N_7766);
or U8421 (N_8421,N_7628,N_7568);
or U8422 (N_8422,N_7541,N_7935);
nor U8423 (N_8423,N_7604,N_7766);
and U8424 (N_8424,N_7702,N_7984);
xor U8425 (N_8425,N_7599,N_7638);
nand U8426 (N_8426,N_7601,N_7608);
nor U8427 (N_8427,N_7644,N_7526);
xnor U8428 (N_8428,N_7702,N_7540);
or U8429 (N_8429,N_7849,N_7562);
xnor U8430 (N_8430,N_7549,N_7508);
or U8431 (N_8431,N_7851,N_7615);
and U8432 (N_8432,N_7834,N_7769);
or U8433 (N_8433,N_7775,N_7961);
and U8434 (N_8434,N_7597,N_7741);
nor U8435 (N_8435,N_7728,N_7875);
or U8436 (N_8436,N_7758,N_7645);
and U8437 (N_8437,N_7983,N_7813);
nand U8438 (N_8438,N_7585,N_7588);
nand U8439 (N_8439,N_7721,N_7729);
or U8440 (N_8440,N_7908,N_7636);
nand U8441 (N_8441,N_7760,N_7816);
xor U8442 (N_8442,N_7765,N_7795);
nor U8443 (N_8443,N_7694,N_7712);
and U8444 (N_8444,N_7601,N_7801);
and U8445 (N_8445,N_7995,N_7702);
or U8446 (N_8446,N_7858,N_7966);
and U8447 (N_8447,N_7967,N_7902);
nand U8448 (N_8448,N_7597,N_7717);
or U8449 (N_8449,N_7563,N_7885);
or U8450 (N_8450,N_7993,N_7811);
xnor U8451 (N_8451,N_7500,N_7581);
nand U8452 (N_8452,N_7991,N_7691);
or U8453 (N_8453,N_7843,N_7589);
and U8454 (N_8454,N_7672,N_7557);
nand U8455 (N_8455,N_7771,N_7801);
or U8456 (N_8456,N_7569,N_7905);
nor U8457 (N_8457,N_7512,N_7978);
or U8458 (N_8458,N_7691,N_7900);
or U8459 (N_8459,N_7853,N_7567);
and U8460 (N_8460,N_7845,N_7662);
and U8461 (N_8461,N_7900,N_7860);
nand U8462 (N_8462,N_7749,N_7968);
nor U8463 (N_8463,N_7938,N_7621);
xnor U8464 (N_8464,N_7670,N_7825);
or U8465 (N_8465,N_7853,N_7916);
and U8466 (N_8466,N_7909,N_7697);
xor U8467 (N_8467,N_7983,N_7569);
xnor U8468 (N_8468,N_7537,N_7810);
and U8469 (N_8469,N_7590,N_7679);
or U8470 (N_8470,N_7661,N_7923);
and U8471 (N_8471,N_7797,N_7922);
nand U8472 (N_8472,N_7712,N_7865);
nand U8473 (N_8473,N_7998,N_7941);
nor U8474 (N_8474,N_7845,N_7935);
and U8475 (N_8475,N_7737,N_7641);
or U8476 (N_8476,N_7667,N_7755);
or U8477 (N_8477,N_7691,N_7931);
or U8478 (N_8478,N_7787,N_7625);
nor U8479 (N_8479,N_7957,N_7634);
or U8480 (N_8480,N_7750,N_7847);
or U8481 (N_8481,N_7862,N_7995);
nand U8482 (N_8482,N_7963,N_7751);
nand U8483 (N_8483,N_7967,N_7546);
or U8484 (N_8484,N_7803,N_7537);
and U8485 (N_8485,N_7983,N_7545);
and U8486 (N_8486,N_7654,N_7681);
or U8487 (N_8487,N_7519,N_7787);
nand U8488 (N_8488,N_7500,N_7982);
and U8489 (N_8489,N_7757,N_7580);
nor U8490 (N_8490,N_7786,N_7501);
xnor U8491 (N_8491,N_7826,N_7703);
nor U8492 (N_8492,N_7943,N_7973);
xor U8493 (N_8493,N_7856,N_7709);
xor U8494 (N_8494,N_7689,N_7590);
or U8495 (N_8495,N_7703,N_7902);
xnor U8496 (N_8496,N_7533,N_7694);
xor U8497 (N_8497,N_7736,N_7682);
and U8498 (N_8498,N_7512,N_7513);
or U8499 (N_8499,N_7747,N_7569);
xor U8500 (N_8500,N_8324,N_8301);
or U8501 (N_8501,N_8236,N_8174);
nand U8502 (N_8502,N_8012,N_8279);
and U8503 (N_8503,N_8345,N_8285);
xor U8504 (N_8504,N_8258,N_8460);
nand U8505 (N_8505,N_8342,N_8153);
and U8506 (N_8506,N_8384,N_8106);
nor U8507 (N_8507,N_8134,N_8125);
nor U8508 (N_8508,N_8095,N_8377);
nand U8509 (N_8509,N_8178,N_8351);
nand U8510 (N_8510,N_8235,N_8437);
nor U8511 (N_8511,N_8193,N_8272);
nand U8512 (N_8512,N_8195,N_8312);
and U8513 (N_8513,N_8109,N_8024);
xnor U8514 (N_8514,N_8292,N_8217);
or U8515 (N_8515,N_8197,N_8485);
nor U8516 (N_8516,N_8154,N_8383);
or U8517 (N_8517,N_8090,N_8323);
and U8518 (N_8518,N_8439,N_8287);
xor U8519 (N_8519,N_8492,N_8418);
or U8520 (N_8520,N_8348,N_8189);
nor U8521 (N_8521,N_8476,N_8468);
xor U8522 (N_8522,N_8014,N_8206);
nor U8523 (N_8523,N_8071,N_8433);
nand U8524 (N_8524,N_8310,N_8443);
nor U8525 (N_8525,N_8023,N_8117);
nand U8526 (N_8526,N_8202,N_8188);
or U8527 (N_8527,N_8094,N_8474);
nor U8528 (N_8528,N_8123,N_8388);
xor U8529 (N_8529,N_8159,N_8131);
or U8530 (N_8530,N_8009,N_8083);
and U8531 (N_8531,N_8403,N_8151);
and U8532 (N_8532,N_8479,N_8074);
xor U8533 (N_8533,N_8302,N_8232);
nor U8534 (N_8534,N_8214,N_8179);
xor U8535 (N_8535,N_8166,N_8004);
nor U8536 (N_8536,N_8011,N_8340);
and U8537 (N_8537,N_8170,N_8026);
xor U8538 (N_8538,N_8239,N_8390);
nor U8539 (N_8539,N_8252,N_8102);
nor U8540 (N_8540,N_8201,N_8008);
nor U8541 (N_8541,N_8475,N_8380);
and U8542 (N_8542,N_8070,N_8286);
nand U8543 (N_8543,N_8404,N_8129);
nor U8544 (N_8544,N_8163,N_8311);
nand U8545 (N_8545,N_8213,N_8007);
nand U8546 (N_8546,N_8414,N_8341);
xor U8547 (N_8547,N_8181,N_8168);
or U8548 (N_8548,N_8415,N_8013);
and U8549 (N_8549,N_8167,N_8079);
nor U8550 (N_8550,N_8470,N_8190);
or U8551 (N_8551,N_8049,N_8489);
nor U8552 (N_8552,N_8427,N_8169);
and U8553 (N_8553,N_8097,N_8028);
xor U8554 (N_8554,N_8056,N_8277);
nand U8555 (N_8555,N_8077,N_8382);
or U8556 (N_8556,N_8454,N_8171);
nor U8557 (N_8557,N_8314,N_8005);
nor U8558 (N_8558,N_8486,N_8135);
or U8559 (N_8559,N_8051,N_8156);
or U8560 (N_8560,N_8172,N_8091);
and U8561 (N_8561,N_8127,N_8021);
and U8562 (N_8562,N_8379,N_8267);
nand U8563 (N_8563,N_8347,N_8034);
xnor U8564 (N_8564,N_8205,N_8303);
or U8565 (N_8565,N_8290,N_8173);
nor U8566 (N_8566,N_8350,N_8374);
or U8567 (N_8567,N_8257,N_8065);
nand U8568 (N_8568,N_8096,N_8488);
nand U8569 (N_8569,N_8221,N_8280);
xnor U8570 (N_8570,N_8422,N_8062);
nor U8571 (N_8571,N_8376,N_8082);
nor U8572 (N_8572,N_8420,N_8080);
and U8573 (N_8573,N_8448,N_8480);
or U8574 (N_8574,N_8118,N_8491);
nand U8575 (N_8575,N_8183,N_8053);
and U8576 (N_8576,N_8473,N_8396);
and U8577 (N_8577,N_8104,N_8234);
nand U8578 (N_8578,N_8325,N_8025);
xnor U8579 (N_8579,N_8140,N_8275);
nor U8580 (N_8580,N_8144,N_8224);
nand U8581 (N_8581,N_8229,N_8246);
or U8582 (N_8582,N_8299,N_8136);
xnor U8583 (N_8583,N_8157,N_8278);
nor U8584 (N_8584,N_8318,N_8450);
nand U8585 (N_8585,N_8200,N_8084);
nand U8586 (N_8586,N_8438,N_8274);
xor U8587 (N_8587,N_8499,N_8288);
nand U8588 (N_8588,N_8133,N_8255);
and U8589 (N_8589,N_8464,N_8164);
nor U8590 (N_8590,N_8319,N_8497);
and U8591 (N_8591,N_8000,N_8216);
xor U8592 (N_8592,N_8250,N_8260);
nand U8593 (N_8593,N_8078,N_8329);
xnor U8594 (N_8594,N_8461,N_8268);
xor U8595 (N_8595,N_8101,N_8281);
nand U8596 (N_8596,N_8247,N_8478);
and U8597 (N_8597,N_8098,N_8225);
or U8598 (N_8598,N_8191,N_8110);
nand U8599 (N_8599,N_8442,N_8316);
xnor U8600 (N_8600,N_8322,N_8240);
nand U8601 (N_8601,N_8033,N_8463);
and U8602 (N_8602,N_8068,N_8370);
nor U8603 (N_8603,N_8054,N_8243);
xor U8604 (N_8604,N_8208,N_8389);
nor U8605 (N_8605,N_8297,N_8435);
nand U8606 (N_8606,N_8270,N_8063);
nand U8607 (N_8607,N_8482,N_8293);
or U8608 (N_8608,N_8385,N_8425);
nand U8609 (N_8609,N_8148,N_8483);
xor U8610 (N_8610,N_8320,N_8241);
nor U8611 (N_8611,N_8269,N_8006);
and U8612 (N_8612,N_8371,N_8199);
nand U8613 (N_8613,N_8328,N_8251);
xor U8614 (N_8614,N_8198,N_8146);
nor U8615 (N_8615,N_8089,N_8030);
and U8616 (N_8616,N_8405,N_8399);
nor U8617 (N_8617,N_8002,N_8059);
and U8618 (N_8618,N_8362,N_8037);
or U8619 (N_8619,N_8363,N_8245);
or U8620 (N_8620,N_8132,N_8203);
nor U8621 (N_8621,N_8185,N_8387);
nand U8622 (N_8622,N_8233,N_8067);
and U8623 (N_8623,N_8400,N_8349);
and U8624 (N_8624,N_8044,N_8394);
and U8625 (N_8625,N_8061,N_8262);
and U8626 (N_8626,N_8451,N_8050);
nand U8627 (N_8627,N_8308,N_8165);
and U8628 (N_8628,N_8452,N_8326);
xor U8629 (N_8629,N_8048,N_8402);
nand U8630 (N_8630,N_8375,N_8114);
and U8631 (N_8631,N_8466,N_8259);
xor U8632 (N_8632,N_8103,N_8226);
and U8633 (N_8633,N_8364,N_8411);
and U8634 (N_8634,N_8313,N_8088);
xnor U8635 (N_8635,N_8130,N_8343);
nand U8636 (N_8636,N_8219,N_8256);
or U8637 (N_8637,N_8058,N_8423);
or U8638 (N_8638,N_8458,N_8176);
nand U8639 (N_8639,N_8001,N_8043);
or U8640 (N_8640,N_8042,N_8115);
nand U8641 (N_8641,N_8421,N_8227);
xor U8642 (N_8642,N_8352,N_8365);
nand U8643 (N_8643,N_8398,N_8177);
nor U8644 (N_8644,N_8338,N_8212);
nand U8645 (N_8645,N_8253,N_8413);
nand U8646 (N_8646,N_8498,N_8108);
or U8647 (N_8647,N_8107,N_8361);
xnor U8648 (N_8648,N_8472,N_8186);
xor U8649 (N_8649,N_8180,N_8099);
nand U8650 (N_8650,N_8052,N_8471);
nor U8651 (N_8651,N_8294,N_8495);
and U8652 (N_8652,N_8357,N_8066);
and U8653 (N_8653,N_8228,N_8330);
or U8654 (N_8654,N_8069,N_8391);
and U8655 (N_8655,N_8242,N_8223);
nand U8656 (N_8656,N_8073,N_8018);
and U8657 (N_8657,N_8032,N_8453);
and U8658 (N_8658,N_8113,N_8010);
nand U8659 (N_8659,N_8428,N_8211);
and U8660 (N_8660,N_8417,N_8017);
or U8661 (N_8661,N_8112,N_8477);
xnor U8662 (N_8662,N_8149,N_8358);
xor U8663 (N_8663,N_8353,N_8335);
or U8664 (N_8664,N_8003,N_8244);
and U8665 (N_8665,N_8386,N_8120);
nor U8666 (N_8666,N_8344,N_8332);
xor U8667 (N_8667,N_8138,N_8465);
nand U8668 (N_8668,N_8055,N_8087);
xnor U8669 (N_8669,N_8487,N_8126);
nand U8670 (N_8670,N_8484,N_8029);
nand U8671 (N_8671,N_8462,N_8248);
nor U8672 (N_8672,N_8305,N_8038);
nor U8673 (N_8673,N_8237,N_8295);
nand U8674 (N_8674,N_8230,N_8254);
and U8675 (N_8675,N_8076,N_8218);
xnor U8676 (N_8676,N_8020,N_8416);
nor U8677 (N_8677,N_8204,N_8446);
nor U8678 (N_8678,N_8457,N_8222);
or U8679 (N_8679,N_8031,N_8467);
nor U8680 (N_8680,N_8441,N_8022);
or U8681 (N_8681,N_8147,N_8336);
and U8682 (N_8682,N_8496,N_8047);
or U8683 (N_8683,N_8092,N_8161);
xor U8684 (N_8684,N_8081,N_8354);
nor U8685 (N_8685,N_8265,N_8284);
or U8686 (N_8686,N_8321,N_8261);
and U8687 (N_8687,N_8209,N_8162);
and U8688 (N_8688,N_8333,N_8494);
nand U8689 (N_8689,N_8152,N_8298);
nand U8690 (N_8690,N_8412,N_8045);
xor U8691 (N_8691,N_8215,N_8128);
xor U8692 (N_8692,N_8016,N_8440);
and U8693 (N_8693,N_8447,N_8137);
nand U8694 (N_8694,N_8306,N_8493);
or U8695 (N_8695,N_8184,N_8327);
and U8696 (N_8696,N_8220,N_8369);
and U8697 (N_8697,N_8431,N_8368);
nand U8698 (N_8698,N_8426,N_8158);
nor U8699 (N_8699,N_8139,N_8296);
and U8700 (N_8700,N_8100,N_8490);
nor U8701 (N_8701,N_8035,N_8249);
and U8702 (N_8702,N_8116,N_8445);
or U8703 (N_8703,N_8397,N_8432);
and U8704 (N_8704,N_8355,N_8430);
and U8705 (N_8705,N_8367,N_8105);
nand U8706 (N_8706,N_8283,N_8392);
and U8707 (N_8707,N_8060,N_8150);
nand U8708 (N_8708,N_8291,N_8409);
or U8709 (N_8709,N_8019,N_8309);
nand U8710 (N_8710,N_8429,N_8040);
or U8711 (N_8711,N_8406,N_8373);
xnor U8712 (N_8712,N_8273,N_8111);
and U8713 (N_8713,N_8238,N_8444);
xor U8714 (N_8714,N_8036,N_8145);
or U8715 (N_8715,N_8155,N_8393);
nand U8716 (N_8716,N_8160,N_8317);
nand U8717 (N_8717,N_8331,N_8192);
xor U8718 (N_8718,N_8378,N_8271);
nand U8719 (N_8719,N_8057,N_8041);
xnor U8720 (N_8720,N_8395,N_8264);
nor U8721 (N_8721,N_8266,N_8424);
nand U8722 (N_8722,N_8182,N_8086);
or U8723 (N_8723,N_8359,N_8210);
and U8724 (N_8724,N_8456,N_8276);
and U8725 (N_8725,N_8124,N_8315);
xor U8726 (N_8726,N_8436,N_8410);
nand U8727 (N_8727,N_8372,N_8039);
and U8728 (N_8728,N_8346,N_8141);
or U8729 (N_8729,N_8187,N_8282);
or U8730 (N_8730,N_8434,N_8339);
or U8731 (N_8731,N_8263,N_8356);
nand U8732 (N_8732,N_8027,N_8459);
nand U8733 (N_8733,N_8143,N_8366);
and U8734 (N_8734,N_8064,N_8072);
nand U8735 (N_8735,N_8455,N_8142);
and U8736 (N_8736,N_8304,N_8046);
or U8737 (N_8737,N_8231,N_8360);
nand U8738 (N_8738,N_8085,N_8015);
nand U8739 (N_8739,N_8408,N_8481);
nand U8740 (N_8740,N_8196,N_8093);
and U8741 (N_8741,N_8419,N_8381);
nand U8742 (N_8742,N_8307,N_8300);
and U8743 (N_8743,N_8289,N_8401);
nor U8744 (N_8744,N_8207,N_8119);
and U8745 (N_8745,N_8194,N_8122);
nor U8746 (N_8746,N_8075,N_8337);
nor U8747 (N_8747,N_8449,N_8407);
nor U8748 (N_8748,N_8334,N_8469);
or U8749 (N_8749,N_8121,N_8175);
nor U8750 (N_8750,N_8294,N_8189);
nand U8751 (N_8751,N_8217,N_8427);
or U8752 (N_8752,N_8049,N_8174);
nor U8753 (N_8753,N_8451,N_8171);
and U8754 (N_8754,N_8489,N_8444);
nand U8755 (N_8755,N_8486,N_8179);
and U8756 (N_8756,N_8220,N_8113);
nor U8757 (N_8757,N_8111,N_8145);
xnor U8758 (N_8758,N_8375,N_8178);
or U8759 (N_8759,N_8265,N_8015);
and U8760 (N_8760,N_8169,N_8395);
and U8761 (N_8761,N_8285,N_8042);
nand U8762 (N_8762,N_8194,N_8429);
and U8763 (N_8763,N_8010,N_8486);
xnor U8764 (N_8764,N_8019,N_8073);
nand U8765 (N_8765,N_8271,N_8021);
or U8766 (N_8766,N_8426,N_8329);
nand U8767 (N_8767,N_8037,N_8050);
nor U8768 (N_8768,N_8137,N_8485);
nand U8769 (N_8769,N_8450,N_8209);
and U8770 (N_8770,N_8005,N_8299);
and U8771 (N_8771,N_8089,N_8484);
nand U8772 (N_8772,N_8041,N_8166);
nand U8773 (N_8773,N_8051,N_8116);
nand U8774 (N_8774,N_8320,N_8174);
nand U8775 (N_8775,N_8075,N_8054);
and U8776 (N_8776,N_8009,N_8020);
nand U8777 (N_8777,N_8148,N_8105);
xnor U8778 (N_8778,N_8351,N_8079);
nor U8779 (N_8779,N_8216,N_8254);
and U8780 (N_8780,N_8232,N_8409);
nand U8781 (N_8781,N_8049,N_8041);
nand U8782 (N_8782,N_8047,N_8229);
and U8783 (N_8783,N_8016,N_8408);
and U8784 (N_8784,N_8152,N_8424);
and U8785 (N_8785,N_8122,N_8178);
or U8786 (N_8786,N_8288,N_8404);
nand U8787 (N_8787,N_8066,N_8219);
and U8788 (N_8788,N_8443,N_8438);
or U8789 (N_8789,N_8295,N_8452);
nor U8790 (N_8790,N_8010,N_8222);
and U8791 (N_8791,N_8022,N_8195);
nor U8792 (N_8792,N_8408,N_8300);
xnor U8793 (N_8793,N_8058,N_8314);
xor U8794 (N_8794,N_8228,N_8043);
nand U8795 (N_8795,N_8397,N_8424);
nor U8796 (N_8796,N_8367,N_8089);
and U8797 (N_8797,N_8408,N_8332);
nand U8798 (N_8798,N_8321,N_8179);
xnor U8799 (N_8799,N_8423,N_8340);
xnor U8800 (N_8800,N_8372,N_8471);
or U8801 (N_8801,N_8047,N_8089);
nand U8802 (N_8802,N_8411,N_8256);
and U8803 (N_8803,N_8344,N_8307);
nand U8804 (N_8804,N_8080,N_8275);
and U8805 (N_8805,N_8495,N_8321);
xnor U8806 (N_8806,N_8086,N_8110);
nand U8807 (N_8807,N_8188,N_8026);
or U8808 (N_8808,N_8088,N_8101);
nand U8809 (N_8809,N_8254,N_8460);
and U8810 (N_8810,N_8439,N_8000);
xnor U8811 (N_8811,N_8137,N_8153);
nor U8812 (N_8812,N_8182,N_8489);
nor U8813 (N_8813,N_8223,N_8481);
xor U8814 (N_8814,N_8287,N_8001);
or U8815 (N_8815,N_8310,N_8202);
nand U8816 (N_8816,N_8092,N_8188);
nor U8817 (N_8817,N_8325,N_8349);
or U8818 (N_8818,N_8495,N_8476);
nor U8819 (N_8819,N_8339,N_8134);
nor U8820 (N_8820,N_8115,N_8472);
or U8821 (N_8821,N_8254,N_8210);
and U8822 (N_8822,N_8461,N_8216);
and U8823 (N_8823,N_8084,N_8428);
nor U8824 (N_8824,N_8247,N_8089);
nor U8825 (N_8825,N_8313,N_8429);
xor U8826 (N_8826,N_8027,N_8207);
or U8827 (N_8827,N_8372,N_8434);
or U8828 (N_8828,N_8191,N_8044);
and U8829 (N_8829,N_8137,N_8460);
or U8830 (N_8830,N_8010,N_8327);
nor U8831 (N_8831,N_8024,N_8194);
xnor U8832 (N_8832,N_8076,N_8210);
nor U8833 (N_8833,N_8407,N_8413);
and U8834 (N_8834,N_8172,N_8243);
nand U8835 (N_8835,N_8039,N_8209);
or U8836 (N_8836,N_8257,N_8125);
nor U8837 (N_8837,N_8262,N_8442);
nor U8838 (N_8838,N_8367,N_8019);
nor U8839 (N_8839,N_8203,N_8421);
and U8840 (N_8840,N_8033,N_8413);
nor U8841 (N_8841,N_8137,N_8173);
xnor U8842 (N_8842,N_8292,N_8321);
xor U8843 (N_8843,N_8102,N_8448);
xor U8844 (N_8844,N_8294,N_8066);
or U8845 (N_8845,N_8171,N_8059);
and U8846 (N_8846,N_8313,N_8004);
and U8847 (N_8847,N_8012,N_8310);
nor U8848 (N_8848,N_8326,N_8094);
nand U8849 (N_8849,N_8434,N_8165);
and U8850 (N_8850,N_8467,N_8096);
and U8851 (N_8851,N_8172,N_8388);
or U8852 (N_8852,N_8442,N_8015);
and U8853 (N_8853,N_8303,N_8063);
nor U8854 (N_8854,N_8143,N_8093);
nand U8855 (N_8855,N_8300,N_8475);
and U8856 (N_8856,N_8009,N_8452);
nor U8857 (N_8857,N_8423,N_8372);
and U8858 (N_8858,N_8036,N_8004);
and U8859 (N_8859,N_8406,N_8024);
and U8860 (N_8860,N_8072,N_8494);
or U8861 (N_8861,N_8219,N_8490);
nand U8862 (N_8862,N_8251,N_8026);
or U8863 (N_8863,N_8108,N_8167);
or U8864 (N_8864,N_8311,N_8062);
nor U8865 (N_8865,N_8435,N_8148);
and U8866 (N_8866,N_8061,N_8056);
nor U8867 (N_8867,N_8090,N_8327);
nor U8868 (N_8868,N_8030,N_8402);
and U8869 (N_8869,N_8064,N_8214);
nor U8870 (N_8870,N_8460,N_8417);
nor U8871 (N_8871,N_8026,N_8444);
nor U8872 (N_8872,N_8247,N_8192);
nand U8873 (N_8873,N_8347,N_8184);
xor U8874 (N_8874,N_8487,N_8390);
and U8875 (N_8875,N_8000,N_8153);
or U8876 (N_8876,N_8383,N_8147);
or U8877 (N_8877,N_8497,N_8376);
xor U8878 (N_8878,N_8286,N_8366);
xor U8879 (N_8879,N_8238,N_8162);
or U8880 (N_8880,N_8157,N_8131);
xor U8881 (N_8881,N_8144,N_8154);
and U8882 (N_8882,N_8034,N_8171);
nand U8883 (N_8883,N_8071,N_8498);
or U8884 (N_8884,N_8122,N_8464);
and U8885 (N_8885,N_8403,N_8051);
nor U8886 (N_8886,N_8378,N_8344);
nor U8887 (N_8887,N_8257,N_8364);
nand U8888 (N_8888,N_8046,N_8082);
and U8889 (N_8889,N_8223,N_8391);
nand U8890 (N_8890,N_8272,N_8144);
nand U8891 (N_8891,N_8094,N_8050);
xnor U8892 (N_8892,N_8438,N_8308);
nand U8893 (N_8893,N_8219,N_8307);
nor U8894 (N_8894,N_8193,N_8381);
xnor U8895 (N_8895,N_8258,N_8250);
or U8896 (N_8896,N_8365,N_8466);
xnor U8897 (N_8897,N_8245,N_8114);
nor U8898 (N_8898,N_8431,N_8009);
and U8899 (N_8899,N_8023,N_8209);
xor U8900 (N_8900,N_8015,N_8436);
xnor U8901 (N_8901,N_8431,N_8132);
or U8902 (N_8902,N_8375,N_8478);
xnor U8903 (N_8903,N_8332,N_8183);
or U8904 (N_8904,N_8256,N_8284);
nor U8905 (N_8905,N_8463,N_8468);
xor U8906 (N_8906,N_8287,N_8283);
xnor U8907 (N_8907,N_8132,N_8451);
xor U8908 (N_8908,N_8353,N_8111);
xnor U8909 (N_8909,N_8140,N_8395);
or U8910 (N_8910,N_8432,N_8112);
xor U8911 (N_8911,N_8262,N_8049);
or U8912 (N_8912,N_8112,N_8016);
and U8913 (N_8913,N_8481,N_8129);
or U8914 (N_8914,N_8074,N_8125);
nand U8915 (N_8915,N_8001,N_8088);
nand U8916 (N_8916,N_8083,N_8139);
nor U8917 (N_8917,N_8477,N_8102);
or U8918 (N_8918,N_8349,N_8357);
and U8919 (N_8919,N_8133,N_8377);
xnor U8920 (N_8920,N_8175,N_8265);
nand U8921 (N_8921,N_8462,N_8372);
and U8922 (N_8922,N_8358,N_8267);
nand U8923 (N_8923,N_8190,N_8244);
nand U8924 (N_8924,N_8006,N_8081);
and U8925 (N_8925,N_8371,N_8344);
nor U8926 (N_8926,N_8106,N_8242);
nor U8927 (N_8927,N_8312,N_8000);
nor U8928 (N_8928,N_8179,N_8204);
nand U8929 (N_8929,N_8026,N_8247);
nor U8930 (N_8930,N_8438,N_8404);
xor U8931 (N_8931,N_8047,N_8002);
xor U8932 (N_8932,N_8320,N_8494);
nand U8933 (N_8933,N_8123,N_8396);
xor U8934 (N_8934,N_8237,N_8349);
or U8935 (N_8935,N_8057,N_8441);
nand U8936 (N_8936,N_8043,N_8123);
xor U8937 (N_8937,N_8274,N_8305);
xnor U8938 (N_8938,N_8434,N_8026);
or U8939 (N_8939,N_8387,N_8294);
and U8940 (N_8940,N_8372,N_8337);
xor U8941 (N_8941,N_8025,N_8462);
xor U8942 (N_8942,N_8043,N_8476);
and U8943 (N_8943,N_8177,N_8418);
xor U8944 (N_8944,N_8461,N_8438);
nand U8945 (N_8945,N_8110,N_8088);
nor U8946 (N_8946,N_8331,N_8419);
nor U8947 (N_8947,N_8190,N_8387);
nor U8948 (N_8948,N_8410,N_8081);
nand U8949 (N_8949,N_8062,N_8263);
nand U8950 (N_8950,N_8051,N_8404);
nor U8951 (N_8951,N_8415,N_8396);
nor U8952 (N_8952,N_8169,N_8174);
xor U8953 (N_8953,N_8065,N_8078);
or U8954 (N_8954,N_8302,N_8155);
nor U8955 (N_8955,N_8058,N_8291);
nand U8956 (N_8956,N_8465,N_8121);
xnor U8957 (N_8957,N_8066,N_8245);
nor U8958 (N_8958,N_8233,N_8374);
and U8959 (N_8959,N_8002,N_8123);
nand U8960 (N_8960,N_8462,N_8345);
and U8961 (N_8961,N_8171,N_8249);
nor U8962 (N_8962,N_8290,N_8484);
nand U8963 (N_8963,N_8232,N_8074);
xnor U8964 (N_8964,N_8146,N_8057);
nand U8965 (N_8965,N_8356,N_8140);
and U8966 (N_8966,N_8273,N_8343);
and U8967 (N_8967,N_8370,N_8164);
and U8968 (N_8968,N_8107,N_8359);
xnor U8969 (N_8969,N_8374,N_8299);
and U8970 (N_8970,N_8190,N_8440);
xnor U8971 (N_8971,N_8123,N_8413);
or U8972 (N_8972,N_8036,N_8178);
nor U8973 (N_8973,N_8376,N_8170);
and U8974 (N_8974,N_8419,N_8002);
nor U8975 (N_8975,N_8160,N_8155);
and U8976 (N_8976,N_8013,N_8028);
and U8977 (N_8977,N_8338,N_8469);
nand U8978 (N_8978,N_8035,N_8340);
nor U8979 (N_8979,N_8493,N_8339);
nand U8980 (N_8980,N_8265,N_8463);
or U8981 (N_8981,N_8437,N_8362);
and U8982 (N_8982,N_8269,N_8479);
nand U8983 (N_8983,N_8020,N_8475);
or U8984 (N_8984,N_8490,N_8278);
xor U8985 (N_8985,N_8342,N_8045);
xnor U8986 (N_8986,N_8236,N_8197);
or U8987 (N_8987,N_8044,N_8251);
and U8988 (N_8988,N_8213,N_8065);
nor U8989 (N_8989,N_8468,N_8192);
xnor U8990 (N_8990,N_8267,N_8457);
xnor U8991 (N_8991,N_8249,N_8177);
and U8992 (N_8992,N_8365,N_8200);
and U8993 (N_8993,N_8454,N_8287);
nor U8994 (N_8994,N_8139,N_8396);
nand U8995 (N_8995,N_8188,N_8401);
and U8996 (N_8996,N_8441,N_8216);
xor U8997 (N_8997,N_8303,N_8074);
or U8998 (N_8998,N_8345,N_8230);
or U8999 (N_8999,N_8151,N_8134);
and U9000 (N_9000,N_8634,N_8838);
xnor U9001 (N_9001,N_8784,N_8641);
and U9002 (N_9002,N_8741,N_8608);
nand U9003 (N_9003,N_8789,N_8625);
and U9004 (N_9004,N_8756,N_8669);
or U9005 (N_9005,N_8824,N_8623);
or U9006 (N_9006,N_8512,N_8963);
and U9007 (N_9007,N_8762,N_8597);
xor U9008 (N_9008,N_8667,N_8939);
and U9009 (N_9009,N_8966,N_8653);
and U9010 (N_9010,N_8964,N_8632);
xor U9011 (N_9011,N_8660,N_8984);
and U9012 (N_9012,N_8593,N_8907);
and U9013 (N_9013,N_8734,N_8574);
xnor U9014 (N_9014,N_8813,N_8547);
xnor U9015 (N_9015,N_8771,N_8913);
or U9016 (N_9016,N_8884,N_8621);
and U9017 (N_9017,N_8742,N_8721);
nor U9018 (N_9018,N_8924,N_8639);
or U9019 (N_9019,N_8686,N_8816);
nand U9020 (N_9020,N_8754,N_8798);
nor U9021 (N_9021,N_8891,N_8647);
nand U9022 (N_9022,N_8659,N_8804);
nor U9023 (N_9023,N_8875,N_8548);
nand U9024 (N_9024,N_8949,N_8562);
nor U9025 (N_9025,N_8751,N_8604);
and U9026 (N_9026,N_8703,N_8753);
xor U9027 (N_9027,N_8672,N_8509);
nand U9028 (N_9028,N_8515,N_8823);
and U9029 (N_9029,N_8769,N_8976);
xnor U9030 (N_9030,N_8561,N_8550);
nand U9031 (N_9031,N_8673,N_8989);
xor U9032 (N_9032,N_8542,N_8802);
and U9033 (N_9033,N_8900,N_8882);
xnor U9034 (N_9034,N_8591,N_8782);
and U9035 (N_9035,N_8956,N_8527);
nand U9036 (N_9036,N_8567,N_8654);
nand U9037 (N_9037,N_8849,N_8968);
nor U9038 (N_9038,N_8776,N_8658);
or U9039 (N_9039,N_8503,N_8555);
and U9040 (N_9040,N_8827,N_8755);
xor U9041 (N_9041,N_8998,N_8601);
nand U9042 (N_9042,N_8916,N_8705);
nor U9043 (N_9043,N_8965,N_8874);
nor U9044 (N_9044,N_8517,N_8828);
xor U9045 (N_9045,N_8731,N_8644);
and U9046 (N_9046,N_8841,N_8817);
or U9047 (N_9047,N_8911,N_8952);
or U9048 (N_9048,N_8925,N_8545);
nor U9049 (N_9049,N_8991,N_8699);
nand U9050 (N_9050,N_8788,N_8738);
xor U9051 (N_9051,N_8941,N_8612);
and U9052 (N_9052,N_8812,N_8611);
xor U9053 (N_9053,N_8583,N_8851);
or U9054 (N_9054,N_8622,N_8847);
nor U9055 (N_9055,N_8945,N_8981);
and U9056 (N_9056,N_8957,N_8848);
xor U9057 (N_9057,N_8843,N_8662);
nand U9058 (N_9058,N_8711,N_8930);
nor U9059 (N_9059,N_8932,N_8779);
nor U9060 (N_9060,N_8839,N_8682);
xnor U9061 (N_9061,N_8960,N_8858);
nand U9062 (N_9062,N_8893,N_8767);
xnor U9063 (N_9063,N_8842,N_8533);
xnor U9064 (N_9064,N_8571,N_8556);
or U9065 (N_9065,N_8748,N_8657);
and U9066 (N_9066,N_8743,N_8563);
xnor U9067 (N_9067,N_8852,N_8580);
nor U9068 (N_9068,N_8931,N_8894);
nor U9069 (N_9069,N_8559,N_8954);
nor U9070 (N_9070,N_8709,N_8724);
and U9071 (N_9071,N_8665,N_8857);
xnor U9072 (N_9072,N_8922,N_8640);
and U9073 (N_9073,N_8810,N_8959);
and U9074 (N_9074,N_8727,N_8706);
nor U9075 (N_9075,N_8615,N_8821);
nor U9076 (N_9076,N_8543,N_8978);
or U9077 (N_9077,N_8683,N_8720);
nor U9078 (N_9078,N_8850,N_8607);
or U9079 (N_9079,N_8783,N_8750);
xor U9080 (N_9080,N_8935,N_8766);
and U9081 (N_9081,N_8862,N_8938);
nand U9082 (N_9082,N_8970,N_8871);
or U9083 (N_9083,N_8504,N_8633);
xor U9084 (N_9084,N_8713,N_8708);
or U9085 (N_9085,N_8596,N_8565);
and U9086 (N_9086,N_8836,N_8890);
nor U9087 (N_9087,N_8902,N_8629);
nand U9088 (N_9088,N_8927,N_8829);
or U9089 (N_9089,N_8818,N_8951);
nand U9090 (N_9090,N_8903,N_8560);
nor U9091 (N_9091,N_8786,N_8923);
nand U9092 (N_9092,N_8661,N_8879);
xor U9093 (N_9093,N_8655,N_8689);
and U9094 (N_9094,N_8860,N_8704);
xor U9095 (N_9095,N_8777,N_8800);
and U9096 (N_9096,N_8814,N_8557);
and U9097 (N_9097,N_8844,N_8746);
nor U9098 (N_9098,N_8915,N_8510);
or U9099 (N_9099,N_8715,N_8757);
nor U9100 (N_9100,N_8877,N_8541);
and U9101 (N_9101,N_8628,N_8716);
and U9102 (N_9102,N_8516,N_8861);
nand U9103 (N_9103,N_8943,N_8797);
xor U9104 (N_9104,N_8570,N_8866);
and U9105 (N_9105,N_8564,N_8588);
or U9106 (N_9106,N_8651,N_8589);
or U9107 (N_9107,N_8575,N_8733);
nor U9108 (N_9108,N_8676,N_8522);
xor U9109 (N_9109,N_8582,N_8992);
or U9110 (N_9110,N_8736,N_8990);
or U9111 (N_9111,N_8552,N_8936);
xor U9112 (N_9112,N_8958,N_8807);
or U9113 (N_9113,N_8864,N_8546);
or U9114 (N_9114,N_8540,N_8679);
nand U9115 (N_9115,N_8648,N_8725);
or U9116 (N_9116,N_8723,N_8791);
and U9117 (N_9117,N_8645,N_8530);
xnor U9118 (N_9118,N_8626,N_8538);
and U9119 (N_9119,N_8520,N_8681);
or U9120 (N_9120,N_8975,N_8697);
and U9121 (N_9121,N_8718,N_8962);
nand U9122 (N_9122,N_8873,N_8885);
or U9123 (N_9123,N_8785,N_8868);
nor U9124 (N_9124,N_8506,N_8898);
and U9125 (N_9125,N_8773,N_8982);
and U9126 (N_9126,N_8664,N_8707);
xor U9127 (N_9127,N_8688,N_8605);
nand U9128 (N_9128,N_8803,N_8642);
nor U9129 (N_9129,N_8770,N_8796);
nand U9130 (N_9130,N_8764,N_8537);
xor U9131 (N_9131,N_8529,N_8896);
nor U9132 (N_9132,N_8880,N_8690);
xor U9133 (N_9133,N_8692,N_8831);
or U9134 (N_9134,N_8906,N_8801);
or U9135 (N_9135,N_8780,N_8942);
nor U9136 (N_9136,N_8729,N_8531);
nor U9137 (N_9137,N_8940,N_8854);
or U9138 (N_9138,N_8815,N_8793);
and U9139 (N_9139,N_8737,N_8977);
or U9140 (N_9140,N_8650,N_8603);
or U9141 (N_9141,N_8630,N_8532);
or U9142 (N_9142,N_8983,N_8830);
or U9143 (N_9143,N_8678,N_8549);
and U9144 (N_9144,N_8521,N_8993);
xnor U9145 (N_9145,N_8886,N_8505);
nand U9146 (N_9146,N_8535,N_8508);
xor U9147 (N_9147,N_8996,N_8616);
and U9148 (N_9148,N_8811,N_8918);
or U9149 (N_9149,N_8609,N_8507);
nor U9150 (N_9150,N_8635,N_8675);
nor U9151 (N_9151,N_8663,N_8888);
nor U9152 (N_9152,N_8614,N_8536);
nor U9153 (N_9153,N_8594,N_8624);
nor U9154 (N_9154,N_8602,N_8671);
and U9155 (N_9155,N_8514,N_8759);
or U9156 (N_9156,N_8761,N_8572);
or U9157 (N_9157,N_8558,N_8863);
nor U9158 (N_9158,N_8677,N_8585);
nand U9159 (N_9159,N_8578,N_8592);
xor U9160 (N_9160,N_8590,N_8502);
nand U9161 (N_9161,N_8528,N_8835);
or U9162 (N_9162,N_8855,N_8889);
nand U9163 (N_9163,N_8787,N_8895);
and U9164 (N_9164,N_8795,N_8969);
nand U9165 (N_9165,N_8670,N_8576);
xor U9166 (N_9166,N_8710,N_8955);
nor U9167 (N_9167,N_8910,N_8832);
xor U9168 (N_9168,N_8887,N_8837);
or U9169 (N_9169,N_8573,N_8775);
xnor U9170 (N_9170,N_8980,N_8749);
and U9171 (N_9171,N_8599,N_8730);
nand U9172 (N_9172,N_8631,N_8961);
xor U9173 (N_9173,N_8695,N_8778);
and U9174 (N_9174,N_8948,N_8618);
nand U9175 (N_9175,N_8909,N_8772);
nand U9176 (N_9176,N_8539,N_8919);
and U9177 (N_9177,N_8953,N_8833);
or U9178 (N_9178,N_8825,N_8834);
and U9179 (N_9179,N_8867,N_8619);
or U9180 (N_9180,N_8735,N_8840);
and U9181 (N_9181,N_8740,N_8525);
nand U9182 (N_9182,N_8666,N_8714);
nor U9183 (N_9183,N_8950,N_8921);
xnor U9184 (N_9184,N_8646,N_8806);
or U9185 (N_9185,N_8584,N_8513);
nand U9186 (N_9186,N_8872,N_8846);
xor U9187 (N_9187,N_8883,N_8912);
and U9188 (N_9188,N_8792,N_8700);
xor U9189 (N_9189,N_8758,N_8995);
nor U9190 (N_9190,N_8869,N_8760);
nand U9191 (N_9191,N_8967,N_8856);
or U9192 (N_9192,N_8933,N_8997);
nand U9193 (N_9193,N_8620,N_8698);
nor U9194 (N_9194,N_8822,N_8518);
nor U9195 (N_9195,N_8586,N_8617);
xor U9196 (N_9196,N_8971,N_8627);
nor U9197 (N_9197,N_8765,N_8702);
or U9198 (N_9198,N_8638,N_8914);
nor U9199 (N_9199,N_8974,N_8696);
nor U9200 (N_9200,N_8568,N_8544);
and U9201 (N_9201,N_8799,N_8901);
xor U9202 (N_9202,N_8701,N_8878);
xor U9203 (N_9203,N_8722,N_8579);
and U9204 (N_9204,N_8994,N_8781);
nor U9205 (N_9205,N_8845,N_8691);
or U9206 (N_9206,N_8587,N_8881);
nor U9207 (N_9207,N_8551,N_8728);
or U9208 (N_9208,N_8908,N_8636);
or U9209 (N_9209,N_8668,N_8649);
or U9210 (N_9210,N_8554,N_8768);
and U9211 (N_9211,N_8892,N_8674);
nand U9212 (N_9212,N_8577,N_8598);
or U9213 (N_9213,N_8917,N_8944);
nand U9214 (N_9214,N_8988,N_8972);
and U9215 (N_9215,N_8680,N_8712);
or U9216 (N_9216,N_8685,N_8744);
or U9217 (N_9217,N_8986,N_8745);
and U9218 (N_9218,N_8929,N_8763);
and U9219 (N_9219,N_8920,N_8519);
and U9220 (N_9220,N_8534,N_8524);
or U9221 (N_9221,N_8500,N_8739);
or U9222 (N_9222,N_8934,N_8747);
xnor U9223 (N_9223,N_8600,N_8694);
or U9224 (N_9224,N_8899,N_8905);
xnor U9225 (N_9225,N_8523,N_8794);
nand U9226 (N_9226,N_8820,N_8752);
nor U9227 (N_9227,N_8973,N_8946);
and U9228 (N_9228,N_8606,N_8684);
or U9229 (N_9229,N_8719,N_8876);
xnor U9230 (N_9230,N_8904,N_8979);
nand U9231 (N_9231,N_8947,N_8808);
xor U9232 (N_9232,N_8637,N_8595);
nand U9233 (N_9233,N_8526,N_8897);
or U9234 (N_9234,N_8826,N_8501);
xor U9235 (N_9235,N_8652,N_8987);
or U9236 (N_9236,N_8928,N_8687);
xnor U9237 (N_9237,N_8859,N_8566);
nor U9238 (N_9238,N_8809,N_8693);
nor U9239 (N_9239,N_8999,N_8643);
nor U9240 (N_9240,N_8610,N_8865);
nand U9241 (N_9241,N_8790,N_8569);
nand U9242 (N_9242,N_8511,N_8732);
or U9243 (N_9243,N_8937,N_8726);
or U9244 (N_9244,N_8870,N_8926);
and U9245 (N_9245,N_8853,N_8805);
xnor U9246 (N_9246,N_8553,N_8717);
xor U9247 (N_9247,N_8985,N_8581);
or U9248 (N_9248,N_8656,N_8819);
nor U9249 (N_9249,N_8774,N_8613);
nand U9250 (N_9250,N_8540,N_8700);
or U9251 (N_9251,N_8701,N_8905);
xor U9252 (N_9252,N_8932,N_8726);
nand U9253 (N_9253,N_8890,N_8791);
or U9254 (N_9254,N_8549,N_8573);
xor U9255 (N_9255,N_8601,N_8742);
and U9256 (N_9256,N_8609,N_8565);
nor U9257 (N_9257,N_8754,N_8878);
or U9258 (N_9258,N_8681,N_8603);
nor U9259 (N_9259,N_8956,N_8611);
nor U9260 (N_9260,N_8903,N_8669);
nand U9261 (N_9261,N_8520,N_8894);
xor U9262 (N_9262,N_8637,N_8932);
or U9263 (N_9263,N_8909,N_8722);
or U9264 (N_9264,N_8583,N_8555);
nor U9265 (N_9265,N_8699,N_8883);
xnor U9266 (N_9266,N_8570,N_8648);
and U9267 (N_9267,N_8684,N_8521);
nor U9268 (N_9268,N_8927,N_8514);
or U9269 (N_9269,N_8569,N_8961);
nor U9270 (N_9270,N_8830,N_8892);
xnor U9271 (N_9271,N_8892,N_8519);
or U9272 (N_9272,N_8654,N_8527);
and U9273 (N_9273,N_8825,N_8929);
nor U9274 (N_9274,N_8879,N_8558);
xor U9275 (N_9275,N_8969,N_8687);
nor U9276 (N_9276,N_8941,N_8589);
or U9277 (N_9277,N_8769,N_8916);
xor U9278 (N_9278,N_8945,N_8641);
nor U9279 (N_9279,N_8696,N_8929);
or U9280 (N_9280,N_8796,N_8563);
nand U9281 (N_9281,N_8865,N_8930);
xnor U9282 (N_9282,N_8903,N_8778);
xor U9283 (N_9283,N_8623,N_8624);
or U9284 (N_9284,N_8646,N_8997);
nand U9285 (N_9285,N_8890,N_8571);
and U9286 (N_9286,N_8910,N_8711);
nand U9287 (N_9287,N_8855,N_8781);
or U9288 (N_9288,N_8670,N_8558);
or U9289 (N_9289,N_8503,N_8908);
or U9290 (N_9290,N_8520,N_8946);
nand U9291 (N_9291,N_8923,N_8538);
and U9292 (N_9292,N_8972,N_8791);
or U9293 (N_9293,N_8764,N_8677);
and U9294 (N_9294,N_8727,N_8759);
xnor U9295 (N_9295,N_8845,N_8614);
and U9296 (N_9296,N_8736,N_8944);
nand U9297 (N_9297,N_8945,N_8561);
or U9298 (N_9298,N_8961,N_8754);
nand U9299 (N_9299,N_8580,N_8880);
and U9300 (N_9300,N_8723,N_8983);
xnor U9301 (N_9301,N_8897,N_8971);
nor U9302 (N_9302,N_8780,N_8928);
nand U9303 (N_9303,N_8835,N_8739);
and U9304 (N_9304,N_8757,N_8770);
xnor U9305 (N_9305,N_8645,N_8575);
or U9306 (N_9306,N_8684,N_8718);
xnor U9307 (N_9307,N_8958,N_8775);
or U9308 (N_9308,N_8775,N_8893);
nor U9309 (N_9309,N_8649,N_8582);
xor U9310 (N_9310,N_8647,N_8718);
and U9311 (N_9311,N_8669,N_8642);
or U9312 (N_9312,N_8536,N_8788);
nand U9313 (N_9313,N_8812,N_8827);
or U9314 (N_9314,N_8538,N_8966);
or U9315 (N_9315,N_8547,N_8703);
and U9316 (N_9316,N_8858,N_8831);
xor U9317 (N_9317,N_8719,N_8940);
or U9318 (N_9318,N_8982,N_8989);
or U9319 (N_9319,N_8974,N_8731);
xor U9320 (N_9320,N_8581,N_8848);
nand U9321 (N_9321,N_8538,N_8618);
nand U9322 (N_9322,N_8529,N_8579);
nor U9323 (N_9323,N_8730,N_8762);
or U9324 (N_9324,N_8953,N_8571);
xnor U9325 (N_9325,N_8554,N_8997);
nand U9326 (N_9326,N_8980,N_8797);
nand U9327 (N_9327,N_8874,N_8539);
nor U9328 (N_9328,N_8756,N_8559);
xor U9329 (N_9329,N_8783,N_8932);
xnor U9330 (N_9330,N_8910,N_8729);
nor U9331 (N_9331,N_8626,N_8649);
nand U9332 (N_9332,N_8846,N_8866);
nor U9333 (N_9333,N_8543,N_8834);
and U9334 (N_9334,N_8607,N_8863);
xor U9335 (N_9335,N_8742,N_8568);
nand U9336 (N_9336,N_8511,N_8852);
and U9337 (N_9337,N_8929,N_8952);
xor U9338 (N_9338,N_8804,N_8779);
xor U9339 (N_9339,N_8552,N_8958);
nor U9340 (N_9340,N_8528,N_8802);
or U9341 (N_9341,N_8713,N_8894);
or U9342 (N_9342,N_8910,N_8957);
nor U9343 (N_9343,N_8864,N_8938);
or U9344 (N_9344,N_8974,N_8820);
and U9345 (N_9345,N_8987,N_8993);
or U9346 (N_9346,N_8940,N_8646);
and U9347 (N_9347,N_8912,N_8763);
nand U9348 (N_9348,N_8635,N_8917);
nand U9349 (N_9349,N_8702,N_8675);
xnor U9350 (N_9350,N_8857,N_8873);
nand U9351 (N_9351,N_8880,N_8608);
nor U9352 (N_9352,N_8657,N_8686);
and U9353 (N_9353,N_8879,N_8552);
or U9354 (N_9354,N_8529,N_8715);
and U9355 (N_9355,N_8661,N_8521);
nand U9356 (N_9356,N_8931,N_8604);
xor U9357 (N_9357,N_8709,N_8974);
and U9358 (N_9358,N_8819,N_8769);
nor U9359 (N_9359,N_8944,N_8521);
or U9360 (N_9360,N_8671,N_8636);
and U9361 (N_9361,N_8655,N_8864);
or U9362 (N_9362,N_8824,N_8632);
nand U9363 (N_9363,N_8782,N_8633);
xor U9364 (N_9364,N_8817,N_8673);
and U9365 (N_9365,N_8709,N_8687);
nand U9366 (N_9366,N_8868,N_8530);
and U9367 (N_9367,N_8643,N_8537);
or U9368 (N_9368,N_8515,N_8624);
and U9369 (N_9369,N_8753,N_8740);
nand U9370 (N_9370,N_8606,N_8970);
and U9371 (N_9371,N_8989,N_8822);
xnor U9372 (N_9372,N_8962,N_8864);
or U9373 (N_9373,N_8736,N_8896);
nand U9374 (N_9374,N_8986,N_8517);
xnor U9375 (N_9375,N_8699,N_8862);
xnor U9376 (N_9376,N_8722,N_8532);
nand U9377 (N_9377,N_8662,N_8642);
or U9378 (N_9378,N_8576,N_8621);
nor U9379 (N_9379,N_8654,N_8669);
or U9380 (N_9380,N_8783,N_8680);
or U9381 (N_9381,N_8719,N_8594);
or U9382 (N_9382,N_8558,N_8823);
xor U9383 (N_9383,N_8903,N_8842);
nor U9384 (N_9384,N_8554,N_8806);
xnor U9385 (N_9385,N_8520,N_8560);
and U9386 (N_9386,N_8671,N_8781);
or U9387 (N_9387,N_8516,N_8725);
nand U9388 (N_9388,N_8676,N_8778);
and U9389 (N_9389,N_8600,N_8786);
xor U9390 (N_9390,N_8634,N_8969);
or U9391 (N_9391,N_8568,N_8786);
or U9392 (N_9392,N_8588,N_8825);
or U9393 (N_9393,N_8926,N_8586);
nand U9394 (N_9394,N_8667,N_8734);
nand U9395 (N_9395,N_8749,N_8901);
xnor U9396 (N_9396,N_8884,N_8544);
and U9397 (N_9397,N_8897,N_8768);
or U9398 (N_9398,N_8819,N_8785);
and U9399 (N_9399,N_8627,N_8786);
nor U9400 (N_9400,N_8563,N_8666);
nor U9401 (N_9401,N_8651,N_8856);
or U9402 (N_9402,N_8664,N_8734);
nor U9403 (N_9403,N_8542,N_8715);
and U9404 (N_9404,N_8769,N_8650);
xor U9405 (N_9405,N_8692,N_8803);
nor U9406 (N_9406,N_8652,N_8551);
and U9407 (N_9407,N_8840,N_8995);
xnor U9408 (N_9408,N_8606,N_8680);
nor U9409 (N_9409,N_8651,N_8642);
or U9410 (N_9410,N_8936,N_8772);
xor U9411 (N_9411,N_8914,N_8771);
and U9412 (N_9412,N_8857,N_8861);
xnor U9413 (N_9413,N_8559,N_8987);
nor U9414 (N_9414,N_8566,N_8894);
and U9415 (N_9415,N_8556,N_8962);
and U9416 (N_9416,N_8573,N_8823);
and U9417 (N_9417,N_8871,N_8859);
and U9418 (N_9418,N_8827,N_8726);
nor U9419 (N_9419,N_8577,N_8931);
and U9420 (N_9420,N_8547,N_8820);
nand U9421 (N_9421,N_8531,N_8965);
xor U9422 (N_9422,N_8971,N_8737);
and U9423 (N_9423,N_8511,N_8570);
and U9424 (N_9424,N_8932,N_8944);
nor U9425 (N_9425,N_8750,N_8643);
xor U9426 (N_9426,N_8900,N_8631);
xnor U9427 (N_9427,N_8580,N_8501);
nor U9428 (N_9428,N_8579,N_8821);
or U9429 (N_9429,N_8717,N_8908);
nor U9430 (N_9430,N_8899,N_8557);
and U9431 (N_9431,N_8710,N_8698);
or U9432 (N_9432,N_8836,N_8534);
xor U9433 (N_9433,N_8854,N_8531);
or U9434 (N_9434,N_8690,N_8959);
and U9435 (N_9435,N_8926,N_8729);
nor U9436 (N_9436,N_8540,N_8558);
nand U9437 (N_9437,N_8723,N_8812);
and U9438 (N_9438,N_8961,N_8922);
and U9439 (N_9439,N_8712,N_8905);
nand U9440 (N_9440,N_8744,N_8729);
nor U9441 (N_9441,N_8503,N_8560);
nor U9442 (N_9442,N_8674,N_8782);
nand U9443 (N_9443,N_8507,N_8700);
nor U9444 (N_9444,N_8820,N_8749);
and U9445 (N_9445,N_8507,N_8845);
and U9446 (N_9446,N_8608,N_8503);
nand U9447 (N_9447,N_8912,N_8675);
xor U9448 (N_9448,N_8812,N_8803);
xor U9449 (N_9449,N_8906,N_8550);
and U9450 (N_9450,N_8583,N_8975);
or U9451 (N_9451,N_8828,N_8751);
xor U9452 (N_9452,N_8980,N_8896);
nand U9453 (N_9453,N_8937,N_8660);
xor U9454 (N_9454,N_8708,N_8748);
nor U9455 (N_9455,N_8979,N_8881);
or U9456 (N_9456,N_8773,N_8880);
nor U9457 (N_9457,N_8609,N_8804);
nand U9458 (N_9458,N_8840,N_8719);
nor U9459 (N_9459,N_8517,N_8567);
and U9460 (N_9460,N_8648,N_8807);
xor U9461 (N_9461,N_8932,N_8601);
or U9462 (N_9462,N_8994,N_8869);
nand U9463 (N_9463,N_8895,N_8821);
xor U9464 (N_9464,N_8777,N_8559);
nand U9465 (N_9465,N_8749,N_8908);
and U9466 (N_9466,N_8774,N_8749);
or U9467 (N_9467,N_8518,N_8605);
nand U9468 (N_9468,N_8769,N_8550);
nor U9469 (N_9469,N_8714,N_8530);
and U9470 (N_9470,N_8583,N_8686);
or U9471 (N_9471,N_8743,N_8808);
or U9472 (N_9472,N_8983,N_8596);
or U9473 (N_9473,N_8887,N_8667);
nor U9474 (N_9474,N_8679,N_8664);
or U9475 (N_9475,N_8832,N_8547);
nor U9476 (N_9476,N_8947,N_8716);
nand U9477 (N_9477,N_8810,N_8699);
xnor U9478 (N_9478,N_8602,N_8519);
nor U9479 (N_9479,N_8800,N_8668);
or U9480 (N_9480,N_8834,N_8609);
and U9481 (N_9481,N_8778,N_8987);
and U9482 (N_9482,N_8517,N_8503);
nand U9483 (N_9483,N_8903,N_8952);
nor U9484 (N_9484,N_8523,N_8805);
nor U9485 (N_9485,N_8984,N_8688);
nor U9486 (N_9486,N_8621,N_8619);
nand U9487 (N_9487,N_8673,N_8960);
xor U9488 (N_9488,N_8858,N_8678);
xor U9489 (N_9489,N_8799,N_8927);
or U9490 (N_9490,N_8901,N_8515);
and U9491 (N_9491,N_8967,N_8684);
nand U9492 (N_9492,N_8576,N_8513);
nor U9493 (N_9493,N_8754,N_8875);
xnor U9494 (N_9494,N_8609,N_8808);
nor U9495 (N_9495,N_8911,N_8550);
and U9496 (N_9496,N_8708,N_8683);
nand U9497 (N_9497,N_8524,N_8923);
nand U9498 (N_9498,N_8618,N_8836);
and U9499 (N_9499,N_8683,N_8693);
or U9500 (N_9500,N_9388,N_9250);
xor U9501 (N_9501,N_9286,N_9288);
and U9502 (N_9502,N_9271,N_9387);
xnor U9503 (N_9503,N_9279,N_9383);
nand U9504 (N_9504,N_9043,N_9304);
and U9505 (N_9505,N_9010,N_9320);
nand U9506 (N_9506,N_9321,N_9448);
or U9507 (N_9507,N_9216,N_9183);
nand U9508 (N_9508,N_9020,N_9494);
or U9509 (N_9509,N_9422,N_9102);
nand U9510 (N_9510,N_9351,N_9088);
xnor U9511 (N_9511,N_9352,N_9360);
xnor U9512 (N_9512,N_9218,N_9457);
nand U9513 (N_9513,N_9394,N_9212);
nand U9514 (N_9514,N_9372,N_9246);
or U9515 (N_9515,N_9342,N_9385);
xnor U9516 (N_9516,N_9478,N_9176);
xnor U9517 (N_9517,N_9065,N_9228);
or U9518 (N_9518,N_9204,N_9337);
or U9519 (N_9519,N_9235,N_9244);
nor U9520 (N_9520,N_9135,N_9336);
nor U9521 (N_9521,N_9042,N_9488);
xnor U9522 (N_9522,N_9446,N_9081);
or U9523 (N_9523,N_9089,N_9078);
and U9524 (N_9524,N_9048,N_9358);
and U9525 (N_9525,N_9229,N_9301);
and U9526 (N_9526,N_9150,N_9164);
xnor U9527 (N_9527,N_9289,N_9362);
nor U9528 (N_9528,N_9124,N_9057);
nor U9529 (N_9529,N_9261,N_9409);
nand U9530 (N_9530,N_9361,N_9155);
nor U9531 (N_9531,N_9047,N_9171);
nand U9532 (N_9532,N_9044,N_9364);
nor U9533 (N_9533,N_9412,N_9177);
and U9534 (N_9534,N_9230,N_9157);
or U9535 (N_9535,N_9138,N_9455);
or U9536 (N_9536,N_9029,N_9463);
and U9537 (N_9537,N_9474,N_9077);
xor U9538 (N_9538,N_9069,N_9175);
nand U9539 (N_9539,N_9083,N_9438);
or U9540 (N_9540,N_9419,N_9114);
or U9541 (N_9541,N_9298,N_9126);
xnor U9542 (N_9542,N_9379,N_9240);
or U9543 (N_9543,N_9134,N_9172);
and U9544 (N_9544,N_9009,N_9169);
xnor U9545 (N_9545,N_9079,N_9315);
xor U9546 (N_9546,N_9165,N_9384);
nor U9547 (N_9547,N_9130,N_9295);
and U9548 (N_9548,N_9190,N_9005);
nand U9549 (N_9549,N_9436,N_9146);
nor U9550 (N_9550,N_9003,N_9173);
nand U9551 (N_9551,N_9015,N_9461);
xor U9552 (N_9552,N_9382,N_9260);
nor U9553 (N_9553,N_9162,N_9205);
and U9554 (N_9554,N_9050,N_9203);
and U9555 (N_9555,N_9011,N_9008);
xor U9556 (N_9556,N_9071,N_9450);
xnor U9557 (N_9557,N_9002,N_9255);
nand U9558 (N_9558,N_9267,N_9073);
nor U9559 (N_9559,N_9094,N_9392);
nor U9560 (N_9560,N_9442,N_9101);
nand U9561 (N_9561,N_9366,N_9319);
or U9562 (N_9562,N_9152,N_9431);
xnor U9563 (N_9563,N_9327,N_9119);
xor U9564 (N_9564,N_9282,N_9389);
nand U9565 (N_9565,N_9132,N_9391);
nand U9566 (N_9566,N_9443,N_9437);
nand U9567 (N_9567,N_9340,N_9468);
nor U9568 (N_9568,N_9280,N_9377);
xnor U9569 (N_9569,N_9410,N_9420);
nor U9570 (N_9570,N_9493,N_9178);
xnor U9571 (N_9571,N_9247,N_9117);
nand U9572 (N_9572,N_9381,N_9365);
or U9573 (N_9573,N_9041,N_9125);
nor U9574 (N_9574,N_9118,N_9451);
or U9575 (N_9575,N_9287,N_9181);
nand U9576 (N_9576,N_9056,N_9241);
xnor U9577 (N_9577,N_9158,N_9332);
and U9578 (N_9578,N_9033,N_9215);
and U9579 (N_9579,N_9371,N_9245);
or U9580 (N_9580,N_9021,N_9100);
nor U9581 (N_9581,N_9060,N_9309);
and U9582 (N_9582,N_9355,N_9080);
or U9583 (N_9583,N_9004,N_9482);
nor U9584 (N_9584,N_9294,N_9166);
and U9585 (N_9585,N_9471,N_9254);
nand U9586 (N_9586,N_9022,N_9053);
nor U9587 (N_9587,N_9236,N_9122);
nand U9588 (N_9588,N_9328,N_9091);
or U9589 (N_9589,N_9445,N_9311);
and U9590 (N_9590,N_9268,N_9202);
xnor U9591 (N_9591,N_9227,N_9490);
nor U9592 (N_9592,N_9075,N_9434);
and U9593 (N_9593,N_9061,N_9472);
xnor U9594 (N_9594,N_9108,N_9313);
and U9595 (N_9595,N_9338,N_9092);
or U9596 (N_9596,N_9395,N_9017);
xor U9597 (N_9597,N_9226,N_9322);
or U9598 (N_9598,N_9481,N_9334);
xnor U9599 (N_9599,N_9019,N_9055);
or U9600 (N_9600,N_9234,N_9084);
and U9601 (N_9601,N_9037,N_9428);
nand U9602 (N_9602,N_9263,N_9459);
xor U9603 (N_9603,N_9099,N_9120);
nand U9604 (N_9604,N_9142,N_9034);
and U9605 (N_9605,N_9277,N_9207);
nor U9606 (N_9606,N_9310,N_9303);
nor U9607 (N_9607,N_9112,N_9486);
xnor U9608 (N_9608,N_9344,N_9014);
or U9609 (N_9609,N_9390,N_9262);
or U9610 (N_9610,N_9469,N_9074);
nand U9611 (N_9611,N_9188,N_9432);
nand U9612 (N_9612,N_9477,N_9440);
nor U9613 (N_9613,N_9098,N_9470);
or U9614 (N_9614,N_9145,N_9306);
nor U9615 (N_9615,N_9483,N_9411);
nand U9616 (N_9616,N_9375,N_9049);
nor U9617 (N_9617,N_9148,N_9035);
and U9618 (N_9618,N_9233,N_9144);
nor U9619 (N_9619,N_9492,N_9040);
xnor U9620 (N_9620,N_9425,N_9012);
xnor U9621 (N_9621,N_9479,N_9269);
and U9622 (N_9622,N_9453,N_9484);
nor U9623 (N_9623,N_9182,N_9249);
or U9624 (N_9624,N_9160,N_9059);
and U9625 (N_9625,N_9219,N_9072);
and U9626 (N_9626,N_9128,N_9025);
xnor U9627 (N_9627,N_9210,N_9464);
nand U9628 (N_9628,N_9110,N_9376);
xor U9629 (N_9629,N_9189,N_9300);
xnor U9630 (N_9630,N_9184,N_9283);
nand U9631 (N_9631,N_9347,N_9127);
or U9632 (N_9632,N_9259,N_9076);
xnor U9633 (N_9633,N_9285,N_9386);
nor U9634 (N_9634,N_9416,N_9105);
and U9635 (N_9635,N_9113,N_9350);
xnor U9636 (N_9636,N_9496,N_9213);
nand U9637 (N_9637,N_9414,N_9317);
and U9638 (N_9638,N_9027,N_9222);
nor U9639 (N_9639,N_9497,N_9238);
or U9640 (N_9640,N_9103,N_9220);
xnor U9641 (N_9641,N_9307,N_9147);
and U9642 (N_9642,N_9449,N_9380);
and U9643 (N_9643,N_9357,N_9243);
and U9644 (N_9644,N_9368,N_9179);
and U9645 (N_9645,N_9064,N_9131);
nor U9646 (N_9646,N_9403,N_9199);
and U9647 (N_9647,N_9324,N_9123);
xor U9648 (N_9648,N_9167,N_9133);
xnor U9649 (N_9649,N_9097,N_9096);
nand U9650 (N_9650,N_9136,N_9067);
nand U9651 (N_9651,N_9281,N_9062);
or U9652 (N_9652,N_9153,N_9404);
nor U9653 (N_9653,N_9149,N_9297);
or U9654 (N_9654,N_9276,N_9242);
or U9655 (N_9655,N_9168,N_9341);
or U9656 (N_9656,N_9185,N_9429);
xor U9657 (N_9657,N_9139,N_9001);
or U9658 (N_9658,N_9367,N_9209);
xnor U9659 (N_9659,N_9023,N_9460);
nor U9660 (N_9660,N_9353,N_9423);
nand U9661 (N_9661,N_9273,N_9191);
xor U9662 (N_9662,N_9396,N_9095);
or U9663 (N_9663,N_9299,N_9121);
nor U9664 (N_9664,N_9346,N_9402);
and U9665 (N_9665,N_9196,N_9331);
xor U9666 (N_9666,N_9417,N_9054);
or U9667 (N_9667,N_9430,N_9441);
or U9668 (N_9668,N_9284,N_9109);
or U9669 (N_9669,N_9296,N_9480);
xor U9670 (N_9670,N_9323,N_9456);
nor U9671 (N_9671,N_9225,N_9454);
nand U9672 (N_9672,N_9433,N_9292);
nor U9673 (N_9673,N_9266,N_9485);
or U9674 (N_9674,N_9406,N_9330);
or U9675 (N_9675,N_9031,N_9413);
xnor U9676 (N_9676,N_9143,N_9264);
or U9677 (N_9677,N_9329,N_9293);
xnor U9678 (N_9678,N_9195,N_9275);
nor U9679 (N_9679,N_9270,N_9418);
and U9680 (N_9680,N_9192,N_9174);
nand U9681 (N_9681,N_9265,N_9051);
nor U9682 (N_9682,N_9200,N_9415);
xnor U9683 (N_9683,N_9013,N_9087);
xnor U9684 (N_9684,N_9038,N_9107);
or U9685 (N_9685,N_9217,N_9349);
and U9686 (N_9686,N_9186,N_9070);
and U9687 (N_9687,N_9066,N_9316);
nand U9688 (N_9688,N_9489,N_9248);
nor U9689 (N_9689,N_9405,N_9326);
nand U9690 (N_9690,N_9163,N_9274);
xnor U9691 (N_9691,N_9198,N_9032);
or U9692 (N_9692,N_9024,N_9398);
or U9693 (N_9693,N_9039,N_9252);
xor U9694 (N_9694,N_9272,N_9221);
nand U9695 (N_9695,N_9487,N_9399);
nand U9696 (N_9696,N_9104,N_9239);
xnor U9697 (N_9697,N_9028,N_9116);
or U9698 (N_9698,N_9256,N_9278);
nor U9699 (N_9699,N_9251,N_9231);
nand U9700 (N_9700,N_9427,N_9063);
xor U9701 (N_9701,N_9421,N_9090);
and U9702 (N_9702,N_9086,N_9036);
or U9703 (N_9703,N_9465,N_9335);
nor U9704 (N_9704,N_9206,N_9348);
nand U9705 (N_9705,N_9466,N_9214);
xnor U9706 (N_9706,N_9141,N_9154);
nand U9707 (N_9707,N_9016,N_9237);
or U9708 (N_9708,N_9211,N_9170);
and U9709 (N_9709,N_9302,N_9452);
and U9710 (N_9710,N_9068,N_9426);
or U9711 (N_9711,N_9318,N_9082);
or U9712 (N_9712,N_9193,N_9224);
nand U9713 (N_9713,N_9491,N_9018);
nand U9714 (N_9714,N_9499,N_9444);
and U9715 (N_9715,N_9354,N_9339);
xor U9716 (N_9716,N_9314,N_9129);
xnor U9717 (N_9717,N_9111,N_9106);
and U9718 (N_9718,N_9058,N_9151);
or U9719 (N_9719,N_9046,N_9253);
nor U9720 (N_9720,N_9258,N_9201);
xor U9721 (N_9721,N_9397,N_9333);
nand U9722 (N_9722,N_9208,N_9393);
nand U9723 (N_9723,N_9378,N_9439);
and U9724 (N_9724,N_9356,N_9407);
or U9725 (N_9725,N_9290,N_9363);
and U9726 (N_9726,N_9291,N_9401);
and U9727 (N_9727,N_9312,N_9475);
and U9728 (N_9728,N_9159,N_9369);
nor U9729 (N_9729,N_9400,N_9085);
nand U9730 (N_9730,N_9345,N_9498);
or U9731 (N_9731,N_9000,N_9045);
and U9732 (N_9732,N_9180,N_9156);
nand U9733 (N_9733,N_9030,N_9458);
nand U9734 (N_9734,N_9161,N_9374);
nand U9735 (N_9735,N_9197,N_9476);
or U9736 (N_9736,N_9140,N_9447);
and U9737 (N_9737,N_9408,N_9435);
nand U9738 (N_9738,N_9495,N_9137);
nor U9739 (N_9739,N_9308,N_9232);
xor U9740 (N_9740,N_9325,N_9370);
and U9741 (N_9741,N_9343,N_9467);
nor U9742 (N_9742,N_9006,N_9093);
and U9743 (N_9743,N_9359,N_9187);
or U9744 (N_9744,N_9194,N_9026);
or U9745 (N_9745,N_9052,N_9007);
nand U9746 (N_9746,N_9257,N_9305);
and U9747 (N_9747,N_9373,N_9115);
or U9748 (N_9748,N_9223,N_9473);
nor U9749 (N_9749,N_9424,N_9462);
or U9750 (N_9750,N_9178,N_9367);
nand U9751 (N_9751,N_9134,N_9474);
nand U9752 (N_9752,N_9279,N_9345);
nand U9753 (N_9753,N_9429,N_9193);
nand U9754 (N_9754,N_9108,N_9024);
or U9755 (N_9755,N_9159,N_9191);
or U9756 (N_9756,N_9296,N_9129);
nor U9757 (N_9757,N_9209,N_9423);
xor U9758 (N_9758,N_9478,N_9166);
nand U9759 (N_9759,N_9024,N_9450);
nor U9760 (N_9760,N_9194,N_9156);
or U9761 (N_9761,N_9414,N_9382);
nor U9762 (N_9762,N_9172,N_9379);
nor U9763 (N_9763,N_9432,N_9114);
nand U9764 (N_9764,N_9363,N_9282);
nor U9765 (N_9765,N_9292,N_9104);
or U9766 (N_9766,N_9446,N_9057);
or U9767 (N_9767,N_9164,N_9454);
nand U9768 (N_9768,N_9097,N_9296);
nand U9769 (N_9769,N_9183,N_9417);
nand U9770 (N_9770,N_9321,N_9218);
xnor U9771 (N_9771,N_9418,N_9481);
nor U9772 (N_9772,N_9001,N_9016);
and U9773 (N_9773,N_9131,N_9188);
and U9774 (N_9774,N_9317,N_9025);
nand U9775 (N_9775,N_9359,N_9499);
nor U9776 (N_9776,N_9332,N_9100);
nand U9777 (N_9777,N_9391,N_9033);
xnor U9778 (N_9778,N_9148,N_9276);
nor U9779 (N_9779,N_9082,N_9439);
and U9780 (N_9780,N_9484,N_9366);
xor U9781 (N_9781,N_9269,N_9206);
and U9782 (N_9782,N_9349,N_9138);
nand U9783 (N_9783,N_9010,N_9146);
nand U9784 (N_9784,N_9285,N_9457);
xnor U9785 (N_9785,N_9465,N_9069);
and U9786 (N_9786,N_9380,N_9122);
nor U9787 (N_9787,N_9444,N_9120);
nor U9788 (N_9788,N_9297,N_9185);
and U9789 (N_9789,N_9188,N_9465);
xor U9790 (N_9790,N_9035,N_9341);
and U9791 (N_9791,N_9369,N_9047);
and U9792 (N_9792,N_9175,N_9281);
and U9793 (N_9793,N_9101,N_9478);
and U9794 (N_9794,N_9173,N_9228);
and U9795 (N_9795,N_9431,N_9023);
and U9796 (N_9796,N_9190,N_9209);
nor U9797 (N_9797,N_9094,N_9120);
nor U9798 (N_9798,N_9242,N_9009);
and U9799 (N_9799,N_9163,N_9246);
nand U9800 (N_9800,N_9071,N_9429);
and U9801 (N_9801,N_9212,N_9192);
nand U9802 (N_9802,N_9237,N_9454);
xnor U9803 (N_9803,N_9265,N_9066);
nor U9804 (N_9804,N_9140,N_9146);
nor U9805 (N_9805,N_9345,N_9217);
nand U9806 (N_9806,N_9080,N_9354);
xnor U9807 (N_9807,N_9395,N_9259);
and U9808 (N_9808,N_9354,N_9136);
or U9809 (N_9809,N_9257,N_9162);
and U9810 (N_9810,N_9119,N_9069);
xor U9811 (N_9811,N_9222,N_9295);
nor U9812 (N_9812,N_9420,N_9108);
and U9813 (N_9813,N_9226,N_9220);
or U9814 (N_9814,N_9354,N_9279);
xor U9815 (N_9815,N_9420,N_9312);
nor U9816 (N_9816,N_9239,N_9043);
and U9817 (N_9817,N_9415,N_9342);
and U9818 (N_9818,N_9292,N_9029);
and U9819 (N_9819,N_9370,N_9338);
and U9820 (N_9820,N_9181,N_9302);
nand U9821 (N_9821,N_9002,N_9491);
and U9822 (N_9822,N_9448,N_9366);
and U9823 (N_9823,N_9394,N_9008);
or U9824 (N_9824,N_9169,N_9363);
xor U9825 (N_9825,N_9463,N_9459);
or U9826 (N_9826,N_9018,N_9240);
nand U9827 (N_9827,N_9118,N_9142);
nor U9828 (N_9828,N_9064,N_9407);
nor U9829 (N_9829,N_9229,N_9190);
xor U9830 (N_9830,N_9441,N_9484);
nor U9831 (N_9831,N_9047,N_9305);
and U9832 (N_9832,N_9300,N_9223);
nand U9833 (N_9833,N_9196,N_9465);
nand U9834 (N_9834,N_9288,N_9112);
nor U9835 (N_9835,N_9382,N_9340);
nor U9836 (N_9836,N_9219,N_9489);
nand U9837 (N_9837,N_9172,N_9033);
nor U9838 (N_9838,N_9187,N_9286);
nor U9839 (N_9839,N_9131,N_9492);
nor U9840 (N_9840,N_9485,N_9174);
or U9841 (N_9841,N_9119,N_9106);
and U9842 (N_9842,N_9313,N_9000);
nand U9843 (N_9843,N_9220,N_9323);
xnor U9844 (N_9844,N_9190,N_9402);
or U9845 (N_9845,N_9463,N_9292);
xor U9846 (N_9846,N_9401,N_9484);
or U9847 (N_9847,N_9476,N_9139);
and U9848 (N_9848,N_9146,N_9434);
nor U9849 (N_9849,N_9498,N_9414);
nand U9850 (N_9850,N_9259,N_9234);
or U9851 (N_9851,N_9245,N_9133);
nand U9852 (N_9852,N_9080,N_9476);
nand U9853 (N_9853,N_9020,N_9275);
nor U9854 (N_9854,N_9224,N_9389);
or U9855 (N_9855,N_9100,N_9000);
or U9856 (N_9856,N_9466,N_9054);
nor U9857 (N_9857,N_9412,N_9044);
nor U9858 (N_9858,N_9147,N_9329);
nor U9859 (N_9859,N_9442,N_9134);
nand U9860 (N_9860,N_9437,N_9486);
or U9861 (N_9861,N_9356,N_9396);
xnor U9862 (N_9862,N_9335,N_9409);
xnor U9863 (N_9863,N_9182,N_9067);
and U9864 (N_9864,N_9395,N_9352);
nor U9865 (N_9865,N_9230,N_9215);
nand U9866 (N_9866,N_9394,N_9415);
xnor U9867 (N_9867,N_9265,N_9251);
xor U9868 (N_9868,N_9487,N_9056);
nand U9869 (N_9869,N_9407,N_9328);
nor U9870 (N_9870,N_9477,N_9197);
xnor U9871 (N_9871,N_9265,N_9184);
and U9872 (N_9872,N_9085,N_9100);
nand U9873 (N_9873,N_9191,N_9003);
xnor U9874 (N_9874,N_9389,N_9398);
nand U9875 (N_9875,N_9497,N_9387);
xor U9876 (N_9876,N_9051,N_9007);
xor U9877 (N_9877,N_9085,N_9283);
nand U9878 (N_9878,N_9140,N_9342);
nand U9879 (N_9879,N_9135,N_9152);
or U9880 (N_9880,N_9169,N_9408);
and U9881 (N_9881,N_9002,N_9390);
nor U9882 (N_9882,N_9321,N_9289);
nor U9883 (N_9883,N_9058,N_9392);
nor U9884 (N_9884,N_9381,N_9169);
or U9885 (N_9885,N_9311,N_9491);
nand U9886 (N_9886,N_9074,N_9459);
xnor U9887 (N_9887,N_9426,N_9296);
xnor U9888 (N_9888,N_9498,N_9122);
xnor U9889 (N_9889,N_9377,N_9123);
nor U9890 (N_9890,N_9450,N_9185);
and U9891 (N_9891,N_9180,N_9292);
or U9892 (N_9892,N_9358,N_9302);
or U9893 (N_9893,N_9160,N_9329);
or U9894 (N_9894,N_9166,N_9219);
xnor U9895 (N_9895,N_9344,N_9086);
nand U9896 (N_9896,N_9370,N_9132);
nand U9897 (N_9897,N_9328,N_9147);
xor U9898 (N_9898,N_9199,N_9369);
nor U9899 (N_9899,N_9335,N_9015);
or U9900 (N_9900,N_9037,N_9148);
nor U9901 (N_9901,N_9218,N_9432);
or U9902 (N_9902,N_9044,N_9372);
nand U9903 (N_9903,N_9349,N_9213);
xor U9904 (N_9904,N_9007,N_9340);
and U9905 (N_9905,N_9318,N_9467);
and U9906 (N_9906,N_9034,N_9433);
or U9907 (N_9907,N_9451,N_9369);
xor U9908 (N_9908,N_9108,N_9359);
and U9909 (N_9909,N_9115,N_9170);
or U9910 (N_9910,N_9214,N_9408);
and U9911 (N_9911,N_9256,N_9143);
nand U9912 (N_9912,N_9074,N_9207);
or U9913 (N_9913,N_9309,N_9335);
and U9914 (N_9914,N_9407,N_9379);
nor U9915 (N_9915,N_9470,N_9176);
xnor U9916 (N_9916,N_9285,N_9401);
xor U9917 (N_9917,N_9151,N_9176);
or U9918 (N_9918,N_9273,N_9117);
xnor U9919 (N_9919,N_9359,N_9290);
xnor U9920 (N_9920,N_9400,N_9196);
xor U9921 (N_9921,N_9010,N_9283);
xnor U9922 (N_9922,N_9020,N_9368);
and U9923 (N_9923,N_9478,N_9490);
and U9924 (N_9924,N_9234,N_9231);
nand U9925 (N_9925,N_9148,N_9071);
nor U9926 (N_9926,N_9452,N_9007);
and U9927 (N_9927,N_9181,N_9310);
and U9928 (N_9928,N_9274,N_9308);
nor U9929 (N_9929,N_9402,N_9264);
nand U9930 (N_9930,N_9475,N_9196);
or U9931 (N_9931,N_9490,N_9316);
or U9932 (N_9932,N_9305,N_9312);
and U9933 (N_9933,N_9037,N_9292);
nor U9934 (N_9934,N_9161,N_9067);
and U9935 (N_9935,N_9286,N_9236);
and U9936 (N_9936,N_9021,N_9184);
xnor U9937 (N_9937,N_9153,N_9226);
nor U9938 (N_9938,N_9060,N_9408);
nand U9939 (N_9939,N_9406,N_9208);
nor U9940 (N_9940,N_9022,N_9075);
nor U9941 (N_9941,N_9037,N_9352);
or U9942 (N_9942,N_9361,N_9241);
and U9943 (N_9943,N_9041,N_9009);
nand U9944 (N_9944,N_9493,N_9125);
nor U9945 (N_9945,N_9115,N_9117);
nand U9946 (N_9946,N_9232,N_9483);
nand U9947 (N_9947,N_9027,N_9046);
or U9948 (N_9948,N_9395,N_9243);
nand U9949 (N_9949,N_9227,N_9027);
nand U9950 (N_9950,N_9330,N_9087);
nor U9951 (N_9951,N_9022,N_9183);
nand U9952 (N_9952,N_9398,N_9175);
and U9953 (N_9953,N_9282,N_9210);
nand U9954 (N_9954,N_9261,N_9023);
or U9955 (N_9955,N_9337,N_9278);
and U9956 (N_9956,N_9408,N_9242);
nand U9957 (N_9957,N_9031,N_9129);
nand U9958 (N_9958,N_9400,N_9392);
xnor U9959 (N_9959,N_9390,N_9130);
nor U9960 (N_9960,N_9034,N_9175);
xnor U9961 (N_9961,N_9010,N_9027);
nor U9962 (N_9962,N_9202,N_9065);
nand U9963 (N_9963,N_9253,N_9358);
nor U9964 (N_9964,N_9192,N_9374);
and U9965 (N_9965,N_9267,N_9492);
xor U9966 (N_9966,N_9397,N_9337);
xnor U9967 (N_9967,N_9249,N_9130);
or U9968 (N_9968,N_9059,N_9251);
nand U9969 (N_9969,N_9119,N_9433);
nand U9970 (N_9970,N_9330,N_9092);
or U9971 (N_9971,N_9313,N_9335);
nand U9972 (N_9972,N_9322,N_9256);
and U9973 (N_9973,N_9255,N_9082);
nor U9974 (N_9974,N_9272,N_9417);
xor U9975 (N_9975,N_9170,N_9438);
xnor U9976 (N_9976,N_9482,N_9204);
xnor U9977 (N_9977,N_9351,N_9016);
xnor U9978 (N_9978,N_9374,N_9034);
and U9979 (N_9979,N_9365,N_9423);
nor U9980 (N_9980,N_9211,N_9026);
or U9981 (N_9981,N_9198,N_9058);
xor U9982 (N_9982,N_9064,N_9352);
xor U9983 (N_9983,N_9099,N_9424);
and U9984 (N_9984,N_9017,N_9346);
nand U9985 (N_9985,N_9162,N_9391);
nor U9986 (N_9986,N_9100,N_9055);
or U9987 (N_9987,N_9497,N_9403);
and U9988 (N_9988,N_9367,N_9432);
or U9989 (N_9989,N_9089,N_9411);
or U9990 (N_9990,N_9121,N_9152);
xnor U9991 (N_9991,N_9071,N_9076);
nor U9992 (N_9992,N_9283,N_9344);
xnor U9993 (N_9993,N_9367,N_9030);
nor U9994 (N_9994,N_9028,N_9173);
nand U9995 (N_9995,N_9034,N_9323);
xnor U9996 (N_9996,N_9353,N_9405);
xnor U9997 (N_9997,N_9457,N_9265);
nor U9998 (N_9998,N_9383,N_9140);
xnor U9999 (N_9999,N_9489,N_9184);
nand U10000 (N_10000,N_9871,N_9604);
or U10001 (N_10001,N_9898,N_9990);
nand U10002 (N_10002,N_9673,N_9717);
or U10003 (N_10003,N_9869,N_9992);
and U10004 (N_10004,N_9585,N_9667);
nor U10005 (N_10005,N_9998,N_9653);
nor U10006 (N_10006,N_9515,N_9841);
or U10007 (N_10007,N_9605,N_9862);
nor U10008 (N_10008,N_9509,N_9546);
xnor U10009 (N_10009,N_9867,N_9937);
xor U10010 (N_10010,N_9792,N_9510);
and U10011 (N_10011,N_9989,N_9684);
nand U10012 (N_10012,N_9743,N_9544);
or U10013 (N_10013,N_9908,N_9996);
and U10014 (N_10014,N_9583,N_9629);
nor U10015 (N_10015,N_9507,N_9560);
or U10016 (N_10016,N_9789,N_9947);
nand U10017 (N_10017,N_9567,N_9540);
nor U10018 (N_10018,N_9536,N_9534);
nor U10019 (N_10019,N_9819,N_9859);
nand U10020 (N_10020,N_9638,N_9704);
nand U10021 (N_10021,N_9844,N_9550);
xnor U10022 (N_10022,N_9516,N_9801);
xnor U10023 (N_10023,N_9821,N_9942);
or U10024 (N_10024,N_9580,N_9883);
and U10025 (N_10025,N_9590,N_9525);
nand U10026 (N_10026,N_9678,N_9562);
nor U10027 (N_10027,N_9565,N_9770);
nand U10028 (N_10028,N_9838,N_9995);
and U10029 (N_10029,N_9651,N_9827);
or U10030 (N_10030,N_9663,N_9648);
xor U10031 (N_10031,N_9620,N_9596);
or U10032 (N_10032,N_9724,N_9729);
and U10033 (N_10033,N_9705,N_9745);
and U10034 (N_10034,N_9710,N_9785);
nand U10035 (N_10035,N_9985,N_9670);
nor U10036 (N_10036,N_9647,N_9698);
and U10037 (N_10037,N_9689,N_9504);
and U10038 (N_10038,N_9796,N_9781);
nor U10039 (N_10039,N_9601,N_9628);
nor U10040 (N_10040,N_9748,N_9921);
and U10041 (N_10041,N_9674,N_9623);
xnor U10042 (N_10042,N_9617,N_9696);
and U10043 (N_10043,N_9733,N_9640);
or U10044 (N_10044,N_9813,N_9881);
xnor U10045 (N_10045,N_9965,N_9764);
nor U10046 (N_10046,N_9830,N_9706);
xor U10047 (N_10047,N_9870,N_9609);
or U10048 (N_10048,N_9902,N_9794);
nand U10049 (N_10049,N_9750,N_9826);
xnor U10050 (N_10050,N_9784,N_9731);
xor U10051 (N_10051,N_9872,N_9941);
or U10052 (N_10052,N_9740,N_9727);
xor U10053 (N_10053,N_9524,N_9966);
xor U10054 (N_10054,N_9887,N_9688);
xnor U10055 (N_10055,N_9527,N_9660);
and U10056 (N_10056,N_9805,N_9514);
nor U10057 (N_10057,N_9849,N_9914);
xnor U10058 (N_10058,N_9880,N_9650);
xnor U10059 (N_10059,N_9850,N_9878);
and U10060 (N_10060,N_9817,N_9814);
and U10061 (N_10061,N_9642,N_9641);
xor U10062 (N_10062,N_9861,N_9708);
or U10063 (N_10063,N_9954,N_9910);
nor U10064 (N_10064,N_9557,N_9734);
xor U10065 (N_10065,N_9940,N_9918);
nand U10066 (N_10066,N_9882,N_9915);
and U10067 (N_10067,N_9800,N_9926);
nor U10068 (N_10068,N_9588,N_9953);
or U10069 (N_10069,N_9969,N_9759);
nor U10070 (N_10070,N_9503,N_9677);
nand U10071 (N_10071,N_9532,N_9854);
nand U10072 (N_10072,N_9686,N_9665);
and U10073 (N_10073,N_9597,N_9829);
xnor U10074 (N_10074,N_9551,N_9719);
or U10075 (N_10075,N_9807,N_9951);
or U10076 (N_10076,N_9783,N_9751);
nand U10077 (N_10077,N_9886,N_9528);
nor U10078 (N_10078,N_9755,N_9857);
xor U10079 (N_10079,N_9575,N_9948);
xnor U10080 (N_10080,N_9676,N_9701);
or U10081 (N_10081,N_9925,N_9636);
nor U10082 (N_10082,N_9702,N_9936);
nor U10083 (N_10083,N_9797,N_9505);
and U10084 (N_10084,N_9892,N_9522);
and U10085 (N_10085,N_9659,N_9868);
nor U10086 (N_10086,N_9610,N_9891);
or U10087 (N_10087,N_9960,N_9763);
nand U10088 (N_10088,N_9820,N_9711);
nor U10089 (N_10089,N_9737,N_9831);
xor U10090 (N_10090,N_9978,N_9556);
nand U10091 (N_10091,N_9526,N_9888);
nand U10092 (N_10092,N_9833,N_9714);
nor U10093 (N_10093,N_9691,N_9955);
and U10094 (N_10094,N_9832,N_9591);
xnor U10095 (N_10095,N_9626,N_9592);
nand U10096 (N_10096,N_9874,N_9683);
nor U10097 (N_10097,N_9757,N_9928);
nand U10098 (N_10098,N_9811,N_9793);
nor U10099 (N_10099,N_9924,N_9579);
nor U10100 (N_10100,N_9856,N_9900);
nor U10101 (N_10101,N_9720,N_9988);
xor U10102 (N_10102,N_9637,N_9839);
or U10103 (N_10103,N_9541,N_9973);
nand U10104 (N_10104,N_9905,N_9533);
or U10105 (N_10105,N_9549,N_9855);
nand U10106 (N_10106,N_9558,N_9538);
and U10107 (N_10107,N_9961,N_9916);
xor U10108 (N_10108,N_9746,N_9968);
or U10109 (N_10109,N_9958,N_9920);
xor U10110 (N_10110,N_9625,N_9622);
nand U10111 (N_10111,N_9790,N_9952);
or U10112 (N_10112,N_9699,N_9694);
or U10113 (N_10113,N_9788,N_9779);
or U10114 (N_10114,N_9984,N_9912);
and U10115 (N_10115,N_9901,N_9675);
nand U10116 (N_10116,N_9885,N_9631);
nor U10117 (N_10117,N_9837,N_9884);
or U10118 (N_10118,N_9695,N_9846);
nand U10119 (N_10119,N_9842,N_9767);
or U10120 (N_10120,N_9923,N_9661);
nor U10121 (N_10121,N_9501,N_9741);
nor U10122 (N_10122,N_9964,N_9762);
and U10123 (N_10123,N_9634,N_9722);
nand U10124 (N_10124,N_9749,N_9753);
nor U10125 (N_10125,N_9975,N_9569);
and U10126 (N_10126,N_9709,N_9654);
and U10127 (N_10127,N_9851,N_9530);
nor U10128 (N_10128,N_9899,N_9555);
nand U10129 (N_10129,N_9618,N_9598);
and U10130 (N_10130,N_9806,N_9639);
and U10131 (N_10131,N_9697,N_9679);
and U10132 (N_10132,N_9935,N_9715);
nand U10133 (N_10133,N_9627,N_9777);
nand U10134 (N_10134,N_9502,N_9982);
nand U10135 (N_10135,N_9758,N_9561);
and U10136 (N_10136,N_9950,N_9782);
and U10137 (N_10137,N_9977,N_9582);
nor U10138 (N_10138,N_9644,N_9687);
nand U10139 (N_10139,N_9766,N_9619);
nand U10140 (N_10140,N_9939,N_9840);
or U10141 (N_10141,N_9879,N_9774);
xnor U10142 (N_10142,N_9692,N_9513);
nor U10143 (N_10143,N_9865,N_9547);
or U10144 (N_10144,N_9621,N_9570);
xor U10145 (N_10145,N_9922,N_9907);
nor U10146 (N_10146,N_9930,N_9738);
nor U10147 (N_10147,N_9962,N_9615);
nor U10148 (N_10148,N_9539,N_9822);
and U10149 (N_10149,N_9852,N_9890);
or U10150 (N_10150,N_9776,N_9836);
xnor U10151 (N_10151,N_9906,N_9559);
and U10152 (N_10152,N_9889,N_9716);
and U10153 (N_10153,N_9537,N_9594);
nor U10154 (N_10154,N_9944,N_9681);
xnor U10155 (N_10155,N_9835,N_9587);
and U10156 (N_10156,N_9574,N_9736);
xnor U10157 (N_10157,N_9703,N_9742);
xor U10158 (N_10158,N_9972,N_9664);
nand U10159 (N_10159,N_9818,N_9876);
nor U10160 (N_10160,N_9730,N_9595);
nor U10161 (N_10161,N_9863,N_9860);
nor U10162 (N_10162,N_9877,N_9643);
or U10163 (N_10163,N_9894,N_9873);
xnor U10164 (N_10164,N_9542,N_9608);
nor U10165 (N_10165,N_9512,N_9991);
nand U10166 (N_10166,N_9957,N_9671);
xnor U10167 (N_10167,N_9816,N_9929);
and U10168 (N_10168,N_9531,N_9732);
and U10169 (N_10169,N_9932,N_9721);
nor U10170 (N_10170,N_9798,N_9812);
nor U10171 (N_10171,N_9529,N_9553);
and U10172 (N_10172,N_9739,N_9848);
or U10173 (N_10173,N_9645,N_9787);
and U10174 (N_10174,N_9646,N_9786);
nor U10175 (N_10175,N_9949,N_9586);
nor U10176 (N_10176,N_9564,N_9974);
and U10177 (N_10177,N_9672,N_9927);
nand U10178 (N_10178,N_9548,N_9934);
and U10179 (N_10179,N_9971,N_9834);
nand U10180 (N_10180,N_9919,N_9690);
xor U10181 (N_10181,N_9773,N_9999);
and U10182 (N_10182,N_9632,N_9726);
xnor U10183 (N_10183,N_9795,N_9810);
and U10184 (N_10184,N_9771,N_9566);
nor U10185 (N_10185,N_9896,N_9804);
nor U10186 (N_10186,N_9700,N_9980);
and U10187 (N_10187,N_9723,N_9607);
and U10188 (N_10188,N_9780,N_9535);
xor U10189 (N_10189,N_9603,N_9772);
nand U10190 (N_10190,N_9847,N_9571);
nand U10191 (N_10191,N_9668,N_9769);
xor U10192 (N_10192,N_9931,N_9602);
nand U10193 (N_10193,N_9843,N_9903);
or U10194 (N_10194,N_9511,N_9768);
or U10195 (N_10195,N_9573,N_9652);
and U10196 (N_10196,N_9523,N_9600);
or U10197 (N_10197,N_9828,N_9599);
and U10198 (N_10198,N_9728,N_9589);
and U10199 (N_10199,N_9893,N_9845);
nand U10200 (N_10200,N_9987,N_9669);
and U10201 (N_10201,N_9864,N_9635);
nor U10202 (N_10202,N_9754,N_9520);
or U10203 (N_10203,N_9803,N_9979);
and U10204 (N_10204,N_9760,N_9508);
and U10205 (N_10205,N_9997,N_9761);
and U10206 (N_10206,N_9959,N_9713);
nor U10207 (N_10207,N_9718,N_9680);
or U10208 (N_10208,N_9707,N_9858);
and U10209 (N_10209,N_9614,N_9943);
xor U10210 (N_10210,N_9981,N_9866);
or U10211 (N_10211,N_9506,N_9606);
xor U10212 (N_10212,N_9976,N_9593);
nor U10213 (N_10213,N_9649,N_9808);
nand U10214 (N_10214,N_9578,N_9744);
nand U10215 (N_10215,N_9823,N_9577);
nand U10216 (N_10216,N_9983,N_9518);
nor U10217 (N_10217,N_9735,N_9809);
or U10218 (N_10218,N_9956,N_9909);
nand U10219 (N_10219,N_9612,N_9897);
nand U10220 (N_10220,N_9682,N_9917);
or U10221 (N_10221,N_9895,N_9775);
nor U10222 (N_10222,N_9613,N_9747);
nand U10223 (N_10223,N_9986,N_9552);
or U10224 (N_10224,N_9911,N_9824);
nor U10225 (N_10225,N_9967,N_9500);
nor U10226 (N_10226,N_9611,N_9685);
nand U10227 (N_10227,N_9802,N_9563);
and U10228 (N_10228,N_9799,N_9825);
nand U10229 (N_10229,N_9904,N_9756);
and U10230 (N_10230,N_9970,N_9875);
or U10231 (N_10231,N_9616,N_9791);
nor U10232 (N_10232,N_9656,N_9554);
or U10233 (N_10233,N_9994,N_9521);
nand U10234 (N_10234,N_9752,N_9543);
and U10235 (N_10235,N_9963,N_9517);
or U10236 (N_10236,N_9765,N_9933);
and U10237 (N_10237,N_9913,N_9712);
xnor U10238 (N_10238,N_9853,N_9938);
xor U10239 (N_10239,N_9581,N_9624);
nor U10240 (N_10240,N_9584,N_9657);
xor U10241 (N_10241,N_9946,N_9945);
and U10242 (N_10242,N_9519,N_9545);
and U10243 (N_10243,N_9655,N_9568);
nor U10244 (N_10244,N_9658,N_9630);
or U10245 (N_10245,N_9666,N_9725);
and U10246 (N_10246,N_9993,N_9633);
xor U10247 (N_10247,N_9693,N_9778);
or U10248 (N_10248,N_9572,N_9815);
xnor U10249 (N_10249,N_9662,N_9576);
and U10250 (N_10250,N_9613,N_9584);
or U10251 (N_10251,N_9667,N_9745);
nand U10252 (N_10252,N_9634,N_9588);
and U10253 (N_10253,N_9704,N_9622);
or U10254 (N_10254,N_9690,N_9682);
and U10255 (N_10255,N_9567,N_9908);
xnor U10256 (N_10256,N_9835,N_9768);
nor U10257 (N_10257,N_9927,N_9823);
or U10258 (N_10258,N_9980,N_9624);
and U10259 (N_10259,N_9717,N_9584);
nand U10260 (N_10260,N_9808,N_9892);
or U10261 (N_10261,N_9621,N_9895);
nor U10262 (N_10262,N_9505,N_9723);
nor U10263 (N_10263,N_9955,N_9996);
nand U10264 (N_10264,N_9605,N_9565);
and U10265 (N_10265,N_9995,N_9942);
nand U10266 (N_10266,N_9630,N_9606);
xor U10267 (N_10267,N_9629,N_9984);
nand U10268 (N_10268,N_9856,N_9631);
and U10269 (N_10269,N_9590,N_9604);
nand U10270 (N_10270,N_9519,N_9975);
or U10271 (N_10271,N_9744,N_9521);
and U10272 (N_10272,N_9974,N_9936);
nand U10273 (N_10273,N_9801,N_9844);
nand U10274 (N_10274,N_9799,N_9522);
xor U10275 (N_10275,N_9721,N_9996);
or U10276 (N_10276,N_9508,N_9854);
or U10277 (N_10277,N_9766,N_9632);
nand U10278 (N_10278,N_9617,N_9781);
nand U10279 (N_10279,N_9522,N_9847);
nor U10280 (N_10280,N_9562,N_9585);
or U10281 (N_10281,N_9985,N_9719);
nand U10282 (N_10282,N_9747,N_9551);
or U10283 (N_10283,N_9573,N_9532);
or U10284 (N_10284,N_9874,N_9625);
nor U10285 (N_10285,N_9731,N_9825);
or U10286 (N_10286,N_9862,N_9749);
or U10287 (N_10287,N_9750,N_9875);
nand U10288 (N_10288,N_9866,N_9902);
or U10289 (N_10289,N_9614,N_9536);
nor U10290 (N_10290,N_9582,N_9905);
xor U10291 (N_10291,N_9940,N_9727);
and U10292 (N_10292,N_9616,N_9899);
and U10293 (N_10293,N_9645,N_9883);
nor U10294 (N_10294,N_9868,N_9690);
nor U10295 (N_10295,N_9812,N_9722);
nor U10296 (N_10296,N_9961,N_9685);
nand U10297 (N_10297,N_9697,N_9560);
and U10298 (N_10298,N_9960,N_9620);
or U10299 (N_10299,N_9615,N_9891);
nand U10300 (N_10300,N_9723,N_9916);
nand U10301 (N_10301,N_9884,N_9814);
or U10302 (N_10302,N_9517,N_9787);
and U10303 (N_10303,N_9673,N_9957);
nand U10304 (N_10304,N_9797,N_9687);
nand U10305 (N_10305,N_9542,N_9892);
nor U10306 (N_10306,N_9856,N_9667);
xor U10307 (N_10307,N_9908,N_9783);
and U10308 (N_10308,N_9564,N_9649);
and U10309 (N_10309,N_9610,N_9851);
nand U10310 (N_10310,N_9640,N_9966);
and U10311 (N_10311,N_9839,N_9878);
nor U10312 (N_10312,N_9912,N_9952);
xor U10313 (N_10313,N_9542,N_9958);
and U10314 (N_10314,N_9771,N_9880);
nor U10315 (N_10315,N_9594,N_9506);
and U10316 (N_10316,N_9541,N_9876);
and U10317 (N_10317,N_9990,N_9932);
nand U10318 (N_10318,N_9631,N_9825);
and U10319 (N_10319,N_9573,N_9742);
and U10320 (N_10320,N_9620,N_9704);
nand U10321 (N_10321,N_9511,N_9836);
nor U10322 (N_10322,N_9915,N_9542);
xnor U10323 (N_10323,N_9751,N_9913);
xnor U10324 (N_10324,N_9964,N_9996);
or U10325 (N_10325,N_9577,N_9955);
or U10326 (N_10326,N_9781,N_9678);
nand U10327 (N_10327,N_9677,N_9903);
and U10328 (N_10328,N_9815,N_9883);
and U10329 (N_10329,N_9716,N_9984);
or U10330 (N_10330,N_9900,N_9917);
nand U10331 (N_10331,N_9617,N_9975);
xor U10332 (N_10332,N_9734,N_9545);
nor U10333 (N_10333,N_9705,N_9861);
or U10334 (N_10334,N_9884,N_9905);
nand U10335 (N_10335,N_9535,N_9603);
nor U10336 (N_10336,N_9526,N_9947);
or U10337 (N_10337,N_9535,N_9708);
nor U10338 (N_10338,N_9671,N_9837);
nor U10339 (N_10339,N_9654,N_9921);
and U10340 (N_10340,N_9839,N_9971);
or U10341 (N_10341,N_9584,N_9570);
and U10342 (N_10342,N_9945,N_9750);
and U10343 (N_10343,N_9562,N_9667);
and U10344 (N_10344,N_9627,N_9704);
or U10345 (N_10345,N_9786,N_9623);
or U10346 (N_10346,N_9539,N_9764);
nand U10347 (N_10347,N_9791,N_9718);
nor U10348 (N_10348,N_9693,N_9837);
and U10349 (N_10349,N_9957,N_9709);
or U10350 (N_10350,N_9643,N_9849);
nand U10351 (N_10351,N_9837,N_9989);
or U10352 (N_10352,N_9837,N_9992);
nor U10353 (N_10353,N_9716,N_9578);
nand U10354 (N_10354,N_9874,N_9689);
and U10355 (N_10355,N_9534,N_9518);
or U10356 (N_10356,N_9694,N_9888);
and U10357 (N_10357,N_9723,N_9875);
or U10358 (N_10358,N_9936,N_9516);
nand U10359 (N_10359,N_9697,N_9711);
nor U10360 (N_10360,N_9706,N_9663);
nor U10361 (N_10361,N_9842,N_9716);
or U10362 (N_10362,N_9514,N_9528);
and U10363 (N_10363,N_9871,N_9983);
xnor U10364 (N_10364,N_9800,N_9842);
or U10365 (N_10365,N_9521,N_9705);
nand U10366 (N_10366,N_9724,N_9917);
and U10367 (N_10367,N_9976,N_9610);
xnor U10368 (N_10368,N_9586,N_9982);
xor U10369 (N_10369,N_9687,N_9855);
and U10370 (N_10370,N_9707,N_9819);
or U10371 (N_10371,N_9620,N_9889);
xor U10372 (N_10372,N_9862,N_9908);
xor U10373 (N_10373,N_9824,N_9600);
nand U10374 (N_10374,N_9508,N_9510);
xor U10375 (N_10375,N_9983,N_9875);
nor U10376 (N_10376,N_9544,N_9701);
or U10377 (N_10377,N_9715,N_9828);
xor U10378 (N_10378,N_9840,N_9837);
and U10379 (N_10379,N_9969,N_9565);
or U10380 (N_10380,N_9886,N_9671);
and U10381 (N_10381,N_9944,N_9675);
or U10382 (N_10382,N_9695,N_9670);
or U10383 (N_10383,N_9728,N_9626);
or U10384 (N_10384,N_9717,N_9821);
or U10385 (N_10385,N_9755,N_9849);
or U10386 (N_10386,N_9538,N_9592);
nand U10387 (N_10387,N_9848,N_9966);
and U10388 (N_10388,N_9791,N_9945);
nor U10389 (N_10389,N_9866,N_9898);
and U10390 (N_10390,N_9637,N_9707);
nand U10391 (N_10391,N_9935,N_9635);
and U10392 (N_10392,N_9973,N_9943);
and U10393 (N_10393,N_9533,N_9830);
nor U10394 (N_10394,N_9607,N_9926);
or U10395 (N_10395,N_9827,N_9578);
and U10396 (N_10396,N_9852,N_9774);
or U10397 (N_10397,N_9871,N_9512);
and U10398 (N_10398,N_9908,N_9669);
nand U10399 (N_10399,N_9524,N_9528);
xnor U10400 (N_10400,N_9944,N_9867);
nand U10401 (N_10401,N_9593,N_9654);
xnor U10402 (N_10402,N_9957,N_9793);
xor U10403 (N_10403,N_9991,N_9504);
nand U10404 (N_10404,N_9785,N_9762);
nand U10405 (N_10405,N_9558,N_9986);
nor U10406 (N_10406,N_9611,N_9911);
nand U10407 (N_10407,N_9607,N_9737);
nand U10408 (N_10408,N_9787,N_9572);
nor U10409 (N_10409,N_9532,N_9949);
and U10410 (N_10410,N_9626,N_9831);
and U10411 (N_10411,N_9700,N_9879);
xor U10412 (N_10412,N_9673,N_9891);
nand U10413 (N_10413,N_9766,N_9773);
xnor U10414 (N_10414,N_9782,N_9619);
or U10415 (N_10415,N_9757,N_9851);
xnor U10416 (N_10416,N_9648,N_9624);
or U10417 (N_10417,N_9944,N_9866);
or U10418 (N_10418,N_9749,N_9871);
nor U10419 (N_10419,N_9531,N_9695);
nand U10420 (N_10420,N_9858,N_9997);
xnor U10421 (N_10421,N_9635,N_9704);
xnor U10422 (N_10422,N_9708,N_9695);
nor U10423 (N_10423,N_9724,N_9854);
xnor U10424 (N_10424,N_9544,N_9666);
or U10425 (N_10425,N_9931,N_9789);
or U10426 (N_10426,N_9855,N_9904);
xor U10427 (N_10427,N_9820,N_9792);
nor U10428 (N_10428,N_9862,N_9942);
and U10429 (N_10429,N_9537,N_9623);
nor U10430 (N_10430,N_9821,N_9774);
and U10431 (N_10431,N_9843,N_9722);
nor U10432 (N_10432,N_9704,N_9727);
nand U10433 (N_10433,N_9875,N_9994);
nand U10434 (N_10434,N_9517,N_9791);
nand U10435 (N_10435,N_9814,N_9765);
xnor U10436 (N_10436,N_9666,N_9703);
nor U10437 (N_10437,N_9703,N_9978);
and U10438 (N_10438,N_9877,N_9853);
or U10439 (N_10439,N_9658,N_9561);
nor U10440 (N_10440,N_9857,N_9884);
and U10441 (N_10441,N_9935,N_9582);
nor U10442 (N_10442,N_9865,N_9548);
nor U10443 (N_10443,N_9869,N_9577);
nand U10444 (N_10444,N_9729,N_9854);
xnor U10445 (N_10445,N_9664,N_9611);
and U10446 (N_10446,N_9579,N_9551);
or U10447 (N_10447,N_9853,N_9707);
nand U10448 (N_10448,N_9510,N_9661);
nor U10449 (N_10449,N_9685,N_9655);
and U10450 (N_10450,N_9936,N_9876);
nor U10451 (N_10451,N_9590,N_9663);
and U10452 (N_10452,N_9781,N_9534);
nand U10453 (N_10453,N_9778,N_9985);
xnor U10454 (N_10454,N_9659,N_9830);
nor U10455 (N_10455,N_9767,N_9646);
nor U10456 (N_10456,N_9510,N_9683);
and U10457 (N_10457,N_9522,N_9825);
xor U10458 (N_10458,N_9891,N_9620);
xor U10459 (N_10459,N_9515,N_9671);
nor U10460 (N_10460,N_9962,N_9712);
nand U10461 (N_10461,N_9757,N_9989);
and U10462 (N_10462,N_9814,N_9692);
nand U10463 (N_10463,N_9558,N_9726);
nor U10464 (N_10464,N_9871,N_9600);
and U10465 (N_10465,N_9911,N_9917);
nor U10466 (N_10466,N_9567,N_9826);
and U10467 (N_10467,N_9958,N_9791);
nand U10468 (N_10468,N_9538,N_9554);
nand U10469 (N_10469,N_9797,N_9575);
nand U10470 (N_10470,N_9586,N_9553);
nor U10471 (N_10471,N_9711,N_9901);
nor U10472 (N_10472,N_9920,N_9922);
or U10473 (N_10473,N_9592,N_9584);
or U10474 (N_10474,N_9955,N_9790);
nand U10475 (N_10475,N_9604,N_9515);
nor U10476 (N_10476,N_9872,N_9712);
nor U10477 (N_10477,N_9947,N_9657);
nand U10478 (N_10478,N_9994,N_9983);
or U10479 (N_10479,N_9689,N_9594);
or U10480 (N_10480,N_9937,N_9693);
or U10481 (N_10481,N_9566,N_9969);
and U10482 (N_10482,N_9781,N_9600);
or U10483 (N_10483,N_9554,N_9642);
xnor U10484 (N_10484,N_9795,N_9783);
or U10485 (N_10485,N_9873,N_9718);
or U10486 (N_10486,N_9863,N_9831);
or U10487 (N_10487,N_9795,N_9817);
nand U10488 (N_10488,N_9827,N_9537);
and U10489 (N_10489,N_9697,N_9587);
xor U10490 (N_10490,N_9585,N_9619);
or U10491 (N_10491,N_9624,N_9599);
xnor U10492 (N_10492,N_9715,N_9946);
xor U10493 (N_10493,N_9641,N_9897);
nand U10494 (N_10494,N_9948,N_9588);
nor U10495 (N_10495,N_9505,N_9585);
xor U10496 (N_10496,N_9902,N_9731);
nand U10497 (N_10497,N_9792,N_9694);
xnor U10498 (N_10498,N_9802,N_9863);
nor U10499 (N_10499,N_9796,N_9932);
or U10500 (N_10500,N_10398,N_10180);
or U10501 (N_10501,N_10041,N_10172);
and U10502 (N_10502,N_10390,N_10472);
and U10503 (N_10503,N_10017,N_10415);
xor U10504 (N_10504,N_10067,N_10037);
or U10505 (N_10505,N_10346,N_10272);
nor U10506 (N_10506,N_10466,N_10051);
xnor U10507 (N_10507,N_10444,N_10433);
nand U10508 (N_10508,N_10064,N_10489);
xnor U10509 (N_10509,N_10100,N_10093);
or U10510 (N_10510,N_10063,N_10341);
and U10511 (N_10511,N_10487,N_10254);
xnor U10512 (N_10512,N_10265,N_10068);
or U10513 (N_10513,N_10091,N_10404);
or U10514 (N_10514,N_10192,N_10416);
or U10515 (N_10515,N_10476,N_10214);
nor U10516 (N_10516,N_10130,N_10053);
nand U10517 (N_10517,N_10249,N_10021);
xnor U10518 (N_10518,N_10028,N_10434);
nor U10519 (N_10519,N_10426,N_10245);
xor U10520 (N_10520,N_10428,N_10105);
and U10521 (N_10521,N_10137,N_10314);
and U10522 (N_10522,N_10166,N_10473);
xnor U10523 (N_10523,N_10417,N_10394);
and U10524 (N_10524,N_10084,N_10264);
xnor U10525 (N_10525,N_10389,N_10150);
xor U10526 (N_10526,N_10116,N_10221);
nand U10527 (N_10527,N_10162,N_10218);
nand U10528 (N_10528,N_10143,N_10169);
nand U10529 (N_10529,N_10370,N_10108);
nand U10530 (N_10530,N_10261,N_10047);
nor U10531 (N_10531,N_10383,N_10029);
and U10532 (N_10532,N_10075,N_10361);
nor U10533 (N_10533,N_10322,N_10027);
nor U10534 (N_10534,N_10200,N_10234);
xor U10535 (N_10535,N_10419,N_10395);
and U10536 (N_10536,N_10163,N_10277);
or U10537 (N_10537,N_10311,N_10279);
or U10538 (N_10538,N_10193,N_10388);
or U10539 (N_10539,N_10276,N_10345);
xnor U10540 (N_10540,N_10482,N_10152);
and U10541 (N_10541,N_10464,N_10182);
nand U10542 (N_10542,N_10004,N_10313);
nor U10543 (N_10543,N_10158,N_10074);
and U10544 (N_10544,N_10055,N_10160);
and U10545 (N_10545,N_10363,N_10088);
xor U10546 (N_10546,N_10283,N_10439);
nand U10547 (N_10547,N_10220,N_10478);
and U10548 (N_10548,N_10039,N_10087);
and U10549 (N_10549,N_10046,N_10140);
and U10550 (N_10550,N_10127,N_10251);
or U10551 (N_10551,N_10080,N_10229);
nand U10552 (N_10552,N_10364,N_10256);
nand U10553 (N_10553,N_10461,N_10362);
and U10554 (N_10554,N_10292,N_10131);
and U10555 (N_10555,N_10386,N_10176);
nand U10556 (N_10556,N_10173,N_10114);
nor U10557 (N_10557,N_10151,N_10452);
and U10558 (N_10558,N_10358,N_10441);
nor U10559 (N_10559,N_10297,N_10414);
or U10560 (N_10560,N_10379,N_10278);
nand U10561 (N_10561,N_10209,N_10223);
nand U10562 (N_10562,N_10164,N_10081);
or U10563 (N_10563,N_10174,N_10185);
nand U10564 (N_10564,N_10418,N_10125);
nand U10565 (N_10565,N_10121,N_10274);
or U10566 (N_10566,N_10486,N_10134);
nand U10567 (N_10567,N_10050,N_10492);
or U10568 (N_10568,N_10213,N_10204);
nor U10569 (N_10569,N_10456,N_10094);
or U10570 (N_10570,N_10212,N_10157);
nor U10571 (N_10571,N_10305,N_10230);
and U10572 (N_10572,N_10049,N_10436);
xor U10573 (N_10573,N_10083,N_10432);
xnor U10574 (N_10574,N_10449,N_10138);
or U10575 (N_10575,N_10145,N_10246);
nand U10576 (N_10576,N_10061,N_10179);
nand U10577 (N_10577,N_10167,N_10040);
or U10578 (N_10578,N_10126,N_10253);
or U10579 (N_10579,N_10186,N_10302);
and U10580 (N_10580,N_10202,N_10147);
xor U10581 (N_10581,N_10109,N_10219);
nor U10582 (N_10582,N_10000,N_10260);
and U10583 (N_10583,N_10409,N_10488);
nor U10584 (N_10584,N_10119,N_10215);
nand U10585 (N_10585,N_10371,N_10038);
xnor U10586 (N_10586,N_10071,N_10224);
xor U10587 (N_10587,N_10124,N_10453);
and U10588 (N_10588,N_10287,N_10233);
xnor U10589 (N_10589,N_10216,N_10319);
or U10590 (N_10590,N_10378,N_10353);
nor U10591 (N_10591,N_10340,N_10024);
and U10592 (N_10592,N_10285,N_10303);
nand U10593 (N_10593,N_10066,N_10493);
nand U10594 (N_10594,N_10092,N_10210);
nor U10595 (N_10595,N_10400,N_10380);
nand U10596 (N_10596,N_10070,N_10026);
and U10597 (N_10597,N_10065,N_10442);
or U10598 (N_10598,N_10463,N_10023);
or U10599 (N_10599,N_10307,N_10333);
nor U10600 (N_10600,N_10351,N_10184);
nor U10601 (N_10601,N_10443,N_10168);
nand U10602 (N_10602,N_10339,N_10144);
nand U10603 (N_10603,N_10481,N_10368);
nor U10604 (N_10604,N_10106,N_10490);
or U10605 (N_10605,N_10183,N_10191);
nor U10606 (N_10606,N_10240,N_10465);
xor U10607 (N_10607,N_10112,N_10329);
or U10608 (N_10608,N_10032,N_10089);
or U10609 (N_10609,N_10247,N_10077);
xor U10610 (N_10610,N_10429,N_10460);
xnor U10611 (N_10611,N_10446,N_10290);
or U10612 (N_10612,N_10033,N_10455);
nor U10613 (N_10613,N_10048,N_10448);
nand U10614 (N_10614,N_10325,N_10059);
or U10615 (N_10615,N_10289,N_10052);
xor U10616 (N_10616,N_10284,N_10308);
nand U10617 (N_10617,N_10072,N_10217);
xor U10618 (N_10618,N_10142,N_10248);
nor U10619 (N_10619,N_10365,N_10331);
nor U10620 (N_10620,N_10069,N_10205);
xor U10621 (N_10621,N_10499,N_10043);
xor U10622 (N_10622,N_10420,N_10470);
and U10623 (N_10623,N_10451,N_10117);
nor U10624 (N_10624,N_10111,N_10252);
or U10625 (N_10625,N_10236,N_10467);
xnor U10626 (N_10626,N_10425,N_10471);
nor U10627 (N_10627,N_10270,N_10058);
nand U10628 (N_10628,N_10073,N_10014);
and U10629 (N_10629,N_10375,N_10045);
and U10630 (N_10630,N_10267,N_10475);
nor U10631 (N_10631,N_10299,N_10301);
xnor U10632 (N_10632,N_10201,N_10239);
nand U10633 (N_10633,N_10086,N_10360);
nand U10634 (N_10634,N_10104,N_10129);
or U10635 (N_10635,N_10403,N_10320);
nand U10636 (N_10636,N_10232,N_10231);
and U10637 (N_10637,N_10318,N_10397);
nor U10638 (N_10638,N_10008,N_10025);
or U10639 (N_10639,N_10009,N_10005);
or U10640 (N_10640,N_10382,N_10042);
xnor U10641 (N_10641,N_10194,N_10141);
and U10642 (N_10642,N_10298,N_10165);
or U10643 (N_10643,N_10110,N_10396);
or U10644 (N_10644,N_10355,N_10016);
nor U10645 (N_10645,N_10374,N_10323);
nor U10646 (N_10646,N_10342,N_10095);
nor U10647 (N_10647,N_10413,N_10227);
and U10648 (N_10648,N_10149,N_10096);
nand U10649 (N_10649,N_10334,N_10002);
nor U10650 (N_10650,N_10243,N_10120);
or U10651 (N_10651,N_10424,N_10352);
nor U10652 (N_10652,N_10139,N_10238);
nor U10653 (N_10653,N_10310,N_10188);
and U10654 (N_10654,N_10317,N_10410);
nor U10655 (N_10655,N_10458,N_10427);
xnor U10656 (N_10656,N_10031,N_10187);
and U10657 (N_10657,N_10135,N_10161);
nand U10658 (N_10658,N_10196,N_10288);
and U10659 (N_10659,N_10468,N_10263);
or U10660 (N_10660,N_10480,N_10373);
or U10661 (N_10661,N_10459,N_10338);
xor U10662 (N_10662,N_10381,N_10423);
nor U10663 (N_10663,N_10122,N_10469);
nand U10664 (N_10664,N_10136,N_10079);
and U10665 (N_10665,N_10401,N_10402);
and U10666 (N_10666,N_10491,N_10098);
xor U10667 (N_10667,N_10155,N_10326);
nor U10668 (N_10668,N_10359,N_10372);
or U10669 (N_10669,N_10132,N_10437);
nor U10670 (N_10670,N_10327,N_10477);
xor U10671 (N_10671,N_10019,N_10078);
nor U10672 (N_10672,N_10101,N_10022);
or U10673 (N_10673,N_10348,N_10153);
xnor U10674 (N_10674,N_10203,N_10128);
and U10675 (N_10675,N_10268,N_10035);
and U10676 (N_10676,N_10332,N_10343);
nand U10677 (N_10677,N_10496,N_10123);
xnor U10678 (N_10678,N_10495,N_10387);
xor U10679 (N_10679,N_10498,N_10408);
nor U10680 (N_10680,N_10321,N_10337);
and U10681 (N_10681,N_10330,N_10244);
or U10682 (N_10682,N_10350,N_10060);
or U10683 (N_10683,N_10349,N_10367);
nand U10684 (N_10684,N_10421,N_10377);
xor U10685 (N_10685,N_10007,N_10271);
nand U10686 (N_10686,N_10103,N_10454);
xnor U10687 (N_10687,N_10090,N_10296);
xnor U10688 (N_10688,N_10097,N_10181);
or U10689 (N_10689,N_10175,N_10336);
nand U10690 (N_10690,N_10281,N_10282);
or U10691 (N_10691,N_10430,N_10309);
nand U10692 (N_10692,N_10391,N_10286);
nand U10693 (N_10693,N_10479,N_10300);
and U10694 (N_10694,N_10294,N_10189);
nand U10695 (N_10695,N_10056,N_10054);
xnor U10696 (N_10696,N_10324,N_10034);
or U10697 (N_10697,N_10369,N_10003);
xor U10698 (N_10698,N_10412,N_10497);
and U10699 (N_10699,N_10484,N_10177);
or U10700 (N_10700,N_10356,N_10291);
xnor U10701 (N_10701,N_10036,N_10393);
nand U10702 (N_10702,N_10347,N_10405);
and U10703 (N_10703,N_10118,N_10206);
nand U10704 (N_10704,N_10199,N_10197);
xnor U10705 (N_10705,N_10146,N_10198);
and U10706 (N_10706,N_10485,N_10159);
nor U10707 (N_10707,N_10392,N_10411);
nand U10708 (N_10708,N_10357,N_10013);
xor U10709 (N_10709,N_10113,N_10328);
xnor U10710 (N_10710,N_10315,N_10269);
xor U10711 (N_10711,N_10241,N_10250);
or U10712 (N_10712,N_10222,N_10450);
nor U10713 (N_10713,N_10435,N_10259);
nor U10714 (N_10714,N_10102,N_10440);
nor U10715 (N_10715,N_10447,N_10462);
xnor U10716 (N_10716,N_10407,N_10438);
xnor U10717 (N_10717,N_10266,N_10316);
or U10718 (N_10718,N_10406,N_10306);
nand U10719 (N_10719,N_10242,N_10006);
nand U10720 (N_10720,N_10483,N_10190);
and U10721 (N_10721,N_10376,N_10255);
nor U10722 (N_10722,N_10422,N_10258);
nor U10723 (N_10723,N_10012,N_10085);
xor U10724 (N_10724,N_10170,N_10366);
or U10725 (N_10725,N_10445,N_10099);
and U10726 (N_10726,N_10257,N_10156);
and U10727 (N_10727,N_10457,N_10207);
nand U10728 (N_10728,N_10133,N_10082);
and U10729 (N_10729,N_10280,N_10211);
or U10730 (N_10730,N_10107,N_10384);
or U10731 (N_10731,N_10262,N_10010);
xor U10732 (N_10732,N_10171,N_10154);
nand U10733 (N_10733,N_10273,N_10431);
or U10734 (N_10734,N_10020,N_10335);
and U10735 (N_10735,N_10385,N_10354);
nor U10736 (N_10736,N_10030,N_10293);
and U10737 (N_10737,N_10062,N_10474);
xor U10738 (N_10738,N_10076,N_10225);
or U10739 (N_10739,N_10226,N_10237);
nand U10740 (N_10740,N_10148,N_10011);
or U10741 (N_10741,N_10195,N_10057);
nor U10742 (N_10742,N_10399,N_10178);
xnor U10743 (N_10743,N_10295,N_10304);
xnor U10744 (N_10744,N_10018,N_10312);
nor U10745 (N_10745,N_10235,N_10275);
nand U10746 (N_10746,N_10344,N_10015);
xnor U10747 (N_10747,N_10115,N_10208);
nor U10748 (N_10748,N_10044,N_10228);
or U10749 (N_10749,N_10494,N_10001);
or U10750 (N_10750,N_10151,N_10008);
xnor U10751 (N_10751,N_10499,N_10289);
or U10752 (N_10752,N_10017,N_10255);
and U10753 (N_10753,N_10392,N_10408);
nand U10754 (N_10754,N_10134,N_10057);
or U10755 (N_10755,N_10138,N_10252);
and U10756 (N_10756,N_10282,N_10343);
and U10757 (N_10757,N_10030,N_10333);
nand U10758 (N_10758,N_10468,N_10416);
nor U10759 (N_10759,N_10271,N_10087);
nor U10760 (N_10760,N_10010,N_10326);
xor U10761 (N_10761,N_10320,N_10137);
xor U10762 (N_10762,N_10109,N_10077);
xor U10763 (N_10763,N_10345,N_10166);
nand U10764 (N_10764,N_10091,N_10438);
nor U10765 (N_10765,N_10059,N_10056);
xnor U10766 (N_10766,N_10374,N_10465);
nor U10767 (N_10767,N_10384,N_10188);
and U10768 (N_10768,N_10297,N_10487);
and U10769 (N_10769,N_10282,N_10390);
xor U10770 (N_10770,N_10134,N_10086);
nand U10771 (N_10771,N_10347,N_10480);
nor U10772 (N_10772,N_10119,N_10350);
nor U10773 (N_10773,N_10396,N_10370);
nand U10774 (N_10774,N_10378,N_10323);
xnor U10775 (N_10775,N_10196,N_10074);
xor U10776 (N_10776,N_10484,N_10023);
xor U10777 (N_10777,N_10214,N_10239);
xnor U10778 (N_10778,N_10277,N_10286);
and U10779 (N_10779,N_10393,N_10494);
or U10780 (N_10780,N_10175,N_10482);
xnor U10781 (N_10781,N_10124,N_10155);
nor U10782 (N_10782,N_10279,N_10032);
nor U10783 (N_10783,N_10309,N_10109);
nand U10784 (N_10784,N_10498,N_10198);
nor U10785 (N_10785,N_10401,N_10329);
or U10786 (N_10786,N_10225,N_10350);
or U10787 (N_10787,N_10404,N_10202);
and U10788 (N_10788,N_10484,N_10048);
nor U10789 (N_10789,N_10075,N_10167);
nor U10790 (N_10790,N_10430,N_10369);
xnor U10791 (N_10791,N_10497,N_10298);
xor U10792 (N_10792,N_10225,N_10237);
and U10793 (N_10793,N_10360,N_10259);
or U10794 (N_10794,N_10278,N_10210);
nand U10795 (N_10795,N_10251,N_10263);
nor U10796 (N_10796,N_10455,N_10398);
xnor U10797 (N_10797,N_10096,N_10208);
nand U10798 (N_10798,N_10291,N_10210);
and U10799 (N_10799,N_10156,N_10341);
nor U10800 (N_10800,N_10471,N_10384);
or U10801 (N_10801,N_10320,N_10328);
and U10802 (N_10802,N_10109,N_10210);
nor U10803 (N_10803,N_10474,N_10149);
and U10804 (N_10804,N_10074,N_10200);
nand U10805 (N_10805,N_10344,N_10198);
nor U10806 (N_10806,N_10059,N_10491);
nand U10807 (N_10807,N_10384,N_10232);
xor U10808 (N_10808,N_10116,N_10162);
xor U10809 (N_10809,N_10411,N_10046);
nand U10810 (N_10810,N_10474,N_10145);
nand U10811 (N_10811,N_10179,N_10236);
and U10812 (N_10812,N_10180,N_10380);
nor U10813 (N_10813,N_10243,N_10317);
or U10814 (N_10814,N_10412,N_10490);
xor U10815 (N_10815,N_10325,N_10231);
nand U10816 (N_10816,N_10319,N_10377);
or U10817 (N_10817,N_10169,N_10235);
or U10818 (N_10818,N_10304,N_10191);
nor U10819 (N_10819,N_10247,N_10452);
nor U10820 (N_10820,N_10123,N_10081);
and U10821 (N_10821,N_10009,N_10004);
nand U10822 (N_10822,N_10319,N_10351);
nor U10823 (N_10823,N_10357,N_10311);
xnor U10824 (N_10824,N_10213,N_10037);
or U10825 (N_10825,N_10043,N_10380);
xor U10826 (N_10826,N_10469,N_10002);
and U10827 (N_10827,N_10258,N_10444);
xor U10828 (N_10828,N_10114,N_10369);
and U10829 (N_10829,N_10246,N_10018);
or U10830 (N_10830,N_10112,N_10267);
nor U10831 (N_10831,N_10096,N_10318);
nand U10832 (N_10832,N_10097,N_10461);
and U10833 (N_10833,N_10275,N_10108);
and U10834 (N_10834,N_10212,N_10002);
and U10835 (N_10835,N_10275,N_10002);
or U10836 (N_10836,N_10073,N_10397);
and U10837 (N_10837,N_10277,N_10296);
nor U10838 (N_10838,N_10066,N_10104);
nor U10839 (N_10839,N_10084,N_10349);
nor U10840 (N_10840,N_10109,N_10324);
or U10841 (N_10841,N_10016,N_10343);
xnor U10842 (N_10842,N_10315,N_10273);
and U10843 (N_10843,N_10476,N_10382);
nor U10844 (N_10844,N_10322,N_10264);
nor U10845 (N_10845,N_10336,N_10188);
or U10846 (N_10846,N_10054,N_10466);
and U10847 (N_10847,N_10053,N_10241);
or U10848 (N_10848,N_10452,N_10239);
and U10849 (N_10849,N_10045,N_10460);
and U10850 (N_10850,N_10411,N_10404);
and U10851 (N_10851,N_10289,N_10433);
and U10852 (N_10852,N_10324,N_10322);
and U10853 (N_10853,N_10117,N_10298);
xnor U10854 (N_10854,N_10028,N_10414);
nor U10855 (N_10855,N_10115,N_10426);
xnor U10856 (N_10856,N_10227,N_10268);
nor U10857 (N_10857,N_10166,N_10288);
nand U10858 (N_10858,N_10327,N_10474);
or U10859 (N_10859,N_10241,N_10019);
nor U10860 (N_10860,N_10467,N_10485);
xor U10861 (N_10861,N_10178,N_10398);
nor U10862 (N_10862,N_10441,N_10134);
or U10863 (N_10863,N_10211,N_10070);
nand U10864 (N_10864,N_10251,N_10116);
or U10865 (N_10865,N_10225,N_10466);
and U10866 (N_10866,N_10455,N_10426);
and U10867 (N_10867,N_10426,N_10248);
or U10868 (N_10868,N_10302,N_10121);
nand U10869 (N_10869,N_10017,N_10240);
nor U10870 (N_10870,N_10300,N_10175);
nor U10871 (N_10871,N_10009,N_10123);
nand U10872 (N_10872,N_10019,N_10421);
and U10873 (N_10873,N_10373,N_10136);
or U10874 (N_10874,N_10477,N_10206);
xnor U10875 (N_10875,N_10353,N_10398);
nor U10876 (N_10876,N_10094,N_10038);
or U10877 (N_10877,N_10444,N_10039);
xnor U10878 (N_10878,N_10393,N_10058);
nand U10879 (N_10879,N_10032,N_10412);
and U10880 (N_10880,N_10142,N_10305);
xnor U10881 (N_10881,N_10340,N_10084);
and U10882 (N_10882,N_10250,N_10177);
nor U10883 (N_10883,N_10459,N_10274);
or U10884 (N_10884,N_10372,N_10045);
or U10885 (N_10885,N_10028,N_10161);
nand U10886 (N_10886,N_10230,N_10165);
or U10887 (N_10887,N_10434,N_10156);
or U10888 (N_10888,N_10275,N_10120);
and U10889 (N_10889,N_10065,N_10132);
or U10890 (N_10890,N_10000,N_10459);
nand U10891 (N_10891,N_10467,N_10444);
nor U10892 (N_10892,N_10459,N_10015);
nor U10893 (N_10893,N_10344,N_10298);
and U10894 (N_10894,N_10146,N_10445);
and U10895 (N_10895,N_10378,N_10219);
xor U10896 (N_10896,N_10124,N_10476);
nand U10897 (N_10897,N_10398,N_10084);
xor U10898 (N_10898,N_10196,N_10352);
nand U10899 (N_10899,N_10025,N_10036);
xnor U10900 (N_10900,N_10257,N_10080);
or U10901 (N_10901,N_10456,N_10107);
and U10902 (N_10902,N_10451,N_10174);
and U10903 (N_10903,N_10083,N_10049);
or U10904 (N_10904,N_10315,N_10226);
and U10905 (N_10905,N_10396,N_10426);
nand U10906 (N_10906,N_10117,N_10200);
and U10907 (N_10907,N_10233,N_10134);
or U10908 (N_10908,N_10136,N_10000);
nor U10909 (N_10909,N_10335,N_10159);
and U10910 (N_10910,N_10200,N_10394);
xor U10911 (N_10911,N_10184,N_10026);
xnor U10912 (N_10912,N_10472,N_10097);
or U10913 (N_10913,N_10395,N_10376);
and U10914 (N_10914,N_10334,N_10081);
or U10915 (N_10915,N_10303,N_10119);
nor U10916 (N_10916,N_10301,N_10316);
nand U10917 (N_10917,N_10104,N_10048);
xor U10918 (N_10918,N_10480,N_10471);
nor U10919 (N_10919,N_10361,N_10467);
or U10920 (N_10920,N_10212,N_10229);
nor U10921 (N_10921,N_10020,N_10211);
nor U10922 (N_10922,N_10247,N_10192);
xnor U10923 (N_10923,N_10399,N_10407);
nor U10924 (N_10924,N_10126,N_10293);
nor U10925 (N_10925,N_10107,N_10412);
nand U10926 (N_10926,N_10425,N_10171);
or U10927 (N_10927,N_10145,N_10184);
or U10928 (N_10928,N_10179,N_10396);
nor U10929 (N_10929,N_10171,N_10191);
xnor U10930 (N_10930,N_10414,N_10134);
nand U10931 (N_10931,N_10027,N_10033);
and U10932 (N_10932,N_10334,N_10367);
or U10933 (N_10933,N_10021,N_10178);
nand U10934 (N_10934,N_10323,N_10214);
xnor U10935 (N_10935,N_10401,N_10319);
xnor U10936 (N_10936,N_10212,N_10220);
nor U10937 (N_10937,N_10043,N_10119);
xor U10938 (N_10938,N_10144,N_10345);
or U10939 (N_10939,N_10170,N_10232);
or U10940 (N_10940,N_10017,N_10199);
and U10941 (N_10941,N_10168,N_10441);
xnor U10942 (N_10942,N_10085,N_10294);
nor U10943 (N_10943,N_10036,N_10430);
nor U10944 (N_10944,N_10081,N_10194);
nand U10945 (N_10945,N_10321,N_10277);
xor U10946 (N_10946,N_10167,N_10233);
xor U10947 (N_10947,N_10194,N_10067);
or U10948 (N_10948,N_10303,N_10358);
xnor U10949 (N_10949,N_10142,N_10277);
xor U10950 (N_10950,N_10268,N_10078);
and U10951 (N_10951,N_10410,N_10065);
nand U10952 (N_10952,N_10090,N_10366);
or U10953 (N_10953,N_10465,N_10090);
nor U10954 (N_10954,N_10340,N_10499);
or U10955 (N_10955,N_10307,N_10496);
or U10956 (N_10956,N_10062,N_10464);
and U10957 (N_10957,N_10351,N_10425);
nor U10958 (N_10958,N_10035,N_10358);
xnor U10959 (N_10959,N_10213,N_10136);
and U10960 (N_10960,N_10089,N_10071);
nand U10961 (N_10961,N_10291,N_10062);
xor U10962 (N_10962,N_10179,N_10042);
or U10963 (N_10963,N_10240,N_10021);
or U10964 (N_10964,N_10158,N_10002);
nand U10965 (N_10965,N_10411,N_10050);
xor U10966 (N_10966,N_10386,N_10380);
and U10967 (N_10967,N_10158,N_10369);
nor U10968 (N_10968,N_10022,N_10402);
or U10969 (N_10969,N_10043,N_10452);
nor U10970 (N_10970,N_10042,N_10078);
xnor U10971 (N_10971,N_10039,N_10234);
and U10972 (N_10972,N_10220,N_10211);
xor U10973 (N_10973,N_10471,N_10099);
or U10974 (N_10974,N_10163,N_10028);
or U10975 (N_10975,N_10145,N_10259);
nor U10976 (N_10976,N_10430,N_10499);
or U10977 (N_10977,N_10453,N_10493);
xor U10978 (N_10978,N_10242,N_10119);
nand U10979 (N_10979,N_10460,N_10333);
and U10980 (N_10980,N_10410,N_10270);
and U10981 (N_10981,N_10276,N_10496);
and U10982 (N_10982,N_10037,N_10363);
nor U10983 (N_10983,N_10054,N_10215);
nor U10984 (N_10984,N_10111,N_10457);
or U10985 (N_10985,N_10040,N_10095);
and U10986 (N_10986,N_10449,N_10273);
xor U10987 (N_10987,N_10316,N_10289);
xnor U10988 (N_10988,N_10427,N_10473);
nand U10989 (N_10989,N_10409,N_10192);
and U10990 (N_10990,N_10171,N_10010);
or U10991 (N_10991,N_10405,N_10232);
nor U10992 (N_10992,N_10260,N_10105);
or U10993 (N_10993,N_10491,N_10246);
and U10994 (N_10994,N_10395,N_10321);
and U10995 (N_10995,N_10468,N_10363);
nor U10996 (N_10996,N_10479,N_10084);
and U10997 (N_10997,N_10398,N_10392);
nand U10998 (N_10998,N_10058,N_10081);
nor U10999 (N_10999,N_10011,N_10222);
nor U11000 (N_11000,N_10578,N_10517);
xnor U11001 (N_11001,N_10857,N_10814);
and U11002 (N_11002,N_10920,N_10762);
nand U11003 (N_11003,N_10876,N_10829);
nand U11004 (N_11004,N_10951,N_10816);
nor U11005 (N_11005,N_10990,N_10932);
nor U11006 (N_11006,N_10635,N_10620);
and U11007 (N_11007,N_10786,N_10668);
nor U11008 (N_11008,N_10794,N_10708);
xor U11009 (N_11009,N_10864,N_10834);
and U11010 (N_11010,N_10712,N_10541);
nor U11011 (N_11011,N_10874,N_10839);
and U11012 (N_11012,N_10875,N_10883);
xor U11013 (N_11013,N_10580,N_10664);
xnor U11014 (N_11014,N_10858,N_10774);
nand U11015 (N_11015,N_10837,N_10566);
or U11016 (N_11016,N_10583,N_10943);
nor U11017 (N_11017,N_10624,N_10775);
nor U11018 (N_11018,N_10614,N_10910);
xnor U11019 (N_11019,N_10863,N_10529);
nor U11020 (N_11020,N_10944,N_10561);
xnor U11021 (N_11021,N_10528,N_10594);
and U11022 (N_11022,N_10637,N_10592);
nor U11023 (N_11023,N_10731,N_10766);
nor U11024 (N_11024,N_10821,N_10714);
xor U11025 (N_11025,N_10523,N_10573);
xor U11026 (N_11026,N_10900,N_10652);
xor U11027 (N_11027,N_10743,N_10749);
xnor U11028 (N_11028,N_10812,N_10658);
or U11029 (N_11029,N_10723,N_10878);
or U11030 (N_11030,N_10512,N_10880);
and U11031 (N_11031,N_10865,N_10842);
xor U11032 (N_11032,N_10942,N_10901);
nor U11033 (N_11033,N_10520,N_10680);
and U11034 (N_11034,N_10755,N_10673);
xnor U11035 (N_11035,N_10830,N_10947);
xnor U11036 (N_11036,N_10725,N_10805);
xnor U11037 (N_11037,N_10789,N_10584);
or U11038 (N_11038,N_10741,N_10683);
nand U11039 (N_11039,N_10732,N_10778);
or U11040 (N_11040,N_10539,N_10899);
or U11041 (N_11041,N_10911,N_10844);
nand U11042 (N_11042,N_10895,N_10507);
or U11043 (N_11043,N_10540,N_10701);
and U11044 (N_11044,N_10933,N_10846);
nand U11045 (N_11045,N_10519,N_10560);
or U11046 (N_11046,N_10927,N_10660);
nand U11047 (N_11047,N_10610,N_10745);
nor U11048 (N_11048,N_10619,N_10695);
nor U11049 (N_11049,N_10736,N_10969);
or U11050 (N_11050,N_10767,N_10593);
and U11051 (N_11051,N_10729,N_10893);
nor U11052 (N_11052,N_10675,N_10963);
nand U11053 (N_11053,N_10502,N_10815);
nor U11054 (N_11054,N_10717,N_10728);
xnor U11055 (N_11055,N_10831,N_10706);
or U11056 (N_11056,N_10793,N_10980);
or U11057 (N_11057,N_10615,N_10681);
xor U11058 (N_11058,N_10948,N_10656);
nand U11059 (N_11059,N_10824,N_10500);
and U11060 (N_11060,N_10532,N_10785);
xor U11061 (N_11061,N_10609,N_10966);
xor U11062 (N_11062,N_10912,N_10887);
nor U11063 (N_11063,N_10960,N_10935);
or U11064 (N_11064,N_10676,N_10569);
and U11065 (N_11065,N_10562,N_10546);
and U11066 (N_11066,N_10801,N_10626);
nor U11067 (N_11067,N_10853,N_10779);
or U11068 (N_11068,N_10993,N_10738);
nand U11069 (N_11069,N_10945,N_10939);
and U11070 (N_11070,N_10733,N_10894);
and U11071 (N_11071,N_10665,N_10633);
nand U11072 (N_11072,N_10551,N_10661);
nand U11073 (N_11073,N_10559,N_10828);
and U11074 (N_11074,N_10744,N_10757);
nor U11075 (N_11075,N_10555,N_10836);
nor U11076 (N_11076,N_10649,N_10719);
nand U11077 (N_11077,N_10671,N_10697);
xnor U11078 (N_11078,N_10525,N_10672);
or U11079 (N_11079,N_10579,N_10638);
nor U11080 (N_11080,N_10501,N_10711);
nor U11081 (N_11081,N_10538,N_10804);
nand U11082 (N_11082,N_10787,N_10552);
and U11083 (N_11083,N_10575,N_10634);
xor U11084 (N_11084,N_10772,N_10617);
nor U11085 (N_11085,N_10784,N_10913);
nor U11086 (N_11086,N_10931,N_10854);
nand U11087 (N_11087,N_10964,N_10759);
nor U11088 (N_11088,N_10631,N_10760);
xnor U11089 (N_11089,N_10926,N_10896);
nor U11090 (N_11090,N_10897,N_10869);
xor U11091 (N_11091,N_10589,N_10504);
nor U11092 (N_11092,N_10710,N_10817);
nand U11093 (N_11093,N_10563,N_10645);
nor U11094 (N_11094,N_10856,N_10601);
nand U11095 (N_11095,N_10898,N_10915);
nor U11096 (N_11096,N_10696,N_10974);
nor U11097 (N_11097,N_10907,N_10871);
nor U11098 (N_11098,N_10946,N_10768);
and U11099 (N_11099,N_10603,N_10983);
and U11100 (N_11100,N_10748,N_10790);
xor U11101 (N_11101,N_10923,N_10632);
xor U11102 (N_11102,N_10642,N_10536);
nand U11103 (N_11103,N_10999,N_10527);
xnor U11104 (N_11104,N_10773,N_10904);
xnor U11105 (N_11105,N_10859,N_10855);
nand U11106 (N_11106,N_10654,N_10582);
xnor U11107 (N_11107,N_10687,N_10950);
nor U11108 (N_11108,N_10808,N_10798);
nor U11109 (N_11109,N_10550,N_10722);
nand U11110 (N_11110,N_10870,N_10841);
or U11111 (N_11111,N_10558,N_10727);
or U11112 (N_11112,N_10800,N_10758);
nor U11113 (N_11113,N_10991,N_10862);
or U11114 (N_11114,N_10835,N_10694);
and U11115 (N_11115,N_10953,N_10524);
xor U11116 (N_11116,N_10567,N_10505);
and U11117 (N_11117,N_10908,N_10813);
xnor U11118 (N_11118,N_10781,N_10833);
xor U11119 (N_11119,N_10850,N_10998);
nor U11120 (N_11120,N_10522,N_10685);
xnor U11121 (N_11121,N_10674,N_10726);
or U11122 (N_11122,N_10761,N_10995);
or U11123 (N_11123,N_10852,N_10713);
and U11124 (N_11124,N_10616,N_10576);
xor U11125 (N_11125,N_10984,N_10688);
nand U11126 (N_11126,N_10707,N_10678);
nor U11127 (N_11127,N_10892,N_10669);
or U11128 (N_11128,N_10585,N_10699);
or U11129 (N_11129,N_10782,N_10693);
nor U11130 (N_11130,N_10959,N_10845);
xnor U11131 (N_11131,N_10640,N_10659);
nand U11132 (N_11132,N_10613,N_10916);
nand U11133 (N_11133,N_10606,N_10648);
nand U11134 (N_11134,N_10989,N_10735);
xor U11135 (N_11135,N_10849,N_10534);
nand U11136 (N_11136,N_10958,N_10737);
and U11137 (N_11137,N_10508,N_10700);
nand U11138 (N_11138,N_10992,N_10739);
and U11139 (N_11139,N_10509,N_10962);
nor U11140 (N_11140,N_10605,N_10811);
or U11141 (N_11141,N_10791,N_10919);
and U11142 (N_11142,N_10720,N_10590);
nand U11143 (N_11143,N_10877,N_10666);
nand U11144 (N_11144,N_10639,N_10802);
nand U11145 (N_11145,N_10806,N_10771);
nand U11146 (N_11146,N_10868,N_10721);
nor U11147 (N_11147,N_10611,N_10533);
and U11148 (N_11148,N_10882,N_10903);
and U11149 (N_11149,N_10977,N_10651);
nand U11150 (N_11150,N_10703,N_10928);
nor U11151 (N_11151,N_10832,N_10747);
and U11152 (N_11152,N_10797,N_10600);
or U11153 (N_11153,N_10574,N_10776);
nor U11154 (N_11154,N_10577,N_10742);
and U11155 (N_11155,N_10572,N_10885);
and U11156 (N_11156,N_10657,N_10543);
nand U11157 (N_11157,N_10607,N_10556);
nand U11158 (N_11158,N_10702,N_10588);
or U11159 (N_11159,N_10750,N_10765);
or U11160 (N_11160,N_10571,N_10888);
nor U11161 (N_11161,N_10650,N_10819);
nor U11162 (N_11162,N_10630,N_10596);
xnor U11163 (N_11163,N_10861,N_10918);
nor U11164 (N_11164,N_10682,N_10783);
nand U11165 (N_11165,N_10860,N_10746);
and U11166 (N_11166,N_10526,N_10965);
nor U11167 (N_11167,N_10934,N_10866);
nor U11168 (N_11168,N_10810,N_10780);
or U11169 (N_11169,N_10510,N_10840);
nor U11170 (N_11170,N_10752,N_10636);
nor U11171 (N_11171,N_10623,N_10591);
xor U11172 (N_11172,N_10715,N_10604);
xnor U11173 (N_11173,N_10570,N_10602);
nor U11174 (N_11174,N_10655,N_10826);
or U11175 (N_11175,N_10891,N_10647);
nor U11176 (N_11176,N_10629,N_10981);
xor U11177 (N_11177,N_10936,N_10568);
and U11178 (N_11178,N_10518,N_10967);
xor U11179 (N_11179,N_10994,N_10954);
nor U11180 (N_11180,N_10704,N_10734);
nand U11181 (N_11181,N_10922,N_10598);
and U11182 (N_11182,N_10938,N_10586);
nand U11183 (N_11183,N_10564,N_10662);
xor U11184 (N_11184,N_10709,N_10690);
and U11185 (N_11185,N_10553,N_10979);
nor U11186 (N_11186,N_10531,N_10955);
nand U11187 (N_11187,N_10513,N_10957);
and U11188 (N_11188,N_10521,N_10952);
nand U11189 (N_11189,N_10684,N_10881);
nor U11190 (N_11190,N_10547,N_10511);
and U11191 (N_11191,N_10587,N_10925);
xor U11192 (N_11192,N_10986,N_10795);
xor U11193 (N_11193,N_10968,N_10764);
nor U11194 (N_11194,N_10554,N_10971);
or U11195 (N_11195,N_10822,N_10906);
nor U11196 (N_11196,N_10530,N_10996);
and U11197 (N_11197,N_10718,N_10515);
nand U11198 (N_11198,N_10641,N_10843);
xnor U11199 (N_11199,N_10988,N_10941);
nand U11200 (N_11200,N_10879,N_10961);
nand U11201 (N_11201,N_10796,N_10930);
nor U11202 (N_11202,N_10608,N_10982);
xnor U11203 (N_11203,N_10581,N_10730);
nand U11204 (N_11204,N_10970,N_10818);
and U11205 (N_11205,N_10973,N_10917);
nor U11206 (N_11206,N_10646,N_10769);
or U11207 (N_11207,N_10643,N_10848);
xnor U11208 (N_11208,N_10751,N_10788);
or U11209 (N_11209,N_10545,N_10905);
or U11210 (N_11210,N_10825,N_10565);
xor U11211 (N_11211,N_10807,N_10621);
and U11212 (N_11212,N_10987,N_10985);
or U11213 (N_11213,N_10667,N_10686);
nand U11214 (N_11214,N_10777,N_10689);
nor U11215 (N_11215,N_10890,N_10557);
nand U11216 (N_11216,N_10770,N_10653);
nand U11217 (N_11217,N_10909,N_10599);
nand U11218 (N_11218,N_10516,N_10799);
nand U11219 (N_11219,N_10618,N_10625);
and U11220 (N_11220,N_10972,N_10872);
nand U11221 (N_11221,N_10503,N_10692);
nand U11222 (N_11222,N_10940,N_10756);
xor U11223 (N_11223,N_10597,N_10975);
xnor U11224 (N_11224,N_10679,N_10595);
nand U11225 (N_11225,N_10886,N_10716);
nor U11226 (N_11226,N_10754,N_10867);
nand U11227 (N_11227,N_10884,N_10549);
or U11228 (N_11228,N_10997,N_10823);
or U11229 (N_11229,N_10924,N_10544);
xnor U11230 (N_11230,N_10622,N_10514);
nand U11231 (N_11231,N_10691,N_10820);
or U11232 (N_11232,N_10698,N_10792);
nor U11233 (N_11233,N_10644,N_10978);
nand U11234 (N_11234,N_10763,N_10677);
or U11235 (N_11235,N_10506,N_10740);
nor U11236 (N_11236,N_10847,N_10921);
or U11237 (N_11237,N_10535,N_10724);
and U11238 (N_11238,N_10537,N_10670);
xor U11239 (N_11239,N_10914,N_10976);
xnor U11240 (N_11240,N_10548,N_10873);
nand U11241 (N_11241,N_10827,N_10949);
and U11242 (N_11242,N_10628,N_10753);
nand U11243 (N_11243,N_10851,N_10929);
nor U11244 (N_11244,N_10838,N_10809);
and U11245 (N_11245,N_10889,N_10542);
nand U11246 (N_11246,N_10627,N_10612);
nand U11247 (N_11247,N_10705,N_10803);
xnor U11248 (N_11248,N_10902,N_10937);
or U11249 (N_11249,N_10956,N_10663);
nor U11250 (N_11250,N_10808,N_10908);
nor U11251 (N_11251,N_10931,N_10875);
nor U11252 (N_11252,N_10932,N_10724);
nand U11253 (N_11253,N_10927,N_10673);
and U11254 (N_11254,N_10730,N_10743);
nor U11255 (N_11255,N_10749,N_10675);
or U11256 (N_11256,N_10522,N_10912);
nor U11257 (N_11257,N_10646,N_10919);
nand U11258 (N_11258,N_10613,N_10792);
xor U11259 (N_11259,N_10655,N_10687);
nand U11260 (N_11260,N_10671,N_10805);
xor U11261 (N_11261,N_10840,N_10796);
nor U11262 (N_11262,N_10538,N_10721);
nor U11263 (N_11263,N_10835,N_10911);
nand U11264 (N_11264,N_10994,N_10885);
nor U11265 (N_11265,N_10502,N_10681);
xor U11266 (N_11266,N_10869,N_10594);
or U11267 (N_11267,N_10657,N_10735);
or U11268 (N_11268,N_10948,N_10571);
or U11269 (N_11269,N_10539,N_10960);
nor U11270 (N_11270,N_10998,N_10570);
xnor U11271 (N_11271,N_10646,N_10552);
xor U11272 (N_11272,N_10981,N_10761);
and U11273 (N_11273,N_10860,N_10749);
or U11274 (N_11274,N_10646,N_10715);
xor U11275 (N_11275,N_10624,N_10657);
xor U11276 (N_11276,N_10835,N_10939);
or U11277 (N_11277,N_10811,N_10913);
xor U11278 (N_11278,N_10797,N_10585);
xnor U11279 (N_11279,N_10959,N_10798);
nand U11280 (N_11280,N_10684,N_10742);
and U11281 (N_11281,N_10725,N_10869);
or U11282 (N_11282,N_10987,N_10926);
nor U11283 (N_11283,N_10708,N_10959);
or U11284 (N_11284,N_10558,N_10702);
nor U11285 (N_11285,N_10871,N_10529);
nand U11286 (N_11286,N_10670,N_10705);
nor U11287 (N_11287,N_10680,N_10786);
and U11288 (N_11288,N_10891,N_10754);
nand U11289 (N_11289,N_10877,N_10651);
xor U11290 (N_11290,N_10796,N_10581);
nor U11291 (N_11291,N_10778,N_10957);
nor U11292 (N_11292,N_10530,N_10962);
nand U11293 (N_11293,N_10976,N_10663);
nor U11294 (N_11294,N_10593,N_10802);
xnor U11295 (N_11295,N_10745,N_10812);
xor U11296 (N_11296,N_10829,N_10740);
and U11297 (N_11297,N_10934,N_10802);
and U11298 (N_11298,N_10945,N_10858);
nor U11299 (N_11299,N_10815,N_10529);
nor U11300 (N_11300,N_10635,N_10754);
nor U11301 (N_11301,N_10609,N_10980);
or U11302 (N_11302,N_10902,N_10976);
or U11303 (N_11303,N_10776,N_10835);
or U11304 (N_11304,N_10864,N_10546);
xnor U11305 (N_11305,N_10557,N_10704);
nand U11306 (N_11306,N_10617,N_10773);
and U11307 (N_11307,N_10921,N_10628);
and U11308 (N_11308,N_10581,N_10587);
or U11309 (N_11309,N_10943,N_10556);
or U11310 (N_11310,N_10905,N_10568);
and U11311 (N_11311,N_10745,N_10922);
nor U11312 (N_11312,N_10579,N_10885);
nand U11313 (N_11313,N_10747,N_10581);
nand U11314 (N_11314,N_10606,N_10967);
xnor U11315 (N_11315,N_10662,N_10671);
and U11316 (N_11316,N_10920,N_10881);
xor U11317 (N_11317,N_10576,N_10622);
xor U11318 (N_11318,N_10645,N_10635);
nor U11319 (N_11319,N_10535,N_10854);
or U11320 (N_11320,N_10842,N_10784);
or U11321 (N_11321,N_10692,N_10987);
nand U11322 (N_11322,N_10602,N_10704);
and U11323 (N_11323,N_10867,N_10805);
or U11324 (N_11324,N_10781,N_10920);
or U11325 (N_11325,N_10500,N_10619);
or U11326 (N_11326,N_10688,N_10827);
or U11327 (N_11327,N_10758,N_10527);
and U11328 (N_11328,N_10580,N_10968);
xor U11329 (N_11329,N_10616,N_10721);
and U11330 (N_11330,N_10670,N_10596);
xnor U11331 (N_11331,N_10773,N_10856);
or U11332 (N_11332,N_10684,N_10767);
or U11333 (N_11333,N_10957,N_10700);
xor U11334 (N_11334,N_10896,N_10756);
and U11335 (N_11335,N_10715,N_10796);
and U11336 (N_11336,N_10954,N_10741);
xor U11337 (N_11337,N_10812,N_10531);
or U11338 (N_11338,N_10611,N_10892);
xor U11339 (N_11339,N_10793,N_10518);
nor U11340 (N_11340,N_10805,N_10755);
nor U11341 (N_11341,N_10582,N_10818);
or U11342 (N_11342,N_10722,N_10850);
nand U11343 (N_11343,N_10735,N_10731);
and U11344 (N_11344,N_10956,N_10812);
xnor U11345 (N_11345,N_10924,N_10737);
or U11346 (N_11346,N_10699,N_10834);
or U11347 (N_11347,N_10701,N_10792);
xor U11348 (N_11348,N_10834,N_10576);
xnor U11349 (N_11349,N_10815,N_10538);
xnor U11350 (N_11350,N_10509,N_10833);
xnor U11351 (N_11351,N_10953,N_10888);
nor U11352 (N_11352,N_10533,N_10577);
nor U11353 (N_11353,N_10783,N_10760);
or U11354 (N_11354,N_10921,N_10682);
nand U11355 (N_11355,N_10966,N_10911);
nor U11356 (N_11356,N_10651,N_10964);
nand U11357 (N_11357,N_10533,N_10864);
nor U11358 (N_11358,N_10915,N_10689);
or U11359 (N_11359,N_10660,N_10625);
xnor U11360 (N_11360,N_10678,N_10872);
and U11361 (N_11361,N_10786,N_10859);
nor U11362 (N_11362,N_10943,N_10572);
or U11363 (N_11363,N_10521,N_10549);
nor U11364 (N_11364,N_10665,N_10610);
xnor U11365 (N_11365,N_10916,N_10566);
and U11366 (N_11366,N_10818,N_10766);
xnor U11367 (N_11367,N_10664,N_10666);
or U11368 (N_11368,N_10958,N_10985);
or U11369 (N_11369,N_10540,N_10599);
and U11370 (N_11370,N_10644,N_10554);
nand U11371 (N_11371,N_10648,N_10866);
xnor U11372 (N_11372,N_10543,N_10508);
or U11373 (N_11373,N_10517,N_10759);
nand U11374 (N_11374,N_10828,N_10731);
and U11375 (N_11375,N_10937,N_10889);
nor U11376 (N_11376,N_10546,N_10727);
or U11377 (N_11377,N_10798,N_10593);
nand U11378 (N_11378,N_10501,N_10839);
and U11379 (N_11379,N_10789,N_10886);
nand U11380 (N_11380,N_10531,N_10764);
xnor U11381 (N_11381,N_10869,N_10643);
and U11382 (N_11382,N_10984,N_10924);
xor U11383 (N_11383,N_10950,N_10548);
xor U11384 (N_11384,N_10580,N_10593);
and U11385 (N_11385,N_10581,N_10669);
or U11386 (N_11386,N_10855,N_10706);
nand U11387 (N_11387,N_10554,N_10964);
xnor U11388 (N_11388,N_10730,N_10640);
nand U11389 (N_11389,N_10683,N_10583);
nand U11390 (N_11390,N_10923,N_10555);
nor U11391 (N_11391,N_10858,N_10989);
or U11392 (N_11392,N_10667,N_10543);
nand U11393 (N_11393,N_10847,N_10969);
nand U11394 (N_11394,N_10919,N_10502);
or U11395 (N_11395,N_10657,N_10704);
xnor U11396 (N_11396,N_10603,N_10673);
xor U11397 (N_11397,N_10946,N_10971);
nor U11398 (N_11398,N_10918,N_10699);
and U11399 (N_11399,N_10671,N_10715);
and U11400 (N_11400,N_10806,N_10555);
nor U11401 (N_11401,N_10720,N_10568);
and U11402 (N_11402,N_10861,N_10550);
nand U11403 (N_11403,N_10797,N_10552);
nor U11404 (N_11404,N_10779,N_10759);
and U11405 (N_11405,N_10765,N_10622);
or U11406 (N_11406,N_10840,N_10799);
nor U11407 (N_11407,N_10898,N_10950);
nand U11408 (N_11408,N_10942,N_10663);
or U11409 (N_11409,N_10995,N_10911);
nor U11410 (N_11410,N_10780,N_10513);
xor U11411 (N_11411,N_10912,N_10503);
nand U11412 (N_11412,N_10984,N_10995);
nand U11413 (N_11413,N_10744,N_10580);
or U11414 (N_11414,N_10731,N_10754);
or U11415 (N_11415,N_10874,N_10948);
nand U11416 (N_11416,N_10814,N_10800);
xnor U11417 (N_11417,N_10626,N_10509);
xnor U11418 (N_11418,N_10612,N_10591);
and U11419 (N_11419,N_10678,N_10841);
nand U11420 (N_11420,N_10767,N_10541);
and U11421 (N_11421,N_10932,N_10576);
and U11422 (N_11422,N_10804,N_10682);
xor U11423 (N_11423,N_10569,N_10621);
or U11424 (N_11424,N_10516,N_10562);
or U11425 (N_11425,N_10858,N_10863);
xor U11426 (N_11426,N_10635,N_10999);
xnor U11427 (N_11427,N_10580,N_10777);
xor U11428 (N_11428,N_10850,N_10961);
or U11429 (N_11429,N_10874,N_10687);
nand U11430 (N_11430,N_10950,N_10723);
nor U11431 (N_11431,N_10652,N_10654);
xnor U11432 (N_11432,N_10873,N_10835);
nand U11433 (N_11433,N_10649,N_10510);
and U11434 (N_11434,N_10929,N_10524);
or U11435 (N_11435,N_10886,N_10931);
and U11436 (N_11436,N_10902,N_10985);
nor U11437 (N_11437,N_10554,N_10926);
nor U11438 (N_11438,N_10575,N_10608);
and U11439 (N_11439,N_10926,N_10718);
nor U11440 (N_11440,N_10822,N_10965);
nor U11441 (N_11441,N_10585,N_10577);
xor U11442 (N_11442,N_10608,N_10708);
and U11443 (N_11443,N_10705,N_10721);
and U11444 (N_11444,N_10746,N_10975);
or U11445 (N_11445,N_10971,N_10684);
nor U11446 (N_11446,N_10942,N_10781);
nor U11447 (N_11447,N_10735,N_10676);
xor U11448 (N_11448,N_10851,N_10679);
or U11449 (N_11449,N_10994,N_10567);
nor U11450 (N_11450,N_10615,N_10519);
nor U11451 (N_11451,N_10779,N_10755);
nand U11452 (N_11452,N_10886,N_10698);
nor U11453 (N_11453,N_10764,N_10917);
and U11454 (N_11454,N_10669,N_10781);
xnor U11455 (N_11455,N_10717,N_10953);
or U11456 (N_11456,N_10655,N_10849);
nand U11457 (N_11457,N_10673,N_10914);
nand U11458 (N_11458,N_10773,N_10514);
and U11459 (N_11459,N_10671,N_10767);
nand U11460 (N_11460,N_10736,N_10918);
or U11461 (N_11461,N_10688,N_10563);
nand U11462 (N_11462,N_10561,N_10825);
nor U11463 (N_11463,N_10641,N_10861);
nor U11464 (N_11464,N_10836,N_10953);
xnor U11465 (N_11465,N_10919,N_10531);
nand U11466 (N_11466,N_10895,N_10885);
xnor U11467 (N_11467,N_10554,N_10729);
nor U11468 (N_11468,N_10767,N_10781);
and U11469 (N_11469,N_10741,N_10780);
or U11470 (N_11470,N_10654,N_10581);
nand U11471 (N_11471,N_10605,N_10549);
or U11472 (N_11472,N_10818,N_10868);
or U11473 (N_11473,N_10820,N_10989);
nor U11474 (N_11474,N_10694,N_10684);
nor U11475 (N_11475,N_10823,N_10707);
nand U11476 (N_11476,N_10604,N_10599);
nand U11477 (N_11477,N_10539,N_10686);
xor U11478 (N_11478,N_10685,N_10906);
or U11479 (N_11479,N_10791,N_10822);
nand U11480 (N_11480,N_10879,N_10661);
and U11481 (N_11481,N_10893,N_10920);
nand U11482 (N_11482,N_10733,N_10685);
and U11483 (N_11483,N_10798,N_10963);
nor U11484 (N_11484,N_10660,N_10878);
or U11485 (N_11485,N_10709,N_10693);
nor U11486 (N_11486,N_10519,N_10870);
or U11487 (N_11487,N_10797,N_10589);
or U11488 (N_11488,N_10514,N_10908);
xnor U11489 (N_11489,N_10881,N_10978);
nor U11490 (N_11490,N_10533,N_10928);
and U11491 (N_11491,N_10584,N_10966);
nor U11492 (N_11492,N_10976,N_10560);
nor U11493 (N_11493,N_10869,N_10872);
xor U11494 (N_11494,N_10577,N_10601);
xnor U11495 (N_11495,N_10990,N_10923);
and U11496 (N_11496,N_10566,N_10824);
and U11497 (N_11497,N_10630,N_10837);
xnor U11498 (N_11498,N_10610,N_10824);
and U11499 (N_11499,N_10745,N_10505);
xnor U11500 (N_11500,N_11353,N_11082);
or U11501 (N_11501,N_11260,N_11072);
and U11502 (N_11502,N_11471,N_11302);
and U11503 (N_11503,N_11381,N_11480);
or U11504 (N_11504,N_11290,N_11374);
or U11505 (N_11505,N_11363,N_11130);
xor U11506 (N_11506,N_11410,N_11437);
or U11507 (N_11507,N_11311,N_11236);
and U11508 (N_11508,N_11203,N_11074);
and U11509 (N_11509,N_11132,N_11219);
and U11510 (N_11510,N_11150,N_11270);
nor U11511 (N_11511,N_11498,N_11327);
xnor U11512 (N_11512,N_11169,N_11456);
and U11513 (N_11513,N_11326,N_11265);
nand U11514 (N_11514,N_11099,N_11312);
and U11515 (N_11515,N_11070,N_11445);
nand U11516 (N_11516,N_11221,N_11448);
nand U11517 (N_11517,N_11494,N_11035);
xor U11518 (N_11518,N_11458,N_11159);
or U11519 (N_11519,N_11325,N_11249);
xnor U11520 (N_11520,N_11168,N_11447);
or U11521 (N_11521,N_11075,N_11131);
nor U11522 (N_11522,N_11129,N_11235);
or U11523 (N_11523,N_11332,N_11063);
and U11524 (N_11524,N_11313,N_11330);
nand U11525 (N_11525,N_11020,N_11419);
nor U11526 (N_11526,N_11119,N_11222);
nand U11527 (N_11527,N_11194,N_11039);
xor U11528 (N_11528,N_11286,N_11014);
or U11529 (N_11529,N_11041,N_11422);
xor U11530 (N_11530,N_11397,N_11375);
or U11531 (N_11531,N_11308,N_11036);
nor U11532 (N_11532,N_11090,N_11151);
xnor U11533 (N_11533,N_11412,N_11100);
xor U11534 (N_11534,N_11413,N_11011);
nand U11535 (N_11535,N_11238,N_11124);
or U11536 (N_11536,N_11182,N_11495);
and U11537 (N_11537,N_11097,N_11190);
xor U11538 (N_11538,N_11256,N_11479);
or U11539 (N_11539,N_11152,N_11490);
nand U11540 (N_11540,N_11186,N_11263);
xnor U11541 (N_11541,N_11395,N_11078);
or U11542 (N_11542,N_11010,N_11389);
and U11543 (N_11543,N_11394,N_11002);
or U11544 (N_11544,N_11218,N_11300);
xor U11545 (N_11545,N_11154,N_11466);
xnor U11546 (N_11546,N_11291,N_11009);
xor U11547 (N_11547,N_11289,N_11157);
nor U11548 (N_11548,N_11279,N_11003);
nand U11549 (N_11549,N_11320,N_11367);
or U11550 (N_11550,N_11175,N_11391);
and U11551 (N_11551,N_11296,N_11434);
xor U11552 (N_11552,N_11066,N_11319);
nor U11553 (N_11553,N_11259,N_11250);
and U11554 (N_11554,N_11164,N_11161);
or U11555 (N_11555,N_11461,N_11073);
nor U11556 (N_11556,N_11133,N_11085);
nor U11557 (N_11557,N_11209,N_11406);
and U11558 (N_11558,N_11470,N_11442);
and U11559 (N_11559,N_11147,N_11370);
nor U11560 (N_11560,N_11081,N_11053);
nor U11561 (N_11561,N_11000,N_11191);
nand U11562 (N_11562,N_11188,N_11115);
nand U11563 (N_11563,N_11058,N_11087);
nor U11564 (N_11564,N_11452,N_11455);
nor U11565 (N_11565,N_11226,N_11364);
or U11566 (N_11566,N_11469,N_11369);
and U11567 (N_11567,N_11460,N_11232);
nor U11568 (N_11568,N_11478,N_11059);
and U11569 (N_11569,N_11243,N_11481);
and U11570 (N_11570,N_11262,N_11379);
nand U11571 (N_11571,N_11040,N_11276);
nand U11572 (N_11572,N_11254,N_11165);
xor U11573 (N_11573,N_11231,N_11468);
or U11574 (N_11574,N_11069,N_11107);
or U11575 (N_11575,N_11368,N_11359);
nor U11576 (N_11576,N_11033,N_11184);
and U11577 (N_11577,N_11068,N_11148);
and U11578 (N_11578,N_11025,N_11357);
or U11579 (N_11579,N_11143,N_11083);
or U11580 (N_11580,N_11292,N_11449);
and U11581 (N_11581,N_11163,N_11344);
nand U11582 (N_11582,N_11427,N_11376);
or U11583 (N_11583,N_11299,N_11295);
xor U11584 (N_11584,N_11287,N_11323);
nand U11585 (N_11585,N_11465,N_11398);
or U11586 (N_11586,N_11060,N_11217);
xor U11587 (N_11587,N_11104,N_11421);
nor U11588 (N_11588,N_11179,N_11120);
xnor U11589 (N_11589,N_11360,N_11430);
and U11590 (N_11590,N_11021,N_11354);
or U11591 (N_11591,N_11482,N_11281);
or U11592 (N_11592,N_11349,N_11228);
nor U11593 (N_11593,N_11028,N_11185);
nand U11594 (N_11594,N_11472,N_11122);
nor U11595 (N_11595,N_11230,N_11372);
and U11596 (N_11596,N_11183,N_11212);
xnor U11597 (N_11597,N_11089,N_11170);
nand U11598 (N_11598,N_11392,N_11283);
or U11599 (N_11599,N_11453,N_11441);
or U11600 (N_11600,N_11192,N_11264);
nand U11601 (N_11601,N_11483,N_11172);
nand U11602 (N_11602,N_11019,N_11001);
xnor U11603 (N_11603,N_11196,N_11269);
or U11604 (N_11604,N_11024,N_11318);
nand U11605 (N_11605,N_11493,N_11136);
nand U11606 (N_11606,N_11213,N_11390);
or U11607 (N_11607,N_11285,N_11373);
or U11608 (N_11608,N_11486,N_11110);
nor U11609 (N_11609,N_11403,N_11111);
and U11610 (N_11610,N_11464,N_11298);
xor U11611 (N_11611,N_11012,N_11239);
xor U11612 (N_11612,N_11223,N_11337);
nor U11613 (N_11613,N_11436,N_11140);
or U11614 (N_11614,N_11432,N_11492);
and U11615 (N_11615,N_11252,N_11386);
nand U11616 (N_11616,N_11034,N_11102);
nor U11617 (N_11617,N_11303,N_11361);
xor U11618 (N_11618,N_11229,N_11206);
nor U11619 (N_11619,N_11031,N_11489);
and U11620 (N_11620,N_11261,N_11418);
nand U11621 (N_11621,N_11329,N_11310);
or U11622 (N_11622,N_11103,N_11399);
nor U11623 (N_11623,N_11156,N_11016);
nand U11624 (N_11624,N_11384,N_11193);
nor U11625 (N_11625,N_11268,N_11027);
nor U11626 (N_11626,N_11258,N_11348);
nor U11627 (N_11627,N_11155,N_11056);
nand U11628 (N_11628,N_11114,N_11116);
nand U11629 (N_11629,N_11401,N_11038);
or U11630 (N_11630,N_11255,N_11091);
or U11631 (N_11631,N_11008,N_11022);
xor U11632 (N_11632,N_11032,N_11315);
or U11633 (N_11633,N_11121,N_11439);
nand U11634 (N_11634,N_11433,N_11144);
and U11635 (N_11635,N_11267,N_11273);
nand U11636 (N_11636,N_11309,N_11065);
and U11637 (N_11637,N_11429,N_11146);
nand U11638 (N_11638,N_11197,N_11109);
nor U11639 (N_11639,N_11352,N_11180);
nand U11640 (N_11640,N_11079,N_11350);
nor U11641 (N_11641,N_11378,N_11037);
or U11642 (N_11642,N_11201,N_11257);
or U11643 (N_11643,N_11029,N_11057);
nor U11644 (N_11644,N_11338,N_11076);
nor U11645 (N_11645,N_11476,N_11496);
nand U11646 (N_11646,N_11048,N_11380);
xor U11647 (N_11647,N_11139,N_11205);
or U11648 (N_11648,N_11137,N_11307);
and U11649 (N_11649,N_11088,N_11431);
nor U11650 (N_11650,N_11142,N_11280);
and U11651 (N_11651,N_11225,N_11328);
and U11652 (N_11652,N_11108,N_11198);
nand U11653 (N_11653,N_11297,N_11451);
and U11654 (N_11654,N_11177,N_11178);
and U11655 (N_11655,N_11084,N_11026);
nor U11656 (N_11656,N_11336,N_11207);
and U11657 (N_11657,N_11202,N_11126);
or U11658 (N_11658,N_11341,N_11485);
or U11659 (N_11659,N_11450,N_11007);
xnor U11660 (N_11660,N_11400,N_11061);
nand U11661 (N_11661,N_11416,N_11105);
or U11662 (N_11662,N_11017,N_11050);
nor U11663 (N_11663,N_11098,N_11118);
nand U11664 (N_11664,N_11162,N_11306);
and U11665 (N_11665,N_11405,N_11342);
nand U11666 (N_11666,N_11459,N_11404);
and U11667 (N_11667,N_11055,N_11467);
or U11668 (N_11668,N_11117,N_11135);
nor U11669 (N_11669,N_11444,N_11095);
or U11670 (N_11670,N_11062,N_11317);
or U11671 (N_11671,N_11324,N_11284);
nand U11672 (N_11672,N_11385,N_11211);
or U11673 (N_11673,N_11425,N_11477);
nor U11674 (N_11674,N_11340,N_11424);
and U11675 (N_11675,N_11475,N_11294);
or U11676 (N_11676,N_11153,N_11371);
and U11677 (N_11677,N_11387,N_11123);
nor U11678 (N_11678,N_11195,N_11176);
and U11679 (N_11679,N_11339,N_11042);
xor U11680 (N_11680,N_11094,N_11051);
nor U11681 (N_11681,N_11277,N_11138);
nand U11682 (N_11682,N_11288,N_11167);
nor U11683 (N_11683,N_11015,N_11077);
and U11684 (N_11684,N_11345,N_11047);
nand U11685 (N_11685,N_11305,N_11388);
xnor U11686 (N_11686,N_11272,N_11365);
xor U11687 (N_11687,N_11141,N_11210);
or U11688 (N_11688,N_11301,N_11127);
and U11689 (N_11689,N_11244,N_11491);
nand U11690 (N_11690,N_11488,N_11484);
or U11691 (N_11691,N_11145,N_11187);
or U11692 (N_11692,N_11420,N_11086);
and U11693 (N_11693,N_11160,N_11358);
xor U11694 (N_11694,N_11253,N_11242);
xnor U11695 (N_11695,N_11064,N_11247);
or U11696 (N_11696,N_11174,N_11474);
or U11697 (N_11697,N_11473,N_11149);
xor U11698 (N_11698,N_11233,N_11393);
nor U11699 (N_11699,N_11248,N_11049);
xnor U11700 (N_11700,N_11227,N_11234);
xor U11701 (N_11701,N_11125,N_11215);
and U11702 (N_11702,N_11246,N_11383);
nor U11703 (N_11703,N_11356,N_11106);
xnor U11704 (N_11704,N_11237,N_11414);
xor U11705 (N_11705,N_11457,N_11266);
nand U11706 (N_11706,N_11045,N_11046);
or U11707 (N_11707,N_11101,N_11463);
and U11708 (N_11708,N_11171,N_11173);
nand U11709 (N_11709,N_11275,N_11402);
xor U11710 (N_11710,N_11181,N_11426);
and U11711 (N_11711,N_11415,N_11052);
nand U11712 (N_11712,N_11335,N_11497);
or U11713 (N_11713,N_11351,N_11487);
xor U11714 (N_11714,N_11321,N_11271);
nand U11715 (N_11715,N_11013,N_11134);
xor U11716 (N_11716,N_11018,N_11274);
nor U11717 (N_11717,N_11366,N_11417);
xnor U11718 (N_11718,N_11023,N_11220);
nor U11719 (N_11719,N_11128,N_11362);
nor U11720 (N_11720,N_11454,N_11006);
xor U11721 (N_11721,N_11440,N_11216);
and U11722 (N_11722,N_11343,N_11446);
or U11723 (N_11723,N_11240,N_11499);
and U11724 (N_11724,N_11204,N_11093);
or U11725 (N_11725,N_11408,N_11331);
or U11726 (N_11726,N_11438,N_11282);
xnor U11727 (N_11727,N_11005,N_11428);
xor U11728 (N_11728,N_11241,N_11158);
nand U11729 (N_11729,N_11314,N_11199);
xor U11730 (N_11730,N_11054,N_11278);
xor U11731 (N_11731,N_11347,N_11334);
xnor U11732 (N_11732,N_11245,N_11409);
nand U11733 (N_11733,N_11435,N_11346);
xnor U11734 (N_11734,N_11443,N_11214);
or U11735 (N_11735,N_11113,N_11316);
nor U11736 (N_11736,N_11293,N_11200);
xnor U11737 (N_11737,N_11377,N_11396);
nand U11738 (N_11738,N_11251,N_11411);
nor U11739 (N_11739,N_11030,N_11423);
and U11740 (N_11740,N_11096,N_11166);
nor U11741 (N_11741,N_11044,N_11112);
nor U11742 (N_11742,N_11071,N_11208);
or U11743 (N_11743,N_11067,N_11322);
nor U11744 (N_11744,N_11333,N_11224);
nand U11745 (N_11745,N_11080,N_11462);
nor U11746 (N_11746,N_11407,N_11004);
nand U11747 (N_11747,N_11043,N_11382);
or U11748 (N_11748,N_11355,N_11092);
or U11749 (N_11749,N_11189,N_11304);
xnor U11750 (N_11750,N_11483,N_11218);
nor U11751 (N_11751,N_11293,N_11313);
xor U11752 (N_11752,N_11469,N_11313);
or U11753 (N_11753,N_11218,N_11001);
nor U11754 (N_11754,N_11280,N_11351);
xnor U11755 (N_11755,N_11195,N_11077);
and U11756 (N_11756,N_11011,N_11415);
xor U11757 (N_11757,N_11458,N_11309);
or U11758 (N_11758,N_11290,N_11107);
or U11759 (N_11759,N_11389,N_11148);
nand U11760 (N_11760,N_11184,N_11339);
xor U11761 (N_11761,N_11468,N_11145);
xor U11762 (N_11762,N_11033,N_11292);
nand U11763 (N_11763,N_11420,N_11440);
and U11764 (N_11764,N_11185,N_11410);
or U11765 (N_11765,N_11348,N_11320);
or U11766 (N_11766,N_11014,N_11298);
nor U11767 (N_11767,N_11291,N_11089);
or U11768 (N_11768,N_11252,N_11139);
and U11769 (N_11769,N_11446,N_11027);
nor U11770 (N_11770,N_11449,N_11348);
and U11771 (N_11771,N_11417,N_11095);
nor U11772 (N_11772,N_11265,N_11173);
xnor U11773 (N_11773,N_11330,N_11417);
nand U11774 (N_11774,N_11299,N_11422);
or U11775 (N_11775,N_11303,N_11360);
xor U11776 (N_11776,N_11064,N_11157);
xor U11777 (N_11777,N_11458,N_11479);
xnor U11778 (N_11778,N_11326,N_11349);
nor U11779 (N_11779,N_11325,N_11083);
and U11780 (N_11780,N_11302,N_11199);
or U11781 (N_11781,N_11385,N_11182);
nor U11782 (N_11782,N_11251,N_11011);
nand U11783 (N_11783,N_11202,N_11433);
xnor U11784 (N_11784,N_11257,N_11242);
xnor U11785 (N_11785,N_11219,N_11142);
and U11786 (N_11786,N_11272,N_11299);
nor U11787 (N_11787,N_11095,N_11278);
and U11788 (N_11788,N_11309,N_11446);
nor U11789 (N_11789,N_11020,N_11472);
nand U11790 (N_11790,N_11163,N_11251);
nand U11791 (N_11791,N_11293,N_11089);
xnor U11792 (N_11792,N_11115,N_11259);
and U11793 (N_11793,N_11489,N_11202);
and U11794 (N_11794,N_11333,N_11087);
or U11795 (N_11795,N_11053,N_11336);
and U11796 (N_11796,N_11484,N_11074);
xor U11797 (N_11797,N_11002,N_11462);
xnor U11798 (N_11798,N_11100,N_11172);
nand U11799 (N_11799,N_11206,N_11015);
and U11800 (N_11800,N_11420,N_11352);
and U11801 (N_11801,N_11105,N_11292);
nor U11802 (N_11802,N_11245,N_11108);
or U11803 (N_11803,N_11253,N_11461);
nor U11804 (N_11804,N_11451,N_11015);
nor U11805 (N_11805,N_11089,N_11335);
and U11806 (N_11806,N_11168,N_11088);
or U11807 (N_11807,N_11452,N_11037);
and U11808 (N_11808,N_11221,N_11019);
nor U11809 (N_11809,N_11183,N_11030);
and U11810 (N_11810,N_11492,N_11291);
xor U11811 (N_11811,N_11312,N_11231);
xor U11812 (N_11812,N_11108,N_11428);
xnor U11813 (N_11813,N_11313,N_11182);
nor U11814 (N_11814,N_11053,N_11422);
and U11815 (N_11815,N_11459,N_11152);
nand U11816 (N_11816,N_11065,N_11422);
nand U11817 (N_11817,N_11369,N_11230);
xnor U11818 (N_11818,N_11413,N_11024);
xnor U11819 (N_11819,N_11046,N_11014);
xor U11820 (N_11820,N_11044,N_11260);
xor U11821 (N_11821,N_11092,N_11053);
xor U11822 (N_11822,N_11226,N_11135);
nor U11823 (N_11823,N_11462,N_11040);
xnor U11824 (N_11824,N_11413,N_11318);
nand U11825 (N_11825,N_11205,N_11376);
xor U11826 (N_11826,N_11249,N_11297);
xnor U11827 (N_11827,N_11276,N_11157);
xnor U11828 (N_11828,N_11269,N_11078);
nand U11829 (N_11829,N_11382,N_11481);
xor U11830 (N_11830,N_11154,N_11031);
xnor U11831 (N_11831,N_11255,N_11415);
xor U11832 (N_11832,N_11071,N_11338);
or U11833 (N_11833,N_11247,N_11437);
or U11834 (N_11834,N_11423,N_11366);
nand U11835 (N_11835,N_11443,N_11070);
or U11836 (N_11836,N_11138,N_11043);
or U11837 (N_11837,N_11225,N_11181);
nor U11838 (N_11838,N_11145,N_11273);
nand U11839 (N_11839,N_11245,N_11063);
or U11840 (N_11840,N_11401,N_11340);
or U11841 (N_11841,N_11405,N_11061);
and U11842 (N_11842,N_11423,N_11207);
nand U11843 (N_11843,N_11453,N_11012);
and U11844 (N_11844,N_11475,N_11143);
nand U11845 (N_11845,N_11159,N_11232);
nor U11846 (N_11846,N_11105,N_11396);
or U11847 (N_11847,N_11230,N_11330);
nor U11848 (N_11848,N_11176,N_11083);
xnor U11849 (N_11849,N_11068,N_11122);
and U11850 (N_11850,N_11380,N_11243);
and U11851 (N_11851,N_11156,N_11368);
nand U11852 (N_11852,N_11169,N_11182);
and U11853 (N_11853,N_11413,N_11395);
or U11854 (N_11854,N_11269,N_11210);
and U11855 (N_11855,N_11035,N_11443);
and U11856 (N_11856,N_11401,N_11225);
xnor U11857 (N_11857,N_11431,N_11096);
xor U11858 (N_11858,N_11161,N_11325);
or U11859 (N_11859,N_11006,N_11066);
nor U11860 (N_11860,N_11492,N_11268);
and U11861 (N_11861,N_11128,N_11224);
xor U11862 (N_11862,N_11492,N_11093);
and U11863 (N_11863,N_11125,N_11390);
nor U11864 (N_11864,N_11271,N_11241);
and U11865 (N_11865,N_11476,N_11343);
xnor U11866 (N_11866,N_11331,N_11277);
nand U11867 (N_11867,N_11231,N_11496);
xnor U11868 (N_11868,N_11030,N_11346);
nand U11869 (N_11869,N_11254,N_11067);
nor U11870 (N_11870,N_11416,N_11296);
nor U11871 (N_11871,N_11060,N_11320);
xnor U11872 (N_11872,N_11118,N_11478);
nor U11873 (N_11873,N_11488,N_11347);
nand U11874 (N_11874,N_11031,N_11221);
xor U11875 (N_11875,N_11462,N_11118);
nor U11876 (N_11876,N_11467,N_11294);
nand U11877 (N_11877,N_11053,N_11056);
nand U11878 (N_11878,N_11468,N_11170);
or U11879 (N_11879,N_11032,N_11483);
xor U11880 (N_11880,N_11074,N_11154);
nor U11881 (N_11881,N_11102,N_11366);
or U11882 (N_11882,N_11288,N_11125);
nor U11883 (N_11883,N_11258,N_11455);
nand U11884 (N_11884,N_11260,N_11384);
nor U11885 (N_11885,N_11349,N_11189);
nor U11886 (N_11886,N_11210,N_11377);
nand U11887 (N_11887,N_11064,N_11262);
or U11888 (N_11888,N_11313,N_11149);
or U11889 (N_11889,N_11479,N_11201);
nand U11890 (N_11890,N_11241,N_11034);
and U11891 (N_11891,N_11370,N_11242);
or U11892 (N_11892,N_11416,N_11080);
xnor U11893 (N_11893,N_11104,N_11403);
nand U11894 (N_11894,N_11354,N_11120);
or U11895 (N_11895,N_11230,N_11172);
and U11896 (N_11896,N_11185,N_11412);
nand U11897 (N_11897,N_11256,N_11424);
and U11898 (N_11898,N_11462,N_11427);
xnor U11899 (N_11899,N_11080,N_11081);
or U11900 (N_11900,N_11082,N_11463);
xor U11901 (N_11901,N_11232,N_11174);
nand U11902 (N_11902,N_11470,N_11324);
and U11903 (N_11903,N_11048,N_11412);
or U11904 (N_11904,N_11169,N_11131);
xor U11905 (N_11905,N_11307,N_11331);
xnor U11906 (N_11906,N_11313,N_11080);
xnor U11907 (N_11907,N_11016,N_11190);
nor U11908 (N_11908,N_11315,N_11330);
nor U11909 (N_11909,N_11231,N_11333);
nor U11910 (N_11910,N_11479,N_11010);
xnor U11911 (N_11911,N_11316,N_11133);
nor U11912 (N_11912,N_11336,N_11031);
nand U11913 (N_11913,N_11438,N_11212);
and U11914 (N_11914,N_11186,N_11297);
xor U11915 (N_11915,N_11032,N_11142);
and U11916 (N_11916,N_11212,N_11034);
nor U11917 (N_11917,N_11279,N_11236);
xor U11918 (N_11918,N_11272,N_11397);
xor U11919 (N_11919,N_11262,N_11463);
xor U11920 (N_11920,N_11052,N_11346);
nand U11921 (N_11921,N_11255,N_11005);
nor U11922 (N_11922,N_11084,N_11216);
xor U11923 (N_11923,N_11082,N_11150);
nand U11924 (N_11924,N_11293,N_11425);
and U11925 (N_11925,N_11225,N_11114);
xor U11926 (N_11926,N_11027,N_11117);
nand U11927 (N_11927,N_11279,N_11169);
and U11928 (N_11928,N_11426,N_11262);
nand U11929 (N_11929,N_11266,N_11099);
nand U11930 (N_11930,N_11336,N_11379);
nand U11931 (N_11931,N_11133,N_11044);
xor U11932 (N_11932,N_11373,N_11345);
or U11933 (N_11933,N_11185,N_11132);
or U11934 (N_11934,N_11448,N_11166);
and U11935 (N_11935,N_11286,N_11450);
or U11936 (N_11936,N_11489,N_11062);
or U11937 (N_11937,N_11045,N_11219);
xor U11938 (N_11938,N_11428,N_11213);
nor U11939 (N_11939,N_11092,N_11151);
nand U11940 (N_11940,N_11140,N_11494);
nand U11941 (N_11941,N_11140,N_11121);
and U11942 (N_11942,N_11202,N_11414);
nand U11943 (N_11943,N_11274,N_11061);
nor U11944 (N_11944,N_11119,N_11341);
nor U11945 (N_11945,N_11400,N_11423);
nor U11946 (N_11946,N_11427,N_11438);
xnor U11947 (N_11947,N_11352,N_11254);
and U11948 (N_11948,N_11196,N_11352);
nor U11949 (N_11949,N_11447,N_11477);
xnor U11950 (N_11950,N_11111,N_11134);
nor U11951 (N_11951,N_11429,N_11155);
or U11952 (N_11952,N_11470,N_11386);
and U11953 (N_11953,N_11153,N_11188);
and U11954 (N_11954,N_11214,N_11128);
and U11955 (N_11955,N_11162,N_11013);
or U11956 (N_11956,N_11293,N_11145);
xnor U11957 (N_11957,N_11407,N_11081);
and U11958 (N_11958,N_11476,N_11458);
or U11959 (N_11959,N_11358,N_11109);
xor U11960 (N_11960,N_11412,N_11176);
or U11961 (N_11961,N_11490,N_11047);
and U11962 (N_11962,N_11047,N_11343);
or U11963 (N_11963,N_11254,N_11331);
xor U11964 (N_11964,N_11469,N_11202);
or U11965 (N_11965,N_11467,N_11115);
nor U11966 (N_11966,N_11011,N_11378);
nand U11967 (N_11967,N_11242,N_11180);
xor U11968 (N_11968,N_11362,N_11048);
xnor U11969 (N_11969,N_11241,N_11341);
or U11970 (N_11970,N_11335,N_11496);
or U11971 (N_11971,N_11192,N_11301);
nand U11972 (N_11972,N_11350,N_11400);
or U11973 (N_11973,N_11448,N_11110);
or U11974 (N_11974,N_11076,N_11455);
or U11975 (N_11975,N_11125,N_11219);
nor U11976 (N_11976,N_11363,N_11196);
nand U11977 (N_11977,N_11272,N_11425);
xnor U11978 (N_11978,N_11457,N_11392);
xor U11979 (N_11979,N_11034,N_11161);
xnor U11980 (N_11980,N_11067,N_11325);
and U11981 (N_11981,N_11074,N_11213);
xnor U11982 (N_11982,N_11436,N_11295);
xor U11983 (N_11983,N_11167,N_11405);
or U11984 (N_11984,N_11296,N_11064);
and U11985 (N_11985,N_11315,N_11448);
or U11986 (N_11986,N_11274,N_11414);
or U11987 (N_11987,N_11223,N_11460);
and U11988 (N_11988,N_11350,N_11411);
nand U11989 (N_11989,N_11175,N_11053);
or U11990 (N_11990,N_11188,N_11487);
nor U11991 (N_11991,N_11267,N_11250);
and U11992 (N_11992,N_11052,N_11183);
nand U11993 (N_11993,N_11492,N_11180);
and U11994 (N_11994,N_11233,N_11252);
nor U11995 (N_11995,N_11285,N_11276);
and U11996 (N_11996,N_11422,N_11291);
and U11997 (N_11997,N_11274,N_11022);
and U11998 (N_11998,N_11330,N_11408);
xor U11999 (N_11999,N_11389,N_11140);
or U12000 (N_12000,N_11977,N_11557);
nand U12001 (N_12001,N_11582,N_11518);
nor U12002 (N_12002,N_11645,N_11816);
xor U12003 (N_12003,N_11549,N_11906);
nor U12004 (N_12004,N_11693,N_11605);
xnor U12005 (N_12005,N_11710,N_11677);
or U12006 (N_12006,N_11650,N_11587);
and U12007 (N_12007,N_11546,N_11961);
nor U12008 (N_12008,N_11809,N_11715);
xnor U12009 (N_12009,N_11731,N_11827);
or U12010 (N_12010,N_11661,N_11714);
xor U12011 (N_12011,N_11717,N_11740);
xor U12012 (N_12012,N_11843,N_11959);
or U12013 (N_12013,N_11745,N_11849);
nand U12014 (N_12014,N_11613,N_11761);
and U12015 (N_12015,N_11951,N_11531);
or U12016 (N_12016,N_11874,N_11835);
or U12017 (N_12017,N_11929,N_11644);
xnor U12018 (N_12018,N_11727,N_11628);
nor U12019 (N_12019,N_11797,N_11592);
nand U12020 (N_12020,N_11668,N_11830);
or U12021 (N_12021,N_11947,N_11516);
and U12022 (N_12022,N_11735,N_11764);
nor U12023 (N_12023,N_11692,N_11974);
or U12024 (N_12024,N_11982,N_11919);
or U12025 (N_12025,N_11676,N_11918);
nand U12026 (N_12026,N_11954,N_11716);
and U12027 (N_12027,N_11766,N_11739);
nor U12028 (N_12028,N_11870,N_11752);
xor U12029 (N_12029,N_11725,N_11864);
or U12030 (N_12030,N_11704,N_11780);
xor U12031 (N_12031,N_11858,N_11878);
xnor U12032 (N_12032,N_11850,N_11633);
nand U12033 (N_12033,N_11896,N_11622);
or U12034 (N_12034,N_11544,N_11917);
nor U12035 (N_12035,N_11892,N_11523);
and U12036 (N_12036,N_11563,N_11660);
nor U12037 (N_12037,N_11672,N_11762);
nand U12038 (N_12038,N_11823,N_11980);
and U12039 (N_12039,N_11701,N_11979);
nor U12040 (N_12040,N_11552,N_11756);
xor U12041 (N_12041,N_11769,N_11584);
or U12042 (N_12042,N_11742,N_11926);
or U12043 (N_12043,N_11601,N_11839);
and U12044 (N_12044,N_11653,N_11884);
and U12045 (N_12045,N_11876,N_11519);
xor U12046 (N_12046,N_11834,N_11734);
and U12047 (N_12047,N_11948,N_11925);
xnor U12048 (N_12048,N_11726,N_11807);
nand U12049 (N_12049,N_11685,N_11895);
nand U12050 (N_12050,N_11658,N_11547);
or U12051 (N_12051,N_11792,N_11664);
nor U12052 (N_12052,N_11789,N_11565);
nor U12053 (N_12053,N_11504,N_11524);
xnor U12054 (N_12054,N_11875,N_11686);
or U12055 (N_12055,N_11904,N_11617);
or U12056 (N_12056,N_11619,N_11998);
nor U12057 (N_12057,N_11551,N_11750);
nor U12058 (N_12058,N_11942,N_11890);
nand U12059 (N_12059,N_11675,N_11515);
or U12060 (N_12060,N_11817,N_11651);
or U12061 (N_12061,N_11641,N_11699);
xnor U12062 (N_12062,N_11831,N_11674);
or U12063 (N_12063,N_11879,N_11861);
xor U12064 (N_12064,N_11970,N_11513);
xnor U12065 (N_12065,N_11869,N_11665);
xor U12066 (N_12066,N_11541,N_11682);
or U12067 (N_12067,N_11567,N_11581);
and U12068 (N_12068,N_11569,N_11845);
and U12069 (N_12069,N_11743,N_11841);
nand U12070 (N_12070,N_11548,N_11796);
or U12071 (N_12071,N_11818,N_11754);
xor U12072 (N_12072,N_11590,N_11678);
or U12073 (N_12073,N_11775,N_11732);
nor U12074 (N_12074,N_11991,N_11700);
and U12075 (N_12075,N_11744,N_11785);
or U12076 (N_12076,N_11530,N_11673);
or U12077 (N_12077,N_11848,N_11705);
xnor U12078 (N_12078,N_11642,N_11736);
nor U12079 (N_12079,N_11969,N_11814);
nor U12080 (N_12080,N_11570,N_11810);
nor U12081 (N_12081,N_11684,N_11966);
xnor U12082 (N_12082,N_11934,N_11965);
and U12083 (N_12083,N_11938,N_11773);
or U12084 (N_12084,N_11638,N_11707);
or U12085 (N_12085,N_11671,N_11542);
and U12086 (N_12086,N_11772,N_11598);
and U12087 (N_12087,N_11629,N_11709);
nand U12088 (N_12088,N_11564,N_11595);
and U12089 (N_12089,N_11536,N_11865);
or U12090 (N_12090,N_11972,N_11688);
xor U12091 (N_12091,N_11526,N_11822);
or U12092 (N_12092,N_11903,N_11691);
or U12093 (N_12093,N_11657,N_11503);
xnor U12094 (N_12094,N_11939,N_11631);
and U12095 (N_12095,N_11930,N_11507);
and U12096 (N_12096,N_11973,N_11680);
xnor U12097 (N_12097,N_11958,N_11620);
and U12098 (N_12098,N_11637,N_11801);
or U12099 (N_12099,N_11888,N_11517);
nand U12100 (N_12100,N_11602,N_11640);
nor U12101 (N_12101,N_11683,N_11609);
xnor U12102 (N_12102,N_11522,N_11989);
nor U12103 (N_12103,N_11920,N_11558);
and U12104 (N_12104,N_11813,N_11828);
nand U12105 (N_12105,N_11616,N_11799);
or U12106 (N_12106,N_11885,N_11837);
xnor U12107 (N_12107,N_11936,N_11997);
or U12108 (N_12108,N_11514,N_11916);
and U12109 (N_12109,N_11774,N_11795);
nor U12110 (N_12110,N_11832,N_11990);
xnor U12111 (N_12111,N_11776,N_11603);
and U12112 (N_12112,N_11634,N_11535);
or U12113 (N_12113,N_11778,N_11931);
nand U12114 (N_12114,N_11912,N_11612);
and U12115 (N_12115,N_11525,N_11532);
xnor U12116 (N_12116,N_11953,N_11679);
nand U12117 (N_12117,N_11550,N_11655);
and U12118 (N_12118,N_11950,N_11741);
xor U12119 (N_12119,N_11844,N_11749);
nand U12120 (N_12120,N_11600,N_11747);
or U12121 (N_12121,N_11702,N_11967);
and U12122 (N_12122,N_11527,N_11815);
and U12123 (N_12123,N_11505,N_11654);
or U12124 (N_12124,N_11868,N_11593);
nand U12125 (N_12125,N_11572,N_11511);
and U12126 (N_12126,N_11730,N_11933);
nor U12127 (N_12127,N_11763,N_11838);
and U12128 (N_12128,N_11639,N_11591);
nand U12129 (N_12129,N_11922,N_11806);
nand U12130 (N_12130,N_11647,N_11502);
and U12131 (N_12131,N_11706,N_11720);
nand U12132 (N_12132,N_11757,N_11580);
nor U12133 (N_12133,N_11893,N_11994);
nand U12134 (N_12134,N_11553,N_11538);
and U12135 (N_12135,N_11646,N_11826);
and U12136 (N_12136,N_11694,N_11891);
xnor U12137 (N_12137,N_11910,N_11908);
or U12138 (N_12138,N_11625,N_11777);
nand U12139 (N_12139,N_11539,N_11872);
xor U12140 (N_12140,N_11941,N_11871);
nor U12141 (N_12141,N_11956,N_11652);
and U12142 (N_12142,N_11798,N_11556);
xnor U12143 (N_12143,N_11555,N_11880);
nor U12144 (N_12144,N_11887,N_11574);
xor U12145 (N_12145,N_11636,N_11867);
nand U12146 (N_12146,N_11981,N_11537);
or U12147 (N_12147,N_11689,N_11854);
nor U12148 (N_12148,N_11696,N_11968);
and U12149 (N_12149,N_11765,N_11862);
and U12150 (N_12150,N_11554,N_11669);
nand U12151 (N_12151,N_11794,N_11866);
nand U12152 (N_12152,N_11976,N_11729);
nand U12153 (N_12153,N_11984,N_11886);
nand U12154 (N_12154,N_11578,N_11803);
nor U12155 (N_12155,N_11690,N_11963);
or U12156 (N_12156,N_11898,N_11728);
xor U12157 (N_12157,N_11995,N_11955);
nand U12158 (N_12158,N_11852,N_11945);
nand U12159 (N_12159,N_11779,N_11860);
and U12160 (N_12160,N_11708,N_11566);
nand U12161 (N_12161,N_11562,N_11975);
nor U12162 (N_12162,N_11604,N_11666);
nand U12163 (N_12163,N_11855,N_11847);
or U12164 (N_12164,N_11506,N_11545);
or U12165 (N_12165,N_11944,N_11533);
xnor U12166 (N_12166,N_11851,N_11663);
and U12167 (N_12167,N_11840,N_11579);
nor U12168 (N_12168,N_11643,N_11594);
nor U12169 (N_12169,N_11615,N_11649);
nor U12170 (N_12170,N_11577,N_11996);
nor U12171 (N_12171,N_11882,N_11771);
and U12172 (N_12172,N_11993,N_11923);
nor U12173 (N_12173,N_11836,N_11829);
nand U12174 (N_12174,N_11897,N_11820);
and U12175 (N_12175,N_11586,N_11819);
or U12176 (N_12176,N_11711,N_11811);
xnor U12177 (N_12177,N_11733,N_11859);
and U12178 (N_12178,N_11568,N_11724);
or U12179 (N_12179,N_11928,N_11500);
or U12180 (N_12180,N_11627,N_11783);
nor U12181 (N_12181,N_11755,N_11738);
xor U12182 (N_12182,N_11805,N_11821);
and U12183 (N_12183,N_11846,N_11589);
xor U12184 (N_12184,N_11790,N_11662);
or U12185 (N_12185,N_11781,N_11902);
nor U12186 (N_12186,N_11608,N_11753);
and U12187 (N_12187,N_11949,N_11804);
and U12188 (N_12188,N_11667,N_11964);
nand U12189 (N_12189,N_11812,N_11787);
xor U12190 (N_12190,N_11758,N_11983);
nor U12191 (N_12191,N_11863,N_11784);
nand U12192 (N_12192,N_11857,N_11632);
and U12193 (N_12193,N_11712,N_11509);
or U12194 (N_12194,N_11960,N_11978);
nor U12195 (N_12195,N_11681,N_11927);
or U12196 (N_12196,N_11881,N_11824);
and U12197 (N_12197,N_11610,N_11883);
nor U12198 (N_12198,N_11611,N_11915);
and U12199 (N_12199,N_11992,N_11946);
or U12200 (N_12200,N_11521,N_11924);
xnor U12201 (N_12201,N_11529,N_11659);
or U12202 (N_12202,N_11943,N_11914);
or U12203 (N_12203,N_11648,N_11833);
xnor U12204 (N_12204,N_11767,N_11697);
and U12205 (N_12205,N_11842,N_11971);
nand U12206 (N_12206,N_11957,N_11932);
xor U12207 (N_12207,N_11560,N_11687);
nor U12208 (N_12208,N_11585,N_11999);
nor U12209 (N_12209,N_11656,N_11800);
xnor U12210 (N_12210,N_11900,N_11623);
xnor U12211 (N_12211,N_11907,N_11721);
xor U12212 (N_12212,N_11751,N_11528);
nor U12213 (N_12213,N_11559,N_11508);
nor U12214 (N_12214,N_11759,N_11635);
and U12215 (N_12215,N_11940,N_11962);
nor U12216 (N_12216,N_11913,N_11695);
nand U12217 (N_12217,N_11520,N_11873);
nand U12218 (N_12218,N_11737,N_11576);
nand U12219 (N_12219,N_11540,N_11596);
nand U12220 (N_12220,N_11614,N_11588);
and U12221 (N_12221,N_11808,N_11768);
nand U12222 (N_12222,N_11985,N_11786);
nor U12223 (N_12223,N_11952,N_11573);
or U12224 (N_12224,N_11899,N_11782);
nor U12225 (N_12225,N_11760,N_11791);
and U12226 (N_12226,N_11856,N_11510);
or U12227 (N_12227,N_11698,N_11988);
nor U12228 (N_12228,N_11561,N_11606);
or U12229 (N_12229,N_11624,N_11986);
and U12230 (N_12230,N_11599,N_11853);
nor U12231 (N_12231,N_11802,N_11543);
nor U12232 (N_12232,N_11618,N_11770);
and U12233 (N_12233,N_11703,N_11901);
and U12234 (N_12234,N_11723,N_11583);
xnor U12235 (N_12235,N_11746,N_11921);
nand U12236 (N_12236,N_11713,N_11607);
or U12237 (N_12237,N_11905,N_11718);
xnor U12238 (N_12238,N_11825,N_11793);
xor U12239 (N_12239,N_11626,N_11877);
and U12240 (N_12240,N_11935,N_11894);
nor U12241 (N_12241,N_11571,N_11501);
nor U12242 (N_12242,N_11512,N_11575);
nand U12243 (N_12243,N_11621,N_11670);
and U12244 (N_12244,N_11630,N_11889);
xnor U12245 (N_12245,N_11597,N_11911);
or U12246 (N_12246,N_11722,N_11748);
or U12247 (N_12247,N_11987,N_11788);
and U12248 (N_12248,N_11909,N_11719);
and U12249 (N_12249,N_11534,N_11937);
and U12250 (N_12250,N_11688,N_11862);
and U12251 (N_12251,N_11837,N_11758);
and U12252 (N_12252,N_11524,N_11906);
nor U12253 (N_12253,N_11849,N_11972);
xor U12254 (N_12254,N_11544,N_11640);
or U12255 (N_12255,N_11778,N_11782);
and U12256 (N_12256,N_11852,N_11508);
nor U12257 (N_12257,N_11959,N_11635);
nor U12258 (N_12258,N_11598,N_11508);
nand U12259 (N_12259,N_11735,N_11721);
nand U12260 (N_12260,N_11941,N_11847);
or U12261 (N_12261,N_11741,N_11914);
nand U12262 (N_12262,N_11844,N_11804);
nand U12263 (N_12263,N_11773,N_11811);
and U12264 (N_12264,N_11719,N_11758);
or U12265 (N_12265,N_11794,N_11907);
and U12266 (N_12266,N_11645,N_11541);
xnor U12267 (N_12267,N_11602,N_11502);
or U12268 (N_12268,N_11945,N_11642);
or U12269 (N_12269,N_11607,N_11649);
nor U12270 (N_12270,N_11902,N_11634);
nor U12271 (N_12271,N_11794,N_11639);
xor U12272 (N_12272,N_11951,N_11730);
or U12273 (N_12273,N_11844,N_11554);
and U12274 (N_12274,N_11546,N_11621);
nand U12275 (N_12275,N_11774,N_11845);
and U12276 (N_12276,N_11963,N_11520);
nor U12277 (N_12277,N_11919,N_11546);
or U12278 (N_12278,N_11645,N_11867);
xnor U12279 (N_12279,N_11591,N_11503);
or U12280 (N_12280,N_11676,N_11525);
nand U12281 (N_12281,N_11913,N_11801);
xor U12282 (N_12282,N_11606,N_11508);
xor U12283 (N_12283,N_11650,N_11986);
and U12284 (N_12284,N_11922,N_11690);
or U12285 (N_12285,N_11874,N_11637);
xnor U12286 (N_12286,N_11977,N_11514);
and U12287 (N_12287,N_11512,N_11884);
nand U12288 (N_12288,N_11899,N_11767);
nand U12289 (N_12289,N_11802,N_11781);
or U12290 (N_12290,N_11669,N_11756);
nor U12291 (N_12291,N_11951,N_11852);
and U12292 (N_12292,N_11902,N_11630);
and U12293 (N_12293,N_11576,N_11864);
xor U12294 (N_12294,N_11969,N_11819);
or U12295 (N_12295,N_11580,N_11674);
and U12296 (N_12296,N_11754,N_11931);
or U12297 (N_12297,N_11725,N_11996);
nor U12298 (N_12298,N_11919,N_11774);
and U12299 (N_12299,N_11691,N_11626);
nand U12300 (N_12300,N_11749,N_11912);
and U12301 (N_12301,N_11880,N_11962);
or U12302 (N_12302,N_11577,N_11977);
nor U12303 (N_12303,N_11934,N_11695);
xnor U12304 (N_12304,N_11666,N_11702);
nor U12305 (N_12305,N_11954,N_11506);
and U12306 (N_12306,N_11990,N_11676);
nor U12307 (N_12307,N_11659,N_11716);
or U12308 (N_12308,N_11689,N_11676);
nor U12309 (N_12309,N_11696,N_11541);
xor U12310 (N_12310,N_11588,N_11801);
nor U12311 (N_12311,N_11526,N_11837);
nor U12312 (N_12312,N_11792,N_11590);
nand U12313 (N_12313,N_11628,N_11631);
or U12314 (N_12314,N_11842,N_11954);
and U12315 (N_12315,N_11843,N_11886);
or U12316 (N_12316,N_11524,N_11566);
or U12317 (N_12317,N_11684,N_11788);
nand U12318 (N_12318,N_11516,N_11845);
or U12319 (N_12319,N_11716,N_11801);
xnor U12320 (N_12320,N_11890,N_11947);
or U12321 (N_12321,N_11942,N_11973);
xor U12322 (N_12322,N_11959,N_11510);
nand U12323 (N_12323,N_11975,N_11824);
and U12324 (N_12324,N_11682,N_11649);
nor U12325 (N_12325,N_11814,N_11670);
and U12326 (N_12326,N_11955,N_11885);
xor U12327 (N_12327,N_11529,N_11856);
and U12328 (N_12328,N_11900,N_11743);
nor U12329 (N_12329,N_11895,N_11673);
and U12330 (N_12330,N_11743,N_11903);
xnor U12331 (N_12331,N_11965,N_11874);
and U12332 (N_12332,N_11915,N_11788);
xor U12333 (N_12333,N_11569,N_11640);
and U12334 (N_12334,N_11750,N_11586);
or U12335 (N_12335,N_11920,N_11503);
xor U12336 (N_12336,N_11955,N_11591);
and U12337 (N_12337,N_11853,N_11798);
or U12338 (N_12338,N_11669,N_11882);
xnor U12339 (N_12339,N_11600,N_11502);
xor U12340 (N_12340,N_11573,N_11913);
xor U12341 (N_12341,N_11513,N_11727);
or U12342 (N_12342,N_11579,N_11540);
nor U12343 (N_12343,N_11750,N_11759);
nor U12344 (N_12344,N_11991,N_11822);
xor U12345 (N_12345,N_11533,N_11804);
or U12346 (N_12346,N_11821,N_11658);
nand U12347 (N_12347,N_11577,N_11911);
nor U12348 (N_12348,N_11548,N_11717);
or U12349 (N_12349,N_11750,N_11655);
nand U12350 (N_12350,N_11769,N_11919);
and U12351 (N_12351,N_11609,N_11990);
or U12352 (N_12352,N_11785,N_11712);
xor U12353 (N_12353,N_11951,N_11855);
xnor U12354 (N_12354,N_11657,N_11615);
xnor U12355 (N_12355,N_11652,N_11546);
or U12356 (N_12356,N_11530,N_11728);
and U12357 (N_12357,N_11887,N_11680);
nor U12358 (N_12358,N_11725,N_11812);
or U12359 (N_12359,N_11625,N_11903);
xor U12360 (N_12360,N_11730,N_11981);
and U12361 (N_12361,N_11564,N_11796);
or U12362 (N_12362,N_11521,N_11647);
nor U12363 (N_12363,N_11737,N_11913);
nand U12364 (N_12364,N_11871,N_11900);
nand U12365 (N_12365,N_11764,N_11747);
nand U12366 (N_12366,N_11698,N_11589);
xor U12367 (N_12367,N_11698,N_11642);
or U12368 (N_12368,N_11935,N_11722);
nand U12369 (N_12369,N_11782,N_11909);
xor U12370 (N_12370,N_11989,N_11822);
nand U12371 (N_12371,N_11517,N_11724);
nor U12372 (N_12372,N_11945,N_11807);
xor U12373 (N_12373,N_11542,N_11593);
and U12374 (N_12374,N_11697,N_11584);
xnor U12375 (N_12375,N_11503,N_11573);
or U12376 (N_12376,N_11849,N_11660);
xnor U12377 (N_12377,N_11953,N_11579);
nand U12378 (N_12378,N_11670,N_11759);
or U12379 (N_12379,N_11976,N_11954);
xor U12380 (N_12380,N_11603,N_11848);
nor U12381 (N_12381,N_11917,N_11923);
nand U12382 (N_12382,N_11850,N_11558);
xor U12383 (N_12383,N_11659,N_11971);
nand U12384 (N_12384,N_11964,N_11587);
nor U12385 (N_12385,N_11747,N_11561);
and U12386 (N_12386,N_11596,N_11622);
nand U12387 (N_12387,N_11725,N_11665);
xor U12388 (N_12388,N_11726,N_11895);
or U12389 (N_12389,N_11960,N_11815);
nor U12390 (N_12390,N_11885,N_11847);
nor U12391 (N_12391,N_11835,N_11909);
or U12392 (N_12392,N_11954,N_11688);
nor U12393 (N_12393,N_11692,N_11557);
nand U12394 (N_12394,N_11892,N_11810);
and U12395 (N_12395,N_11733,N_11520);
xnor U12396 (N_12396,N_11899,N_11952);
nand U12397 (N_12397,N_11754,N_11822);
or U12398 (N_12398,N_11800,N_11651);
or U12399 (N_12399,N_11866,N_11670);
or U12400 (N_12400,N_11536,N_11521);
and U12401 (N_12401,N_11858,N_11922);
and U12402 (N_12402,N_11732,N_11796);
nor U12403 (N_12403,N_11604,N_11945);
or U12404 (N_12404,N_11716,N_11601);
and U12405 (N_12405,N_11889,N_11519);
or U12406 (N_12406,N_11685,N_11620);
xnor U12407 (N_12407,N_11960,N_11768);
or U12408 (N_12408,N_11944,N_11806);
nor U12409 (N_12409,N_11857,N_11965);
nor U12410 (N_12410,N_11607,N_11528);
nand U12411 (N_12411,N_11608,N_11634);
and U12412 (N_12412,N_11663,N_11801);
nor U12413 (N_12413,N_11800,N_11726);
and U12414 (N_12414,N_11744,N_11981);
and U12415 (N_12415,N_11500,N_11737);
and U12416 (N_12416,N_11993,N_11559);
or U12417 (N_12417,N_11554,N_11994);
xor U12418 (N_12418,N_11797,N_11838);
nor U12419 (N_12419,N_11608,N_11919);
and U12420 (N_12420,N_11764,N_11561);
xor U12421 (N_12421,N_11986,N_11763);
and U12422 (N_12422,N_11816,N_11965);
or U12423 (N_12423,N_11560,N_11774);
xnor U12424 (N_12424,N_11580,N_11623);
xnor U12425 (N_12425,N_11917,N_11586);
nand U12426 (N_12426,N_11588,N_11823);
or U12427 (N_12427,N_11702,N_11905);
and U12428 (N_12428,N_11565,N_11535);
and U12429 (N_12429,N_11579,N_11549);
nor U12430 (N_12430,N_11555,N_11615);
or U12431 (N_12431,N_11601,N_11703);
nand U12432 (N_12432,N_11948,N_11814);
or U12433 (N_12433,N_11772,N_11579);
nand U12434 (N_12434,N_11713,N_11626);
or U12435 (N_12435,N_11838,N_11734);
or U12436 (N_12436,N_11693,N_11881);
nand U12437 (N_12437,N_11730,N_11953);
and U12438 (N_12438,N_11770,N_11813);
nor U12439 (N_12439,N_11564,N_11925);
and U12440 (N_12440,N_11716,N_11672);
or U12441 (N_12441,N_11881,N_11870);
xor U12442 (N_12442,N_11653,N_11984);
nand U12443 (N_12443,N_11724,N_11995);
or U12444 (N_12444,N_11790,N_11885);
or U12445 (N_12445,N_11602,N_11671);
xnor U12446 (N_12446,N_11807,N_11846);
and U12447 (N_12447,N_11759,N_11788);
xnor U12448 (N_12448,N_11624,N_11655);
xor U12449 (N_12449,N_11597,N_11821);
nor U12450 (N_12450,N_11690,N_11651);
nand U12451 (N_12451,N_11849,N_11595);
nand U12452 (N_12452,N_11561,N_11621);
nor U12453 (N_12453,N_11654,N_11708);
or U12454 (N_12454,N_11701,N_11587);
and U12455 (N_12455,N_11612,N_11582);
or U12456 (N_12456,N_11949,N_11519);
nor U12457 (N_12457,N_11984,N_11943);
or U12458 (N_12458,N_11898,N_11809);
or U12459 (N_12459,N_11594,N_11625);
or U12460 (N_12460,N_11521,N_11510);
xnor U12461 (N_12461,N_11672,N_11882);
and U12462 (N_12462,N_11935,N_11537);
xnor U12463 (N_12463,N_11932,N_11782);
nor U12464 (N_12464,N_11548,N_11789);
nand U12465 (N_12465,N_11644,N_11892);
nor U12466 (N_12466,N_11753,N_11614);
and U12467 (N_12467,N_11663,N_11860);
nand U12468 (N_12468,N_11869,N_11597);
nand U12469 (N_12469,N_11532,N_11911);
xor U12470 (N_12470,N_11679,N_11894);
xnor U12471 (N_12471,N_11522,N_11500);
xnor U12472 (N_12472,N_11503,N_11604);
nor U12473 (N_12473,N_11654,N_11516);
xor U12474 (N_12474,N_11630,N_11780);
nand U12475 (N_12475,N_11776,N_11905);
nor U12476 (N_12476,N_11771,N_11997);
nand U12477 (N_12477,N_11715,N_11944);
and U12478 (N_12478,N_11656,N_11671);
nand U12479 (N_12479,N_11963,N_11784);
or U12480 (N_12480,N_11814,N_11583);
nor U12481 (N_12481,N_11520,N_11766);
and U12482 (N_12482,N_11697,N_11619);
nand U12483 (N_12483,N_11937,N_11525);
nand U12484 (N_12484,N_11578,N_11668);
nor U12485 (N_12485,N_11870,N_11913);
nand U12486 (N_12486,N_11532,N_11999);
and U12487 (N_12487,N_11856,N_11610);
nand U12488 (N_12488,N_11982,N_11679);
and U12489 (N_12489,N_11762,N_11950);
nand U12490 (N_12490,N_11666,N_11904);
xnor U12491 (N_12491,N_11736,N_11765);
and U12492 (N_12492,N_11954,N_11822);
and U12493 (N_12493,N_11592,N_11684);
nor U12494 (N_12494,N_11999,N_11578);
and U12495 (N_12495,N_11845,N_11836);
and U12496 (N_12496,N_11958,N_11652);
nand U12497 (N_12497,N_11656,N_11922);
nand U12498 (N_12498,N_11617,N_11770);
xor U12499 (N_12499,N_11649,N_11856);
or U12500 (N_12500,N_12058,N_12024);
nand U12501 (N_12501,N_12463,N_12198);
xnor U12502 (N_12502,N_12216,N_12369);
nor U12503 (N_12503,N_12037,N_12021);
nand U12504 (N_12504,N_12049,N_12084);
xnor U12505 (N_12505,N_12493,N_12467);
xnor U12506 (N_12506,N_12470,N_12047);
and U12507 (N_12507,N_12119,N_12337);
or U12508 (N_12508,N_12309,N_12341);
and U12509 (N_12509,N_12320,N_12067);
and U12510 (N_12510,N_12459,N_12453);
xnor U12511 (N_12511,N_12207,N_12436);
xor U12512 (N_12512,N_12439,N_12231);
xor U12513 (N_12513,N_12124,N_12315);
and U12514 (N_12514,N_12193,N_12053);
or U12515 (N_12515,N_12336,N_12062);
nor U12516 (N_12516,N_12005,N_12095);
nand U12517 (N_12517,N_12134,N_12013);
nor U12518 (N_12518,N_12178,N_12366);
xnor U12519 (N_12519,N_12399,N_12461);
or U12520 (N_12520,N_12370,N_12474);
nand U12521 (N_12521,N_12215,N_12057);
or U12522 (N_12522,N_12250,N_12044);
nor U12523 (N_12523,N_12194,N_12290);
or U12524 (N_12524,N_12222,N_12078);
nor U12525 (N_12525,N_12238,N_12322);
and U12526 (N_12526,N_12196,N_12180);
nor U12527 (N_12527,N_12043,N_12432);
nand U12528 (N_12528,N_12495,N_12425);
nand U12529 (N_12529,N_12148,N_12170);
nand U12530 (N_12530,N_12421,N_12131);
or U12531 (N_12531,N_12318,N_12045);
nor U12532 (N_12532,N_12168,N_12055);
or U12533 (N_12533,N_12208,N_12423);
and U12534 (N_12534,N_12165,N_12099);
nor U12535 (N_12535,N_12275,N_12481);
and U12536 (N_12536,N_12116,N_12327);
nand U12537 (N_12537,N_12257,N_12025);
nand U12538 (N_12538,N_12225,N_12262);
nor U12539 (N_12539,N_12303,N_12412);
xnor U12540 (N_12540,N_12097,N_12073);
nor U12541 (N_12541,N_12172,N_12301);
nand U12542 (N_12542,N_12200,N_12100);
nand U12543 (N_12543,N_12496,N_12085);
nor U12544 (N_12544,N_12107,N_12307);
nand U12545 (N_12545,N_12071,N_12205);
or U12546 (N_12546,N_12312,N_12498);
nor U12547 (N_12547,N_12380,N_12145);
nand U12548 (N_12548,N_12104,N_12343);
xnor U12549 (N_12549,N_12183,N_12296);
and U12550 (N_12550,N_12008,N_12373);
nor U12551 (N_12551,N_12326,N_12305);
xor U12552 (N_12552,N_12035,N_12036);
or U12553 (N_12553,N_12435,N_12192);
or U12554 (N_12554,N_12394,N_12235);
or U12555 (N_12555,N_12228,N_12219);
nand U12556 (N_12556,N_12471,N_12094);
nor U12557 (N_12557,N_12065,N_12454);
nor U12558 (N_12558,N_12427,N_12297);
xnor U12559 (N_12559,N_12022,N_12018);
nor U12560 (N_12560,N_12384,N_12351);
and U12561 (N_12561,N_12147,N_12137);
or U12562 (N_12562,N_12347,N_12114);
and U12563 (N_12563,N_12087,N_12237);
nand U12564 (N_12564,N_12151,N_12437);
and U12565 (N_12565,N_12382,N_12082);
and U12566 (N_12566,N_12484,N_12141);
xor U12567 (N_12567,N_12175,N_12034);
or U12568 (N_12568,N_12408,N_12265);
and U12569 (N_12569,N_12346,N_12450);
xnor U12570 (N_12570,N_12039,N_12052);
nor U12571 (N_12571,N_12383,N_12187);
or U12572 (N_12572,N_12203,N_12096);
nor U12573 (N_12573,N_12294,N_12110);
xor U12574 (N_12574,N_12077,N_12186);
or U12575 (N_12575,N_12224,N_12433);
or U12576 (N_12576,N_12229,N_12368);
and U12577 (N_12577,N_12393,N_12146);
and U12578 (N_12578,N_12121,N_12251);
nor U12579 (N_12579,N_12163,N_12051);
or U12580 (N_12580,N_12418,N_12009);
xor U12581 (N_12581,N_12220,N_12092);
nor U12582 (N_12582,N_12190,N_12345);
or U12583 (N_12583,N_12029,N_12348);
and U12584 (N_12584,N_12046,N_12266);
and U12585 (N_12585,N_12001,N_12226);
nor U12586 (N_12586,N_12469,N_12388);
nand U12587 (N_12587,N_12404,N_12031);
xnor U12588 (N_12588,N_12491,N_12431);
nand U12589 (N_12589,N_12221,N_12392);
nand U12590 (N_12590,N_12189,N_12456);
xnor U12591 (N_12591,N_12160,N_12492);
and U12592 (N_12592,N_12117,N_12111);
xnor U12593 (N_12593,N_12448,N_12455);
nor U12594 (N_12594,N_12422,N_12335);
or U12595 (N_12595,N_12443,N_12245);
nor U12596 (N_12596,N_12088,N_12365);
nand U12597 (N_12597,N_12473,N_12376);
xnor U12598 (N_12598,N_12386,N_12342);
nor U12599 (N_12599,N_12156,N_12329);
nand U12600 (N_12600,N_12089,N_12304);
xnor U12601 (N_12601,N_12179,N_12390);
xor U12602 (N_12602,N_12401,N_12164);
or U12603 (N_12603,N_12234,N_12494);
xor U12604 (N_12604,N_12015,N_12325);
or U12605 (N_12605,N_12478,N_12441);
or U12606 (N_12606,N_12387,N_12197);
or U12607 (N_12607,N_12103,N_12379);
xnor U12608 (N_12608,N_12123,N_12214);
xor U12609 (N_12609,N_12472,N_12217);
or U12610 (N_12610,N_12218,N_12069);
xor U12611 (N_12611,N_12310,N_12158);
nor U12612 (N_12612,N_12152,N_12352);
xor U12613 (N_12613,N_12182,N_12264);
nand U12614 (N_12614,N_12210,N_12483);
nand U12615 (N_12615,N_12113,N_12277);
nor U12616 (N_12616,N_12091,N_12149);
nand U12617 (N_12617,N_12201,N_12293);
xnor U12618 (N_12618,N_12389,N_12497);
and U12619 (N_12619,N_12012,N_12188);
nand U12620 (N_12620,N_12402,N_12291);
nand U12621 (N_12621,N_12153,N_12283);
nor U12622 (N_12622,N_12490,N_12256);
nand U12623 (N_12623,N_12429,N_12177);
xnor U12624 (N_12624,N_12269,N_12438);
or U12625 (N_12625,N_12048,N_12199);
nand U12626 (N_12626,N_12072,N_12068);
and U12627 (N_12627,N_12406,N_12233);
nor U12628 (N_12628,N_12236,N_12263);
or U12629 (N_12629,N_12122,N_12241);
nor U12630 (N_12630,N_12460,N_12059);
xnor U12631 (N_12631,N_12367,N_12061);
nand U12632 (N_12632,N_12129,N_12362);
or U12633 (N_12633,N_12167,N_12360);
xnor U12634 (N_12634,N_12209,N_12133);
nand U12635 (N_12635,N_12157,N_12042);
xnor U12636 (N_12636,N_12181,N_12247);
nor U12637 (N_12637,N_12356,N_12255);
nand U12638 (N_12638,N_12174,N_12298);
and U12639 (N_12639,N_12434,N_12041);
and U12640 (N_12640,N_12244,N_12105);
xnor U12641 (N_12641,N_12249,N_12282);
xnor U12642 (N_12642,N_12017,N_12206);
or U12643 (N_12643,N_12324,N_12391);
nand U12644 (N_12644,N_12344,N_12426);
or U12645 (N_12645,N_12054,N_12279);
and U12646 (N_12646,N_12306,N_12195);
and U12647 (N_12647,N_12419,N_12278);
xor U12648 (N_12648,N_12028,N_12477);
nor U12649 (N_12649,N_12125,N_12020);
nor U12650 (N_12650,N_12011,N_12106);
and U12651 (N_12651,N_12288,N_12440);
or U12652 (N_12652,N_12355,N_12120);
and U12653 (N_12653,N_12004,N_12374);
or U12654 (N_12654,N_12268,N_12359);
xnor U12655 (N_12655,N_12447,N_12444);
xnor U12656 (N_12656,N_12254,N_12098);
xor U12657 (N_12657,N_12138,N_12162);
and U12658 (N_12658,N_12377,N_12284);
nand U12659 (N_12659,N_12246,N_12191);
nor U12660 (N_12660,N_12417,N_12489);
nor U12661 (N_12661,N_12033,N_12010);
xor U12662 (N_12662,N_12060,N_12130);
or U12663 (N_12663,N_12213,N_12185);
nand U12664 (N_12664,N_12300,N_12354);
and U12665 (N_12665,N_12385,N_12211);
or U12666 (N_12666,N_12480,N_12428);
xor U12667 (N_12667,N_12272,N_12023);
nor U12668 (N_12668,N_12006,N_12016);
nor U12669 (N_12669,N_12451,N_12333);
and U12670 (N_12670,N_12398,N_12281);
xor U12671 (N_12671,N_12202,N_12350);
or U12672 (N_12672,N_12108,N_12128);
or U12673 (N_12673,N_12232,N_12287);
and U12674 (N_12674,N_12361,N_12285);
xor U12675 (N_12675,N_12040,N_12349);
nand U12676 (N_12676,N_12499,N_12458);
and U12677 (N_12677,N_12184,N_12323);
xnor U12678 (N_12678,N_12204,N_12364);
nor U12679 (N_12679,N_12169,N_12173);
or U12680 (N_12680,N_12405,N_12430);
xor U12681 (N_12681,N_12446,N_12409);
nand U12682 (N_12682,N_12075,N_12050);
nand U12683 (N_12683,N_12395,N_12413);
xnor U12684 (N_12684,N_12063,N_12081);
xnor U12685 (N_12685,N_12479,N_12295);
xor U12686 (N_12686,N_12248,N_12090);
xnor U12687 (N_12687,N_12136,N_12358);
nor U12688 (N_12688,N_12372,N_12271);
nand U12689 (N_12689,N_12155,N_12452);
nand U12690 (N_12690,N_12259,N_12396);
xnor U12691 (N_12691,N_12118,N_12371);
nor U12692 (N_12692,N_12038,N_12330);
or U12693 (N_12693,N_12115,N_12466);
and U12694 (N_12694,N_12171,N_12242);
xor U12695 (N_12695,N_12258,N_12328);
nand U12696 (N_12696,N_12161,N_12007);
nor U12697 (N_12697,N_12317,N_12411);
nand U12698 (N_12698,N_12101,N_12485);
xnor U12699 (N_12699,N_12019,N_12465);
and U12700 (N_12700,N_12074,N_12449);
or U12701 (N_12701,N_12261,N_12166);
and U12702 (N_12702,N_12286,N_12076);
nand U12703 (N_12703,N_12363,N_12027);
nor U12704 (N_12704,N_12420,N_12002);
and U12705 (N_12705,N_12457,N_12488);
xnor U12706 (N_12706,N_12086,N_12487);
or U12707 (N_12707,N_12482,N_12064);
nand U12708 (N_12708,N_12280,N_12445);
or U12709 (N_12709,N_12292,N_12273);
nand U12710 (N_12710,N_12407,N_12400);
nand U12711 (N_12711,N_12416,N_12338);
nor U12712 (N_12712,N_12003,N_12140);
xnor U12713 (N_12713,N_12302,N_12410);
xnor U12714 (N_12714,N_12132,N_12227);
nand U12715 (N_12715,N_12274,N_12414);
and U12716 (N_12716,N_12313,N_12308);
nor U12717 (N_12717,N_12243,N_12139);
xor U12718 (N_12718,N_12462,N_12464);
or U12719 (N_12719,N_12230,N_12468);
and U12720 (N_12720,N_12154,N_12276);
and U12721 (N_12721,N_12253,N_12334);
nor U12722 (N_12722,N_12311,N_12340);
and U12723 (N_12723,N_12375,N_12331);
xnor U12724 (N_12724,N_12056,N_12403);
nor U12725 (N_12725,N_12357,N_12112);
or U12726 (N_12726,N_12316,N_12442);
xnor U12727 (N_12727,N_12127,N_12321);
and U12728 (N_12728,N_12270,N_12424);
nor U12729 (N_12729,N_12135,N_12176);
nand U12730 (N_12730,N_12397,N_12299);
and U12731 (N_12731,N_12223,N_12030);
or U12732 (N_12732,N_12339,N_12252);
nand U12733 (N_12733,N_12150,N_12289);
xnor U12734 (N_12734,N_12080,N_12319);
and U12735 (N_12735,N_12126,N_12032);
and U12736 (N_12736,N_12332,N_12026);
or U12737 (N_12737,N_12381,N_12415);
xor U12738 (N_12738,N_12353,N_12102);
or U12739 (N_12739,N_12000,N_12142);
and U12740 (N_12740,N_12070,N_12159);
xnor U12741 (N_12741,N_12260,N_12093);
or U12742 (N_12742,N_12079,N_12378);
xnor U12743 (N_12743,N_12267,N_12212);
nand U12744 (N_12744,N_12476,N_12144);
and U12745 (N_12745,N_12083,N_12240);
and U12746 (N_12746,N_12486,N_12066);
xnor U12747 (N_12747,N_12143,N_12239);
or U12748 (N_12748,N_12314,N_12109);
nor U12749 (N_12749,N_12014,N_12475);
or U12750 (N_12750,N_12197,N_12183);
and U12751 (N_12751,N_12025,N_12214);
nand U12752 (N_12752,N_12042,N_12195);
xor U12753 (N_12753,N_12329,N_12084);
and U12754 (N_12754,N_12355,N_12308);
or U12755 (N_12755,N_12449,N_12350);
nand U12756 (N_12756,N_12013,N_12474);
and U12757 (N_12757,N_12454,N_12326);
and U12758 (N_12758,N_12493,N_12241);
nand U12759 (N_12759,N_12389,N_12407);
and U12760 (N_12760,N_12319,N_12352);
and U12761 (N_12761,N_12218,N_12314);
or U12762 (N_12762,N_12344,N_12393);
or U12763 (N_12763,N_12142,N_12460);
nor U12764 (N_12764,N_12061,N_12146);
nand U12765 (N_12765,N_12041,N_12406);
nand U12766 (N_12766,N_12129,N_12119);
or U12767 (N_12767,N_12415,N_12154);
nand U12768 (N_12768,N_12072,N_12262);
and U12769 (N_12769,N_12351,N_12409);
nor U12770 (N_12770,N_12116,N_12167);
xnor U12771 (N_12771,N_12335,N_12170);
nand U12772 (N_12772,N_12333,N_12093);
nand U12773 (N_12773,N_12094,N_12001);
nor U12774 (N_12774,N_12264,N_12314);
nor U12775 (N_12775,N_12287,N_12360);
nor U12776 (N_12776,N_12279,N_12202);
or U12777 (N_12777,N_12210,N_12476);
and U12778 (N_12778,N_12409,N_12018);
nor U12779 (N_12779,N_12202,N_12418);
and U12780 (N_12780,N_12073,N_12187);
nor U12781 (N_12781,N_12226,N_12038);
or U12782 (N_12782,N_12341,N_12455);
xnor U12783 (N_12783,N_12317,N_12414);
xnor U12784 (N_12784,N_12249,N_12015);
nand U12785 (N_12785,N_12326,N_12082);
nand U12786 (N_12786,N_12015,N_12330);
xnor U12787 (N_12787,N_12054,N_12108);
nor U12788 (N_12788,N_12227,N_12072);
and U12789 (N_12789,N_12126,N_12299);
nand U12790 (N_12790,N_12489,N_12283);
nand U12791 (N_12791,N_12191,N_12438);
or U12792 (N_12792,N_12075,N_12341);
or U12793 (N_12793,N_12358,N_12043);
nand U12794 (N_12794,N_12428,N_12406);
nor U12795 (N_12795,N_12443,N_12423);
and U12796 (N_12796,N_12128,N_12230);
or U12797 (N_12797,N_12486,N_12227);
nand U12798 (N_12798,N_12027,N_12148);
xnor U12799 (N_12799,N_12227,N_12049);
nand U12800 (N_12800,N_12368,N_12124);
nor U12801 (N_12801,N_12276,N_12439);
and U12802 (N_12802,N_12279,N_12371);
and U12803 (N_12803,N_12347,N_12111);
xnor U12804 (N_12804,N_12123,N_12010);
nor U12805 (N_12805,N_12094,N_12134);
nand U12806 (N_12806,N_12361,N_12075);
xnor U12807 (N_12807,N_12418,N_12019);
xor U12808 (N_12808,N_12101,N_12228);
and U12809 (N_12809,N_12484,N_12380);
xor U12810 (N_12810,N_12139,N_12249);
or U12811 (N_12811,N_12157,N_12464);
nand U12812 (N_12812,N_12331,N_12104);
and U12813 (N_12813,N_12487,N_12262);
and U12814 (N_12814,N_12390,N_12005);
nand U12815 (N_12815,N_12293,N_12354);
or U12816 (N_12816,N_12128,N_12472);
xor U12817 (N_12817,N_12182,N_12332);
nor U12818 (N_12818,N_12065,N_12344);
xor U12819 (N_12819,N_12063,N_12410);
nor U12820 (N_12820,N_12299,N_12218);
nor U12821 (N_12821,N_12262,N_12397);
or U12822 (N_12822,N_12367,N_12417);
or U12823 (N_12823,N_12159,N_12167);
xor U12824 (N_12824,N_12193,N_12245);
xnor U12825 (N_12825,N_12347,N_12055);
nand U12826 (N_12826,N_12361,N_12181);
and U12827 (N_12827,N_12482,N_12253);
or U12828 (N_12828,N_12067,N_12060);
nand U12829 (N_12829,N_12004,N_12338);
and U12830 (N_12830,N_12184,N_12094);
and U12831 (N_12831,N_12113,N_12149);
xor U12832 (N_12832,N_12444,N_12176);
and U12833 (N_12833,N_12069,N_12003);
nand U12834 (N_12834,N_12015,N_12357);
nor U12835 (N_12835,N_12116,N_12145);
or U12836 (N_12836,N_12470,N_12133);
xnor U12837 (N_12837,N_12144,N_12494);
nor U12838 (N_12838,N_12409,N_12102);
nor U12839 (N_12839,N_12037,N_12126);
and U12840 (N_12840,N_12009,N_12102);
nor U12841 (N_12841,N_12155,N_12246);
nor U12842 (N_12842,N_12329,N_12237);
or U12843 (N_12843,N_12420,N_12424);
nand U12844 (N_12844,N_12001,N_12430);
xor U12845 (N_12845,N_12487,N_12020);
xor U12846 (N_12846,N_12345,N_12072);
or U12847 (N_12847,N_12263,N_12213);
or U12848 (N_12848,N_12054,N_12457);
nand U12849 (N_12849,N_12008,N_12470);
and U12850 (N_12850,N_12346,N_12385);
xor U12851 (N_12851,N_12441,N_12059);
and U12852 (N_12852,N_12402,N_12363);
or U12853 (N_12853,N_12176,N_12158);
xor U12854 (N_12854,N_12129,N_12283);
or U12855 (N_12855,N_12418,N_12067);
or U12856 (N_12856,N_12467,N_12469);
or U12857 (N_12857,N_12348,N_12340);
and U12858 (N_12858,N_12276,N_12190);
xnor U12859 (N_12859,N_12494,N_12076);
and U12860 (N_12860,N_12006,N_12173);
nand U12861 (N_12861,N_12140,N_12489);
xor U12862 (N_12862,N_12384,N_12407);
and U12863 (N_12863,N_12227,N_12168);
or U12864 (N_12864,N_12062,N_12152);
or U12865 (N_12865,N_12065,N_12341);
and U12866 (N_12866,N_12303,N_12400);
and U12867 (N_12867,N_12428,N_12282);
and U12868 (N_12868,N_12315,N_12033);
nor U12869 (N_12869,N_12241,N_12270);
and U12870 (N_12870,N_12309,N_12302);
nor U12871 (N_12871,N_12092,N_12325);
xnor U12872 (N_12872,N_12157,N_12164);
or U12873 (N_12873,N_12336,N_12214);
xnor U12874 (N_12874,N_12007,N_12362);
nor U12875 (N_12875,N_12470,N_12182);
and U12876 (N_12876,N_12367,N_12226);
or U12877 (N_12877,N_12109,N_12377);
nor U12878 (N_12878,N_12449,N_12091);
nor U12879 (N_12879,N_12498,N_12270);
nor U12880 (N_12880,N_12286,N_12484);
or U12881 (N_12881,N_12499,N_12440);
and U12882 (N_12882,N_12293,N_12238);
xnor U12883 (N_12883,N_12188,N_12209);
nor U12884 (N_12884,N_12248,N_12142);
nand U12885 (N_12885,N_12060,N_12038);
and U12886 (N_12886,N_12328,N_12217);
nand U12887 (N_12887,N_12209,N_12359);
nand U12888 (N_12888,N_12312,N_12337);
and U12889 (N_12889,N_12361,N_12053);
nand U12890 (N_12890,N_12485,N_12039);
and U12891 (N_12891,N_12394,N_12261);
or U12892 (N_12892,N_12278,N_12339);
nor U12893 (N_12893,N_12016,N_12317);
and U12894 (N_12894,N_12024,N_12144);
and U12895 (N_12895,N_12323,N_12467);
and U12896 (N_12896,N_12193,N_12380);
and U12897 (N_12897,N_12138,N_12206);
and U12898 (N_12898,N_12175,N_12075);
nand U12899 (N_12899,N_12217,N_12363);
nor U12900 (N_12900,N_12311,N_12418);
and U12901 (N_12901,N_12415,N_12367);
or U12902 (N_12902,N_12407,N_12481);
or U12903 (N_12903,N_12098,N_12195);
nand U12904 (N_12904,N_12455,N_12369);
and U12905 (N_12905,N_12130,N_12380);
nand U12906 (N_12906,N_12433,N_12290);
nor U12907 (N_12907,N_12114,N_12019);
nor U12908 (N_12908,N_12326,N_12179);
nand U12909 (N_12909,N_12018,N_12026);
nand U12910 (N_12910,N_12351,N_12467);
nand U12911 (N_12911,N_12494,N_12052);
and U12912 (N_12912,N_12076,N_12415);
xor U12913 (N_12913,N_12045,N_12031);
and U12914 (N_12914,N_12237,N_12059);
nor U12915 (N_12915,N_12199,N_12107);
xor U12916 (N_12916,N_12133,N_12156);
and U12917 (N_12917,N_12367,N_12387);
xor U12918 (N_12918,N_12145,N_12263);
nor U12919 (N_12919,N_12431,N_12197);
nand U12920 (N_12920,N_12231,N_12380);
xor U12921 (N_12921,N_12141,N_12308);
xor U12922 (N_12922,N_12005,N_12141);
and U12923 (N_12923,N_12181,N_12034);
nor U12924 (N_12924,N_12442,N_12384);
and U12925 (N_12925,N_12077,N_12096);
nand U12926 (N_12926,N_12000,N_12208);
nand U12927 (N_12927,N_12391,N_12422);
or U12928 (N_12928,N_12288,N_12072);
nand U12929 (N_12929,N_12276,N_12246);
nand U12930 (N_12930,N_12028,N_12247);
nor U12931 (N_12931,N_12176,N_12070);
xor U12932 (N_12932,N_12428,N_12117);
or U12933 (N_12933,N_12260,N_12145);
nor U12934 (N_12934,N_12481,N_12227);
xor U12935 (N_12935,N_12486,N_12438);
xor U12936 (N_12936,N_12411,N_12016);
xor U12937 (N_12937,N_12300,N_12381);
and U12938 (N_12938,N_12062,N_12055);
and U12939 (N_12939,N_12249,N_12372);
or U12940 (N_12940,N_12368,N_12181);
nand U12941 (N_12941,N_12316,N_12270);
nor U12942 (N_12942,N_12424,N_12450);
nor U12943 (N_12943,N_12370,N_12468);
xor U12944 (N_12944,N_12039,N_12383);
nor U12945 (N_12945,N_12302,N_12009);
xnor U12946 (N_12946,N_12090,N_12167);
or U12947 (N_12947,N_12186,N_12288);
nand U12948 (N_12948,N_12082,N_12357);
nor U12949 (N_12949,N_12122,N_12176);
nand U12950 (N_12950,N_12438,N_12418);
or U12951 (N_12951,N_12318,N_12339);
xor U12952 (N_12952,N_12316,N_12254);
nand U12953 (N_12953,N_12362,N_12240);
and U12954 (N_12954,N_12341,N_12385);
nor U12955 (N_12955,N_12338,N_12036);
nor U12956 (N_12956,N_12242,N_12403);
xor U12957 (N_12957,N_12209,N_12405);
nor U12958 (N_12958,N_12130,N_12302);
or U12959 (N_12959,N_12385,N_12033);
nor U12960 (N_12960,N_12195,N_12177);
xnor U12961 (N_12961,N_12443,N_12124);
or U12962 (N_12962,N_12312,N_12082);
xnor U12963 (N_12963,N_12223,N_12240);
nor U12964 (N_12964,N_12026,N_12049);
nor U12965 (N_12965,N_12169,N_12098);
xnor U12966 (N_12966,N_12453,N_12394);
xor U12967 (N_12967,N_12111,N_12279);
nor U12968 (N_12968,N_12327,N_12081);
xnor U12969 (N_12969,N_12343,N_12115);
and U12970 (N_12970,N_12480,N_12347);
nor U12971 (N_12971,N_12010,N_12031);
or U12972 (N_12972,N_12267,N_12328);
xor U12973 (N_12973,N_12014,N_12213);
nor U12974 (N_12974,N_12360,N_12482);
or U12975 (N_12975,N_12116,N_12258);
nor U12976 (N_12976,N_12374,N_12367);
nand U12977 (N_12977,N_12236,N_12051);
or U12978 (N_12978,N_12415,N_12009);
nand U12979 (N_12979,N_12371,N_12194);
nor U12980 (N_12980,N_12327,N_12138);
and U12981 (N_12981,N_12073,N_12286);
nor U12982 (N_12982,N_12145,N_12017);
and U12983 (N_12983,N_12046,N_12150);
nor U12984 (N_12984,N_12318,N_12133);
and U12985 (N_12985,N_12314,N_12106);
and U12986 (N_12986,N_12104,N_12405);
and U12987 (N_12987,N_12442,N_12031);
or U12988 (N_12988,N_12260,N_12125);
nand U12989 (N_12989,N_12370,N_12199);
and U12990 (N_12990,N_12089,N_12227);
nand U12991 (N_12991,N_12259,N_12236);
and U12992 (N_12992,N_12231,N_12060);
and U12993 (N_12993,N_12286,N_12240);
xnor U12994 (N_12994,N_12315,N_12186);
xnor U12995 (N_12995,N_12281,N_12163);
or U12996 (N_12996,N_12192,N_12260);
nor U12997 (N_12997,N_12380,N_12211);
nand U12998 (N_12998,N_12011,N_12122);
nor U12999 (N_12999,N_12061,N_12012);
and U13000 (N_13000,N_12710,N_12996);
xnor U13001 (N_13001,N_12883,N_12741);
nor U13002 (N_13002,N_12993,N_12685);
and U13003 (N_13003,N_12540,N_12732);
and U13004 (N_13004,N_12946,N_12785);
and U13005 (N_13005,N_12765,N_12771);
nand U13006 (N_13006,N_12565,N_12523);
nand U13007 (N_13007,N_12768,N_12649);
or U13008 (N_13008,N_12794,N_12812);
xor U13009 (N_13009,N_12893,N_12999);
and U13010 (N_13010,N_12693,N_12642);
nand U13011 (N_13011,N_12778,N_12677);
nor U13012 (N_13012,N_12575,N_12655);
nand U13013 (N_13013,N_12942,N_12774);
xor U13014 (N_13014,N_12604,N_12740);
nor U13015 (N_13015,N_12660,N_12966);
and U13016 (N_13016,N_12998,N_12869);
nand U13017 (N_13017,N_12967,N_12504);
xor U13018 (N_13018,N_12757,N_12628);
xor U13019 (N_13019,N_12758,N_12580);
nor U13020 (N_13020,N_12776,N_12853);
nor U13021 (N_13021,N_12916,N_12514);
or U13022 (N_13022,N_12895,N_12991);
or U13023 (N_13023,N_12703,N_12976);
nor U13024 (N_13024,N_12557,N_12933);
nand U13025 (N_13025,N_12592,N_12688);
xnor U13026 (N_13026,N_12760,N_12657);
nand U13027 (N_13027,N_12558,N_12726);
nand U13028 (N_13028,N_12922,N_12725);
nor U13029 (N_13029,N_12852,N_12746);
or U13030 (N_13030,N_12845,N_12890);
xor U13031 (N_13031,N_12803,N_12879);
xnor U13032 (N_13032,N_12975,N_12682);
nand U13033 (N_13033,N_12616,N_12752);
xor U13034 (N_13034,N_12730,N_12738);
or U13035 (N_13035,N_12934,N_12526);
and U13036 (N_13036,N_12601,N_12903);
nand U13037 (N_13037,N_12536,N_12638);
xnor U13038 (N_13038,N_12925,N_12500);
nor U13039 (N_13039,N_12621,N_12539);
or U13040 (N_13040,N_12817,N_12722);
nor U13041 (N_13041,N_12992,N_12661);
and U13042 (N_13042,N_12945,N_12714);
nor U13043 (N_13043,N_12844,N_12995);
and U13044 (N_13044,N_12786,N_12915);
nor U13045 (N_13045,N_12877,N_12856);
or U13046 (N_13046,N_12961,N_12985);
xnor U13047 (N_13047,N_12653,N_12644);
and U13048 (N_13048,N_12633,N_12931);
xnor U13049 (N_13049,N_12764,N_12582);
or U13050 (N_13050,N_12734,N_12891);
and U13051 (N_13051,N_12620,N_12591);
or U13052 (N_13052,N_12737,N_12824);
nor U13053 (N_13053,N_12864,N_12566);
nor U13054 (N_13054,N_12751,N_12646);
xor U13055 (N_13055,N_12594,N_12910);
and U13056 (N_13056,N_12980,N_12599);
xnor U13057 (N_13057,N_12784,N_12613);
nor U13058 (N_13058,N_12749,N_12836);
or U13059 (N_13059,N_12637,N_12927);
xnor U13060 (N_13060,N_12678,N_12887);
and U13061 (N_13061,N_12551,N_12850);
xor U13062 (N_13062,N_12807,N_12574);
or U13063 (N_13063,N_12894,N_12607);
xnor U13064 (N_13064,N_12917,N_12981);
nor U13065 (N_13065,N_12796,N_12762);
and U13066 (N_13066,N_12899,N_12605);
nor U13067 (N_13067,N_12986,N_12559);
nor U13068 (N_13068,N_12783,N_12567);
nand U13069 (N_13069,N_12520,N_12861);
and U13070 (N_13070,N_12948,N_12990);
and U13071 (N_13071,N_12742,N_12772);
or U13072 (N_13072,N_12808,N_12549);
or U13073 (N_13073,N_12518,N_12862);
nor U13074 (N_13074,N_12609,N_12795);
nor U13075 (N_13075,N_12564,N_12516);
or U13076 (N_13076,N_12667,N_12619);
and U13077 (N_13077,N_12718,N_12799);
and U13078 (N_13078,N_12503,N_12907);
and U13079 (N_13079,N_12831,N_12712);
nor U13080 (N_13080,N_12550,N_12709);
nor U13081 (N_13081,N_12878,N_12805);
or U13082 (N_13082,N_12792,N_12519);
and U13083 (N_13083,N_12555,N_12588);
and U13084 (N_13084,N_12859,N_12909);
nor U13085 (N_13085,N_12970,N_12675);
and U13086 (N_13086,N_12790,N_12533);
or U13087 (N_13087,N_12911,N_12791);
or U13088 (N_13088,N_12548,N_12806);
or U13089 (N_13089,N_12953,N_12651);
xor U13090 (N_13090,N_12534,N_12502);
nor U13091 (N_13091,N_12640,N_12973);
nor U13092 (N_13092,N_12700,N_12971);
xor U13093 (N_13093,N_12511,N_12882);
nand U13094 (N_13094,N_12979,N_12597);
xor U13095 (N_13095,N_12809,N_12721);
or U13096 (N_13096,N_12913,N_12957);
or U13097 (N_13097,N_12668,N_12950);
nand U13098 (N_13098,N_12881,N_12600);
xnor U13099 (N_13099,N_12754,N_12684);
and U13100 (N_13100,N_12848,N_12816);
or U13101 (N_13101,N_12524,N_12531);
nor U13102 (N_13102,N_12696,N_12645);
nor U13103 (N_13103,N_12835,N_12800);
xor U13104 (N_13104,N_12802,N_12572);
and U13105 (N_13105,N_12673,N_12963);
nor U13106 (N_13106,N_12687,N_12811);
xnor U13107 (N_13107,N_12941,N_12804);
nand U13108 (N_13108,N_12552,N_12527);
or U13109 (N_13109,N_12964,N_12629);
xnor U13110 (N_13110,N_12560,N_12728);
nor U13111 (N_13111,N_12855,N_12625);
nor U13112 (N_13112,N_12918,N_12822);
and U13113 (N_13113,N_12716,N_12501);
or U13114 (N_13114,N_12690,N_12720);
or U13115 (N_13115,N_12537,N_12779);
and U13116 (N_13116,N_12930,N_12873);
xor U13117 (N_13117,N_12830,N_12868);
nand U13118 (N_13118,N_12956,N_12603);
nor U13119 (N_13119,N_12538,N_12639);
or U13120 (N_13120,N_12876,N_12884);
nand U13121 (N_13121,N_12698,N_12775);
nand U13122 (N_13122,N_12929,N_12641);
nor U13123 (N_13123,N_12529,N_12729);
xor U13124 (N_13124,N_12612,N_12648);
and U13125 (N_13125,N_12589,N_12590);
and U13126 (N_13126,N_12727,N_12820);
xnor U13127 (N_13127,N_12631,N_12770);
nand U13128 (N_13128,N_12949,N_12837);
or U13129 (N_13129,N_12715,N_12573);
or U13130 (N_13130,N_12507,N_12984);
xor U13131 (N_13131,N_12959,N_12920);
xor U13132 (N_13132,N_12767,N_12650);
nand U13133 (N_13133,N_12706,N_12602);
xnor U13134 (N_13134,N_12701,N_12505);
xor U13135 (N_13135,N_12854,N_12828);
nand U13136 (N_13136,N_12935,N_12542);
nand U13137 (N_13137,N_12522,N_12926);
or U13138 (N_13138,N_12704,N_12626);
or U13139 (N_13139,N_12671,N_12821);
nor U13140 (N_13140,N_12823,N_12875);
nor U13141 (N_13141,N_12595,N_12571);
and U13142 (N_13142,N_12872,N_12928);
or U13143 (N_13143,N_12825,N_12744);
or U13144 (N_13144,N_12506,N_12988);
and U13145 (N_13145,N_12952,N_12829);
and U13146 (N_13146,N_12686,N_12826);
nor U13147 (N_13147,N_12632,N_12663);
and U13148 (N_13148,N_12798,N_12750);
and U13149 (N_13149,N_12969,N_12618);
or U13150 (N_13150,N_12691,N_12793);
or U13151 (N_13151,N_12892,N_12561);
xor U13152 (N_13152,N_12944,N_12579);
xor U13153 (N_13153,N_12978,N_12908);
nor U13154 (N_13154,N_12766,N_12939);
xnor U13155 (N_13155,N_12581,N_12905);
or U13156 (N_13156,N_12997,N_12545);
or U13157 (N_13157,N_12654,N_12960);
xor U13158 (N_13158,N_12577,N_12797);
nor U13159 (N_13159,N_12692,N_12955);
nor U13160 (N_13160,N_12846,N_12919);
nor U13161 (N_13161,N_12598,N_12841);
nor U13162 (N_13162,N_12583,N_12611);
nand U13163 (N_13163,N_12513,N_12745);
and U13164 (N_13164,N_12815,N_12994);
xnor U13165 (N_13165,N_12521,N_12748);
nand U13166 (N_13166,N_12719,N_12936);
or U13167 (N_13167,N_12896,N_12665);
or U13168 (N_13168,N_12938,N_12880);
nand U13169 (N_13169,N_12723,N_12867);
and U13170 (N_13170,N_12761,N_12832);
and U13171 (N_13171,N_12681,N_12711);
xor U13172 (N_13172,N_12888,N_12622);
and U13173 (N_13173,N_12553,N_12914);
nor U13174 (N_13174,N_12724,N_12525);
nand U13175 (N_13175,N_12635,N_12586);
xnor U13176 (N_13176,N_12987,N_12554);
or U13177 (N_13177,N_12556,N_12530);
nor U13178 (N_13178,N_12563,N_12623);
or U13179 (N_13179,N_12568,N_12819);
or U13180 (N_13180,N_12617,N_12906);
or U13181 (N_13181,N_12814,N_12865);
nor U13182 (N_13182,N_12900,N_12827);
xnor U13183 (N_13183,N_12656,N_12773);
nand U13184 (N_13184,N_12659,N_12593);
nor U13185 (N_13185,N_12889,N_12874);
xor U13186 (N_13186,N_12843,N_12983);
and U13187 (N_13187,N_12839,N_12932);
and U13188 (N_13188,N_12669,N_12858);
or U13189 (N_13189,N_12810,N_12596);
nand U13190 (N_13190,N_12782,N_12652);
and U13191 (N_13191,N_12544,N_12679);
nand U13192 (N_13192,N_12897,N_12780);
nor U13193 (N_13193,N_12512,N_12705);
or U13194 (N_13194,N_12543,N_12777);
xor U13195 (N_13195,N_12756,N_12863);
and U13196 (N_13196,N_12755,N_12666);
nor U13197 (N_13197,N_12958,N_12643);
nand U13198 (N_13198,N_12870,N_12610);
nand U13199 (N_13199,N_12912,N_12731);
and U13200 (N_13200,N_12947,N_12515);
nand U13201 (N_13201,N_12707,N_12940);
nor U13202 (N_13202,N_12871,N_12951);
and U13203 (N_13203,N_12840,N_12689);
nor U13204 (N_13204,N_12697,N_12924);
or U13205 (N_13205,N_12965,N_12974);
xnor U13206 (N_13206,N_12695,N_12833);
xor U13207 (N_13207,N_12627,N_12789);
or U13208 (N_13208,N_12717,N_12781);
nor U13209 (N_13209,N_12636,N_12662);
nor U13210 (N_13210,N_12509,N_12676);
and U13211 (N_13211,N_12528,N_12851);
and U13212 (N_13212,N_12860,N_12672);
nor U13213 (N_13213,N_12541,N_12921);
and U13214 (N_13214,N_12923,N_12743);
or U13215 (N_13215,N_12532,N_12683);
and U13216 (N_13216,N_12834,N_12647);
and U13217 (N_13217,N_12813,N_12937);
nor U13218 (N_13218,N_12585,N_12508);
nand U13219 (N_13219,N_12634,N_12866);
nand U13220 (N_13220,N_12753,N_12702);
nand U13221 (N_13221,N_12838,N_12674);
xor U13222 (N_13222,N_12699,N_12818);
nor U13223 (N_13223,N_12977,N_12547);
xor U13224 (N_13224,N_12759,N_12569);
nand U13225 (N_13225,N_12576,N_12630);
nor U13226 (N_13226,N_12982,N_12736);
nor U13227 (N_13227,N_12747,N_12788);
nor U13228 (N_13228,N_12562,N_12801);
nand U13229 (N_13229,N_12763,N_12680);
or U13230 (N_13230,N_12587,N_12885);
and U13231 (N_13231,N_12842,N_12904);
and U13232 (N_13232,N_12708,N_12733);
and U13233 (N_13233,N_12943,N_12901);
nor U13234 (N_13234,N_12857,N_12739);
nand U13235 (N_13235,N_12713,N_12694);
nor U13236 (N_13236,N_12658,N_12615);
nor U13237 (N_13237,N_12902,N_12769);
nand U13238 (N_13238,N_12847,N_12886);
and U13239 (N_13239,N_12608,N_12787);
nand U13240 (N_13240,N_12510,N_12664);
xor U13241 (N_13241,N_12954,N_12606);
nand U13242 (N_13242,N_12972,N_12584);
or U13243 (N_13243,N_12570,N_12535);
or U13244 (N_13244,N_12578,N_12898);
xnor U13245 (N_13245,N_12517,N_12968);
xor U13246 (N_13246,N_12962,N_12849);
and U13247 (N_13247,N_12670,N_12989);
or U13248 (N_13248,N_12735,N_12546);
nand U13249 (N_13249,N_12614,N_12624);
nor U13250 (N_13250,N_12862,N_12526);
nand U13251 (N_13251,N_12991,N_12759);
or U13252 (N_13252,N_12676,N_12745);
nor U13253 (N_13253,N_12624,N_12911);
or U13254 (N_13254,N_12683,N_12691);
and U13255 (N_13255,N_12940,N_12946);
nand U13256 (N_13256,N_12620,N_12864);
nand U13257 (N_13257,N_12727,N_12849);
or U13258 (N_13258,N_12643,N_12501);
xnor U13259 (N_13259,N_12990,N_12764);
or U13260 (N_13260,N_12688,N_12864);
nand U13261 (N_13261,N_12914,N_12933);
and U13262 (N_13262,N_12779,N_12970);
xnor U13263 (N_13263,N_12680,N_12517);
nor U13264 (N_13264,N_12807,N_12601);
nor U13265 (N_13265,N_12795,N_12837);
xor U13266 (N_13266,N_12804,N_12642);
nand U13267 (N_13267,N_12802,N_12613);
or U13268 (N_13268,N_12908,N_12964);
xnor U13269 (N_13269,N_12897,N_12888);
nor U13270 (N_13270,N_12807,N_12729);
nand U13271 (N_13271,N_12652,N_12817);
or U13272 (N_13272,N_12967,N_12601);
or U13273 (N_13273,N_12770,N_12636);
nand U13274 (N_13274,N_12530,N_12507);
or U13275 (N_13275,N_12655,N_12580);
or U13276 (N_13276,N_12685,N_12932);
and U13277 (N_13277,N_12517,N_12730);
xor U13278 (N_13278,N_12848,N_12901);
nor U13279 (N_13279,N_12949,N_12640);
or U13280 (N_13280,N_12805,N_12840);
nand U13281 (N_13281,N_12686,N_12870);
nand U13282 (N_13282,N_12646,N_12993);
and U13283 (N_13283,N_12969,N_12578);
or U13284 (N_13284,N_12598,N_12766);
nor U13285 (N_13285,N_12648,N_12537);
and U13286 (N_13286,N_12923,N_12998);
or U13287 (N_13287,N_12654,N_12578);
and U13288 (N_13288,N_12957,N_12880);
nor U13289 (N_13289,N_12860,N_12906);
nor U13290 (N_13290,N_12881,N_12724);
or U13291 (N_13291,N_12685,N_12693);
xor U13292 (N_13292,N_12891,N_12854);
xnor U13293 (N_13293,N_12925,N_12945);
nor U13294 (N_13294,N_12953,N_12975);
and U13295 (N_13295,N_12673,N_12807);
nor U13296 (N_13296,N_12589,N_12917);
nand U13297 (N_13297,N_12560,N_12879);
xnor U13298 (N_13298,N_12830,N_12716);
and U13299 (N_13299,N_12923,N_12905);
and U13300 (N_13300,N_12611,N_12709);
nor U13301 (N_13301,N_12809,N_12823);
or U13302 (N_13302,N_12833,N_12725);
xnor U13303 (N_13303,N_12697,N_12936);
nor U13304 (N_13304,N_12502,N_12682);
nor U13305 (N_13305,N_12700,N_12992);
or U13306 (N_13306,N_12750,N_12616);
nand U13307 (N_13307,N_12715,N_12918);
xor U13308 (N_13308,N_12970,N_12814);
xnor U13309 (N_13309,N_12768,N_12659);
nor U13310 (N_13310,N_12643,N_12727);
and U13311 (N_13311,N_12914,N_12566);
nor U13312 (N_13312,N_12818,N_12985);
or U13313 (N_13313,N_12895,N_12813);
xnor U13314 (N_13314,N_12724,N_12988);
xor U13315 (N_13315,N_12533,N_12605);
and U13316 (N_13316,N_12537,N_12531);
and U13317 (N_13317,N_12817,N_12916);
or U13318 (N_13318,N_12625,N_12666);
nand U13319 (N_13319,N_12949,N_12875);
nor U13320 (N_13320,N_12801,N_12540);
xnor U13321 (N_13321,N_12612,N_12987);
and U13322 (N_13322,N_12511,N_12955);
nand U13323 (N_13323,N_12917,N_12735);
nand U13324 (N_13324,N_12866,N_12905);
and U13325 (N_13325,N_12862,N_12748);
nand U13326 (N_13326,N_12750,N_12902);
xor U13327 (N_13327,N_12673,N_12728);
nand U13328 (N_13328,N_12612,N_12587);
nand U13329 (N_13329,N_12965,N_12929);
xnor U13330 (N_13330,N_12566,N_12831);
and U13331 (N_13331,N_12609,N_12831);
or U13332 (N_13332,N_12681,N_12818);
or U13333 (N_13333,N_12894,N_12644);
and U13334 (N_13334,N_12578,N_12680);
nor U13335 (N_13335,N_12664,N_12566);
nor U13336 (N_13336,N_12583,N_12629);
and U13337 (N_13337,N_12731,N_12657);
nand U13338 (N_13338,N_12889,N_12679);
nand U13339 (N_13339,N_12799,N_12526);
xor U13340 (N_13340,N_12962,N_12793);
or U13341 (N_13341,N_12870,N_12852);
nor U13342 (N_13342,N_12962,N_12511);
or U13343 (N_13343,N_12550,N_12971);
or U13344 (N_13344,N_12693,N_12559);
nor U13345 (N_13345,N_12877,N_12912);
nand U13346 (N_13346,N_12878,N_12777);
or U13347 (N_13347,N_12520,N_12637);
nand U13348 (N_13348,N_12935,N_12650);
and U13349 (N_13349,N_12992,N_12825);
and U13350 (N_13350,N_12573,N_12544);
nand U13351 (N_13351,N_12626,N_12779);
nor U13352 (N_13352,N_12764,N_12523);
and U13353 (N_13353,N_12762,N_12874);
xor U13354 (N_13354,N_12921,N_12688);
nand U13355 (N_13355,N_12702,N_12751);
or U13356 (N_13356,N_12957,N_12681);
or U13357 (N_13357,N_12857,N_12874);
and U13358 (N_13358,N_12962,N_12563);
nor U13359 (N_13359,N_12579,N_12857);
xor U13360 (N_13360,N_12798,N_12602);
or U13361 (N_13361,N_12732,N_12520);
xnor U13362 (N_13362,N_12697,N_12738);
nand U13363 (N_13363,N_12673,N_12967);
nand U13364 (N_13364,N_12817,N_12574);
nand U13365 (N_13365,N_12529,N_12763);
nor U13366 (N_13366,N_12990,N_12627);
and U13367 (N_13367,N_12843,N_12900);
and U13368 (N_13368,N_12501,N_12852);
xnor U13369 (N_13369,N_12668,N_12522);
nand U13370 (N_13370,N_12660,N_12600);
xnor U13371 (N_13371,N_12817,N_12963);
and U13372 (N_13372,N_12500,N_12702);
or U13373 (N_13373,N_12988,N_12711);
nor U13374 (N_13374,N_12668,N_12880);
and U13375 (N_13375,N_12803,N_12919);
and U13376 (N_13376,N_12619,N_12722);
and U13377 (N_13377,N_12687,N_12930);
and U13378 (N_13378,N_12908,N_12817);
and U13379 (N_13379,N_12917,N_12501);
xnor U13380 (N_13380,N_12644,N_12919);
nand U13381 (N_13381,N_12555,N_12584);
xnor U13382 (N_13382,N_12663,N_12502);
nor U13383 (N_13383,N_12792,N_12566);
xnor U13384 (N_13384,N_12794,N_12567);
xor U13385 (N_13385,N_12976,N_12797);
or U13386 (N_13386,N_12851,N_12644);
and U13387 (N_13387,N_12536,N_12781);
or U13388 (N_13388,N_12513,N_12503);
or U13389 (N_13389,N_12892,N_12843);
and U13390 (N_13390,N_12824,N_12836);
nor U13391 (N_13391,N_12945,N_12901);
nor U13392 (N_13392,N_12652,N_12919);
or U13393 (N_13393,N_12934,N_12721);
nor U13394 (N_13394,N_12660,N_12824);
or U13395 (N_13395,N_12656,N_12726);
and U13396 (N_13396,N_12541,N_12802);
and U13397 (N_13397,N_12939,N_12627);
and U13398 (N_13398,N_12742,N_12751);
and U13399 (N_13399,N_12617,N_12542);
xor U13400 (N_13400,N_12724,N_12667);
nor U13401 (N_13401,N_12919,N_12712);
and U13402 (N_13402,N_12634,N_12532);
nand U13403 (N_13403,N_12928,N_12516);
nor U13404 (N_13404,N_12600,N_12999);
xor U13405 (N_13405,N_12947,N_12501);
and U13406 (N_13406,N_12678,N_12749);
or U13407 (N_13407,N_12675,N_12840);
xor U13408 (N_13408,N_12863,N_12938);
nor U13409 (N_13409,N_12642,N_12956);
nand U13410 (N_13410,N_12789,N_12610);
nand U13411 (N_13411,N_12637,N_12843);
xnor U13412 (N_13412,N_12930,N_12876);
xnor U13413 (N_13413,N_12900,N_12527);
nor U13414 (N_13414,N_12945,N_12805);
or U13415 (N_13415,N_12824,N_12711);
xor U13416 (N_13416,N_12810,N_12889);
xor U13417 (N_13417,N_12649,N_12570);
nor U13418 (N_13418,N_12893,N_12936);
nand U13419 (N_13419,N_12587,N_12705);
nand U13420 (N_13420,N_12820,N_12909);
nand U13421 (N_13421,N_12677,N_12726);
or U13422 (N_13422,N_12747,N_12706);
xor U13423 (N_13423,N_12774,N_12853);
nand U13424 (N_13424,N_12792,N_12730);
or U13425 (N_13425,N_12546,N_12538);
xor U13426 (N_13426,N_12541,N_12841);
nand U13427 (N_13427,N_12822,N_12613);
xnor U13428 (N_13428,N_12569,N_12915);
nand U13429 (N_13429,N_12885,N_12591);
xnor U13430 (N_13430,N_12819,N_12942);
nand U13431 (N_13431,N_12919,N_12975);
nand U13432 (N_13432,N_12889,N_12947);
and U13433 (N_13433,N_12682,N_12892);
and U13434 (N_13434,N_12892,N_12722);
and U13435 (N_13435,N_12521,N_12859);
nand U13436 (N_13436,N_12794,N_12895);
nand U13437 (N_13437,N_12629,N_12893);
nand U13438 (N_13438,N_12613,N_12992);
and U13439 (N_13439,N_12883,N_12709);
nor U13440 (N_13440,N_12779,N_12951);
nand U13441 (N_13441,N_12798,N_12800);
nand U13442 (N_13442,N_12524,N_12610);
nand U13443 (N_13443,N_12762,N_12991);
and U13444 (N_13444,N_12916,N_12658);
xor U13445 (N_13445,N_12503,N_12643);
and U13446 (N_13446,N_12817,N_12803);
and U13447 (N_13447,N_12611,N_12517);
nor U13448 (N_13448,N_12773,N_12899);
xor U13449 (N_13449,N_12930,N_12797);
nor U13450 (N_13450,N_12639,N_12742);
nor U13451 (N_13451,N_12813,N_12943);
and U13452 (N_13452,N_12818,N_12634);
or U13453 (N_13453,N_12773,N_12837);
and U13454 (N_13454,N_12625,N_12713);
nand U13455 (N_13455,N_12593,N_12797);
nor U13456 (N_13456,N_12769,N_12781);
or U13457 (N_13457,N_12974,N_12766);
or U13458 (N_13458,N_12781,N_12777);
or U13459 (N_13459,N_12953,N_12520);
and U13460 (N_13460,N_12694,N_12852);
or U13461 (N_13461,N_12761,N_12577);
xnor U13462 (N_13462,N_12714,N_12541);
and U13463 (N_13463,N_12809,N_12840);
xor U13464 (N_13464,N_12779,N_12591);
or U13465 (N_13465,N_12589,N_12765);
nor U13466 (N_13466,N_12863,N_12796);
nand U13467 (N_13467,N_12937,N_12870);
nand U13468 (N_13468,N_12679,N_12752);
or U13469 (N_13469,N_12823,N_12933);
nand U13470 (N_13470,N_12686,N_12748);
or U13471 (N_13471,N_12864,N_12856);
nand U13472 (N_13472,N_12539,N_12700);
or U13473 (N_13473,N_12703,N_12674);
and U13474 (N_13474,N_12745,N_12590);
nand U13475 (N_13475,N_12553,N_12772);
xnor U13476 (N_13476,N_12695,N_12933);
nand U13477 (N_13477,N_12799,N_12689);
nand U13478 (N_13478,N_12884,N_12837);
xor U13479 (N_13479,N_12820,N_12809);
and U13480 (N_13480,N_12615,N_12807);
and U13481 (N_13481,N_12730,N_12968);
and U13482 (N_13482,N_12631,N_12811);
nand U13483 (N_13483,N_12722,N_12584);
xor U13484 (N_13484,N_12803,N_12530);
xnor U13485 (N_13485,N_12970,N_12994);
nor U13486 (N_13486,N_12966,N_12702);
nor U13487 (N_13487,N_12873,N_12987);
and U13488 (N_13488,N_12945,N_12801);
nand U13489 (N_13489,N_12649,N_12554);
nor U13490 (N_13490,N_12640,N_12647);
and U13491 (N_13491,N_12992,N_12665);
xnor U13492 (N_13492,N_12616,N_12738);
and U13493 (N_13493,N_12707,N_12614);
and U13494 (N_13494,N_12915,N_12760);
nand U13495 (N_13495,N_12517,N_12787);
nand U13496 (N_13496,N_12930,N_12576);
or U13497 (N_13497,N_12764,N_12849);
xnor U13498 (N_13498,N_12952,N_12998);
and U13499 (N_13499,N_12783,N_12726);
nor U13500 (N_13500,N_13072,N_13459);
and U13501 (N_13501,N_13385,N_13313);
and U13502 (N_13502,N_13286,N_13057);
nand U13503 (N_13503,N_13298,N_13239);
nor U13504 (N_13504,N_13254,N_13299);
xnor U13505 (N_13505,N_13377,N_13292);
xor U13506 (N_13506,N_13097,N_13091);
nor U13507 (N_13507,N_13346,N_13386);
xor U13508 (N_13508,N_13441,N_13053);
and U13509 (N_13509,N_13045,N_13479);
xnor U13510 (N_13510,N_13174,N_13063);
nand U13511 (N_13511,N_13396,N_13328);
or U13512 (N_13512,N_13167,N_13276);
xor U13513 (N_13513,N_13090,N_13223);
xnor U13514 (N_13514,N_13327,N_13410);
nor U13515 (N_13515,N_13234,N_13211);
and U13516 (N_13516,N_13071,N_13061);
xnor U13517 (N_13517,N_13191,N_13403);
or U13518 (N_13518,N_13028,N_13249);
nand U13519 (N_13519,N_13026,N_13336);
nor U13520 (N_13520,N_13092,N_13088);
nand U13521 (N_13521,N_13078,N_13205);
or U13522 (N_13522,N_13388,N_13378);
or U13523 (N_13523,N_13348,N_13280);
or U13524 (N_13524,N_13259,N_13204);
xor U13525 (N_13525,N_13374,N_13151);
xnor U13526 (N_13526,N_13193,N_13447);
nand U13527 (N_13527,N_13435,N_13210);
nand U13528 (N_13528,N_13450,N_13414);
or U13529 (N_13529,N_13290,N_13323);
and U13530 (N_13530,N_13436,N_13007);
and U13531 (N_13531,N_13251,N_13423);
xnor U13532 (N_13532,N_13464,N_13296);
xnor U13533 (N_13533,N_13149,N_13489);
and U13534 (N_13534,N_13017,N_13331);
nand U13535 (N_13535,N_13206,N_13418);
xnor U13536 (N_13536,N_13340,N_13256);
nand U13537 (N_13537,N_13409,N_13006);
or U13538 (N_13538,N_13356,N_13482);
or U13539 (N_13539,N_13132,N_13443);
and U13540 (N_13540,N_13085,N_13067);
xnor U13541 (N_13541,N_13069,N_13173);
or U13542 (N_13542,N_13080,N_13042);
or U13543 (N_13543,N_13220,N_13333);
and U13544 (N_13544,N_13082,N_13359);
nor U13545 (N_13545,N_13355,N_13363);
nor U13546 (N_13546,N_13165,N_13121);
nand U13547 (N_13547,N_13314,N_13177);
nand U13548 (N_13548,N_13473,N_13122);
xnor U13549 (N_13549,N_13209,N_13446);
and U13550 (N_13550,N_13487,N_13406);
or U13551 (N_13551,N_13233,N_13214);
nor U13552 (N_13552,N_13189,N_13154);
nand U13553 (N_13553,N_13319,N_13253);
or U13554 (N_13554,N_13390,N_13188);
nor U13555 (N_13555,N_13245,N_13094);
or U13556 (N_13556,N_13486,N_13027);
and U13557 (N_13557,N_13244,N_13427);
nor U13558 (N_13558,N_13279,N_13415);
and U13559 (N_13559,N_13420,N_13407);
and U13560 (N_13560,N_13162,N_13039);
or U13561 (N_13561,N_13268,N_13303);
or U13562 (N_13562,N_13275,N_13324);
or U13563 (N_13563,N_13004,N_13339);
nor U13564 (N_13564,N_13195,N_13203);
nand U13565 (N_13565,N_13170,N_13497);
and U13566 (N_13566,N_13466,N_13389);
or U13567 (N_13567,N_13412,N_13438);
xor U13568 (N_13568,N_13467,N_13140);
nor U13569 (N_13569,N_13023,N_13460);
xnor U13570 (N_13570,N_13117,N_13202);
nor U13571 (N_13571,N_13086,N_13477);
xor U13572 (N_13572,N_13016,N_13156);
nor U13573 (N_13573,N_13228,N_13105);
and U13574 (N_13574,N_13498,N_13136);
xnor U13575 (N_13575,N_13011,N_13181);
nor U13576 (N_13576,N_13432,N_13133);
nor U13577 (N_13577,N_13469,N_13293);
xnor U13578 (N_13578,N_13106,N_13369);
nor U13579 (N_13579,N_13083,N_13169);
or U13580 (N_13580,N_13131,N_13213);
or U13581 (N_13581,N_13076,N_13231);
and U13582 (N_13582,N_13095,N_13046);
or U13583 (N_13583,N_13014,N_13087);
xor U13584 (N_13584,N_13033,N_13431);
nand U13585 (N_13585,N_13036,N_13257);
and U13586 (N_13586,N_13393,N_13287);
nand U13587 (N_13587,N_13190,N_13212);
nand U13588 (N_13588,N_13449,N_13305);
and U13589 (N_13589,N_13222,N_13332);
nand U13590 (N_13590,N_13000,N_13391);
or U13591 (N_13591,N_13098,N_13029);
xor U13592 (N_13592,N_13421,N_13186);
nor U13593 (N_13593,N_13301,N_13208);
or U13594 (N_13594,N_13445,N_13242);
nand U13595 (N_13595,N_13454,N_13059);
xor U13596 (N_13596,N_13005,N_13178);
nor U13597 (N_13597,N_13325,N_13411);
nor U13598 (N_13598,N_13395,N_13089);
nand U13599 (N_13599,N_13401,N_13093);
nor U13600 (N_13600,N_13232,N_13003);
nor U13601 (N_13601,N_13426,N_13134);
xor U13602 (N_13602,N_13144,N_13399);
nor U13603 (N_13603,N_13175,N_13269);
or U13604 (N_13604,N_13020,N_13491);
nor U13605 (N_13605,N_13316,N_13031);
or U13606 (N_13606,N_13044,N_13141);
and U13607 (N_13607,N_13338,N_13265);
or U13608 (N_13608,N_13096,N_13066);
nand U13609 (N_13609,N_13272,N_13052);
xor U13610 (N_13610,N_13152,N_13428);
nor U13611 (N_13611,N_13456,N_13297);
or U13612 (N_13612,N_13019,N_13326);
nor U13613 (N_13613,N_13452,N_13488);
or U13614 (N_13614,N_13372,N_13074);
nand U13615 (N_13615,N_13103,N_13010);
and U13616 (N_13616,N_13110,N_13495);
nand U13617 (N_13617,N_13476,N_13168);
xor U13618 (N_13618,N_13264,N_13439);
nand U13619 (N_13619,N_13371,N_13358);
and U13620 (N_13620,N_13442,N_13444);
nor U13621 (N_13621,N_13382,N_13049);
nor U13622 (N_13622,N_13183,N_13365);
xor U13623 (N_13623,N_13367,N_13274);
nand U13624 (N_13624,N_13062,N_13047);
or U13625 (N_13625,N_13038,N_13184);
and U13626 (N_13626,N_13229,N_13224);
xor U13627 (N_13627,N_13381,N_13109);
or U13628 (N_13628,N_13343,N_13468);
nand U13629 (N_13629,N_13041,N_13375);
or U13630 (N_13630,N_13102,N_13058);
nand U13631 (N_13631,N_13425,N_13334);
and U13632 (N_13632,N_13392,N_13304);
nor U13633 (N_13633,N_13187,N_13250);
xnor U13634 (N_13634,N_13267,N_13157);
or U13635 (N_13635,N_13252,N_13079);
or U13636 (N_13636,N_13379,N_13101);
and U13637 (N_13637,N_13260,N_13176);
or U13638 (N_13638,N_13135,N_13200);
nand U13639 (N_13639,N_13361,N_13337);
and U13640 (N_13640,N_13362,N_13164);
xnor U13641 (N_13641,N_13376,N_13322);
or U13642 (N_13642,N_13373,N_13430);
xnor U13643 (N_13643,N_13398,N_13283);
and U13644 (N_13644,N_13277,N_13463);
nor U13645 (N_13645,N_13417,N_13002);
nand U13646 (N_13646,N_13113,N_13320);
nor U13647 (N_13647,N_13353,N_13125);
or U13648 (N_13648,N_13349,N_13318);
or U13649 (N_13649,N_13118,N_13284);
xnor U13650 (N_13650,N_13060,N_13345);
or U13651 (N_13651,N_13147,N_13111);
nand U13652 (N_13652,N_13015,N_13306);
and U13653 (N_13653,N_13461,N_13050);
xnor U13654 (N_13654,N_13448,N_13009);
nand U13655 (N_13655,N_13230,N_13143);
nor U13656 (N_13656,N_13470,N_13317);
nor U13657 (N_13657,N_13351,N_13383);
nand U13658 (N_13658,N_13455,N_13243);
xor U13659 (N_13659,N_13309,N_13051);
and U13660 (N_13660,N_13483,N_13226);
and U13661 (N_13661,N_13494,N_13278);
nand U13662 (N_13662,N_13240,N_13241);
nor U13663 (N_13663,N_13018,N_13030);
nor U13664 (N_13664,N_13453,N_13295);
and U13665 (N_13665,N_13273,N_13022);
nand U13666 (N_13666,N_13070,N_13370);
and U13667 (N_13667,N_13148,N_13413);
and U13668 (N_13668,N_13237,N_13380);
nand U13669 (N_13669,N_13166,N_13159);
xnor U13670 (N_13670,N_13225,N_13262);
nand U13671 (N_13671,N_13481,N_13099);
or U13672 (N_13672,N_13311,N_13137);
nand U13673 (N_13673,N_13075,N_13416);
xor U13674 (N_13674,N_13227,N_13160);
and U13675 (N_13675,N_13307,N_13219);
or U13676 (N_13676,N_13451,N_13116);
nor U13677 (N_13677,N_13302,N_13255);
and U13678 (N_13678,N_13215,N_13024);
or U13679 (N_13679,N_13107,N_13040);
xor U13680 (N_13680,N_13402,N_13138);
and U13681 (N_13681,N_13179,N_13480);
nand U13682 (N_13682,N_13185,N_13248);
nand U13683 (N_13683,N_13238,N_13246);
xor U13684 (N_13684,N_13115,N_13043);
or U13685 (N_13685,N_13150,N_13073);
nand U13686 (N_13686,N_13218,N_13270);
or U13687 (N_13687,N_13457,N_13490);
and U13688 (N_13688,N_13342,N_13261);
and U13689 (N_13689,N_13180,N_13437);
nor U13690 (N_13690,N_13081,N_13155);
and U13691 (N_13691,N_13124,N_13397);
xnor U13692 (N_13692,N_13104,N_13424);
or U13693 (N_13693,N_13440,N_13266);
and U13694 (N_13694,N_13294,N_13034);
and U13695 (N_13695,N_13408,N_13108);
nor U13696 (N_13696,N_13285,N_13054);
xnor U13697 (N_13697,N_13321,N_13496);
nand U13698 (N_13698,N_13128,N_13474);
nand U13699 (N_13699,N_13130,N_13289);
or U13700 (N_13700,N_13308,N_13350);
and U13701 (N_13701,N_13433,N_13127);
xnor U13702 (N_13702,N_13217,N_13329);
and U13703 (N_13703,N_13025,N_13126);
nor U13704 (N_13704,N_13037,N_13100);
xnor U13705 (N_13705,N_13112,N_13485);
nor U13706 (N_13706,N_13064,N_13300);
or U13707 (N_13707,N_13387,N_13499);
or U13708 (N_13708,N_13129,N_13145);
and U13709 (N_13709,N_13282,N_13405);
nor U13710 (N_13710,N_13196,N_13236);
or U13711 (N_13711,N_13035,N_13344);
xor U13712 (N_13712,N_13493,N_13008);
and U13713 (N_13713,N_13422,N_13458);
nor U13714 (N_13714,N_13310,N_13171);
nor U13715 (N_13715,N_13366,N_13434);
and U13716 (N_13716,N_13368,N_13384);
or U13717 (N_13717,N_13032,N_13492);
and U13718 (N_13718,N_13077,N_13247);
nand U13719 (N_13719,N_13013,N_13199);
or U13720 (N_13720,N_13001,N_13352);
xor U13721 (N_13721,N_13341,N_13400);
xor U13722 (N_13722,N_13330,N_13281);
and U13723 (N_13723,N_13161,N_13429);
and U13724 (N_13724,N_13065,N_13146);
or U13725 (N_13725,N_13315,N_13347);
nor U13726 (N_13726,N_13216,N_13258);
nand U13727 (N_13727,N_13207,N_13153);
nor U13728 (N_13728,N_13194,N_13360);
nor U13729 (N_13729,N_13084,N_13055);
and U13730 (N_13730,N_13182,N_13475);
nor U13731 (N_13731,N_13068,N_13119);
nor U13732 (N_13732,N_13021,N_13192);
or U13733 (N_13733,N_13139,N_13056);
nand U13734 (N_13734,N_13288,N_13335);
or U13735 (N_13735,N_13142,N_13394);
xnor U13736 (N_13736,N_13465,N_13357);
nand U13737 (N_13737,N_13163,N_13235);
and U13738 (N_13738,N_13114,N_13364);
xnor U13739 (N_13739,N_13048,N_13123);
nor U13740 (N_13740,N_13478,N_13484);
and U13741 (N_13741,N_13221,N_13419);
or U13742 (N_13742,N_13471,N_13271);
and U13743 (N_13743,N_13404,N_13472);
xor U13744 (N_13744,N_13263,N_13198);
and U13745 (N_13745,N_13120,N_13312);
and U13746 (N_13746,N_13201,N_13197);
xor U13747 (N_13747,N_13012,N_13291);
nand U13748 (N_13748,N_13158,N_13462);
xnor U13749 (N_13749,N_13172,N_13354);
and U13750 (N_13750,N_13499,N_13016);
and U13751 (N_13751,N_13347,N_13372);
and U13752 (N_13752,N_13056,N_13429);
nor U13753 (N_13753,N_13328,N_13323);
xnor U13754 (N_13754,N_13022,N_13272);
or U13755 (N_13755,N_13494,N_13208);
and U13756 (N_13756,N_13183,N_13171);
nor U13757 (N_13757,N_13194,N_13228);
and U13758 (N_13758,N_13433,N_13182);
xnor U13759 (N_13759,N_13101,N_13290);
nand U13760 (N_13760,N_13112,N_13384);
nand U13761 (N_13761,N_13485,N_13309);
nand U13762 (N_13762,N_13065,N_13492);
nand U13763 (N_13763,N_13094,N_13435);
nand U13764 (N_13764,N_13398,N_13213);
and U13765 (N_13765,N_13046,N_13127);
and U13766 (N_13766,N_13399,N_13035);
or U13767 (N_13767,N_13466,N_13141);
nor U13768 (N_13768,N_13351,N_13453);
and U13769 (N_13769,N_13442,N_13368);
and U13770 (N_13770,N_13196,N_13148);
or U13771 (N_13771,N_13138,N_13236);
nand U13772 (N_13772,N_13358,N_13136);
nand U13773 (N_13773,N_13444,N_13043);
nor U13774 (N_13774,N_13369,N_13326);
xnor U13775 (N_13775,N_13258,N_13366);
or U13776 (N_13776,N_13370,N_13035);
or U13777 (N_13777,N_13225,N_13304);
xnor U13778 (N_13778,N_13108,N_13377);
nand U13779 (N_13779,N_13451,N_13411);
or U13780 (N_13780,N_13031,N_13340);
nor U13781 (N_13781,N_13313,N_13475);
and U13782 (N_13782,N_13416,N_13387);
or U13783 (N_13783,N_13276,N_13112);
nand U13784 (N_13784,N_13437,N_13031);
or U13785 (N_13785,N_13048,N_13169);
xnor U13786 (N_13786,N_13462,N_13427);
xor U13787 (N_13787,N_13223,N_13317);
and U13788 (N_13788,N_13404,N_13120);
and U13789 (N_13789,N_13221,N_13258);
nor U13790 (N_13790,N_13171,N_13398);
nor U13791 (N_13791,N_13392,N_13155);
nor U13792 (N_13792,N_13078,N_13464);
or U13793 (N_13793,N_13408,N_13206);
xnor U13794 (N_13794,N_13160,N_13193);
or U13795 (N_13795,N_13479,N_13110);
xnor U13796 (N_13796,N_13145,N_13044);
xnor U13797 (N_13797,N_13071,N_13257);
nand U13798 (N_13798,N_13183,N_13332);
or U13799 (N_13799,N_13321,N_13333);
xnor U13800 (N_13800,N_13115,N_13081);
or U13801 (N_13801,N_13123,N_13058);
and U13802 (N_13802,N_13086,N_13079);
xnor U13803 (N_13803,N_13088,N_13086);
nand U13804 (N_13804,N_13290,N_13319);
nand U13805 (N_13805,N_13353,N_13406);
nor U13806 (N_13806,N_13000,N_13067);
and U13807 (N_13807,N_13234,N_13243);
nand U13808 (N_13808,N_13440,N_13258);
and U13809 (N_13809,N_13229,N_13027);
nand U13810 (N_13810,N_13275,N_13360);
nand U13811 (N_13811,N_13355,N_13050);
or U13812 (N_13812,N_13370,N_13423);
and U13813 (N_13813,N_13316,N_13314);
nor U13814 (N_13814,N_13130,N_13022);
xor U13815 (N_13815,N_13240,N_13379);
and U13816 (N_13816,N_13192,N_13494);
xnor U13817 (N_13817,N_13358,N_13158);
and U13818 (N_13818,N_13330,N_13323);
nand U13819 (N_13819,N_13169,N_13020);
or U13820 (N_13820,N_13209,N_13292);
nand U13821 (N_13821,N_13202,N_13046);
and U13822 (N_13822,N_13025,N_13172);
xnor U13823 (N_13823,N_13154,N_13131);
and U13824 (N_13824,N_13306,N_13339);
nor U13825 (N_13825,N_13193,N_13387);
nand U13826 (N_13826,N_13157,N_13219);
or U13827 (N_13827,N_13346,N_13075);
nand U13828 (N_13828,N_13037,N_13478);
and U13829 (N_13829,N_13161,N_13324);
nor U13830 (N_13830,N_13307,N_13004);
and U13831 (N_13831,N_13444,N_13328);
nand U13832 (N_13832,N_13039,N_13293);
and U13833 (N_13833,N_13359,N_13354);
xnor U13834 (N_13834,N_13048,N_13162);
nor U13835 (N_13835,N_13008,N_13031);
nand U13836 (N_13836,N_13285,N_13432);
or U13837 (N_13837,N_13036,N_13326);
nand U13838 (N_13838,N_13115,N_13116);
or U13839 (N_13839,N_13080,N_13116);
or U13840 (N_13840,N_13262,N_13012);
nand U13841 (N_13841,N_13039,N_13210);
nor U13842 (N_13842,N_13079,N_13387);
xor U13843 (N_13843,N_13201,N_13314);
nand U13844 (N_13844,N_13476,N_13028);
nand U13845 (N_13845,N_13275,N_13294);
or U13846 (N_13846,N_13339,N_13065);
nand U13847 (N_13847,N_13240,N_13194);
xor U13848 (N_13848,N_13359,N_13272);
nand U13849 (N_13849,N_13200,N_13336);
and U13850 (N_13850,N_13488,N_13245);
and U13851 (N_13851,N_13217,N_13005);
xnor U13852 (N_13852,N_13266,N_13490);
xor U13853 (N_13853,N_13476,N_13090);
or U13854 (N_13854,N_13490,N_13329);
nor U13855 (N_13855,N_13289,N_13443);
and U13856 (N_13856,N_13432,N_13127);
or U13857 (N_13857,N_13283,N_13445);
or U13858 (N_13858,N_13321,N_13227);
or U13859 (N_13859,N_13325,N_13422);
nand U13860 (N_13860,N_13130,N_13458);
nor U13861 (N_13861,N_13138,N_13306);
xor U13862 (N_13862,N_13391,N_13063);
xor U13863 (N_13863,N_13419,N_13076);
and U13864 (N_13864,N_13305,N_13003);
or U13865 (N_13865,N_13116,N_13050);
nand U13866 (N_13866,N_13256,N_13288);
nor U13867 (N_13867,N_13450,N_13384);
nor U13868 (N_13868,N_13237,N_13163);
and U13869 (N_13869,N_13283,N_13368);
or U13870 (N_13870,N_13207,N_13136);
xor U13871 (N_13871,N_13151,N_13246);
xnor U13872 (N_13872,N_13471,N_13383);
and U13873 (N_13873,N_13195,N_13423);
and U13874 (N_13874,N_13263,N_13338);
or U13875 (N_13875,N_13157,N_13274);
or U13876 (N_13876,N_13060,N_13055);
or U13877 (N_13877,N_13180,N_13178);
nor U13878 (N_13878,N_13469,N_13216);
xor U13879 (N_13879,N_13275,N_13303);
nor U13880 (N_13880,N_13377,N_13345);
and U13881 (N_13881,N_13177,N_13339);
nor U13882 (N_13882,N_13083,N_13475);
nand U13883 (N_13883,N_13275,N_13083);
nand U13884 (N_13884,N_13252,N_13099);
nand U13885 (N_13885,N_13292,N_13410);
and U13886 (N_13886,N_13425,N_13210);
xor U13887 (N_13887,N_13113,N_13134);
nor U13888 (N_13888,N_13381,N_13017);
nor U13889 (N_13889,N_13484,N_13144);
xor U13890 (N_13890,N_13330,N_13399);
nand U13891 (N_13891,N_13479,N_13143);
and U13892 (N_13892,N_13157,N_13210);
or U13893 (N_13893,N_13040,N_13256);
nand U13894 (N_13894,N_13348,N_13088);
xnor U13895 (N_13895,N_13349,N_13145);
and U13896 (N_13896,N_13384,N_13258);
xnor U13897 (N_13897,N_13359,N_13161);
or U13898 (N_13898,N_13347,N_13002);
xor U13899 (N_13899,N_13131,N_13424);
xor U13900 (N_13900,N_13358,N_13054);
or U13901 (N_13901,N_13081,N_13274);
or U13902 (N_13902,N_13025,N_13100);
xor U13903 (N_13903,N_13477,N_13126);
and U13904 (N_13904,N_13101,N_13413);
or U13905 (N_13905,N_13175,N_13003);
xnor U13906 (N_13906,N_13413,N_13368);
xor U13907 (N_13907,N_13118,N_13163);
nor U13908 (N_13908,N_13495,N_13485);
xnor U13909 (N_13909,N_13390,N_13377);
nor U13910 (N_13910,N_13362,N_13134);
and U13911 (N_13911,N_13112,N_13274);
nand U13912 (N_13912,N_13490,N_13117);
and U13913 (N_13913,N_13072,N_13268);
nor U13914 (N_13914,N_13437,N_13135);
xnor U13915 (N_13915,N_13433,N_13485);
xor U13916 (N_13916,N_13246,N_13323);
and U13917 (N_13917,N_13190,N_13325);
nand U13918 (N_13918,N_13283,N_13192);
nand U13919 (N_13919,N_13107,N_13312);
nor U13920 (N_13920,N_13331,N_13031);
nor U13921 (N_13921,N_13098,N_13071);
or U13922 (N_13922,N_13106,N_13166);
xnor U13923 (N_13923,N_13252,N_13214);
and U13924 (N_13924,N_13245,N_13285);
nor U13925 (N_13925,N_13350,N_13049);
and U13926 (N_13926,N_13244,N_13159);
nor U13927 (N_13927,N_13472,N_13024);
nor U13928 (N_13928,N_13349,N_13330);
nor U13929 (N_13929,N_13492,N_13167);
or U13930 (N_13930,N_13158,N_13082);
nand U13931 (N_13931,N_13472,N_13128);
and U13932 (N_13932,N_13020,N_13225);
xor U13933 (N_13933,N_13182,N_13003);
nand U13934 (N_13934,N_13120,N_13492);
and U13935 (N_13935,N_13471,N_13402);
and U13936 (N_13936,N_13247,N_13002);
nand U13937 (N_13937,N_13408,N_13436);
and U13938 (N_13938,N_13191,N_13309);
nand U13939 (N_13939,N_13053,N_13481);
and U13940 (N_13940,N_13172,N_13167);
nor U13941 (N_13941,N_13346,N_13224);
nor U13942 (N_13942,N_13000,N_13107);
and U13943 (N_13943,N_13069,N_13066);
nand U13944 (N_13944,N_13486,N_13145);
and U13945 (N_13945,N_13353,N_13023);
and U13946 (N_13946,N_13126,N_13310);
and U13947 (N_13947,N_13446,N_13004);
and U13948 (N_13948,N_13222,N_13275);
or U13949 (N_13949,N_13203,N_13350);
xor U13950 (N_13950,N_13063,N_13140);
nor U13951 (N_13951,N_13002,N_13342);
nand U13952 (N_13952,N_13092,N_13110);
and U13953 (N_13953,N_13248,N_13227);
and U13954 (N_13954,N_13207,N_13346);
xnor U13955 (N_13955,N_13344,N_13309);
nand U13956 (N_13956,N_13498,N_13333);
xnor U13957 (N_13957,N_13067,N_13075);
nand U13958 (N_13958,N_13231,N_13359);
or U13959 (N_13959,N_13329,N_13169);
and U13960 (N_13960,N_13438,N_13462);
nand U13961 (N_13961,N_13259,N_13459);
and U13962 (N_13962,N_13113,N_13477);
and U13963 (N_13963,N_13389,N_13013);
xnor U13964 (N_13964,N_13371,N_13342);
nand U13965 (N_13965,N_13388,N_13327);
and U13966 (N_13966,N_13434,N_13287);
nand U13967 (N_13967,N_13406,N_13418);
and U13968 (N_13968,N_13430,N_13461);
and U13969 (N_13969,N_13028,N_13240);
or U13970 (N_13970,N_13294,N_13419);
nand U13971 (N_13971,N_13083,N_13151);
and U13972 (N_13972,N_13322,N_13141);
xnor U13973 (N_13973,N_13030,N_13373);
nor U13974 (N_13974,N_13429,N_13231);
nand U13975 (N_13975,N_13248,N_13212);
or U13976 (N_13976,N_13333,N_13432);
or U13977 (N_13977,N_13279,N_13204);
nand U13978 (N_13978,N_13078,N_13074);
xnor U13979 (N_13979,N_13077,N_13213);
nand U13980 (N_13980,N_13057,N_13481);
and U13981 (N_13981,N_13327,N_13067);
xnor U13982 (N_13982,N_13372,N_13044);
xnor U13983 (N_13983,N_13043,N_13274);
and U13984 (N_13984,N_13180,N_13360);
xnor U13985 (N_13985,N_13035,N_13400);
nand U13986 (N_13986,N_13225,N_13201);
nand U13987 (N_13987,N_13470,N_13230);
and U13988 (N_13988,N_13045,N_13067);
xnor U13989 (N_13989,N_13165,N_13406);
nand U13990 (N_13990,N_13163,N_13024);
nor U13991 (N_13991,N_13189,N_13147);
nand U13992 (N_13992,N_13478,N_13424);
or U13993 (N_13993,N_13229,N_13198);
or U13994 (N_13994,N_13017,N_13105);
xor U13995 (N_13995,N_13432,N_13302);
nand U13996 (N_13996,N_13183,N_13322);
xnor U13997 (N_13997,N_13043,N_13492);
and U13998 (N_13998,N_13497,N_13041);
nor U13999 (N_13999,N_13252,N_13331);
and U14000 (N_14000,N_13591,N_13799);
nand U14001 (N_14001,N_13550,N_13642);
nor U14002 (N_14002,N_13569,N_13778);
nor U14003 (N_14003,N_13938,N_13983);
and U14004 (N_14004,N_13653,N_13795);
and U14005 (N_14005,N_13792,N_13524);
nand U14006 (N_14006,N_13730,N_13510);
or U14007 (N_14007,N_13600,N_13726);
or U14008 (N_14008,N_13901,N_13568);
xor U14009 (N_14009,N_13800,N_13880);
or U14010 (N_14010,N_13749,N_13863);
xnor U14011 (N_14011,N_13574,N_13849);
and U14012 (N_14012,N_13713,N_13545);
and U14013 (N_14013,N_13665,N_13556);
nand U14014 (N_14014,N_13514,N_13715);
nor U14015 (N_14015,N_13826,N_13626);
and U14016 (N_14016,N_13567,N_13807);
or U14017 (N_14017,N_13821,N_13531);
and U14018 (N_14018,N_13672,N_13752);
and U14019 (N_14019,N_13994,N_13644);
and U14020 (N_14020,N_13618,N_13595);
xnor U14021 (N_14021,N_13991,N_13534);
nor U14022 (N_14022,N_13903,N_13918);
or U14023 (N_14023,N_13636,N_13561);
nand U14024 (N_14024,N_13937,N_13558);
nand U14025 (N_14025,N_13537,N_13695);
nand U14026 (N_14026,N_13520,N_13746);
or U14027 (N_14027,N_13607,N_13592);
xnor U14028 (N_14028,N_13835,N_13815);
xnor U14029 (N_14029,N_13980,N_13616);
xor U14030 (N_14030,N_13624,N_13861);
nor U14031 (N_14031,N_13608,N_13717);
xor U14032 (N_14032,N_13610,N_13984);
or U14033 (N_14033,N_13614,N_13620);
nand U14034 (N_14034,N_13544,N_13963);
xor U14035 (N_14035,N_13612,N_13705);
nor U14036 (N_14036,N_13742,N_13660);
xnor U14037 (N_14037,N_13707,N_13874);
and U14038 (N_14038,N_13511,N_13629);
or U14039 (N_14039,N_13602,N_13768);
and U14040 (N_14040,N_13504,N_13690);
nor U14041 (N_14041,N_13968,N_13704);
xnor U14042 (N_14042,N_13725,N_13748);
and U14043 (N_14043,N_13606,N_13936);
and U14044 (N_14044,N_13577,N_13522);
nand U14045 (N_14045,N_13689,N_13883);
and U14046 (N_14046,N_13621,N_13506);
or U14047 (N_14047,N_13663,N_13895);
xor U14048 (N_14048,N_13584,N_13623);
or U14049 (N_14049,N_13759,N_13528);
and U14050 (N_14050,N_13908,N_13915);
xnor U14051 (N_14051,N_13617,N_13747);
nor U14052 (N_14052,N_13942,N_13944);
or U14053 (N_14053,N_13559,N_13879);
xnor U14054 (N_14054,N_13538,N_13836);
xor U14055 (N_14055,N_13886,N_13519);
and U14056 (N_14056,N_13875,N_13699);
and U14057 (N_14057,N_13666,N_13535);
xor U14058 (N_14058,N_13590,N_13774);
or U14059 (N_14059,N_13987,N_13572);
nor U14060 (N_14060,N_13667,N_13896);
or U14061 (N_14061,N_13654,N_13831);
or U14062 (N_14062,N_13700,N_13714);
nand U14063 (N_14063,N_13685,N_13563);
and U14064 (N_14064,N_13503,N_13662);
and U14065 (N_14065,N_13767,N_13952);
and U14066 (N_14066,N_13913,N_13683);
nor U14067 (N_14067,N_13619,N_13775);
and U14068 (N_14068,N_13907,N_13884);
nor U14069 (N_14069,N_13583,N_13659);
xnor U14070 (N_14070,N_13854,N_13540);
xnor U14071 (N_14071,N_13601,N_13694);
or U14072 (N_14072,N_13817,N_13744);
nand U14073 (N_14073,N_13736,N_13575);
nand U14074 (N_14074,N_13548,N_13627);
or U14075 (N_14075,N_13541,N_13904);
xor U14076 (N_14076,N_13931,N_13939);
nor U14077 (N_14077,N_13959,N_13684);
or U14078 (N_14078,N_13894,N_13703);
nand U14079 (N_14079,N_13679,N_13811);
and U14080 (N_14080,N_13961,N_13677);
nand U14081 (N_14081,N_13993,N_13941);
nand U14082 (N_14082,N_13737,N_13738);
and U14083 (N_14083,N_13710,N_13878);
or U14084 (N_14084,N_13518,N_13929);
and U14085 (N_14085,N_13691,N_13582);
or U14086 (N_14086,N_13765,N_13631);
and U14087 (N_14087,N_13755,N_13926);
or U14088 (N_14088,N_13822,N_13841);
xor U14089 (N_14089,N_13740,N_13638);
and U14090 (N_14090,N_13928,N_13674);
or U14091 (N_14091,N_13647,N_13932);
and U14092 (N_14092,N_13507,N_13851);
xor U14093 (N_14093,N_13566,N_13789);
and U14094 (N_14094,N_13523,N_13825);
nand U14095 (N_14095,N_13787,N_13578);
nor U14096 (N_14096,N_13530,N_13870);
and U14097 (N_14097,N_13508,N_13852);
and U14098 (N_14098,N_13943,N_13670);
or U14099 (N_14099,N_13734,N_13933);
or U14100 (N_14100,N_13656,N_13900);
or U14101 (N_14101,N_13948,N_13827);
and U14102 (N_14102,N_13697,N_13971);
or U14103 (N_14103,N_13598,N_13946);
and U14104 (N_14104,N_13754,N_13805);
or U14105 (N_14105,N_13760,N_13888);
and U14106 (N_14106,N_13719,N_13573);
and U14107 (N_14107,N_13887,N_13848);
or U14108 (N_14108,N_13988,N_13945);
nand U14109 (N_14109,N_13824,N_13844);
or U14110 (N_14110,N_13625,N_13965);
nor U14111 (N_14111,N_13500,N_13972);
xnor U14112 (N_14112,N_13655,N_13585);
nor U14113 (N_14113,N_13910,N_13532);
xnor U14114 (N_14114,N_13909,N_13557);
nand U14115 (N_14115,N_13846,N_13711);
nor U14116 (N_14116,N_13635,N_13833);
and U14117 (N_14117,N_13688,N_13978);
xnor U14118 (N_14118,N_13989,N_13969);
nand U14119 (N_14119,N_13889,N_13814);
xnor U14120 (N_14120,N_13505,N_13513);
nor U14121 (N_14121,N_13798,N_13763);
xnor U14122 (N_14122,N_13935,N_13858);
xnor U14123 (N_14123,N_13893,N_13772);
xor U14124 (N_14124,N_13553,N_13560);
nor U14125 (N_14125,N_13562,N_13862);
or U14126 (N_14126,N_13839,N_13735);
nor U14127 (N_14127,N_13727,N_13751);
nor U14128 (N_14128,N_13588,N_13554);
or U14129 (N_14129,N_13603,N_13790);
nor U14130 (N_14130,N_13865,N_13641);
nor U14131 (N_14131,N_13784,N_13985);
nand U14132 (N_14132,N_13581,N_13974);
or U14133 (N_14133,N_13834,N_13917);
nor U14134 (N_14134,N_13611,N_13533);
nor U14135 (N_14135,N_13649,N_13840);
nand U14136 (N_14136,N_13958,N_13867);
xnor U14137 (N_14137,N_13664,N_13905);
nor U14138 (N_14138,N_13501,N_13823);
nor U14139 (N_14139,N_13812,N_13853);
and U14140 (N_14140,N_13843,N_13990);
xnor U14141 (N_14141,N_13552,N_13709);
nand U14142 (N_14142,N_13829,N_13813);
nor U14143 (N_14143,N_13605,N_13995);
or U14144 (N_14144,N_13922,N_13962);
nand U14145 (N_14145,N_13783,N_13919);
xnor U14146 (N_14146,N_13809,N_13599);
or U14147 (N_14147,N_13830,N_13788);
nor U14148 (N_14148,N_13766,N_13847);
nand U14149 (N_14149,N_13973,N_13930);
and U14150 (N_14150,N_13956,N_13819);
xor U14151 (N_14151,N_13837,N_13885);
or U14152 (N_14152,N_13587,N_13576);
or U14153 (N_14153,N_13701,N_13925);
nand U14154 (N_14154,N_13687,N_13871);
nor U14155 (N_14155,N_13923,N_13542);
and U14156 (N_14156,N_13992,N_13640);
nor U14157 (N_14157,N_13634,N_13845);
nand U14158 (N_14158,N_13881,N_13977);
or U14159 (N_14159,N_13982,N_13517);
nand U14160 (N_14160,N_13756,N_13571);
and U14161 (N_14161,N_13912,N_13949);
and U14162 (N_14162,N_13536,N_13806);
nand U14163 (N_14163,N_13579,N_13820);
xnor U14164 (N_14164,N_13782,N_13686);
nor U14165 (N_14165,N_13914,N_13981);
xnor U14166 (N_14166,N_13764,N_13745);
xnor U14167 (N_14167,N_13869,N_13650);
xor U14168 (N_14168,N_13724,N_13967);
and U14169 (N_14169,N_13543,N_13779);
and U14170 (N_14170,N_13892,N_13808);
nor U14171 (N_14171,N_13791,N_13786);
nand U14172 (N_14172,N_13741,N_13777);
nand U14173 (N_14173,N_13856,N_13780);
or U14174 (N_14174,N_13934,N_13776);
or U14175 (N_14175,N_13630,N_13570);
xor U14176 (N_14176,N_13906,N_13940);
nand U14177 (N_14177,N_13521,N_13639);
or U14178 (N_14178,N_13743,N_13793);
xor U14179 (N_14179,N_13722,N_13996);
xnor U14180 (N_14180,N_13872,N_13997);
nand U14181 (N_14181,N_13731,N_13979);
or U14182 (N_14182,N_13729,N_13866);
nor U14183 (N_14183,N_13753,N_13525);
nand U14184 (N_14184,N_13868,N_13646);
nor U14185 (N_14185,N_13970,N_13564);
and U14186 (N_14186,N_13678,N_13950);
and U14187 (N_14187,N_13960,N_13924);
nand U14188 (N_14188,N_13897,N_13613);
nor U14189 (N_14189,N_13964,N_13502);
nand U14190 (N_14190,N_13515,N_13549);
or U14191 (N_14191,N_13916,N_13551);
xnor U14192 (N_14192,N_13951,N_13953);
nand U14193 (N_14193,N_13976,N_13658);
nand U14194 (N_14194,N_13668,N_13516);
nor U14195 (N_14195,N_13716,N_13855);
nand U14196 (N_14196,N_13721,N_13891);
nor U14197 (N_14197,N_13632,N_13604);
xor U14198 (N_14198,N_13818,N_13651);
nor U14199 (N_14199,N_13920,N_13850);
xnor U14200 (N_14200,N_13860,N_13758);
nand U14201 (N_14201,N_13899,N_13794);
nand U14202 (N_14202,N_13802,N_13999);
xnor U14203 (N_14203,N_13539,N_13546);
or U14204 (N_14204,N_13857,N_13615);
and U14205 (N_14205,N_13681,N_13586);
or U14206 (N_14206,N_13637,N_13609);
or U14207 (N_14207,N_13773,N_13547);
or U14208 (N_14208,N_13921,N_13902);
nand U14209 (N_14209,N_13770,N_13733);
xor U14210 (N_14210,N_13702,N_13810);
or U14211 (N_14211,N_13529,N_13565);
and U14212 (N_14212,N_13698,N_13757);
or U14213 (N_14213,N_13986,N_13652);
and U14214 (N_14214,N_13643,N_13890);
nor U14215 (N_14215,N_13512,N_13873);
or U14216 (N_14216,N_13526,N_13645);
xnor U14217 (N_14217,N_13859,N_13580);
nand U14218 (N_14218,N_13877,N_13955);
and U14219 (N_14219,N_13750,N_13696);
or U14220 (N_14220,N_13712,N_13594);
or U14221 (N_14221,N_13720,N_13803);
nor U14222 (N_14222,N_13828,N_13628);
or U14223 (N_14223,N_13954,N_13781);
and U14224 (N_14224,N_13975,N_13769);
and U14225 (N_14225,N_13801,N_13927);
nor U14226 (N_14226,N_13739,N_13680);
and U14227 (N_14227,N_13706,N_13596);
xnor U14228 (N_14228,N_13555,N_13796);
and U14229 (N_14229,N_13676,N_13797);
nor U14230 (N_14230,N_13723,N_13728);
and U14231 (N_14231,N_13657,N_13898);
and U14232 (N_14232,N_13673,N_13661);
or U14233 (N_14233,N_13771,N_13947);
nor U14234 (N_14234,N_13589,N_13911);
nand U14235 (N_14235,N_13671,N_13762);
xor U14236 (N_14236,N_13998,N_13882);
nand U14237 (N_14237,N_13597,N_13876);
or U14238 (N_14238,N_13648,N_13633);
and U14239 (N_14239,N_13838,N_13842);
and U14240 (N_14240,N_13957,N_13708);
and U14241 (N_14241,N_13527,N_13622);
or U14242 (N_14242,N_13509,N_13761);
and U14243 (N_14243,N_13816,N_13966);
or U14244 (N_14244,N_13593,N_13804);
nand U14245 (N_14245,N_13692,N_13732);
or U14246 (N_14246,N_13693,N_13669);
nand U14247 (N_14247,N_13785,N_13718);
and U14248 (N_14248,N_13864,N_13675);
nand U14249 (N_14249,N_13832,N_13682);
or U14250 (N_14250,N_13957,N_13513);
or U14251 (N_14251,N_13739,N_13508);
and U14252 (N_14252,N_13531,N_13999);
and U14253 (N_14253,N_13834,N_13634);
and U14254 (N_14254,N_13886,N_13677);
nor U14255 (N_14255,N_13594,N_13659);
nor U14256 (N_14256,N_13683,N_13729);
xnor U14257 (N_14257,N_13524,N_13544);
xnor U14258 (N_14258,N_13726,N_13573);
nor U14259 (N_14259,N_13692,N_13672);
nor U14260 (N_14260,N_13667,N_13551);
or U14261 (N_14261,N_13783,N_13889);
and U14262 (N_14262,N_13932,N_13876);
nor U14263 (N_14263,N_13995,N_13641);
nand U14264 (N_14264,N_13503,N_13816);
xor U14265 (N_14265,N_13988,N_13859);
nor U14266 (N_14266,N_13662,N_13936);
and U14267 (N_14267,N_13857,N_13874);
nand U14268 (N_14268,N_13949,N_13544);
nand U14269 (N_14269,N_13617,N_13784);
nor U14270 (N_14270,N_13561,N_13968);
or U14271 (N_14271,N_13620,N_13622);
nand U14272 (N_14272,N_13942,N_13974);
and U14273 (N_14273,N_13711,N_13952);
nand U14274 (N_14274,N_13611,N_13526);
and U14275 (N_14275,N_13809,N_13792);
or U14276 (N_14276,N_13649,N_13832);
or U14277 (N_14277,N_13977,N_13785);
nor U14278 (N_14278,N_13952,N_13915);
nand U14279 (N_14279,N_13888,N_13940);
nand U14280 (N_14280,N_13560,N_13642);
or U14281 (N_14281,N_13609,N_13639);
xor U14282 (N_14282,N_13875,N_13587);
xnor U14283 (N_14283,N_13866,N_13827);
and U14284 (N_14284,N_13798,N_13676);
and U14285 (N_14285,N_13501,N_13616);
and U14286 (N_14286,N_13972,N_13942);
nor U14287 (N_14287,N_13999,N_13513);
nand U14288 (N_14288,N_13937,N_13670);
nand U14289 (N_14289,N_13752,N_13930);
or U14290 (N_14290,N_13961,N_13796);
xnor U14291 (N_14291,N_13507,N_13972);
nor U14292 (N_14292,N_13679,N_13742);
and U14293 (N_14293,N_13788,N_13626);
and U14294 (N_14294,N_13565,N_13731);
and U14295 (N_14295,N_13523,N_13605);
nand U14296 (N_14296,N_13921,N_13972);
or U14297 (N_14297,N_13790,N_13526);
xor U14298 (N_14298,N_13991,N_13963);
and U14299 (N_14299,N_13760,N_13660);
and U14300 (N_14300,N_13998,N_13607);
nand U14301 (N_14301,N_13999,N_13594);
nand U14302 (N_14302,N_13792,N_13991);
nor U14303 (N_14303,N_13657,N_13979);
xnor U14304 (N_14304,N_13643,N_13917);
or U14305 (N_14305,N_13825,N_13577);
nor U14306 (N_14306,N_13772,N_13797);
nand U14307 (N_14307,N_13804,N_13890);
nand U14308 (N_14308,N_13598,N_13747);
nand U14309 (N_14309,N_13627,N_13777);
xnor U14310 (N_14310,N_13704,N_13828);
nor U14311 (N_14311,N_13744,N_13583);
nor U14312 (N_14312,N_13956,N_13929);
and U14313 (N_14313,N_13534,N_13953);
nor U14314 (N_14314,N_13925,N_13751);
and U14315 (N_14315,N_13686,N_13875);
and U14316 (N_14316,N_13500,N_13521);
and U14317 (N_14317,N_13576,N_13817);
nor U14318 (N_14318,N_13966,N_13885);
nor U14319 (N_14319,N_13577,N_13518);
xor U14320 (N_14320,N_13752,N_13502);
xor U14321 (N_14321,N_13911,N_13779);
nand U14322 (N_14322,N_13826,N_13615);
and U14323 (N_14323,N_13676,N_13984);
xnor U14324 (N_14324,N_13671,N_13644);
xnor U14325 (N_14325,N_13881,N_13643);
and U14326 (N_14326,N_13692,N_13778);
or U14327 (N_14327,N_13526,N_13878);
nand U14328 (N_14328,N_13828,N_13565);
nand U14329 (N_14329,N_13718,N_13771);
or U14330 (N_14330,N_13734,N_13818);
and U14331 (N_14331,N_13929,N_13546);
or U14332 (N_14332,N_13962,N_13964);
or U14333 (N_14333,N_13934,N_13528);
xor U14334 (N_14334,N_13680,N_13888);
or U14335 (N_14335,N_13645,N_13852);
or U14336 (N_14336,N_13953,N_13947);
nand U14337 (N_14337,N_13946,N_13836);
nor U14338 (N_14338,N_13853,N_13769);
xnor U14339 (N_14339,N_13549,N_13851);
or U14340 (N_14340,N_13673,N_13964);
nor U14341 (N_14341,N_13739,N_13671);
nor U14342 (N_14342,N_13810,N_13800);
nand U14343 (N_14343,N_13572,N_13959);
nor U14344 (N_14344,N_13702,N_13880);
nand U14345 (N_14345,N_13692,N_13972);
xnor U14346 (N_14346,N_13540,N_13568);
xor U14347 (N_14347,N_13545,N_13572);
and U14348 (N_14348,N_13814,N_13709);
xnor U14349 (N_14349,N_13823,N_13876);
xnor U14350 (N_14350,N_13810,N_13779);
xor U14351 (N_14351,N_13990,N_13981);
xnor U14352 (N_14352,N_13770,N_13785);
and U14353 (N_14353,N_13822,N_13928);
or U14354 (N_14354,N_13816,N_13887);
and U14355 (N_14355,N_13859,N_13983);
xnor U14356 (N_14356,N_13724,N_13953);
nand U14357 (N_14357,N_13691,N_13591);
or U14358 (N_14358,N_13706,N_13717);
xnor U14359 (N_14359,N_13867,N_13724);
nor U14360 (N_14360,N_13808,N_13536);
nor U14361 (N_14361,N_13800,N_13663);
and U14362 (N_14362,N_13614,N_13973);
xor U14363 (N_14363,N_13750,N_13700);
or U14364 (N_14364,N_13984,N_13849);
nor U14365 (N_14365,N_13938,N_13788);
and U14366 (N_14366,N_13951,N_13794);
nand U14367 (N_14367,N_13643,N_13951);
and U14368 (N_14368,N_13682,N_13544);
nor U14369 (N_14369,N_13896,N_13582);
nand U14370 (N_14370,N_13951,N_13725);
xor U14371 (N_14371,N_13500,N_13724);
or U14372 (N_14372,N_13769,N_13761);
xnor U14373 (N_14373,N_13894,N_13828);
nand U14374 (N_14374,N_13883,N_13701);
and U14375 (N_14375,N_13562,N_13743);
nor U14376 (N_14376,N_13868,N_13802);
and U14377 (N_14377,N_13609,N_13682);
nand U14378 (N_14378,N_13511,N_13772);
or U14379 (N_14379,N_13528,N_13918);
nor U14380 (N_14380,N_13827,N_13685);
nor U14381 (N_14381,N_13621,N_13829);
or U14382 (N_14382,N_13571,N_13994);
or U14383 (N_14383,N_13866,N_13764);
and U14384 (N_14384,N_13643,N_13929);
or U14385 (N_14385,N_13621,N_13945);
xor U14386 (N_14386,N_13670,N_13628);
or U14387 (N_14387,N_13560,N_13927);
nand U14388 (N_14388,N_13744,N_13675);
nand U14389 (N_14389,N_13579,N_13615);
nand U14390 (N_14390,N_13613,N_13964);
nand U14391 (N_14391,N_13873,N_13584);
nand U14392 (N_14392,N_13848,N_13927);
and U14393 (N_14393,N_13911,N_13635);
and U14394 (N_14394,N_13638,N_13546);
nand U14395 (N_14395,N_13761,N_13873);
nor U14396 (N_14396,N_13878,N_13839);
nor U14397 (N_14397,N_13675,N_13814);
xnor U14398 (N_14398,N_13599,N_13876);
nor U14399 (N_14399,N_13971,N_13571);
xnor U14400 (N_14400,N_13939,N_13532);
xor U14401 (N_14401,N_13901,N_13823);
nor U14402 (N_14402,N_13779,N_13613);
nand U14403 (N_14403,N_13933,N_13930);
nor U14404 (N_14404,N_13762,N_13770);
or U14405 (N_14405,N_13692,N_13844);
nand U14406 (N_14406,N_13738,N_13995);
and U14407 (N_14407,N_13899,N_13809);
or U14408 (N_14408,N_13557,N_13550);
nor U14409 (N_14409,N_13759,N_13993);
nand U14410 (N_14410,N_13982,N_13661);
xor U14411 (N_14411,N_13705,N_13591);
nand U14412 (N_14412,N_13862,N_13735);
and U14413 (N_14413,N_13573,N_13659);
nand U14414 (N_14414,N_13601,N_13714);
xor U14415 (N_14415,N_13873,N_13733);
or U14416 (N_14416,N_13510,N_13585);
nand U14417 (N_14417,N_13889,N_13539);
and U14418 (N_14418,N_13500,N_13743);
xnor U14419 (N_14419,N_13720,N_13701);
nor U14420 (N_14420,N_13827,N_13864);
nor U14421 (N_14421,N_13952,N_13585);
and U14422 (N_14422,N_13625,N_13948);
nand U14423 (N_14423,N_13541,N_13693);
or U14424 (N_14424,N_13641,N_13566);
or U14425 (N_14425,N_13810,N_13716);
or U14426 (N_14426,N_13788,N_13721);
nand U14427 (N_14427,N_13940,N_13920);
or U14428 (N_14428,N_13928,N_13631);
nand U14429 (N_14429,N_13616,N_13599);
and U14430 (N_14430,N_13934,N_13971);
nor U14431 (N_14431,N_13693,N_13915);
or U14432 (N_14432,N_13906,N_13844);
xnor U14433 (N_14433,N_13761,N_13739);
and U14434 (N_14434,N_13723,N_13680);
nand U14435 (N_14435,N_13910,N_13974);
or U14436 (N_14436,N_13879,N_13744);
or U14437 (N_14437,N_13863,N_13703);
nor U14438 (N_14438,N_13860,N_13718);
or U14439 (N_14439,N_13865,N_13629);
and U14440 (N_14440,N_13700,N_13518);
nor U14441 (N_14441,N_13596,N_13855);
and U14442 (N_14442,N_13550,N_13687);
xnor U14443 (N_14443,N_13691,N_13800);
or U14444 (N_14444,N_13989,N_13948);
nand U14445 (N_14445,N_13960,N_13829);
nor U14446 (N_14446,N_13848,N_13766);
xnor U14447 (N_14447,N_13525,N_13572);
nand U14448 (N_14448,N_13994,N_13639);
or U14449 (N_14449,N_13669,N_13608);
nor U14450 (N_14450,N_13576,N_13654);
nor U14451 (N_14451,N_13526,N_13977);
nand U14452 (N_14452,N_13820,N_13780);
xor U14453 (N_14453,N_13864,N_13586);
nor U14454 (N_14454,N_13711,N_13621);
and U14455 (N_14455,N_13656,N_13523);
nand U14456 (N_14456,N_13850,N_13674);
and U14457 (N_14457,N_13835,N_13728);
nand U14458 (N_14458,N_13940,N_13545);
xor U14459 (N_14459,N_13562,N_13674);
xnor U14460 (N_14460,N_13597,N_13810);
nor U14461 (N_14461,N_13741,N_13935);
xor U14462 (N_14462,N_13957,N_13915);
nand U14463 (N_14463,N_13780,N_13880);
or U14464 (N_14464,N_13837,N_13798);
nand U14465 (N_14465,N_13965,N_13984);
nor U14466 (N_14466,N_13561,N_13923);
nand U14467 (N_14467,N_13682,N_13751);
nand U14468 (N_14468,N_13909,N_13569);
or U14469 (N_14469,N_13689,N_13590);
xnor U14470 (N_14470,N_13915,N_13704);
xor U14471 (N_14471,N_13517,N_13651);
or U14472 (N_14472,N_13570,N_13876);
xnor U14473 (N_14473,N_13864,N_13926);
or U14474 (N_14474,N_13553,N_13659);
or U14475 (N_14475,N_13958,N_13807);
or U14476 (N_14476,N_13743,N_13894);
or U14477 (N_14477,N_13697,N_13517);
nand U14478 (N_14478,N_13684,N_13941);
xnor U14479 (N_14479,N_13548,N_13614);
or U14480 (N_14480,N_13854,N_13798);
and U14481 (N_14481,N_13598,N_13550);
and U14482 (N_14482,N_13844,N_13527);
nand U14483 (N_14483,N_13839,N_13817);
nor U14484 (N_14484,N_13701,N_13764);
nor U14485 (N_14485,N_13959,N_13784);
nand U14486 (N_14486,N_13993,N_13916);
nand U14487 (N_14487,N_13735,N_13924);
and U14488 (N_14488,N_13801,N_13618);
xor U14489 (N_14489,N_13661,N_13616);
or U14490 (N_14490,N_13699,N_13592);
or U14491 (N_14491,N_13980,N_13969);
nor U14492 (N_14492,N_13540,N_13589);
xor U14493 (N_14493,N_13617,N_13526);
xnor U14494 (N_14494,N_13956,N_13874);
or U14495 (N_14495,N_13778,N_13531);
or U14496 (N_14496,N_13860,N_13909);
nand U14497 (N_14497,N_13560,N_13599);
nand U14498 (N_14498,N_13905,N_13779);
and U14499 (N_14499,N_13820,N_13704);
and U14500 (N_14500,N_14319,N_14392);
and U14501 (N_14501,N_14484,N_14083);
nor U14502 (N_14502,N_14120,N_14329);
nor U14503 (N_14503,N_14087,N_14433);
nor U14504 (N_14504,N_14119,N_14448);
or U14505 (N_14505,N_14275,N_14345);
or U14506 (N_14506,N_14487,N_14341);
nand U14507 (N_14507,N_14270,N_14452);
xnor U14508 (N_14508,N_14092,N_14358);
and U14509 (N_14509,N_14113,N_14179);
xor U14510 (N_14510,N_14372,N_14408);
xor U14511 (N_14511,N_14430,N_14055);
nand U14512 (N_14512,N_14272,N_14035);
or U14513 (N_14513,N_14236,N_14114);
or U14514 (N_14514,N_14378,N_14042);
nand U14515 (N_14515,N_14160,N_14432);
and U14516 (N_14516,N_14200,N_14024);
nor U14517 (N_14517,N_14065,N_14108);
and U14518 (N_14518,N_14306,N_14124);
xor U14519 (N_14519,N_14205,N_14324);
xnor U14520 (N_14520,N_14285,N_14493);
nand U14521 (N_14521,N_14420,N_14398);
xor U14522 (N_14522,N_14362,N_14370);
or U14523 (N_14523,N_14048,N_14170);
or U14524 (N_14524,N_14497,N_14422);
and U14525 (N_14525,N_14058,N_14063);
nor U14526 (N_14526,N_14038,N_14053);
nor U14527 (N_14527,N_14061,N_14472);
nor U14528 (N_14528,N_14116,N_14198);
and U14529 (N_14529,N_14017,N_14415);
and U14530 (N_14530,N_14254,N_14054);
and U14531 (N_14531,N_14327,N_14330);
xor U14532 (N_14532,N_14246,N_14070);
nand U14533 (N_14533,N_14308,N_14156);
or U14534 (N_14534,N_14383,N_14148);
and U14535 (N_14535,N_14044,N_14269);
and U14536 (N_14536,N_14013,N_14001);
or U14537 (N_14537,N_14421,N_14371);
and U14538 (N_14538,N_14296,N_14142);
and U14539 (N_14539,N_14458,N_14043);
and U14540 (N_14540,N_14218,N_14459);
nor U14541 (N_14541,N_14460,N_14334);
and U14542 (N_14542,N_14299,N_14344);
nor U14543 (N_14543,N_14000,N_14014);
and U14544 (N_14544,N_14413,N_14313);
and U14545 (N_14545,N_14105,N_14090);
nand U14546 (N_14546,N_14078,N_14264);
nand U14547 (N_14547,N_14332,N_14258);
or U14548 (N_14548,N_14088,N_14248);
or U14549 (N_14549,N_14139,N_14361);
and U14550 (N_14550,N_14434,N_14294);
and U14551 (N_14551,N_14117,N_14208);
nand U14552 (N_14552,N_14195,N_14107);
nor U14553 (N_14553,N_14134,N_14436);
nand U14554 (N_14554,N_14473,N_14266);
xnor U14555 (N_14555,N_14225,N_14149);
and U14556 (N_14556,N_14192,N_14260);
nor U14557 (N_14557,N_14032,N_14278);
nor U14558 (N_14558,N_14019,N_14445);
nor U14559 (N_14559,N_14424,N_14310);
xnor U14560 (N_14560,N_14118,N_14396);
nand U14561 (N_14561,N_14253,N_14367);
nand U14562 (N_14562,N_14171,N_14315);
and U14563 (N_14563,N_14033,N_14259);
xnor U14564 (N_14564,N_14305,N_14402);
nand U14565 (N_14565,N_14106,N_14005);
nand U14566 (N_14566,N_14244,N_14464);
nand U14567 (N_14567,N_14261,N_14166);
nor U14568 (N_14568,N_14185,N_14293);
nand U14569 (N_14569,N_14158,N_14159);
xnor U14570 (N_14570,N_14303,N_14084);
or U14571 (N_14571,N_14176,N_14164);
xnor U14572 (N_14572,N_14110,N_14256);
nand U14573 (N_14573,N_14165,N_14197);
nand U14574 (N_14574,N_14446,N_14191);
nor U14575 (N_14575,N_14199,N_14438);
and U14576 (N_14576,N_14190,N_14414);
nand U14577 (N_14577,N_14389,N_14470);
nor U14578 (N_14578,N_14346,N_14444);
nand U14579 (N_14579,N_14382,N_14123);
or U14580 (N_14580,N_14461,N_14290);
xor U14581 (N_14581,N_14411,N_14468);
nor U14582 (N_14582,N_14137,N_14373);
nand U14583 (N_14583,N_14262,N_14220);
nand U14584 (N_14584,N_14209,N_14125);
nand U14585 (N_14585,N_14485,N_14477);
nand U14586 (N_14586,N_14186,N_14079);
xnor U14587 (N_14587,N_14064,N_14004);
or U14588 (N_14588,N_14219,N_14016);
or U14589 (N_14589,N_14152,N_14012);
nor U14590 (N_14590,N_14386,N_14251);
or U14591 (N_14591,N_14009,N_14155);
or U14592 (N_14592,N_14489,N_14126);
nand U14593 (N_14593,N_14034,N_14040);
or U14594 (N_14594,N_14355,N_14416);
and U14595 (N_14595,N_14214,N_14273);
xor U14596 (N_14596,N_14181,N_14026);
nor U14597 (N_14597,N_14075,N_14302);
nor U14598 (N_14598,N_14453,N_14011);
xnor U14599 (N_14599,N_14095,N_14428);
and U14600 (N_14600,N_14304,N_14404);
and U14601 (N_14601,N_14059,N_14103);
nand U14602 (N_14602,N_14437,N_14006);
xor U14603 (N_14603,N_14368,N_14284);
xor U14604 (N_14604,N_14224,N_14109);
or U14605 (N_14605,N_14086,N_14425);
nand U14606 (N_14606,N_14222,N_14154);
nor U14607 (N_14607,N_14474,N_14322);
and U14608 (N_14608,N_14068,N_14049);
nand U14609 (N_14609,N_14442,N_14057);
and U14610 (N_14610,N_14223,N_14463);
xor U14611 (N_14611,N_14317,N_14307);
and U14612 (N_14612,N_14288,N_14478);
nor U14613 (N_14613,N_14074,N_14394);
nand U14614 (N_14614,N_14077,N_14471);
and U14615 (N_14615,N_14316,N_14390);
and U14616 (N_14616,N_14029,N_14245);
and U14617 (N_14617,N_14216,N_14099);
nand U14618 (N_14618,N_14136,N_14320);
xor U14619 (N_14619,N_14406,N_14435);
and U14620 (N_14620,N_14357,N_14381);
xor U14621 (N_14621,N_14052,N_14080);
or U14622 (N_14622,N_14204,N_14311);
nand U14623 (N_14623,N_14169,N_14349);
nor U14624 (N_14624,N_14279,N_14265);
or U14625 (N_14625,N_14151,N_14462);
nand U14626 (N_14626,N_14291,N_14111);
nor U14627 (N_14627,N_14274,N_14309);
nor U14628 (N_14628,N_14020,N_14071);
nand U14629 (N_14629,N_14140,N_14342);
nand U14630 (N_14630,N_14187,N_14295);
or U14631 (N_14631,N_14393,N_14297);
nand U14632 (N_14632,N_14335,N_14115);
nor U14633 (N_14633,N_14096,N_14379);
or U14634 (N_14634,N_14385,N_14483);
nand U14635 (N_14635,N_14491,N_14359);
xor U14636 (N_14636,N_14128,N_14229);
xor U14637 (N_14637,N_14352,N_14351);
nor U14638 (N_14638,N_14321,N_14369);
nand U14639 (N_14639,N_14130,N_14069);
nor U14640 (N_14640,N_14135,N_14407);
nand U14641 (N_14641,N_14280,N_14364);
and U14642 (N_14642,N_14081,N_14097);
and U14643 (N_14643,N_14377,N_14481);
nor U14644 (N_14644,N_14289,N_14380);
nor U14645 (N_14645,N_14331,N_14237);
and U14646 (N_14646,N_14353,N_14443);
and U14647 (N_14647,N_14238,N_14467);
xnor U14648 (N_14648,N_14230,N_14374);
xnor U14649 (N_14649,N_14173,N_14091);
nand U14650 (N_14650,N_14363,N_14450);
or U14651 (N_14651,N_14384,N_14027);
nand U14652 (N_14652,N_14226,N_14480);
xnor U14653 (N_14653,N_14021,N_14490);
or U14654 (N_14654,N_14400,N_14283);
and U14655 (N_14655,N_14486,N_14131);
and U14656 (N_14656,N_14333,N_14066);
or U14657 (N_14657,N_14082,N_14440);
nand U14658 (N_14658,N_14465,N_14194);
nand U14659 (N_14659,N_14388,N_14073);
and U14660 (N_14660,N_14062,N_14039);
nand U14661 (N_14661,N_14180,N_14174);
nor U14662 (N_14662,N_14456,N_14144);
nand U14663 (N_14663,N_14401,N_14405);
xnor U14664 (N_14664,N_14498,N_14449);
nor U14665 (N_14665,N_14072,N_14045);
nand U14666 (N_14666,N_14277,N_14133);
or U14667 (N_14667,N_14231,N_14267);
and U14668 (N_14668,N_14094,N_14228);
nand U14669 (N_14669,N_14177,N_14161);
nand U14670 (N_14670,N_14469,N_14050);
nor U14671 (N_14671,N_14276,N_14494);
and U14672 (N_14672,N_14143,N_14201);
xnor U14673 (N_14673,N_14060,N_14010);
nor U14674 (N_14674,N_14356,N_14041);
and U14675 (N_14675,N_14350,N_14093);
or U14676 (N_14676,N_14112,N_14215);
nand U14677 (N_14677,N_14239,N_14046);
nand U14678 (N_14678,N_14211,N_14121);
nor U14679 (N_14679,N_14418,N_14429);
or U14680 (N_14680,N_14234,N_14475);
nor U14681 (N_14681,N_14292,N_14212);
or U14682 (N_14682,N_14492,N_14360);
and U14683 (N_14683,N_14188,N_14210);
nor U14684 (N_14684,N_14249,N_14347);
or U14685 (N_14685,N_14252,N_14221);
and U14686 (N_14686,N_14100,N_14202);
nand U14687 (N_14687,N_14397,N_14495);
nand U14688 (N_14688,N_14447,N_14240);
nand U14689 (N_14689,N_14376,N_14104);
nand U14690 (N_14690,N_14030,N_14287);
nor U14691 (N_14691,N_14184,N_14153);
and U14692 (N_14692,N_14089,N_14286);
xnor U14693 (N_14693,N_14337,N_14243);
or U14694 (N_14694,N_14301,N_14206);
or U14695 (N_14695,N_14051,N_14023);
nand U14696 (N_14696,N_14036,N_14399);
nand U14697 (N_14697,N_14423,N_14127);
nand U14698 (N_14698,N_14193,N_14003);
nand U14699 (N_14699,N_14348,N_14403);
and U14700 (N_14700,N_14235,N_14300);
or U14701 (N_14701,N_14076,N_14207);
and U14702 (N_14702,N_14325,N_14145);
or U14703 (N_14703,N_14085,N_14354);
or U14704 (N_14704,N_14499,N_14439);
nand U14705 (N_14705,N_14129,N_14168);
nor U14706 (N_14706,N_14451,N_14338);
xor U14707 (N_14707,N_14482,N_14203);
and U14708 (N_14708,N_14122,N_14183);
or U14709 (N_14709,N_14328,N_14141);
nor U14710 (N_14710,N_14028,N_14242);
xnor U14711 (N_14711,N_14454,N_14281);
nor U14712 (N_14712,N_14419,N_14326);
or U14713 (N_14713,N_14157,N_14025);
and U14714 (N_14714,N_14178,N_14182);
and U14715 (N_14715,N_14196,N_14189);
nand U14716 (N_14716,N_14412,N_14018);
or U14717 (N_14717,N_14339,N_14257);
and U14718 (N_14718,N_14431,N_14476);
xor U14719 (N_14719,N_14227,N_14015);
xor U14720 (N_14720,N_14255,N_14318);
or U14721 (N_14721,N_14479,N_14340);
or U14722 (N_14722,N_14008,N_14366);
and U14723 (N_14723,N_14213,N_14263);
or U14724 (N_14724,N_14175,N_14163);
xor U14725 (N_14725,N_14056,N_14037);
nor U14726 (N_14726,N_14047,N_14098);
or U14727 (N_14727,N_14336,N_14496);
nor U14728 (N_14728,N_14314,N_14375);
xor U14729 (N_14729,N_14323,N_14233);
nor U14730 (N_14730,N_14312,N_14007);
or U14731 (N_14731,N_14488,N_14391);
and U14732 (N_14732,N_14298,N_14167);
nand U14733 (N_14733,N_14146,N_14365);
nand U14734 (N_14734,N_14441,N_14247);
xor U14735 (N_14735,N_14101,N_14067);
or U14736 (N_14736,N_14162,N_14387);
and U14737 (N_14737,N_14150,N_14343);
nand U14738 (N_14738,N_14147,N_14022);
and U14739 (N_14739,N_14426,N_14031);
nand U14740 (N_14740,N_14250,N_14002);
xnor U14741 (N_14741,N_14282,N_14417);
nand U14742 (N_14742,N_14466,N_14172);
and U14743 (N_14743,N_14232,N_14268);
and U14744 (N_14744,N_14427,N_14395);
xor U14745 (N_14745,N_14410,N_14102);
nand U14746 (N_14746,N_14409,N_14271);
and U14747 (N_14747,N_14457,N_14241);
nand U14748 (N_14748,N_14132,N_14217);
or U14749 (N_14749,N_14138,N_14455);
nand U14750 (N_14750,N_14009,N_14300);
and U14751 (N_14751,N_14229,N_14194);
nor U14752 (N_14752,N_14434,N_14385);
and U14753 (N_14753,N_14278,N_14412);
nand U14754 (N_14754,N_14020,N_14286);
or U14755 (N_14755,N_14489,N_14322);
and U14756 (N_14756,N_14105,N_14452);
or U14757 (N_14757,N_14308,N_14006);
and U14758 (N_14758,N_14371,N_14175);
xor U14759 (N_14759,N_14449,N_14446);
and U14760 (N_14760,N_14221,N_14192);
and U14761 (N_14761,N_14393,N_14132);
or U14762 (N_14762,N_14402,N_14163);
and U14763 (N_14763,N_14118,N_14252);
xor U14764 (N_14764,N_14313,N_14143);
nand U14765 (N_14765,N_14077,N_14283);
xnor U14766 (N_14766,N_14017,N_14357);
and U14767 (N_14767,N_14027,N_14119);
nand U14768 (N_14768,N_14151,N_14129);
nor U14769 (N_14769,N_14013,N_14209);
xnor U14770 (N_14770,N_14128,N_14172);
xor U14771 (N_14771,N_14358,N_14437);
nand U14772 (N_14772,N_14443,N_14372);
or U14773 (N_14773,N_14082,N_14192);
or U14774 (N_14774,N_14319,N_14099);
nand U14775 (N_14775,N_14186,N_14295);
and U14776 (N_14776,N_14185,N_14102);
or U14777 (N_14777,N_14433,N_14042);
or U14778 (N_14778,N_14125,N_14033);
xnor U14779 (N_14779,N_14421,N_14217);
nand U14780 (N_14780,N_14071,N_14168);
xnor U14781 (N_14781,N_14223,N_14027);
nand U14782 (N_14782,N_14373,N_14221);
nor U14783 (N_14783,N_14003,N_14457);
nand U14784 (N_14784,N_14153,N_14355);
nor U14785 (N_14785,N_14206,N_14046);
and U14786 (N_14786,N_14088,N_14409);
nor U14787 (N_14787,N_14228,N_14379);
nor U14788 (N_14788,N_14183,N_14306);
or U14789 (N_14789,N_14123,N_14498);
or U14790 (N_14790,N_14441,N_14437);
nand U14791 (N_14791,N_14027,N_14177);
xnor U14792 (N_14792,N_14044,N_14334);
xor U14793 (N_14793,N_14325,N_14253);
and U14794 (N_14794,N_14294,N_14132);
nor U14795 (N_14795,N_14362,N_14366);
xor U14796 (N_14796,N_14344,N_14233);
xor U14797 (N_14797,N_14290,N_14434);
xor U14798 (N_14798,N_14030,N_14401);
nor U14799 (N_14799,N_14218,N_14196);
nor U14800 (N_14800,N_14107,N_14366);
xnor U14801 (N_14801,N_14083,N_14027);
or U14802 (N_14802,N_14150,N_14392);
or U14803 (N_14803,N_14091,N_14140);
or U14804 (N_14804,N_14160,N_14294);
nor U14805 (N_14805,N_14482,N_14217);
and U14806 (N_14806,N_14410,N_14012);
xnor U14807 (N_14807,N_14062,N_14077);
nand U14808 (N_14808,N_14422,N_14237);
nand U14809 (N_14809,N_14222,N_14336);
nand U14810 (N_14810,N_14087,N_14308);
or U14811 (N_14811,N_14387,N_14451);
and U14812 (N_14812,N_14273,N_14020);
and U14813 (N_14813,N_14208,N_14259);
and U14814 (N_14814,N_14013,N_14122);
nor U14815 (N_14815,N_14086,N_14052);
xor U14816 (N_14816,N_14266,N_14493);
nor U14817 (N_14817,N_14239,N_14391);
nor U14818 (N_14818,N_14156,N_14283);
or U14819 (N_14819,N_14418,N_14094);
and U14820 (N_14820,N_14090,N_14106);
nor U14821 (N_14821,N_14452,N_14159);
nor U14822 (N_14822,N_14426,N_14400);
or U14823 (N_14823,N_14150,N_14492);
xor U14824 (N_14824,N_14358,N_14436);
nand U14825 (N_14825,N_14020,N_14090);
nor U14826 (N_14826,N_14097,N_14078);
or U14827 (N_14827,N_14239,N_14357);
or U14828 (N_14828,N_14187,N_14105);
nand U14829 (N_14829,N_14360,N_14442);
nor U14830 (N_14830,N_14337,N_14197);
nor U14831 (N_14831,N_14242,N_14402);
or U14832 (N_14832,N_14329,N_14135);
or U14833 (N_14833,N_14442,N_14078);
and U14834 (N_14834,N_14351,N_14100);
nand U14835 (N_14835,N_14358,N_14047);
or U14836 (N_14836,N_14386,N_14327);
nor U14837 (N_14837,N_14257,N_14249);
nand U14838 (N_14838,N_14453,N_14402);
or U14839 (N_14839,N_14497,N_14489);
nand U14840 (N_14840,N_14066,N_14267);
nor U14841 (N_14841,N_14119,N_14223);
and U14842 (N_14842,N_14154,N_14103);
nor U14843 (N_14843,N_14070,N_14422);
nand U14844 (N_14844,N_14081,N_14437);
and U14845 (N_14845,N_14477,N_14102);
xnor U14846 (N_14846,N_14452,N_14173);
xnor U14847 (N_14847,N_14175,N_14019);
nor U14848 (N_14848,N_14181,N_14172);
nand U14849 (N_14849,N_14480,N_14159);
xor U14850 (N_14850,N_14109,N_14213);
or U14851 (N_14851,N_14405,N_14116);
nor U14852 (N_14852,N_14092,N_14405);
or U14853 (N_14853,N_14433,N_14459);
nor U14854 (N_14854,N_14454,N_14202);
or U14855 (N_14855,N_14242,N_14408);
and U14856 (N_14856,N_14217,N_14467);
or U14857 (N_14857,N_14144,N_14321);
and U14858 (N_14858,N_14408,N_14346);
xor U14859 (N_14859,N_14080,N_14397);
and U14860 (N_14860,N_14158,N_14022);
and U14861 (N_14861,N_14357,N_14263);
xor U14862 (N_14862,N_14045,N_14077);
and U14863 (N_14863,N_14446,N_14403);
nor U14864 (N_14864,N_14169,N_14201);
nand U14865 (N_14865,N_14414,N_14204);
nand U14866 (N_14866,N_14387,N_14083);
or U14867 (N_14867,N_14276,N_14095);
nor U14868 (N_14868,N_14157,N_14001);
nor U14869 (N_14869,N_14312,N_14271);
and U14870 (N_14870,N_14063,N_14352);
nand U14871 (N_14871,N_14337,N_14041);
nand U14872 (N_14872,N_14352,N_14381);
nor U14873 (N_14873,N_14300,N_14153);
nor U14874 (N_14874,N_14215,N_14447);
or U14875 (N_14875,N_14031,N_14065);
and U14876 (N_14876,N_14410,N_14266);
or U14877 (N_14877,N_14017,N_14366);
nor U14878 (N_14878,N_14450,N_14228);
nand U14879 (N_14879,N_14147,N_14134);
xor U14880 (N_14880,N_14220,N_14092);
nor U14881 (N_14881,N_14224,N_14156);
nand U14882 (N_14882,N_14175,N_14126);
nor U14883 (N_14883,N_14343,N_14186);
and U14884 (N_14884,N_14297,N_14324);
or U14885 (N_14885,N_14390,N_14338);
xor U14886 (N_14886,N_14328,N_14288);
nand U14887 (N_14887,N_14283,N_14014);
xnor U14888 (N_14888,N_14202,N_14043);
nand U14889 (N_14889,N_14295,N_14390);
nor U14890 (N_14890,N_14075,N_14398);
nand U14891 (N_14891,N_14358,N_14381);
nand U14892 (N_14892,N_14081,N_14024);
and U14893 (N_14893,N_14237,N_14344);
or U14894 (N_14894,N_14176,N_14452);
or U14895 (N_14895,N_14159,N_14050);
or U14896 (N_14896,N_14075,N_14497);
xor U14897 (N_14897,N_14137,N_14468);
or U14898 (N_14898,N_14234,N_14173);
nor U14899 (N_14899,N_14145,N_14279);
or U14900 (N_14900,N_14035,N_14256);
xor U14901 (N_14901,N_14410,N_14365);
and U14902 (N_14902,N_14454,N_14116);
nor U14903 (N_14903,N_14494,N_14018);
nor U14904 (N_14904,N_14274,N_14490);
and U14905 (N_14905,N_14199,N_14284);
nand U14906 (N_14906,N_14372,N_14138);
xnor U14907 (N_14907,N_14191,N_14145);
nor U14908 (N_14908,N_14008,N_14051);
xnor U14909 (N_14909,N_14044,N_14276);
nand U14910 (N_14910,N_14299,N_14484);
nor U14911 (N_14911,N_14359,N_14128);
nor U14912 (N_14912,N_14435,N_14426);
nand U14913 (N_14913,N_14143,N_14401);
and U14914 (N_14914,N_14287,N_14065);
nand U14915 (N_14915,N_14418,N_14470);
or U14916 (N_14916,N_14309,N_14289);
nor U14917 (N_14917,N_14246,N_14003);
nor U14918 (N_14918,N_14459,N_14200);
nor U14919 (N_14919,N_14479,N_14141);
and U14920 (N_14920,N_14466,N_14363);
or U14921 (N_14921,N_14128,N_14444);
nor U14922 (N_14922,N_14440,N_14436);
or U14923 (N_14923,N_14461,N_14427);
nand U14924 (N_14924,N_14374,N_14119);
nand U14925 (N_14925,N_14375,N_14052);
or U14926 (N_14926,N_14486,N_14283);
xor U14927 (N_14927,N_14063,N_14286);
nand U14928 (N_14928,N_14235,N_14440);
and U14929 (N_14929,N_14049,N_14228);
nand U14930 (N_14930,N_14130,N_14101);
nand U14931 (N_14931,N_14009,N_14411);
and U14932 (N_14932,N_14287,N_14350);
nand U14933 (N_14933,N_14060,N_14253);
nand U14934 (N_14934,N_14354,N_14292);
xor U14935 (N_14935,N_14084,N_14313);
nor U14936 (N_14936,N_14068,N_14150);
nor U14937 (N_14937,N_14191,N_14048);
nand U14938 (N_14938,N_14044,N_14466);
nand U14939 (N_14939,N_14332,N_14207);
nand U14940 (N_14940,N_14079,N_14137);
nand U14941 (N_14941,N_14419,N_14435);
or U14942 (N_14942,N_14357,N_14050);
nor U14943 (N_14943,N_14039,N_14063);
nor U14944 (N_14944,N_14311,N_14435);
or U14945 (N_14945,N_14285,N_14066);
nor U14946 (N_14946,N_14477,N_14412);
and U14947 (N_14947,N_14327,N_14356);
nand U14948 (N_14948,N_14326,N_14288);
nand U14949 (N_14949,N_14309,N_14294);
and U14950 (N_14950,N_14084,N_14046);
nand U14951 (N_14951,N_14362,N_14257);
or U14952 (N_14952,N_14416,N_14409);
nand U14953 (N_14953,N_14457,N_14042);
or U14954 (N_14954,N_14013,N_14307);
and U14955 (N_14955,N_14105,N_14242);
nand U14956 (N_14956,N_14053,N_14410);
nand U14957 (N_14957,N_14218,N_14030);
and U14958 (N_14958,N_14250,N_14210);
nor U14959 (N_14959,N_14177,N_14261);
nand U14960 (N_14960,N_14038,N_14112);
xnor U14961 (N_14961,N_14465,N_14329);
and U14962 (N_14962,N_14262,N_14025);
xor U14963 (N_14963,N_14374,N_14450);
or U14964 (N_14964,N_14484,N_14087);
or U14965 (N_14965,N_14256,N_14034);
or U14966 (N_14966,N_14090,N_14212);
or U14967 (N_14967,N_14490,N_14246);
and U14968 (N_14968,N_14052,N_14157);
nor U14969 (N_14969,N_14430,N_14020);
nor U14970 (N_14970,N_14192,N_14228);
or U14971 (N_14971,N_14318,N_14193);
and U14972 (N_14972,N_14047,N_14105);
or U14973 (N_14973,N_14210,N_14180);
or U14974 (N_14974,N_14419,N_14252);
and U14975 (N_14975,N_14375,N_14093);
xnor U14976 (N_14976,N_14423,N_14292);
and U14977 (N_14977,N_14131,N_14035);
nand U14978 (N_14978,N_14105,N_14133);
or U14979 (N_14979,N_14162,N_14498);
and U14980 (N_14980,N_14238,N_14044);
and U14981 (N_14981,N_14193,N_14097);
or U14982 (N_14982,N_14076,N_14138);
and U14983 (N_14983,N_14419,N_14034);
nand U14984 (N_14984,N_14237,N_14192);
or U14985 (N_14985,N_14327,N_14455);
nand U14986 (N_14986,N_14440,N_14083);
or U14987 (N_14987,N_14182,N_14411);
and U14988 (N_14988,N_14252,N_14393);
xnor U14989 (N_14989,N_14268,N_14091);
or U14990 (N_14990,N_14357,N_14208);
nand U14991 (N_14991,N_14159,N_14306);
nand U14992 (N_14992,N_14404,N_14328);
or U14993 (N_14993,N_14498,N_14148);
and U14994 (N_14994,N_14475,N_14406);
and U14995 (N_14995,N_14278,N_14109);
and U14996 (N_14996,N_14466,N_14457);
xnor U14997 (N_14997,N_14316,N_14038);
nor U14998 (N_14998,N_14490,N_14145);
nand U14999 (N_14999,N_14470,N_14294);
nand U15000 (N_15000,N_14835,N_14985);
or U15001 (N_15001,N_14947,N_14945);
nand U15002 (N_15002,N_14654,N_14899);
xor U15003 (N_15003,N_14935,N_14674);
or U15004 (N_15004,N_14570,N_14611);
xnor U15005 (N_15005,N_14821,N_14605);
and U15006 (N_15006,N_14824,N_14582);
or U15007 (N_15007,N_14556,N_14744);
or U15008 (N_15008,N_14549,N_14711);
xnor U15009 (N_15009,N_14586,N_14970);
nand U15010 (N_15010,N_14538,N_14953);
and U15011 (N_15011,N_14708,N_14598);
xor U15012 (N_15012,N_14734,N_14660);
xor U15013 (N_15013,N_14907,N_14606);
nor U15014 (N_15014,N_14775,N_14941);
xnor U15015 (N_15015,N_14689,N_14546);
or U15016 (N_15016,N_14933,N_14998);
nand U15017 (N_15017,N_14676,N_14569);
xnor U15018 (N_15018,N_14680,N_14709);
nand U15019 (N_15019,N_14866,N_14509);
and U15020 (N_15020,N_14838,N_14865);
nor U15021 (N_15021,N_14579,N_14560);
and U15022 (N_15022,N_14514,N_14594);
and U15023 (N_15023,N_14664,N_14741);
and U15024 (N_15024,N_14743,N_14553);
nor U15025 (N_15025,N_14784,N_14858);
nand U15026 (N_15026,N_14703,N_14531);
nor U15027 (N_15027,N_14652,N_14980);
nand U15028 (N_15028,N_14891,N_14547);
or U15029 (N_15029,N_14515,N_14615);
and U15030 (N_15030,N_14507,N_14673);
or U15031 (N_15031,N_14565,N_14942);
or U15032 (N_15032,N_14996,N_14796);
xor U15033 (N_15033,N_14620,N_14874);
nand U15034 (N_15034,N_14792,N_14966);
nand U15035 (N_15035,N_14690,N_14931);
xnor U15036 (N_15036,N_14927,N_14596);
nor U15037 (N_15037,N_14505,N_14618);
and U15038 (N_15038,N_14897,N_14829);
xor U15039 (N_15039,N_14712,N_14639);
xnor U15040 (N_15040,N_14552,N_14526);
nor U15041 (N_15041,N_14626,N_14906);
or U15042 (N_15042,N_14677,N_14994);
or U15043 (N_15043,N_14642,N_14767);
and U15044 (N_15044,N_14661,N_14789);
and U15045 (N_15045,N_14679,N_14869);
nor U15046 (N_15046,N_14956,N_14727);
nand U15047 (N_15047,N_14644,N_14561);
or U15048 (N_15048,N_14978,N_14532);
or U15049 (N_15049,N_14613,N_14862);
nor U15050 (N_15050,N_14848,N_14732);
nor U15051 (N_15051,N_14663,N_14969);
xnor U15052 (N_15052,N_14748,N_14668);
nor U15053 (N_15053,N_14993,N_14809);
and U15054 (N_15054,N_14923,N_14894);
or U15055 (N_15055,N_14577,N_14905);
nand U15056 (N_15056,N_14908,N_14593);
or U15057 (N_15057,N_14916,N_14873);
or U15058 (N_15058,N_14995,N_14856);
or U15059 (N_15059,N_14887,N_14769);
or U15060 (N_15060,N_14782,N_14982);
nand U15061 (N_15061,N_14754,N_14802);
nor U15062 (N_15062,N_14601,N_14511);
xor U15063 (N_15063,N_14752,N_14818);
or U15064 (N_15064,N_14742,N_14563);
nand U15065 (N_15065,N_14839,N_14772);
nand U15066 (N_15066,N_14859,N_14881);
xnor U15067 (N_15067,N_14675,N_14877);
nand U15068 (N_15068,N_14999,N_14946);
xnor U15069 (N_15069,N_14595,N_14659);
xor U15070 (N_15070,N_14909,N_14760);
nor U15071 (N_15071,N_14501,N_14517);
nand U15072 (N_15072,N_14631,N_14692);
nand U15073 (N_15073,N_14527,N_14901);
or U15074 (N_15074,N_14610,N_14841);
and U15075 (N_15075,N_14851,N_14831);
nand U15076 (N_15076,N_14603,N_14648);
nor U15077 (N_15077,N_14846,N_14948);
and U15078 (N_15078,N_14700,N_14814);
nand U15079 (N_15079,N_14799,N_14600);
or U15080 (N_15080,N_14997,N_14807);
xor U15081 (N_15081,N_14888,N_14518);
or U15082 (N_15082,N_14584,N_14612);
and U15083 (N_15083,N_14926,N_14559);
xor U15084 (N_15084,N_14896,N_14885);
nand U15085 (N_15085,N_14840,N_14961);
xnor U15086 (N_15086,N_14629,N_14646);
and U15087 (N_15087,N_14950,N_14981);
or U15088 (N_15088,N_14804,N_14836);
nor U15089 (N_15089,N_14794,N_14702);
nor U15090 (N_15090,N_14850,N_14681);
nand U15091 (N_15091,N_14832,N_14695);
and U15092 (N_15092,N_14903,N_14588);
or U15093 (N_15093,N_14863,N_14637);
or U15094 (N_15094,N_14710,N_14638);
xnor U15095 (N_15095,N_14714,N_14774);
nor U15096 (N_15096,N_14658,N_14979);
nor U15097 (N_15097,N_14973,N_14820);
nand U15098 (N_15098,N_14576,N_14653);
and U15099 (N_15099,N_14834,N_14954);
nor U15100 (N_15100,N_14550,N_14694);
xnor U15101 (N_15101,N_14825,N_14949);
nand U15102 (N_15102,N_14587,N_14591);
xor U15103 (N_15103,N_14977,N_14808);
xnor U15104 (N_15104,N_14705,N_14911);
and U15105 (N_15105,N_14771,N_14793);
and U15106 (N_15106,N_14707,N_14750);
and U15107 (N_15107,N_14649,N_14542);
nor U15108 (N_15108,N_14880,N_14790);
or U15109 (N_15109,N_14893,N_14928);
nand U15110 (N_15110,N_14967,N_14720);
and U15111 (N_15111,N_14619,N_14854);
nand U15112 (N_15112,N_14934,N_14568);
and U15113 (N_15113,N_14762,N_14861);
nand U15114 (N_15114,N_14987,N_14730);
or U15115 (N_15115,N_14573,N_14766);
nor U15116 (N_15116,N_14847,N_14915);
xnor U15117 (N_15117,N_14806,N_14965);
or U15118 (N_15118,N_14686,N_14844);
xnor U15119 (N_15119,N_14544,N_14882);
nand U15120 (N_15120,N_14910,N_14914);
xnor U15121 (N_15121,N_14955,N_14578);
nor U15122 (N_15122,N_14738,N_14656);
nor U15123 (N_15123,N_14698,N_14651);
nand U15124 (N_15124,N_14722,N_14951);
xnor U15125 (N_15125,N_14974,N_14622);
or U15126 (N_15126,N_14780,N_14512);
and U15127 (N_15127,N_14528,N_14585);
or U15128 (N_15128,N_14545,N_14759);
nor U15129 (N_15129,N_14886,N_14878);
nand U15130 (N_15130,N_14548,N_14571);
nor U15131 (N_15131,N_14616,N_14657);
and U15132 (N_15132,N_14739,N_14699);
and U15133 (N_15133,N_14683,N_14687);
or U15134 (N_15134,N_14904,N_14813);
xnor U15135 (N_15135,N_14716,N_14621);
nand U15136 (N_15136,N_14617,N_14643);
nand U15137 (N_15137,N_14819,N_14747);
xor U15138 (N_15138,N_14715,N_14597);
and U15139 (N_15139,N_14922,N_14917);
nor U15140 (N_15140,N_14581,N_14721);
and U15141 (N_15141,N_14826,N_14930);
or U15142 (N_15142,N_14785,N_14816);
and U15143 (N_15143,N_14608,N_14736);
or U15144 (N_15144,N_14855,N_14539);
nand U15145 (N_15145,N_14671,N_14876);
nor U15146 (N_15146,N_14920,N_14731);
or U15147 (N_15147,N_14756,N_14860);
nand U15148 (N_15148,N_14519,N_14520);
xor U15149 (N_15149,N_14589,N_14890);
and U15150 (N_15150,N_14669,N_14609);
nand U15151 (N_15151,N_14823,N_14892);
or U15152 (N_15152,N_14830,N_14575);
or U15153 (N_15153,N_14857,N_14845);
or U15154 (N_15154,N_14939,N_14728);
and U15155 (N_15155,N_14729,N_14919);
xnor U15156 (N_15156,N_14691,N_14773);
nand U15157 (N_15157,N_14937,N_14765);
nand U15158 (N_15158,N_14770,N_14758);
nor U15159 (N_15159,N_14696,N_14628);
nand U15160 (N_15160,N_14898,N_14952);
xnor U15161 (N_15161,N_14627,N_14795);
or U15162 (N_15162,N_14636,N_14929);
nor U15163 (N_15163,N_14875,N_14884);
nor U15164 (N_15164,N_14853,N_14801);
nand U15165 (N_15165,N_14530,N_14522);
nor U15166 (N_15166,N_14555,N_14537);
and U15167 (N_15167,N_14564,N_14986);
nand U15168 (N_15168,N_14684,N_14755);
and U15169 (N_15169,N_14924,N_14533);
and U15170 (N_15170,N_14912,N_14957);
xnor U15171 (N_15171,N_14602,N_14701);
xnor U15172 (N_15172,N_14670,N_14843);
nand U15173 (N_15173,N_14726,N_14828);
nor U15174 (N_15174,N_14574,N_14724);
and U15175 (N_15175,N_14833,N_14786);
nand U15176 (N_15176,N_14879,N_14554);
nor U15177 (N_15177,N_14719,N_14817);
nand U15178 (N_15178,N_14717,N_14870);
nand U15179 (N_15179,N_14815,N_14913);
nand U15180 (N_15180,N_14972,N_14940);
or U15181 (N_15181,N_14614,N_14751);
xor U15182 (N_15182,N_14811,N_14842);
or U15183 (N_15183,N_14635,N_14718);
or U15184 (N_15184,N_14849,N_14976);
xnor U15185 (N_15185,N_14810,N_14740);
nand U15186 (N_15186,N_14990,N_14529);
nor U15187 (N_15187,N_14523,N_14962);
xnor U15188 (N_15188,N_14685,N_14513);
xnor U15189 (N_15189,N_14641,N_14746);
nand U15190 (N_15190,N_14540,N_14607);
nand U15191 (N_15191,N_14918,N_14557);
nor U15192 (N_15192,N_14634,N_14500);
or U15193 (N_15193,N_14989,N_14778);
nand U15194 (N_15194,N_14704,N_14852);
nand U15195 (N_15195,N_14788,N_14590);
nor U15196 (N_15196,N_14943,N_14524);
or U15197 (N_15197,N_14580,N_14936);
xor U15198 (N_15198,N_14535,N_14889);
xor U15199 (N_15199,N_14650,N_14991);
nand U15200 (N_15200,N_14733,N_14666);
nor U15201 (N_15201,N_14693,N_14800);
xor U15202 (N_15202,N_14983,N_14803);
nor U15203 (N_15203,N_14723,N_14959);
or U15204 (N_15204,N_14583,N_14791);
nor U15205 (N_15205,N_14902,N_14988);
nor U15206 (N_15206,N_14763,N_14900);
and U15207 (N_15207,N_14682,N_14779);
or U15208 (N_15208,N_14932,N_14783);
xor U15209 (N_15209,N_14633,N_14777);
xor U15210 (N_15210,N_14764,N_14944);
nand U15211 (N_15211,N_14787,N_14655);
nand U15212 (N_15212,N_14812,N_14567);
xor U15213 (N_15213,N_14632,N_14776);
nor U15214 (N_15214,N_14623,N_14975);
xor U15215 (N_15215,N_14757,N_14798);
and U15216 (N_15216,N_14968,N_14566);
nand U15217 (N_15217,N_14665,N_14960);
and U15218 (N_15218,N_14883,N_14630);
nand U15219 (N_15219,N_14895,N_14536);
nand U15220 (N_15220,N_14735,N_14805);
or U15221 (N_15221,N_14510,N_14558);
or U15222 (N_15222,N_14713,N_14504);
nand U15223 (N_15223,N_14871,N_14506);
nand U15224 (N_15224,N_14958,N_14781);
nor U15225 (N_15225,N_14592,N_14761);
xnor U15226 (N_15226,N_14737,N_14543);
xor U15227 (N_15227,N_14521,N_14541);
and U15228 (N_15228,N_14645,N_14867);
nor U15229 (N_15229,N_14562,N_14672);
and U15230 (N_15230,N_14647,N_14525);
xor U15231 (N_15231,N_14502,N_14662);
and U15232 (N_15232,N_14534,N_14837);
nand U15233 (N_15233,N_14984,N_14868);
or U15234 (N_15234,N_14678,N_14688);
and U15235 (N_15235,N_14697,N_14963);
xnor U15236 (N_15236,N_14864,N_14640);
and U15237 (N_15237,N_14625,N_14624);
nor U15238 (N_15238,N_14964,N_14971);
and U15239 (N_15239,N_14516,N_14753);
or U15240 (N_15240,N_14921,N_14508);
nor U15241 (N_15241,N_14551,N_14745);
or U15242 (N_15242,N_14768,N_14822);
nor U15243 (N_15243,N_14749,N_14872);
and U15244 (N_15244,N_14992,N_14604);
and U15245 (N_15245,N_14827,N_14503);
and U15246 (N_15246,N_14938,N_14667);
nor U15247 (N_15247,N_14706,N_14599);
nand U15248 (N_15248,N_14572,N_14725);
or U15249 (N_15249,N_14797,N_14925);
xnor U15250 (N_15250,N_14664,N_14514);
nor U15251 (N_15251,N_14914,N_14768);
or U15252 (N_15252,N_14839,N_14704);
and U15253 (N_15253,N_14958,N_14551);
and U15254 (N_15254,N_14624,N_14854);
or U15255 (N_15255,N_14598,N_14837);
nand U15256 (N_15256,N_14798,N_14639);
or U15257 (N_15257,N_14829,N_14758);
xor U15258 (N_15258,N_14508,N_14775);
nor U15259 (N_15259,N_14747,N_14545);
or U15260 (N_15260,N_14679,N_14661);
xnor U15261 (N_15261,N_14846,N_14735);
or U15262 (N_15262,N_14909,N_14775);
and U15263 (N_15263,N_14825,N_14974);
and U15264 (N_15264,N_14871,N_14883);
or U15265 (N_15265,N_14975,N_14693);
or U15266 (N_15266,N_14565,N_14844);
or U15267 (N_15267,N_14646,N_14553);
or U15268 (N_15268,N_14949,N_14822);
nand U15269 (N_15269,N_14737,N_14678);
or U15270 (N_15270,N_14616,N_14634);
nand U15271 (N_15271,N_14714,N_14988);
nor U15272 (N_15272,N_14616,N_14886);
nor U15273 (N_15273,N_14599,N_14511);
or U15274 (N_15274,N_14831,N_14873);
nor U15275 (N_15275,N_14674,N_14538);
nand U15276 (N_15276,N_14726,N_14519);
and U15277 (N_15277,N_14521,N_14966);
or U15278 (N_15278,N_14623,N_14931);
nand U15279 (N_15279,N_14569,N_14576);
or U15280 (N_15280,N_14890,N_14637);
xor U15281 (N_15281,N_14971,N_14691);
nor U15282 (N_15282,N_14563,N_14575);
xnor U15283 (N_15283,N_14725,N_14965);
nor U15284 (N_15284,N_14720,N_14728);
xnor U15285 (N_15285,N_14664,N_14904);
and U15286 (N_15286,N_14676,N_14657);
and U15287 (N_15287,N_14756,N_14733);
and U15288 (N_15288,N_14705,N_14631);
nor U15289 (N_15289,N_14695,N_14778);
xnor U15290 (N_15290,N_14996,N_14665);
xor U15291 (N_15291,N_14560,N_14929);
and U15292 (N_15292,N_14685,N_14520);
nor U15293 (N_15293,N_14870,N_14871);
xor U15294 (N_15294,N_14610,N_14667);
nor U15295 (N_15295,N_14966,N_14880);
nor U15296 (N_15296,N_14975,N_14534);
or U15297 (N_15297,N_14978,N_14671);
nor U15298 (N_15298,N_14742,N_14646);
nor U15299 (N_15299,N_14822,N_14568);
and U15300 (N_15300,N_14554,N_14938);
or U15301 (N_15301,N_14650,N_14553);
nand U15302 (N_15302,N_14724,N_14923);
xnor U15303 (N_15303,N_14581,N_14812);
nor U15304 (N_15304,N_14895,N_14778);
and U15305 (N_15305,N_14787,N_14843);
xnor U15306 (N_15306,N_14648,N_14730);
and U15307 (N_15307,N_14513,N_14929);
xnor U15308 (N_15308,N_14651,N_14714);
or U15309 (N_15309,N_14528,N_14955);
nand U15310 (N_15310,N_14999,N_14526);
nand U15311 (N_15311,N_14961,N_14560);
and U15312 (N_15312,N_14725,N_14656);
or U15313 (N_15313,N_14644,N_14773);
or U15314 (N_15314,N_14740,N_14998);
nand U15315 (N_15315,N_14931,N_14701);
and U15316 (N_15316,N_14900,N_14503);
xor U15317 (N_15317,N_14618,N_14917);
nand U15318 (N_15318,N_14943,N_14675);
or U15319 (N_15319,N_14801,N_14876);
or U15320 (N_15320,N_14941,N_14591);
and U15321 (N_15321,N_14926,N_14742);
xnor U15322 (N_15322,N_14528,N_14882);
nand U15323 (N_15323,N_14584,N_14720);
nand U15324 (N_15324,N_14507,N_14818);
nand U15325 (N_15325,N_14662,N_14691);
nor U15326 (N_15326,N_14668,N_14926);
xor U15327 (N_15327,N_14905,N_14507);
and U15328 (N_15328,N_14992,N_14629);
nand U15329 (N_15329,N_14813,N_14639);
xor U15330 (N_15330,N_14665,N_14778);
xnor U15331 (N_15331,N_14658,N_14780);
xor U15332 (N_15332,N_14933,N_14838);
xor U15333 (N_15333,N_14934,N_14872);
and U15334 (N_15334,N_14916,N_14580);
and U15335 (N_15335,N_14651,N_14835);
xor U15336 (N_15336,N_14908,N_14632);
xnor U15337 (N_15337,N_14884,N_14559);
and U15338 (N_15338,N_14696,N_14557);
xnor U15339 (N_15339,N_14876,N_14782);
nor U15340 (N_15340,N_14536,N_14963);
and U15341 (N_15341,N_14791,N_14595);
and U15342 (N_15342,N_14586,N_14557);
or U15343 (N_15343,N_14875,N_14824);
or U15344 (N_15344,N_14813,N_14998);
nand U15345 (N_15345,N_14710,N_14865);
or U15346 (N_15346,N_14608,N_14794);
nor U15347 (N_15347,N_14843,N_14701);
or U15348 (N_15348,N_14650,N_14823);
and U15349 (N_15349,N_14742,N_14732);
xnor U15350 (N_15350,N_14992,N_14755);
nand U15351 (N_15351,N_14634,N_14908);
nand U15352 (N_15352,N_14790,N_14973);
and U15353 (N_15353,N_14934,N_14500);
nand U15354 (N_15354,N_14781,N_14945);
nor U15355 (N_15355,N_14556,N_14677);
nand U15356 (N_15356,N_14735,N_14982);
xnor U15357 (N_15357,N_14814,N_14764);
nor U15358 (N_15358,N_14802,N_14720);
xnor U15359 (N_15359,N_14837,N_14706);
and U15360 (N_15360,N_14896,N_14611);
and U15361 (N_15361,N_14580,N_14538);
nor U15362 (N_15362,N_14502,N_14839);
xnor U15363 (N_15363,N_14646,N_14675);
nor U15364 (N_15364,N_14764,N_14758);
xor U15365 (N_15365,N_14957,N_14625);
nor U15366 (N_15366,N_14537,N_14744);
xor U15367 (N_15367,N_14570,N_14721);
and U15368 (N_15368,N_14515,N_14673);
nand U15369 (N_15369,N_14606,N_14827);
xor U15370 (N_15370,N_14641,N_14721);
and U15371 (N_15371,N_14753,N_14814);
xor U15372 (N_15372,N_14687,N_14745);
or U15373 (N_15373,N_14534,N_14971);
and U15374 (N_15374,N_14525,N_14970);
xnor U15375 (N_15375,N_14820,N_14898);
nand U15376 (N_15376,N_14775,N_14668);
or U15377 (N_15377,N_14983,N_14634);
nand U15378 (N_15378,N_14729,N_14979);
or U15379 (N_15379,N_14870,N_14546);
and U15380 (N_15380,N_14548,N_14588);
xor U15381 (N_15381,N_14894,N_14654);
xnor U15382 (N_15382,N_14707,N_14962);
and U15383 (N_15383,N_14850,N_14637);
or U15384 (N_15384,N_14979,N_14815);
nor U15385 (N_15385,N_14920,N_14916);
and U15386 (N_15386,N_14610,N_14860);
and U15387 (N_15387,N_14539,N_14994);
or U15388 (N_15388,N_14513,N_14519);
nor U15389 (N_15389,N_14514,N_14737);
xor U15390 (N_15390,N_14902,N_14756);
nor U15391 (N_15391,N_14843,N_14986);
or U15392 (N_15392,N_14657,N_14690);
xnor U15393 (N_15393,N_14942,N_14761);
xor U15394 (N_15394,N_14539,N_14826);
xor U15395 (N_15395,N_14883,N_14672);
nor U15396 (N_15396,N_14809,N_14797);
and U15397 (N_15397,N_14602,N_14575);
and U15398 (N_15398,N_14830,N_14711);
nor U15399 (N_15399,N_14649,N_14587);
nor U15400 (N_15400,N_14571,N_14635);
nand U15401 (N_15401,N_14540,N_14797);
and U15402 (N_15402,N_14621,N_14749);
xnor U15403 (N_15403,N_14538,N_14966);
and U15404 (N_15404,N_14721,N_14784);
and U15405 (N_15405,N_14921,N_14630);
xor U15406 (N_15406,N_14857,N_14538);
nand U15407 (N_15407,N_14686,N_14635);
xor U15408 (N_15408,N_14854,N_14799);
nor U15409 (N_15409,N_14922,N_14758);
and U15410 (N_15410,N_14535,N_14684);
nor U15411 (N_15411,N_14896,N_14761);
or U15412 (N_15412,N_14906,N_14597);
xor U15413 (N_15413,N_14573,N_14631);
xnor U15414 (N_15414,N_14767,N_14883);
nor U15415 (N_15415,N_14504,N_14634);
xor U15416 (N_15416,N_14876,N_14999);
xor U15417 (N_15417,N_14843,N_14894);
nor U15418 (N_15418,N_14649,N_14977);
and U15419 (N_15419,N_14995,N_14970);
and U15420 (N_15420,N_14599,N_14568);
nor U15421 (N_15421,N_14667,N_14734);
xnor U15422 (N_15422,N_14824,N_14645);
nor U15423 (N_15423,N_14589,N_14984);
xor U15424 (N_15424,N_14614,N_14798);
xor U15425 (N_15425,N_14805,N_14864);
xnor U15426 (N_15426,N_14813,N_14876);
nor U15427 (N_15427,N_14777,N_14510);
nand U15428 (N_15428,N_14636,N_14747);
xor U15429 (N_15429,N_14698,N_14600);
nor U15430 (N_15430,N_14573,N_14575);
and U15431 (N_15431,N_14968,N_14908);
nand U15432 (N_15432,N_14791,N_14809);
or U15433 (N_15433,N_14537,N_14530);
and U15434 (N_15434,N_14854,N_14977);
nand U15435 (N_15435,N_14558,N_14826);
nor U15436 (N_15436,N_14683,N_14601);
xnor U15437 (N_15437,N_14742,N_14982);
nand U15438 (N_15438,N_14916,N_14877);
and U15439 (N_15439,N_14796,N_14573);
nor U15440 (N_15440,N_14775,N_14845);
or U15441 (N_15441,N_14987,N_14517);
or U15442 (N_15442,N_14803,N_14839);
nor U15443 (N_15443,N_14870,N_14701);
xnor U15444 (N_15444,N_14717,N_14957);
nor U15445 (N_15445,N_14893,N_14649);
and U15446 (N_15446,N_14712,N_14810);
and U15447 (N_15447,N_14679,N_14729);
and U15448 (N_15448,N_14969,N_14649);
nand U15449 (N_15449,N_14838,N_14937);
nand U15450 (N_15450,N_14872,N_14823);
nand U15451 (N_15451,N_14523,N_14702);
and U15452 (N_15452,N_14704,N_14597);
and U15453 (N_15453,N_14749,N_14842);
nand U15454 (N_15454,N_14879,N_14740);
xnor U15455 (N_15455,N_14750,N_14634);
xnor U15456 (N_15456,N_14894,N_14817);
xor U15457 (N_15457,N_14528,N_14599);
or U15458 (N_15458,N_14658,N_14903);
nor U15459 (N_15459,N_14584,N_14907);
nand U15460 (N_15460,N_14920,N_14553);
or U15461 (N_15461,N_14517,N_14938);
and U15462 (N_15462,N_14738,N_14709);
xnor U15463 (N_15463,N_14631,N_14934);
or U15464 (N_15464,N_14742,N_14572);
nor U15465 (N_15465,N_14723,N_14508);
nor U15466 (N_15466,N_14777,N_14685);
nor U15467 (N_15467,N_14983,N_14615);
xnor U15468 (N_15468,N_14758,N_14783);
xor U15469 (N_15469,N_14755,N_14930);
and U15470 (N_15470,N_14975,N_14523);
nand U15471 (N_15471,N_14901,N_14757);
and U15472 (N_15472,N_14749,N_14526);
nor U15473 (N_15473,N_14591,N_14829);
xnor U15474 (N_15474,N_14511,N_14593);
or U15475 (N_15475,N_14596,N_14840);
xor U15476 (N_15476,N_14612,N_14508);
nand U15477 (N_15477,N_14715,N_14726);
and U15478 (N_15478,N_14953,N_14710);
nor U15479 (N_15479,N_14736,N_14745);
or U15480 (N_15480,N_14790,N_14799);
and U15481 (N_15481,N_14872,N_14516);
nand U15482 (N_15482,N_14852,N_14844);
xnor U15483 (N_15483,N_14837,N_14810);
nand U15484 (N_15484,N_14572,N_14884);
nand U15485 (N_15485,N_14763,N_14958);
nor U15486 (N_15486,N_14908,N_14913);
and U15487 (N_15487,N_14700,N_14547);
nand U15488 (N_15488,N_14554,N_14872);
nand U15489 (N_15489,N_14520,N_14575);
nand U15490 (N_15490,N_14670,N_14651);
xor U15491 (N_15491,N_14785,N_14914);
xnor U15492 (N_15492,N_14705,N_14903);
or U15493 (N_15493,N_14966,N_14535);
nor U15494 (N_15494,N_14773,N_14885);
and U15495 (N_15495,N_14998,N_14738);
nor U15496 (N_15496,N_14828,N_14723);
and U15497 (N_15497,N_14797,N_14565);
or U15498 (N_15498,N_14800,N_14849);
or U15499 (N_15499,N_14817,N_14613);
nand U15500 (N_15500,N_15127,N_15188);
or U15501 (N_15501,N_15007,N_15051);
or U15502 (N_15502,N_15053,N_15244);
nor U15503 (N_15503,N_15418,N_15406);
nand U15504 (N_15504,N_15357,N_15466);
or U15505 (N_15505,N_15265,N_15093);
nor U15506 (N_15506,N_15035,N_15427);
and U15507 (N_15507,N_15399,N_15270);
nor U15508 (N_15508,N_15046,N_15088);
nor U15509 (N_15509,N_15227,N_15212);
or U15510 (N_15510,N_15442,N_15283);
nand U15511 (N_15511,N_15237,N_15006);
xor U15512 (N_15512,N_15463,N_15459);
xnor U15513 (N_15513,N_15339,N_15488);
or U15514 (N_15514,N_15172,N_15091);
xor U15515 (N_15515,N_15003,N_15061);
or U15516 (N_15516,N_15347,N_15178);
or U15517 (N_15517,N_15079,N_15487);
or U15518 (N_15518,N_15390,N_15369);
and U15519 (N_15519,N_15101,N_15142);
xnor U15520 (N_15520,N_15461,N_15361);
and U15521 (N_15521,N_15438,N_15349);
nor U15522 (N_15522,N_15489,N_15001);
xnor U15523 (N_15523,N_15010,N_15113);
xnor U15524 (N_15524,N_15310,N_15037);
nand U15525 (N_15525,N_15315,N_15126);
or U15526 (N_15526,N_15253,N_15081);
or U15527 (N_15527,N_15462,N_15191);
xnor U15528 (N_15528,N_15471,N_15258);
or U15529 (N_15529,N_15481,N_15193);
nor U15530 (N_15530,N_15054,N_15065);
nor U15531 (N_15531,N_15385,N_15116);
or U15532 (N_15532,N_15002,N_15450);
or U15533 (N_15533,N_15386,N_15082);
or U15534 (N_15534,N_15411,N_15419);
or U15535 (N_15535,N_15200,N_15394);
or U15536 (N_15536,N_15202,N_15161);
or U15537 (N_15537,N_15375,N_15423);
and U15538 (N_15538,N_15073,N_15320);
nand U15539 (N_15539,N_15210,N_15284);
nor U15540 (N_15540,N_15495,N_15132);
and U15541 (N_15541,N_15206,N_15058);
or U15542 (N_15542,N_15312,N_15222);
nor U15543 (N_15543,N_15134,N_15441);
nor U15544 (N_15544,N_15345,N_15299);
nor U15545 (N_15545,N_15092,N_15179);
nand U15546 (N_15546,N_15074,N_15140);
nand U15547 (N_15547,N_15122,N_15041);
or U15548 (N_15548,N_15297,N_15359);
xnor U15549 (N_15549,N_15292,N_15175);
nor U15550 (N_15550,N_15255,N_15384);
nor U15551 (N_15551,N_15008,N_15391);
and U15552 (N_15552,N_15393,N_15430);
and U15553 (N_15553,N_15224,N_15447);
xor U15554 (N_15554,N_15023,N_15036);
nor U15555 (N_15555,N_15440,N_15346);
nor U15556 (N_15556,N_15165,N_15186);
and U15557 (N_15557,N_15236,N_15263);
xor U15558 (N_15558,N_15448,N_15434);
nor U15559 (N_15559,N_15313,N_15412);
or U15560 (N_15560,N_15445,N_15314);
or U15561 (N_15561,N_15039,N_15205);
nor U15562 (N_15562,N_15392,N_15473);
or U15563 (N_15563,N_15018,N_15323);
nand U15564 (N_15564,N_15107,N_15135);
nand U15565 (N_15565,N_15217,N_15425);
xor U15566 (N_15566,N_15366,N_15112);
xor U15567 (N_15567,N_15497,N_15278);
xor U15568 (N_15568,N_15408,N_15052);
xor U15569 (N_15569,N_15211,N_15398);
nand U15570 (N_15570,N_15443,N_15176);
nand U15571 (N_15571,N_15477,N_15060);
xnor U15572 (N_15572,N_15275,N_15376);
nor U15573 (N_15573,N_15141,N_15121);
nor U15574 (N_15574,N_15492,N_15195);
nor U15575 (N_15575,N_15012,N_15029);
nor U15576 (N_15576,N_15261,N_15137);
or U15577 (N_15577,N_15120,N_15262);
xnor U15578 (N_15578,N_15031,N_15334);
nand U15579 (N_15579,N_15213,N_15301);
xor U15580 (N_15580,N_15154,N_15281);
and U15581 (N_15581,N_15019,N_15469);
and U15582 (N_15582,N_15364,N_15279);
xor U15583 (N_15583,N_15353,N_15449);
nand U15584 (N_15584,N_15421,N_15389);
or U15585 (N_15585,N_15221,N_15118);
or U15586 (N_15586,N_15420,N_15063);
nand U15587 (N_15587,N_15096,N_15405);
nand U15588 (N_15588,N_15152,N_15038);
and U15589 (N_15589,N_15341,N_15280);
nand U15590 (N_15590,N_15336,N_15470);
nand U15591 (N_15591,N_15250,N_15454);
nand U15592 (N_15592,N_15057,N_15407);
and U15593 (N_15593,N_15242,N_15467);
nand U15594 (N_15594,N_15291,N_15247);
and U15595 (N_15595,N_15215,N_15371);
nor U15596 (N_15596,N_15174,N_15214);
xnor U15597 (N_15597,N_15017,N_15468);
or U15598 (N_15598,N_15269,N_15256);
xnor U15599 (N_15599,N_15155,N_15180);
xnor U15600 (N_15600,N_15072,N_15095);
or U15601 (N_15601,N_15271,N_15327);
nor U15602 (N_15602,N_15431,N_15160);
or U15603 (N_15603,N_15226,N_15304);
xnor U15604 (N_15604,N_15167,N_15335);
nand U15605 (N_15605,N_15138,N_15196);
and U15606 (N_15606,N_15111,N_15311);
xnor U15607 (N_15607,N_15429,N_15254);
and U15608 (N_15608,N_15047,N_15109);
and U15609 (N_15609,N_15128,N_15344);
nand U15610 (N_15610,N_15373,N_15043);
xnor U15611 (N_15611,N_15050,N_15189);
nand U15612 (N_15612,N_15040,N_15192);
nand U15613 (N_15613,N_15474,N_15444);
nand U15614 (N_15614,N_15048,N_15169);
xnor U15615 (N_15615,N_15294,N_15499);
nor U15616 (N_15616,N_15356,N_15231);
and U15617 (N_15617,N_15337,N_15240);
nand U15618 (N_15618,N_15124,N_15319);
nor U15619 (N_15619,N_15485,N_15087);
xor U15620 (N_15620,N_15415,N_15322);
xor U15621 (N_15621,N_15317,N_15168);
nand U15622 (N_15622,N_15378,N_15402);
xor U15623 (N_15623,N_15171,N_15309);
nor U15624 (N_15624,N_15153,N_15325);
and U15625 (N_15625,N_15077,N_15354);
or U15626 (N_15626,N_15277,N_15187);
nor U15627 (N_15627,N_15055,N_15351);
nor U15628 (N_15628,N_15290,N_15476);
nor U15629 (N_15629,N_15451,N_15252);
or U15630 (N_15630,N_15316,N_15099);
nand U15631 (N_15631,N_15208,N_15021);
nand U15632 (N_15632,N_15108,N_15318);
and U15633 (N_15633,N_15422,N_15225);
nor U15634 (N_15634,N_15194,N_15251);
and U15635 (N_15635,N_15076,N_15044);
or U15636 (N_15636,N_15433,N_15005);
and U15637 (N_15637,N_15228,N_15472);
nor U15638 (N_15638,N_15401,N_15381);
or U15639 (N_15639,N_15395,N_15158);
xnor U15640 (N_15640,N_15143,N_15117);
and U15641 (N_15641,N_15136,N_15151);
nand U15642 (N_15642,N_15230,N_15400);
and U15643 (N_15643,N_15370,N_15287);
xnor U15644 (N_15644,N_15177,N_15289);
and U15645 (N_15645,N_15148,N_15484);
and U15646 (N_15646,N_15350,N_15182);
nor U15647 (N_15647,N_15083,N_15159);
nand U15648 (N_15648,N_15146,N_15098);
nand U15649 (N_15649,N_15348,N_15062);
or U15650 (N_15650,N_15028,N_15331);
or U15651 (N_15651,N_15343,N_15330);
and U15652 (N_15652,N_15358,N_15372);
and U15653 (N_15653,N_15004,N_15374);
nor U15654 (N_15654,N_15000,N_15272);
and U15655 (N_15655,N_15446,N_15110);
nand U15656 (N_15656,N_15413,N_15479);
or U15657 (N_15657,N_15388,N_15102);
and U15658 (N_15658,N_15465,N_15363);
nor U15659 (N_15659,N_15305,N_15367);
xor U15660 (N_15660,N_15298,N_15241);
nand U15661 (N_15661,N_15145,N_15303);
and U15662 (N_15662,N_15166,N_15295);
and U15663 (N_15663,N_15268,N_15204);
nand U15664 (N_15664,N_15486,N_15494);
or U15665 (N_15665,N_15382,N_15483);
xor U15666 (N_15666,N_15094,N_15173);
or U15667 (N_15667,N_15078,N_15266);
nor U15668 (N_15668,N_15246,N_15377);
xor U15669 (N_15669,N_15199,N_15306);
and U15670 (N_15670,N_15034,N_15426);
nand U15671 (N_15671,N_15307,N_15439);
and U15672 (N_15672,N_15286,N_15020);
nand U15673 (N_15673,N_15260,N_15219);
nor U15674 (N_15674,N_15308,N_15387);
nor U15675 (N_15675,N_15328,N_15380);
nor U15676 (N_15676,N_15480,N_15243);
xor U15677 (N_15677,N_15342,N_15106);
and U15678 (N_15678,N_15059,N_15404);
nor U15679 (N_15679,N_15379,N_15285);
nor U15680 (N_15680,N_15115,N_15482);
or U15681 (N_15681,N_15080,N_15070);
nor U15682 (N_15682,N_15455,N_15209);
nor U15683 (N_15683,N_15332,N_15201);
nor U15684 (N_15684,N_15119,N_15066);
and U15685 (N_15685,N_15259,N_15162);
xnor U15686 (N_15686,N_15144,N_15452);
or U15687 (N_15687,N_15282,N_15264);
xnor U15688 (N_15688,N_15475,N_15293);
or U15689 (N_15689,N_15435,N_15056);
xnor U15690 (N_15690,N_15300,N_15410);
nand U15691 (N_15691,N_15185,N_15338);
and U15692 (N_15692,N_15009,N_15245);
and U15693 (N_15693,N_15086,N_15014);
and U15694 (N_15694,N_15249,N_15491);
xor U15695 (N_15695,N_15170,N_15460);
and U15696 (N_15696,N_15015,N_15183);
nand U15697 (N_15697,N_15355,N_15248);
nor U15698 (N_15698,N_15493,N_15011);
nor U15699 (N_15699,N_15016,N_15045);
xnor U15700 (N_15700,N_15218,N_15097);
xnor U15701 (N_15701,N_15233,N_15417);
nand U15702 (N_15702,N_15064,N_15030);
and U15703 (N_15703,N_15383,N_15129);
xnor U15704 (N_15704,N_15184,N_15416);
nor U15705 (N_15705,N_15321,N_15133);
and U15706 (N_15706,N_15302,N_15027);
and U15707 (N_15707,N_15414,N_15288);
or U15708 (N_15708,N_15464,N_15432);
xor U15709 (N_15709,N_15157,N_15163);
and U15710 (N_15710,N_15147,N_15197);
nand U15711 (N_15711,N_15024,N_15090);
nand U15712 (N_15712,N_15409,N_15239);
nand U15713 (N_15713,N_15326,N_15232);
nand U15714 (N_15714,N_15352,N_15273);
and U15715 (N_15715,N_15100,N_15084);
and U15716 (N_15716,N_15105,N_15013);
xor U15717 (N_15717,N_15456,N_15025);
and U15718 (N_15718,N_15032,N_15296);
xor U15719 (N_15719,N_15458,N_15104);
nand U15720 (N_15720,N_15437,N_15125);
and U15721 (N_15721,N_15069,N_15234);
nand U15722 (N_15722,N_15216,N_15340);
nand U15723 (N_15723,N_15049,N_15457);
or U15724 (N_15724,N_15164,N_15220);
nor U15725 (N_15725,N_15257,N_15198);
nor U15726 (N_15726,N_15453,N_15203);
xor U15727 (N_15727,N_15362,N_15139);
and U15728 (N_15728,N_15207,N_15190);
xnor U15729 (N_15729,N_15103,N_15396);
xnor U15730 (N_15730,N_15114,N_15033);
or U15731 (N_15731,N_15365,N_15130);
and U15732 (N_15732,N_15324,N_15068);
nand U15733 (N_15733,N_15267,N_15156);
nand U15734 (N_15734,N_15498,N_15089);
or U15735 (N_15735,N_15424,N_15150);
nand U15736 (N_15736,N_15071,N_15403);
or U15737 (N_15737,N_15131,N_15397);
xor U15738 (N_15738,N_15042,N_15022);
nor U15739 (N_15739,N_15478,N_15026);
and U15740 (N_15740,N_15149,N_15368);
or U15741 (N_15741,N_15496,N_15428);
nand U15742 (N_15742,N_15329,N_15436);
nand U15743 (N_15743,N_15490,N_15229);
xor U15744 (N_15744,N_15223,N_15333);
xnor U15745 (N_15745,N_15276,N_15123);
nor U15746 (N_15746,N_15235,N_15360);
nand U15747 (N_15747,N_15075,N_15274);
nor U15748 (N_15748,N_15085,N_15181);
nand U15749 (N_15749,N_15238,N_15067);
nor U15750 (N_15750,N_15167,N_15416);
or U15751 (N_15751,N_15365,N_15131);
xor U15752 (N_15752,N_15117,N_15471);
and U15753 (N_15753,N_15033,N_15305);
or U15754 (N_15754,N_15100,N_15466);
nand U15755 (N_15755,N_15489,N_15358);
xor U15756 (N_15756,N_15296,N_15018);
xnor U15757 (N_15757,N_15127,N_15305);
xnor U15758 (N_15758,N_15476,N_15367);
xnor U15759 (N_15759,N_15076,N_15027);
xnor U15760 (N_15760,N_15062,N_15030);
nand U15761 (N_15761,N_15172,N_15076);
or U15762 (N_15762,N_15312,N_15480);
nand U15763 (N_15763,N_15345,N_15215);
nor U15764 (N_15764,N_15037,N_15001);
and U15765 (N_15765,N_15160,N_15209);
xnor U15766 (N_15766,N_15148,N_15274);
nand U15767 (N_15767,N_15111,N_15063);
or U15768 (N_15768,N_15299,N_15466);
xnor U15769 (N_15769,N_15039,N_15246);
nand U15770 (N_15770,N_15428,N_15401);
nor U15771 (N_15771,N_15260,N_15114);
and U15772 (N_15772,N_15265,N_15280);
and U15773 (N_15773,N_15403,N_15381);
xnor U15774 (N_15774,N_15074,N_15277);
and U15775 (N_15775,N_15111,N_15410);
and U15776 (N_15776,N_15047,N_15250);
and U15777 (N_15777,N_15269,N_15376);
or U15778 (N_15778,N_15239,N_15218);
or U15779 (N_15779,N_15296,N_15150);
and U15780 (N_15780,N_15351,N_15251);
nor U15781 (N_15781,N_15019,N_15242);
and U15782 (N_15782,N_15043,N_15369);
or U15783 (N_15783,N_15317,N_15272);
nand U15784 (N_15784,N_15386,N_15266);
nor U15785 (N_15785,N_15394,N_15077);
xnor U15786 (N_15786,N_15421,N_15400);
nor U15787 (N_15787,N_15320,N_15241);
nor U15788 (N_15788,N_15243,N_15200);
xor U15789 (N_15789,N_15018,N_15292);
nand U15790 (N_15790,N_15208,N_15058);
nor U15791 (N_15791,N_15032,N_15312);
nor U15792 (N_15792,N_15129,N_15206);
and U15793 (N_15793,N_15198,N_15494);
and U15794 (N_15794,N_15222,N_15356);
nor U15795 (N_15795,N_15245,N_15371);
and U15796 (N_15796,N_15002,N_15312);
or U15797 (N_15797,N_15221,N_15285);
and U15798 (N_15798,N_15241,N_15453);
or U15799 (N_15799,N_15087,N_15163);
nand U15800 (N_15800,N_15231,N_15164);
nor U15801 (N_15801,N_15114,N_15139);
nand U15802 (N_15802,N_15020,N_15365);
nand U15803 (N_15803,N_15385,N_15097);
and U15804 (N_15804,N_15144,N_15362);
nand U15805 (N_15805,N_15084,N_15220);
xnor U15806 (N_15806,N_15263,N_15456);
nand U15807 (N_15807,N_15104,N_15303);
or U15808 (N_15808,N_15276,N_15328);
and U15809 (N_15809,N_15315,N_15286);
xor U15810 (N_15810,N_15392,N_15209);
or U15811 (N_15811,N_15319,N_15141);
nand U15812 (N_15812,N_15495,N_15224);
nor U15813 (N_15813,N_15074,N_15276);
nor U15814 (N_15814,N_15247,N_15456);
nand U15815 (N_15815,N_15337,N_15325);
xnor U15816 (N_15816,N_15334,N_15274);
nand U15817 (N_15817,N_15463,N_15149);
nand U15818 (N_15818,N_15309,N_15351);
and U15819 (N_15819,N_15315,N_15316);
or U15820 (N_15820,N_15446,N_15361);
nand U15821 (N_15821,N_15208,N_15270);
nand U15822 (N_15822,N_15088,N_15096);
nor U15823 (N_15823,N_15349,N_15254);
nand U15824 (N_15824,N_15074,N_15375);
nor U15825 (N_15825,N_15020,N_15041);
or U15826 (N_15826,N_15319,N_15090);
and U15827 (N_15827,N_15498,N_15446);
or U15828 (N_15828,N_15257,N_15083);
xor U15829 (N_15829,N_15394,N_15420);
xnor U15830 (N_15830,N_15008,N_15044);
nor U15831 (N_15831,N_15177,N_15093);
nor U15832 (N_15832,N_15165,N_15303);
xnor U15833 (N_15833,N_15407,N_15442);
nand U15834 (N_15834,N_15145,N_15163);
nor U15835 (N_15835,N_15017,N_15446);
nand U15836 (N_15836,N_15292,N_15057);
nand U15837 (N_15837,N_15081,N_15171);
and U15838 (N_15838,N_15108,N_15219);
and U15839 (N_15839,N_15295,N_15281);
nand U15840 (N_15840,N_15056,N_15336);
nand U15841 (N_15841,N_15477,N_15387);
nand U15842 (N_15842,N_15017,N_15294);
nand U15843 (N_15843,N_15106,N_15103);
nand U15844 (N_15844,N_15148,N_15283);
nand U15845 (N_15845,N_15199,N_15422);
nor U15846 (N_15846,N_15201,N_15198);
nor U15847 (N_15847,N_15101,N_15264);
nor U15848 (N_15848,N_15240,N_15313);
and U15849 (N_15849,N_15187,N_15051);
xor U15850 (N_15850,N_15497,N_15048);
and U15851 (N_15851,N_15243,N_15004);
and U15852 (N_15852,N_15342,N_15202);
and U15853 (N_15853,N_15272,N_15135);
nor U15854 (N_15854,N_15353,N_15128);
and U15855 (N_15855,N_15337,N_15458);
and U15856 (N_15856,N_15202,N_15488);
nor U15857 (N_15857,N_15217,N_15064);
xnor U15858 (N_15858,N_15186,N_15391);
xnor U15859 (N_15859,N_15417,N_15430);
xnor U15860 (N_15860,N_15488,N_15256);
nor U15861 (N_15861,N_15140,N_15484);
nor U15862 (N_15862,N_15477,N_15452);
or U15863 (N_15863,N_15021,N_15430);
and U15864 (N_15864,N_15389,N_15455);
and U15865 (N_15865,N_15445,N_15247);
or U15866 (N_15866,N_15249,N_15288);
nor U15867 (N_15867,N_15422,N_15480);
nor U15868 (N_15868,N_15467,N_15280);
and U15869 (N_15869,N_15428,N_15346);
xor U15870 (N_15870,N_15449,N_15355);
xnor U15871 (N_15871,N_15229,N_15336);
xor U15872 (N_15872,N_15407,N_15084);
nand U15873 (N_15873,N_15131,N_15243);
xnor U15874 (N_15874,N_15353,N_15070);
xnor U15875 (N_15875,N_15143,N_15476);
xor U15876 (N_15876,N_15342,N_15431);
nor U15877 (N_15877,N_15437,N_15323);
nand U15878 (N_15878,N_15435,N_15327);
xor U15879 (N_15879,N_15471,N_15223);
nor U15880 (N_15880,N_15009,N_15273);
or U15881 (N_15881,N_15406,N_15407);
or U15882 (N_15882,N_15180,N_15257);
and U15883 (N_15883,N_15345,N_15019);
or U15884 (N_15884,N_15021,N_15401);
xnor U15885 (N_15885,N_15256,N_15048);
or U15886 (N_15886,N_15357,N_15494);
and U15887 (N_15887,N_15221,N_15054);
nor U15888 (N_15888,N_15243,N_15023);
and U15889 (N_15889,N_15275,N_15374);
nand U15890 (N_15890,N_15144,N_15282);
nand U15891 (N_15891,N_15012,N_15251);
xnor U15892 (N_15892,N_15091,N_15422);
xor U15893 (N_15893,N_15064,N_15171);
xnor U15894 (N_15894,N_15264,N_15092);
xor U15895 (N_15895,N_15076,N_15446);
or U15896 (N_15896,N_15146,N_15297);
xnor U15897 (N_15897,N_15320,N_15211);
or U15898 (N_15898,N_15381,N_15043);
nand U15899 (N_15899,N_15488,N_15388);
nand U15900 (N_15900,N_15252,N_15032);
nor U15901 (N_15901,N_15048,N_15026);
nand U15902 (N_15902,N_15301,N_15142);
nand U15903 (N_15903,N_15264,N_15211);
xnor U15904 (N_15904,N_15312,N_15087);
xor U15905 (N_15905,N_15320,N_15051);
and U15906 (N_15906,N_15246,N_15047);
xnor U15907 (N_15907,N_15025,N_15406);
nor U15908 (N_15908,N_15311,N_15020);
nand U15909 (N_15909,N_15109,N_15052);
nand U15910 (N_15910,N_15212,N_15312);
nand U15911 (N_15911,N_15400,N_15432);
or U15912 (N_15912,N_15077,N_15180);
nor U15913 (N_15913,N_15175,N_15328);
xnor U15914 (N_15914,N_15159,N_15454);
nand U15915 (N_15915,N_15243,N_15467);
or U15916 (N_15916,N_15351,N_15223);
and U15917 (N_15917,N_15261,N_15136);
nor U15918 (N_15918,N_15337,N_15334);
or U15919 (N_15919,N_15012,N_15304);
nand U15920 (N_15920,N_15336,N_15343);
nor U15921 (N_15921,N_15332,N_15469);
xnor U15922 (N_15922,N_15081,N_15469);
and U15923 (N_15923,N_15291,N_15488);
xnor U15924 (N_15924,N_15492,N_15033);
nand U15925 (N_15925,N_15017,N_15214);
nor U15926 (N_15926,N_15105,N_15373);
and U15927 (N_15927,N_15057,N_15394);
and U15928 (N_15928,N_15184,N_15279);
nand U15929 (N_15929,N_15266,N_15315);
nand U15930 (N_15930,N_15234,N_15324);
or U15931 (N_15931,N_15217,N_15372);
nor U15932 (N_15932,N_15044,N_15258);
xnor U15933 (N_15933,N_15084,N_15269);
or U15934 (N_15934,N_15148,N_15125);
or U15935 (N_15935,N_15416,N_15362);
nand U15936 (N_15936,N_15147,N_15397);
nor U15937 (N_15937,N_15345,N_15067);
and U15938 (N_15938,N_15455,N_15217);
nand U15939 (N_15939,N_15068,N_15408);
or U15940 (N_15940,N_15051,N_15053);
nor U15941 (N_15941,N_15469,N_15186);
xnor U15942 (N_15942,N_15285,N_15401);
nor U15943 (N_15943,N_15062,N_15248);
nand U15944 (N_15944,N_15006,N_15258);
nor U15945 (N_15945,N_15013,N_15178);
nand U15946 (N_15946,N_15431,N_15483);
xnor U15947 (N_15947,N_15046,N_15108);
xnor U15948 (N_15948,N_15094,N_15344);
or U15949 (N_15949,N_15290,N_15154);
and U15950 (N_15950,N_15014,N_15391);
xnor U15951 (N_15951,N_15036,N_15026);
or U15952 (N_15952,N_15199,N_15241);
nand U15953 (N_15953,N_15191,N_15363);
xor U15954 (N_15954,N_15074,N_15129);
and U15955 (N_15955,N_15048,N_15488);
nand U15956 (N_15956,N_15379,N_15038);
xor U15957 (N_15957,N_15295,N_15250);
xor U15958 (N_15958,N_15459,N_15209);
nor U15959 (N_15959,N_15100,N_15411);
and U15960 (N_15960,N_15405,N_15122);
nand U15961 (N_15961,N_15298,N_15207);
xnor U15962 (N_15962,N_15455,N_15060);
or U15963 (N_15963,N_15216,N_15385);
xor U15964 (N_15964,N_15064,N_15237);
xor U15965 (N_15965,N_15034,N_15086);
and U15966 (N_15966,N_15319,N_15126);
xnor U15967 (N_15967,N_15074,N_15041);
nor U15968 (N_15968,N_15392,N_15192);
and U15969 (N_15969,N_15075,N_15417);
and U15970 (N_15970,N_15074,N_15359);
and U15971 (N_15971,N_15081,N_15312);
nand U15972 (N_15972,N_15229,N_15008);
nand U15973 (N_15973,N_15061,N_15085);
nand U15974 (N_15974,N_15109,N_15320);
nand U15975 (N_15975,N_15394,N_15339);
or U15976 (N_15976,N_15372,N_15429);
nor U15977 (N_15977,N_15479,N_15116);
and U15978 (N_15978,N_15124,N_15052);
xnor U15979 (N_15979,N_15494,N_15131);
nor U15980 (N_15980,N_15463,N_15176);
xor U15981 (N_15981,N_15216,N_15001);
and U15982 (N_15982,N_15257,N_15028);
nand U15983 (N_15983,N_15479,N_15168);
xor U15984 (N_15984,N_15215,N_15425);
nor U15985 (N_15985,N_15259,N_15380);
nor U15986 (N_15986,N_15087,N_15493);
xnor U15987 (N_15987,N_15401,N_15189);
or U15988 (N_15988,N_15262,N_15196);
or U15989 (N_15989,N_15275,N_15264);
and U15990 (N_15990,N_15202,N_15136);
nor U15991 (N_15991,N_15024,N_15119);
or U15992 (N_15992,N_15250,N_15069);
xnor U15993 (N_15993,N_15135,N_15442);
nor U15994 (N_15994,N_15235,N_15321);
or U15995 (N_15995,N_15405,N_15482);
and U15996 (N_15996,N_15182,N_15079);
nand U15997 (N_15997,N_15164,N_15476);
nor U15998 (N_15998,N_15221,N_15323);
nand U15999 (N_15999,N_15019,N_15490);
and U16000 (N_16000,N_15784,N_15976);
xnor U16001 (N_16001,N_15850,N_15759);
nor U16002 (N_16002,N_15582,N_15694);
nor U16003 (N_16003,N_15924,N_15898);
and U16004 (N_16004,N_15527,N_15584);
or U16005 (N_16005,N_15516,N_15608);
xor U16006 (N_16006,N_15579,N_15642);
nor U16007 (N_16007,N_15792,N_15842);
and U16008 (N_16008,N_15502,N_15816);
nor U16009 (N_16009,N_15671,N_15514);
nand U16010 (N_16010,N_15674,N_15625);
or U16011 (N_16011,N_15756,N_15830);
nor U16012 (N_16012,N_15847,N_15856);
nand U16013 (N_16013,N_15628,N_15989);
nor U16014 (N_16014,N_15656,N_15611);
xor U16015 (N_16015,N_15602,N_15869);
and U16016 (N_16016,N_15963,N_15787);
nor U16017 (N_16017,N_15509,N_15624);
or U16018 (N_16018,N_15866,N_15889);
xnor U16019 (N_16019,N_15843,N_15603);
nor U16020 (N_16020,N_15743,N_15551);
and U16021 (N_16021,N_15685,N_15931);
nor U16022 (N_16022,N_15814,N_15712);
and U16023 (N_16023,N_15553,N_15948);
and U16024 (N_16024,N_15996,N_15960);
and U16025 (N_16025,N_15583,N_15926);
nand U16026 (N_16026,N_15728,N_15880);
xor U16027 (N_16027,N_15914,N_15615);
xnor U16028 (N_16028,N_15886,N_15975);
and U16029 (N_16029,N_15910,N_15723);
or U16030 (N_16030,N_15557,N_15770);
and U16031 (N_16031,N_15697,N_15987);
nor U16032 (N_16032,N_15979,N_15892);
xnor U16033 (N_16033,N_15760,N_15517);
nor U16034 (N_16034,N_15610,N_15523);
nor U16035 (N_16035,N_15537,N_15581);
and U16036 (N_16036,N_15844,N_15765);
nand U16037 (N_16037,N_15675,N_15563);
and U16038 (N_16038,N_15994,N_15676);
or U16039 (N_16039,N_15564,N_15706);
nand U16040 (N_16040,N_15797,N_15600);
xor U16041 (N_16041,N_15936,N_15790);
nor U16042 (N_16042,N_15710,N_15887);
or U16043 (N_16043,N_15609,N_15932);
or U16044 (N_16044,N_15807,N_15549);
nand U16045 (N_16045,N_15782,N_15944);
and U16046 (N_16046,N_15741,N_15541);
or U16047 (N_16047,N_15641,N_15801);
xor U16048 (N_16048,N_15578,N_15607);
and U16049 (N_16049,N_15528,N_15973);
nand U16050 (N_16050,N_15995,N_15550);
and U16051 (N_16051,N_15588,N_15845);
xnor U16052 (N_16052,N_15954,N_15916);
xnor U16053 (N_16053,N_15907,N_15824);
nor U16054 (N_16054,N_15992,N_15623);
and U16055 (N_16055,N_15590,N_15655);
nand U16056 (N_16056,N_15829,N_15882);
nand U16057 (N_16057,N_15902,N_15651);
nor U16058 (N_16058,N_15638,N_15700);
and U16059 (N_16059,N_15868,N_15633);
and U16060 (N_16060,N_15769,N_15719);
and U16061 (N_16061,N_15666,N_15725);
or U16062 (N_16062,N_15983,N_15632);
or U16063 (N_16063,N_15956,N_15731);
and U16064 (N_16064,N_15503,N_15810);
nor U16065 (N_16065,N_15661,N_15925);
and U16066 (N_16066,N_15640,N_15893);
nor U16067 (N_16067,N_15978,N_15779);
xnor U16068 (N_16068,N_15965,N_15945);
and U16069 (N_16069,N_15686,N_15970);
nand U16070 (N_16070,N_15576,N_15605);
nand U16071 (N_16071,N_15542,N_15683);
xor U16072 (N_16072,N_15967,N_15870);
nand U16073 (N_16073,N_15680,N_15750);
or U16074 (N_16074,N_15653,N_15938);
nand U16075 (N_16075,N_15739,N_15935);
or U16076 (N_16076,N_15665,N_15981);
xor U16077 (N_16077,N_15749,N_15789);
and U16078 (N_16078,N_15679,N_15885);
xnor U16079 (N_16079,N_15668,N_15500);
nor U16080 (N_16080,N_15891,N_15753);
xnor U16081 (N_16081,N_15764,N_15639);
xnor U16082 (N_16082,N_15918,N_15812);
or U16083 (N_16083,N_15673,N_15693);
and U16084 (N_16084,N_15781,N_15606);
nor U16085 (N_16085,N_15861,N_15566);
nand U16086 (N_16086,N_15813,N_15803);
and U16087 (N_16087,N_15835,N_15928);
or U16088 (N_16088,N_15863,N_15802);
xor U16089 (N_16089,N_15592,N_15644);
nor U16090 (N_16090,N_15986,N_15904);
xnor U16091 (N_16091,N_15552,N_15934);
nor U16092 (N_16092,N_15777,N_15630);
and U16093 (N_16093,N_15717,N_15672);
nand U16094 (N_16094,N_15682,N_15727);
or U16095 (N_16095,N_15939,N_15919);
or U16096 (N_16096,N_15718,N_15940);
or U16097 (N_16097,N_15574,N_15993);
and U16098 (N_16098,N_15852,N_15699);
and U16099 (N_16099,N_15800,N_15691);
nand U16100 (N_16100,N_15714,N_15968);
xor U16101 (N_16101,N_15927,N_15732);
and U16102 (N_16102,N_15822,N_15670);
and U16103 (N_16103,N_15874,N_15876);
and U16104 (N_16104,N_15649,N_15601);
nor U16105 (N_16105,N_15821,N_15715);
or U16106 (N_16106,N_15513,N_15833);
or U16107 (N_16107,N_15660,N_15622);
nand U16108 (N_16108,N_15846,N_15867);
nor U16109 (N_16109,N_15818,N_15820);
xnor U16110 (N_16110,N_15562,N_15988);
nor U16111 (N_16111,N_15798,N_15959);
or U16112 (N_16112,N_15937,N_15828);
xnor U16113 (N_16113,N_15594,N_15569);
or U16114 (N_16114,N_15546,N_15524);
or U16115 (N_16115,N_15540,N_15722);
or U16116 (N_16116,N_15751,N_15678);
nor U16117 (N_16117,N_15556,N_15747);
xnor U16118 (N_16118,N_15841,N_15793);
nand U16119 (N_16119,N_15774,N_15883);
or U16120 (N_16120,N_15859,N_15535);
or U16121 (N_16121,N_15646,N_15984);
nand U16122 (N_16122,N_15763,N_15703);
xnor U16123 (N_16123,N_15506,N_15692);
nand U16124 (N_16124,N_15840,N_15571);
or U16125 (N_16125,N_15766,N_15853);
nor U16126 (N_16126,N_15738,N_15545);
nand U16127 (N_16127,N_15532,N_15695);
nor U16128 (N_16128,N_15547,N_15791);
and U16129 (N_16129,N_15626,N_15512);
nor U16130 (N_16130,N_15613,N_15909);
and U16131 (N_16131,N_15966,N_15720);
xnor U16132 (N_16132,N_15754,N_15521);
nand U16133 (N_16133,N_15690,N_15543);
nor U16134 (N_16134,N_15857,N_15554);
xor U16135 (N_16135,N_15825,N_15786);
xor U16136 (N_16136,N_15534,N_15913);
or U16137 (N_16137,N_15999,N_15511);
nor U16138 (N_16138,N_15768,N_15617);
xnor U16139 (N_16139,N_15637,N_15687);
xnor U16140 (N_16140,N_15884,N_15531);
xor U16141 (N_16141,N_15771,N_15575);
xnor U16142 (N_16142,N_15567,N_15930);
and U16143 (N_16143,N_15669,N_15831);
or U16144 (N_16144,N_15878,N_15593);
or U16145 (N_16145,N_15903,N_15808);
and U16146 (N_16146,N_15659,N_15744);
nor U16147 (N_16147,N_15708,N_15775);
nand U16148 (N_16148,N_15538,N_15890);
nor U16149 (N_16149,N_15972,N_15507);
and U16150 (N_16150,N_15619,N_15848);
nand U16151 (N_16151,N_15901,N_15953);
and U16152 (N_16152,N_15572,N_15908);
xnor U16153 (N_16153,N_15565,N_15711);
and U16154 (N_16154,N_15871,N_15614);
nand U16155 (N_16155,N_15520,N_15952);
nor U16156 (N_16156,N_15780,N_15681);
and U16157 (N_16157,N_15804,N_15895);
nand U16158 (N_16158,N_15636,N_15688);
and U16159 (N_16159,N_15875,N_15597);
nor U16160 (N_16160,N_15980,N_15530);
nand U16161 (N_16161,N_15740,N_15746);
and U16162 (N_16162,N_15865,N_15580);
nand U16163 (N_16163,N_15817,N_15709);
nor U16164 (N_16164,N_15839,N_15823);
and U16165 (N_16165,N_15985,N_15595);
nand U16166 (N_16166,N_15634,N_15539);
and U16167 (N_16167,N_15652,N_15618);
nor U16168 (N_16168,N_15827,N_15872);
nand U16169 (N_16169,N_15941,N_15881);
or U16170 (N_16170,N_15604,N_15877);
nor U16171 (N_16171,N_15568,N_15648);
or U16172 (N_16172,N_15589,N_15977);
nor U16173 (N_16173,N_15997,N_15698);
and U16174 (N_16174,N_15947,N_15635);
nor U16175 (N_16175,N_15773,N_15888);
or U16176 (N_16176,N_15742,N_15855);
xnor U16177 (N_16177,N_15707,N_15762);
xnor U16178 (N_16178,N_15923,N_15647);
xor U16179 (N_16179,N_15776,N_15501);
and U16180 (N_16180,N_15806,N_15663);
xnor U16181 (N_16181,N_15561,N_15505);
and U16182 (N_16182,N_15586,N_15677);
nor U16183 (N_16183,N_15555,N_15836);
and U16184 (N_16184,N_15783,N_15849);
and U16185 (N_16185,N_15548,N_15896);
and U16186 (N_16186,N_15757,N_15796);
nor U16187 (N_16187,N_15858,N_15854);
or U16188 (N_16188,N_15826,N_15758);
and U16189 (N_16189,N_15990,N_15544);
xnor U16190 (N_16190,N_15911,N_15529);
nand U16191 (N_16191,N_15974,N_15795);
and U16192 (N_16192,N_15788,N_15522);
nand U16193 (N_16193,N_15658,N_15721);
nor U16194 (N_16194,N_15736,N_15667);
or U16195 (N_16195,N_15819,N_15922);
and U16196 (N_16196,N_15654,N_15929);
xor U16197 (N_16197,N_15864,N_15696);
nor U16198 (N_16198,N_15643,N_15533);
and U16199 (N_16199,N_15778,N_15612);
or U16200 (N_16200,N_15900,N_15573);
nand U16201 (N_16201,N_15942,N_15964);
nor U16202 (N_16202,N_15745,N_15689);
xor U16203 (N_16203,N_15621,N_15799);
or U16204 (N_16204,N_15724,N_15950);
or U16205 (N_16205,N_15519,N_15794);
and U16206 (N_16206,N_15525,N_15627);
nor U16207 (N_16207,N_15917,N_15933);
nor U16208 (N_16208,N_15591,N_15832);
or U16209 (N_16209,N_15899,N_15815);
xnor U16210 (N_16210,N_15838,N_15599);
or U16211 (N_16211,N_15958,N_15915);
and U16212 (N_16212,N_15596,N_15716);
nor U16213 (N_16213,N_15704,N_15734);
and U16214 (N_16214,N_15735,N_15726);
nand U16215 (N_16215,N_15920,N_15657);
xnor U16216 (N_16216,N_15905,N_15730);
xor U16217 (N_16217,N_15733,N_15961);
and U16218 (N_16218,N_15629,N_15862);
nand U16219 (N_16219,N_15515,N_15631);
nor U16220 (N_16220,N_15684,N_15752);
or U16221 (N_16221,N_15748,N_15587);
nand U16222 (N_16222,N_15897,N_15616);
nand U16223 (N_16223,N_15526,N_15921);
and U16224 (N_16224,N_15664,N_15620);
nand U16225 (N_16225,N_15701,N_15772);
or U16226 (N_16226,N_15971,N_15949);
and U16227 (N_16227,N_15645,N_15510);
nor U16228 (N_16228,N_15508,N_15577);
and U16229 (N_16229,N_15851,N_15504);
or U16230 (N_16230,N_15834,N_15705);
or U16231 (N_16231,N_15873,N_15957);
xor U16232 (N_16232,N_15906,N_15946);
nand U16233 (N_16233,N_15809,N_15991);
nor U16234 (N_16234,N_15598,N_15650);
or U16235 (N_16235,N_15761,N_15837);
and U16236 (N_16236,N_15955,N_15570);
xor U16237 (N_16237,N_15785,N_15951);
xnor U16238 (N_16238,N_15894,N_15962);
xnor U16239 (N_16239,N_15879,N_15982);
or U16240 (N_16240,N_15811,N_15805);
nor U16241 (N_16241,N_15713,N_15860);
and U16242 (N_16242,N_15518,N_15662);
nor U16243 (N_16243,N_15998,N_15559);
xnor U16244 (N_16244,N_15702,N_15536);
and U16245 (N_16245,N_15912,N_15755);
nand U16246 (N_16246,N_15943,N_15585);
or U16247 (N_16247,N_15729,N_15969);
or U16248 (N_16248,N_15767,N_15560);
or U16249 (N_16249,N_15558,N_15737);
and U16250 (N_16250,N_15929,N_15676);
nor U16251 (N_16251,N_15621,N_15726);
nand U16252 (N_16252,N_15630,N_15628);
xnor U16253 (N_16253,N_15986,N_15532);
xor U16254 (N_16254,N_15727,N_15557);
xnor U16255 (N_16255,N_15568,N_15563);
nor U16256 (N_16256,N_15641,N_15745);
or U16257 (N_16257,N_15855,N_15686);
nand U16258 (N_16258,N_15535,N_15903);
nor U16259 (N_16259,N_15858,N_15504);
nor U16260 (N_16260,N_15802,N_15919);
xor U16261 (N_16261,N_15848,N_15957);
or U16262 (N_16262,N_15648,N_15959);
nand U16263 (N_16263,N_15843,N_15812);
nor U16264 (N_16264,N_15655,N_15899);
nand U16265 (N_16265,N_15786,N_15910);
nor U16266 (N_16266,N_15858,N_15933);
nor U16267 (N_16267,N_15665,N_15835);
or U16268 (N_16268,N_15638,N_15663);
nor U16269 (N_16269,N_15649,N_15820);
nor U16270 (N_16270,N_15876,N_15653);
and U16271 (N_16271,N_15568,N_15912);
xnor U16272 (N_16272,N_15901,N_15793);
and U16273 (N_16273,N_15809,N_15931);
nand U16274 (N_16274,N_15861,N_15799);
or U16275 (N_16275,N_15516,N_15856);
or U16276 (N_16276,N_15597,N_15909);
or U16277 (N_16277,N_15722,N_15721);
nor U16278 (N_16278,N_15802,N_15635);
nor U16279 (N_16279,N_15902,N_15733);
nand U16280 (N_16280,N_15802,N_15850);
nand U16281 (N_16281,N_15615,N_15664);
and U16282 (N_16282,N_15859,N_15884);
or U16283 (N_16283,N_15765,N_15583);
and U16284 (N_16284,N_15899,N_15838);
nor U16285 (N_16285,N_15619,N_15935);
nor U16286 (N_16286,N_15529,N_15742);
nand U16287 (N_16287,N_15646,N_15848);
nand U16288 (N_16288,N_15623,N_15718);
nand U16289 (N_16289,N_15806,N_15936);
nor U16290 (N_16290,N_15679,N_15716);
nand U16291 (N_16291,N_15856,N_15845);
xor U16292 (N_16292,N_15681,N_15750);
nor U16293 (N_16293,N_15544,N_15944);
nand U16294 (N_16294,N_15844,N_15856);
nand U16295 (N_16295,N_15683,N_15525);
and U16296 (N_16296,N_15643,N_15874);
nor U16297 (N_16297,N_15508,N_15532);
and U16298 (N_16298,N_15786,N_15923);
and U16299 (N_16299,N_15717,N_15686);
or U16300 (N_16300,N_15940,N_15550);
nor U16301 (N_16301,N_15924,N_15698);
nor U16302 (N_16302,N_15827,N_15957);
or U16303 (N_16303,N_15673,N_15887);
or U16304 (N_16304,N_15815,N_15529);
nor U16305 (N_16305,N_15844,N_15978);
or U16306 (N_16306,N_15939,N_15665);
or U16307 (N_16307,N_15888,N_15601);
nor U16308 (N_16308,N_15819,N_15635);
xnor U16309 (N_16309,N_15588,N_15722);
or U16310 (N_16310,N_15681,N_15707);
xnor U16311 (N_16311,N_15775,N_15685);
and U16312 (N_16312,N_15588,N_15728);
xor U16313 (N_16313,N_15646,N_15559);
nor U16314 (N_16314,N_15512,N_15798);
nand U16315 (N_16315,N_15736,N_15746);
or U16316 (N_16316,N_15744,N_15848);
nand U16317 (N_16317,N_15877,N_15636);
nor U16318 (N_16318,N_15951,N_15982);
and U16319 (N_16319,N_15666,N_15862);
and U16320 (N_16320,N_15798,N_15671);
nand U16321 (N_16321,N_15651,N_15940);
and U16322 (N_16322,N_15766,N_15633);
nor U16323 (N_16323,N_15611,N_15781);
nand U16324 (N_16324,N_15829,N_15526);
xnor U16325 (N_16325,N_15758,N_15835);
xor U16326 (N_16326,N_15690,N_15963);
or U16327 (N_16327,N_15923,N_15506);
xnor U16328 (N_16328,N_15549,N_15895);
xnor U16329 (N_16329,N_15516,N_15640);
and U16330 (N_16330,N_15542,N_15841);
and U16331 (N_16331,N_15546,N_15826);
nor U16332 (N_16332,N_15521,N_15801);
xnor U16333 (N_16333,N_15901,N_15516);
and U16334 (N_16334,N_15988,N_15638);
and U16335 (N_16335,N_15781,N_15830);
xnor U16336 (N_16336,N_15856,N_15514);
nor U16337 (N_16337,N_15565,N_15680);
xor U16338 (N_16338,N_15985,N_15602);
or U16339 (N_16339,N_15775,N_15521);
or U16340 (N_16340,N_15791,N_15984);
and U16341 (N_16341,N_15662,N_15957);
and U16342 (N_16342,N_15914,N_15589);
or U16343 (N_16343,N_15667,N_15689);
nand U16344 (N_16344,N_15731,N_15888);
nor U16345 (N_16345,N_15732,N_15829);
nand U16346 (N_16346,N_15717,N_15893);
and U16347 (N_16347,N_15906,N_15793);
nor U16348 (N_16348,N_15569,N_15505);
and U16349 (N_16349,N_15855,N_15565);
or U16350 (N_16350,N_15833,N_15737);
xnor U16351 (N_16351,N_15584,N_15978);
or U16352 (N_16352,N_15879,N_15685);
nor U16353 (N_16353,N_15586,N_15986);
xnor U16354 (N_16354,N_15669,N_15687);
or U16355 (N_16355,N_15667,N_15709);
xor U16356 (N_16356,N_15547,N_15970);
or U16357 (N_16357,N_15513,N_15655);
xnor U16358 (N_16358,N_15774,N_15871);
nand U16359 (N_16359,N_15814,N_15975);
nor U16360 (N_16360,N_15870,N_15738);
nand U16361 (N_16361,N_15749,N_15752);
nand U16362 (N_16362,N_15868,N_15937);
or U16363 (N_16363,N_15978,N_15586);
and U16364 (N_16364,N_15720,N_15866);
nor U16365 (N_16365,N_15783,N_15822);
and U16366 (N_16366,N_15718,N_15916);
xor U16367 (N_16367,N_15814,N_15521);
nand U16368 (N_16368,N_15982,N_15662);
nand U16369 (N_16369,N_15677,N_15856);
or U16370 (N_16370,N_15637,N_15780);
or U16371 (N_16371,N_15638,N_15670);
nor U16372 (N_16372,N_15817,N_15593);
nor U16373 (N_16373,N_15673,N_15800);
or U16374 (N_16374,N_15671,N_15527);
xnor U16375 (N_16375,N_15902,N_15668);
nand U16376 (N_16376,N_15553,N_15589);
xnor U16377 (N_16377,N_15714,N_15980);
nor U16378 (N_16378,N_15533,N_15627);
nand U16379 (N_16379,N_15700,N_15869);
or U16380 (N_16380,N_15520,N_15950);
nor U16381 (N_16381,N_15989,N_15583);
nand U16382 (N_16382,N_15889,N_15693);
or U16383 (N_16383,N_15576,N_15767);
and U16384 (N_16384,N_15626,N_15848);
and U16385 (N_16385,N_15878,N_15889);
nor U16386 (N_16386,N_15825,N_15741);
or U16387 (N_16387,N_15948,N_15776);
xor U16388 (N_16388,N_15896,N_15525);
nor U16389 (N_16389,N_15729,N_15586);
nand U16390 (N_16390,N_15671,N_15512);
xor U16391 (N_16391,N_15811,N_15920);
nand U16392 (N_16392,N_15803,N_15700);
or U16393 (N_16393,N_15567,N_15524);
and U16394 (N_16394,N_15590,N_15561);
nand U16395 (N_16395,N_15522,N_15961);
nand U16396 (N_16396,N_15602,N_15921);
nand U16397 (N_16397,N_15928,N_15791);
nand U16398 (N_16398,N_15735,N_15756);
xnor U16399 (N_16399,N_15752,N_15963);
nor U16400 (N_16400,N_15707,N_15720);
nand U16401 (N_16401,N_15696,N_15673);
nand U16402 (N_16402,N_15797,N_15746);
and U16403 (N_16403,N_15817,N_15715);
or U16404 (N_16404,N_15593,N_15583);
xor U16405 (N_16405,N_15926,N_15652);
nand U16406 (N_16406,N_15588,N_15781);
or U16407 (N_16407,N_15579,N_15634);
xor U16408 (N_16408,N_15794,N_15952);
xor U16409 (N_16409,N_15776,N_15992);
nor U16410 (N_16410,N_15914,N_15748);
xnor U16411 (N_16411,N_15563,N_15853);
xnor U16412 (N_16412,N_15879,N_15551);
nand U16413 (N_16413,N_15918,N_15927);
nand U16414 (N_16414,N_15713,N_15715);
or U16415 (N_16415,N_15516,N_15545);
nand U16416 (N_16416,N_15589,N_15605);
nor U16417 (N_16417,N_15991,N_15553);
or U16418 (N_16418,N_15887,N_15508);
nand U16419 (N_16419,N_15694,N_15653);
and U16420 (N_16420,N_15974,N_15880);
nor U16421 (N_16421,N_15934,N_15619);
and U16422 (N_16422,N_15832,N_15818);
nor U16423 (N_16423,N_15515,N_15936);
xor U16424 (N_16424,N_15675,N_15933);
nor U16425 (N_16425,N_15929,N_15825);
nor U16426 (N_16426,N_15553,N_15852);
nor U16427 (N_16427,N_15765,N_15947);
or U16428 (N_16428,N_15708,N_15568);
xnor U16429 (N_16429,N_15870,N_15700);
nand U16430 (N_16430,N_15768,N_15518);
nor U16431 (N_16431,N_15901,N_15847);
nor U16432 (N_16432,N_15567,N_15902);
and U16433 (N_16433,N_15899,N_15560);
nand U16434 (N_16434,N_15639,N_15892);
nand U16435 (N_16435,N_15621,N_15879);
nand U16436 (N_16436,N_15958,N_15880);
nand U16437 (N_16437,N_15897,N_15531);
and U16438 (N_16438,N_15706,N_15521);
nor U16439 (N_16439,N_15621,N_15500);
nor U16440 (N_16440,N_15889,N_15611);
xor U16441 (N_16441,N_15581,N_15561);
nand U16442 (N_16442,N_15927,N_15504);
nor U16443 (N_16443,N_15991,N_15536);
nor U16444 (N_16444,N_15708,N_15834);
or U16445 (N_16445,N_15511,N_15988);
and U16446 (N_16446,N_15722,N_15966);
or U16447 (N_16447,N_15695,N_15789);
nand U16448 (N_16448,N_15915,N_15988);
and U16449 (N_16449,N_15546,N_15586);
nor U16450 (N_16450,N_15852,N_15640);
nand U16451 (N_16451,N_15670,N_15737);
xor U16452 (N_16452,N_15813,N_15883);
nor U16453 (N_16453,N_15625,N_15556);
or U16454 (N_16454,N_15751,N_15612);
xor U16455 (N_16455,N_15746,N_15791);
or U16456 (N_16456,N_15613,N_15792);
xnor U16457 (N_16457,N_15670,N_15754);
nand U16458 (N_16458,N_15574,N_15648);
and U16459 (N_16459,N_15557,N_15691);
xnor U16460 (N_16460,N_15927,N_15707);
xnor U16461 (N_16461,N_15971,N_15614);
xnor U16462 (N_16462,N_15674,N_15586);
nand U16463 (N_16463,N_15918,N_15923);
nand U16464 (N_16464,N_15922,N_15716);
nor U16465 (N_16465,N_15750,N_15592);
or U16466 (N_16466,N_15571,N_15597);
xor U16467 (N_16467,N_15554,N_15831);
nand U16468 (N_16468,N_15991,N_15512);
xor U16469 (N_16469,N_15895,N_15539);
nand U16470 (N_16470,N_15542,N_15949);
nor U16471 (N_16471,N_15770,N_15627);
xor U16472 (N_16472,N_15790,N_15969);
and U16473 (N_16473,N_15725,N_15536);
and U16474 (N_16474,N_15601,N_15698);
nand U16475 (N_16475,N_15546,N_15722);
xnor U16476 (N_16476,N_15793,N_15747);
nor U16477 (N_16477,N_15551,N_15947);
nand U16478 (N_16478,N_15585,N_15876);
nand U16479 (N_16479,N_15959,N_15976);
nand U16480 (N_16480,N_15732,N_15790);
and U16481 (N_16481,N_15880,N_15532);
nor U16482 (N_16482,N_15788,N_15665);
xnor U16483 (N_16483,N_15880,N_15690);
nand U16484 (N_16484,N_15764,N_15664);
or U16485 (N_16485,N_15629,N_15877);
and U16486 (N_16486,N_15935,N_15906);
nor U16487 (N_16487,N_15657,N_15553);
nand U16488 (N_16488,N_15581,N_15618);
nand U16489 (N_16489,N_15829,N_15635);
and U16490 (N_16490,N_15505,N_15970);
nand U16491 (N_16491,N_15619,N_15603);
and U16492 (N_16492,N_15724,N_15647);
nor U16493 (N_16493,N_15789,N_15697);
and U16494 (N_16494,N_15761,N_15762);
or U16495 (N_16495,N_15524,N_15846);
or U16496 (N_16496,N_15907,N_15713);
nand U16497 (N_16497,N_15729,N_15607);
nand U16498 (N_16498,N_15932,N_15667);
and U16499 (N_16499,N_15673,N_15741);
and U16500 (N_16500,N_16129,N_16448);
and U16501 (N_16501,N_16303,N_16413);
nor U16502 (N_16502,N_16223,N_16384);
nor U16503 (N_16503,N_16302,N_16251);
or U16504 (N_16504,N_16188,N_16086);
xor U16505 (N_16505,N_16265,N_16433);
nand U16506 (N_16506,N_16155,N_16245);
xor U16507 (N_16507,N_16292,N_16009);
xnor U16508 (N_16508,N_16332,N_16197);
xor U16509 (N_16509,N_16154,N_16180);
nand U16510 (N_16510,N_16478,N_16297);
or U16511 (N_16511,N_16058,N_16014);
xor U16512 (N_16512,N_16134,N_16263);
nor U16513 (N_16513,N_16078,N_16214);
xor U16514 (N_16514,N_16125,N_16296);
nor U16515 (N_16515,N_16207,N_16015);
nor U16516 (N_16516,N_16108,N_16010);
and U16517 (N_16517,N_16314,N_16228);
or U16518 (N_16518,N_16226,N_16375);
or U16519 (N_16519,N_16218,N_16311);
nor U16520 (N_16520,N_16221,N_16242);
xor U16521 (N_16521,N_16183,N_16318);
or U16522 (N_16522,N_16094,N_16415);
and U16523 (N_16523,N_16334,N_16372);
or U16524 (N_16524,N_16304,N_16471);
nand U16525 (N_16525,N_16392,N_16167);
nor U16526 (N_16526,N_16117,N_16428);
or U16527 (N_16527,N_16411,N_16164);
nor U16528 (N_16528,N_16212,N_16294);
xor U16529 (N_16529,N_16241,N_16450);
or U16530 (N_16530,N_16016,N_16036);
nor U16531 (N_16531,N_16008,N_16257);
nor U16532 (N_16532,N_16160,N_16333);
or U16533 (N_16533,N_16383,N_16374);
xor U16534 (N_16534,N_16491,N_16140);
or U16535 (N_16535,N_16170,N_16441);
nor U16536 (N_16536,N_16031,N_16176);
nor U16537 (N_16537,N_16330,N_16429);
or U16538 (N_16538,N_16012,N_16208);
xnor U16539 (N_16539,N_16153,N_16168);
and U16540 (N_16540,N_16186,N_16277);
nor U16541 (N_16541,N_16109,N_16427);
xor U16542 (N_16542,N_16486,N_16021);
and U16543 (N_16543,N_16146,N_16145);
nor U16544 (N_16544,N_16071,N_16192);
nor U16545 (N_16545,N_16095,N_16271);
and U16546 (N_16546,N_16417,N_16191);
nor U16547 (N_16547,N_16141,N_16293);
nor U16548 (N_16548,N_16481,N_16085);
or U16549 (N_16549,N_16477,N_16003);
xor U16550 (N_16550,N_16258,N_16139);
xnor U16551 (N_16551,N_16389,N_16060);
nor U16552 (N_16552,N_16329,N_16128);
nor U16553 (N_16553,N_16136,N_16088);
or U16554 (N_16554,N_16361,N_16324);
nor U16555 (N_16555,N_16269,N_16456);
nor U16556 (N_16556,N_16340,N_16222);
xor U16557 (N_16557,N_16284,N_16034);
xnor U16558 (N_16558,N_16341,N_16199);
or U16559 (N_16559,N_16414,N_16490);
nand U16560 (N_16560,N_16252,N_16081);
xnor U16561 (N_16561,N_16150,N_16487);
nand U16562 (N_16562,N_16325,N_16373);
or U16563 (N_16563,N_16469,N_16110);
or U16564 (N_16564,N_16067,N_16326);
xor U16565 (N_16565,N_16460,N_16102);
xor U16566 (N_16566,N_16111,N_16463);
xnor U16567 (N_16567,N_16407,N_16217);
or U16568 (N_16568,N_16026,N_16045);
xnor U16569 (N_16569,N_16187,N_16358);
nor U16570 (N_16570,N_16057,N_16410);
nor U16571 (N_16571,N_16184,N_16126);
nand U16572 (N_16572,N_16204,N_16308);
nand U16573 (N_16573,N_16219,N_16476);
nand U16574 (N_16574,N_16363,N_16113);
xnor U16575 (N_16575,N_16458,N_16143);
or U16576 (N_16576,N_16432,N_16209);
and U16577 (N_16577,N_16062,N_16200);
nand U16578 (N_16578,N_16305,N_16425);
or U16579 (N_16579,N_16457,N_16005);
or U16580 (N_16580,N_16181,N_16416);
or U16581 (N_16581,N_16398,N_16073);
xor U16582 (N_16582,N_16349,N_16243);
or U16583 (N_16583,N_16482,N_16210);
nand U16584 (N_16584,N_16001,N_16017);
nand U16585 (N_16585,N_16230,N_16461);
or U16586 (N_16586,N_16421,N_16422);
nand U16587 (N_16587,N_16420,N_16193);
and U16588 (N_16588,N_16104,N_16087);
and U16589 (N_16589,N_16404,N_16464);
and U16590 (N_16590,N_16229,N_16234);
nor U16591 (N_16591,N_16177,N_16403);
or U16592 (N_16592,N_16352,N_16006);
and U16593 (N_16593,N_16216,N_16494);
xnor U16594 (N_16594,N_16366,N_16479);
xor U16595 (N_16595,N_16118,N_16142);
xnor U16596 (N_16596,N_16247,N_16497);
nor U16597 (N_16597,N_16100,N_16350);
xnor U16598 (N_16598,N_16048,N_16371);
nor U16599 (N_16599,N_16344,N_16198);
xor U16600 (N_16600,N_16158,N_16347);
nand U16601 (N_16601,N_16114,N_16130);
xor U16602 (N_16602,N_16261,N_16260);
or U16603 (N_16603,N_16055,N_16270);
nor U16604 (N_16604,N_16121,N_16038);
xnor U16605 (N_16605,N_16290,N_16443);
nor U16606 (N_16606,N_16323,N_16220);
nand U16607 (N_16607,N_16203,N_16097);
xor U16608 (N_16608,N_16040,N_16238);
and U16609 (N_16609,N_16235,N_16285);
or U16610 (N_16610,N_16054,N_16019);
xnor U16611 (N_16611,N_16339,N_16098);
or U16612 (N_16612,N_16368,N_16163);
nor U16613 (N_16613,N_16262,N_16179);
xor U16614 (N_16614,N_16291,N_16075);
nand U16615 (N_16615,N_16282,N_16107);
nand U16616 (N_16616,N_16239,N_16424);
nand U16617 (N_16617,N_16419,N_16488);
xnor U16618 (N_16618,N_16063,N_16434);
and U16619 (N_16619,N_16059,N_16313);
nand U16620 (N_16620,N_16148,N_16051);
nor U16621 (N_16621,N_16496,N_16056);
nor U16622 (N_16622,N_16231,N_16385);
or U16623 (N_16623,N_16149,N_16091);
nor U16624 (N_16624,N_16024,N_16156);
nor U16625 (N_16625,N_16405,N_16387);
and U16626 (N_16626,N_16236,N_16030);
and U16627 (N_16627,N_16215,N_16233);
and U16628 (N_16628,N_16328,N_16119);
and U16629 (N_16629,N_16396,N_16211);
xor U16630 (N_16630,N_16319,N_16483);
and U16631 (N_16631,N_16072,N_16127);
nor U16632 (N_16632,N_16189,N_16240);
nand U16633 (N_16633,N_16439,N_16224);
nor U16634 (N_16634,N_16190,N_16386);
nor U16635 (N_16635,N_16171,N_16064);
and U16636 (N_16636,N_16336,N_16307);
nand U16637 (N_16637,N_16338,N_16152);
or U16638 (N_16638,N_16266,N_16037);
nand U16639 (N_16639,N_16489,N_16335);
and U16640 (N_16640,N_16409,N_16053);
or U16641 (N_16641,N_16470,N_16165);
nand U16642 (N_16642,N_16213,N_16043);
and U16643 (N_16643,N_16131,N_16356);
and U16644 (N_16644,N_16380,N_16317);
nor U16645 (N_16645,N_16112,N_16011);
nand U16646 (N_16646,N_16173,N_16322);
and U16647 (N_16647,N_16175,N_16096);
and U16648 (N_16648,N_16355,N_16082);
nand U16649 (N_16649,N_16227,N_16115);
nor U16650 (N_16650,N_16312,N_16280);
xor U16651 (N_16651,N_16367,N_16159);
nor U16652 (N_16652,N_16196,N_16103);
nand U16653 (N_16653,N_16437,N_16364);
xor U16654 (N_16654,N_16066,N_16225);
nor U16655 (N_16655,N_16455,N_16378);
or U16656 (N_16656,N_16138,N_16185);
or U16657 (N_16657,N_16089,N_16306);
or U16658 (N_16658,N_16331,N_16452);
or U16659 (N_16659,N_16327,N_16084);
xor U16660 (N_16660,N_16423,N_16298);
xnor U16661 (N_16661,N_16345,N_16273);
or U16662 (N_16662,N_16178,N_16289);
or U16663 (N_16663,N_16388,N_16028);
and U16664 (N_16664,N_16315,N_16157);
xnor U16665 (N_16665,N_16074,N_16281);
xor U16666 (N_16666,N_16249,N_16259);
or U16667 (N_16667,N_16390,N_16246);
nor U16668 (N_16668,N_16474,N_16172);
or U16669 (N_16669,N_16248,N_16473);
and U16670 (N_16670,N_16359,N_16077);
and U16671 (N_16671,N_16357,N_16065);
and U16672 (N_16672,N_16206,N_16391);
xor U16673 (N_16673,N_16162,N_16412);
or U16674 (N_16674,N_16499,N_16498);
xnor U16675 (N_16675,N_16151,N_16124);
xor U16676 (N_16676,N_16083,N_16069);
xnor U16677 (N_16677,N_16309,N_16360);
nand U16678 (N_16678,N_16278,N_16122);
or U16679 (N_16679,N_16301,N_16080);
nor U16680 (N_16680,N_16052,N_16268);
or U16681 (N_16681,N_16394,N_16430);
and U16682 (N_16682,N_16133,N_16046);
nand U16683 (N_16683,N_16254,N_16316);
nand U16684 (N_16684,N_16070,N_16068);
nand U16685 (N_16685,N_16493,N_16022);
or U16686 (N_16686,N_16376,N_16253);
nand U16687 (N_16687,N_16007,N_16406);
nand U16688 (N_16688,N_16274,N_16000);
nand U16689 (N_16689,N_16343,N_16467);
and U16690 (N_16690,N_16029,N_16013);
or U16691 (N_16691,N_16061,N_16279);
or U16692 (N_16692,N_16020,N_16288);
nor U16693 (N_16693,N_16395,N_16362);
nor U16694 (N_16694,N_16342,N_16451);
or U16695 (N_16695,N_16300,N_16050);
and U16696 (N_16696,N_16264,N_16351);
nor U16697 (N_16697,N_16244,N_16093);
and U16698 (N_16698,N_16079,N_16275);
nor U16699 (N_16699,N_16272,N_16166);
nand U16700 (N_16700,N_16436,N_16337);
or U16701 (N_16701,N_16459,N_16431);
nor U16702 (N_16702,N_16426,N_16287);
nand U16703 (N_16703,N_16237,N_16418);
nor U16704 (N_16704,N_16033,N_16480);
nand U16705 (N_16705,N_16047,N_16092);
xnor U16706 (N_16706,N_16381,N_16468);
and U16707 (N_16707,N_16256,N_16018);
nand U16708 (N_16708,N_16002,N_16466);
nor U16709 (N_16709,N_16447,N_16299);
and U16710 (N_16710,N_16472,N_16435);
and U16711 (N_16711,N_16346,N_16377);
nand U16712 (N_16712,N_16397,N_16400);
nor U16713 (N_16713,N_16401,N_16147);
or U16714 (N_16714,N_16202,N_16438);
nor U16715 (N_16715,N_16041,N_16382);
xor U16716 (N_16716,N_16232,N_16025);
and U16717 (N_16717,N_16090,N_16027);
and U16718 (N_16718,N_16123,N_16137);
or U16719 (N_16719,N_16161,N_16169);
nor U16720 (N_16720,N_16379,N_16076);
xor U16721 (N_16721,N_16444,N_16495);
or U16722 (N_16722,N_16408,N_16201);
and U16723 (N_16723,N_16484,N_16320);
or U16724 (N_16724,N_16354,N_16370);
nor U16725 (N_16725,N_16365,N_16250);
and U16726 (N_16726,N_16099,N_16492);
and U16727 (N_16727,N_16120,N_16462);
or U16728 (N_16728,N_16454,N_16485);
or U16729 (N_16729,N_16182,N_16144);
or U16730 (N_16730,N_16004,N_16132);
or U16731 (N_16731,N_16049,N_16348);
and U16732 (N_16732,N_16399,N_16393);
or U16733 (N_16733,N_16035,N_16286);
or U16734 (N_16734,N_16276,N_16174);
nor U16735 (N_16735,N_16295,N_16042);
nand U16736 (N_16736,N_16032,N_16369);
or U16737 (N_16737,N_16255,N_16475);
and U16738 (N_16738,N_16321,N_16106);
or U16739 (N_16739,N_16310,N_16194);
xor U16740 (N_16740,N_16205,N_16267);
nor U16741 (N_16741,N_16442,N_16453);
xor U16742 (N_16742,N_16135,N_16105);
and U16743 (N_16743,N_16402,N_16449);
nand U16744 (N_16744,N_16101,N_16283);
nor U16745 (N_16745,N_16446,N_16440);
nand U16746 (N_16746,N_16039,N_16465);
and U16747 (N_16747,N_16044,N_16116);
or U16748 (N_16748,N_16353,N_16195);
or U16749 (N_16749,N_16445,N_16023);
or U16750 (N_16750,N_16402,N_16130);
or U16751 (N_16751,N_16476,N_16472);
xnor U16752 (N_16752,N_16322,N_16447);
or U16753 (N_16753,N_16028,N_16386);
and U16754 (N_16754,N_16366,N_16290);
nand U16755 (N_16755,N_16345,N_16304);
or U16756 (N_16756,N_16382,N_16132);
nand U16757 (N_16757,N_16403,N_16303);
and U16758 (N_16758,N_16123,N_16126);
and U16759 (N_16759,N_16480,N_16065);
nand U16760 (N_16760,N_16084,N_16282);
and U16761 (N_16761,N_16326,N_16177);
or U16762 (N_16762,N_16386,N_16281);
and U16763 (N_16763,N_16324,N_16137);
xnor U16764 (N_16764,N_16452,N_16329);
and U16765 (N_16765,N_16046,N_16395);
xnor U16766 (N_16766,N_16176,N_16043);
nand U16767 (N_16767,N_16181,N_16461);
nand U16768 (N_16768,N_16129,N_16429);
xnor U16769 (N_16769,N_16294,N_16492);
xnor U16770 (N_16770,N_16418,N_16310);
or U16771 (N_16771,N_16132,N_16138);
and U16772 (N_16772,N_16231,N_16132);
xor U16773 (N_16773,N_16241,N_16246);
and U16774 (N_16774,N_16202,N_16375);
and U16775 (N_16775,N_16288,N_16373);
and U16776 (N_16776,N_16182,N_16422);
or U16777 (N_16777,N_16029,N_16472);
xnor U16778 (N_16778,N_16380,N_16451);
nor U16779 (N_16779,N_16031,N_16040);
and U16780 (N_16780,N_16097,N_16208);
and U16781 (N_16781,N_16214,N_16260);
and U16782 (N_16782,N_16280,N_16472);
nand U16783 (N_16783,N_16079,N_16332);
nand U16784 (N_16784,N_16246,N_16499);
nand U16785 (N_16785,N_16198,N_16249);
nor U16786 (N_16786,N_16491,N_16252);
nor U16787 (N_16787,N_16092,N_16188);
or U16788 (N_16788,N_16012,N_16454);
xor U16789 (N_16789,N_16198,N_16360);
nand U16790 (N_16790,N_16473,N_16358);
nand U16791 (N_16791,N_16397,N_16042);
nand U16792 (N_16792,N_16425,N_16040);
or U16793 (N_16793,N_16214,N_16304);
and U16794 (N_16794,N_16007,N_16015);
xor U16795 (N_16795,N_16442,N_16435);
nand U16796 (N_16796,N_16411,N_16493);
or U16797 (N_16797,N_16449,N_16419);
xor U16798 (N_16798,N_16364,N_16468);
and U16799 (N_16799,N_16259,N_16346);
xor U16800 (N_16800,N_16433,N_16471);
and U16801 (N_16801,N_16485,N_16276);
and U16802 (N_16802,N_16479,N_16150);
or U16803 (N_16803,N_16266,N_16313);
nand U16804 (N_16804,N_16031,N_16008);
and U16805 (N_16805,N_16268,N_16458);
xor U16806 (N_16806,N_16081,N_16416);
and U16807 (N_16807,N_16413,N_16294);
or U16808 (N_16808,N_16461,N_16115);
and U16809 (N_16809,N_16318,N_16018);
and U16810 (N_16810,N_16014,N_16020);
nand U16811 (N_16811,N_16076,N_16498);
or U16812 (N_16812,N_16210,N_16432);
nor U16813 (N_16813,N_16208,N_16315);
xnor U16814 (N_16814,N_16055,N_16451);
nand U16815 (N_16815,N_16472,N_16091);
nand U16816 (N_16816,N_16265,N_16130);
or U16817 (N_16817,N_16310,N_16107);
nand U16818 (N_16818,N_16126,N_16216);
nor U16819 (N_16819,N_16281,N_16202);
and U16820 (N_16820,N_16498,N_16333);
or U16821 (N_16821,N_16267,N_16060);
nand U16822 (N_16822,N_16036,N_16008);
or U16823 (N_16823,N_16313,N_16116);
nor U16824 (N_16824,N_16168,N_16177);
or U16825 (N_16825,N_16085,N_16191);
or U16826 (N_16826,N_16139,N_16244);
nor U16827 (N_16827,N_16472,N_16356);
nand U16828 (N_16828,N_16380,N_16009);
nand U16829 (N_16829,N_16414,N_16261);
and U16830 (N_16830,N_16306,N_16095);
nor U16831 (N_16831,N_16057,N_16174);
xor U16832 (N_16832,N_16078,N_16373);
xnor U16833 (N_16833,N_16167,N_16347);
nor U16834 (N_16834,N_16297,N_16346);
and U16835 (N_16835,N_16088,N_16478);
nor U16836 (N_16836,N_16451,N_16037);
and U16837 (N_16837,N_16373,N_16281);
and U16838 (N_16838,N_16281,N_16177);
nor U16839 (N_16839,N_16270,N_16249);
or U16840 (N_16840,N_16372,N_16252);
nand U16841 (N_16841,N_16351,N_16012);
and U16842 (N_16842,N_16111,N_16327);
xnor U16843 (N_16843,N_16135,N_16469);
nor U16844 (N_16844,N_16420,N_16123);
or U16845 (N_16845,N_16435,N_16477);
and U16846 (N_16846,N_16433,N_16409);
nand U16847 (N_16847,N_16178,N_16120);
or U16848 (N_16848,N_16293,N_16046);
nor U16849 (N_16849,N_16111,N_16060);
nand U16850 (N_16850,N_16417,N_16187);
nand U16851 (N_16851,N_16115,N_16220);
or U16852 (N_16852,N_16372,N_16416);
nor U16853 (N_16853,N_16255,N_16355);
nor U16854 (N_16854,N_16079,N_16411);
nor U16855 (N_16855,N_16183,N_16349);
or U16856 (N_16856,N_16200,N_16269);
or U16857 (N_16857,N_16335,N_16277);
nand U16858 (N_16858,N_16253,N_16076);
and U16859 (N_16859,N_16035,N_16177);
and U16860 (N_16860,N_16421,N_16447);
xor U16861 (N_16861,N_16117,N_16493);
or U16862 (N_16862,N_16162,N_16493);
nor U16863 (N_16863,N_16119,N_16143);
xor U16864 (N_16864,N_16310,N_16049);
xnor U16865 (N_16865,N_16051,N_16090);
nand U16866 (N_16866,N_16237,N_16394);
nor U16867 (N_16867,N_16353,N_16485);
or U16868 (N_16868,N_16225,N_16248);
and U16869 (N_16869,N_16294,N_16053);
xor U16870 (N_16870,N_16294,N_16182);
nand U16871 (N_16871,N_16187,N_16498);
nor U16872 (N_16872,N_16360,N_16231);
xor U16873 (N_16873,N_16443,N_16132);
and U16874 (N_16874,N_16003,N_16447);
nand U16875 (N_16875,N_16027,N_16294);
or U16876 (N_16876,N_16108,N_16274);
and U16877 (N_16877,N_16487,N_16249);
or U16878 (N_16878,N_16102,N_16147);
nor U16879 (N_16879,N_16217,N_16276);
nand U16880 (N_16880,N_16217,N_16352);
or U16881 (N_16881,N_16088,N_16489);
or U16882 (N_16882,N_16345,N_16241);
or U16883 (N_16883,N_16168,N_16354);
xnor U16884 (N_16884,N_16224,N_16213);
nor U16885 (N_16885,N_16321,N_16177);
xor U16886 (N_16886,N_16089,N_16489);
nand U16887 (N_16887,N_16453,N_16062);
xnor U16888 (N_16888,N_16453,N_16252);
xor U16889 (N_16889,N_16242,N_16061);
and U16890 (N_16890,N_16214,N_16138);
xnor U16891 (N_16891,N_16416,N_16385);
xnor U16892 (N_16892,N_16409,N_16194);
xnor U16893 (N_16893,N_16467,N_16104);
nor U16894 (N_16894,N_16012,N_16061);
and U16895 (N_16895,N_16266,N_16152);
nor U16896 (N_16896,N_16308,N_16397);
and U16897 (N_16897,N_16069,N_16027);
or U16898 (N_16898,N_16169,N_16082);
xor U16899 (N_16899,N_16446,N_16058);
or U16900 (N_16900,N_16483,N_16377);
nor U16901 (N_16901,N_16213,N_16255);
nand U16902 (N_16902,N_16280,N_16440);
nor U16903 (N_16903,N_16152,N_16088);
xnor U16904 (N_16904,N_16142,N_16412);
or U16905 (N_16905,N_16306,N_16398);
and U16906 (N_16906,N_16018,N_16483);
nand U16907 (N_16907,N_16135,N_16155);
or U16908 (N_16908,N_16071,N_16460);
xor U16909 (N_16909,N_16342,N_16260);
and U16910 (N_16910,N_16269,N_16008);
and U16911 (N_16911,N_16008,N_16062);
or U16912 (N_16912,N_16289,N_16466);
xor U16913 (N_16913,N_16120,N_16071);
nand U16914 (N_16914,N_16390,N_16427);
or U16915 (N_16915,N_16346,N_16268);
or U16916 (N_16916,N_16396,N_16317);
and U16917 (N_16917,N_16363,N_16299);
nor U16918 (N_16918,N_16253,N_16342);
nor U16919 (N_16919,N_16225,N_16042);
xor U16920 (N_16920,N_16146,N_16041);
nor U16921 (N_16921,N_16307,N_16251);
and U16922 (N_16922,N_16273,N_16076);
nand U16923 (N_16923,N_16202,N_16240);
nor U16924 (N_16924,N_16461,N_16014);
nor U16925 (N_16925,N_16153,N_16348);
xnor U16926 (N_16926,N_16027,N_16219);
nand U16927 (N_16927,N_16019,N_16079);
and U16928 (N_16928,N_16340,N_16129);
and U16929 (N_16929,N_16041,N_16044);
and U16930 (N_16930,N_16128,N_16434);
and U16931 (N_16931,N_16186,N_16143);
and U16932 (N_16932,N_16019,N_16394);
nand U16933 (N_16933,N_16013,N_16106);
nor U16934 (N_16934,N_16162,N_16113);
nor U16935 (N_16935,N_16214,N_16048);
or U16936 (N_16936,N_16136,N_16339);
nor U16937 (N_16937,N_16470,N_16072);
or U16938 (N_16938,N_16192,N_16088);
nand U16939 (N_16939,N_16154,N_16282);
and U16940 (N_16940,N_16184,N_16042);
or U16941 (N_16941,N_16313,N_16415);
and U16942 (N_16942,N_16250,N_16371);
nand U16943 (N_16943,N_16095,N_16460);
xor U16944 (N_16944,N_16367,N_16278);
xnor U16945 (N_16945,N_16419,N_16198);
nor U16946 (N_16946,N_16084,N_16054);
and U16947 (N_16947,N_16170,N_16380);
nand U16948 (N_16948,N_16073,N_16322);
nand U16949 (N_16949,N_16080,N_16363);
or U16950 (N_16950,N_16040,N_16304);
and U16951 (N_16951,N_16013,N_16480);
nand U16952 (N_16952,N_16019,N_16478);
xnor U16953 (N_16953,N_16346,N_16452);
nor U16954 (N_16954,N_16406,N_16353);
and U16955 (N_16955,N_16042,N_16027);
xnor U16956 (N_16956,N_16343,N_16216);
or U16957 (N_16957,N_16355,N_16450);
and U16958 (N_16958,N_16365,N_16196);
and U16959 (N_16959,N_16254,N_16095);
nor U16960 (N_16960,N_16176,N_16053);
or U16961 (N_16961,N_16193,N_16257);
nor U16962 (N_16962,N_16152,N_16075);
nand U16963 (N_16963,N_16355,N_16138);
or U16964 (N_16964,N_16451,N_16371);
or U16965 (N_16965,N_16275,N_16089);
nand U16966 (N_16966,N_16434,N_16174);
nor U16967 (N_16967,N_16357,N_16397);
or U16968 (N_16968,N_16363,N_16200);
xor U16969 (N_16969,N_16394,N_16222);
nor U16970 (N_16970,N_16331,N_16325);
and U16971 (N_16971,N_16479,N_16312);
and U16972 (N_16972,N_16009,N_16148);
nor U16973 (N_16973,N_16037,N_16141);
nor U16974 (N_16974,N_16284,N_16222);
and U16975 (N_16975,N_16454,N_16387);
nand U16976 (N_16976,N_16263,N_16470);
xnor U16977 (N_16977,N_16016,N_16348);
and U16978 (N_16978,N_16099,N_16330);
and U16979 (N_16979,N_16323,N_16335);
or U16980 (N_16980,N_16383,N_16347);
xor U16981 (N_16981,N_16438,N_16412);
xor U16982 (N_16982,N_16055,N_16479);
xnor U16983 (N_16983,N_16498,N_16357);
or U16984 (N_16984,N_16374,N_16440);
nand U16985 (N_16985,N_16268,N_16071);
or U16986 (N_16986,N_16126,N_16354);
nor U16987 (N_16987,N_16494,N_16044);
nor U16988 (N_16988,N_16300,N_16079);
and U16989 (N_16989,N_16171,N_16057);
or U16990 (N_16990,N_16038,N_16088);
or U16991 (N_16991,N_16217,N_16258);
and U16992 (N_16992,N_16050,N_16036);
and U16993 (N_16993,N_16019,N_16253);
nor U16994 (N_16994,N_16494,N_16126);
nand U16995 (N_16995,N_16067,N_16209);
nand U16996 (N_16996,N_16194,N_16469);
or U16997 (N_16997,N_16380,N_16068);
and U16998 (N_16998,N_16142,N_16472);
nor U16999 (N_16999,N_16150,N_16239);
nor U17000 (N_17000,N_16506,N_16637);
and U17001 (N_17001,N_16688,N_16683);
or U17002 (N_17002,N_16949,N_16664);
or U17003 (N_17003,N_16565,N_16734);
and U17004 (N_17004,N_16988,N_16904);
nand U17005 (N_17005,N_16790,N_16969);
nand U17006 (N_17006,N_16566,N_16987);
nand U17007 (N_17007,N_16890,N_16586);
and U17008 (N_17008,N_16797,N_16658);
xor U17009 (N_17009,N_16524,N_16621);
nor U17010 (N_17010,N_16922,N_16775);
and U17011 (N_17011,N_16919,N_16612);
nor U17012 (N_17012,N_16707,N_16542);
nand U17013 (N_17013,N_16980,N_16924);
nand U17014 (N_17014,N_16968,N_16930);
nor U17015 (N_17015,N_16893,N_16654);
xnor U17016 (N_17016,N_16818,N_16653);
nand U17017 (N_17017,N_16527,N_16941);
nand U17018 (N_17018,N_16902,N_16788);
nor U17019 (N_17019,N_16720,N_16856);
nor U17020 (N_17020,N_16846,N_16884);
nor U17021 (N_17021,N_16717,N_16757);
xor U17022 (N_17022,N_16889,N_16912);
xor U17023 (N_17023,N_16598,N_16872);
and U17024 (N_17024,N_16713,N_16859);
xor U17025 (N_17025,N_16594,N_16644);
nand U17026 (N_17026,N_16748,N_16714);
and U17027 (N_17027,N_16840,N_16505);
and U17028 (N_17028,N_16662,N_16845);
nor U17029 (N_17029,N_16557,N_16711);
nor U17030 (N_17030,N_16769,N_16963);
or U17031 (N_17031,N_16920,N_16923);
nor U17032 (N_17032,N_16588,N_16504);
and U17033 (N_17033,N_16752,N_16817);
xor U17034 (N_17034,N_16740,N_16806);
nand U17035 (N_17035,N_16606,N_16511);
xor U17036 (N_17036,N_16521,N_16873);
xor U17037 (N_17037,N_16756,N_16607);
or U17038 (N_17038,N_16648,N_16743);
nor U17039 (N_17039,N_16863,N_16899);
and U17040 (N_17040,N_16955,N_16555);
nor U17041 (N_17041,N_16871,N_16680);
or U17042 (N_17042,N_16731,N_16804);
nand U17043 (N_17043,N_16879,N_16529);
nand U17044 (N_17044,N_16631,N_16992);
and U17045 (N_17045,N_16885,N_16706);
or U17046 (N_17046,N_16967,N_16633);
xnor U17047 (N_17047,N_16576,N_16808);
xor U17048 (N_17048,N_16541,N_16568);
nor U17049 (N_17049,N_16903,N_16772);
nand U17050 (N_17050,N_16852,N_16905);
and U17051 (N_17051,N_16800,N_16767);
nand U17052 (N_17052,N_16689,N_16589);
nor U17053 (N_17053,N_16940,N_16936);
or U17054 (N_17054,N_16866,N_16876);
nand U17055 (N_17055,N_16974,N_16726);
nor U17056 (N_17056,N_16700,N_16661);
and U17057 (N_17057,N_16690,N_16829);
nor U17058 (N_17058,N_16887,N_16552);
nand U17059 (N_17059,N_16971,N_16609);
and U17060 (N_17060,N_16768,N_16815);
nor U17061 (N_17061,N_16771,N_16781);
and U17062 (N_17062,N_16805,N_16533);
nor U17063 (N_17063,N_16693,N_16608);
nor U17064 (N_17064,N_16755,N_16639);
nand U17065 (N_17065,N_16513,N_16641);
xor U17066 (N_17066,N_16675,N_16892);
or U17067 (N_17067,N_16823,N_16735);
and U17068 (N_17068,N_16519,N_16858);
or U17069 (N_17069,N_16616,N_16832);
nor U17070 (N_17070,N_16652,N_16821);
nand U17071 (N_17071,N_16831,N_16710);
nand U17072 (N_17072,N_16684,N_16867);
and U17073 (N_17073,N_16824,N_16965);
and U17074 (N_17074,N_16763,N_16875);
or U17075 (N_17075,N_16750,N_16833);
or U17076 (N_17076,N_16702,N_16766);
nand U17077 (N_17077,N_16929,N_16986);
nand U17078 (N_17078,N_16921,N_16749);
and U17079 (N_17079,N_16628,N_16679);
or U17080 (N_17080,N_16909,N_16878);
nand U17081 (N_17081,N_16956,N_16585);
xnor U17082 (N_17082,N_16843,N_16794);
and U17083 (N_17083,N_16860,N_16786);
and U17084 (N_17084,N_16895,N_16522);
xnor U17085 (N_17085,N_16647,N_16976);
nor U17086 (N_17086,N_16646,N_16877);
nand U17087 (N_17087,N_16593,N_16862);
or U17088 (N_17088,N_16952,N_16882);
nor U17089 (N_17089,N_16869,N_16623);
or U17090 (N_17090,N_16841,N_16667);
nor U17091 (N_17091,N_16881,N_16514);
nor U17092 (N_17092,N_16681,N_16825);
nand U17093 (N_17093,N_16659,N_16666);
nand U17094 (N_17094,N_16914,N_16716);
and U17095 (N_17095,N_16539,N_16729);
and U17096 (N_17096,N_16996,N_16697);
nor U17097 (N_17097,N_16933,N_16886);
and U17098 (N_17098,N_16503,N_16728);
or U17099 (N_17099,N_16855,N_16809);
xor U17100 (N_17100,N_16820,N_16550);
and U17101 (N_17101,N_16709,N_16730);
nor U17102 (N_17102,N_16674,N_16799);
and U17103 (N_17103,N_16977,N_16678);
and U17104 (N_17104,N_16548,N_16959);
or U17105 (N_17105,N_16792,N_16698);
or U17106 (N_17106,N_16634,N_16981);
nand U17107 (N_17107,N_16798,N_16719);
xnor U17108 (N_17108,N_16844,N_16512);
nand U17109 (N_17109,N_16842,N_16906);
nand U17110 (N_17110,N_16642,N_16508);
and U17111 (N_17111,N_16957,N_16701);
or U17112 (N_17112,N_16943,N_16880);
and U17113 (N_17113,N_16733,N_16671);
nor U17114 (N_17114,N_16764,N_16618);
nor U17115 (N_17115,N_16682,N_16838);
and U17116 (N_17116,N_16615,N_16564);
nand U17117 (N_17117,N_16556,N_16962);
xnor U17118 (N_17118,N_16656,N_16970);
and U17119 (N_17119,N_16857,N_16789);
nand U17120 (N_17120,N_16650,N_16972);
nand U17121 (N_17121,N_16934,N_16861);
or U17122 (N_17122,N_16668,N_16783);
or U17123 (N_17123,N_16896,N_16915);
nor U17124 (N_17124,N_16810,N_16526);
nor U17125 (N_17125,N_16651,N_16724);
nand U17126 (N_17126,N_16935,N_16830);
and U17127 (N_17127,N_16629,N_16549);
nand U17128 (N_17128,N_16692,N_16950);
nor U17129 (N_17129,N_16758,N_16672);
xor U17130 (N_17130,N_16649,N_16828);
or U17131 (N_17131,N_16746,N_16907);
nand U17132 (N_17132,N_16993,N_16617);
xnor U17133 (N_17133,N_16534,N_16708);
nor U17134 (N_17134,N_16762,N_16624);
nand U17135 (N_17135,N_16925,N_16500);
and U17136 (N_17136,N_16570,N_16718);
and U17137 (N_17137,N_16520,N_16543);
and U17138 (N_17138,N_16753,N_16917);
nand U17139 (N_17139,N_16677,N_16721);
xnor U17140 (N_17140,N_16747,N_16803);
xor U17141 (N_17141,N_16583,N_16515);
nand U17142 (N_17142,N_16827,N_16793);
xor U17143 (N_17143,N_16913,N_16951);
and U17144 (N_17144,N_16737,N_16540);
and U17145 (N_17145,N_16578,N_16742);
nor U17146 (N_17146,N_16574,N_16632);
and U17147 (N_17147,N_16655,N_16779);
nand U17148 (N_17148,N_16562,N_16791);
nor U17149 (N_17149,N_16625,N_16532);
and U17150 (N_17150,N_16865,N_16979);
nand U17151 (N_17151,N_16812,N_16847);
and U17152 (N_17152,N_16712,N_16501);
and U17153 (N_17153,N_16874,N_16695);
nor U17154 (N_17154,N_16964,N_16705);
nor U17155 (N_17155,N_16989,N_16722);
and U17156 (N_17156,N_16691,N_16638);
and U17157 (N_17157,N_16926,N_16854);
and U17158 (N_17158,N_16911,N_16944);
nand U17159 (N_17159,N_16732,N_16942);
and U17160 (N_17160,N_16599,N_16547);
or U17161 (N_17161,N_16908,N_16813);
xnor U17162 (N_17162,N_16973,N_16814);
nand U17163 (N_17163,N_16773,N_16900);
nand U17164 (N_17164,N_16643,N_16894);
xor U17165 (N_17165,N_16834,N_16745);
or U17166 (N_17166,N_16910,N_16531);
nand U17167 (N_17167,N_16635,N_16751);
nor U17168 (N_17168,N_16960,N_16610);
or U17169 (N_17169,N_16984,N_16961);
xor U17170 (N_17170,N_16560,N_16736);
or U17171 (N_17171,N_16597,N_16850);
or U17172 (N_17172,N_16518,N_16999);
nor U17173 (N_17173,N_16525,N_16928);
xor U17174 (N_17174,N_16581,N_16774);
or U17175 (N_17175,N_16660,N_16580);
xor U17176 (N_17176,N_16554,N_16901);
or U17177 (N_17177,N_16537,N_16613);
xor U17178 (N_17178,N_16620,N_16897);
xnor U17179 (N_17179,N_16538,N_16782);
nand U17180 (N_17180,N_16918,N_16528);
xnor U17181 (N_17181,N_16811,N_16535);
and U17182 (N_17182,N_16777,N_16946);
xnor U17183 (N_17183,N_16727,N_16725);
or U17184 (N_17184,N_16669,N_16738);
and U17185 (N_17185,N_16509,N_16611);
nand U17186 (N_17186,N_16739,N_16851);
nand U17187 (N_17187,N_16559,N_16636);
or U17188 (N_17188,N_16826,N_16523);
xor U17189 (N_17189,N_16600,N_16575);
or U17190 (N_17190,N_16760,N_16807);
or U17191 (N_17191,N_16507,N_16985);
nand U17192 (N_17192,N_16604,N_16948);
nand U17193 (N_17193,N_16868,N_16640);
nand U17194 (N_17194,N_16835,N_16572);
nor U17195 (N_17195,N_16761,N_16978);
or U17196 (N_17196,N_16898,N_16995);
and U17197 (N_17197,N_16991,N_16997);
nor U17198 (N_17198,N_16927,N_16696);
nand U17199 (N_17199,N_16626,N_16590);
nand U17200 (N_17200,N_16770,N_16596);
nand U17201 (N_17201,N_16754,N_16994);
nand U17202 (N_17202,N_16561,N_16787);
or U17203 (N_17203,N_16573,N_16795);
and U17204 (N_17204,N_16545,N_16741);
nand U17205 (N_17205,N_16785,N_16744);
and U17206 (N_17206,N_16990,N_16665);
nor U17207 (N_17207,N_16780,N_16849);
xor U17208 (N_17208,N_16975,N_16853);
or U17209 (N_17209,N_16558,N_16983);
nand U17210 (N_17210,N_16888,N_16546);
and U17211 (N_17211,N_16544,N_16602);
xor U17212 (N_17212,N_16592,N_16802);
and U17213 (N_17213,N_16839,N_16516);
nor U17214 (N_17214,N_16663,N_16510);
nor U17215 (N_17215,N_16954,N_16577);
nand U17216 (N_17216,N_16603,N_16657);
and U17217 (N_17217,N_16703,N_16723);
nor U17218 (N_17218,N_16848,N_16953);
nor U17219 (N_17219,N_16836,N_16982);
nor U17220 (N_17220,N_16605,N_16686);
and U17221 (N_17221,N_16685,N_16776);
and U17222 (N_17222,N_16801,N_16819);
and U17223 (N_17223,N_16816,N_16704);
and U17224 (N_17224,N_16796,N_16587);
nand U17225 (N_17225,N_16567,N_16670);
nand U17226 (N_17226,N_16579,N_16765);
nor U17227 (N_17227,N_16551,N_16939);
nand U17228 (N_17228,N_16931,N_16601);
xor U17229 (N_17229,N_16563,N_16645);
nand U17230 (N_17230,N_16530,N_16571);
xor U17231 (N_17231,N_16947,N_16870);
and U17232 (N_17232,N_16536,N_16627);
xnor U17233 (N_17233,N_16502,N_16864);
nor U17234 (N_17234,N_16595,N_16584);
xnor U17235 (N_17235,N_16673,N_16891);
or U17236 (N_17236,N_16622,N_16937);
nand U17237 (N_17237,N_16619,N_16998);
xor U17238 (N_17238,N_16582,N_16822);
nand U17239 (N_17239,N_16778,N_16694);
and U17240 (N_17240,N_16759,N_16553);
nor U17241 (N_17241,N_16687,N_16715);
xnor U17242 (N_17242,N_16916,N_16958);
nor U17243 (N_17243,N_16591,N_16883);
or U17244 (N_17244,N_16932,N_16630);
nand U17245 (N_17245,N_16966,N_16614);
nor U17246 (N_17246,N_16517,N_16837);
nor U17247 (N_17247,N_16676,N_16699);
nor U17248 (N_17248,N_16569,N_16938);
or U17249 (N_17249,N_16945,N_16784);
xnor U17250 (N_17250,N_16579,N_16507);
xor U17251 (N_17251,N_16577,N_16619);
xnor U17252 (N_17252,N_16667,N_16718);
nand U17253 (N_17253,N_16996,N_16574);
nor U17254 (N_17254,N_16691,N_16883);
or U17255 (N_17255,N_16663,N_16831);
xnor U17256 (N_17256,N_16671,N_16687);
or U17257 (N_17257,N_16660,N_16765);
or U17258 (N_17258,N_16918,N_16549);
xnor U17259 (N_17259,N_16959,N_16843);
nor U17260 (N_17260,N_16526,N_16863);
xor U17261 (N_17261,N_16640,N_16768);
xnor U17262 (N_17262,N_16999,N_16576);
and U17263 (N_17263,N_16751,N_16569);
nor U17264 (N_17264,N_16642,N_16551);
and U17265 (N_17265,N_16572,N_16711);
xnor U17266 (N_17266,N_16804,N_16951);
and U17267 (N_17267,N_16819,N_16908);
xnor U17268 (N_17268,N_16615,N_16995);
and U17269 (N_17269,N_16701,N_16545);
nand U17270 (N_17270,N_16543,N_16771);
or U17271 (N_17271,N_16870,N_16622);
xnor U17272 (N_17272,N_16922,N_16800);
nor U17273 (N_17273,N_16789,N_16815);
or U17274 (N_17274,N_16525,N_16552);
nor U17275 (N_17275,N_16864,N_16836);
nor U17276 (N_17276,N_16855,N_16815);
and U17277 (N_17277,N_16959,N_16674);
nor U17278 (N_17278,N_16930,N_16697);
and U17279 (N_17279,N_16528,N_16991);
nor U17280 (N_17280,N_16829,N_16700);
or U17281 (N_17281,N_16560,N_16886);
or U17282 (N_17282,N_16687,N_16948);
and U17283 (N_17283,N_16674,N_16621);
nand U17284 (N_17284,N_16838,N_16809);
nor U17285 (N_17285,N_16567,N_16541);
nand U17286 (N_17286,N_16839,N_16725);
and U17287 (N_17287,N_16643,N_16723);
nor U17288 (N_17288,N_16910,N_16729);
and U17289 (N_17289,N_16509,N_16827);
xor U17290 (N_17290,N_16822,N_16669);
nor U17291 (N_17291,N_16663,N_16846);
or U17292 (N_17292,N_16915,N_16919);
or U17293 (N_17293,N_16591,N_16929);
nand U17294 (N_17294,N_16733,N_16555);
or U17295 (N_17295,N_16991,N_16587);
and U17296 (N_17296,N_16939,N_16934);
and U17297 (N_17297,N_16649,N_16950);
nor U17298 (N_17298,N_16811,N_16512);
xor U17299 (N_17299,N_16600,N_16621);
or U17300 (N_17300,N_16711,N_16838);
xnor U17301 (N_17301,N_16753,N_16920);
nand U17302 (N_17302,N_16565,N_16778);
xor U17303 (N_17303,N_16965,N_16688);
nor U17304 (N_17304,N_16568,N_16740);
nor U17305 (N_17305,N_16956,N_16903);
nand U17306 (N_17306,N_16619,N_16534);
nor U17307 (N_17307,N_16850,N_16631);
and U17308 (N_17308,N_16607,N_16589);
and U17309 (N_17309,N_16501,N_16650);
nor U17310 (N_17310,N_16926,N_16881);
nor U17311 (N_17311,N_16939,N_16683);
nor U17312 (N_17312,N_16772,N_16672);
and U17313 (N_17313,N_16991,N_16946);
or U17314 (N_17314,N_16799,N_16694);
nor U17315 (N_17315,N_16921,N_16667);
and U17316 (N_17316,N_16823,N_16513);
or U17317 (N_17317,N_16774,N_16559);
nand U17318 (N_17318,N_16523,N_16673);
xnor U17319 (N_17319,N_16724,N_16625);
nor U17320 (N_17320,N_16795,N_16785);
or U17321 (N_17321,N_16685,N_16552);
or U17322 (N_17322,N_16521,N_16973);
or U17323 (N_17323,N_16982,N_16537);
or U17324 (N_17324,N_16581,N_16546);
xnor U17325 (N_17325,N_16514,N_16747);
nand U17326 (N_17326,N_16916,N_16636);
and U17327 (N_17327,N_16907,N_16510);
nand U17328 (N_17328,N_16729,N_16698);
nor U17329 (N_17329,N_16730,N_16560);
xor U17330 (N_17330,N_16845,N_16549);
nor U17331 (N_17331,N_16550,N_16707);
xor U17332 (N_17332,N_16781,N_16520);
nor U17333 (N_17333,N_16559,N_16860);
or U17334 (N_17334,N_16696,N_16817);
or U17335 (N_17335,N_16595,N_16657);
nor U17336 (N_17336,N_16841,N_16611);
nand U17337 (N_17337,N_16871,N_16776);
xor U17338 (N_17338,N_16884,N_16853);
xor U17339 (N_17339,N_16993,N_16642);
nand U17340 (N_17340,N_16816,N_16892);
or U17341 (N_17341,N_16882,N_16913);
nand U17342 (N_17342,N_16872,N_16964);
nand U17343 (N_17343,N_16938,N_16745);
and U17344 (N_17344,N_16530,N_16550);
or U17345 (N_17345,N_16878,N_16949);
and U17346 (N_17346,N_16581,N_16929);
nand U17347 (N_17347,N_16709,N_16640);
and U17348 (N_17348,N_16918,N_16570);
or U17349 (N_17349,N_16903,N_16848);
nand U17350 (N_17350,N_16605,N_16834);
or U17351 (N_17351,N_16727,N_16853);
nand U17352 (N_17352,N_16929,N_16695);
or U17353 (N_17353,N_16852,N_16794);
and U17354 (N_17354,N_16691,N_16927);
nor U17355 (N_17355,N_16884,N_16861);
xor U17356 (N_17356,N_16525,N_16590);
and U17357 (N_17357,N_16869,N_16682);
nor U17358 (N_17358,N_16699,N_16557);
and U17359 (N_17359,N_16886,N_16780);
xnor U17360 (N_17360,N_16811,N_16863);
nand U17361 (N_17361,N_16899,N_16971);
nor U17362 (N_17362,N_16812,N_16900);
nand U17363 (N_17363,N_16614,N_16739);
nand U17364 (N_17364,N_16719,N_16609);
or U17365 (N_17365,N_16916,N_16583);
and U17366 (N_17366,N_16727,N_16571);
or U17367 (N_17367,N_16547,N_16582);
xor U17368 (N_17368,N_16671,N_16710);
xor U17369 (N_17369,N_16950,N_16639);
nor U17370 (N_17370,N_16518,N_16873);
nor U17371 (N_17371,N_16787,N_16993);
or U17372 (N_17372,N_16550,N_16998);
xnor U17373 (N_17373,N_16608,N_16528);
nor U17374 (N_17374,N_16870,N_16966);
nand U17375 (N_17375,N_16902,N_16760);
xnor U17376 (N_17376,N_16655,N_16966);
and U17377 (N_17377,N_16958,N_16811);
xor U17378 (N_17378,N_16921,N_16717);
nor U17379 (N_17379,N_16896,N_16561);
nor U17380 (N_17380,N_16536,N_16870);
and U17381 (N_17381,N_16781,N_16630);
xor U17382 (N_17382,N_16582,N_16674);
nand U17383 (N_17383,N_16633,N_16729);
or U17384 (N_17384,N_16764,N_16695);
xor U17385 (N_17385,N_16727,N_16903);
and U17386 (N_17386,N_16546,N_16641);
and U17387 (N_17387,N_16765,N_16545);
xnor U17388 (N_17388,N_16567,N_16629);
nor U17389 (N_17389,N_16891,N_16702);
nand U17390 (N_17390,N_16736,N_16763);
nor U17391 (N_17391,N_16877,N_16536);
xor U17392 (N_17392,N_16647,N_16645);
xor U17393 (N_17393,N_16915,N_16579);
nand U17394 (N_17394,N_16737,N_16599);
and U17395 (N_17395,N_16990,N_16948);
xor U17396 (N_17396,N_16661,N_16883);
or U17397 (N_17397,N_16756,N_16528);
nand U17398 (N_17398,N_16687,N_16874);
nor U17399 (N_17399,N_16601,N_16631);
nor U17400 (N_17400,N_16817,N_16675);
nand U17401 (N_17401,N_16975,N_16722);
or U17402 (N_17402,N_16853,N_16540);
nor U17403 (N_17403,N_16768,N_16983);
nand U17404 (N_17404,N_16521,N_16652);
xor U17405 (N_17405,N_16831,N_16969);
nor U17406 (N_17406,N_16714,N_16839);
xnor U17407 (N_17407,N_16612,N_16935);
nand U17408 (N_17408,N_16582,N_16922);
xor U17409 (N_17409,N_16766,N_16612);
and U17410 (N_17410,N_16722,N_16923);
nand U17411 (N_17411,N_16643,N_16955);
xnor U17412 (N_17412,N_16889,N_16682);
xor U17413 (N_17413,N_16758,N_16986);
xor U17414 (N_17414,N_16580,N_16922);
and U17415 (N_17415,N_16602,N_16987);
nand U17416 (N_17416,N_16813,N_16608);
or U17417 (N_17417,N_16804,N_16941);
xor U17418 (N_17418,N_16524,N_16762);
and U17419 (N_17419,N_16671,N_16975);
or U17420 (N_17420,N_16950,N_16724);
and U17421 (N_17421,N_16790,N_16712);
nor U17422 (N_17422,N_16584,N_16981);
nand U17423 (N_17423,N_16766,N_16593);
and U17424 (N_17424,N_16834,N_16940);
or U17425 (N_17425,N_16711,N_16719);
xnor U17426 (N_17426,N_16995,N_16838);
and U17427 (N_17427,N_16671,N_16855);
nor U17428 (N_17428,N_16547,N_16636);
nand U17429 (N_17429,N_16846,N_16722);
nor U17430 (N_17430,N_16936,N_16558);
nor U17431 (N_17431,N_16718,N_16830);
and U17432 (N_17432,N_16956,N_16865);
or U17433 (N_17433,N_16510,N_16987);
xnor U17434 (N_17434,N_16973,N_16847);
and U17435 (N_17435,N_16534,N_16952);
nand U17436 (N_17436,N_16982,N_16703);
xor U17437 (N_17437,N_16971,N_16783);
or U17438 (N_17438,N_16534,N_16665);
or U17439 (N_17439,N_16641,N_16524);
nor U17440 (N_17440,N_16565,N_16793);
and U17441 (N_17441,N_16772,N_16898);
nor U17442 (N_17442,N_16652,N_16667);
xor U17443 (N_17443,N_16822,N_16624);
or U17444 (N_17444,N_16964,N_16755);
and U17445 (N_17445,N_16792,N_16903);
nand U17446 (N_17446,N_16863,N_16909);
and U17447 (N_17447,N_16971,N_16606);
nor U17448 (N_17448,N_16962,N_16569);
xnor U17449 (N_17449,N_16534,N_16546);
xnor U17450 (N_17450,N_16523,N_16883);
nand U17451 (N_17451,N_16504,N_16965);
and U17452 (N_17452,N_16544,N_16946);
or U17453 (N_17453,N_16944,N_16692);
xor U17454 (N_17454,N_16627,N_16786);
nor U17455 (N_17455,N_16941,N_16830);
and U17456 (N_17456,N_16974,N_16790);
nor U17457 (N_17457,N_16727,N_16957);
or U17458 (N_17458,N_16824,N_16702);
xor U17459 (N_17459,N_16865,N_16618);
and U17460 (N_17460,N_16747,N_16746);
nand U17461 (N_17461,N_16938,N_16962);
and U17462 (N_17462,N_16879,N_16548);
and U17463 (N_17463,N_16617,N_16675);
and U17464 (N_17464,N_16973,N_16640);
nand U17465 (N_17465,N_16864,N_16839);
or U17466 (N_17466,N_16806,N_16938);
or U17467 (N_17467,N_16565,N_16965);
and U17468 (N_17468,N_16673,N_16818);
and U17469 (N_17469,N_16597,N_16858);
nand U17470 (N_17470,N_16878,N_16632);
and U17471 (N_17471,N_16877,N_16557);
and U17472 (N_17472,N_16570,N_16887);
nand U17473 (N_17473,N_16677,N_16839);
nand U17474 (N_17474,N_16710,N_16846);
or U17475 (N_17475,N_16505,N_16805);
xor U17476 (N_17476,N_16633,N_16837);
or U17477 (N_17477,N_16602,N_16704);
nand U17478 (N_17478,N_16978,N_16866);
nand U17479 (N_17479,N_16550,N_16979);
and U17480 (N_17480,N_16905,N_16980);
xor U17481 (N_17481,N_16625,N_16714);
nand U17482 (N_17482,N_16868,N_16719);
nand U17483 (N_17483,N_16724,N_16723);
nand U17484 (N_17484,N_16817,N_16853);
nand U17485 (N_17485,N_16598,N_16995);
nand U17486 (N_17486,N_16730,N_16573);
or U17487 (N_17487,N_16697,N_16651);
and U17488 (N_17488,N_16971,N_16524);
and U17489 (N_17489,N_16532,N_16996);
nand U17490 (N_17490,N_16943,N_16515);
xor U17491 (N_17491,N_16817,N_16758);
or U17492 (N_17492,N_16610,N_16848);
and U17493 (N_17493,N_16941,N_16666);
or U17494 (N_17494,N_16556,N_16721);
and U17495 (N_17495,N_16871,N_16585);
xor U17496 (N_17496,N_16769,N_16695);
nand U17497 (N_17497,N_16864,N_16887);
nand U17498 (N_17498,N_16588,N_16940);
or U17499 (N_17499,N_16862,N_16565);
nand U17500 (N_17500,N_17361,N_17342);
and U17501 (N_17501,N_17146,N_17469);
nand U17502 (N_17502,N_17011,N_17344);
nor U17503 (N_17503,N_17213,N_17373);
nand U17504 (N_17504,N_17403,N_17296);
and U17505 (N_17505,N_17042,N_17204);
xnor U17506 (N_17506,N_17396,N_17125);
nand U17507 (N_17507,N_17270,N_17268);
and U17508 (N_17508,N_17447,N_17421);
or U17509 (N_17509,N_17443,N_17168);
xnor U17510 (N_17510,N_17107,N_17050);
and U17511 (N_17511,N_17008,N_17163);
xor U17512 (N_17512,N_17093,N_17110);
xnor U17513 (N_17513,N_17141,N_17427);
or U17514 (N_17514,N_17186,N_17006);
or U17515 (N_17515,N_17206,N_17167);
or U17516 (N_17516,N_17081,N_17232);
and U17517 (N_17517,N_17169,N_17479);
nor U17518 (N_17518,N_17357,N_17193);
and U17519 (N_17519,N_17085,N_17070);
nor U17520 (N_17520,N_17363,N_17105);
nor U17521 (N_17521,N_17264,N_17409);
or U17522 (N_17522,N_17013,N_17377);
and U17523 (N_17523,N_17267,N_17490);
xnor U17524 (N_17524,N_17441,N_17347);
nor U17525 (N_17525,N_17208,N_17283);
nor U17526 (N_17526,N_17462,N_17231);
or U17527 (N_17527,N_17234,N_17442);
and U17528 (N_17528,N_17028,N_17404);
nand U17529 (N_17529,N_17035,N_17248);
nand U17530 (N_17530,N_17030,N_17422);
xor U17531 (N_17531,N_17184,N_17387);
nor U17532 (N_17532,N_17484,N_17384);
and U17533 (N_17533,N_17196,N_17027);
and U17534 (N_17534,N_17108,N_17021);
xnor U17535 (N_17535,N_17436,N_17138);
and U17536 (N_17536,N_17172,N_17197);
nand U17537 (N_17537,N_17118,N_17445);
nand U17538 (N_17538,N_17372,N_17117);
nor U17539 (N_17539,N_17075,N_17148);
or U17540 (N_17540,N_17461,N_17275);
nand U17541 (N_17541,N_17195,N_17339);
xnor U17542 (N_17542,N_17219,N_17240);
or U17543 (N_17543,N_17455,N_17429);
or U17544 (N_17544,N_17348,N_17049);
xnor U17545 (N_17545,N_17124,N_17350);
or U17546 (N_17546,N_17474,N_17122);
or U17547 (N_17547,N_17487,N_17016);
and U17548 (N_17548,N_17097,N_17279);
xor U17549 (N_17549,N_17173,N_17135);
and U17550 (N_17550,N_17327,N_17091);
and U17551 (N_17551,N_17368,N_17489);
nand U17552 (N_17552,N_17210,N_17079);
nand U17553 (N_17553,N_17343,N_17177);
nand U17554 (N_17554,N_17094,N_17493);
nand U17555 (N_17555,N_17480,N_17115);
nand U17556 (N_17556,N_17444,N_17098);
nand U17557 (N_17557,N_17380,N_17077);
nor U17558 (N_17558,N_17376,N_17180);
nor U17559 (N_17559,N_17149,N_17375);
nor U17560 (N_17560,N_17395,N_17096);
or U17561 (N_17561,N_17014,N_17058);
or U17562 (N_17562,N_17294,N_17494);
nand U17563 (N_17563,N_17450,N_17237);
or U17564 (N_17564,N_17040,N_17015);
and U17565 (N_17565,N_17379,N_17066);
nor U17566 (N_17566,N_17465,N_17316);
nor U17567 (N_17567,N_17383,N_17134);
nand U17568 (N_17568,N_17295,N_17106);
nor U17569 (N_17569,N_17308,N_17119);
and U17570 (N_17570,N_17127,N_17470);
nand U17571 (N_17571,N_17452,N_17340);
nor U17572 (N_17572,N_17290,N_17235);
xor U17573 (N_17573,N_17052,N_17496);
nand U17574 (N_17574,N_17223,N_17055);
or U17575 (N_17575,N_17202,N_17416);
nor U17576 (N_17576,N_17492,N_17498);
nor U17577 (N_17577,N_17104,N_17408);
xor U17578 (N_17578,N_17349,N_17394);
or U17579 (N_17579,N_17174,N_17183);
and U17580 (N_17580,N_17491,N_17103);
and U17581 (N_17581,N_17087,N_17284);
xor U17582 (N_17582,N_17229,N_17392);
and U17583 (N_17583,N_17386,N_17060);
and U17584 (N_17584,N_17150,N_17246);
xor U17585 (N_17585,N_17381,N_17164);
or U17586 (N_17586,N_17269,N_17354);
or U17587 (N_17587,N_17225,N_17092);
xnor U17588 (N_17588,N_17337,N_17084);
xnor U17589 (N_17589,N_17009,N_17100);
xor U17590 (N_17590,N_17448,N_17265);
xnor U17591 (N_17591,N_17488,N_17266);
or U17592 (N_17592,N_17113,N_17326);
or U17593 (N_17593,N_17139,N_17360);
and U17594 (N_17594,N_17407,N_17324);
or U17595 (N_17595,N_17261,N_17282);
nand U17596 (N_17596,N_17067,N_17185);
or U17597 (N_17597,N_17182,N_17086);
and U17598 (N_17598,N_17038,N_17018);
and U17599 (N_17599,N_17147,N_17227);
or U17600 (N_17600,N_17259,N_17287);
or U17601 (N_17601,N_17311,N_17307);
and U17602 (N_17602,N_17002,N_17258);
nor U17603 (N_17603,N_17362,N_17318);
nand U17604 (N_17604,N_17226,N_17424);
xnor U17605 (N_17605,N_17102,N_17338);
nand U17606 (N_17606,N_17260,N_17305);
nor U17607 (N_17607,N_17400,N_17143);
and U17608 (N_17608,N_17000,N_17082);
and U17609 (N_17609,N_17170,N_17405);
or U17610 (N_17610,N_17026,N_17224);
or U17611 (N_17611,N_17053,N_17476);
nor U17612 (N_17612,N_17198,N_17262);
nor U17613 (N_17613,N_17459,N_17365);
nor U17614 (N_17614,N_17353,N_17005);
or U17615 (N_17615,N_17370,N_17056);
xnor U17616 (N_17616,N_17298,N_17304);
and U17617 (N_17617,N_17333,N_17426);
xor U17618 (N_17618,N_17121,N_17310);
nor U17619 (N_17619,N_17222,N_17043);
nor U17620 (N_17620,N_17364,N_17406);
nor U17621 (N_17621,N_17414,N_17257);
or U17622 (N_17622,N_17057,N_17128);
or U17623 (N_17623,N_17288,N_17359);
or U17624 (N_17624,N_17473,N_17194);
and U17625 (N_17625,N_17130,N_17073);
nand U17626 (N_17626,N_17382,N_17320);
or U17627 (N_17627,N_17080,N_17238);
or U17628 (N_17628,N_17061,N_17137);
xor U17629 (N_17629,N_17303,N_17317);
nand U17630 (N_17630,N_17458,N_17366);
xnor U17631 (N_17631,N_17482,N_17218);
xor U17632 (N_17632,N_17034,N_17142);
xnor U17633 (N_17633,N_17435,N_17328);
and U17634 (N_17634,N_17254,N_17044);
or U17635 (N_17635,N_17214,N_17495);
and U17636 (N_17636,N_17432,N_17242);
or U17637 (N_17637,N_17412,N_17292);
nor U17638 (N_17638,N_17249,N_17312);
or U17639 (N_17639,N_17151,N_17123);
or U17640 (N_17640,N_17335,N_17062);
or U17641 (N_17641,N_17176,N_17033);
xor U17642 (N_17642,N_17145,N_17059);
and U17643 (N_17643,N_17341,N_17356);
or U17644 (N_17644,N_17191,N_17181);
xnor U17645 (N_17645,N_17095,N_17160);
or U17646 (N_17646,N_17215,N_17256);
or U17647 (N_17647,N_17300,N_17355);
xnor U17648 (N_17648,N_17467,N_17020);
xor U17649 (N_17649,N_17263,N_17369);
nand U17650 (N_17650,N_17276,N_17090);
xor U17651 (N_17651,N_17289,N_17003);
or U17652 (N_17652,N_17393,N_17385);
or U17653 (N_17653,N_17212,N_17297);
xnor U17654 (N_17654,N_17468,N_17063);
and U17655 (N_17655,N_17031,N_17449);
nand U17656 (N_17656,N_17454,N_17321);
xor U17657 (N_17657,N_17047,N_17140);
or U17658 (N_17658,N_17293,N_17331);
nand U17659 (N_17659,N_17425,N_17345);
or U17660 (N_17660,N_17131,N_17065);
xnor U17661 (N_17661,N_17132,N_17434);
nor U17662 (N_17662,N_17486,N_17078);
nor U17663 (N_17663,N_17358,N_17483);
and U17664 (N_17664,N_17313,N_17023);
and U17665 (N_17665,N_17398,N_17439);
and U17666 (N_17666,N_17374,N_17319);
or U17667 (N_17667,N_17045,N_17054);
nand U17668 (N_17668,N_17253,N_17126);
and U17669 (N_17669,N_17192,N_17475);
xor U17670 (N_17670,N_17472,N_17413);
xnor U17671 (N_17671,N_17207,N_17154);
nor U17672 (N_17672,N_17463,N_17336);
nand U17673 (N_17673,N_17155,N_17162);
or U17674 (N_17674,N_17064,N_17478);
and U17675 (N_17675,N_17460,N_17099);
nand U17676 (N_17676,N_17109,N_17280);
xnor U17677 (N_17677,N_17175,N_17046);
nor U17678 (N_17678,N_17152,N_17423);
and U17679 (N_17679,N_17101,N_17378);
nand U17680 (N_17680,N_17271,N_17171);
nand U17681 (N_17681,N_17007,N_17402);
and U17682 (N_17682,N_17178,N_17440);
nor U17683 (N_17683,N_17438,N_17323);
and U17684 (N_17684,N_17243,N_17471);
and U17685 (N_17685,N_17004,N_17088);
nor U17686 (N_17686,N_17166,N_17071);
xor U17687 (N_17687,N_17286,N_17114);
nor U17688 (N_17688,N_17431,N_17221);
and U17689 (N_17689,N_17241,N_17159);
nand U17690 (N_17690,N_17211,N_17189);
or U17691 (N_17691,N_17325,N_17179);
and U17692 (N_17692,N_17437,N_17401);
or U17693 (N_17693,N_17209,N_17329);
xnor U17694 (N_17694,N_17112,N_17203);
or U17695 (N_17695,N_17036,N_17217);
and U17696 (N_17696,N_17281,N_17291);
nand U17697 (N_17697,N_17161,N_17228);
and U17698 (N_17698,N_17301,N_17165);
nand U17699 (N_17699,N_17251,N_17322);
xnor U17700 (N_17700,N_17144,N_17239);
nand U17701 (N_17701,N_17083,N_17278);
xnor U17702 (N_17702,N_17074,N_17187);
xnor U17703 (N_17703,N_17451,N_17272);
nor U17704 (N_17704,N_17111,N_17024);
nor U17705 (N_17705,N_17285,N_17309);
nor U17706 (N_17706,N_17076,N_17156);
nor U17707 (N_17707,N_17453,N_17497);
nor U17708 (N_17708,N_17029,N_17157);
and U17709 (N_17709,N_17245,N_17068);
xnor U17710 (N_17710,N_17205,N_17273);
nor U17711 (N_17711,N_17220,N_17190);
and U17712 (N_17712,N_17201,N_17477);
xor U17713 (N_17713,N_17200,N_17017);
nand U17714 (N_17714,N_17299,N_17464);
or U17715 (N_17715,N_17371,N_17199);
nand U17716 (N_17716,N_17032,N_17446);
nand U17717 (N_17717,N_17352,N_17315);
xnor U17718 (N_17718,N_17420,N_17069);
or U17719 (N_17719,N_17158,N_17019);
or U17720 (N_17720,N_17153,N_17012);
and U17721 (N_17721,N_17390,N_17332);
or U17722 (N_17722,N_17255,N_17419);
or U17723 (N_17723,N_17418,N_17417);
nor U17724 (N_17724,N_17216,N_17428);
xnor U17725 (N_17725,N_17025,N_17430);
xor U17726 (N_17726,N_17410,N_17399);
xnor U17727 (N_17727,N_17129,N_17397);
xnor U17728 (N_17728,N_17230,N_17274);
nand U17729 (N_17729,N_17136,N_17233);
or U17730 (N_17730,N_17072,N_17120);
and U17731 (N_17731,N_17250,N_17277);
and U17732 (N_17732,N_17039,N_17306);
xnor U17733 (N_17733,N_17456,N_17411);
nand U17734 (N_17734,N_17302,N_17367);
and U17735 (N_17735,N_17481,N_17391);
nand U17736 (N_17736,N_17499,N_17022);
and U17737 (N_17737,N_17334,N_17433);
or U17738 (N_17738,N_17244,N_17116);
or U17739 (N_17739,N_17252,N_17389);
and U17740 (N_17740,N_17314,N_17133);
and U17741 (N_17741,N_17188,N_17010);
and U17742 (N_17742,N_17330,N_17485);
nand U17743 (N_17743,N_17415,N_17048);
or U17744 (N_17744,N_17041,N_17346);
nand U17745 (N_17745,N_17247,N_17001);
xor U17746 (N_17746,N_17051,N_17236);
nor U17747 (N_17747,N_17466,N_17351);
nand U17748 (N_17748,N_17037,N_17089);
or U17749 (N_17749,N_17388,N_17457);
nand U17750 (N_17750,N_17086,N_17254);
and U17751 (N_17751,N_17471,N_17138);
and U17752 (N_17752,N_17124,N_17276);
or U17753 (N_17753,N_17317,N_17221);
nor U17754 (N_17754,N_17269,N_17090);
nor U17755 (N_17755,N_17298,N_17161);
xor U17756 (N_17756,N_17016,N_17258);
nor U17757 (N_17757,N_17303,N_17134);
and U17758 (N_17758,N_17218,N_17411);
nor U17759 (N_17759,N_17313,N_17413);
nand U17760 (N_17760,N_17090,N_17275);
or U17761 (N_17761,N_17235,N_17314);
or U17762 (N_17762,N_17465,N_17496);
nand U17763 (N_17763,N_17068,N_17256);
xor U17764 (N_17764,N_17259,N_17193);
nand U17765 (N_17765,N_17206,N_17459);
nor U17766 (N_17766,N_17375,N_17282);
xor U17767 (N_17767,N_17291,N_17020);
nand U17768 (N_17768,N_17298,N_17301);
nor U17769 (N_17769,N_17357,N_17429);
nand U17770 (N_17770,N_17047,N_17120);
or U17771 (N_17771,N_17083,N_17207);
or U17772 (N_17772,N_17015,N_17072);
or U17773 (N_17773,N_17399,N_17429);
xnor U17774 (N_17774,N_17071,N_17237);
nand U17775 (N_17775,N_17452,N_17158);
or U17776 (N_17776,N_17350,N_17017);
nor U17777 (N_17777,N_17046,N_17060);
and U17778 (N_17778,N_17427,N_17154);
nand U17779 (N_17779,N_17480,N_17284);
or U17780 (N_17780,N_17102,N_17167);
nand U17781 (N_17781,N_17396,N_17155);
and U17782 (N_17782,N_17016,N_17456);
and U17783 (N_17783,N_17151,N_17248);
xnor U17784 (N_17784,N_17434,N_17464);
nor U17785 (N_17785,N_17240,N_17165);
and U17786 (N_17786,N_17467,N_17314);
or U17787 (N_17787,N_17088,N_17470);
and U17788 (N_17788,N_17014,N_17304);
xor U17789 (N_17789,N_17047,N_17229);
or U17790 (N_17790,N_17061,N_17029);
nor U17791 (N_17791,N_17203,N_17173);
nor U17792 (N_17792,N_17165,N_17387);
xor U17793 (N_17793,N_17470,N_17107);
and U17794 (N_17794,N_17349,N_17443);
and U17795 (N_17795,N_17211,N_17132);
or U17796 (N_17796,N_17326,N_17390);
nand U17797 (N_17797,N_17427,N_17323);
or U17798 (N_17798,N_17418,N_17390);
xor U17799 (N_17799,N_17137,N_17275);
or U17800 (N_17800,N_17220,N_17491);
nand U17801 (N_17801,N_17290,N_17260);
nor U17802 (N_17802,N_17428,N_17066);
nand U17803 (N_17803,N_17488,N_17130);
xnor U17804 (N_17804,N_17111,N_17240);
nor U17805 (N_17805,N_17149,N_17257);
or U17806 (N_17806,N_17372,N_17026);
or U17807 (N_17807,N_17082,N_17264);
nand U17808 (N_17808,N_17110,N_17205);
xnor U17809 (N_17809,N_17257,N_17366);
xor U17810 (N_17810,N_17005,N_17171);
nor U17811 (N_17811,N_17206,N_17193);
nand U17812 (N_17812,N_17384,N_17458);
nand U17813 (N_17813,N_17371,N_17127);
xor U17814 (N_17814,N_17228,N_17058);
and U17815 (N_17815,N_17418,N_17402);
nor U17816 (N_17816,N_17186,N_17064);
xnor U17817 (N_17817,N_17082,N_17072);
nand U17818 (N_17818,N_17159,N_17461);
nand U17819 (N_17819,N_17212,N_17470);
xor U17820 (N_17820,N_17421,N_17116);
or U17821 (N_17821,N_17324,N_17347);
xor U17822 (N_17822,N_17047,N_17356);
xnor U17823 (N_17823,N_17088,N_17412);
or U17824 (N_17824,N_17082,N_17488);
xnor U17825 (N_17825,N_17202,N_17138);
xor U17826 (N_17826,N_17224,N_17198);
xnor U17827 (N_17827,N_17251,N_17465);
nor U17828 (N_17828,N_17049,N_17147);
or U17829 (N_17829,N_17048,N_17218);
and U17830 (N_17830,N_17224,N_17434);
xor U17831 (N_17831,N_17370,N_17446);
and U17832 (N_17832,N_17156,N_17240);
and U17833 (N_17833,N_17324,N_17072);
and U17834 (N_17834,N_17418,N_17467);
xor U17835 (N_17835,N_17317,N_17368);
nor U17836 (N_17836,N_17278,N_17320);
nand U17837 (N_17837,N_17088,N_17400);
nand U17838 (N_17838,N_17169,N_17340);
and U17839 (N_17839,N_17492,N_17496);
or U17840 (N_17840,N_17235,N_17013);
nand U17841 (N_17841,N_17379,N_17294);
or U17842 (N_17842,N_17413,N_17323);
nor U17843 (N_17843,N_17379,N_17012);
nand U17844 (N_17844,N_17251,N_17342);
nand U17845 (N_17845,N_17235,N_17379);
and U17846 (N_17846,N_17312,N_17397);
or U17847 (N_17847,N_17264,N_17048);
or U17848 (N_17848,N_17031,N_17248);
xor U17849 (N_17849,N_17096,N_17110);
and U17850 (N_17850,N_17240,N_17057);
and U17851 (N_17851,N_17212,N_17291);
nor U17852 (N_17852,N_17248,N_17026);
xor U17853 (N_17853,N_17384,N_17173);
or U17854 (N_17854,N_17451,N_17300);
nor U17855 (N_17855,N_17052,N_17481);
xnor U17856 (N_17856,N_17096,N_17251);
nor U17857 (N_17857,N_17373,N_17090);
nand U17858 (N_17858,N_17237,N_17370);
or U17859 (N_17859,N_17212,N_17083);
xnor U17860 (N_17860,N_17240,N_17438);
xor U17861 (N_17861,N_17110,N_17168);
xnor U17862 (N_17862,N_17293,N_17241);
xnor U17863 (N_17863,N_17174,N_17105);
nand U17864 (N_17864,N_17115,N_17259);
or U17865 (N_17865,N_17146,N_17066);
nand U17866 (N_17866,N_17138,N_17220);
or U17867 (N_17867,N_17239,N_17067);
and U17868 (N_17868,N_17497,N_17226);
nand U17869 (N_17869,N_17276,N_17065);
nand U17870 (N_17870,N_17138,N_17036);
and U17871 (N_17871,N_17319,N_17035);
or U17872 (N_17872,N_17011,N_17390);
or U17873 (N_17873,N_17419,N_17231);
nand U17874 (N_17874,N_17034,N_17192);
xor U17875 (N_17875,N_17375,N_17015);
xor U17876 (N_17876,N_17016,N_17203);
and U17877 (N_17877,N_17332,N_17011);
or U17878 (N_17878,N_17364,N_17449);
or U17879 (N_17879,N_17267,N_17258);
or U17880 (N_17880,N_17207,N_17110);
nor U17881 (N_17881,N_17006,N_17177);
nor U17882 (N_17882,N_17474,N_17405);
and U17883 (N_17883,N_17185,N_17366);
and U17884 (N_17884,N_17217,N_17178);
or U17885 (N_17885,N_17015,N_17120);
and U17886 (N_17886,N_17234,N_17356);
nor U17887 (N_17887,N_17132,N_17103);
xor U17888 (N_17888,N_17028,N_17346);
xnor U17889 (N_17889,N_17097,N_17358);
nor U17890 (N_17890,N_17268,N_17308);
nor U17891 (N_17891,N_17080,N_17160);
or U17892 (N_17892,N_17383,N_17155);
or U17893 (N_17893,N_17332,N_17371);
xor U17894 (N_17894,N_17447,N_17360);
nand U17895 (N_17895,N_17428,N_17292);
xor U17896 (N_17896,N_17021,N_17113);
nand U17897 (N_17897,N_17212,N_17228);
nand U17898 (N_17898,N_17415,N_17309);
or U17899 (N_17899,N_17205,N_17086);
nor U17900 (N_17900,N_17148,N_17067);
xor U17901 (N_17901,N_17341,N_17384);
nand U17902 (N_17902,N_17413,N_17026);
nand U17903 (N_17903,N_17064,N_17062);
or U17904 (N_17904,N_17322,N_17249);
or U17905 (N_17905,N_17356,N_17174);
nand U17906 (N_17906,N_17387,N_17002);
or U17907 (N_17907,N_17248,N_17034);
xor U17908 (N_17908,N_17409,N_17229);
nor U17909 (N_17909,N_17146,N_17474);
nand U17910 (N_17910,N_17463,N_17071);
nor U17911 (N_17911,N_17375,N_17299);
nor U17912 (N_17912,N_17070,N_17117);
or U17913 (N_17913,N_17097,N_17017);
and U17914 (N_17914,N_17141,N_17434);
nand U17915 (N_17915,N_17417,N_17488);
and U17916 (N_17916,N_17202,N_17387);
nand U17917 (N_17917,N_17289,N_17161);
nor U17918 (N_17918,N_17005,N_17337);
nand U17919 (N_17919,N_17161,N_17333);
and U17920 (N_17920,N_17315,N_17222);
and U17921 (N_17921,N_17048,N_17397);
or U17922 (N_17922,N_17412,N_17455);
or U17923 (N_17923,N_17165,N_17340);
xor U17924 (N_17924,N_17086,N_17400);
and U17925 (N_17925,N_17151,N_17051);
xnor U17926 (N_17926,N_17295,N_17239);
nor U17927 (N_17927,N_17134,N_17399);
and U17928 (N_17928,N_17370,N_17203);
and U17929 (N_17929,N_17118,N_17099);
xor U17930 (N_17930,N_17285,N_17310);
nor U17931 (N_17931,N_17042,N_17302);
and U17932 (N_17932,N_17476,N_17355);
nor U17933 (N_17933,N_17063,N_17374);
nor U17934 (N_17934,N_17449,N_17236);
and U17935 (N_17935,N_17495,N_17177);
xnor U17936 (N_17936,N_17266,N_17007);
nor U17937 (N_17937,N_17250,N_17175);
xnor U17938 (N_17938,N_17091,N_17041);
nand U17939 (N_17939,N_17210,N_17393);
or U17940 (N_17940,N_17495,N_17096);
and U17941 (N_17941,N_17115,N_17151);
nor U17942 (N_17942,N_17128,N_17422);
or U17943 (N_17943,N_17191,N_17211);
nor U17944 (N_17944,N_17108,N_17420);
nor U17945 (N_17945,N_17377,N_17367);
xor U17946 (N_17946,N_17062,N_17249);
and U17947 (N_17947,N_17407,N_17288);
nand U17948 (N_17948,N_17094,N_17455);
nand U17949 (N_17949,N_17265,N_17363);
and U17950 (N_17950,N_17017,N_17383);
xnor U17951 (N_17951,N_17096,N_17485);
and U17952 (N_17952,N_17442,N_17246);
and U17953 (N_17953,N_17200,N_17225);
or U17954 (N_17954,N_17360,N_17064);
and U17955 (N_17955,N_17453,N_17431);
nor U17956 (N_17956,N_17419,N_17456);
xor U17957 (N_17957,N_17273,N_17434);
nor U17958 (N_17958,N_17317,N_17417);
nand U17959 (N_17959,N_17469,N_17436);
nand U17960 (N_17960,N_17010,N_17007);
nor U17961 (N_17961,N_17116,N_17140);
and U17962 (N_17962,N_17203,N_17334);
and U17963 (N_17963,N_17197,N_17151);
xnor U17964 (N_17964,N_17310,N_17194);
nor U17965 (N_17965,N_17061,N_17362);
or U17966 (N_17966,N_17163,N_17105);
or U17967 (N_17967,N_17104,N_17397);
or U17968 (N_17968,N_17261,N_17328);
nor U17969 (N_17969,N_17297,N_17112);
nand U17970 (N_17970,N_17141,N_17263);
xor U17971 (N_17971,N_17325,N_17446);
xnor U17972 (N_17972,N_17032,N_17041);
nor U17973 (N_17973,N_17345,N_17327);
nand U17974 (N_17974,N_17003,N_17359);
xnor U17975 (N_17975,N_17373,N_17378);
or U17976 (N_17976,N_17316,N_17153);
or U17977 (N_17977,N_17180,N_17019);
nand U17978 (N_17978,N_17247,N_17212);
nand U17979 (N_17979,N_17385,N_17262);
or U17980 (N_17980,N_17061,N_17246);
nand U17981 (N_17981,N_17364,N_17254);
or U17982 (N_17982,N_17273,N_17427);
nor U17983 (N_17983,N_17051,N_17475);
and U17984 (N_17984,N_17263,N_17486);
xor U17985 (N_17985,N_17230,N_17314);
and U17986 (N_17986,N_17060,N_17127);
or U17987 (N_17987,N_17397,N_17255);
nand U17988 (N_17988,N_17132,N_17026);
or U17989 (N_17989,N_17020,N_17058);
xnor U17990 (N_17990,N_17440,N_17156);
nor U17991 (N_17991,N_17447,N_17340);
nor U17992 (N_17992,N_17058,N_17494);
nand U17993 (N_17993,N_17450,N_17031);
or U17994 (N_17994,N_17151,N_17011);
and U17995 (N_17995,N_17361,N_17444);
or U17996 (N_17996,N_17491,N_17146);
and U17997 (N_17997,N_17284,N_17214);
nor U17998 (N_17998,N_17450,N_17177);
xnor U17999 (N_17999,N_17217,N_17133);
nand U18000 (N_18000,N_17699,N_17527);
and U18001 (N_18001,N_17783,N_17873);
xor U18002 (N_18002,N_17704,N_17762);
and U18003 (N_18003,N_17551,N_17809);
xnor U18004 (N_18004,N_17858,N_17883);
or U18005 (N_18005,N_17823,N_17707);
nand U18006 (N_18006,N_17628,N_17942);
nand U18007 (N_18007,N_17564,N_17925);
and U18008 (N_18008,N_17961,N_17518);
or U18009 (N_18009,N_17879,N_17862);
and U18010 (N_18010,N_17607,N_17801);
and U18011 (N_18011,N_17740,N_17738);
or U18012 (N_18012,N_17582,N_17763);
xor U18013 (N_18013,N_17833,N_17843);
and U18014 (N_18014,N_17675,N_17727);
and U18015 (N_18015,N_17659,N_17872);
xor U18016 (N_18016,N_17665,N_17746);
and U18017 (N_18017,N_17674,N_17737);
and U18018 (N_18018,N_17671,N_17932);
nor U18019 (N_18019,N_17702,N_17871);
or U18020 (N_18020,N_17690,N_17832);
nor U18021 (N_18021,N_17970,N_17557);
xor U18022 (N_18022,N_17595,N_17505);
or U18023 (N_18023,N_17621,N_17850);
and U18024 (N_18024,N_17842,N_17549);
nor U18025 (N_18025,N_17692,N_17771);
nor U18026 (N_18026,N_17951,N_17870);
or U18027 (N_18027,N_17515,N_17927);
and U18028 (N_18028,N_17941,N_17859);
nor U18029 (N_18029,N_17955,N_17693);
nand U18030 (N_18030,N_17953,N_17876);
nor U18031 (N_18031,N_17547,N_17614);
xnor U18032 (N_18032,N_17922,N_17851);
nand U18033 (N_18033,N_17626,N_17752);
xnor U18034 (N_18034,N_17720,N_17980);
or U18035 (N_18035,N_17630,N_17610);
or U18036 (N_18036,N_17652,N_17716);
nand U18037 (N_18037,N_17543,N_17601);
and U18038 (N_18038,N_17897,N_17660);
xor U18039 (N_18039,N_17683,N_17532);
nor U18040 (N_18040,N_17896,N_17962);
and U18041 (N_18041,N_17826,N_17578);
and U18042 (N_18042,N_17797,N_17540);
nand U18043 (N_18043,N_17829,N_17593);
nor U18044 (N_18044,N_17960,N_17910);
or U18045 (N_18045,N_17625,N_17535);
or U18046 (N_18046,N_17957,N_17567);
and U18047 (N_18047,N_17638,N_17988);
and U18048 (N_18048,N_17937,N_17744);
or U18049 (N_18049,N_17755,N_17701);
nor U18050 (N_18050,N_17722,N_17511);
nand U18051 (N_18051,N_17887,N_17725);
or U18052 (N_18052,N_17987,N_17906);
xnor U18053 (N_18053,N_17637,N_17944);
nor U18054 (N_18054,N_17780,N_17706);
and U18055 (N_18055,N_17898,N_17939);
and U18056 (N_18056,N_17633,N_17837);
or U18057 (N_18057,N_17748,N_17766);
xor U18058 (N_18058,N_17928,N_17577);
or U18059 (N_18059,N_17516,N_17571);
or U18060 (N_18060,N_17513,N_17676);
or U18061 (N_18061,N_17803,N_17892);
nand U18062 (N_18062,N_17849,N_17793);
nand U18063 (N_18063,N_17632,N_17764);
nand U18064 (N_18064,N_17997,N_17992);
xnor U18065 (N_18065,N_17563,N_17681);
or U18066 (N_18066,N_17990,N_17995);
nor U18067 (N_18067,N_17865,N_17560);
nand U18068 (N_18068,N_17684,N_17787);
nand U18069 (N_18069,N_17597,N_17613);
nor U18070 (N_18070,N_17768,N_17821);
and U18071 (N_18071,N_17945,N_17617);
or U18072 (N_18072,N_17680,N_17856);
nand U18073 (N_18073,N_17657,N_17594);
xnor U18074 (N_18074,N_17973,N_17841);
nor U18075 (N_18075,N_17971,N_17667);
xnor U18076 (N_18076,N_17888,N_17544);
nor U18077 (N_18077,N_17866,N_17539);
nand U18078 (N_18078,N_17817,N_17524);
nor U18079 (N_18079,N_17718,N_17743);
xor U18080 (N_18080,N_17635,N_17974);
xnor U18081 (N_18081,N_17816,N_17574);
and U18082 (N_18082,N_17736,N_17982);
nor U18083 (N_18083,N_17696,N_17636);
and U18084 (N_18084,N_17760,N_17891);
xor U18085 (N_18085,N_17519,N_17885);
nor U18086 (N_18086,N_17972,N_17919);
nand U18087 (N_18087,N_17650,N_17869);
xor U18088 (N_18088,N_17996,N_17967);
nor U18089 (N_18089,N_17559,N_17724);
xnor U18090 (N_18090,N_17770,N_17658);
xnor U18091 (N_18091,N_17598,N_17948);
and U18092 (N_18092,N_17900,N_17890);
nand U18093 (N_18093,N_17662,N_17506);
and U18094 (N_18094,N_17978,N_17773);
nor U18095 (N_18095,N_17620,N_17983);
xor U18096 (N_18096,N_17750,N_17694);
and U18097 (N_18097,N_17857,N_17558);
xnor U18098 (N_18098,N_17759,N_17989);
xor U18099 (N_18099,N_17586,N_17827);
nor U18100 (N_18100,N_17572,N_17705);
and U18101 (N_18101,N_17986,N_17999);
and U18102 (N_18102,N_17703,N_17673);
or U18103 (N_18103,N_17569,N_17968);
nor U18104 (N_18104,N_17708,N_17952);
xnor U18105 (N_18105,N_17646,N_17729);
nand U18106 (N_18106,N_17943,N_17845);
xor U18107 (N_18107,N_17711,N_17808);
or U18108 (N_18108,N_17709,N_17730);
xnor U18109 (N_18109,N_17861,N_17698);
or U18110 (N_18110,N_17509,N_17534);
nand U18111 (N_18111,N_17503,N_17697);
nor U18112 (N_18112,N_17774,N_17938);
and U18113 (N_18113,N_17921,N_17507);
xor U18114 (N_18114,N_17687,N_17695);
xor U18115 (N_18115,N_17618,N_17964);
nor U18116 (N_18116,N_17615,N_17649);
or U18117 (N_18117,N_17745,N_17741);
nor U18118 (N_18118,N_17612,N_17596);
nor U18119 (N_18119,N_17965,N_17807);
nor U18120 (N_18120,N_17875,N_17689);
nand U18121 (N_18121,N_17517,N_17556);
and U18122 (N_18122,N_17915,N_17828);
xor U18123 (N_18123,N_17723,N_17624);
nor U18124 (N_18124,N_17895,N_17510);
nand U18125 (N_18125,N_17604,N_17909);
and U18126 (N_18126,N_17786,N_17717);
xnor U18127 (N_18127,N_17512,N_17565);
nor U18128 (N_18128,N_17605,N_17806);
xor U18129 (N_18129,N_17846,N_17661);
nor U18130 (N_18130,N_17712,N_17640);
xnor U18131 (N_18131,N_17568,N_17530);
and U18132 (N_18132,N_17931,N_17575);
and U18133 (N_18133,N_17670,N_17504);
xnor U18134 (N_18134,N_17644,N_17799);
nor U18135 (N_18135,N_17886,N_17867);
and U18136 (N_18136,N_17813,N_17611);
xnor U18137 (N_18137,N_17985,N_17528);
nand U18138 (N_18138,N_17522,N_17753);
and U18139 (N_18139,N_17781,N_17566);
xnor U18140 (N_18140,N_17669,N_17977);
and U18141 (N_18141,N_17769,N_17576);
or U18142 (N_18142,N_17863,N_17903);
or U18143 (N_18143,N_17820,N_17685);
xor U18144 (N_18144,N_17798,N_17538);
or U18145 (N_18145,N_17838,N_17726);
nor U18146 (N_18146,N_17788,N_17682);
xor U18147 (N_18147,N_17553,N_17579);
nor U18148 (N_18148,N_17648,N_17501);
nor U18149 (N_18149,N_17719,N_17508);
or U18150 (N_18150,N_17656,N_17877);
xor U18151 (N_18151,N_17691,N_17592);
nand U18152 (N_18152,N_17537,N_17639);
nand U18153 (N_18153,N_17548,N_17839);
or U18154 (N_18154,N_17880,N_17914);
or U18155 (N_18155,N_17562,N_17778);
and U18156 (N_18156,N_17642,N_17765);
or U18157 (N_18157,N_17521,N_17946);
or U18158 (N_18158,N_17502,N_17934);
nor U18159 (N_18159,N_17795,N_17555);
nand U18160 (N_18160,N_17761,N_17785);
nand U18161 (N_18161,N_17643,N_17523);
nand U18162 (N_18162,N_17590,N_17550);
or U18163 (N_18163,N_17664,N_17836);
xnor U18164 (N_18164,N_17647,N_17917);
and U18165 (N_18165,N_17984,N_17956);
or U18166 (N_18166,N_17603,N_17732);
and U18167 (N_18167,N_17790,N_17700);
nand U18168 (N_18168,N_17822,N_17860);
xor U18169 (N_18169,N_17735,N_17882);
or U18170 (N_18170,N_17926,N_17533);
nand U18171 (N_18171,N_17713,N_17772);
xnor U18172 (N_18172,N_17580,N_17855);
nor U18173 (N_18173,N_17591,N_17634);
and U18174 (N_18174,N_17901,N_17679);
nand U18175 (N_18175,N_17784,N_17733);
nand U18176 (N_18176,N_17545,N_17546);
and U18177 (N_18177,N_17654,N_17606);
xor U18178 (N_18178,N_17905,N_17645);
nor U18179 (N_18179,N_17777,N_17998);
nor U18180 (N_18180,N_17840,N_17570);
nand U18181 (N_18181,N_17520,N_17969);
or U18182 (N_18182,N_17554,N_17758);
xor U18183 (N_18183,N_17963,N_17923);
xor U18184 (N_18184,N_17852,N_17918);
nand U18185 (N_18185,N_17854,N_17608);
or U18186 (N_18186,N_17811,N_17573);
and U18187 (N_18187,N_17976,N_17710);
nor U18188 (N_18188,N_17631,N_17810);
and U18189 (N_18189,N_17831,N_17889);
nor U18190 (N_18190,N_17749,N_17616);
nand U18191 (N_18191,N_17653,N_17904);
nand U18192 (N_18192,N_17847,N_17714);
nor U18193 (N_18193,N_17715,N_17800);
or U18194 (N_18194,N_17791,N_17756);
nand U18195 (N_18195,N_17979,N_17668);
and U18196 (N_18196,N_17819,N_17531);
nand U18197 (N_18197,N_17666,N_17627);
nor U18198 (N_18198,N_17583,N_17881);
and U18199 (N_18199,N_17599,N_17677);
and U18200 (N_18200,N_17864,N_17913);
nand U18201 (N_18201,N_17526,N_17975);
nor U18202 (N_18202,N_17581,N_17686);
nor U18203 (N_18203,N_17950,N_17966);
xnor U18204 (N_18204,N_17920,N_17525);
nand U18205 (N_18205,N_17802,N_17622);
or U18206 (N_18206,N_17994,N_17907);
and U18207 (N_18207,N_17924,N_17815);
or U18208 (N_18208,N_17751,N_17757);
or U18209 (N_18209,N_17782,N_17893);
nor U18210 (N_18210,N_17911,N_17552);
nor U18211 (N_18211,N_17629,N_17804);
or U18212 (N_18212,N_17912,N_17993);
and U18213 (N_18213,N_17902,N_17792);
nand U18214 (N_18214,N_17940,N_17655);
xnor U18215 (N_18215,N_17619,N_17542);
nor U18216 (N_18216,N_17954,N_17651);
and U18217 (N_18217,N_17796,N_17514);
nor U18218 (N_18218,N_17830,N_17868);
and U18219 (N_18219,N_17600,N_17739);
or U18220 (N_18220,N_17825,N_17541);
xnor U18221 (N_18221,N_17754,N_17587);
or U18222 (N_18222,N_17609,N_17688);
xor U18223 (N_18223,N_17731,N_17589);
xnor U18224 (N_18224,N_17958,N_17878);
nand U18225 (N_18225,N_17935,N_17747);
xnor U18226 (N_18226,N_17584,N_17536);
nor U18227 (N_18227,N_17641,N_17834);
nand U18228 (N_18228,N_17776,N_17500);
nand U18229 (N_18229,N_17874,N_17916);
xor U18230 (N_18230,N_17853,N_17794);
or U18231 (N_18231,N_17678,N_17899);
nor U18232 (N_18232,N_17933,N_17663);
and U18233 (N_18233,N_17588,N_17672);
or U18234 (N_18234,N_17949,N_17779);
xnor U18235 (N_18235,N_17884,N_17818);
and U18236 (N_18236,N_17775,N_17742);
nor U18237 (N_18237,N_17908,N_17929);
nand U18238 (N_18238,N_17805,N_17947);
nor U18239 (N_18239,N_17789,N_17936);
or U18240 (N_18240,N_17991,N_17728);
or U18241 (N_18241,N_17844,N_17981);
and U18242 (N_18242,N_17734,N_17959);
and U18243 (N_18243,N_17585,N_17721);
nand U18244 (N_18244,N_17561,N_17894);
or U18245 (N_18245,N_17814,N_17602);
nand U18246 (N_18246,N_17824,N_17812);
xor U18247 (N_18247,N_17835,N_17529);
and U18248 (N_18248,N_17767,N_17623);
nor U18249 (N_18249,N_17930,N_17848);
nor U18250 (N_18250,N_17980,N_17930);
nor U18251 (N_18251,N_17772,N_17689);
nor U18252 (N_18252,N_17980,N_17589);
nor U18253 (N_18253,N_17948,N_17919);
nand U18254 (N_18254,N_17791,N_17894);
nand U18255 (N_18255,N_17561,N_17818);
nor U18256 (N_18256,N_17746,N_17820);
nor U18257 (N_18257,N_17574,N_17614);
and U18258 (N_18258,N_17871,N_17870);
nor U18259 (N_18259,N_17954,N_17879);
nor U18260 (N_18260,N_17816,N_17862);
xor U18261 (N_18261,N_17721,N_17719);
and U18262 (N_18262,N_17772,N_17748);
or U18263 (N_18263,N_17825,N_17834);
xor U18264 (N_18264,N_17808,N_17541);
nor U18265 (N_18265,N_17540,N_17784);
nor U18266 (N_18266,N_17918,N_17741);
and U18267 (N_18267,N_17980,N_17657);
xor U18268 (N_18268,N_17720,N_17808);
and U18269 (N_18269,N_17540,N_17562);
nor U18270 (N_18270,N_17899,N_17992);
and U18271 (N_18271,N_17522,N_17766);
nor U18272 (N_18272,N_17636,N_17513);
or U18273 (N_18273,N_17773,N_17569);
nor U18274 (N_18274,N_17795,N_17596);
nor U18275 (N_18275,N_17838,N_17552);
or U18276 (N_18276,N_17784,N_17721);
nand U18277 (N_18277,N_17584,N_17662);
xnor U18278 (N_18278,N_17696,N_17609);
nand U18279 (N_18279,N_17942,N_17913);
and U18280 (N_18280,N_17605,N_17890);
nand U18281 (N_18281,N_17947,N_17951);
or U18282 (N_18282,N_17676,N_17737);
nand U18283 (N_18283,N_17609,N_17613);
nand U18284 (N_18284,N_17649,N_17856);
or U18285 (N_18285,N_17718,N_17656);
and U18286 (N_18286,N_17848,N_17522);
xor U18287 (N_18287,N_17659,N_17691);
and U18288 (N_18288,N_17923,N_17645);
or U18289 (N_18289,N_17734,N_17825);
and U18290 (N_18290,N_17743,N_17673);
and U18291 (N_18291,N_17623,N_17842);
and U18292 (N_18292,N_17567,N_17729);
or U18293 (N_18293,N_17745,N_17546);
and U18294 (N_18294,N_17825,N_17544);
or U18295 (N_18295,N_17892,N_17723);
xnor U18296 (N_18296,N_17706,N_17713);
nand U18297 (N_18297,N_17540,N_17999);
nand U18298 (N_18298,N_17734,N_17841);
nand U18299 (N_18299,N_17512,N_17808);
xor U18300 (N_18300,N_17724,N_17971);
or U18301 (N_18301,N_17591,N_17968);
and U18302 (N_18302,N_17609,N_17903);
nor U18303 (N_18303,N_17860,N_17624);
xor U18304 (N_18304,N_17626,N_17570);
xnor U18305 (N_18305,N_17764,N_17761);
nor U18306 (N_18306,N_17904,N_17549);
nand U18307 (N_18307,N_17537,N_17673);
xor U18308 (N_18308,N_17656,N_17772);
and U18309 (N_18309,N_17872,N_17790);
and U18310 (N_18310,N_17669,N_17858);
or U18311 (N_18311,N_17960,N_17898);
xnor U18312 (N_18312,N_17606,N_17952);
nand U18313 (N_18313,N_17588,N_17981);
and U18314 (N_18314,N_17967,N_17995);
or U18315 (N_18315,N_17763,N_17662);
nand U18316 (N_18316,N_17549,N_17556);
or U18317 (N_18317,N_17755,N_17528);
nand U18318 (N_18318,N_17979,N_17568);
nand U18319 (N_18319,N_17649,N_17789);
nand U18320 (N_18320,N_17603,N_17573);
and U18321 (N_18321,N_17850,N_17634);
nand U18322 (N_18322,N_17877,N_17750);
nor U18323 (N_18323,N_17720,N_17647);
nand U18324 (N_18324,N_17578,N_17977);
xor U18325 (N_18325,N_17771,N_17525);
nor U18326 (N_18326,N_17685,N_17598);
nand U18327 (N_18327,N_17893,N_17662);
and U18328 (N_18328,N_17990,N_17756);
or U18329 (N_18329,N_17883,N_17581);
or U18330 (N_18330,N_17782,N_17629);
nand U18331 (N_18331,N_17914,N_17511);
nand U18332 (N_18332,N_17888,N_17794);
or U18333 (N_18333,N_17827,N_17763);
nor U18334 (N_18334,N_17626,N_17758);
nor U18335 (N_18335,N_17729,N_17574);
nand U18336 (N_18336,N_17903,N_17628);
and U18337 (N_18337,N_17616,N_17697);
and U18338 (N_18338,N_17850,N_17995);
nor U18339 (N_18339,N_17756,N_17862);
or U18340 (N_18340,N_17950,N_17516);
xor U18341 (N_18341,N_17649,N_17587);
nor U18342 (N_18342,N_17906,N_17933);
nand U18343 (N_18343,N_17749,N_17975);
or U18344 (N_18344,N_17997,N_17759);
nor U18345 (N_18345,N_17875,N_17671);
xnor U18346 (N_18346,N_17854,N_17666);
nand U18347 (N_18347,N_17840,N_17853);
and U18348 (N_18348,N_17702,N_17593);
or U18349 (N_18349,N_17646,N_17591);
nor U18350 (N_18350,N_17935,N_17578);
or U18351 (N_18351,N_17672,N_17831);
and U18352 (N_18352,N_17663,N_17850);
nor U18353 (N_18353,N_17768,N_17514);
or U18354 (N_18354,N_17969,N_17729);
or U18355 (N_18355,N_17574,N_17765);
nor U18356 (N_18356,N_17751,N_17999);
and U18357 (N_18357,N_17610,N_17537);
or U18358 (N_18358,N_17696,N_17678);
nor U18359 (N_18359,N_17989,N_17523);
xnor U18360 (N_18360,N_17645,N_17580);
nand U18361 (N_18361,N_17907,N_17645);
xor U18362 (N_18362,N_17785,N_17709);
nand U18363 (N_18363,N_17891,N_17925);
and U18364 (N_18364,N_17904,N_17754);
nor U18365 (N_18365,N_17757,N_17921);
and U18366 (N_18366,N_17936,N_17595);
xnor U18367 (N_18367,N_17947,N_17686);
xnor U18368 (N_18368,N_17733,N_17671);
or U18369 (N_18369,N_17516,N_17914);
and U18370 (N_18370,N_17637,N_17707);
and U18371 (N_18371,N_17985,N_17926);
nand U18372 (N_18372,N_17908,N_17631);
and U18373 (N_18373,N_17725,N_17767);
xnor U18374 (N_18374,N_17704,N_17745);
nand U18375 (N_18375,N_17776,N_17738);
xor U18376 (N_18376,N_17851,N_17648);
and U18377 (N_18377,N_17969,N_17998);
nand U18378 (N_18378,N_17578,N_17816);
or U18379 (N_18379,N_17935,N_17921);
xnor U18380 (N_18380,N_17581,N_17570);
nand U18381 (N_18381,N_17746,N_17702);
or U18382 (N_18382,N_17595,N_17659);
xor U18383 (N_18383,N_17762,N_17730);
nor U18384 (N_18384,N_17732,N_17837);
nor U18385 (N_18385,N_17990,N_17778);
nor U18386 (N_18386,N_17864,N_17852);
and U18387 (N_18387,N_17556,N_17806);
or U18388 (N_18388,N_17784,N_17589);
xor U18389 (N_18389,N_17645,N_17945);
or U18390 (N_18390,N_17668,N_17822);
nor U18391 (N_18391,N_17593,N_17981);
or U18392 (N_18392,N_17926,N_17555);
nor U18393 (N_18393,N_17976,N_17537);
and U18394 (N_18394,N_17661,N_17696);
xor U18395 (N_18395,N_17904,N_17589);
or U18396 (N_18396,N_17584,N_17840);
nand U18397 (N_18397,N_17915,N_17666);
nand U18398 (N_18398,N_17901,N_17689);
nor U18399 (N_18399,N_17914,N_17871);
or U18400 (N_18400,N_17535,N_17694);
xor U18401 (N_18401,N_17636,N_17947);
and U18402 (N_18402,N_17760,N_17742);
nor U18403 (N_18403,N_17523,N_17686);
and U18404 (N_18404,N_17682,N_17695);
and U18405 (N_18405,N_17983,N_17846);
xor U18406 (N_18406,N_17957,N_17980);
and U18407 (N_18407,N_17513,N_17525);
nand U18408 (N_18408,N_17698,N_17617);
nor U18409 (N_18409,N_17659,N_17962);
or U18410 (N_18410,N_17586,N_17637);
or U18411 (N_18411,N_17911,N_17859);
or U18412 (N_18412,N_17617,N_17574);
or U18413 (N_18413,N_17966,N_17956);
and U18414 (N_18414,N_17918,N_17826);
nor U18415 (N_18415,N_17849,N_17735);
and U18416 (N_18416,N_17501,N_17637);
or U18417 (N_18417,N_17790,N_17520);
or U18418 (N_18418,N_17887,N_17683);
nor U18419 (N_18419,N_17583,N_17516);
nand U18420 (N_18420,N_17890,N_17542);
xnor U18421 (N_18421,N_17584,N_17894);
xor U18422 (N_18422,N_17814,N_17789);
nand U18423 (N_18423,N_17785,N_17776);
and U18424 (N_18424,N_17974,N_17569);
xor U18425 (N_18425,N_17822,N_17874);
nand U18426 (N_18426,N_17608,N_17827);
and U18427 (N_18427,N_17821,N_17914);
and U18428 (N_18428,N_17768,N_17886);
nand U18429 (N_18429,N_17883,N_17548);
nand U18430 (N_18430,N_17925,N_17964);
xnor U18431 (N_18431,N_17677,N_17503);
xor U18432 (N_18432,N_17764,N_17666);
xnor U18433 (N_18433,N_17567,N_17649);
xor U18434 (N_18434,N_17780,N_17864);
nand U18435 (N_18435,N_17572,N_17807);
and U18436 (N_18436,N_17590,N_17887);
or U18437 (N_18437,N_17985,N_17786);
nor U18438 (N_18438,N_17926,N_17913);
xnor U18439 (N_18439,N_17959,N_17986);
or U18440 (N_18440,N_17805,N_17522);
and U18441 (N_18441,N_17629,N_17954);
nand U18442 (N_18442,N_17726,N_17793);
nor U18443 (N_18443,N_17862,N_17831);
nor U18444 (N_18444,N_17923,N_17540);
and U18445 (N_18445,N_17759,N_17792);
nor U18446 (N_18446,N_17955,N_17637);
nand U18447 (N_18447,N_17599,N_17640);
and U18448 (N_18448,N_17707,N_17870);
nand U18449 (N_18449,N_17683,N_17881);
nand U18450 (N_18450,N_17870,N_17989);
nor U18451 (N_18451,N_17584,N_17613);
or U18452 (N_18452,N_17795,N_17617);
or U18453 (N_18453,N_17666,N_17522);
or U18454 (N_18454,N_17708,N_17665);
nand U18455 (N_18455,N_17922,N_17569);
or U18456 (N_18456,N_17504,N_17913);
and U18457 (N_18457,N_17629,N_17692);
or U18458 (N_18458,N_17781,N_17736);
and U18459 (N_18459,N_17816,N_17806);
or U18460 (N_18460,N_17661,N_17873);
nand U18461 (N_18461,N_17867,N_17964);
nor U18462 (N_18462,N_17570,N_17959);
xnor U18463 (N_18463,N_17722,N_17635);
xnor U18464 (N_18464,N_17754,N_17898);
nor U18465 (N_18465,N_17927,N_17757);
or U18466 (N_18466,N_17816,N_17635);
and U18467 (N_18467,N_17948,N_17682);
xnor U18468 (N_18468,N_17652,N_17655);
nor U18469 (N_18469,N_17618,N_17824);
or U18470 (N_18470,N_17733,N_17539);
xnor U18471 (N_18471,N_17871,N_17597);
nand U18472 (N_18472,N_17684,N_17859);
or U18473 (N_18473,N_17596,N_17625);
xor U18474 (N_18474,N_17811,N_17783);
nand U18475 (N_18475,N_17775,N_17630);
xor U18476 (N_18476,N_17998,N_17552);
and U18477 (N_18477,N_17767,N_17735);
nor U18478 (N_18478,N_17884,N_17635);
or U18479 (N_18479,N_17715,N_17913);
nor U18480 (N_18480,N_17935,N_17820);
nand U18481 (N_18481,N_17538,N_17825);
or U18482 (N_18482,N_17998,N_17625);
or U18483 (N_18483,N_17609,N_17775);
nor U18484 (N_18484,N_17768,N_17641);
xor U18485 (N_18485,N_17856,N_17615);
or U18486 (N_18486,N_17508,N_17944);
and U18487 (N_18487,N_17725,N_17891);
and U18488 (N_18488,N_17908,N_17507);
and U18489 (N_18489,N_17575,N_17635);
nor U18490 (N_18490,N_17724,N_17940);
xnor U18491 (N_18491,N_17694,N_17815);
and U18492 (N_18492,N_17512,N_17732);
and U18493 (N_18493,N_17556,N_17559);
and U18494 (N_18494,N_17686,N_17780);
or U18495 (N_18495,N_17513,N_17770);
nor U18496 (N_18496,N_17899,N_17959);
nor U18497 (N_18497,N_17644,N_17933);
nand U18498 (N_18498,N_17691,N_17643);
nor U18499 (N_18499,N_17795,N_17529);
xnor U18500 (N_18500,N_18000,N_18240);
nor U18501 (N_18501,N_18206,N_18024);
xor U18502 (N_18502,N_18214,N_18191);
and U18503 (N_18503,N_18430,N_18138);
nand U18504 (N_18504,N_18385,N_18080);
xnor U18505 (N_18505,N_18381,N_18421);
nand U18506 (N_18506,N_18209,N_18187);
xor U18507 (N_18507,N_18189,N_18038);
or U18508 (N_18508,N_18215,N_18291);
nand U18509 (N_18509,N_18300,N_18217);
or U18510 (N_18510,N_18102,N_18406);
nor U18511 (N_18511,N_18053,N_18134);
or U18512 (N_18512,N_18165,N_18472);
nor U18513 (N_18513,N_18477,N_18235);
nand U18514 (N_18514,N_18241,N_18265);
nand U18515 (N_18515,N_18422,N_18366);
nand U18516 (N_18516,N_18297,N_18070);
and U18517 (N_18517,N_18037,N_18302);
and U18518 (N_18518,N_18137,N_18447);
xor U18519 (N_18519,N_18197,N_18391);
xor U18520 (N_18520,N_18319,N_18463);
xor U18521 (N_18521,N_18237,N_18151);
nand U18522 (N_18522,N_18152,N_18320);
nand U18523 (N_18523,N_18095,N_18365);
and U18524 (N_18524,N_18163,N_18042);
xnor U18525 (N_18525,N_18337,N_18147);
or U18526 (N_18526,N_18234,N_18012);
nor U18527 (N_18527,N_18020,N_18470);
and U18528 (N_18528,N_18104,N_18015);
nor U18529 (N_18529,N_18001,N_18378);
or U18530 (N_18530,N_18060,N_18199);
nor U18531 (N_18531,N_18420,N_18142);
nor U18532 (N_18532,N_18374,N_18039);
or U18533 (N_18533,N_18158,N_18145);
nor U18534 (N_18534,N_18059,N_18269);
and U18535 (N_18535,N_18125,N_18239);
xnor U18536 (N_18536,N_18415,N_18476);
xnor U18537 (N_18537,N_18480,N_18310);
nor U18538 (N_18538,N_18375,N_18127);
nand U18539 (N_18539,N_18164,N_18148);
or U18540 (N_18540,N_18454,N_18332);
and U18541 (N_18541,N_18351,N_18271);
xor U18542 (N_18542,N_18333,N_18350);
xnor U18543 (N_18543,N_18123,N_18090);
nand U18544 (N_18544,N_18110,N_18021);
or U18545 (N_18545,N_18380,N_18071);
nor U18546 (N_18546,N_18065,N_18390);
or U18547 (N_18547,N_18186,N_18219);
xor U18548 (N_18548,N_18352,N_18361);
and U18549 (N_18549,N_18314,N_18008);
xnor U18550 (N_18550,N_18464,N_18451);
and U18551 (N_18551,N_18462,N_18274);
xor U18552 (N_18552,N_18418,N_18093);
and U18553 (N_18553,N_18162,N_18167);
xor U18554 (N_18554,N_18312,N_18136);
nand U18555 (N_18555,N_18201,N_18118);
xor U18556 (N_18556,N_18404,N_18325);
nor U18557 (N_18557,N_18182,N_18175);
nor U18558 (N_18558,N_18455,N_18106);
and U18559 (N_18559,N_18224,N_18135);
and U18560 (N_18560,N_18128,N_18097);
nor U18561 (N_18561,N_18054,N_18003);
xor U18562 (N_18562,N_18452,N_18210);
or U18563 (N_18563,N_18481,N_18270);
nor U18564 (N_18564,N_18105,N_18023);
nor U18565 (N_18565,N_18208,N_18223);
and U18566 (N_18566,N_18119,N_18130);
or U18567 (N_18567,N_18304,N_18260);
and U18568 (N_18568,N_18443,N_18305);
and U18569 (N_18569,N_18216,N_18261);
xor U18570 (N_18570,N_18149,N_18379);
nor U18571 (N_18571,N_18282,N_18027);
nor U18572 (N_18572,N_18245,N_18205);
xor U18573 (N_18573,N_18225,N_18246);
xor U18574 (N_18574,N_18446,N_18335);
xor U18575 (N_18575,N_18459,N_18228);
xnor U18576 (N_18576,N_18308,N_18016);
nand U18577 (N_18577,N_18244,N_18120);
xnor U18578 (N_18578,N_18022,N_18401);
and U18579 (N_18579,N_18079,N_18315);
or U18580 (N_18580,N_18388,N_18184);
nand U18581 (N_18581,N_18359,N_18408);
and U18582 (N_18582,N_18416,N_18345);
nand U18583 (N_18583,N_18334,N_18253);
nor U18584 (N_18584,N_18156,N_18083);
or U18585 (N_18585,N_18153,N_18025);
or U18586 (N_18586,N_18107,N_18252);
nor U18587 (N_18587,N_18203,N_18276);
and U18588 (N_18588,N_18195,N_18433);
or U18589 (N_18589,N_18262,N_18340);
and U18590 (N_18590,N_18382,N_18202);
or U18591 (N_18591,N_18207,N_18400);
nor U18592 (N_18592,N_18045,N_18168);
xor U18593 (N_18593,N_18429,N_18236);
nand U18594 (N_18594,N_18428,N_18435);
and U18595 (N_18595,N_18461,N_18456);
nand U18596 (N_18596,N_18154,N_18295);
or U18597 (N_18597,N_18264,N_18457);
or U18598 (N_18598,N_18268,N_18032);
nor U18599 (N_18599,N_18087,N_18434);
xor U18600 (N_18600,N_18306,N_18288);
or U18601 (N_18601,N_18177,N_18460);
xnor U18602 (N_18602,N_18247,N_18383);
nand U18603 (N_18603,N_18348,N_18041);
nand U18604 (N_18604,N_18399,N_18063);
or U18605 (N_18605,N_18331,N_18084);
xor U18606 (N_18606,N_18094,N_18133);
or U18607 (N_18607,N_18115,N_18188);
nand U18608 (N_18608,N_18036,N_18109);
xor U18609 (N_18609,N_18174,N_18483);
nand U18610 (N_18610,N_18254,N_18081);
or U18611 (N_18611,N_18407,N_18121);
nor U18612 (N_18612,N_18222,N_18307);
and U18613 (N_18613,N_18143,N_18492);
xnor U18614 (N_18614,N_18384,N_18330);
nand U18615 (N_18615,N_18267,N_18285);
nand U18616 (N_18616,N_18495,N_18280);
nand U18617 (N_18617,N_18259,N_18360);
nor U18618 (N_18618,N_18474,N_18086);
nand U18619 (N_18619,N_18413,N_18078);
or U18620 (N_18620,N_18465,N_18371);
nor U18621 (N_18621,N_18448,N_18294);
and U18622 (N_18622,N_18030,N_18067);
nor U18623 (N_18623,N_18101,N_18339);
and U18624 (N_18624,N_18160,N_18144);
nand U18625 (N_18625,N_18243,N_18444);
or U18626 (N_18626,N_18486,N_18410);
nor U18627 (N_18627,N_18373,N_18009);
nand U18628 (N_18628,N_18114,N_18129);
nor U18629 (N_18629,N_18449,N_18198);
or U18630 (N_18630,N_18028,N_18050);
and U18631 (N_18631,N_18303,N_18229);
or U18632 (N_18632,N_18031,N_18044);
or U18633 (N_18633,N_18442,N_18498);
xor U18634 (N_18634,N_18146,N_18226);
or U18635 (N_18635,N_18327,N_18193);
nor U18636 (N_18636,N_18355,N_18321);
or U18637 (N_18637,N_18467,N_18436);
nand U18638 (N_18638,N_18073,N_18317);
nand U18639 (N_18639,N_18347,N_18006);
and U18640 (N_18640,N_18493,N_18393);
nand U18641 (N_18641,N_18033,N_18389);
and U18642 (N_18642,N_18497,N_18341);
xor U18643 (N_18643,N_18412,N_18499);
xor U18644 (N_18644,N_18494,N_18004);
or U18645 (N_18645,N_18281,N_18061);
and U18646 (N_18646,N_18257,N_18103);
and U18647 (N_18647,N_18309,N_18091);
nand U18648 (N_18648,N_18034,N_18190);
nor U18649 (N_18649,N_18040,N_18011);
nand U18650 (N_18650,N_18296,N_18284);
xor U18651 (N_18651,N_18238,N_18290);
nand U18652 (N_18652,N_18438,N_18386);
or U18653 (N_18653,N_18277,N_18453);
nand U18654 (N_18654,N_18139,N_18221);
nor U18655 (N_18655,N_18322,N_18230);
or U18656 (N_18656,N_18369,N_18272);
nor U18657 (N_18657,N_18372,N_18287);
or U18658 (N_18658,N_18218,N_18170);
nand U18659 (N_18659,N_18099,N_18005);
xor U18660 (N_18660,N_18396,N_18298);
or U18661 (N_18661,N_18166,N_18096);
nor U18662 (N_18662,N_18484,N_18113);
and U18663 (N_18663,N_18426,N_18362);
nand U18664 (N_18664,N_18316,N_18204);
xor U18665 (N_18665,N_18176,N_18356);
nand U18666 (N_18666,N_18473,N_18466);
nand U18667 (N_18667,N_18392,N_18157);
xor U18668 (N_18668,N_18403,N_18342);
or U18669 (N_18669,N_18323,N_18211);
nor U18670 (N_18670,N_18122,N_18450);
or U18671 (N_18671,N_18414,N_18266);
or U18672 (N_18672,N_18183,N_18013);
xor U18673 (N_18673,N_18066,N_18485);
nand U18674 (N_18674,N_18417,N_18394);
nor U18675 (N_18675,N_18075,N_18299);
and U18676 (N_18676,N_18035,N_18089);
xor U18677 (N_18677,N_18196,N_18116);
or U18678 (N_18678,N_18251,N_18052);
nand U18679 (N_18679,N_18441,N_18482);
nor U18680 (N_18680,N_18488,N_18377);
xor U18681 (N_18681,N_18301,N_18343);
and U18682 (N_18682,N_18180,N_18098);
xor U18683 (N_18683,N_18049,N_18349);
or U18684 (N_18684,N_18082,N_18431);
nand U18685 (N_18685,N_18108,N_18077);
xor U18686 (N_18686,N_18010,N_18289);
nor U18687 (N_18687,N_18336,N_18076);
nand U18688 (N_18688,N_18256,N_18150);
nand U18689 (N_18689,N_18273,N_18131);
nand U18690 (N_18690,N_18064,N_18074);
or U18691 (N_18691,N_18088,N_18169);
nor U18692 (N_18692,N_18026,N_18017);
nand U18693 (N_18693,N_18437,N_18057);
nand U18694 (N_18694,N_18141,N_18019);
or U18695 (N_18695,N_18058,N_18258);
and U18696 (N_18696,N_18292,N_18124);
and U18697 (N_18697,N_18458,N_18425);
nand U18698 (N_18698,N_18367,N_18427);
xor U18699 (N_18699,N_18018,N_18275);
nand U18700 (N_18700,N_18172,N_18043);
or U18701 (N_18701,N_18376,N_18405);
nor U18702 (N_18702,N_18233,N_18051);
xor U18703 (N_18703,N_18242,N_18368);
or U18704 (N_18704,N_18346,N_18111);
or U18705 (N_18705,N_18293,N_18402);
or U18706 (N_18706,N_18029,N_18048);
nor U18707 (N_18707,N_18255,N_18475);
nand U18708 (N_18708,N_18014,N_18370);
nor U18709 (N_18709,N_18338,N_18212);
xnor U18710 (N_18710,N_18155,N_18479);
xnor U18711 (N_18711,N_18478,N_18328);
nor U18712 (N_18712,N_18248,N_18344);
nand U18713 (N_18713,N_18069,N_18132);
xnor U18714 (N_18714,N_18181,N_18445);
xor U18715 (N_18715,N_18409,N_18179);
nand U18716 (N_18716,N_18468,N_18178);
xnor U18717 (N_18717,N_18398,N_18286);
or U18718 (N_18718,N_18068,N_18440);
and U18719 (N_18719,N_18397,N_18112);
or U18720 (N_18720,N_18192,N_18363);
nor U18721 (N_18721,N_18395,N_18220);
nand U18722 (N_18722,N_18002,N_18364);
nor U18723 (N_18723,N_18318,N_18439);
and U18724 (N_18724,N_18047,N_18326);
and U18725 (N_18725,N_18173,N_18046);
xor U18726 (N_18726,N_18491,N_18055);
xor U18727 (N_18727,N_18185,N_18194);
nand U18728 (N_18728,N_18469,N_18250);
and U18729 (N_18729,N_18171,N_18313);
and U18730 (N_18730,N_18311,N_18213);
nor U18731 (N_18731,N_18487,N_18387);
and U18732 (N_18732,N_18200,N_18279);
nand U18733 (N_18733,N_18140,N_18283);
nand U18734 (N_18734,N_18489,N_18056);
nor U18735 (N_18735,N_18496,N_18411);
nor U18736 (N_18736,N_18357,N_18432);
nand U18737 (N_18737,N_18324,N_18062);
xnor U18738 (N_18738,N_18278,N_18419);
or U18739 (N_18739,N_18126,N_18100);
or U18740 (N_18740,N_18358,N_18159);
nor U18741 (N_18741,N_18092,N_18085);
nor U18742 (N_18742,N_18263,N_18249);
or U18743 (N_18743,N_18007,N_18490);
nor U18744 (N_18744,N_18227,N_18353);
nand U18745 (N_18745,N_18232,N_18329);
and U18746 (N_18746,N_18117,N_18161);
nor U18747 (N_18747,N_18471,N_18424);
xor U18748 (N_18748,N_18072,N_18354);
and U18749 (N_18749,N_18423,N_18231);
or U18750 (N_18750,N_18310,N_18437);
nor U18751 (N_18751,N_18367,N_18216);
and U18752 (N_18752,N_18469,N_18220);
nand U18753 (N_18753,N_18461,N_18465);
nand U18754 (N_18754,N_18404,N_18032);
nand U18755 (N_18755,N_18158,N_18100);
xnor U18756 (N_18756,N_18103,N_18313);
nor U18757 (N_18757,N_18364,N_18047);
xor U18758 (N_18758,N_18169,N_18419);
and U18759 (N_18759,N_18474,N_18388);
or U18760 (N_18760,N_18238,N_18325);
nand U18761 (N_18761,N_18493,N_18167);
nand U18762 (N_18762,N_18103,N_18283);
xnor U18763 (N_18763,N_18039,N_18148);
nor U18764 (N_18764,N_18117,N_18172);
or U18765 (N_18765,N_18422,N_18284);
nor U18766 (N_18766,N_18047,N_18027);
nor U18767 (N_18767,N_18131,N_18321);
or U18768 (N_18768,N_18196,N_18490);
xnor U18769 (N_18769,N_18056,N_18459);
or U18770 (N_18770,N_18228,N_18195);
xnor U18771 (N_18771,N_18178,N_18011);
nor U18772 (N_18772,N_18499,N_18002);
or U18773 (N_18773,N_18329,N_18309);
nand U18774 (N_18774,N_18112,N_18442);
xnor U18775 (N_18775,N_18001,N_18167);
nor U18776 (N_18776,N_18386,N_18317);
and U18777 (N_18777,N_18092,N_18302);
nand U18778 (N_18778,N_18091,N_18417);
or U18779 (N_18779,N_18168,N_18095);
nand U18780 (N_18780,N_18384,N_18106);
or U18781 (N_18781,N_18303,N_18267);
nand U18782 (N_18782,N_18412,N_18403);
nor U18783 (N_18783,N_18422,N_18166);
or U18784 (N_18784,N_18276,N_18331);
or U18785 (N_18785,N_18045,N_18492);
nand U18786 (N_18786,N_18347,N_18398);
nor U18787 (N_18787,N_18389,N_18084);
and U18788 (N_18788,N_18283,N_18329);
nand U18789 (N_18789,N_18451,N_18458);
xnor U18790 (N_18790,N_18191,N_18279);
or U18791 (N_18791,N_18415,N_18063);
or U18792 (N_18792,N_18035,N_18061);
nor U18793 (N_18793,N_18320,N_18127);
nand U18794 (N_18794,N_18195,N_18292);
and U18795 (N_18795,N_18399,N_18208);
xor U18796 (N_18796,N_18119,N_18096);
or U18797 (N_18797,N_18353,N_18032);
or U18798 (N_18798,N_18142,N_18332);
nand U18799 (N_18799,N_18392,N_18162);
nor U18800 (N_18800,N_18074,N_18350);
or U18801 (N_18801,N_18003,N_18408);
nor U18802 (N_18802,N_18126,N_18048);
and U18803 (N_18803,N_18243,N_18461);
nand U18804 (N_18804,N_18008,N_18440);
nor U18805 (N_18805,N_18165,N_18444);
nor U18806 (N_18806,N_18352,N_18334);
nor U18807 (N_18807,N_18321,N_18103);
nand U18808 (N_18808,N_18228,N_18405);
and U18809 (N_18809,N_18456,N_18259);
nand U18810 (N_18810,N_18387,N_18219);
nand U18811 (N_18811,N_18055,N_18327);
or U18812 (N_18812,N_18316,N_18475);
nand U18813 (N_18813,N_18269,N_18068);
and U18814 (N_18814,N_18301,N_18488);
xnor U18815 (N_18815,N_18461,N_18437);
and U18816 (N_18816,N_18197,N_18122);
nand U18817 (N_18817,N_18302,N_18053);
and U18818 (N_18818,N_18470,N_18137);
nand U18819 (N_18819,N_18263,N_18348);
nand U18820 (N_18820,N_18019,N_18413);
nor U18821 (N_18821,N_18189,N_18059);
xor U18822 (N_18822,N_18117,N_18274);
xor U18823 (N_18823,N_18243,N_18100);
nor U18824 (N_18824,N_18344,N_18370);
or U18825 (N_18825,N_18386,N_18142);
and U18826 (N_18826,N_18062,N_18177);
nand U18827 (N_18827,N_18375,N_18403);
and U18828 (N_18828,N_18341,N_18231);
nor U18829 (N_18829,N_18154,N_18141);
or U18830 (N_18830,N_18223,N_18255);
or U18831 (N_18831,N_18268,N_18362);
nand U18832 (N_18832,N_18413,N_18392);
and U18833 (N_18833,N_18226,N_18048);
or U18834 (N_18834,N_18405,N_18471);
or U18835 (N_18835,N_18343,N_18226);
nand U18836 (N_18836,N_18469,N_18334);
and U18837 (N_18837,N_18067,N_18451);
nand U18838 (N_18838,N_18045,N_18434);
nor U18839 (N_18839,N_18476,N_18156);
xnor U18840 (N_18840,N_18490,N_18099);
nand U18841 (N_18841,N_18329,N_18423);
and U18842 (N_18842,N_18475,N_18146);
nand U18843 (N_18843,N_18376,N_18125);
nor U18844 (N_18844,N_18336,N_18212);
nand U18845 (N_18845,N_18327,N_18103);
or U18846 (N_18846,N_18494,N_18206);
nor U18847 (N_18847,N_18069,N_18335);
or U18848 (N_18848,N_18105,N_18073);
xnor U18849 (N_18849,N_18226,N_18457);
nand U18850 (N_18850,N_18362,N_18489);
and U18851 (N_18851,N_18218,N_18422);
nand U18852 (N_18852,N_18398,N_18404);
and U18853 (N_18853,N_18220,N_18123);
or U18854 (N_18854,N_18164,N_18388);
xnor U18855 (N_18855,N_18492,N_18375);
nor U18856 (N_18856,N_18313,N_18256);
xor U18857 (N_18857,N_18309,N_18445);
xnor U18858 (N_18858,N_18061,N_18424);
and U18859 (N_18859,N_18235,N_18090);
and U18860 (N_18860,N_18420,N_18440);
or U18861 (N_18861,N_18465,N_18347);
and U18862 (N_18862,N_18415,N_18058);
nand U18863 (N_18863,N_18322,N_18013);
xor U18864 (N_18864,N_18460,N_18200);
nor U18865 (N_18865,N_18300,N_18323);
nor U18866 (N_18866,N_18184,N_18030);
nand U18867 (N_18867,N_18130,N_18284);
or U18868 (N_18868,N_18340,N_18121);
and U18869 (N_18869,N_18240,N_18146);
nand U18870 (N_18870,N_18340,N_18178);
and U18871 (N_18871,N_18328,N_18332);
or U18872 (N_18872,N_18154,N_18063);
or U18873 (N_18873,N_18151,N_18177);
and U18874 (N_18874,N_18473,N_18024);
or U18875 (N_18875,N_18247,N_18136);
nor U18876 (N_18876,N_18368,N_18364);
and U18877 (N_18877,N_18449,N_18148);
nand U18878 (N_18878,N_18294,N_18154);
or U18879 (N_18879,N_18345,N_18153);
xnor U18880 (N_18880,N_18340,N_18004);
nor U18881 (N_18881,N_18214,N_18464);
nor U18882 (N_18882,N_18065,N_18461);
nor U18883 (N_18883,N_18468,N_18389);
xor U18884 (N_18884,N_18025,N_18123);
nor U18885 (N_18885,N_18031,N_18398);
and U18886 (N_18886,N_18398,N_18351);
xor U18887 (N_18887,N_18331,N_18038);
xor U18888 (N_18888,N_18437,N_18484);
nor U18889 (N_18889,N_18487,N_18242);
xnor U18890 (N_18890,N_18166,N_18001);
xor U18891 (N_18891,N_18350,N_18203);
or U18892 (N_18892,N_18411,N_18041);
xnor U18893 (N_18893,N_18148,N_18469);
nor U18894 (N_18894,N_18451,N_18010);
or U18895 (N_18895,N_18004,N_18193);
and U18896 (N_18896,N_18344,N_18103);
or U18897 (N_18897,N_18306,N_18291);
xnor U18898 (N_18898,N_18461,N_18041);
xnor U18899 (N_18899,N_18006,N_18467);
nand U18900 (N_18900,N_18327,N_18147);
and U18901 (N_18901,N_18255,N_18189);
or U18902 (N_18902,N_18392,N_18184);
nand U18903 (N_18903,N_18213,N_18425);
and U18904 (N_18904,N_18284,N_18228);
or U18905 (N_18905,N_18396,N_18141);
and U18906 (N_18906,N_18187,N_18348);
and U18907 (N_18907,N_18104,N_18167);
and U18908 (N_18908,N_18483,N_18048);
nand U18909 (N_18909,N_18121,N_18053);
or U18910 (N_18910,N_18199,N_18387);
xnor U18911 (N_18911,N_18382,N_18404);
nor U18912 (N_18912,N_18371,N_18262);
nand U18913 (N_18913,N_18389,N_18267);
or U18914 (N_18914,N_18397,N_18205);
or U18915 (N_18915,N_18297,N_18492);
nand U18916 (N_18916,N_18245,N_18433);
nand U18917 (N_18917,N_18425,N_18028);
and U18918 (N_18918,N_18256,N_18495);
xnor U18919 (N_18919,N_18168,N_18058);
and U18920 (N_18920,N_18326,N_18497);
nand U18921 (N_18921,N_18485,N_18138);
xnor U18922 (N_18922,N_18105,N_18295);
xor U18923 (N_18923,N_18175,N_18101);
and U18924 (N_18924,N_18271,N_18346);
and U18925 (N_18925,N_18169,N_18412);
or U18926 (N_18926,N_18477,N_18229);
nand U18927 (N_18927,N_18488,N_18394);
and U18928 (N_18928,N_18363,N_18299);
nand U18929 (N_18929,N_18455,N_18122);
nand U18930 (N_18930,N_18456,N_18037);
nand U18931 (N_18931,N_18466,N_18151);
and U18932 (N_18932,N_18308,N_18119);
nor U18933 (N_18933,N_18039,N_18407);
nand U18934 (N_18934,N_18305,N_18291);
or U18935 (N_18935,N_18173,N_18218);
nor U18936 (N_18936,N_18191,N_18035);
xnor U18937 (N_18937,N_18050,N_18434);
or U18938 (N_18938,N_18221,N_18249);
nand U18939 (N_18939,N_18381,N_18245);
or U18940 (N_18940,N_18256,N_18407);
or U18941 (N_18941,N_18064,N_18444);
nand U18942 (N_18942,N_18379,N_18042);
and U18943 (N_18943,N_18160,N_18088);
nand U18944 (N_18944,N_18484,N_18062);
and U18945 (N_18945,N_18186,N_18090);
or U18946 (N_18946,N_18470,N_18087);
and U18947 (N_18947,N_18049,N_18244);
xnor U18948 (N_18948,N_18402,N_18233);
nand U18949 (N_18949,N_18210,N_18320);
xor U18950 (N_18950,N_18363,N_18449);
and U18951 (N_18951,N_18273,N_18097);
xor U18952 (N_18952,N_18087,N_18402);
nor U18953 (N_18953,N_18361,N_18307);
nor U18954 (N_18954,N_18186,N_18141);
and U18955 (N_18955,N_18174,N_18107);
xnor U18956 (N_18956,N_18481,N_18427);
or U18957 (N_18957,N_18075,N_18275);
nand U18958 (N_18958,N_18401,N_18387);
nand U18959 (N_18959,N_18132,N_18315);
xnor U18960 (N_18960,N_18453,N_18439);
and U18961 (N_18961,N_18041,N_18225);
xnor U18962 (N_18962,N_18276,N_18064);
or U18963 (N_18963,N_18224,N_18432);
nand U18964 (N_18964,N_18218,N_18163);
nand U18965 (N_18965,N_18044,N_18480);
xnor U18966 (N_18966,N_18198,N_18472);
nor U18967 (N_18967,N_18263,N_18319);
nor U18968 (N_18968,N_18264,N_18095);
and U18969 (N_18969,N_18325,N_18112);
nand U18970 (N_18970,N_18182,N_18116);
xnor U18971 (N_18971,N_18400,N_18497);
and U18972 (N_18972,N_18354,N_18207);
nand U18973 (N_18973,N_18155,N_18174);
xor U18974 (N_18974,N_18265,N_18242);
xor U18975 (N_18975,N_18445,N_18489);
and U18976 (N_18976,N_18182,N_18395);
or U18977 (N_18977,N_18137,N_18348);
or U18978 (N_18978,N_18128,N_18465);
nor U18979 (N_18979,N_18310,N_18180);
nand U18980 (N_18980,N_18479,N_18054);
xnor U18981 (N_18981,N_18379,N_18385);
nand U18982 (N_18982,N_18420,N_18320);
or U18983 (N_18983,N_18003,N_18256);
nand U18984 (N_18984,N_18258,N_18397);
and U18985 (N_18985,N_18329,N_18203);
nand U18986 (N_18986,N_18362,N_18192);
or U18987 (N_18987,N_18200,N_18246);
nor U18988 (N_18988,N_18300,N_18123);
or U18989 (N_18989,N_18245,N_18276);
or U18990 (N_18990,N_18044,N_18260);
nand U18991 (N_18991,N_18282,N_18308);
or U18992 (N_18992,N_18314,N_18195);
nor U18993 (N_18993,N_18167,N_18303);
xnor U18994 (N_18994,N_18007,N_18371);
nor U18995 (N_18995,N_18277,N_18098);
and U18996 (N_18996,N_18209,N_18486);
nand U18997 (N_18997,N_18205,N_18189);
or U18998 (N_18998,N_18356,N_18431);
xor U18999 (N_18999,N_18150,N_18060);
xnor U19000 (N_19000,N_18623,N_18990);
nand U19001 (N_19001,N_18538,N_18602);
and U19002 (N_19002,N_18892,N_18649);
xor U19003 (N_19003,N_18918,N_18738);
nor U19004 (N_19004,N_18636,N_18837);
xnor U19005 (N_19005,N_18994,N_18825);
or U19006 (N_19006,N_18520,N_18725);
and U19007 (N_19007,N_18769,N_18693);
xnor U19008 (N_19008,N_18665,N_18827);
nand U19009 (N_19009,N_18529,N_18749);
nor U19010 (N_19010,N_18876,N_18708);
and U19011 (N_19011,N_18977,N_18836);
nand U19012 (N_19012,N_18785,N_18916);
xnor U19013 (N_19013,N_18691,N_18500);
and U19014 (N_19014,N_18878,N_18931);
and U19015 (N_19015,N_18954,N_18597);
nand U19016 (N_19016,N_18546,N_18633);
nor U19017 (N_19017,N_18604,N_18849);
xnor U19018 (N_19018,N_18700,N_18591);
or U19019 (N_19019,N_18800,N_18563);
nand U19020 (N_19020,N_18787,N_18619);
nand U19021 (N_19021,N_18550,N_18777);
nor U19022 (N_19022,N_18618,N_18654);
and U19023 (N_19023,N_18898,N_18944);
xnor U19024 (N_19024,N_18516,N_18941);
nand U19025 (N_19025,N_18624,N_18603);
nand U19026 (N_19026,N_18702,N_18524);
nor U19027 (N_19027,N_18584,N_18780);
and U19028 (N_19028,N_18621,N_18906);
nor U19029 (N_19029,N_18672,N_18804);
and U19030 (N_19030,N_18860,N_18763);
nor U19031 (N_19031,N_18698,N_18686);
or U19032 (N_19032,N_18681,N_18788);
xnor U19033 (N_19033,N_18796,N_18543);
nor U19034 (N_19034,N_18940,N_18542);
and U19035 (N_19035,N_18853,N_18746);
or U19036 (N_19036,N_18679,N_18536);
nor U19037 (N_19037,N_18824,N_18528);
or U19038 (N_19038,N_18645,N_18851);
or U19039 (N_19039,N_18970,N_18730);
or U19040 (N_19040,N_18888,N_18910);
or U19041 (N_19041,N_18856,N_18525);
and U19042 (N_19042,N_18518,N_18705);
xnor U19043 (N_19043,N_18617,N_18963);
xor U19044 (N_19044,N_18660,N_18987);
or U19045 (N_19045,N_18998,N_18807);
nand U19046 (N_19046,N_18894,N_18723);
or U19047 (N_19047,N_18579,N_18883);
nand U19048 (N_19048,N_18687,N_18674);
nand U19049 (N_19049,N_18526,N_18846);
nand U19050 (N_19050,N_18647,N_18710);
nand U19051 (N_19051,N_18507,N_18552);
nor U19052 (N_19052,N_18799,N_18947);
nand U19053 (N_19053,N_18544,N_18783);
or U19054 (N_19054,N_18714,N_18770);
and U19055 (N_19055,N_18775,N_18774);
nand U19056 (N_19056,N_18991,N_18781);
and U19057 (N_19057,N_18611,N_18965);
nand U19058 (N_19058,N_18966,N_18822);
or U19059 (N_19059,N_18872,N_18949);
and U19060 (N_19060,N_18850,N_18881);
nor U19061 (N_19061,N_18841,N_18605);
nand U19062 (N_19062,N_18508,N_18534);
nand U19063 (N_19063,N_18643,N_18820);
nand U19064 (N_19064,N_18974,N_18573);
and U19065 (N_19065,N_18740,N_18964);
xnor U19066 (N_19066,N_18988,N_18968);
nor U19067 (N_19067,N_18902,N_18896);
nor U19068 (N_19068,N_18903,N_18612);
and U19069 (N_19069,N_18720,N_18939);
or U19070 (N_19070,N_18598,N_18690);
xor U19071 (N_19071,N_18831,N_18502);
nand U19072 (N_19072,N_18967,N_18727);
nor U19073 (N_19073,N_18514,N_18874);
nand U19074 (N_19074,N_18628,N_18812);
and U19075 (N_19075,N_18537,N_18762);
nor U19076 (N_19076,N_18829,N_18557);
xor U19077 (N_19077,N_18569,N_18663);
nor U19078 (N_19078,N_18784,N_18900);
nand U19079 (N_19079,N_18639,N_18531);
xnor U19080 (N_19080,N_18759,N_18771);
nor U19081 (N_19081,N_18701,N_18752);
nor U19082 (N_19082,N_18779,N_18521);
and U19083 (N_19083,N_18601,N_18561);
nand U19084 (N_19084,N_18513,N_18957);
nor U19085 (N_19085,N_18745,N_18983);
xor U19086 (N_19086,N_18928,N_18667);
nor U19087 (N_19087,N_18840,N_18657);
xnor U19088 (N_19088,N_18862,N_18515);
nor U19089 (N_19089,N_18540,N_18772);
nor U19090 (N_19090,N_18927,N_18973);
and U19091 (N_19091,N_18950,N_18659);
xnor U19092 (N_19092,N_18697,N_18936);
nor U19093 (N_19093,N_18845,N_18703);
or U19094 (N_19094,N_18562,N_18778);
or U19095 (N_19095,N_18585,N_18713);
or U19096 (N_19096,N_18620,N_18732);
nor U19097 (N_19097,N_18907,N_18652);
xnor U19098 (N_19098,N_18593,N_18934);
and U19099 (N_19099,N_18958,N_18870);
and U19100 (N_19100,N_18889,N_18721);
and U19101 (N_19101,N_18764,N_18982);
xor U19102 (N_19102,N_18935,N_18885);
nor U19103 (N_19103,N_18826,N_18637);
nor U19104 (N_19104,N_18553,N_18993);
xnor U19105 (N_19105,N_18960,N_18979);
and U19106 (N_19106,N_18805,N_18776);
xor U19107 (N_19107,N_18737,N_18635);
and U19108 (N_19108,N_18980,N_18819);
or U19109 (N_19109,N_18678,N_18753);
nor U19110 (N_19110,N_18891,N_18689);
and U19111 (N_19111,N_18914,N_18984);
nor U19112 (N_19112,N_18908,N_18504);
xnor U19113 (N_19113,N_18684,N_18782);
and U19114 (N_19114,N_18739,N_18625);
nand U19115 (N_19115,N_18522,N_18816);
or U19116 (N_19116,N_18580,N_18731);
or U19117 (N_19117,N_18677,N_18981);
and U19118 (N_19118,N_18632,N_18761);
nand U19119 (N_19119,N_18886,N_18661);
nor U19120 (N_19120,N_18995,N_18533);
nor U19121 (N_19121,N_18909,N_18609);
or U19122 (N_19122,N_18666,N_18608);
nand U19123 (N_19123,N_18791,N_18817);
or U19124 (N_19124,N_18638,N_18786);
xor U19125 (N_19125,N_18999,N_18747);
and U19126 (N_19126,N_18879,N_18932);
xnor U19127 (N_19127,N_18863,N_18847);
nor U19128 (N_19128,N_18951,N_18871);
or U19129 (N_19129,N_18716,N_18748);
xnor U19130 (N_19130,N_18578,N_18595);
and U19131 (N_19131,N_18673,N_18583);
and U19132 (N_19132,N_18728,N_18880);
xor U19133 (N_19133,N_18961,N_18726);
nor U19134 (N_19134,N_18848,N_18838);
or U19135 (N_19135,N_18556,N_18839);
xnor U19136 (N_19136,N_18946,N_18530);
nand U19137 (N_19137,N_18616,N_18952);
nor U19138 (N_19138,N_18688,N_18555);
or U19139 (N_19139,N_18589,N_18955);
xnor U19140 (N_19140,N_18629,N_18539);
nand U19141 (N_19141,N_18832,N_18933);
or U19142 (N_19142,N_18717,N_18765);
or U19143 (N_19143,N_18711,N_18712);
xor U19144 (N_19144,N_18794,N_18692);
nor U19145 (N_19145,N_18724,N_18828);
nand U19146 (N_19146,N_18867,N_18795);
and U19147 (N_19147,N_18741,N_18859);
or U19148 (N_19148,N_18613,N_18656);
nor U19149 (N_19149,N_18685,N_18718);
xor U19150 (N_19150,N_18587,N_18615);
nor U19151 (N_19151,N_18877,N_18789);
xor U19152 (N_19152,N_18582,N_18676);
and U19153 (N_19153,N_18890,N_18948);
xor U19154 (N_19154,N_18901,N_18996);
nand U19155 (N_19155,N_18913,N_18869);
nand U19156 (N_19156,N_18986,N_18792);
nor U19157 (N_19157,N_18942,N_18699);
nand U19158 (N_19158,N_18801,N_18924);
or U19159 (N_19159,N_18565,N_18576);
xor U19160 (N_19160,N_18959,N_18581);
and U19161 (N_19161,N_18707,N_18547);
and U19162 (N_19162,N_18842,N_18938);
nand U19163 (N_19163,N_18923,N_18930);
or U19164 (N_19164,N_18943,N_18627);
nand U19165 (N_19165,N_18568,N_18755);
xor U19166 (N_19166,N_18926,N_18564);
or U19167 (N_19167,N_18743,N_18655);
nand U19168 (N_19168,N_18682,N_18921);
xnor U19169 (N_19169,N_18833,N_18919);
or U19170 (N_19170,N_18767,N_18835);
nand U19171 (N_19171,N_18953,N_18857);
nor U19172 (N_19172,N_18945,N_18733);
xnor U19173 (N_19173,N_18830,N_18642);
or U19174 (N_19174,N_18566,N_18742);
nand U19175 (N_19175,N_18917,N_18852);
and U19176 (N_19176,N_18600,N_18962);
xor U19177 (N_19177,N_18814,N_18855);
nor U19178 (N_19178,N_18640,N_18675);
nand U19179 (N_19179,N_18545,N_18815);
and U19180 (N_19180,N_18823,N_18937);
or U19181 (N_19181,N_18868,N_18861);
or U19182 (N_19182,N_18607,N_18882);
and U19183 (N_19183,N_18813,N_18523);
and U19184 (N_19184,N_18736,N_18798);
and U19185 (N_19185,N_18884,N_18558);
or U19186 (N_19186,N_18866,N_18821);
and U19187 (N_19187,N_18806,N_18641);
and U19188 (N_19188,N_18592,N_18843);
nand U19189 (N_19189,N_18997,N_18662);
nand U19190 (N_19190,N_18535,N_18517);
nand U19191 (N_19191,N_18750,N_18634);
and U19192 (N_19192,N_18505,N_18596);
nor U19193 (N_19193,N_18757,N_18735);
nand U19194 (N_19194,N_18811,N_18560);
or U19195 (N_19195,N_18511,N_18744);
nand U19196 (N_19196,N_18873,N_18729);
or U19197 (N_19197,N_18834,N_18956);
or U19198 (N_19198,N_18904,N_18658);
xor U19199 (N_19199,N_18519,N_18709);
xnor U19200 (N_19200,N_18670,N_18695);
nor U19201 (N_19201,N_18864,N_18793);
xor U19202 (N_19202,N_18803,N_18650);
xnor U19203 (N_19203,N_18758,N_18512);
nand U19204 (N_19204,N_18683,N_18577);
nor U19205 (N_19205,N_18754,N_18631);
nor U19206 (N_19206,N_18644,N_18671);
xnor U19207 (N_19207,N_18532,N_18549);
and U19208 (N_19208,N_18810,N_18590);
xor U19209 (N_19209,N_18875,N_18844);
nand U19210 (N_19210,N_18858,N_18905);
or U19211 (N_19211,N_18922,N_18929);
nand U19212 (N_19212,N_18893,N_18694);
and U19213 (N_19213,N_18567,N_18626);
nand U19214 (N_19214,N_18897,N_18760);
and U19215 (N_19215,N_18976,N_18588);
nand U19216 (N_19216,N_18527,N_18985);
xor U19217 (N_19217,N_18809,N_18648);
nand U19218 (N_19218,N_18989,N_18610);
nor U19219 (N_19219,N_18768,N_18975);
xnor U19220 (N_19220,N_18630,N_18972);
nor U19221 (N_19221,N_18510,N_18594);
or U19222 (N_19222,N_18622,N_18586);
or U19223 (N_19223,N_18554,N_18915);
and U19224 (N_19224,N_18912,N_18756);
or U19225 (N_19225,N_18548,N_18808);
nand U19226 (N_19226,N_18559,N_18575);
xnor U19227 (N_19227,N_18978,N_18992);
nand U19228 (N_19228,N_18599,N_18865);
nor U19229 (N_19229,N_18696,N_18887);
nor U19230 (N_19230,N_18509,N_18501);
nand U19231 (N_19231,N_18715,N_18572);
nor U19232 (N_19232,N_18653,N_18541);
and U19233 (N_19233,N_18551,N_18969);
or U19234 (N_19234,N_18680,N_18704);
nor U19235 (N_19235,N_18895,N_18818);
and U19236 (N_19236,N_18802,N_18790);
nor U19237 (N_19237,N_18664,N_18571);
nand U19238 (N_19238,N_18719,N_18773);
and U19239 (N_19239,N_18606,N_18911);
or U19240 (N_19240,N_18751,N_18766);
or U19241 (N_19241,N_18574,N_18646);
nor U19242 (N_19242,N_18925,N_18614);
or U19243 (N_19243,N_18570,N_18669);
or U19244 (N_19244,N_18854,N_18506);
or U19245 (N_19245,N_18899,N_18920);
and U19246 (N_19246,N_18734,N_18668);
nand U19247 (N_19247,N_18706,N_18651);
nor U19248 (N_19248,N_18971,N_18722);
nor U19249 (N_19249,N_18797,N_18503);
or U19250 (N_19250,N_18720,N_18553);
and U19251 (N_19251,N_18623,N_18781);
xnor U19252 (N_19252,N_18614,N_18930);
nand U19253 (N_19253,N_18879,N_18714);
or U19254 (N_19254,N_18646,N_18982);
nor U19255 (N_19255,N_18945,N_18641);
xnor U19256 (N_19256,N_18794,N_18884);
nand U19257 (N_19257,N_18559,N_18938);
or U19258 (N_19258,N_18751,N_18712);
and U19259 (N_19259,N_18721,N_18623);
and U19260 (N_19260,N_18765,N_18590);
or U19261 (N_19261,N_18858,N_18538);
xnor U19262 (N_19262,N_18751,N_18523);
and U19263 (N_19263,N_18504,N_18816);
nor U19264 (N_19264,N_18681,N_18809);
nand U19265 (N_19265,N_18558,N_18777);
nor U19266 (N_19266,N_18503,N_18872);
xnor U19267 (N_19267,N_18995,N_18549);
or U19268 (N_19268,N_18570,N_18832);
nor U19269 (N_19269,N_18529,N_18687);
and U19270 (N_19270,N_18835,N_18763);
nor U19271 (N_19271,N_18510,N_18691);
and U19272 (N_19272,N_18878,N_18934);
nand U19273 (N_19273,N_18509,N_18821);
xor U19274 (N_19274,N_18547,N_18705);
nor U19275 (N_19275,N_18548,N_18798);
nor U19276 (N_19276,N_18613,N_18760);
or U19277 (N_19277,N_18731,N_18885);
nand U19278 (N_19278,N_18747,N_18854);
and U19279 (N_19279,N_18535,N_18635);
nand U19280 (N_19280,N_18813,N_18739);
or U19281 (N_19281,N_18937,N_18739);
nand U19282 (N_19282,N_18783,N_18944);
nand U19283 (N_19283,N_18807,N_18532);
or U19284 (N_19284,N_18521,N_18951);
nor U19285 (N_19285,N_18561,N_18764);
xnor U19286 (N_19286,N_18879,N_18726);
nor U19287 (N_19287,N_18911,N_18693);
xor U19288 (N_19288,N_18613,N_18659);
and U19289 (N_19289,N_18636,N_18838);
nor U19290 (N_19290,N_18597,N_18930);
nand U19291 (N_19291,N_18854,N_18795);
and U19292 (N_19292,N_18791,N_18747);
nand U19293 (N_19293,N_18616,N_18522);
nand U19294 (N_19294,N_18782,N_18736);
nand U19295 (N_19295,N_18973,N_18911);
and U19296 (N_19296,N_18744,N_18835);
xor U19297 (N_19297,N_18981,N_18730);
and U19298 (N_19298,N_18968,N_18830);
nand U19299 (N_19299,N_18754,N_18841);
or U19300 (N_19300,N_18848,N_18882);
and U19301 (N_19301,N_18529,N_18815);
nor U19302 (N_19302,N_18920,N_18518);
nor U19303 (N_19303,N_18893,N_18918);
and U19304 (N_19304,N_18719,N_18749);
xnor U19305 (N_19305,N_18840,N_18678);
xnor U19306 (N_19306,N_18574,N_18621);
nand U19307 (N_19307,N_18504,N_18524);
nor U19308 (N_19308,N_18649,N_18847);
and U19309 (N_19309,N_18652,N_18635);
nor U19310 (N_19310,N_18887,N_18527);
xnor U19311 (N_19311,N_18756,N_18674);
nand U19312 (N_19312,N_18566,N_18876);
xor U19313 (N_19313,N_18944,N_18974);
and U19314 (N_19314,N_18844,N_18778);
xor U19315 (N_19315,N_18890,N_18675);
or U19316 (N_19316,N_18978,N_18544);
xnor U19317 (N_19317,N_18535,N_18627);
xor U19318 (N_19318,N_18997,N_18946);
or U19319 (N_19319,N_18729,N_18694);
or U19320 (N_19320,N_18908,N_18703);
or U19321 (N_19321,N_18939,N_18787);
xnor U19322 (N_19322,N_18549,N_18950);
or U19323 (N_19323,N_18802,N_18811);
and U19324 (N_19324,N_18772,N_18695);
nor U19325 (N_19325,N_18833,N_18872);
and U19326 (N_19326,N_18752,N_18670);
or U19327 (N_19327,N_18776,N_18670);
nor U19328 (N_19328,N_18663,N_18671);
xor U19329 (N_19329,N_18644,N_18709);
xor U19330 (N_19330,N_18662,N_18525);
nand U19331 (N_19331,N_18500,N_18613);
nor U19332 (N_19332,N_18566,N_18595);
xnor U19333 (N_19333,N_18658,N_18568);
or U19334 (N_19334,N_18873,N_18841);
nand U19335 (N_19335,N_18886,N_18601);
nor U19336 (N_19336,N_18595,N_18764);
nand U19337 (N_19337,N_18822,N_18544);
nor U19338 (N_19338,N_18914,N_18737);
nand U19339 (N_19339,N_18616,N_18963);
and U19340 (N_19340,N_18877,N_18676);
xnor U19341 (N_19341,N_18711,N_18617);
nand U19342 (N_19342,N_18524,N_18550);
xor U19343 (N_19343,N_18589,N_18594);
or U19344 (N_19344,N_18560,N_18528);
nand U19345 (N_19345,N_18595,N_18846);
xnor U19346 (N_19346,N_18665,N_18655);
and U19347 (N_19347,N_18617,N_18975);
or U19348 (N_19348,N_18960,N_18506);
and U19349 (N_19349,N_18595,N_18562);
nand U19350 (N_19350,N_18936,N_18951);
and U19351 (N_19351,N_18666,N_18582);
or U19352 (N_19352,N_18606,N_18627);
nor U19353 (N_19353,N_18855,N_18568);
nand U19354 (N_19354,N_18985,N_18930);
and U19355 (N_19355,N_18556,N_18695);
and U19356 (N_19356,N_18613,N_18640);
nand U19357 (N_19357,N_18546,N_18834);
nand U19358 (N_19358,N_18870,N_18904);
and U19359 (N_19359,N_18702,N_18868);
and U19360 (N_19360,N_18879,N_18607);
nand U19361 (N_19361,N_18986,N_18573);
and U19362 (N_19362,N_18502,N_18867);
xnor U19363 (N_19363,N_18948,N_18956);
or U19364 (N_19364,N_18506,N_18750);
nand U19365 (N_19365,N_18848,N_18754);
and U19366 (N_19366,N_18725,N_18689);
xnor U19367 (N_19367,N_18816,N_18828);
nand U19368 (N_19368,N_18903,N_18946);
xnor U19369 (N_19369,N_18935,N_18647);
nor U19370 (N_19370,N_18919,N_18654);
nor U19371 (N_19371,N_18723,N_18846);
nand U19372 (N_19372,N_18633,N_18501);
nand U19373 (N_19373,N_18900,N_18687);
and U19374 (N_19374,N_18971,N_18821);
and U19375 (N_19375,N_18968,N_18965);
nor U19376 (N_19376,N_18751,N_18693);
xnor U19377 (N_19377,N_18819,N_18590);
nor U19378 (N_19378,N_18677,N_18789);
nand U19379 (N_19379,N_18890,N_18631);
or U19380 (N_19380,N_18702,N_18985);
xnor U19381 (N_19381,N_18805,N_18733);
and U19382 (N_19382,N_18644,N_18849);
and U19383 (N_19383,N_18924,N_18553);
nand U19384 (N_19384,N_18553,N_18922);
nor U19385 (N_19385,N_18533,N_18796);
xnor U19386 (N_19386,N_18794,N_18557);
xnor U19387 (N_19387,N_18798,N_18612);
nand U19388 (N_19388,N_18663,N_18648);
nand U19389 (N_19389,N_18888,N_18505);
nand U19390 (N_19390,N_18679,N_18841);
and U19391 (N_19391,N_18523,N_18836);
or U19392 (N_19392,N_18680,N_18625);
or U19393 (N_19393,N_18720,N_18759);
and U19394 (N_19394,N_18959,N_18856);
and U19395 (N_19395,N_18675,N_18683);
and U19396 (N_19396,N_18699,N_18796);
and U19397 (N_19397,N_18769,N_18798);
xnor U19398 (N_19398,N_18585,N_18562);
xor U19399 (N_19399,N_18766,N_18626);
or U19400 (N_19400,N_18620,N_18831);
xnor U19401 (N_19401,N_18667,N_18846);
xor U19402 (N_19402,N_18798,N_18626);
or U19403 (N_19403,N_18789,N_18855);
xor U19404 (N_19404,N_18963,N_18525);
nand U19405 (N_19405,N_18660,N_18575);
or U19406 (N_19406,N_18714,N_18940);
and U19407 (N_19407,N_18649,N_18937);
or U19408 (N_19408,N_18796,N_18676);
nor U19409 (N_19409,N_18762,N_18654);
nor U19410 (N_19410,N_18553,N_18872);
and U19411 (N_19411,N_18861,N_18567);
or U19412 (N_19412,N_18973,N_18680);
xnor U19413 (N_19413,N_18504,N_18912);
or U19414 (N_19414,N_18836,N_18973);
nor U19415 (N_19415,N_18748,N_18896);
xor U19416 (N_19416,N_18895,N_18770);
nor U19417 (N_19417,N_18850,N_18550);
and U19418 (N_19418,N_18614,N_18915);
and U19419 (N_19419,N_18504,N_18772);
or U19420 (N_19420,N_18755,N_18901);
nand U19421 (N_19421,N_18896,N_18742);
and U19422 (N_19422,N_18918,N_18941);
and U19423 (N_19423,N_18674,N_18916);
nand U19424 (N_19424,N_18937,N_18671);
or U19425 (N_19425,N_18703,N_18905);
and U19426 (N_19426,N_18963,N_18809);
xor U19427 (N_19427,N_18849,N_18648);
and U19428 (N_19428,N_18539,N_18737);
or U19429 (N_19429,N_18929,N_18700);
nor U19430 (N_19430,N_18975,N_18833);
or U19431 (N_19431,N_18603,N_18998);
nor U19432 (N_19432,N_18642,N_18804);
and U19433 (N_19433,N_18661,N_18719);
nor U19434 (N_19434,N_18635,N_18804);
nand U19435 (N_19435,N_18529,N_18789);
or U19436 (N_19436,N_18919,N_18643);
nand U19437 (N_19437,N_18812,N_18883);
xor U19438 (N_19438,N_18526,N_18952);
nand U19439 (N_19439,N_18718,N_18508);
or U19440 (N_19440,N_18973,N_18650);
or U19441 (N_19441,N_18693,N_18515);
and U19442 (N_19442,N_18608,N_18837);
or U19443 (N_19443,N_18728,N_18634);
nor U19444 (N_19444,N_18929,N_18640);
or U19445 (N_19445,N_18992,N_18809);
nand U19446 (N_19446,N_18616,N_18694);
xor U19447 (N_19447,N_18604,N_18750);
xor U19448 (N_19448,N_18790,N_18852);
or U19449 (N_19449,N_18992,N_18843);
nor U19450 (N_19450,N_18748,N_18856);
nand U19451 (N_19451,N_18842,N_18599);
and U19452 (N_19452,N_18697,N_18686);
or U19453 (N_19453,N_18739,N_18744);
and U19454 (N_19454,N_18978,N_18920);
and U19455 (N_19455,N_18576,N_18915);
and U19456 (N_19456,N_18678,N_18613);
nand U19457 (N_19457,N_18885,N_18593);
and U19458 (N_19458,N_18563,N_18584);
and U19459 (N_19459,N_18552,N_18703);
nand U19460 (N_19460,N_18752,N_18772);
or U19461 (N_19461,N_18949,N_18831);
nand U19462 (N_19462,N_18656,N_18655);
nand U19463 (N_19463,N_18926,N_18963);
nand U19464 (N_19464,N_18978,N_18557);
nand U19465 (N_19465,N_18655,N_18690);
nand U19466 (N_19466,N_18967,N_18556);
or U19467 (N_19467,N_18928,N_18512);
nor U19468 (N_19468,N_18790,N_18707);
nand U19469 (N_19469,N_18768,N_18620);
or U19470 (N_19470,N_18903,N_18980);
nand U19471 (N_19471,N_18819,N_18727);
nand U19472 (N_19472,N_18877,N_18790);
nor U19473 (N_19473,N_18730,N_18648);
and U19474 (N_19474,N_18773,N_18799);
xnor U19475 (N_19475,N_18618,N_18673);
nand U19476 (N_19476,N_18739,N_18690);
nand U19477 (N_19477,N_18638,N_18862);
and U19478 (N_19478,N_18796,N_18869);
xnor U19479 (N_19479,N_18707,N_18933);
and U19480 (N_19480,N_18628,N_18547);
nor U19481 (N_19481,N_18693,N_18861);
nor U19482 (N_19482,N_18999,N_18882);
nand U19483 (N_19483,N_18683,N_18757);
and U19484 (N_19484,N_18799,N_18744);
nand U19485 (N_19485,N_18621,N_18970);
nand U19486 (N_19486,N_18672,N_18751);
nor U19487 (N_19487,N_18674,N_18823);
nor U19488 (N_19488,N_18964,N_18757);
nand U19489 (N_19489,N_18915,N_18930);
and U19490 (N_19490,N_18511,N_18523);
or U19491 (N_19491,N_18580,N_18850);
and U19492 (N_19492,N_18860,N_18881);
xor U19493 (N_19493,N_18918,N_18625);
nand U19494 (N_19494,N_18502,N_18837);
nor U19495 (N_19495,N_18714,N_18602);
nor U19496 (N_19496,N_18961,N_18538);
nor U19497 (N_19497,N_18783,N_18860);
or U19498 (N_19498,N_18950,N_18778);
nor U19499 (N_19499,N_18730,N_18601);
and U19500 (N_19500,N_19388,N_19083);
xnor U19501 (N_19501,N_19425,N_19216);
or U19502 (N_19502,N_19107,N_19387);
xnor U19503 (N_19503,N_19131,N_19036);
nor U19504 (N_19504,N_19420,N_19471);
nor U19505 (N_19505,N_19209,N_19356);
nor U19506 (N_19506,N_19454,N_19426);
or U19507 (N_19507,N_19057,N_19439);
or U19508 (N_19508,N_19304,N_19381);
and U19509 (N_19509,N_19460,N_19213);
or U19510 (N_19510,N_19328,N_19284);
or U19511 (N_19511,N_19062,N_19244);
nor U19512 (N_19512,N_19455,N_19446);
nor U19513 (N_19513,N_19316,N_19429);
xor U19514 (N_19514,N_19030,N_19151);
nor U19515 (N_19515,N_19177,N_19330);
nand U19516 (N_19516,N_19458,N_19462);
nand U19517 (N_19517,N_19317,N_19155);
nor U19518 (N_19518,N_19363,N_19094);
nand U19519 (N_19519,N_19436,N_19437);
nor U19520 (N_19520,N_19236,N_19310);
xor U19521 (N_19521,N_19185,N_19093);
and U19522 (N_19522,N_19096,N_19366);
nand U19523 (N_19523,N_19005,N_19137);
nor U19524 (N_19524,N_19190,N_19012);
xnor U19525 (N_19525,N_19272,N_19476);
xnor U19526 (N_19526,N_19459,N_19335);
nor U19527 (N_19527,N_19170,N_19283);
and U19528 (N_19528,N_19312,N_19119);
nand U19529 (N_19529,N_19334,N_19331);
xnor U19530 (N_19530,N_19053,N_19218);
or U19531 (N_19531,N_19203,N_19428);
nor U19532 (N_19532,N_19327,N_19480);
xnor U19533 (N_19533,N_19302,N_19435);
and U19534 (N_19534,N_19117,N_19440);
and U19535 (N_19535,N_19291,N_19377);
nor U19536 (N_19536,N_19142,N_19488);
xor U19537 (N_19537,N_19417,N_19208);
or U19538 (N_19538,N_19132,N_19069);
nor U19539 (N_19539,N_19329,N_19163);
nor U19540 (N_19540,N_19063,N_19207);
nor U19541 (N_19541,N_19006,N_19221);
nand U19542 (N_19542,N_19433,N_19411);
xnor U19543 (N_19543,N_19452,N_19072);
nand U19544 (N_19544,N_19368,N_19251);
xor U19545 (N_19545,N_19343,N_19201);
nor U19546 (N_19546,N_19453,N_19182);
nor U19547 (N_19547,N_19038,N_19199);
xnor U19548 (N_19548,N_19285,N_19442);
xor U19549 (N_19549,N_19139,N_19000);
nor U19550 (N_19550,N_19238,N_19263);
nor U19551 (N_19551,N_19065,N_19332);
or U19552 (N_19552,N_19260,N_19373);
xnor U19553 (N_19553,N_19273,N_19074);
nand U19554 (N_19554,N_19194,N_19308);
xnor U19555 (N_19555,N_19295,N_19214);
nor U19556 (N_19556,N_19071,N_19434);
nand U19557 (N_19557,N_19324,N_19148);
and U19558 (N_19558,N_19350,N_19371);
or U19559 (N_19559,N_19192,N_19470);
nor U19560 (N_19560,N_19269,N_19043);
nand U19561 (N_19561,N_19042,N_19009);
and U19562 (N_19562,N_19301,N_19109);
xnor U19563 (N_19563,N_19003,N_19432);
xnor U19564 (N_19564,N_19088,N_19242);
nor U19565 (N_19565,N_19322,N_19020);
or U19566 (N_19566,N_19122,N_19247);
or U19567 (N_19567,N_19372,N_19204);
xnor U19568 (N_19568,N_19211,N_19075);
nor U19569 (N_19569,N_19186,N_19378);
or U19570 (N_19570,N_19278,N_19008);
nor U19571 (N_19571,N_19326,N_19281);
nor U19572 (N_19572,N_19469,N_19015);
xor U19573 (N_19573,N_19487,N_19147);
nand U19574 (N_19574,N_19212,N_19115);
and U19575 (N_19575,N_19073,N_19105);
nor U19576 (N_19576,N_19154,N_19309);
and U19577 (N_19577,N_19023,N_19467);
nand U19578 (N_19578,N_19286,N_19489);
nor U19579 (N_19579,N_19364,N_19473);
and U19580 (N_19580,N_19397,N_19391);
xnor U19581 (N_19581,N_19416,N_19110);
nand U19582 (N_19582,N_19261,N_19392);
and U19583 (N_19583,N_19128,N_19494);
nand U19584 (N_19584,N_19360,N_19362);
or U19585 (N_19585,N_19400,N_19121);
nor U19586 (N_19586,N_19293,N_19232);
nor U19587 (N_19587,N_19159,N_19379);
or U19588 (N_19588,N_19288,N_19376);
and U19589 (N_19589,N_19412,N_19191);
and U19590 (N_19590,N_19033,N_19405);
or U19591 (N_19591,N_19361,N_19246);
xor U19592 (N_19592,N_19479,N_19485);
and U19593 (N_19593,N_19018,N_19415);
and U19594 (N_19594,N_19339,N_19114);
and U19595 (N_19595,N_19183,N_19138);
nand U19596 (N_19596,N_19438,N_19133);
or U19597 (N_19597,N_19380,N_19359);
nor U19598 (N_19598,N_19102,N_19490);
or U19599 (N_19599,N_19079,N_19080);
nor U19600 (N_19600,N_19497,N_19456);
nand U19601 (N_19601,N_19370,N_19172);
nor U19602 (N_19602,N_19058,N_19262);
or U19603 (N_19603,N_19225,N_19457);
nor U19604 (N_19604,N_19315,N_19461);
xor U19605 (N_19605,N_19255,N_19265);
nand U19606 (N_19606,N_19205,N_19101);
and U19607 (N_19607,N_19077,N_19189);
xor U19608 (N_19608,N_19493,N_19385);
nor U19609 (N_19609,N_19064,N_19258);
or U19610 (N_19610,N_19342,N_19045);
nand U19611 (N_19611,N_19025,N_19197);
and U19612 (N_19612,N_19168,N_19399);
nand U19613 (N_19613,N_19389,N_19268);
xnor U19614 (N_19614,N_19341,N_19245);
nand U19615 (N_19615,N_19078,N_19249);
xnor U19616 (N_19616,N_19424,N_19113);
xor U19617 (N_19617,N_19303,N_19034);
nor U19618 (N_19618,N_19321,N_19289);
xor U19619 (N_19619,N_19323,N_19031);
nand U19620 (N_19620,N_19149,N_19252);
and U19621 (N_19621,N_19418,N_19481);
nand U19622 (N_19622,N_19103,N_19085);
nand U19623 (N_19623,N_19338,N_19174);
or U19624 (N_19624,N_19144,N_19024);
or U19625 (N_19625,N_19164,N_19002);
nand U19626 (N_19626,N_19290,N_19407);
nand U19627 (N_19627,N_19318,N_19365);
or U19628 (N_19628,N_19219,N_19052);
nor U19629 (N_19629,N_19448,N_19040);
xor U19630 (N_19630,N_19171,N_19305);
nor U19631 (N_19631,N_19398,N_19431);
and U19632 (N_19632,N_19298,N_19287);
nor U19633 (N_19633,N_19181,N_19230);
nand U19634 (N_19634,N_19141,N_19097);
nand U19635 (N_19635,N_19066,N_19491);
nor U19636 (N_19636,N_19222,N_19382);
and U19637 (N_19637,N_19325,N_19135);
and U19638 (N_19638,N_19019,N_19390);
nor U19639 (N_19639,N_19028,N_19233);
xor U19640 (N_19640,N_19153,N_19130);
xnor U19641 (N_19641,N_19257,N_19237);
and U19642 (N_19642,N_19108,N_19210);
nand U19643 (N_19643,N_19294,N_19050);
or U19644 (N_19644,N_19337,N_19195);
and U19645 (N_19645,N_19313,N_19406);
nand U19646 (N_19646,N_19419,N_19224);
nor U19647 (N_19647,N_19482,N_19145);
nor U19648 (N_19648,N_19167,N_19344);
xnor U19649 (N_19649,N_19266,N_19410);
and U19650 (N_19650,N_19013,N_19044);
xnor U19651 (N_19651,N_19367,N_19220);
and U19652 (N_19652,N_19136,N_19129);
nand U19653 (N_19653,N_19248,N_19270);
nor U19654 (N_19654,N_19127,N_19178);
or U19655 (N_19655,N_19444,N_19158);
nor U19656 (N_19656,N_19175,N_19466);
and U19657 (N_19657,N_19292,N_19187);
and U19658 (N_19658,N_19346,N_19267);
xor U19659 (N_19659,N_19306,N_19047);
nand U19660 (N_19660,N_19095,N_19282);
nor U19661 (N_19661,N_19276,N_19125);
xnor U19662 (N_19662,N_19423,N_19484);
nand U19663 (N_19663,N_19202,N_19051);
and U19664 (N_19664,N_19229,N_19228);
and U19665 (N_19665,N_19451,N_19014);
nand U19666 (N_19666,N_19395,N_19348);
and U19667 (N_19667,N_19166,N_19239);
nor U19668 (N_19668,N_19447,N_19496);
and U19669 (N_19669,N_19374,N_19472);
nor U19670 (N_19670,N_19126,N_19478);
nor U19671 (N_19671,N_19223,N_19347);
nand U19672 (N_19672,N_19413,N_19180);
nor U19673 (N_19673,N_19277,N_19032);
or U19674 (N_19674,N_19100,N_19037);
and U19675 (N_19675,N_19393,N_19234);
nor U19676 (N_19676,N_19320,N_19059);
nor U19677 (N_19677,N_19254,N_19215);
nand U19678 (N_19678,N_19021,N_19235);
and U19679 (N_19679,N_19492,N_19156);
xnor U19680 (N_19680,N_19421,N_19430);
xor U19681 (N_19681,N_19241,N_19081);
xor U19682 (N_19682,N_19314,N_19465);
and U19683 (N_19683,N_19226,N_19243);
nand U19684 (N_19684,N_19396,N_19300);
or U19685 (N_19685,N_19198,N_19001);
nand U19686 (N_19686,N_19082,N_19048);
nand U19687 (N_19687,N_19076,N_19275);
xor U19688 (N_19688,N_19404,N_19146);
xor U19689 (N_19689,N_19296,N_19087);
or U19690 (N_19690,N_19067,N_19422);
xor U19691 (N_19691,N_19427,N_19483);
xnor U19692 (N_19692,N_19055,N_19409);
nand U19693 (N_19693,N_19169,N_19264);
xnor U19694 (N_19694,N_19026,N_19091);
nand U19695 (N_19695,N_19150,N_19477);
xor U19696 (N_19696,N_19084,N_19160);
and U19697 (N_19697,N_19157,N_19061);
xor U19698 (N_19698,N_19319,N_19336);
xor U19699 (N_19699,N_19035,N_19123);
nor U19700 (N_19700,N_19140,N_19092);
and U19701 (N_19701,N_19375,N_19414);
nand U19702 (N_19702,N_19274,N_19162);
nor U19703 (N_19703,N_19253,N_19450);
nor U19704 (N_19704,N_19054,N_19016);
nand U19705 (N_19705,N_19099,N_19299);
nor U19706 (N_19706,N_19217,N_19049);
nor U19707 (N_19707,N_19463,N_19060);
or U19708 (N_19708,N_19124,N_19152);
xnor U19709 (N_19709,N_19120,N_19259);
nand U19710 (N_19710,N_19256,N_19468);
nand U19711 (N_19711,N_19464,N_19352);
nor U19712 (N_19712,N_19475,N_19118);
nand U19713 (N_19713,N_19022,N_19056);
xor U19714 (N_19714,N_19394,N_19089);
nor U19715 (N_19715,N_19474,N_19353);
nor U19716 (N_19716,N_19086,N_19041);
nand U19717 (N_19717,N_19231,N_19499);
nor U19718 (N_19718,N_19345,N_19112);
or U19719 (N_19719,N_19240,N_19271);
nor U19720 (N_19720,N_19486,N_19090);
nor U19721 (N_19721,N_19196,N_19449);
nor U19722 (N_19722,N_19354,N_19227);
xor U19723 (N_19723,N_19403,N_19402);
xnor U19724 (N_19724,N_19176,N_19017);
or U19725 (N_19725,N_19358,N_19401);
nor U19726 (N_19726,N_19029,N_19039);
and U19727 (N_19727,N_19173,N_19386);
and U19728 (N_19728,N_19111,N_19010);
xor U19729 (N_19729,N_19441,N_19070);
nand U19730 (N_19730,N_19349,N_19007);
nor U19731 (N_19731,N_19161,N_19280);
nand U19732 (N_19732,N_19011,N_19068);
xor U19733 (N_19733,N_19200,N_19333);
and U19734 (N_19734,N_19495,N_19134);
xor U19735 (N_19735,N_19369,N_19355);
or U19736 (N_19736,N_19104,N_19307);
nor U19737 (N_19737,N_19250,N_19184);
nor U19738 (N_19738,N_19297,N_19106);
nor U19739 (N_19739,N_19027,N_19143);
and U19740 (N_19740,N_19383,N_19351);
xor U19741 (N_19741,N_19206,N_19445);
nor U19742 (N_19742,N_19165,N_19098);
nand U19743 (N_19743,N_19311,N_19408);
or U19744 (N_19744,N_19498,N_19046);
xnor U19745 (N_19745,N_19443,N_19340);
or U19746 (N_19746,N_19384,N_19357);
or U19747 (N_19747,N_19004,N_19116);
nor U19748 (N_19748,N_19193,N_19279);
nor U19749 (N_19749,N_19188,N_19179);
nor U19750 (N_19750,N_19342,N_19181);
or U19751 (N_19751,N_19392,N_19133);
nand U19752 (N_19752,N_19287,N_19077);
nand U19753 (N_19753,N_19270,N_19459);
xnor U19754 (N_19754,N_19429,N_19238);
nor U19755 (N_19755,N_19081,N_19092);
xnor U19756 (N_19756,N_19207,N_19463);
and U19757 (N_19757,N_19113,N_19020);
xnor U19758 (N_19758,N_19237,N_19354);
nand U19759 (N_19759,N_19262,N_19099);
xor U19760 (N_19760,N_19121,N_19311);
nor U19761 (N_19761,N_19163,N_19254);
nor U19762 (N_19762,N_19336,N_19246);
or U19763 (N_19763,N_19381,N_19177);
and U19764 (N_19764,N_19262,N_19183);
nand U19765 (N_19765,N_19473,N_19393);
and U19766 (N_19766,N_19176,N_19206);
nand U19767 (N_19767,N_19492,N_19446);
xnor U19768 (N_19768,N_19081,N_19286);
or U19769 (N_19769,N_19008,N_19044);
nor U19770 (N_19770,N_19129,N_19273);
or U19771 (N_19771,N_19367,N_19304);
and U19772 (N_19772,N_19263,N_19432);
or U19773 (N_19773,N_19370,N_19287);
and U19774 (N_19774,N_19180,N_19122);
xnor U19775 (N_19775,N_19288,N_19020);
and U19776 (N_19776,N_19148,N_19496);
xnor U19777 (N_19777,N_19150,N_19152);
nor U19778 (N_19778,N_19204,N_19189);
and U19779 (N_19779,N_19444,N_19293);
or U19780 (N_19780,N_19127,N_19334);
nor U19781 (N_19781,N_19409,N_19296);
nor U19782 (N_19782,N_19001,N_19418);
nor U19783 (N_19783,N_19058,N_19304);
nand U19784 (N_19784,N_19451,N_19222);
and U19785 (N_19785,N_19048,N_19250);
nand U19786 (N_19786,N_19400,N_19481);
or U19787 (N_19787,N_19158,N_19438);
xor U19788 (N_19788,N_19035,N_19236);
nand U19789 (N_19789,N_19122,N_19411);
xor U19790 (N_19790,N_19395,N_19376);
nand U19791 (N_19791,N_19136,N_19320);
or U19792 (N_19792,N_19287,N_19393);
and U19793 (N_19793,N_19316,N_19056);
nor U19794 (N_19794,N_19217,N_19363);
and U19795 (N_19795,N_19236,N_19435);
nor U19796 (N_19796,N_19379,N_19051);
xnor U19797 (N_19797,N_19462,N_19414);
xnor U19798 (N_19798,N_19434,N_19159);
nor U19799 (N_19799,N_19373,N_19144);
xnor U19800 (N_19800,N_19473,N_19367);
or U19801 (N_19801,N_19294,N_19217);
nor U19802 (N_19802,N_19359,N_19251);
or U19803 (N_19803,N_19155,N_19395);
and U19804 (N_19804,N_19470,N_19005);
and U19805 (N_19805,N_19270,N_19375);
xor U19806 (N_19806,N_19413,N_19144);
and U19807 (N_19807,N_19212,N_19405);
or U19808 (N_19808,N_19375,N_19316);
nor U19809 (N_19809,N_19471,N_19104);
and U19810 (N_19810,N_19443,N_19485);
xnor U19811 (N_19811,N_19270,N_19472);
nand U19812 (N_19812,N_19015,N_19103);
nand U19813 (N_19813,N_19373,N_19249);
or U19814 (N_19814,N_19136,N_19210);
nor U19815 (N_19815,N_19377,N_19484);
and U19816 (N_19816,N_19035,N_19418);
and U19817 (N_19817,N_19085,N_19097);
and U19818 (N_19818,N_19331,N_19093);
or U19819 (N_19819,N_19470,N_19136);
xnor U19820 (N_19820,N_19462,N_19099);
nand U19821 (N_19821,N_19255,N_19154);
nand U19822 (N_19822,N_19135,N_19182);
and U19823 (N_19823,N_19017,N_19083);
xnor U19824 (N_19824,N_19095,N_19373);
nor U19825 (N_19825,N_19030,N_19493);
xor U19826 (N_19826,N_19264,N_19205);
and U19827 (N_19827,N_19081,N_19341);
nand U19828 (N_19828,N_19063,N_19150);
nand U19829 (N_19829,N_19236,N_19179);
or U19830 (N_19830,N_19328,N_19359);
xor U19831 (N_19831,N_19005,N_19420);
and U19832 (N_19832,N_19472,N_19317);
nand U19833 (N_19833,N_19266,N_19373);
and U19834 (N_19834,N_19052,N_19158);
nor U19835 (N_19835,N_19137,N_19268);
nor U19836 (N_19836,N_19422,N_19065);
nand U19837 (N_19837,N_19018,N_19465);
nor U19838 (N_19838,N_19156,N_19010);
and U19839 (N_19839,N_19013,N_19195);
or U19840 (N_19840,N_19303,N_19473);
xor U19841 (N_19841,N_19467,N_19246);
or U19842 (N_19842,N_19028,N_19218);
or U19843 (N_19843,N_19492,N_19358);
or U19844 (N_19844,N_19454,N_19210);
or U19845 (N_19845,N_19097,N_19267);
nand U19846 (N_19846,N_19057,N_19360);
xor U19847 (N_19847,N_19242,N_19240);
or U19848 (N_19848,N_19148,N_19492);
nand U19849 (N_19849,N_19155,N_19489);
nor U19850 (N_19850,N_19244,N_19477);
or U19851 (N_19851,N_19173,N_19189);
and U19852 (N_19852,N_19300,N_19442);
nand U19853 (N_19853,N_19366,N_19089);
or U19854 (N_19854,N_19086,N_19437);
xnor U19855 (N_19855,N_19133,N_19470);
nor U19856 (N_19856,N_19161,N_19034);
xnor U19857 (N_19857,N_19386,N_19354);
and U19858 (N_19858,N_19490,N_19427);
or U19859 (N_19859,N_19071,N_19288);
xnor U19860 (N_19860,N_19172,N_19427);
xor U19861 (N_19861,N_19357,N_19406);
or U19862 (N_19862,N_19497,N_19157);
or U19863 (N_19863,N_19299,N_19022);
or U19864 (N_19864,N_19061,N_19356);
nor U19865 (N_19865,N_19327,N_19211);
or U19866 (N_19866,N_19104,N_19255);
nand U19867 (N_19867,N_19267,N_19123);
nand U19868 (N_19868,N_19347,N_19173);
xnor U19869 (N_19869,N_19265,N_19103);
xor U19870 (N_19870,N_19006,N_19195);
nor U19871 (N_19871,N_19211,N_19165);
xnor U19872 (N_19872,N_19050,N_19447);
or U19873 (N_19873,N_19148,N_19180);
xnor U19874 (N_19874,N_19367,N_19387);
and U19875 (N_19875,N_19211,N_19269);
nand U19876 (N_19876,N_19461,N_19120);
nor U19877 (N_19877,N_19105,N_19201);
and U19878 (N_19878,N_19124,N_19001);
or U19879 (N_19879,N_19120,N_19473);
and U19880 (N_19880,N_19317,N_19454);
nand U19881 (N_19881,N_19117,N_19330);
nand U19882 (N_19882,N_19290,N_19015);
xor U19883 (N_19883,N_19279,N_19485);
xor U19884 (N_19884,N_19190,N_19187);
nand U19885 (N_19885,N_19405,N_19233);
and U19886 (N_19886,N_19437,N_19246);
nand U19887 (N_19887,N_19274,N_19229);
nor U19888 (N_19888,N_19181,N_19158);
or U19889 (N_19889,N_19212,N_19138);
and U19890 (N_19890,N_19165,N_19237);
nand U19891 (N_19891,N_19343,N_19130);
xor U19892 (N_19892,N_19014,N_19459);
nor U19893 (N_19893,N_19197,N_19296);
xor U19894 (N_19894,N_19368,N_19197);
nand U19895 (N_19895,N_19025,N_19121);
or U19896 (N_19896,N_19358,N_19493);
xnor U19897 (N_19897,N_19060,N_19163);
or U19898 (N_19898,N_19016,N_19346);
and U19899 (N_19899,N_19256,N_19328);
xnor U19900 (N_19900,N_19263,N_19434);
nor U19901 (N_19901,N_19497,N_19284);
xnor U19902 (N_19902,N_19174,N_19398);
nand U19903 (N_19903,N_19101,N_19349);
and U19904 (N_19904,N_19224,N_19156);
and U19905 (N_19905,N_19219,N_19023);
or U19906 (N_19906,N_19308,N_19089);
nor U19907 (N_19907,N_19494,N_19385);
xnor U19908 (N_19908,N_19045,N_19120);
nor U19909 (N_19909,N_19082,N_19407);
xor U19910 (N_19910,N_19452,N_19221);
nand U19911 (N_19911,N_19496,N_19315);
nor U19912 (N_19912,N_19344,N_19147);
or U19913 (N_19913,N_19260,N_19106);
xnor U19914 (N_19914,N_19095,N_19019);
nand U19915 (N_19915,N_19393,N_19178);
and U19916 (N_19916,N_19449,N_19256);
or U19917 (N_19917,N_19377,N_19234);
nand U19918 (N_19918,N_19486,N_19006);
and U19919 (N_19919,N_19016,N_19098);
and U19920 (N_19920,N_19241,N_19086);
and U19921 (N_19921,N_19224,N_19266);
or U19922 (N_19922,N_19087,N_19093);
xor U19923 (N_19923,N_19434,N_19074);
and U19924 (N_19924,N_19402,N_19116);
and U19925 (N_19925,N_19047,N_19459);
or U19926 (N_19926,N_19010,N_19478);
nand U19927 (N_19927,N_19123,N_19357);
xor U19928 (N_19928,N_19036,N_19469);
or U19929 (N_19929,N_19480,N_19273);
or U19930 (N_19930,N_19219,N_19051);
nor U19931 (N_19931,N_19044,N_19146);
and U19932 (N_19932,N_19128,N_19208);
and U19933 (N_19933,N_19315,N_19278);
and U19934 (N_19934,N_19384,N_19170);
nor U19935 (N_19935,N_19330,N_19331);
nor U19936 (N_19936,N_19489,N_19348);
nor U19937 (N_19937,N_19032,N_19251);
and U19938 (N_19938,N_19075,N_19158);
or U19939 (N_19939,N_19224,N_19154);
nor U19940 (N_19940,N_19110,N_19142);
nand U19941 (N_19941,N_19225,N_19487);
or U19942 (N_19942,N_19119,N_19064);
or U19943 (N_19943,N_19171,N_19418);
nor U19944 (N_19944,N_19223,N_19282);
or U19945 (N_19945,N_19158,N_19491);
xor U19946 (N_19946,N_19123,N_19100);
xnor U19947 (N_19947,N_19460,N_19253);
or U19948 (N_19948,N_19426,N_19406);
xnor U19949 (N_19949,N_19156,N_19326);
nor U19950 (N_19950,N_19136,N_19473);
and U19951 (N_19951,N_19074,N_19431);
nor U19952 (N_19952,N_19265,N_19045);
nor U19953 (N_19953,N_19455,N_19140);
or U19954 (N_19954,N_19016,N_19034);
or U19955 (N_19955,N_19120,N_19480);
or U19956 (N_19956,N_19284,N_19485);
xor U19957 (N_19957,N_19064,N_19447);
nor U19958 (N_19958,N_19019,N_19098);
or U19959 (N_19959,N_19043,N_19493);
xnor U19960 (N_19960,N_19471,N_19194);
or U19961 (N_19961,N_19213,N_19027);
nand U19962 (N_19962,N_19474,N_19109);
and U19963 (N_19963,N_19409,N_19186);
and U19964 (N_19964,N_19063,N_19293);
nor U19965 (N_19965,N_19211,N_19031);
xnor U19966 (N_19966,N_19481,N_19128);
nand U19967 (N_19967,N_19191,N_19311);
or U19968 (N_19968,N_19214,N_19170);
xor U19969 (N_19969,N_19319,N_19067);
nand U19970 (N_19970,N_19425,N_19276);
xor U19971 (N_19971,N_19187,N_19412);
nand U19972 (N_19972,N_19075,N_19483);
xor U19973 (N_19973,N_19227,N_19100);
nor U19974 (N_19974,N_19169,N_19057);
or U19975 (N_19975,N_19258,N_19075);
nand U19976 (N_19976,N_19335,N_19162);
nor U19977 (N_19977,N_19400,N_19153);
and U19978 (N_19978,N_19415,N_19488);
or U19979 (N_19979,N_19345,N_19034);
or U19980 (N_19980,N_19152,N_19076);
or U19981 (N_19981,N_19268,N_19122);
nor U19982 (N_19982,N_19406,N_19150);
nor U19983 (N_19983,N_19417,N_19380);
and U19984 (N_19984,N_19081,N_19300);
or U19985 (N_19985,N_19134,N_19334);
xor U19986 (N_19986,N_19116,N_19162);
nor U19987 (N_19987,N_19438,N_19346);
and U19988 (N_19988,N_19079,N_19303);
nand U19989 (N_19989,N_19321,N_19455);
nand U19990 (N_19990,N_19449,N_19319);
nor U19991 (N_19991,N_19095,N_19369);
xor U19992 (N_19992,N_19212,N_19338);
xnor U19993 (N_19993,N_19062,N_19006);
and U19994 (N_19994,N_19114,N_19060);
xnor U19995 (N_19995,N_19283,N_19094);
nand U19996 (N_19996,N_19283,N_19226);
and U19997 (N_19997,N_19056,N_19073);
xor U19998 (N_19998,N_19498,N_19039);
nand U19999 (N_19999,N_19070,N_19359);
and U20000 (N_20000,N_19769,N_19581);
nor U20001 (N_20001,N_19900,N_19676);
nor U20002 (N_20002,N_19990,N_19851);
and U20003 (N_20003,N_19880,N_19584);
or U20004 (N_20004,N_19820,N_19735);
nor U20005 (N_20005,N_19726,N_19641);
or U20006 (N_20006,N_19977,N_19685);
nand U20007 (N_20007,N_19892,N_19833);
or U20008 (N_20008,N_19717,N_19598);
nor U20009 (N_20009,N_19835,N_19810);
or U20010 (N_20010,N_19597,N_19976);
nor U20011 (N_20011,N_19995,N_19682);
xnor U20012 (N_20012,N_19801,N_19629);
nand U20013 (N_20013,N_19754,N_19572);
xnor U20014 (N_20014,N_19909,N_19505);
or U20015 (N_20015,N_19815,N_19924);
nand U20016 (N_20016,N_19780,N_19929);
xor U20017 (N_20017,N_19928,N_19679);
nor U20018 (N_20018,N_19960,N_19906);
nand U20019 (N_20019,N_19839,N_19761);
or U20020 (N_20020,N_19519,N_19999);
and U20021 (N_20021,N_19596,N_19905);
and U20022 (N_20022,N_19746,N_19849);
or U20023 (N_20023,N_19721,N_19850);
or U20024 (N_20024,N_19805,N_19671);
nand U20025 (N_20025,N_19760,N_19785);
xor U20026 (N_20026,N_19954,N_19503);
xor U20027 (N_20027,N_19506,N_19922);
nand U20028 (N_20028,N_19654,N_19628);
nand U20029 (N_20029,N_19707,N_19652);
xor U20030 (N_20030,N_19606,N_19804);
nand U20031 (N_20031,N_19936,N_19718);
xor U20032 (N_20032,N_19670,N_19779);
and U20033 (N_20033,N_19702,N_19994);
xnor U20034 (N_20034,N_19797,N_19813);
nor U20035 (N_20035,N_19555,N_19817);
or U20036 (N_20036,N_19586,N_19799);
or U20037 (N_20037,N_19933,N_19895);
nand U20038 (N_20038,N_19864,N_19631);
nor U20039 (N_20039,N_19877,N_19811);
nand U20040 (N_20040,N_19703,N_19547);
and U20041 (N_20041,N_19668,N_19580);
and U20042 (N_20042,N_19786,N_19768);
or U20043 (N_20043,N_19957,N_19614);
or U20044 (N_20044,N_19619,N_19648);
xor U20045 (N_20045,N_19823,N_19918);
nor U20046 (N_20046,N_19891,N_19605);
xor U20047 (N_20047,N_19621,N_19622);
or U20048 (N_20048,N_19642,N_19512);
nor U20049 (N_20049,N_19940,N_19744);
xnor U20050 (N_20050,N_19727,N_19963);
nand U20051 (N_20051,N_19883,N_19587);
nand U20052 (N_20052,N_19537,N_19788);
xor U20053 (N_20053,N_19912,N_19659);
and U20054 (N_20054,N_19603,N_19569);
xor U20055 (N_20055,N_19790,N_19705);
or U20056 (N_20056,N_19923,N_19948);
or U20057 (N_20057,N_19568,N_19860);
xnor U20058 (N_20058,N_19806,N_19694);
or U20059 (N_20059,N_19508,N_19767);
nor U20060 (N_20060,N_19657,N_19543);
and U20061 (N_20061,N_19870,N_19800);
xnor U20062 (N_20062,N_19879,N_19926);
xnor U20063 (N_20063,N_19573,N_19612);
and U20064 (N_20064,N_19902,N_19638);
or U20065 (N_20065,N_19917,N_19934);
nor U20066 (N_20066,N_19894,N_19983);
nand U20067 (N_20067,N_19561,N_19781);
and U20068 (N_20068,N_19985,N_19826);
or U20069 (N_20069,N_19664,N_19889);
xnor U20070 (N_20070,N_19757,N_19803);
nor U20071 (N_20071,N_19635,N_19509);
and U20072 (N_20072,N_19618,N_19546);
nand U20073 (N_20073,N_19545,N_19549);
or U20074 (N_20074,N_19706,N_19571);
nor U20075 (N_20075,N_19719,N_19697);
or U20076 (N_20076,N_19520,N_19625);
xnor U20077 (N_20077,N_19858,N_19932);
xor U20078 (N_20078,N_19574,N_19558);
or U20079 (N_20079,N_19964,N_19687);
nor U20080 (N_20080,N_19938,N_19861);
nor U20081 (N_20081,N_19959,N_19798);
xnor U20082 (N_20082,N_19920,N_19910);
and U20083 (N_20083,N_19551,N_19966);
nand U20084 (N_20084,N_19930,N_19653);
nor U20085 (N_20085,N_19737,N_19544);
or U20086 (N_20086,N_19740,N_19548);
nor U20087 (N_20087,N_19681,N_19890);
nor U20088 (N_20088,N_19998,N_19617);
or U20089 (N_20089,N_19843,N_19824);
or U20090 (N_20090,N_19680,N_19968);
xnor U20091 (N_20091,N_19557,N_19764);
nor U20092 (N_20092,N_19575,N_19988);
nor U20093 (N_20093,N_19846,N_19911);
nor U20094 (N_20094,N_19728,N_19686);
xor U20095 (N_20095,N_19856,N_19517);
or U20096 (N_20096,N_19973,N_19613);
and U20097 (N_20097,N_19822,N_19853);
nand U20098 (N_20098,N_19540,N_19658);
and U20099 (N_20099,N_19980,N_19749);
or U20100 (N_20100,N_19837,N_19699);
or U20101 (N_20101,N_19626,N_19875);
nor U20102 (N_20102,N_19812,N_19935);
and U20103 (N_20103,N_19755,N_19848);
and U20104 (N_20104,N_19510,N_19634);
nor U20105 (N_20105,N_19828,N_19689);
nor U20106 (N_20106,N_19518,N_19915);
nor U20107 (N_20107,N_19691,N_19770);
and U20108 (N_20108,N_19713,N_19904);
nand U20109 (N_20109,N_19807,N_19742);
nor U20110 (N_20110,N_19762,N_19787);
nor U20111 (N_20111,N_19534,N_19640);
xor U20112 (N_20112,N_19784,N_19766);
and U20113 (N_20113,N_19939,N_19541);
xnor U20114 (N_20114,N_19921,N_19992);
and U20115 (N_20115,N_19971,N_19867);
or U20116 (N_20116,N_19565,N_19886);
nand U20117 (N_20117,N_19996,N_19852);
nand U20118 (N_20118,N_19925,N_19704);
nand U20119 (N_20119,N_19765,N_19620);
xnor U20120 (N_20120,N_19778,N_19599);
xor U20121 (N_20121,N_19608,N_19991);
or U20122 (N_20122,N_19604,N_19834);
nand U20123 (N_20123,N_19554,N_19600);
or U20124 (N_20124,N_19842,N_19979);
nor U20125 (N_20125,N_19528,N_19560);
nand U20126 (N_20126,N_19845,N_19590);
nor U20127 (N_20127,N_19919,N_19756);
nor U20128 (N_20128,N_19644,N_19592);
or U20129 (N_20129,N_19532,N_19637);
nand U20130 (N_20130,N_19821,N_19692);
nand U20131 (N_20131,N_19944,N_19987);
nor U20132 (N_20132,N_19907,N_19516);
or U20133 (N_20133,N_19684,N_19825);
or U20134 (N_20134,N_19738,N_19507);
xor U20135 (N_20135,N_19712,N_19502);
nor U20136 (N_20136,N_19639,N_19723);
xor U20137 (N_20137,N_19792,N_19564);
and U20138 (N_20138,N_19504,N_19552);
or U20139 (N_20139,N_19931,N_19593);
or U20140 (N_20140,N_19868,N_19693);
nor U20141 (N_20141,N_19696,N_19808);
nor U20142 (N_20142,N_19885,N_19969);
xnor U20143 (N_20143,N_19777,N_19666);
nor U20144 (N_20144,N_19533,N_19873);
and U20145 (N_20145,N_19927,N_19750);
xnor U20146 (N_20146,N_19993,N_19615);
nand U20147 (N_20147,N_19576,N_19897);
and U20148 (N_20148,N_19623,N_19630);
xnor U20149 (N_20149,N_19535,N_19859);
or U20150 (N_20150,N_19763,N_19947);
and U20151 (N_20151,N_19690,N_19783);
and U20152 (N_20152,N_19501,N_19952);
or U20153 (N_20153,N_19970,N_19795);
nor U20154 (N_20154,N_19536,N_19847);
or U20155 (N_20155,N_19677,N_19515);
xnor U20156 (N_20156,N_19583,N_19611);
or U20157 (N_20157,N_19863,N_19725);
and U20158 (N_20158,N_19759,N_19831);
nand U20159 (N_20159,N_19708,N_19701);
nand U20160 (N_20160,N_19752,N_19522);
nor U20161 (N_20161,N_19711,N_19730);
or U20162 (N_20162,N_19539,N_19570);
nand U20163 (N_20163,N_19585,N_19660);
and U20164 (N_20164,N_19955,N_19595);
nor U20165 (N_20165,N_19773,N_19945);
and U20166 (N_20166,N_19739,N_19526);
nor U20167 (N_20167,N_19978,N_19589);
nor U20168 (N_20168,N_19743,N_19578);
nand U20169 (N_20169,N_19669,N_19789);
and U20170 (N_20170,N_19700,N_19809);
nand U20171 (N_20171,N_19898,N_19601);
and U20172 (N_20172,N_19771,N_19732);
xnor U20173 (N_20173,N_19525,N_19956);
and U20174 (N_20174,N_19559,N_19782);
or U20175 (N_20175,N_19562,N_19695);
xnor U20176 (N_20176,N_19655,N_19500);
or U20177 (N_20177,N_19633,N_19673);
xor U20178 (N_20178,N_19942,N_19871);
xor U20179 (N_20179,N_19627,N_19530);
nor U20180 (N_20180,N_19674,N_19683);
nor U20181 (N_20181,N_19943,N_19796);
nand U20182 (N_20182,N_19513,N_19866);
nand U20183 (N_20183,N_19916,N_19986);
or U20184 (N_20184,N_19550,N_19899);
and U20185 (N_20185,N_19793,N_19818);
or U20186 (N_20186,N_19588,N_19840);
and U20187 (N_20187,N_19913,N_19714);
and U20188 (N_20188,N_19794,N_19758);
nand U20189 (N_20189,N_19901,N_19903);
nand U20190 (N_20190,N_19962,N_19667);
xor U20191 (N_20191,N_19838,N_19523);
nor U20192 (N_20192,N_19616,N_19646);
nand U20193 (N_20193,N_19511,N_19645);
nor U20194 (N_20194,N_19816,N_19914);
or U20195 (N_20195,N_19567,N_19524);
nor U20196 (N_20196,N_19636,N_19878);
nand U20197 (N_20197,N_19941,N_19937);
and U20198 (N_20198,N_19844,N_19997);
nand U20199 (N_20199,N_19741,N_19722);
and U20200 (N_20200,N_19908,N_19688);
and U20201 (N_20201,N_19745,N_19724);
nor U20202 (N_20202,N_19733,N_19650);
nor U20203 (N_20203,N_19984,N_19814);
nor U20204 (N_20204,N_19874,N_19876);
nor U20205 (N_20205,N_19579,N_19836);
and U20206 (N_20206,N_19531,N_19729);
and U20207 (N_20207,N_19751,N_19678);
xor U20208 (N_20208,N_19881,N_19854);
nand U20209 (N_20209,N_19950,N_19802);
nor U20210 (N_20210,N_19989,N_19949);
xor U20211 (N_20211,N_19582,N_19594);
xor U20212 (N_20212,N_19609,N_19965);
nor U20213 (N_20213,N_19882,N_19632);
and U20214 (N_20214,N_19776,N_19715);
xor U20215 (N_20215,N_19591,N_19961);
and U20216 (N_20216,N_19649,N_19521);
xnor U20217 (N_20217,N_19946,N_19841);
xnor U20218 (N_20218,N_19982,N_19731);
or U20219 (N_20219,N_19869,N_19675);
nor U20220 (N_20220,N_19791,N_19734);
or U20221 (N_20221,N_19872,N_19736);
and U20222 (N_20222,N_19747,N_19720);
nor U20223 (N_20223,N_19884,N_19974);
nand U20224 (N_20224,N_19972,N_19893);
or U20225 (N_20225,N_19832,N_19887);
xnor U20226 (N_20226,N_19967,N_19656);
or U20227 (N_20227,N_19538,N_19896);
nand U20228 (N_20228,N_19529,N_19709);
xor U20229 (N_20229,N_19624,N_19610);
nor U20230 (N_20230,N_19827,N_19953);
nor U20231 (N_20231,N_19662,N_19775);
nand U20232 (N_20232,N_19577,N_19888);
and U20233 (N_20233,N_19865,N_19772);
and U20234 (N_20234,N_19753,N_19607);
xnor U20235 (N_20235,N_19855,N_19566);
nor U20236 (N_20236,N_19698,N_19829);
nor U20237 (N_20237,N_19857,N_19514);
nor U20238 (N_20238,N_19975,N_19527);
nand U20239 (N_20239,N_19830,N_19774);
and U20240 (N_20240,N_19556,N_19647);
or U20241 (N_20241,N_19663,N_19643);
or U20242 (N_20242,N_19951,N_19672);
nor U20243 (N_20243,N_19748,N_19665);
or U20244 (N_20244,N_19553,N_19710);
and U20245 (N_20245,N_19716,N_19862);
xor U20246 (N_20246,N_19563,N_19542);
or U20247 (N_20247,N_19661,N_19602);
or U20248 (N_20248,N_19958,N_19981);
xnor U20249 (N_20249,N_19819,N_19651);
and U20250 (N_20250,N_19864,N_19895);
or U20251 (N_20251,N_19861,N_19990);
and U20252 (N_20252,N_19536,N_19969);
nor U20253 (N_20253,N_19569,N_19955);
xor U20254 (N_20254,N_19514,N_19516);
nand U20255 (N_20255,N_19781,N_19664);
and U20256 (N_20256,N_19657,N_19509);
and U20257 (N_20257,N_19671,N_19883);
nor U20258 (N_20258,N_19764,N_19897);
or U20259 (N_20259,N_19646,N_19906);
and U20260 (N_20260,N_19562,N_19977);
or U20261 (N_20261,N_19793,N_19977);
and U20262 (N_20262,N_19967,N_19628);
nand U20263 (N_20263,N_19687,N_19684);
and U20264 (N_20264,N_19791,N_19875);
xnor U20265 (N_20265,N_19739,N_19602);
nor U20266 (N_20266,N_19576,N_19794);
nor U20267 (N_20267,N_19791,N_19845);
nor U20268 (N_20268,N_19568,N_19707);
or U20269 (N_20269,N_19734,N_19717);
or U20270 (N_20270,N_19859,N_19744);
nand U20271 (N_20271,N_19917,N_19604);
nand U20272 (N_20272,N_19835,N_19808);
or U20273 (N_20273,N_19989,N_19570);
nor U20274 (N_20274,N_19524,N_19898);
and U20275 (N_20275,N_19833,N_19716);
nor U20276 (N_20276,N_19790,N_19756);
nand U20277 (N_20277,N_19871,N_19878);
xnor U20278 (N_20278,N_19918,N_19853);
and U20279 (N_20279,N_19721,N_19858);
and U20280 (N_20280,N_19674,N_19760);
nor U20281 (N_20281,N_19627,N_19582);
xor U20282 (N_20282,N_19712,N_19600);
and U20283 (N_20283,N_19840,N_19504);
nor U20284 (N_20284,N_19523,N_19830);
and U20285 (N_20285,N_19597,N_19607);
xor U20286 (N_20286,N_19505,N_19981);
nand U20287 (N_20287,N_19949,N_19919);
xor U20288 (N_20288,N_19528,N_19692);
and U20289 (N_20289,N_19696,N_19703);
nor U20290 (N_20290,N_19549,N_19915);
nand U20291 (N_20291,N_19662,N_19737);
or U20292 (N_20292,N_19678,N_19997);
nand U20293 (N_20293,N_19688,N_19687);
and U20294 (N_20294,N_19634,N_19817);
xor U20295 (N_20295,N_19683,N_19528);
xnor U20296 (N_20296,N_19723,N_19781);
or U20297 (N_20297,N_19822,N_19864);
nand U20298 (N_20298,N_19638,N_19853);
and U20299 (N_20299,N_19540,N_19851);
or U20300 (N_20300,N_19857,N_19837);
nor U20301 (N_20301,N_19992,N_19804);
xor U20302 (N_20302,N_19736,N_19894);
xnor U20303 (N_20303,N_19963,N_19658);
or U20304 (N_20304,N_19920,N_19726);
nand U20305 (N_20305,N_19711,N_19878);
xnor U20306 (N_20306,N_19697,N_19670);
nor U20307 (N_20307,N_19728,N_19648);
or U20308 (N_20308,N_19741,N_19928);
xnor U20309 (N_20309,N_19930,N_19600);
or U20310 (N_20310,N_19855,N_19714);
or U20311 (N_20311,N_19588,N_19984);
xor U20312 (N_20312,N_19974,N_19678);
xor U20313 (N_20313,N_19824,N_19963);
and U20314 (N_20314,N_19841,N_19838);
or U20315 (N_20315,N_19708,N_19780);
nor U20316 (N_20316,N_19587,N_19907);
nor U20317 (N_20317,N_19855,N_19555);
or U20318 (N_20318,N_19909,N_19519);
nand U20319 (N_20319,N_19664,N_19736);
or U20320 (N_20320,N_19562,N_19550);
nand U20321 (N_20321,N_19521,N_19774);
or U20322 (N_20322,N_19624,N_19908);
nor U20323 (N_20323,N_19827,N_19536);
or U20324 (N_20324,N_19771,N_19785);
nand U20325 (N_20325,N_19503,N_19525);
or U20326 (N_20326,N_19656,N_19761);
and U20327 (N_20327,N_19602,N_19685);
or U20328 (N_20328,N_19622,N_19964);
or U20329 (N_20329,N_19881,N_19879);
xnor U20330 (N_20330,N_19796,N_19777);
and U20331 (N_20331,N_19685,N_19628);
and U20332 (N_20332,N_19936,N_19761);
xnor U20333 (N_20333,N_19590,N_19698);
nand U20334 (N_20334,N_19554,N_19503);
xnor U20335 (N_20335,N_19974,N_19805);
or U20336 (N_20336,N_19712,N_19938);
or U20337 (N_20337,N_19638,N_19771);
or U20338 (N_20338,N_19969,N_19857);
or U20339 (N_20339,N_19504,N_19612);
or U20340 (N_20340,N_19788,N_19927);
or U20341 (N_20341,N_19530,N_19669);
or U20342 (N_20342,N_19560,N_19714);
and U20343 (N_20343,N_19574,N_19658);
xor U20344 (N_20344,N_19689,N_19713);
nand U20345 (N_20345,N_19984,N_19679);
nor U20346 (N_20346,N_19604,N_19963);
or U20347 (N_20347,N_19781,N_19726);
nand U20348 (N_20348,N_19579,N_19596);
or U20349 (N_20349,N_19757,N_19828);
or U20350 (N_20350,N_19810,N_19745);
or U20351 (N_20351,N_19868,N_19705);
nor U20352 (N_20352,N_19625,N_19854);
and U20353 (N_20353,N_19852,N_19665);
and U20354 (N_20354,N_19568,N_19769);
nor U20355 (N_20355,N_19554,N_19594);
nor U20356 (N_20356,N_19923,N_19837);
nor U20357 (N_20357,N_19882,N_19854);
nand U20358 (N_20358,N_19515,N_19552);
nor U20359 (N_20359,N_19694,N_19790);
nand U20360 (N_20360,N_19593,N_19923);
nor U20361 (N_20361,N_19541,N_19659);
xor U20362 (N_20362,N_19711,N_19938);
nor U20363 (N_20363,N_19670,N_19761);
or U20364 (N_20364,N_19503,N_19527);
nand U20365 (N_20365,N_19603,N_19870);
or U20366 (N_20366,N_19585,N_19829);
or U20367 (N_20367,N_19501,N_19546);
nor U20368 (N_20368,N_19781,N_19710);
or U20369 (N_20369,N_19868,N_19676);
and U20370 (N_20370,N_19500,N_19669);
nor U20371 (N_20371,N_19747,N_19714);
nor U20372 (N_20372,N_19672,N_19697);
xnor U20373 (N_20373,N_19990,N_19628);
nand U20374 (N_20374,N_19829,N_19893);
xor U20375 (N_20375,N_19958,N_19866);
nor U20376 (N_20376,N_19533,N_19881);
nor U20377 (N_20377,N_19545,N_19785);
nor U20378 (N_20378,N_19842,N_19852);
nor U20379 (N_20379,N_19659,N_19502);
xor U20380 (N_20380,N_19518,N_19896);
nor U20381 (N_20381,N_19697,N_19626);
and U20382 (N_20382,N_19861,N_19716);
xor U20383 (N_20383,N_19595,N_19968);
nor U20384 (N_20384,N_19795,N_19631);
xor U20385 (N_20385,N_19819,N_19598);
or U20386 (N_20386,N_19864,N_19980);
and U20387 (N_20387,N_19826,N_19627);
xor U20388 (N_20388,N_19889,N_19577);
nand U20389 (N_20389,N_19706,N_19928);
or U20390 (N_20390,N_19692,N_19951);
xnor U20391 (N_20391,N_19857,N_19505);
nor U20392 (N_20392,N_19929,N_19990);
xor U20393 (N_20393,N_19976,N_19615);
or U20394 (N_20394,N_19679,N_19632);
and U20395 (N_20395,N_19890,N_19772);
xor U20396 (N_20396,N_19563,N_19727);
xnor U20397 (N_20397,N_19791,N_19608);
xnor U20398 (N_20398,N_19788,N_19708);
and U20399 (N_20399,N_19627,N_19905);
or U20400 (N_20400,N_19667,N_19848);
nor U20401 (N_20401,N_19971,N_19876);
or U20402 (N_20402,N_19585,N_19864);
nor U20403 (N_20403,N_19687,N_19531);
and U20404 (N_20404,N_19618,N_19762);
nor U20405 (N_20405,N_19967,N_19832);
nand U20406 (N_20406,N_19638,N_19580);
xnor U20407 (N_20407,N_19574,N_19503);
nand U20408 (N_20408,N_19751,N_19591);
nor U20409 (N_20409,N_19792,N_19917);
and U20410 (N_20410,N_19578,N_19525);
or U20411 (N_20411,N_19753,N_19543);
or U20412 (N_20412,N_19971,N_19824);
or U20413 (N_20413,N_19608,N_19816);
xor U20414 (N_20414,N_19807,N_19685);
or U20415 (N_20415,N_19717,N_19868);
xor U20416 (N_20416,N_19558,N_19821);
nand U20417 (N_20417,N_19507,N_19581);
nor U20418 (N_20418,N_19976,N_19732);
and U20419 (N_20419,N_19571,N_19805);
and U20420 (N_20420,N_19569,N_19522);
or U20421 (N_20421,N_19620,N_19913);
nor U20422 (N_20422,N_19503,N_19694);
xnor U20423 (N_20423,N_19842,N_19965);
nor U20424 (N_20424,N_19942,N_19729);
nor U20425 (N_20425,N_19953,N_19741);
nand U20426 (N_20426,N_19897,N_19680);
nor U20427 (N_20427,N_19671,N_19641);
or U20428 (N_20428,N_19814,N_19592);
nor U20429 (N_20429,N_19761,N_19573);
or U20430 (N_20430,N_19920,N_19764);
xnor U20431 (N_20431,N_19882,N_19711);
or U20432 (N_20432,N_19782,N_19934);
nor U20433 (N_20433,N_19644,N_19544);
xor U20434 (N_20434,N_19579,N_19545);
or U20435 (N_20435,N_19559,N_19508);
nor U20436 (N_20436,N_19617,N_19991);
nand U20437 (N_20437,N_19609,N_19572);
or U20438 (N_20438,N_19677,N_19798);
xor U20439 (N_20439,N_19685,N_19730);
and U20440 (N_20440,N_19920,N_19542);
xor U20441 (N_20441,N_19542,N_19858);
and U20442 (N_20442,N_19850,N_19639);
or U20443 (N_20443,N_19519,N_19849);
nand U20444 (N_20444,N_19774,N_19784);
xnor U20445 (N_20445,N_19679,N_19544);
xor U20446 (N_20446,N_19914,N_19674);
nand U20447 (N_20447,N_19688,N_19830);
xor U20448 (N_20448,N_19937,N_19513);
and U20449 (N_20449,N_19716,N_19548);
or U20450 (N_20450,N_19958,N_19556);
and U20451 (N_20451,N_19948,N_19526);
nand U20452 (N_20452,N_19817,N_19800);
and U20453 (N_20453,N_19719,N_19938);
or U20454 (N_20454,N_19572,N_19975);
or U20455 (N_20455,N_19961,N_19603);
and U20456 (N_20456,N_19640,N_19713);
and U20457 (N_20457,N_19902,N_19599);
xnor U20458 (N_20458,N_19693,N_19501);
and U20459 (N_20459,N_19974,N_19511);
xnor U20460 (N_20460,N_19567,N_19741);
and U20461 (N_20461,N_19805,N_19676);
or U20462 (N_20462,N_19872,N_19942);
nand U20463 (N_20463,N_19985,N_19549);
or U20464 (N_20464,N_19957,N_19982);
xnor U20465 (N_20465,N_19962,N_19934);
nand U20466 (N_20466,N_19964,N_19847);
nor U20467 (N_20467,N_19816,N_19858);
nor U20468 (N_20468,N_19616,N_19545);
xnor U20469 (N_20469,N_19745,N_19705);
nand U20470 (N_20470,N_19631,N_19769);
or U20471 (N_20471,N_19730,N_19649);
xnor U20472 (N_20472,N_19986,N_19688);
or U20473 (N_20473,N_19668,N_19907);
and U20474 (N_20474,N_19807,N_19646);
nor U20475 (N_20475,N_19937,N_19759);
nand U20476 (N_20476,N_19710,N_19612);
or U20477 (N_20477,N_19903,N_19730);
and U20478 (N_20478,N_19622,N_19812);
nand U20479 (N_20479,N_19571,N_19845);
xnor U20480 (N_20480,N_19788,N_19844);
xnor U20481 (N_20481,N_19616,N_19989);
xnor U20482 (N_20482,N_19866,N_19947);
xnor U20483 (N_20483,N_19948,N_19742);
xor U20484 (N_20484,N_19881,N_19802);
nand U20485 (N_20485,N_19697,N_19764);
xnor U20486 (N_20486,N_19997,N_19707);
xor U20487 (N_20487,N_19912,N_19712);
xor U20488 (N_20488,N_19635,N_19520);
or U20489 (N_20489,N_19796,N_19576);
nand U20490 (N_20490,N_19850,N_19828);
xor U20491 (N_20491,N_19539,N_19947);
nand U20492 (N_20492,N_19611,N_19898);
or U20493 (N_20493,N_19710,N_19645);
nand U20494 (N_20494,N_19537,N_19617);
and U20495 (N_20495,N_19707,N_19797);
and U20496 (N_20496,N_19506,N_19626);
or U20497 (N_20497,N_19696,N_19660);
or U20498 (N_20498,N_19544,N_19508);
nand U20499 (N_20499,N_19756,N_19773);
nor U20500 (N_20500,N_20317,N_20009);
nand U20501 (N_20501,N_20000,N_20087);
and U20502 (N_20502,N_20246,N_20236);
xnor U20503 (N_20503,N_20218,N_20485);
and U20504 (N_20504,N_20135,N_20415);
or U20505 (N_20505,N_20037,N_20184);
or U20506 (N_20506,N_20042,N_20044);
xnor U20507 (N_20507,N_20123,N_20142);
and U20508 (N_20508,N_20180,N_20474);
nand U20509 (N_20509,N_20328,N_20083);
and U20510 (N_20510,N_20105,N_20173);
xnor U20511 (N_20511,N_20378,N_20162);
xnor U20512 (N_20512,N_20024,N_20472);
xor U20513 (N_20513,N_20279,N_20023);
nand U20514 (N_20514,N_20071,N_20106);
xor U20515 (N_20515,N_20159,N_20222);
and U20516 (N_20516,N_20278,N_20225);
or U20517 (N_20517,N_20147,N_20059);
or U20518 (N_20518,N_20302,N_20019);
or U20519 (N_20519,N_20092,N_20285);
nor U20520 (N_20520,N_20273,N_20304);
nand U20521 (N_20521,N_20397,N_20340);
and U20522 (N_20522,N_20205,N_20161);
nand U20523 (N_20523,N_20309,N_20363);
nor U20524 (N_20524,N_20155,N_20371);
and U20525 (N_20525,N_20431,N_20082);
xnor U20526 (N_20526,N_20212,N_20081);
nand U20527 (N_20527,N_20034,N_20254);
or U20528 (N_20528,N_20354,N_20428);
xor U20529 (N_20529,N_20330,N_20463);
and U20530 (N_20530,N_20005,N_20269);
nor U20531 (N_20531,N_20169,N_20311);
xnor U20532 (N_20532,N_20191,N_20442);
xnor U20533 (N_20533,N_20366,N_20220);
and U20534 (N_20534,N_20486,N_20174);
nand U20535 (N_20535,N_20310,N_20255);
nor U20536 (N_20536,N_20404,N_20445);
nor U20537 (N_20537,N_20067,N_20425);
xor U20538 (N_20538,N_20275,N_20150);
xor U20539 (N_20539,N_20251,N_20232);
or U20540 (N_20540,N_20239,N_20259);
nand U20541 (N_20541,N_20429,N_20073);
or U20542 (N_20542,N_20414,N_20406);
xnor U20543 (N_20543,N_20271,N_20393);
or U20544 (N_20544,N_20226,N_20030);
or U20545 (N_20545,N_20033,N_20470);
xor U20546 (N_20546,N_20158,N_20266);
nand U20547 (N_20547,N_20095,N_20375);
and U20548 (N_20548,N_20418,N_20412);
nand U20549 (N_20549,N_20336,N_20010);
nor U20550 (N_20550,N_20111,N_20172);
nand U20551 (N_20551,N_20368,N_20417);
and U20552 (N_20552,N_20286,N_20408);
nor U20553 (N_20553,N_20139,N_20282);
xnor U20554 (N_20554,N_20197,N_20211);
xnor U20555 (N_20555,N_20333,N_20396);
or U20556 (N_20556,N_20316,N_20342);
and U20557 (N_20557,N_20413,N_20138);
and U20558 (N_20558,N_20498,N_20313);
xnor U20559 (N_20559,N_20410,N_20475);
nand U20560 (N_20560,N_20433,N_20101);
nand U20561 (N_20561,N_20258,N_20494);
xnor U20562 (N_20562,N_20039,N_20061);
and U20563 (N_20563,N_20055,N_20458);
or U20564 (N_20564,N_20341,N_20054);
and U20565 (N_20565,N_20427,N_20240);
or U20566 (N_20566,N_20160,N_20253);
and U20567 (N_20567,N_20086,N_20124);
and U20568 (N_20568,N_20379,N_20383);
xor U20569 (N_20569,N_20080,N_20227);
nand U20570 (N_20570,N_20104,N_20306);
and U20571 (N_20571,N_20457,N_20489);
and U20572 (N_20572,N_20261,N_20423);
and U20573 (N_20573,N_20060,N_20373);
nand U20574 (N_20574,N_20399,N_20032);
and U20575 (N_20575,N_20112,N_20108);
nor U20576 (N_20576,N_20134,N_20116);
and U20577 (N_20577,N_20177,N_20130);
or U20578 (N_20578,N_20094,N_20045);
and U20579 (N_20579,N_20362,N_20332);
nor U20580 (N_20580,N_20281,N_20435);
nor U20581 (N_20581,N_20078,N_20143);
xor U20582 (N_20582,N_20293,N_20451);
nor U20583 (N_20583,N_20127,N_20051);
and U20584 (N_20584,N_20292,N_20125);
or U20585 (N_20585,N_20265,N_20247);
xnor U20586 (N_20586,N_20439,N_20385);
nor U20587 (N_20587,N_20478,N_20016);
nand U20588 (N_20588,N_20062,N_20327);
nor U20589 (N_20589,N_20074,N_20483);
xor U20590 (N_20590,N_20499,N_20260);
nand U20591 (N_20591,N_20455,N_20091);
and U20592 (N_20592,N_20424,N_20201);
nand U20593 (N_20593,N_20118,N_20047);
xor U20594 (N_20594,N_20352,N_20441);
and U20595 (N_20595,N_20377,N_20331);
nand U20596 (N_20596,N_20031,N_20440);
and U20597 (N_20597,N_20338,N_20299);
xor U20598 (N_20598,N_20107,N_20202);
and U20599 (N_20599,N_20267,N_20314);
xor U20600 (N_20600,N_20013,N_20443);
or U20601 (N_20601,N_20221,N_20121);
nand U20602 (N_20602,N_20097,N_20450);
or U20603 (N_20603,N_20151,N_20264);
nand U20604 (N_20604,N_20464,N_20113);
and U20605 (N_20605,N_20098,N_20228);
and U20606 (N_20606,N_20492,N_20318);
or U20607 (N_20607,N_20168,N_20294);
nand U20608 (N_20608,N_20493,N_20387);
nand U20609 (N_20609,N_20350,N_20004);
xor U20610 (N_20610,N_20276,N_20416);
and U20611 (N_20611,N_20145,N_20308);
xnor U20612 (N_20612,N_20206,N_20163);
or U20613 (N_20613,N_20181,N_20358);
nand U20614 (N_20614,N_20085,N_20049);
nand U20615 (N_20615,N_20153,N_20344);
nand U20616 (N_20616,N_20346,N_20021);
xnor U20617 (N_20617,N_20190,N_20167);
nor U20618 (N_20618,N_20224,N_20223);
and U20619 (N_20619,N_20364,N_20090);
nand U20620 (N_20620,N_20403,N_20136);
and U20621 (N_20621,N_20057,N_20434);
nand U20622 (N_20622,N_20476,N_20388);
nor U20623 (N_20623,N_20217,N_20233);
xor U20624 (N_20624,N_20148,N_20384);
or U20625 (N_20625,N_20178,N_20242);
nand U20626 (N_20626,N_20459,N_20015);
or U20627 (N_20627,N_20132,N_20337);
and U20628 (N_20628,N_20003,N_20192);
nand U20629 (N_20629,N_20183,N_20409);
nand U20630 (N_20630,N_20133,N_20072);
xnor U20631 (N_20631,N_20329,N_20088);
and U20632 (N_20632,N_20323,N_20100);
or U20633 (N_20633,N_20477,N_20198);
nand U20634 (N_20634,N_20149,N_20001);
or U20635 (N_20635,N_20339,N_20256);
nand U20636 (N_20636,N_20126,N_20252);
xor U20637 (N_20637,N_20166,N_20165);
xor U20638 (N_20638,N_20011,N_20157);
or U20639 (N_20639,N_20374,N_20050);
nor U20640 (N_20640,N_20064,N_20482);
xor U20641 (N_20641,N_20320,N_20018);
xor U20642 (N_20642,N_20322,N_20186);
nand U20643 (N_20643,N_20296,N_20381);
nand U20644 (N_20644,N_20065,N_20480);
and U20645 (N_20645,N_20359,N_20263);
nor U20646 (N_20646,N_20356,N_20208);
or U20647 (N_20647,N_20012,N_20093);
or U20648 (N_20648,N_20204,N_20456);
nor U20649 (N_20649,N_20250,N_20146);
nor U20650 (N_20650,N_20115,N_20481);
nand U20651 (N_20651,N_20283,N_20070);
nand U20652 (N_20652,N_20029,N_20182);
nand U20653 (N_20653,N_20386,N_20128);
or U20654 (N_20654,N_20119,N_20069);
xor U20655 (N_20655,N_20426,N_20324);
or U20656 (N_20656,N_20196,N_20193);
nand U20657 (N_20657,N_20466,N_20484);
nand U20658 (N_20658,N_20230,N_20297);
xor U20659 (N_20659,N_20195,N_20468);
or U20660 (N_20660,N_20170,N_20084);
nor U20661 (N_20661,N_20274,N_20432);
nand U20662 (N_20662,N_20262,N_20076);
xnor U20663 (N_20663,N_20141,N_20056);
xor U20664 (N_20664,N_20448,N_20453);
nand U20665 (N_20665,N_20401,N_20089);
nor U20666 (N_20666,N_20040,N_20214);
or U20667 (N_20667,N_20353,N_20194);
nor U20668 (N_20668,N_20215,N_20248);
or U20669 (N_20669,N_20312,N_20140);
nand U20670 (N_20670,N_20244,N_20238);
and U20671 (N_20671,N_20473,N_20209);
nor U20672 (N_20672,N_20436,N_20210);
and U20673 (N_20673,N_20411,N_20277);
nand U20674 (N_20674,N_20355,N_20131);
nand U20675 (N_20675,N_20447,N_20245);
and U20676 (N_20676,N_20200,N_20430);
nor U20677 (N_20677,N_20175,N_20300);
or U20678 (N_20678,N_20488,N_20452);
xor U20679 (N_20679,N_20156,N_20189);
and U20680 (N_20680,N_20291,N_20025);
xor U20681 (N_20681,N_20325,N_20203);
nor U20682 (N_20682,N_20400,N_20438);
xor U20683 (N_20683,N_20096,N_20380);
and U20684 (N_20684,N_20022,N_20219);
and U20685 (N_20685,N_20122,N_20491);
or U20686 (N_20686,N_20303,N_20129);
nand U20687 (N_20687,N_20407,N_20079);
and U20688 (N_20688,N_20063,N_20068);
nand U20689 (N_20689,N_20053,N_20361);
xor U20690 (N_20690,N_20365,N_20421);
nand U20691 (N_20691,N_20465,N_20347);
xnor U20692 (N_20692,N_20027,N_20467);
xor U20693 (N_20693,N_20351,N_20295);
and U20694 (N_20694,N_20036,N_20046);
and U20695 (N_20695,N_20497,N_20114);
nand U20696 (N_20696,N_20028,N_20237);
xor U20697 (N_20697,N_20301,N_20234);
nand U20698 (N_20698,N_20020,N_20179);
xor U20699 (N_20699,N_20349,N_20176);
or U20700 (N_20700,N_20469,N_20307);
and U20701 (N_20701,N_20287,N_20376);
nor U20702 (N_20702,N_20315,N_20462);
and U20703 (N_20703,N_20479,N_20357);
or U20704 (N_20704,N_20343,N_20437);
nor U20705 (N_20705,N_20284,N_20335);
and U20706 (N_20706,N_20490,N_20471);
nor U20707 (N_20707,N_20394,N_20035);
nand U20708 (N_20708,N_20213,N_20187);
nand U20709 (N_20709,N_20099,N_20395);
and U20710 (N_20710,N_20372,N_20109);
or U20711 (N_20711,N_20444,N_20334);
nand U20712 (N_20712,N_20446,N_20058);
or U20713 (N_20713,N_20229,N_20017);
or U20714 (N_20714,N_20243,N_20268);
xnor U20715 (N_20715,N_20152,N_20137);
and U20716 (N_20716,N_20487,N_20495);
xor U20717 (N_20717,N_20120,N_20185);
nand U20718 (N_20718,N_20241,N_20207);
and U20719 (N_20719,N_20454,N_20345);
nor U20720 (N_20720,N_20402,N_20103);
or U20721 (N_20721,N_20280,N_20370);
and U20722 (N_20722,N_20461,N_20272);
and U20723 (N_20723,N_20171,N_20290);
and U20724 (N_20724,N_20043,N_20270);
or U20725 (N_20725,N_20188,N_20382);
xor U20726 (N_20726,N_20367,N_20360);
nand U20727 (N_20727,N_20392,N_20038);
and U20728 (N_20728,N_20231,N_20117);
xnor U20729 (N_20729,N_20389,N_20144);
or U20730 (N_20730,N_20420,N_20216);
or U20731 (N_20731,N_20041,N_20199);
nand U20732 (N_20732,N_20026,N_20289);
or U20733 (N_20733,N_20321,N_20419);
xor U20734 (N_20734,N_20288,N_20102);
or U20735 (N_20735,N_20002,N_20066);
nand U20736 (N_20736,N_20348,N_20075);
and U20737 (N_20737,N_20422,N_20235);
xnor U20738 (N_20738,N_20164,N_20154);
nor U20739 (N_20739,N_20449,N_20369);
and U20740 (N_20740,N_20326,N_20496);
xnor U20741 (N_20741,N_20007,N_20014);
nor U20742 (N_20742,N_20249,N_20319);
or U20743 (N_20743,N_20460,N_20257);
nor U20744 (N_20744,N_20006,N_20305);
and U20745 (N_20745,N_20077,N_20048);
nand U20746 (N_20746,N_20390,N_20008);
and U20747 (N_20747,N_20405,N_20052);
nand U20748 (N_20748,N_20110,N_20391);
nor U20749 (N_20749,N_20298,N_20398);
xnor U20750 (N_20750,N_20045,N_20314);
nor U20751 (N_20751,N_20315,N_20302);
nor U20752 (N_20752,N_20247,N_20274);
or U20753 (N_20753,N_20178,N_20449);
or U20754 (N_20754,N_20275,N_20270);
and U20755 (N_20755,N_20199,N_20371);
xor U20756 (N_20756,N_20465,N_20471);
and U20757 (N_20757,N_20396,N_20188);
nor U20758 (N_20758,N_20049,N_20475);
xnor U20759 (N_20759,N_20001,N_20025);
and U20760 (N_20760,N_20212,N_20322);
or U20761 (N_20761,N_20005,N_20075);
nor U20762 (N_20762,N_20263,N_20020);
and U20763 (N_20763,N_20128,N_20209);
and U20764 (N_20764,N_20047,N_20398);
xor U20765 (N_20765,N_20482,N_20180);
nor U20766 (N_20766,N_20279,N_20291);
and U20767 (N_20767,N_20310,N_20033);
or U20768 (N_20768,N_20151,N_20338);
xnor U20769 (N_20769,N_20359,N_20188);
nand U20770 (N_20770,N_20459,N_20109);
or U20771 (N_20771,N_20269,N_20482);
or U20772 (N_20772,N_20081,N_20481);
xor U20773 (N_20773,N_20181,N_20354);
nand U20774 (N_20774,N_20209,N_20378);
or U20775 (N_20775,N_20494,N_20110);
or U20776 (N_20776,N_20436,N_20488);
and U20777 (N_20777,N_20192,N_20410);
and U20778 (N_20778,N_20175,N_20255);
xnor U20779 (N_20779,N_20324,N_20046);
nor U20780 (N_20780,N_20496,N_20260);
and U20781 (N_20781,N_20180,N_20017);
nor U20782 (N_20782,N_20219,N_20344);
and U20783 (N_20783,N_20420,N_20456);
or U20784 (N_20784,N_20234,N_20193);
nand U20785 (N_20785,N_20376,N_20286);
or U20786 (N_20786,N_20089,N_20212);
nor U20787 (N_20787,N_20234,N_20318);
xor U20788 (N_20788,N_20395,N_20251);
nand U20789 (N_20789,N_20237,N_20202);
xor U20790 (N_20790,N_20260,N_20469);
nand U20791 (N_20791,N_20096,N_20204);
and U20792 (N_20792,N_20210,N_20483);
or U20793 (N_20793,N_20271,N_20273);
or U20794 (N_20794,N_20456,N_20492);
or U20795 (N_20795,N_20449,N_20114);
nor U20796 (N_20796,N_20306,N_20417);
nor U20797 (N_20797,N_20064,N_20024);
or U20798 (N_20798,N_20103,N_20398);
and U20799 (N_20799,N_20151,N_20123);
and U20800 (N_20800,N_20371,N_20461);
xnor U20801 (N_20801,N_20059,N_20445);
nand U20802 (N_20802,N_20475,N_20255);
and U20803 (N_20803,N_20404,N_20268);
or U20804 (N_20804,N_20456,N_20467);
nor U20805 (N_20805,N_20217,N_20066);
nand U20806 (N_20806,N_20367,N_20331);
xor U20807 (N_20807,N_20058,N_20440);
xor U20808 (N_20808,N_20261,N_20183);
nor U20809 (N_20809,N_20273,N_20496);
xor U20810 (N_20810,N_20363,N_20299);
and U20811 (N_20811,N_20306,N_20161);
nor U20812 (N_20812,N_20219,N_20135);
or U20813 (N_20813,N_20045,N_20461);
or U20814 (N_20814,N_20265,N_20191);
or U20815 (N_20815,N_20424,N_20471);
xor U20816 (N_20816,N_20064,N_20065);
or U20817 (N_20817,N_20238,N_20012);
nand U20818 (N_20818,N_20141,N_20499);
xor U20819 (N_20819,N_20445,N_20238);
or U20820 (N_20820,N_20251,N_20279);
nand U20821 (N_20821,N_20255,N_20165);
nor U20822 (N_20822,N_20467,N_20157);
or U20823 (N_20823,N_20272,N_20485);
nor U20824 (N_20824,N_20108,N_20262);
nand U20825 (N_20825,N_20460,N_20222);
xor U20826 (N_20826,N_20191,N_20039);
or U20827 (N_20827,N_20024,N_20422);
or U20828 (N_20828,N_20336,N_20404);
xnor U20829 (N_20829,N_20226,N_20083);
nand U20830 (N_20830,N_20072,N_20078);
and U20831 (N_20831,N_20286,N_20167);
or U20832 (N_20832,N_20039,N_20343);
and U20833 (N_20833,N_20265,N_20015);
xnor U20834 (N_20834,N_20492,N_20164);
and U20835 (N_20835,N_20445,N_20488);
and U20836 (N_20836,N_20490,N_20208);
nand U20837 (N_20837,N_20459,N_20439);
xnor U20838 (N_20838,N_20079,N_20242);
nor U20839 (N_20839,N_20101,N_20088);
nor U20840 (N_20840,N_20189,N_20261);
and U20841 (N_20841,N_20135,N_20345);
nand U20842 (N_20842,N_20435,N_20182);
and U20843 (N_20843,N_20223,N_20410);
nor U20844 (N_20844,N_20434,N_20047);
nand U20845 (N_20845,N_20364,N_20203);
or U20846 (N_20846,N_20455,N_20181);
nand U20847 (N_20847,N_20108,N_20339);
xnor U20848 (N_20848,N_20185,N_20341);
xnor U20849 (N_20849,N_20287,N_20155);
xnor U20850 (N_20850,N_20393,N_20048);
nor U20851 (N_20851,N_20466,N_20067);
or U20852 (N_20852,N_20383,N_20205);
or U20853 (N_20853,N_20359,N_20067);
and U20854 (N_20854,N_20016,N_20094);
nand U20855 (N_20855,N_20102,N_20449);
xor U20856 (N_20856,N_20173,N_20078);
nor U20857 (N_20857,N_20332,N_20100);
xor U20858 (N_20858,N_20090,N_20108);
and U20859 (N_20859,N_20198,N_20080);
and U20860 (N_20860,N_20409,N_20456);
and U20861 (N_20861,N_20368,N_20311);
or U20862 (N_20862,N_20291,N_20326);
and U20863 (N_20863,N_20103,N_20373);
and U20864 (N_20864,N_20468,N_20102);
or U20865 (N_20865,N_20304,N_20193);
and U20866 (N_20866,N_20464,N_20454);
and U20867 (N_20867,N_20085,N_20415);
or U20868 (N_20868,N_20428,N_20067);
nand U20869 (N_20869,N_20393,N_20403);
nand U20870 (N_20870,N_20099,N_20163);
and U20871 (N_20871,N_20186,N_20060);
xnor U20872 (N_20872,N_20097,N_20113);
nor U20873 (N_20873,N_20093,N_20008);
or U20874 (N_20874,N_20437,N_20079);
nand U20875 (N_20875,N_20286,N_20382);
xor U20876 (N_20876,N_20295,N_20262);
and U20877 (N_20877,N_20300,N_20186);
or U20878 (N_20878,N_20330,N_20018);
or U20879 (N_20879,N_20194,N_20027);
nand U20880 (N_20880,N_20069,N_20202);
nor U20881 (N_20881,N_20221,N_20095);
and U20882 (N_20882,N_20395,N_20063);
nand U20883 (N_20883,N_20412,N_20058);
nand U20884 (N_20884,N_20038,N_20215);
nor U20885 (N_20885,N_20012,N_20280);
xnor U20886 (N_20886,N_20145,N_20111);
and U20887 (N_20887,N_20456,N_20237);
nand U20888 (N_20888,N_20300,N_20377);
and U20889 (N_20889,N_20285,N_20039);
and U20890 (N_20890,N_20447,N_20478);
nand U20891 (N_20891,N_20101,N_20238);
nor U20892 (N_20892,N_20426,N_20150);
or U20893 (N_20893,N_20466,N_20132);
xor U20894 (N_20894,N_20497,N_20063);
xor U20895 (N_20895,N_20076,N_20093);
or U20896 (N_20896,N_20124,N_20352);
nor U20897 (N_20897,N_20050,N_20446);
and U20898 (N_20898,N_20291,N_20163);
nand U20899 (N_20899,N_20168,N_20077);
and U20900 (N_20900,N_20450,N_20398);
or U20901 (N_20901,N_20386,N_20387);
and U20902 (N_20902,N_20339,N_20059);
nor U20903 (N_20903,N_20147,N_20463);
or U20904 (N_20904,N_20488,N_20208);
nor U20905 (N_20905,N_20359,N_20400);
nand U20906 (N_20906,N_20286,N_20103);
xnor U20907 (N_20907,N_20080,N_20335);
xnor U20908 (N_20908,N_20068,N_20091);
or U20909 (N_20909,N_20149,N_20287);
and U20910 (N_20910,N_20464,N_20166);
nor U20911 (N_20911,N_20144,N_20087);
xor U20912 (N_20912,N_20083,N_20113);
nand U20913 (N_20913,N_20443,N_20065);
and U20914 (N_20914,N_20488,N_20205);
xnor U20915 (N_20915,N_20294,N_20008);
and U20916 (N_20916,N_20422,N_20492);
and U20917 (N_20917,N_20180,N_20095);
nor U20918 (N_20918,N_20231,N_20334);
xnor U20919 (N_20919,N_20127,N_20193);
or U20920 (N_20920,N_20267,N_20260);
nand U20921 (N_20921,N_20310,N_20114);
and U20922 (N_20922,N_20443,N_20166);
xor U20923 (N_20923,N_20036,N_20467);
and U20924 (N_20924,N_20479,N_20306);
nor U20925 (N_20925,N_20011,N_20160);
nand U20926 (N_20926,N_20274,N_20123);
nor U20927 (N_20927,N_20290,N_20031);
or U20928 (N_20928,N_20002,N_20319);
or U20929 (N_20929,N_20344,N_20455);
nor U20930 (N_20930,N_20380,N_20238);
xnor U20931 (N_20931,N_20323,N_20471);
and U20932 (N_20932,N_20320,N_20447);
nand U20933 (N_20933,N_20309,N_20343);
nor U20934 (N_20934,N_20461,N_20319);
nand U20935 (N_20935,N_20154,N_20424);
or U20936 (N_20936,N_20346,N_20341);
or U20937 (N_20937,N_20195,N_20056);
xnor U20938 (N_20938,N_20085,N_20379);
nand U20939 (N_20939,N_20431,N_20484);
nor U20940 (N_20940,N_20106,N_20037);
xnor U20941 (N_20941,N_20318,N_20449);
xnor U20942 (N_20942,N_20350,N_20139);
nand U20943 (N_20943,N_20239,N_20201);
nand U20944 (N_20944,N_20385,N_20321);
xor U20945 (N_20945,N_20403,N_20329);
xnor U20946 (N_20946,N_20102,N_20214);
nand U20947 (N_20947,N_20459,N_20461);
xnor U20948 (N_20948,N_20498,N_20346);
nand U20949 (N_20949,N_20321,N_20004);
and U20950 (N_20950,N_20116,N_20280);
and U20951 (N_20951,N_20061,N_20366);
xor U20952 (N_20952,N_20217,N_20353);
or U20953 (N_20953,N_20047,N_20399);
and U20954 (N_20954,N_20008,N_20097);
nand U20955 (N_20955,N_20275,N_20162);
or U20956 (N_20956,N_20004,N_20449);
xor U20957 (N_20957,N_20370,N_20354);
and U20958 (N_20958,N_20016,N_20233);
nand U20959 (N_20959,N_20441,N_20467);
nor U20960 (N_20960,N_20495,N_20277);
or U20961 (N_20961,N_20305,N_20224);
nor U20962 (N_20962,N_20021,N_20312);
or U20963 (N_20963,N_20028,N_20209);
and U20964 (N_20964,N_20480,N_20189);
nor U20965 (N_20965,N_20029,N_20220);
nor U20966 (N_20966,N_20200,N_20215);
nor U20967 (N_20967,N_20361,N_20415);
nand U20968 (N_20968,N_20311,N_20315);
nor U20969 (N_20969,N_20175,N_20080);
xnor U20970 (N_20970,N_20047,N_20269);
nand U20971 (N_20971,N_20073,N_20045);
xor U20972 (N_20972,N_20479,N_20047);
or U20973 (N_20973,N_20298,N_20138);
nor U20974 (N_20974,N_20056,N_20167);
nand U20975 (N_20975,N_20039,N_20437);
and U20976 (N_20976,N_20187,N_20417);
or U20977 (N_20977,N_20026,N_20059);
or U20978 (N_20978,N_20087,N_20269);
nor U20979 (N_20979,N_20234,N_20368);
and U20980 (N_20980,N_20322,N_20377);
nand U20981 (N_20981,N_20479,N_20120);
nor U20982 (N_20982,N_20293,N_20005);
or U20983 (N_20983,N_20428,N_20158);
nor U20984 (N_20984,N_20347,N_20135);
nor U20985 (N_20985,N_20375,N_20120);
or U20986 (N_20986,N_20480,N_20022);
or U20987 (N_20987,N_20240,N_20213);
or U20988 (N_20988,N_20038,N_20293);
nand U20989 (N_20989,N_20341,N_20452);
xnor U20990 (N_20990,N_20476,N_20173);
or U20991 (N_20991,N_20400,N_20467);
xnor U20992 (N_20992,N_20041,N_20461);
and U20993 (N_20993,N_20453,N_20272);
nand U20994 (N_20994,N_20475,N_20160);
or U20995 (N_20995,N_20216,N_20181);
or U20996 (N_20996,N_20309,N_20176);
nand U20997 (N_20997,N_20349,N_20240);
or U20998 (N_20998,N_20231,N_20023);
nand U20999 (N_20999,N_20476,N_20147);
nand U21000 (N_21000,N_20554,N_20592);
nand U21001 (N_21001,N_20612,N_20782);
nor U21002 (N_21002,N_20688,N_20527);
and U21003 (N_21003,N_20936,N_20606);
and U21004 (N_21004,N_20698,N_20506);
and U21005 (N_21005,N_20515,N_20779);
nor U21006 (N_21006,N_20574,N_20796);
nand U21007 (N_21007,N_20602,N_20898);
nand U21008 (N_21008,N_20939,N_20847);
nand U21009 (N_21009,N_20586,N_20593);
or U21010 (N_21010,N_20821,N_20626);
or U21011 (N_21011,N_20690,N_20599);
or U21012 (N_21012,N_20518,N_20851);
nand U21013 (N_21013,N_20906,N_20877);
and U21014 (N_21014,N_20846,N_20883);
xnor U21015 (N_21015,N_20604,N_20733);
or U21016 (N_21016,N_20943,N_20930);
xnor U21017 (N_21017,N_20966,N_20650);
nor U21018 (N_21018,N_20844,N_20820);
nor U21019 (N_21019,N_20721,N_20636);
xnor U21020 (N_21020,N_20984,N_20584);
xnor U21021 (N_21021,N_20717,N_20627);
nand U21022 (N_21022,N_20770,N_20551);
xor U21023 (N_21023,N_20925,N_20826);
nand U21024 (N_21024,N_20855,N_20668);
or U21025 (N_21025,N_20525,N_20780);
xor U21026 (N_21026,N_20817,N_20608);
nand U21027 (N_21027,N_20792,N_20736);
xor U21028 (N_21028,N_20601,N_20511);
xnor U21029 (N_21029,N_20856,N_20932);
or U21030 (N_21030,N_20542,N_20622);
and U21031 (N_21031,N_20617,N_20910);
or U21032 (N_21032,N_20922,N_20789);
and U21033 (N_21033,N_20833,N_20728);
nand U21034 (N_21034,N_20834,N_20890);
nor U21035 (N_21035,N_20957,N_20775);
nor U21036 (N_21036,N_20711,N_20903);
nor U21037 (N_21037,N_20995,N_20917);
or U21038 (N_21038,N_20894,N_20799);
or U21039 (N_21039,N_20937,N_20940);
nor U21040 (N_21040,N_20578,N_20703);
or U21041 (N_21041,N_20712,N_20755);
or U21042 (N_21042,N_20920,N_20986);
nand U21043 (N_21043,N_20541,N_20563);
nor U21044 (N_21044,N_20837,N_20701);
and U21045 (N_21045,N_20972,N_20929);
and U21046 (N_21046,N_20643,N_20529);
or U21047 (N_21047,N_20651,N_20576);
nor U21048 (N_21048,N_20987,N_20776);
xor U21049 (N_21049,N_20904,N_20706);
or U21050 (N_21050,N_20771,N_20635);
or U21051 (N_21051,N_20528,N_20687);
and U21052 (N_21052,N_20814,N_20561);
and U21053 (N_21053,N_20764,N_20708);
xor U21054 (N_21054,N_20657,N_20951);
nand U21055 (N_21055,N_20848,N_20956);
or U21056 (N_21056,N_20676,N_20689);
and U21057 (N_21057,N_20928,N_20885);
nor U21058 (N_21058,N_20854,N_20559);
nor U21059 (N_21059,N_20667,N_20808);
and U21060 (N_21060,N_20944,N_20621);
nor U21061 (N_21061,N_20996,N_20861);
nand U21062 (N_21062,N_20638,N_20582);
nand U21063 (N_21063,N_20868,N_20693);
xnor U21064 (N_21064,N_20777,N_20546);
or U21065 (N_21065,N_20838,N_20666);
nor U21066 (N_21066,N_20531,N_20514);
nor U21067 (N_21067,N_20884,N_20603);
and U21068 (N_21068,N_20547,N_20824);
nand U21069 (N_21069,N_20634,N_20516);
and U21070 (N_21070,N_20700,N_20908);
and U21071 (N_21071,N_20927,N_20760);
xnor U21072 (N_21072,N_20590,N_20719);
nor U21073 (N_21073,N_20620,N_20993);
nand U21074 (N_21074,N_20614,N_20870);
nor U21075 (N_21075,N_20572,N_20778);
or U21076 (N_21076,N_20998,N_20742);
or U21077 (N_21077,N_20513,N_20954);
xnor U21078 (N_21078,N_20595,N_20562);
and U21079 (N_21079,N_20896,N_20875);
nand U21080 (N_21080,N_20880,N_20653);
xor U21081 (N_21081,N_20677,N_20807);
and U21082 (N_21082,N_20919,N_20611);
nand U21083 (N_21083,N_20704,N_20823);
or U21084 (N_21084,N_20757,N_20619);
nand U21085 (N_21085,N_20675,N_20718);
and U21086 (N_21086,N_20580,N_20683);
or U21087 (N_21087,N_20625,N_20921);
or U21088 (N_21088,N_20945,N_20732);
xor U21089 (N_21089,N_20613,N_20512);
and U21090 (N_21090,N_20933,N_20825);
or U21091 (N_21091,N_20616,N_20905);
xor U21092 (N_21092,N_20685,N_20530);
nand U21093 (N_21093,N_20640,N_20926);
xnor U21094 (N_21094,N_20639,N_20978);
and U21095 (N_21095,N_20686,N_20680);
or U21096 (N_21096,N_20723,N_20953);
and U21097 (N_21097,N_20647,N_20963);
and U21098 (N_21098,N_20869,N_20507);
nand U21099 (N_21099,N_20806,N_20615);
or U21100 (N_21100,N_20669,N_20751);
xor U21101 (N_21101,N_20911,N_20540);
and U21102 (N_21102,N_20748,N_20923);
and U21103 (N_21103,N_20947,N_20598);
nand U21104 (N_21104,N_20988,N_20637);
or U21105 (N_21105,N_20664,N_20508);
nor U21106 (N_21106,N_20801,N_20705);
or U21107 (N_21107,N_20505,N_20959);
and U21108 (N_21108,N_20863,N_20946);
and U21109 (N_21109,N_20845,N_20759);
nand U21110 (N_21110,N_20909,N_20655);
or U21111 (N_21111,N_20767,N_20804);
nand U21112 (N_21112,N_20886,N_20501);
xnor U21113 (N_21113,N_20990,N_20517);
and U21114 (N_21114,N_20850,N_20912);
nor U21115 (N_21115,N_20740,N_20713);
xnor U21116 (N_21116,N_20671,N_20982);
xor U21117 (N_21117,N_20992,N_20548);
xor U21118 (N_21118,N_20899,N_20991);
nor U21119 (N_21119,N_20938,N_20882);
or U21120 (N_21120,N_20752,N_20697);
xor U21121 (N_21121,N_20750,N_20607);
and U21122 (N_21122,N_20661,N_20976);
and U21123 (N_21123,N_20526,N_20624);
nand U21124 (N_21124,N_20630,N_20983);
or U21125 (N_21125,N_20605,N_20522);
and U21126 (N_21126,N_20545,N_20534);
and U21127 (N_21127,N_20691,N_20761);
nor U21128 (N_21128,N_20811,N_20900);
xor U21129 (N_21129,N_20793,N_20556);
xnor U21130 (N_21130,N_20997,N_20549);
nor U21131 (N_21131,N_20857,N_20785);
or U21132 (N_21132,N_20769,N_20743);
or U21133 (N_21133,N_20726,N_20521);
and U21134 (N_21134,N_20597,N_20795);
nand U21135 (N_21135,N_20720,N_20753);
nand U21136 (N_21136,N_20569,N_20980);
or U21137 (N_21137,N_20949,N_20977);
nor U21138 (N_21138,N_20999,N_20577);
and U21139 (N_21139,N_20860,N_20631);
xor U21140 (N_21140,N_20536,N_20813);
or U21141 (N_21141,N_20695,N_20874);
or U21142 (N_21142,N_20891,N_20766);
nand U21143 (N_21143,N_20815,N_20519);
xor U21144 (N_21144,N_20672,N_20892);
xnor U21145 (N_21145,N_20557,N_20942);
or U21146 (N_21146,N_20818,N_20962);
or U21147 (N_21147,N_20571,N_20765);
nor U21148 (N_21148,N_20739,N_20558);
nor U21149 (N_21149,N_20994,N_20692);
or U21150 (N_21150,N_20564,N_20888);
or U21151 (N_21151,N_20809,N_20800);
and U21152 (N_21152,N_20762,N_20594);
xnor U21153 (N_21153,N_20663,N_20968);
xor U21154 (N_21154,N_20862,N_20805);
xor U21155 (N_21155,N_20871,N_20918);
and U21156 (N_21156,N_20539,N_20523);
xnor U21157 (N_21157,N_20915,N_20955);
nand U21158 (N_21158,N_20985,N_20596);
nor U21159 (N_21159,N_20674,N_20830);
and U21160 (N_21160,N_20756,N_20858);
or U21161 (N_21161,N_20935,N_20952);
or U21162 (N_21162,N_20585,N_20763);
nor U21163 (N_21163,N_20843,N_20503);
nor U21164 (N_21164,N_20747,N_20791);
nor U21165 (N_21165,N_20652,N_20787);
nand U21166 (N_21166,N_20537,N_20694);
and U21167 (N_21167,N_20533,N_20646);
nor U21168 (N_21168,N_20974,N_20836);
or U21169 (N_21169,N_20744,N_20566);
nand U21170 (N_21170,N_20914,N_20520);
and U21171 (N_21171,N_20738,N_20950);
nor U21172 (N_21172,N_20786,N_20964);
or U21173 (N_21173,N_20961,N_20729);
nand U21174 (N_21174,N_20618,N_20816);
xor U21175 (N_21175,N_20610,N_20532);
and U21176 (N_21176,N_20975,N_20710);
nor U21177 (N_21177,N_20510,N_20872);
or U21178 (N_21178,N_20901,N_20822);
and U21179 (N_21179,N_20754,N_20958);
or U21180 (N_21180,N_20879,N_20812);
and U21181 (N_21181,N_20831,N_20745);
nor U21182 (N_21182,N_20960,N_20628);
or U21183 (N_21183,N_20581,N_20859);
or U21184 (N_21184,N_20648,N_20781);
and U21185 (N_21185,N_20591,N_20741);
nor U21186 (N_21186,N_20788,N_20727);
nand U21187 (N_21187,N_20575,N_20864);
nor U21188 (N_21188,N_20500,N_20934);
or U21189 (N_21189,N_20524,N_20970);
and U21190 (N_21190,N_20730,N_20979);
nor U21191 (N_21191,N_20588,N_20971);
xor U21192 (N_21192,N_20609,N_20969);
xnor U21193 (N_21193,N_20907,N_20832);
and U21194 (N_21194,N_20924,N_20797);
nor U21195 (N_21195,N_20642,N_20783);
nor U21196 (N_21196,N_20731,N_20560);
nand U21197 (N_21197,N_20749,N_20583);
or U21198 (N_21198,N_20772,N_20893);
xor U21199 (N_21199,N_20654,N_20662);
or U21200 (N_21200,N_20589,N_20841);
or U21201 (N_21201,N_20784,N_20876);
nor U21202 (N_21202,N_20658,N_20768);
nand U21203 (N_21203,N_20881,N_20579);
xnor U21204 (N_21204,N_20897,N_20802);
or U21205 (N_21205,N_20587,N_20916);
xnor U21206 (N_21206,N_20828,N_20790);
nor U21207 (N_21207,N_20570,N_20649);
nor U21208 (N_21208,N_20629,N_20867);
xnor U21209 (N_21209,N_20641,N_20902);
xnor U21210 (N_21210,N_20573,N_20535);
nand U21211 (N_21211,N_20849,N_20509);
nor U21212 (N_21212,N_20699,N_20889);
or U21213 (N_21213,N_20567,N_20734);
and U21214 (N_21214,N_20684,N_20853);
xor U21215 (N_21215,N_20773,N_20873);
nor U21216 (N_21216,N_20839,N_20981);
and U21217 (N_21217,N_20665,N_20746);
or U21218 (N_21218,N_20553,N_20887);
and U21219 (N_21219,N_20819,N_20681);
xor U21220 (N_21220,N_20702,N_20803);
xnor U21221 (N_21221,N_20866,N_20829);
and U21222 (N_21222,N_20644,N_20810);
xnor U21223 (N_21223,N_20948,N_20895);
or U21224 (N_21224,N_20941,N_20724);
and U21225 (N_21225,N_20965,N_20623);
nor U21226 (N_21226,N_20842,N_20504);
and U21227 (N_21227,N_20852,N_20878);
nand U21228 (N_21228,N_20714,N_20758);
nor U21229 (N_21229,N_20709,N_20502);
nand U21230 (N_21230,N_20673,N_20827);
xnor U21231 (N_21231,N_20865,N_20682);
xnor U21232 (N_21232,N_20794,N_20735);
or U21233 (N_21233,N_20600,N_20931);
or U21234 (N_21234,N_20989,N_20550);
xor U21235 (N_21235,N_20716,N_20632);
xor U21236 (N_21236,N_20774,N_20670);
nand U21237 (N_21237,N_20538,N_20707);
or U21238 (N_21238,N_20840,N_20633);
nor U21239 (N_21239,N_20552,N_20565);
nor U21240 (N_21240,N_20715,N_20679);
xor U21241 (N_21241,N_20967,N_20913);
or U21242 (N_21242,N_20555,N_20835);
xor U21243 (N_21243,N_20645,N_20678);
nor U21244 (N_21244,N_20544,N_20660);
nand U21245 (N_21245,N_20656,N_20725);
nand U21246 (N_21246,N_20696,N_20659);
and U21247 (N_21247,N_20722,N_20973);
or U21248 (N_21248,N_20543,N_20568);
nand U21249 (N_21249,N_20737,N_20798);
or U21250 (N_21250,N_20622,N_20510);
and U21251 (N_21251,N_20546,N_20765);
nand U21252 (N_21252,N_20961,N_20863);
xnor U21253 (N_21253,N_20920,N_20828);
nand U21254 (N_21254,N_20842,N_20959);
nand U21255 (N_21255,N_20997,N_20668);
xor U21256 (N_21256,N_20996,N_20794);
nor U21257 (N_21257,N_20881,N_20646);
xor U21258 (N_21258,N_20606,N_20621);
xor U21259 (N_21259,N_20573,N_20660);
or U21260 (N_21260,N_20927,N_20585);
xnor U21261 (N_21261,N_20684,N_20646);
or U21262 (N_21262,N_20676,N_20714);
or U21263 (N_21263,N_20595,N_20884);
or U21264 (N_21264,N_20935,N_20806);
or U21265 (N_21265,N_20534,N_20502);
or U21266 (N_21266,N_20951,N_20886);
nor U21267 (N_21267,N_20769,N_20855);
xnor U21268 (N_21268,N_20770,N_20867);
xnor U21269 (N_21269,N_20515,N_20827);
or U21270 (N_21270,N_20922,N_20615);
nand U21271 (N_21271,N_20503,N_20812);
nor U21272 (N_21272,N_20577,N_20735);
xor U21273 (N_21273,N_20698,N_20895);
nor U21274 (N_21274,N_20825,N_20618);
nand U21275 (N_21275,N_20544,N_20884);
xnor U21276 (N_21276,N_20714,N_20569);
and U21277 (N_21277,N_20766,N_20972);
nor U21278 (N_21278,N_20733,N_20677);
or U21279 (N_21279,N_20535,N_20656);
nor U21280 (N_21280,N_20880,N_20941);
and U21281 (N_21281,N_20644,N_20931);
nand U21282 (N_21282,N_20868,N_20613);
and U21283 (N_21283,N_20770,N_20824);
nor U21284 (N_21284,N_20656,N_20501);
or U21285 (N_21285,N_20525,N_20626);
or U21286 (N_21286,N_20967,N_20514);
nand U21287 (N_21287,N_20602,N_20719);
or U21288 (N_21288,N_20680,N_20740);
nand U21289 (N_21289,N_20996,N_20748);
nand U21290 (N_21290,N_20701,N_20660);
xor U21291 (N_21291,N_20949,N_20781);
and U21292 (N_21292,N_20869,N_20992);
xor U21293 (N_21293,N_20645,N_20520);
nand U21294 (N_21294,N_20868,N_20561);
or U21295 (N_21295,N_20734,N_20892);
or U21296 (N_21296,N_20759,N_20651);
or U21297 (N_21297,N_20575,N_20613);
nor U21298 (N_21298,N_20782,N_20606);
nand U21299 (N_21299,N_20842,N_20506);
nor U21300 (N_21300,N_20696,N_20683);
or U21301 (N_21301,N_20878,N_20868);
or U21302 (N_21302,N_20643,N_20580);
xnor U21303 (N_21303,N_20765,N_20619);
nand U21304 (N_21304,N_20938,N_20507);
xnor U21305 (N_21305,N_20696,N_20599);
nand U21306 (N_21306,N_20655,N_20543);
nand U21307 (N_21307,N_20974,N_20936);
and U21308 (N_21308,N_20893,N_20506);
and U21309 (N_21309,N_20671,N_20545);
nor U21310 (N_21310,N_20902,N_20642);
and U21311 (N_21311,N_20592,N_20581);
xor U21312 (N_21312,N_20895,N_20522);
nand U21313 (N_21313,N_20833,N_20658);
or U21314 (N_21314,N_20515,N_20957);
nand U21315 (N_21315,N_20793,N_20694);
or U21316 (N_21316,N_20710,N_20781);
xnor U21317 (N_21317,N_20519,N_20669);
and U21318 (N_21318,N_20963,N_20855);
nor U21319 (N_21319,N_20766,N_20544);
and U21320 (N_21320,N_20539,N_20607);
nand U21321 (N_21321,N_20741,N_20979);
or U21322 (N_21322,N_20521,N_20639);
and U21323 (N_21323,N_20831,N_20716);
and U21324 (N_21324,N_20730,N_20958);
nand U21325 (N_21325,N_20860,N_20588);
and U21326 (N_21326,N_20588,N_20528);
or U21327 (N_21327,N_20723,N_20707);
xor U21328 (N_21328,N_20653,N_20754);
nand U21329 (N_21329,N_20660,N_20561);
nand U21330 (N_21330,N_20844,N_20856);
xor U21331 (N_21331,N_20617,N_20544);
or U21332 (N_21332,N_20537,N_20572);
nor U21333 (N_21333,N_20791,N_20501);
or U21334 (N_21334,N_20651,N_20577);
or U21335 (N_21335,N_20850,N_20647);
xor U21336 (N_21336,N_20641,N_20563);
nor U21337 (N_21337,N_20700,N_20861);
or U21338 (N_21338,N_20821,N_20906);
and U21339 (N_21339,N_20793,N_20698);
nor U21340 (N_21340,N_20756,N_20986);
nor U21341 (N_21341,N_20638,N_20916);
nand U21342 (N_21342,N_20733,N_20939);
and U21343 (N_21343,N_20898,N_20527);
nor U21344 (N_21344,N_20682,N_20876);
nor U21345 (N_21345,N_20767,N_20686);
nor U21346 (N_21346,N_20642,N_20671);
and U21347 (N_21347,N_20638,N_20644);
nand U21348 (N_21348,N_20872,N_20894);
or U21349 (N_21349,N_20772,N_20938);
xnor U21350 (N_21350,N_20824,N_20725);
and U21351 (N_21351,N_20815,N_20652);
and U21352 (N_21352,N_20775,N_20997);
nand U21353 (N_21353,N_20711,N_20768);
nor U21354 (N_21354,N_20924,N_20917);
xnor U21355 (N_21355,N_20800,N_20938);
and U21356 (N_21356,N_20715,N_20978);
nor U21357 (N_21357,N_20592,N_20985);
nor U21358 (N_21358,N_20915,N_20506);
nand U21359 (N_21359,N_20621,N_20520);
and U21360 (N_21360,N_20648,N_20528);
or U21361 (N_21361,N_20712,N_20691);
xnor U21362 (N_21362,N_20568,N_20813);
or U21363 (N_21363,N_20907,N_20713);
or U21364 (N_21364,N_20792,N_20778);
or U21365 (N_21365,N_20808,N_20976);
xnor U21366 (N_21366,N_20527,N_20822);
nand U21367 (N_21367,N_20646,N_20804);
and U21368 (N_21368,N_20910,N_20995);
nor U21369 (N_21369,N_20689,N_20579);
nor U21370 (N_21370,N_20607,N_20746);
or U21371 (N_21371,N_20670,N_20726);
nand U21372 (N_21372,N_20896,N_20915);
xor U21373 (N_21373,N_20584,N_20852);
xor U21374 (N_21374,N_20559,N_20857);
nor U21375 (N_21375,N_20800,N_20878);
and U21376 (N_21376,N_20591,N_20514);
nor U21377 (N_21377,N_20835,N_20962);
nor U21378 (N_21378,N_20850,N_20867);
xnor U21379 (N_21379,N_20687,N_20770);
or U21380 (N_21380,N_20898,N_20712);
nand U21381 (N_21381,N_20877,N_20642);
nor U21382 (N_21382,N_20897,N_20654);
xnor U21383 (N_21383,N_20873,N_20507);
or U21384 (N_21384,N_20760,N_20881);
nand U21385 (N_21385,N_20571,N_20800);
or U21386 (N_21386,N_20580,N_20682);
xor U21387 (N_21387,N_20575,N_20787);
nor U21388 (N_21388,N_20669,N_20573);
xor U21389 (N_21389,N_20924,N_20910);
or U21390 (N_21390,N_20969,N_20948);
or U21391 (N_21391,N_20626,N_20934);
xor U21392 (N_21392,N_20618,N_20978);
nand U21393 (N_21393,N_20842,N_20613);
nor U21394 (N_21394,N_20504,N_20542);
xor U21395 (N_21395,N_20689,N_20517);
and U21396 (N_21396,N_20965,N_20986);
nor U21397 (N_21397,N_20584,N_20868);
xnor U21398 (N_21398,N_20929,N_20549);
xnor U21399 (N_21399,N_20709,N_20686);
nor U21400 (N_21400,N_20801,N_20566);
nand U21401 (N_21401,N_20823,N_20972);
nand U21402 (N_21402,N_20503,N_20697);
nor U21403 (N_21403,N_20613,N_20947);
or U21404 (N_21404,N_20653,N_20637);
and U21405 (N_21405,N_20952,N_20555);
nand U21406 (N_21406,N_20708,N_20746);
and U21407 (N_21407,N_20681,N_20737);
xnor U21408 (N_21408,N_20795,N_20714);
xor U21409 (N_21409,N_20597,N_20916);
nand U21410 (N_21410,N_20778,N_20748);
nand U21411 (N_21411,N_20761,N_20890);
or U21412 (N_21412,N_20819,N_20582);
and U21413 (N_21413,N_20629,N_20790);
nand U21414 (N_21414,N_20571,N_20972);
nor U21415 (N_21415,N_20858,N_20586);
nor U21416 (N_21416,N_20529,N_20582);
xor U21417 (N_21417,N_20827,N_20529);
xor U21418 (N_21418,N_20575,N_20942);
or U21419 (N_21419,N_20700,N_20599);
and U21420 (N_21420,N_20994,N_20714);
nand U21421 (N_21421,N_20911,N_20715);
xor U21422 (N_21422,N_20730,N_20953);
and U21423 (N_21423,N_20873,N_20595);
xnor U21424 (N_21424,N_20561,N_20939);
xnor U21425 (N_21425,N_20903,N_20581);
xor U21426 (N_21426,N_20658,N_20749);
and U21427 (N_21427,N_20962,N_20593);
or U21428 (N_21428,N_20917,N_20886);
xnor U21429 (N_21429,N_20761,N_20645);
xor U21430 (N_21430,N_20988,N_20788);
nand U21431 (N_21431,N_20925,N_20970);
nand U21432 (N_21432,N_20802,N_20615);
nor U21433 (N_21433,N_20930,N_20924);
and U21434 (N_21434,N_20593,N_20918);
xor U21435 (N_21435,N_20811,N_20535);
or U21436 (N_21436,N_20665,N_20731);
and U21437 (N_21437,N_20725,N_20870);
nor U21438 (N_21438,N_20871,N_20956);
nand U21439 (N_21439,N_20566,N_20629);
nand U21440 (N_21440,N_20769,N_20781);
and U21441 (N_21441,N_20904,N_20555);
or U21442 (N_21442,N_20906,N_20564);
and U21443 (N_21443,N_20864,N_20957);
xnor U21444 (N_21444,N_20622,N_20832);
or U21445 (N_21445,N_20629,N_20868);
nor U21446 (N_21446,N_20798,N_20712);
or U21447 (N_21447,N_20695,N_20899);
and U21448 (N_21448,N_20766,N_20765);
nand U21449 (N_21449,N_20514,N_20612);
nor U21450 (N_21450,N_20994,N_20651);
xnor U21451 (N_21451,N_20789,N_20998);
xor U21452 (N_21452,N_20682,N_20793);
or U21453 (N_21453,N_20698,N_20908);
nand U21454 (N_21454,N_20653,N_20694);
nor U21455 (N_21455,N_20522,N_20693);
xnor U21456 (N_21456,N_20734,N_20659);
nor U21457 (N_21457,N_20973,N_20859);
nor U21458 (N_21458,N_20670,N_20662);
xnor U21459 (N_21459,N_20647,N_20678);
nand U21460 (N_21460,N_20815,N_20630);
and U21461 (N_21461,N_20976,N_20951);
xnor U21462 (N_21462,N_20847,N_20819);
and U21463 (N_21463,N_20807,N_20922);
or U21464 (N_21464,N_20970,N_20562);
and U21465 (N_21465,N_20643,N_20680);
xnor U21466 (N_21466,N_20740,N_20681);
xnor U21467 (N_21467,N_20812,N_20642);
and U21468 (N_21468,N_20901,N_20989);
nand U21469 (N_21469,N_20537,N_20736);
nor U21470 (N_21470,N_20505,N_20934);
xor U21471 (N_21471,N_20773,N_20601);
or U21472 (N_21472,N_20932,N_20983);
nand U21473 (N_21473,N_20981,N_20567);
or U21474 (N_21474,N_20685,N_20907);
and U21475 (N_21475,N_20971,N_20998);
and U21476 (N_21476,N_20584,N_20782);
or U21477 (N_21477,N_20684,N_20791);
nand U21478 (N_21478,N_20533,N_20691);
or U21479 (N_21479,N_20598,N_20874);
xnor U21480 (N_21480,N_20813,N_20848);
and U21481 (N_21481,N_20721,N_20575);
nor U21482 (N_21482,N_20666,N_20948);
nor U21483 (N_21483,N_20900,N_20647);
nor U21484 (N_21484,N_20915,N_20838);
nand U21485 (N_21485,N_20617,N_20962);
or U21486 (N_21486,N_20567,N_20768);
nand U21487 (N_21487,N_20739,N_20515);
and U21488 (N_21488,N_20620,N_20916);
xnor U21489 (N_21489,N_20803,N_20799);
or U21490 (N_21490,N_20838,N_20879);
xnor U21491 (N_21491,N_20694,N_20762);
or U21492 (N_21492,N_20806,N_20519);
nand U21493 (N_21493,N_20633,N_20598);
and U21494 (N_21494,N_20789,N_20646);
nor U21495 (N_21495,N_20696,N_20684);
nor U21496 (N_21496,N_20605,N_20819);
nor U21497 (N_21497,N_20592,N_20631);
or U21498 (N_21498,N_20735,N_20629);
nand U21499 (N_21499,N_20985,N_20861);
nand U21500 (N_21500,N_21083,N_21424);
xnor U21501 (N_21501,N_21345,N_21162);
or U21502 (N_21502,N_21129,N_21431);
xnor U21503 (N_21503,N_21216,N_21050);
nor U21504 (N_21504,N_21228,N_21114);
xnor U21505 (N_21505,N_21446,N_21080);
and U21506 (N_21506,N_21309,N_21176);
xor U21507 (N_21507,N_21220,N_21331);
or U21508 (N_21508,N_21429,N_21163);
nand U21509 (N_21509,N_21039,N_21440);
nand U21510 (N_21510,N_21200,N_21274);
nand U21511 (N_21511,N_21231,N_21277);
and U21512 (N_21512,N_21323,N_21320);
and U21513 (N_21513,N_21386,N_21079);
xnor U21514 (N_21514,N_21142,N_21249);
nor U21515 (N_21515,N_21393,N_21020);
and U21516 (N_21516,N_21361,N_21019);
xor U21517 (N_21517,N_21290,N_21418);
and U21518 (N_21518,N_21430,N_21230);
and U21519 (N_21519,N_21270,N_21475);
and U21520 (N_21520,N_21049,N_21375);
nor U21521 (N_21521,N_21089,N_21296);
nor U21522 (N_21522,N_21466,N_21155);
or U21523 (N_21523,N_21093,N_21340);
nand U21524 (N_21524,N_21141,N_21445);
nor U21525 (N_21525,N_21333,N_21243);
nor U21526 (N_21526,N_21450,N_21472);
nor U21527 (N_21527,N_21364,N_21409);
xor U21528 (N_21528,N_21298,N_21017);
xnor U21529 (N_21529,N_21315,N_21332);
nor U21530 (N_21530,N_21421,N_21169);
nand U21531 (N_21531,N_21058,N_21159);
xnor U21532 (N_21532,N_21091,N_21282);
xor U21533 (N_21533,N_21023,N_21301);
nand U21534 (N_21534,N_21411,N_21343);
nor U21535 (N_21535,N_21314,N_21160);
or U21536 (N_21536,N_21405,N_21355);
nand U21537 (N_21537,N_21130,N_21491);
nand U21538 (N_21538,N_21383,N_21040);
xnor U21539 (N_21539,N_21000,N_21497);
nor U21540 (N_21540,N_21055,N_21347);
nor U21541 (N_21541,N_21027,N_21225);
xnor U21542 (N_21542,N_21257,N_21478);
nor U21543 (N_21543,N_21457,N_21154);
xor U21544 (N_21544,N_21006,N_21490);
or U21545 (N_21545,N_21232,N_21145);
xor U21546 (N_21546,N_21030,N_21338);
nor U21547 (N_21547,N_21380,N_21035);
or U21548 (N_21548,N_21062,N_21453);
and U21549 (N_21549,N_21013,N_21413);
nor U21550 (N_21550,N_21212,N_21100);
nor U21551 (N_21551,N_21010,N_21188);
nor U21552 (N_21552,N_21346,N_21066);
nor U21553 (N_21553,N_21102,N_21121);
or U21554 (N_21554,N_21423,N_21117);
and U21555 (N_21555,N_21451,N_21455);
nor U21556 (N_21556,N_21064,N_21172);
or U21557 (N_21557,N_21038,N_21353);
nand U21558 (N_21558,N_21488,N_21495);
nand U21559 (N_21559,N_21279,N_21113);
xor U21560 (N_21560,N_21029,N_21311);
nor U21561 (N_21561,N_21492,N_21218);
nor U21562 (N_21562,N_21138,N_21428);
xnor U21563 (N_21563,N_21021,N_21085);
nor U21564 (N_21564,N_21187,N_21362);
xnor U21565 (N_21565,N_21056,N_21244);
xor U21566 (N_21566,N_21042,N_21069);
or U21567 (N_21567,N_21389,N_21151);
xor U21568 (N_21568,N_21369,N_21449);
and U21569 (N_21569,N_21496,N_21097);
and U21570 (N_21570,N_21047,N_21268);
xor U21571 (N_21571,N_21482,N_21476);
and U21572 (N_21572,N_21272,N_21190);
or U21573 (N_21573,N_21334,N_21258);
or U21574 (N_21574,N_21084,N_21378);
nand U21575 (N_21575,N_21112,N_21381);
nor U21576 (N_21576,N_21276,N_21173);
nand U21577 (N_21577,N_21061,N_21132);
nand U21578 (N_21578,N_21376,N_21137);
nand U21579 (N_21579,N_21307,N_21266);
or U21580 (N_21580,N_21417,N_21330);
xor U21581 (N_21581,N_21358,N_21278);
nand U21582 (N_21582,N_21480,N_21167);
and U21583 (N_21583,N_21305,N_21441);
or U21584 (N_21584,N_21054,N_21177);
or U21585 (N_21585,N_21240,N_21374);
xor U21586 (N_21586,N_21014,N_21170);
nor U21587 (N_21587,N_21094,N_21452);
and U21588 (N_21588,N_21204,N_21394);
or U21589 (N_21589,N_21146,N_21260);
xnor U21590 (N_21590,N_21245,N_21438);
nor U21591 (N_21591,N_21032,N_21107);
nor U21592 (N_21592,N_21165,N_21227);
or U21593 (N_21593,N_21373,N_21456);
xnor U21594 (N_21594,N_21289,N_21148);
xor U21595 (N_21595,N_21426,N_21072);
and U21596 (N_21596,N_21484,N_21003);
nor U21597 (N_21597,N_21057,N_21180);
or U21598 (N_21598,N_21067,N_21237);
xnor U21599 (N_21599,N_21007,N_21202);
and U21600 (N_21600,N_21341,N_21203);
and U21601 (N_21601,N_21081,N_21463);
nor U21602 (N_21602,N_21224,N_21250);
or U21603 (N_21603,N_21462,N_21001);
nor U21604 (N_21604,N_21025,N_21256);
or U21605 (N_21605,N_21174,N_21168);
or U21606 (N_21606,N_21179,N_21269);
xor U21607 (N_21607,N_21372,N_21087);
nor U21608 (N_21608,N_21422,N_21494);
xor U21609 (N_21609,N_21267,N_21403);
or U21610 (N_21610,N_21086,N_21280);
nor U21611 (N_21611,N_21195,N_21499);
nor U21612 (N_21612,N_21184,N_21226);
and U21613 (N_21613,N_21291,N_21099);
and U21614 (N_21614,N_21234,N_21248);
or U21615 (N_21615,N_21458,N_21120);
or U21616 (N_21616,N_21005,N_21400);
nor U21617 (N_21617,N_21390,N_21461);
or U21618 (N_21618,N_21308,N_21398);
xor U21619 (N_21619,N_21473,N_21359);
nand U21620 (N_21620,N_21391,N_21209);
and U21621 (N_21621,N_21396,N_21063);
and U21622 (N_21622,N_21486,N_21365);
nor U21623 (N_21623,N_21263,N_21485);
and U21624 (N_21624,N_21073,N_21175);
xor U21625 (N_21625,N_21354,N_21349);
and U21626 (N_21626,N_21071,N_21414);
and U21627 (N_21627,N_21026,N_21329);
or U21628 (N_21628,N_21316,N_21217);
xor U21629 (N_21629,N_21284,N_21402);
nand U21630 (N_21630,N_21467,N_21447);
xnor U21631 (N_21631,N_21356,N_21205);
and U21632 (N_21632,N_21233,N_21382);
and U21633 (N_21633,N_21285,N_21420);
and U21634 (N_21634,N_21498,N_21344);
and U21635 (N_21635,N_21186,N_21041);
nand U21636 (N_21636,N_21252,N_21281);
xnor U21637 (N_21637,N_21408,N_21493);
nand U21638 (N_21638,N_21191,N_21322);
nor U21639 (N_21639,N_21024,N_21147);
nor U21640 (N_21640,N_21127,N_21051);
nor U21641 (N_21641,N_21299,N_21109);
nor U21642 (N_21642,N_21339,N_21335);
xor U21643 (N_21643,N_21407,N_21479);
nand U21644 (N_21644,N_21034,N_21406);
or U21645 (N_21645,N_21255,N_21131);
xnor U21646 (N_21646,N_21008,N_21351);
nor U21647 (N_21647,N_21262,N_21192);
and U21648 (N_21648,N_21294,N_21292);
or U21649 (N_21649,N_21325,N_21443);
and U21650 (N_21650,N_21033,N_21101);
or U21651 (N_21651,N_21370,N_21367);
nand U21652 (N_21652,N_21213,N_21004);
or U21653 (N_21653,N_21348,N_21223);
xnor U21654 (N_21654,N_21385,N_21412);
and U21655 (N_21655,N_21327,N_21208);
nand U21656 (N_21656,N_21321,N_21253);
and U21657 (N_21657,N_21247,N_21219);
or U21658 (N_21658,N_21324,N_21283);
nand U21659 (N_21659,N_21106,N_21222);
or U21660 (N_21660,N_21483,N_21286);
or U21661 (N_21661,N_21002,N_21074);
or U21662 (N_21662,N_21388,N_21293);
xnor U21663 (N_21663,N_21241,N_21031);
nor U21664 (N_21664,N_21448,N_21210);
or U21665 (N_21665,N_21288,N_21312);
xnor U21666 (N_21666,N_21110,N_21350);
nand U21667 (N_21667,N_21152,N_21236);
and U21668 (N_21668,N_21206,N_21300);
nand U21669 (N_21669,N_21119,N_21487);
nand U21670 (N_21670,N_21427,N_21239);
or U21671 (N_21671,N_21149,N_21157);
or U21672 (N_21672,N_21379,N_21442);
nor U21673 (N_21673,N_21181,N_21489);
or U21674 (N_21674,N_21095,N_21016);
nor U21675 (N_21675,N_21158,N_21028);
xor U21676 (N_21676,N_21434,N_21171);
and U21677 (N_21677,N_21363,N_21082);
and U21678 (N_21678,N_21077,N_21092);
or U21679 (N_21679,N_21317,N_21022);
or U21680 (N_21680,N_21377,N_21433);
or U21681 (N_21681,N_21437,N_21122);
nor U21682 (N_21682,N_21435,N_21215);
or U21683 (N_21683,N_21143,N_21133);
and U21684 (N_21684,N_21139,N_21328);
or U21685 (N_21685,N_21297,N_21135);
xor U21686 (N_21686,N_21153,N_21326);
nor U21687 (N_21687,N_21271,N_21235);
and U21688 (N_21688,N_21183,N_21425);
xnor U21689 (N_21689,N_21126,N_21404);
nand U21690 (N_21690,N_21392,N_21018);
or U21691 (N_21691,N_21465,N_21295);
nor U21692 (N_21692,N_21287,N_21009);
nor U21693 (N_21693,N_21125,N_21161);
and U21694 (N_21694,N_21460,N_21468);
nand U21695 (N_21695,N_21470,N_21189);
xor U21696 (N_21696,N_21124,N_21166);
nand U21697 (N_21697,N_21459,N_21144);
xnor U21698 (N_21698,N_21196,N_21432);
nor U21699 (N_21699,N_21318,N_21128);
and U21700 (N_21700,N_21104,N_21384);
nand U21701 (N_21701,N_21469,N_21078);
xnor U21702 (N_21702,N_21261,N_21156);
and U21703 (N_21703,N_21088,N_21242);
or U21704 (N_21704,N_21352,N_21045);
xor U21705 (N_21705,N_21123,N_21419);
and U21706 (N_21706,N_21342,N_21471);
xor U21707 (N_21707,N_21319,N_21015);
nand U21708 (N_21708,N_21108,N_21090);
nand U21709 (N_21709,N_21313,N_21068);
nor U21710 (N_21710,N_21150,N_21366);
xnor U21711 (N_21711,N_21052,N_21194);
xor U21712 (N_21712,N_21229,N_21360);
xnor U21713 (N_21713,N_21306,N_21444);
xor U21714 (N_21714,N_21115,N_21439);
nand U21715 (N_21715,N_21048,N_21037);
or U21716 (N_21716,N_21436,N_21197);
nand U21717 (N_21717,N_21046,N_21454);
or U21718 (N_21718,N_21302,N_21207);
nand U21719 (N_21719,N_21201,N_21103);
xnor U21720 (N_21720,N_21111,N_21273);
nor U21721 (N_21721,N_21185,N_21410);
xor U21722 (N_21722,N_21199,N_21304);
nor U21723 (N_21723,N_21477,N_21105);
and U21724 (N_21724,N_21310,N_21251);
xnor U21725 (N_21725,N_21134,N_21474);
and U21726 (N_21726,N_21065,N_21011);
xor U21727 (N_21727,N_21481,N_21044);
nand U21728 (N_21728,N_21043,N_21399);
xnor U21729 (N_21729,N_21140,N_21098);
or U21730 (N_21730,N_21012,N_21337);
nand U21731 (N_21731,N_21060,N_21182);
nand U21732 (N_21732,N_21395,N_21357);
nand U21733 (N_21733,N_21464,N_21336);
nor U21734 (N_21734,N_21368,N_21036);
nand U21735 (N_21735,N_21164,N_21116);
or U21736 (N_21736,N_21371,N_21076);
nand U21737 (N_21737,N_21118,N_21238);
or U21738 (N_21738,N_21259,N_21070);
nor U21739 (N_21739,N_21265,N_21193);
xor U21740 (N_21740,N_21096,N_21059);
nor U21741 (N_21741,N_21246,N_21415);
and U21742 (N_21742,N_21198,N_21075);
nand U21743 (N_21743,N_21387,N_21397);
or U21744 (N_21744,N_21178,N_21053);
xnor U21745 (N_21745,N_21416,N_21275);
or U21746 (N_21746,N_21214,N_21401);
nand U21747 (N_21747,N_21254,N_21264);
nor U21748 (N_21748,N_21221,N_21136);
xnor U21749 (N_21749,N_21303,N_21211);
and U21750 (N_21750,N_21141,N_21180);
or U21751 (N_21751,N_21266,N_21462);
or U21752 (N_21752,N_21059,N_21293);
nand U21753 (N_21753,N_21210,N_21457);
nor U21754 (N_21754,N_21210,N_21150);
or U21755 (N_21755,N_21204,N_21459);
nand U21756 (N_21756,N_21138,N_21290);
nor U21757 (N_21757,N_21159,N_21084);
and U21758 (N_21758,N_21329,N_21159);
xnor U21759 (N_21759,N_21235,N_21286);
nand U21760 (N_21760,N_21458,N_21241);
nand U21761 (N_21761,N_21316,N_21444);
nand U21762 (N_21762,N_21150,N_21083);
nand U21763 (N_21763,N_21300,N_21489);
nor U21764 (N_21764,N_21451,N_21471);
and U21765 (N_21765,N_21020,N_21060);
and U21766 (N_21766,N_21307,N_21458);
nand U21767 (N_21767,N_21254,N_21198);
xor U21768 (N_21768,N_21094,N_21459);
nand U21769 (N_21769,N_21322,N_21472);
or U21770 (N_21770,N_21225,N_21276);
nor U21771 (N_21771,N_21267,N_21279);
xor U21772 (N_21772,N_21104,N_21291);
nor U21773 (N_21773,N_21267,N_21413);
xnor U21774 (N_21774,N_21418,N_21111);
and U21775 (N_21775,N_21295,N_21093);
nor U21776 (N_21776,N_21043,N_21333);
nand U21777 (N_21777,N_21257,N_21434);
and U21778 (N_21778,N_21246,N_21000);
xor U21779 (N_21779,N_21432,N_21352);
or U21780 (N_21780,N_21393,N_21465);
or U21781 (N_21781,N_21268,N_21393);
or U21782 (N_21782,N_21238,N_21489);
xnor U21783 (N_21783,N_21023,N_21411);
or U21784 (N_21784,N_21464,N_21071);
or U21785 (N_21785,N_21357,N_21291);
nand U21786 (N_21786,N_21351,N_21126);
nand U21787 (N_21787,N_21251,N_21169);
and U21788 (N_21788,N_21001,N_21067);
nand U21789 (N_21789,N_21310,N_21093);
xnor U21790 (N_21790,N_21379,N_21006);
or U21791 (N_21791,N_21456,N_21341);
xor U21792 (N_21792,N_21294,N_21058);
nand U21793 (N_21793,N_21259,N_21209);
or U21794 (N_21794,N_21145,N_21064);
and U21795 (N_21795,N_21024,N_21210);
xor U21796 (N_21796,N_21013,N_21287);
or U21797 (N_21797,N_21303,N_21044);
nand U21798 (N_21798,N_21203,N_21058);
or U21799 (N_21799,N_21232,N_21354);
nand U21800 (N_21800,N_21486,N_21436);
nor U21801 (N_21801,N_21258,N_21239);
and U21802 (N_21802,N_21168,N_21092);
xor U21803 (N_21803,N_21042,N_21239);
xor U21804 (N_21804,N_21468,N_21215);
nor U21805 (N_21805,N_21123,N_21465);
xor U21806 (N_21806,N_21292,N_21329);
xor U21807 (N_21807,N_21460,N_21231);
or U21808 (N_21808,N_21390,N_21200);
nor U21809 (N_21809,N_21435,N_21259);
nand U21810 (N_21810,N_21024,N_21183);
nor U21811 (N_21811,N_21217,N_21196);
xnor U21812 (N_21812,N_21395,N_21086);
or U21813 (N_21813,N_21254,N_21210);
and U21814 (N_21814,N_21323,N_21450);
or U21815 (N_21815,N_21028,N_21489);
nand U21816 (N_21816,N_21246,N_21332);
and U21817 (N_21817,N_21003,N_21412);
nor U21818 (N_21818,N_21476,N_21398);
xor U21819 (N_21819,N_21202,N_21392);
nor U21820 (N_21820,N_21359,N_21385);
nor U21821 (N_21821,N_21185,N_21064);
or U21822 (N_21822,N_21226,N_21096);
nand U21823 (N_21823,N_21344,N_21365);
xnor U21824 (N_21824,N_21499,N_21328);
or U21825 (N_21825,N_21219,N_21384);
nand U21826 (N_21826,N_21119,N_21442);
and U21827 (N_21827,N_21437,N_21024);
xor U21828 (N_21828,N_21139,N_21164);
and U21829 (N_21829,N_21202,N_21153);
or U21830 (N_21830,N_21045,N_21196);
xor U21831 (N_21831,N_21148,N_21161);
nand U21832 (N_21832,N_21323,N_21298);
xor U21833 (N_21833,N_21457,N_21016);
and U21834 (N_21834,N_21076,N_21441);
and U21835 (N_21835,N_21371,N_21083);
xor U21836 (N_21836,N_21421,N_21106);
nor U21837 (N_21837,N_21430,N_21177);
nand U21838 (N_21838,N_21481,N_21364);
and U21839 (N_21839,N_21111,N_21256);
nor U21840 (N_21840,N_21189,N_21108);
nor U21841 (N_21841,N_21190,N_21256);
and U21842 (N_21842,N_21279,N_21080);
xor U21843 (N_21843,N_21480,N_21379);
xnor U21844 (N_21844,N_21395,N_21215);
xor U21845 (N_21845,N_21404,N_21313);
or U21846 (N_21846,N_21038,N_21098);
nor U21847 (N_21847,N_21491,N_21364);
and U21848 (N_21848,N_21350,N_21252);
or U21849 (N_21849,N_21074,N_21496);
xnor U21850 (N_21850,N_21337,N_21100);
nor U21851 (N_21851,N_21383,N_21278);
xor U21852 (N_21852,N_21309,N_21204);
nand U21853 (N_21853,N_21449,N_21492);
or U21854 (N_21854,N_21384,N_21312);
nor U21855 (N_21855,N_21226,N_21156);
xor U21856 (N_21856,N_21027,N_21043);
nand U21857 (N_21857,N_21063,N_21225);
xor U21858 (N_21858,N_21452,N_21030);
or U21859 (N_21859,N_21035,N_21473);
and U21860 (N_21860,N_21455,N_21005);
and U21861 (N_21861,N_21030,N_21349);
and U21862 (N_21862,N_21442,N_21005);
nand U21863 (N_21863,N_21451,N_21414);
and U21864 (N_21864,N_21290,N_21341);
or U21865 (N_21865,N_21321,N_21478);
or U21866 (N_21866,N_21174,N_21430);
and U21867 (N_21867,N_21109,N_21160);
nand U21868 (N_21868,N_21407,N_21423);
or U21869 (N_21869,N_21248,N_21358);
and U21870 (N_21870,N_21361,N_21350);
nand U21871 (N_21871,N_21269,N_21050);
nand U21872 (N_21872,N_21358,N_21489);
nand U21873 (N_21873,N_21179,N_21280);
xnor U21874 (N_21874,N_21185,N_21260);
or U21875 (N_21875,N_21477,N_21082);
nand U21876 (N_21876,N_21421,N_21131);
nand U21877 (N_21877,N_21168,N_21150);
xnor U21878 (N_21878,N_21419,N_21066);
or U21879 (N_21879,N_21288,N_21403);
or U21880 (N_21880,N_21018,N_21440);
nand U21881 (N_21881,N_21455,N_21033);
and U21882 (N_21882,N_21271,N_21455);
or U21883 (N_21883,N_21185,N_21246);
and U21884 (N_21884,N_21352,N_21268);
and U21885 (N_21885,N_21088,N_21408);
nand U21886 (N_21886,N_21439,N_21468);
and U21887 (N_21887,N_21167,N_21023);
nand U21888 (N_21888,N_21097,N_21352);
nor U21889 (N_21889,N_21327,N_21283);
xor U21890 (N_21890,N_21383,N_21227);
and U21891 (N_21891,N_21304,N_21211);
or U21892 (N_21892,N_21278,N_21347);
or U21893 (N_21893,N_21483,N_21050);
xnor U21894 (N_21894,N_21485,N_21071);
nor U21895 (N_21895,N_21230,N_21492);
xnor U21896 (N_21896,N_21275,N_21394);
and U21897 (N_21897,N_21158,N_21010);
and U21898 (N_21898,N_21168,N_21052);
nand U21899 (N_21899,N_21025,N_21454);
or U21900 (N_21900,N_21349,N_21098);
and U21901 (N_21901,N_21373,N_21155);
or U21902 (N_21902,N_21208,N_21446);
and U21903 (N_21903,N_21136,N_21319);
and U21904 (N_21904,N_21454,N_21182);
or U21905 (N_21905,N_21093,N_21446);
nand U21906 (N_21906,N_21101,N_21062);
nor U21907 (N_21907,N_21425,N_21352);
nand U21908 (N_21908,N_21181,N_21151);
xnor U21909 (N_21909,N_21469,N_21081);
or U21910 (N_21910,N_21104,N_21110);
and U21911 (N_21911,N_21467,N_21480);
nand U21912 (N_21912,N_21220,N_21103);
and U21913 (N_21913,N_21110,N_21126);
xor U21914 (N_21914,N_21215,N_21441);
and U21915 (N_21915,N_21087,N_21097);
and U21916 (N_21916,N_21214,N_21315);
nand U21917 (N_21917,N_21180,N_21136);
nor U21918 (N_21918,N_21026,N_21172);
nor U21919 (N_21919,N_21209,N_21419);
nor U21920 (N_21920,N_21018,N_21133);
nor U21921 (N_21921,N_21437,N_21452);
nand U21922 (N_21922,N_21282,N_21229);
and U21923 (N_21923,N_21267,N_21263);
nor U21924 (N_21924,N_21174,N_21377);
or U21925 (N_21925,N_21413,N_21167);
or U21926 (N_21926,N_21078,N_21230);
nor U21927 (N_21927,N_21086,N_21027);
or U21928 (N_21928,N_21283,N_21064);
xnor U21929 (N_21929,N_21369,N_21013);
or U21930 (N_21930,N_21248,N_21325);
or U21931 (N_21931,N_21297,N_21250);
nor U21932 (N_21932,N_21137,N_21097);
and U21933 (N_21933,N_21218,N_21159);
and U21934 (N_21934,N_21474,N_21386);
or U21935 (N_21935,N_21343,N_21372);
and U21936 (N_21936,N_21179,N_21058);
nand U21937 (N_21937,N_21462,N_21093);
or U21938 (N_21938,N_21486,N_21080);
xnor U21939 (N_21939,N_21254,N_21341);
xnor U21940 (N_21940,N_21109,N_21178);
or U21941 (N_21941,N_21196,N_21242);
nand U21942 (N_21942,N_21200,N_21232);
nand U21943 (N_21943,N_21360,N_21137);
or U21944 (N_21944,N_21119,N_21294);
xnor U21945 (N_21945,N_21346,N_21474);
nand U21946 (N_21946,N_21123,N_21093);
xnor U21947 (N_21947,N_21320,N_21217);
nand U21948 (N_21948,N_21049,N_21405);
or U21949 (N_21949,N_21256,N_21091);
and U21950 (N_21950,N_21248,N_21408);
nor U21951 (N_21951,N_21347,N_21419);
nor U21952 (N_21952,N_21074,N_21420);
nor U21953 (N_21953,N_21312,N_21309);
or U21954 (N_21954,N_21436,N_21339);
or U21955 (N_21955,N_21108,N_21070);
xor U21956 (N_21956,N_21443,N_21315);
or U21957 (N_21957,N_21358,N_21454);
xnor U21958 (N_21958,N_21468,N_21076);
and U21959 (N_21959,N_21180,N_21039);
xor U21960 (N_21960,N_21431,N_21445);
and U21961 (N_21961,N_21105,N_21376);
and U21962 (N_21962,N_21160,N_21392);
xor U21963 (N_21963,N_21254,N_21246);
and U21964 (N_21964,N_21060,N_21380);
nor U21965 (N_21965,N_21055,N_21468);
and U21966 (N_21966,N_21038,N_21345);
and U21967 (N_21967,N_21374,N_21424);
xnor U21968 (N_21968,N_21351,N_21233);
nand U21969 (N_21969,N_21039,N_21447);
or U21970 (N_21970,N_21499,N_21494);
and U21971 (N_21971,N_21323,N_21170);
nor U21972 (N_21972,N_21253,N_21265);
or U21973 (N_21973,N_21469,N_21372);
nand U21974 (N_21974,N_21029,N_21261);
nand U21975 (N_21975,N_21049,N_21372);
nand U21976 (N_21976,N_21310,N_21151);
and U21977 (N_21977,N_21355,N_21163);
or U21978 (N_21978,N_21264,N_21388);
or U21979 (N_21979,N_21346,N_21216);
and U21980 (N_21980,N_21065,N_21103);
nand U21981 (N_21981,N_21110,N_21477);
or U21982 (N_21982,N_21267,N_21081);
or U21983 (N_21983,N_21462,N_21169);
or U21984 (N_21984,N_21276,N_21194);
nand U21985 (N_21985,N_21222,N_21033);
or U21986 (N_21986,N_21454,N_21042);
nand U21987 (N_21987,N_21393,N_21157);
xor U21988 (N_21988,N_21229,N_21154);
and U21989 (N_21989,N_21086,N_21196);
xor U21990 (N_21990,N_21371,N_21356);
and U21991 (N_21991,N_21440,N_21360);
nor U21992 (N_21992,N_21358,N_21009);
and U21993 (N_21993,N_21445,N_21137);
xor U21994 (N_21994,N_21494,N_21373);
nor U21995 (N_21995,N_21042,N_21484);
or U21996 (N_21996,N_21173,N_21121);
or U21997 (N_21997,N_21158,N_21267);
nand U21998 (N_21998,N_21434,N_21397);
nor U21999 (N_21999,N_21498,N_21191);
nor U22000 (N_22000,N_21997,N_21835);
nand U22001 (N_22001,N_21687,N_21829);
nor U22002 (N_22002,N_21524,N_21656);
nor U22003 (N_22003,N_21973,N_21659);
nor U22004 (N_22004,N_21534,N_21544);
nor U22005 (N_22005,N_21844,N_21560);
nor U22006 (N_22006,N_21916,N_21870);
nand U22007 (N_22007,N_21837,N_21709);
xnor U22008 (N_22008,N_21507,N_21741);
xnor U22009 (N_22009,N_21630,N_21721);
or U22010 (N_22010,N_21777,N_21954);
xnor U22011 (N_22011,N_21909,N_21712);
or U22012 (N_22012,N_21778,N_21776);
xnor U22013 (N_22013,N_21750,N_21617);
nor U22014 (N_22014,N_21807,N_21886);
and U22015 (N_22015,N_21917,N_21629);
nor U22016 (N_22016,N_21640,N_21736);
nor U22017 (N_22017,N_21615,N_21998);
and U22018 (N_22018,N_21670,N_21865);
xnor U22019 (N_22019,N_21848,N_21590);
or U22020 (N_22020,N_21546,N_21825);
and U22021 (N_22021,N_21627,N_21708);
nor U22022 (N_22022,N_21999,N_21566);
nor U22023 (N_22023,N_21834,N_21734);
or U22024 (N_22024,N_21793,N_21550);
nor U22025 (N_22025,N_21786,N_21822);
xnor U22026 (N_22026,N_21919,N_21592);
and U22027 (N_22027,N_21811,N_21842);
nand U22028 (N_22028,N_21542,N_21730);
or U22029 (N_22029,N_21691,N_21717);
and U22030 (N_22030,N_21828,N_21802);
xor U22031 (N_22031,N_21703,N_21685);
nor U22032 (N_22032,N_21962,N_21573);
xor U22033 (N_22033,N_21826,N_21924);
and U22034 (N_22034,N_21767,N_21985);
nand U22035 (N_22035,N_21603,N_21645);
or U22036 (N_22036,N_21654,N_21693);
nor U22037 (N_22037,N_21583,N_21795);
and U22038 (N_22038,N_21780,N_21894);
or U22039 (N_22039,N_21641,N_21902);
nor U22040 (N_22040,N_21788,N_21801);
or U22041 (N_22041,N_21791,N_21614);
or U22042 (N_22042,N_21591,N_21881);
or U22043 (N_22043,N_21984,N_21664);
and U22044 (N_22044,N_21686,N_21503);
and U22045 (N_22045,N_21612,N_21940);
nor U22046 (N_22046,N_21775,N_21876);
nor U22047 (N_22047,N_21809,N_21638);
xnor U22048 (N_22048,N_21574,N_21548);
xor U22049 (N_22049,N_21990,N_21994);
nand U22050 (N_22050,N_21789,N_21831);
nor U22051 (N_22051,N_21599,N_21637);
nor U22052 (N_22052,N_21509,N_21991);
and U22053 (N_22053,N_21996,N_21972);
nor U22054 (N_22054,N_21680,N_21711);
and U22055 (N_22055,N_21514,N_21500);
nand U22056 (N_22056,N_21506,N_21600);
or U22057 (N_22057,N_21959,N_21849);
nor U22058 (N_22058,N_21974,N_21915);
or U22059 (N_22059,N_21678,N_21636);
nand U22060 (N_22060,N_21947,N_21867);
nand U22061 (N_22061,N_21593,N_21563);
nor U22062 (N_22062,N_21633,N_21679);
nor U22063 (N_22063,N_21861,N_21960);
or U22064 (N_22064,N_21675,N_21946);
and U22065 (N_22065,N_21905,N_21850);
or U22066 (N_22066,N_21648,N_21758);
xor U22067 (N_22067,N_21812,N_21677);
nand U22068 (N_22068,N_21597,N_21732);
and U22069 (N_22069,N_21774,N_21816);
xnor U22070 (N_22070,N_21933,N_21644);
nor U22071 (N_22071,N_21950,N_21935);
nand U22072 (N_22072,N_21521,N_21983);
and U22073 (N_22073,N_21653,N_21926);
xor U22074 (N_22074,N_21803,N_21893);
nand U22075 (N_22075,N_21530,N_21879);
nand U22076 (N_22076,N_21971,N_21862);
nor U22077 (N_22077,N_21810,N_21863);
or U22078 (N_22078,N_21626,N_21604);
xor U22079 (N_22079,N_21925,N_21649);
and U22080 (N_22080,N_21657,N_21769);
xnor U22081 (N_22081,N_21525,N_21818);
xnor U22082 (N_22082,N_21745,N_21873);
xor U22083 (N_22083,N_21541,N_21569);
and U22084 (N_22084,N_21505,N_21901);
or U22085 (N_22085,N_21557,N_21661);
xor U22086 (N_22086,N_21864,N_21673);
nor U22087 (N_22087,N_21531,N_21535);
nand U22088 (N_22088,N_21790,N_21771);
xnor U22089 (N_22089,N_21662,N_21719);
nand U22090 (N_22090,N_21938,N_21552);
nand U22091 (N_22091,N_21911,N_21949);
xor U22092 (N_22092,N_21572,N_21526);
and U22093 (N_22093,N_21781,N_21533);
or U22094 (N_22094,N_21756,N_21692);
and U22095 (N_22095,N_21658,N_21581);
xor U22096 (N_22096,N_21773,N_21930);
nor U22097 (N_22097,N_21968,N_21596);
xnor U22098 (N_22098,N_21969,N_21737);
nor U22099 (N_22099,N_21868,N_21619);
and U22100 (N_22100,N_21532,N_21515);
and U22101 (N_22101,N_21878,N_21823);
xor U22102 (N_22102,N_21553,N_21609);
nor U22103 (N_22103,N_21527,N_21714);
nand U22104 (N_22104,N_21502,N_21900);
and U22105 (N_22105,N_21965,N_21508);
nand U22106 (N_22106,N_21547,N_21671);
or U22107 (N_22107,N_21877,N_21704);
or U22108 (N_22108,N_21551,N_21976);
and U22109 (N_22109,N_21602,N_21753);
xnor U22110 (N_22110,N_21883,N_21880);
xnor U22111 (N_22111,N_21945,N_21549);
nor U22112 (N_22112,N_21872,N_21833);
and U22113 (N_22113,N_21631,N_21565);
xnor U22114 (N_22114,N_21855,N_21815);
or U22115 (N_22115,N_21797,N_21707);
or U22116 (N_22116,N_21857,N_21808);
and U22117 (N_22117,N_21763,N_21896);
and U22118 (N_22118,N_21501,N_21794);
or U22119 (N_22119,N_21696,N_21610);
and U22120 (N_22120,N_21989,N_21706);
nor U22121 (N_22121,N_21922,N_21655);
xor U22122 (N_22122,N_21884,N_21622);
nand U22123 (N_22123,N_21580,N_21598);
nand U22124 (N_22124,N_21529,N_21699);
and U22125 (N_22125,N_21585,N_21584);
or U22126 (N_22126,N_21956,N_21571);
and U22127 (N_22127,N_21830,N_21683);
and U22128 (N_22128,N_21827,N_21513);
xnor U22129 (N_22129,N_21840,N_21952);
or U22130 (N_22130,N_21860,N_21986);
or U22131 (N_22131,N_21931,N_21504);
xnor U22132 (N_22132,N_21701,N_21616);
xor U22133 (N_22133,N_21582,N_21889);
nand U22134 (N_22134,N_21943,N_21824);
nand U22135 (N_22135,N_21854,N_21921);
nor U22136 (N_22136,N_21611,N_21620);
and U22137 (N_22137,N_21770,N_21682);
and U22138 (N_22138,N_21601,N_21684);
nor U22139 (N_22139,N_21647,N_21747);
and U22140 (N_22140,N_21606,N_21937);
nor U22141 (N_22141,N_21910,N_21804);
xnor U22142 (N_22142,N_21715,N_21512);
xor U22143 (N_22143,N_21888,N_21895);
or U22144 (N_22144,N_21594,N_21744);
or U22145 (N_22145,N_21847,N_21559);
nand U22146 (N_22146,N_21705,N_21543);
nand U22147 (N_22147,N_21843,N_21676);
xor U22148 (N_22148,N_21729,N_21672);
nor U22149 (N_22149,N_21817,N_21595);
xor U22150 (N_22150,N_21785,N_21784);
nor U22151 (N_22151,N_21740,N_21927);
nor U22152 (N_22152,N_21934,N_21652);
xor U22153 (N_22153,N_21733,N_21993);
and U22154 (N_22154,N_21511,N_21698);
xor U22155 (N_22155,N_21832,N_21754);
or U22156 (N_22156,N_21588,N_21912);
nor U22157 (N_22157,N_21779,N_21942);
nand U22158 (N_22158,N_21528,N_21751);
nor U22159 (N_22159,N_21575,N_21787);
nand U22160 (N_22160,N_21975,N_21702);
and U22161 (N_22161,N_21759,N_21891);
xnor U22162 (N_22162,N_21977,N_21836);
or U22163 (N_22163,N_21806,N_21562);
xor U22164 (N_22164,N_21689,N_21713);
and U22165 (N_22165,N_21518,N_21948);
or U22166 (N_22166,N_21718,N_21982);
or U22167 (N_22167,N_21918,N_21743);
or U22168 (N_22168,N_21970,N_21887);
and U22169 (N_22169,N_21735,N_21568);
nor U22170 (N_22170,N_21522,N_21517);
nand U22171 (N_22171,N_21716,N_21853);
and U22172 (N_22172,N_21936,N_21782);
nand U22173 (N_22173,N_21760,N_21967);
xnor U22174 (N_22174,N_21914,N_21814);
or U22175 (N_22175,N_21725,N_21663);
nor U22176 (N_22176,N_21749,N_21667);
nor U22177 (N_22177,N_21539,N_21607);
nor U22178 (N_22178,N_21646,N_21987);
or U22179 (N_22179,N_21869,N_21981);
nor U22180 (N_22180,N_21783,N_21755);
and U22181 (N_22181,N_21536,N_21624);
nor U22182 (N_22182,N_21694,N_21966);
or U22183 (N_22183,N_21746,N_21964);
and U22184 (N_22184,N_21913,N_21766);
nor U22185 (N_22185,N_21564,N_21537);
nand U22186 (N_22186,N_21738,N_21839);
nor U22187 (N_22187,N_21761,N_21669);
xnor U22188 (N_22188,N_21625,N_21700);
xnor U22189 (N_22189,N_21858,N_21613);
nor U22190 (N_22190,N_21742,N_21772);
xor U22191 (N_22191,N_21866,N_21856);
xnor U22192 (N_22192,N_21906,N_21519);
nor U22193 (N_22193,N_21752,N_21556);
nand U22194 (N_22194,N_21540,N_21567);
or U22195 (N_22195,N_21897,N_21903);
nor U22196 (N_22196,N_21578,N_21796);
nor U22197 (N_22197,N_21632,N_21577);
and U22198 (N_22198,N_21576,N_21634);
or U22199 (N_22199,N_21643,N_21890);
xnor U22200 (N_22200,N_21988,N_21621);
or U22201 (N_22201,N_21845,N_21852);
nor U22202 (N_22202,N_21798,N_21642);
xnor U22203 (N_22203,N_21764,N_21805);
xnor U22204 (N_22204,N_21618,N_21668);
and U22205 (N_22205,N_21978,N_21681);
nand U22206 (N_22206,N_21765,N_21875);
nand U22207 (N_22207,N_21586,N_21688);
xor U22208 (N_22208,N_21874,N_21819);
nor U22209 (N_22209,N_21941,N_21695);
nor U22210 (N_22210,N_21800,N_21768);
nand U22211 (N_22211,N_21792,N_21762);
and U22212 (N_22212,N_21813,N_21963);
nor U22213 (N_22213,N_21538,N_21674);
nand U22214 (N_22214,N_21651,N_21841);
xnor U22215 (N_22215,N_21570,N_21958);
nor U22216 (N_22216,N_21923,N_21838);
and U22217 (N_22217,N_21710,N_21720);
or U22218 (N_22218,N_21799,N_21820);
nor U22219 (N_22219,N_21623,N_21665);
or U22220 (N_22220,N_21929,N_21660);
nand U22221 (N_22221,N_21545,N_21635);
nor U22222 (N_22222,N_21979,N_21904);
or U22223 (N_22223,N_21523,N_21589);
or U22224 (N_22224,N_21885,N_21520);
nand U22225 (N_22225,N_21892,N_21961);
or U22226 (N_22226,N_21723,N_21726);
or U22227 (N_22227,N_21561,N_21899);
or U22228 (N_22228,N_21579,N_21722);
xnor U22229 (N_22229,N_21846,N_21932);
nor U22230 (N_22230,N_21558,N_21953);
nand U22231 (N_22231,N_21605,N_21980);
xnor U22232 (N_22232,N_21944,N_21666);
nor U22233 (N_22233,N_21920,N_21821);
xor U22234 (N_22234,N_21587,N_21690);
nand U22235 (N_22235,N_21951,N_21992);
nor U22236 (N_22236,N_21871,N_21510);
xnor U22237 (N_22237,N_21724,N_21650);
xor U22238 (N_22238,N_21639,N_21939);
nand U22239 (N_22239,N_21757,N_21955);
or U22240 (N_22240,N_21928,N_21516);
nand U22241 (N_22241,N_21628,N_21555);
and U22242 (N_22242,N_21697,N_21748);
or U22243 (N_22243,N_21727,N_21907);
nor U22244 (N_22244,N_21731,N_21957);
and U22245 (N_22245,N_21882,N_21851);
nand U22246 (N_22246,N_21898,N_21554);
or U22247 (N_22247,N_21728,N_21995);
and U22248 (N_22248,N_21908,N_21739);
nand U22249 (N_22249,N_21859,N_21608);
or U22250 (N_22250,N_21568,N_21884);
nand U22251 (N_22251,N_21850,N_21825);
and U22252 (N_22252,N_21871,N_21704);
and U22253 (N_22253,N_21897,N_21990);
and U22254 (N_22254,N_21791,N_21656);
nor U22255 (N_22255,N_21829,N_21889);
nand U22256 (N_22256,N_21810,N_21958);
xnor U22257 (N_22257,N_21765,N_21927);
or U22258 (N_22258,N_21749,N_21563);
nor U22259 (N_22259,N_21940,N_21539);
and U22260 (N_22260,N_21792,N_21822);
and U22261 (N_22261,N_21907,N_21928);
nor U22262 (N_22262,N_21752,N_21822);
xor U22263 (N_22263,N_21517,N_21950);
and U22264 (N_22264,N_21866,N_21621);
xor U22265 (N_22265,N_21961,N_21568);
and U22266 (N_22266,N_21861,N_21959);
or U22267 (N_22267,N_21702,N_21544);
nor U22268 (N_22268,N_21562,N_21773);
xor U22269 (N_22269,N_21754,N_21516);
nor U22270 (N_22270,N_21940,N_21977);
nand U22271 (N_22271,N_21617,N_21805);
nand U22272 (N_22272,N_21818,N_21560);
nand U22273 (N_22273,N_21539,N_21722);
xor U22274 (N_22274,N_21607,N_21952);
xnor U22275 (N_22275,N_21937,N_21806);
nand U22276 (N_22276,N_21749,N_21566);
nor U22277 (N_22277,N_21587,N_21914);
xnor U22278 (N_22278,N_21757,N_21730);
or U22279 (N_22279,N_21535,N_21998);
nand U22280 (N_22280,N_21784,N_21835);
xnor U22281 (N_22281,N_21997,N_21862);
xnor U22282 (N_22282,N_21867,N_21957);
or U22283 (N_22283,N_21998,N_21519);
xor U22284 (N_22284,N_21862,N_21789);
xnor U22285 (N_22285,N_21832,N_21714);
nor U22286 (N_22286,N_21580,N_21921);
xnor U22287 (N_22287,N_21770,N_21871);
or U22288 (N_22288,N_21513,N_21865);
and U22289 (N_22289,N_21744,N_21693);
nand U22290 (N_22290,N_21510,N_21545);
or U22291 (N_22291,N_21705,N_21905);
or U22292 (N_22292,N_21716,N_21564);
xnor U22293 (N_22293,N_21568,N_21947);
nor U22294 (N_22294,N_21853,N_21634);
xnor U22295 (N_22295,N_21572,N_21651);
nand U22296 (N_22296,N_21944,N_21888);
nand U22297 (N_22297,N_21647,N_21923);
and U22298 (N_22298,N_21747,N_21517);
nand U22299 (N_22299,N_21616,N_21587);
xnor U22300 (N_22300,N_21513,N_21854);
nand U22301 (N_22301,N_21845,N_21678);
nor U22302 (N_22302,N_21855,N_21800);
xnor U22303 (N_22303,N_21797,N_21740);
nand U22304 (N_22304,N_21928,N_21950);
xnor U22305 (N_22305,N_21574,N_21516);
nand U22306 (N_22306,N_21628,N_21948);
nor U22307 (N_22307,N_21869,N_21831);
or U22308 (N_22308,N_21783,N_21641);
and U22309 (N_22309,N_21985,N_21638);
and U22310 (N_22310,N_21792,N_21761);
xor U22311 (N_22311,N_21775,N_21982);
or U22312 (N_22312,N_21649,N_21935);
xor U22313 (N_22313,N_21853,N_21977);
xnor U22314 (N_22314,N_21963,N_21936);
nand U22315 (N_22315,N_21754,N_21759);
nor U22316 (N_22316,N_21995,N_21757);
and U22317 (N_22317,N_21736,N_21805);
xnor U22318 (N_22318,N_21813,N_21681);
xnor U22319 (N_22319,N_21807,N_21940);
nand U22320 (N_22320,N_21668,N_21685);
xor U22321 (N_22321,N_21951,N_21568);
nand U22322 (N_22322,N_21735,N_21863);
nor U22323 (N_22323,N_21894,N_21656);
nand U22324 (N_22324,N_21566,N_21836);
xnor U22325 (N_22325,N_21733,N_21694);
or U22326 (N_22326,N_21548,N_21881);
or U22327 (N_22327,N_21780,N_21869);
and U22328 (N_22328,N_21778,N_21585);
xnor U22329 (N_22329,N_21760,N_21588);
nor U22330 (N_22330,N_21721,N_21854);
nand U22331 (N_22331,N_21723,N_21536);
nor U22332 (N_22332,N_21923,N_21679);
nand U22333 (N_22333,N_21921,N_21827);
xor U22334 (N_22334,N_21988,N_21932);
or U22335 (N_22335,N_21791,N_21758);
or U22336 (N_22336,N_21630,N_21545);
nor U22337 (N_22337,N_21613,N_21612);
or U22338 (N_22338,N_21962,N_21540);
nand U22339 (N_22339,N_21706,N_21720);
nor U22340 (N_22340,N_21831,N_21879);
nor U22341 (N_22341,N_21551,N_21684);
xor U22342 (N_22342,N_21918,N_21871);
and U22343 (N_22343,N_21691,N_21722);
nor U22344 (N_22344,N_21974,N_21841);
xnor U22345 (N_22345,N_21771,N_21547);
xor U22346 (N_22346,N_21988,N_21916);
xnor U22347 (N_22347,N_21534,N_21573);
or U22348 (N_22348,N_21996,N_21810);
nor U22349 (N_22349,N_21805,N_21993);
nor U22350 (N_22350,N_21884,N_21731);
xnor U22351 (N_22351,N_21930,N_21915);
nor U22352 (N_22352,N_21544,N_21807);
nand U22353 (N_22353,N_21767,N_21534);
nand U22354 (N_22354,N_21774,N_21666);
and U22355 (N_22355,N_21554,N_21641);
xnor U22356 (N_22356,N_21563,N_21854);
nor U22357 (N_22357,N_21790,N_21788);
xor U22358 (N_22358,N_21784,N_21510);
and U22359 (N_22359,N_21510,N_21531);
nor U22360 (N_22360,N_21641,N_21736);
or U22361 (N_22361,N_21676,N_21629);
xor U22362 (N_22362,N_21800,N_21888);
xnor U22363 (N_22363,N_21585,N_21885);
nor U22364 (N_22364,N_21710,N_21688);
xor U22365 (N_22365,N_21768,N_21554);
or U22366 (N_22366,N_21809,N_21938);
nor U22367 (N_22367,N_21903,N_21539);
nor U22368 (N_22368,N_21583,N_21959);
nand U22369 (N_22369,N_21661,N_21563);
nor U22370 (N_22370,N_21894,N_21751);
nand U22371 (N_22371,N_21659,N_21545);
nand U22372 (N_22372,N_21782,N_21572);
or U22373 (N_22373,N_21742,N_21589);
nor U22374 (N_22374,N_21833,N_21675);
and U22375 (N_22375,N_21693,N_21688);
nand U22376 (N_22376,N_21709,N_21983);
nor U22377 (N_22377,N_21525,N_21881);
nand U22378 (N_22378,N_21626,N_21941);
nor U22379 (N_22379,N_21587,N_21783);
and U22380 (N_22380,N_21870,N_21938);
or U22381 (N_22381,N_21658,N_21736);
nor U22382 (N_22382,N_21933,N_21576);
or U22383 (N_22383,N_21646,N_21720);
and U22384 (N_22384,N_21719,N_21521);
nand U22385 (N_22385,N_21618,N_21549);
nor U22386 (N_22386,N_21800,N_21569);
and U22387 (N_22387,N_21566,N_21771);
nor U22388 (N_22388,N_21643,N_21865);
and U22389 (N_22389,N_21831,N_21827);
and U22390 (N_22390,N_21625,N_21765);
nor U22391 (N_22391,N_21869,N_21942);
nand U22392 (N_22392,N_21639,N_21569);
or U22393 (N_22393,N_21597,N_21500);
or U22394 (N_22394,N_21966,N_21969);
or U22395 (N_22395,N_21805,N_21567);
nand U22396 (N_22396,N_21969,N_21675);
and U22397 (N_22397,N_21990,N_21746);
nand U22398 (N_22398,N_21619,N_21977);
xnor U22399 (N_22399,N_21950,N_21696);
nor U22400 (N_22400,N_21745,N_21575);
xnor U22401 (N_22401,N_21863,N_21813);
xor U22402 (N_22402,N_21825,N_21982);
nor U22403 (N_22403,N_21735,N_21971);
xor U22404 (N_22404,N_21707,N_21907);
or U22405 (N_22405,N_21884,N_21505);
nand U22406 (N_22406,N_21941,N_21592);
nand U22407 (N_22407,N_21916,N_21940);
nor U22408 (N_22408,N_21557,N_21914);
nor U22409 (N_22409,N_21587,N_21517);
and U22410 (N_22410,N_21540,N_21549);
nand U22411 (N_22411,N_21581,N_21915);
nor U22412 (N_22412,N_21527,N_21711);
and U22413 (N_22413,N_21809,N_21776);
nand U22414 (N_22414,N_21608,N_21942);
or U22415 (N_22415,N_21786,N_21700);
nand U22416 (N_22416,N_21989,N_21997);
and U22417 (N_22417,N_21889,N_21995);
and U22418 (N_22418,N_21710,N_21636);
or U22419 (N_22419,N_21794,N_21955);
nor U22420 (N_22420,N_21973,N_21833);
nor U22421 (N_22421,N_21842,N_21892);
nor U22422 (N_22422,N_21728,N_21544);
or U22423 (N_22423,N_21587,N_21710);
xnor U22424 (N_22424,N_21971,N_21893);
or U22425 (N_22425,N_21613,N_21840);
nor U22426 (N_22426,N_21755,N_21636);
and U22427 (N_22427,N_21548,N_21924);
and U22428 (N_22428,N_21765,N_21565);
nand U22429 (N_22429,N_21844,N_21935);
xor U22430 (N_22430,N_21705,N_21861);
or U22431 (N_22431,N_21637,N_21680);
nor U22432 (N_22432,N_21512,N_21962);
nor U22433 (N_22433,N_21789,N_21653);
and U22434 (N_22434,N_21733,N_21510);
and U22435 (N_22435,N_21722,N_21840);
and U22436 (N_22436,N_21611,N_21855);
and U22437 (N_22437,N_21785,N_21662);
nor U22438 (N_22438,N_21670,N_21615);
or U22439 (N_22439,N_21729,N_21536);
and U22440 (N_22440,N_21798,N_21614);
or U22441 (N_22441,N_21839,N_21838);
or U22442 (N_22442,N_21524,N_21546);
or U22443 (N_22443,N_21565,N_21789);
nand U22444 (N_22444,N_21509,N_21752);
xor U22445 (N_22445,N_21889,N_21685);
nor U22446 (N_22446,N_21822,N_21970);
nor U22447 (N_22447,N_21536,N_21628);
or U22448 (N_22448,N_21646,N_21855);
and U22449 (N_22449,N_21842,N_21669);
or U22450 (N_22450,N_21537,N_21563);
nor U22451 (N_22451,N_21711,N_21842);
or U22452 (N_22452,N_21802,N_21957);
xnor U22453 (N_22453,N_21745,N_21867);
and U22454 (N_22454,N_21800,N_21930);
xnor U22455 (N_22455,N_21536,N_21688);
and U22456 (N_22456,N_21635,N_21810);
nand U22457 (N_22457,N_21760,N_21968);
xor U22458 (N_22458,N_21670,N_21862);
nor U22459 (N_22459,N_21756,N_21501);
nor U22460 (N_22460,N_21946,N_21798);
xor U22461 (N_22461,N_21893,N_21901);
nor U22462 (N_22462,N_21860,N_21769);
and U22463 (N_22463,N_21858,N_21835);
or U22464 (N_22464,N_21694,N_21998);
nor U22465 (N_22465,N_21549,N_21639);
and U22466 (N_22466,N_21534,N_21871);
nand U22467 (N_22467,N_21933,N_21716);
or U22468 (N_22468,N_21825,N_21669);
or U22469 (N_22469,N_21968,N_21644);
nor U22470 (N_22470,N_21790,N_21548);
xnor U22471 (N_22471,N_21693,N_21922);
nand U22472 (N_22472,N_21759,N_21762);
nand U22473 (N_22473,N_21760,N_21851);
nor U22474 (N_22474,N_21939,N_21754);
and U22475 (N_22475,N_21823,N_21779);
and U22476 (N_22476,N_21615,N_21828);
or U22477 (N_22477,N_21938,N_21775);
or U22478 (N_22478,N_21796,N_21589);
and U22479 (N_22479,N_21872,N_21636);
nand U22480 (N_22480,N_21700,N_21922);
nor U22481 (N_22481,N_21699,N_21600);
or U22482 (N_22482,N_21517,N_21741);
xor U22483 (N_22483,N_21966,N_21618);
and U22484 (N_22484,N_21648,N_21675);
and U22485 (N_22485,N_21699,N_21576);
or U22486 (N_22486,N_21959,N_21960);
xor U22487 (N_22487,N_21539,N_21945);
and U22488 (N_22488,N_21511,N_21651);
nand U22489 (N_22489,N_21715,N_21986);
nand U22490 (N_22490,N_21677,N_21510);
and U22491 (N_22491,N_21752,N_21517);
or U22492 (N_22492,N_21995,N_21960);
xnor U22493 (N_22493,N_21768,N_21765);
nor U22494 (N_22494,N_21827,N_21751);
nand U22495 (N_22495,N_21789,N_21930);
and U22496 (N_22496,N_21959,N_21770);
and U22497 (N_22497,N_21611,N_21504);
xnor U22498 (N_22498,N_21682,N_21786);
nor U22499 (N_22499,N_21887,N_21876);
nor U22500 (N_22500,N_22117,N_22250);
and U22501 (N_22501,N_22150,N_22194);
or U22502 (N_22502,N_22335,N_22091);
or U22503 (N_22503,N_22306,N_22222);
and U22504 (N_22504,N_22493,N_22039);
xor U22505 (N_22505,N_22234,N_22143);
nand U22506 (N_22506,N_22040,N_22427);
and U22507 (N_22507,N_22063,N_22497);
xnor U22508 (N_22508,N_22221,N_22456);
or U22509 (N_22509,N_22321,N_22320);
xor U22510 (N_22510,N_22113,N_22011);
xor U22511 (N_22511,N_22488,N_22440);
xor U22512 (N_22512,N_22359,N_22027);
nor U22513 (N_22513,N_22471,N_22316);
and U22514 (N_22514,N_22036,N_22002);
xor U22515 (N_22515,N_22298,N_22302);
xor U22516 (N_22516,N_22024,N_22156);
xor U22517 (N_22517,N_22209,N_22429);
nor U22518 (N_22518,N_22311,N_22420);
xor U22519 (N_22519,N_22430,N_22025);
and U22520 (N_22520,N_22394,N_22152);
xnor U22521 (N_22521,N_22477,N_22189);
nand U22522 (N_22522,N_22075,N_22203);
and U22523 (N_22523,N_22325,N_22148);
and U22524 (N_22524,N_22305,N_22214);
nand U22525 (N_22525,N_22317,N_22399);
nand U22526 (N_22526,N_22049,N_22242);
and U22527 (N_22527,N_22251,N_22193);
or U22528 (N_22528,N_22228,N_22092);
xnor U22529 (N_22529,N_22386,N_22123);
and U22530 (N_22530,N_22205,N_22131);
nand U22531 (N_22531,N_22391,N_22437);
xnor U22532 (N_22532,N_22147,N_22486);
and U22533 (N_22533,N_22196,N_22366);
or U22534 (N_22534,N_22031,N_22277);
nand U22535 (N_22535,N_22385,N_22243);
or U22536 (N_22536,N_22273,N_22454);
xor U22537 (N_22537,N_22238,N_22411);
xor U22538 (N_22538,N_22248,N_22389);
and U22539 (N_22539,N_22047,N_22481);
xnor U22540 (N_22540,N_22354,N_22499);
or U22541 (N_22541,N_22278,N_22169);
or U22542 (N_22542,N_22183,N_22216);
nand U22543 (N_22543,N_22101,N_22443);
nand U22544 (N_22544,N_22431,N_22478);
and U22545 (N_22545,N_22457,N_22281);
nor U22546 (N_22546,N_22037,N_22467);
or U22547 (N_22547,N_22190,N_22247);
or U22548 (N_22548,N_22496,N_22022);
and U22549 (N_22549,N_22262,N_22107);
and U22550 (N_22550,N_22468,N_22142);
nand U22551 (N_22551,N_22406,N_22367);
nor U22552 (N_22552,N_22404,N_22177);
or U22553 (N_22553,N_22065,N_22292);
nand U22554 (N_22554,N_22276,N_22180);
nor U22555 (N_22555,N_22265,N_22151);
nand U22556 (N_22556,N_22185,N_22097);
nand U22557 (N_22557,N_22034,N_22163);
and U22558 (N_22558,N_22108,N_22257);
nand U22559 (N_22559,N_22446,N_22327);
nor U22560 (N_22560,N_22412,N_22450);
xor U22561 (N_22561,N_22199,N_22057);
nand U22562 (N_22562,N_22046,N_22200);
and U22563 (N_22563,N_22170,N_22332);
and U22564 (N_22564,N_22013,N_22353);
or U22565 (N_22565,N_22224,N_22361);
or U22566 (N_22566,N_22282,N_22048);
and U22567 (N_22567,N_22043,N_22233);
xnor U22568 (N_22568,N_22225,N_22279);
or U22569 (N_22569,N_22266,N_22198);
nor U22570 (N_22570,N_22307,N_22355);
and U22571 (N_22571,N_22470,N_22283);
nand U22572 (N_22572,N_22474,N_22186);
xor U22573 (N_22573,N_22280,N_22442);
nor U22574 (N_22574,N_22270,N_22241);
xnor U22575 (N_22575,N_22181,N_22017);
or U22576 (N_22576,N_22398,N_22349);
nand U22577 (N_22577,N_22469,N_22275);
nand U22578 (N_22578,N_22121,N_22313);
and U22579 (N_22579,N_22329,N_22340);
xnor U22580 (N_22580,N_22094,N_22319);
nand U22581 (N_22581,N_22338,N_22295);
nand U22582 (N_22582,N_22482,N_22415);
nor U22583 (N_22583,N_22370,N_22378);
nor U22584 (N_22584,N_22004,N_22284);
nor U22585 (N_22585,N_22447,N_22333);
and U22586 (N_22586,N_22328,N_22105);
xor U22587 (N_22587,N_22259,N_22462);
xnor U22588 (N_22588,N_22168,N_22347);
or U22589 (N_22589,N_22083,N_22124);
nand U22590 (N_22590,N_22115,N_22051);
or U22591 (N_22591,N_22261,N_22165);
xnor U22592 (N_22592,N_22035,N_22171);
nand U22593 (N_22593,N_22345,N_22155);
xnor U22594 (N_22594,N_22461,N_22357);
nor U22595 (N_22595,N_22096,N_22324);
and U22596 (N_22596,N_22393,N_22245);
nand U22597 (N_22597,N_22045,N_22291);
nor U22598 (N_22598,N_22483,N_22460);
nor U22599 (N_22599,N_22387,N_22237);
xnor U22600 (N_22600,N_22087,N_22294);
xor U22601 (N_22601,N_22009,N_22079);
or U22602 (N_22602,N_22490,N_22230);
xor U22603 (N_22603,N_22111,N_22114);
nor U22604 (N_22604,N_22217,N_22435);
nor U22605 (N_22605,N_22133,N_22487);
nor U22606 (N_22606,N_22000,N_22479);
nand U22607 (N_22607,N_22498,N_22289);
or U22608 (N_22608,N_22365,N_22069);
xor U22609 (N_22609,N_22167,N_22402);
xnor U22610 (N_22610,N_22020,N_22272);
nor U22611 (N_22611,N_22158,N_22119);
and U22612 (N_22612,N_22060,N_22232);
and U22613 (N_22613,N_22129,N_22323);
and U22614 (N_22614,N_22231,N_22130);
and U22615 (N_22615,N_22244,N_22380);
nor U22616 (N_22616,N_22226,N_22064);
and U22617 (N_22617,N_22463,N_22179);
or U22618 (N_22618,N_22016,N_22010);
nand U22619 (N_22619,N_22356,N_22384);
xnor U22620 (N_22620,N_22476,N_22297);
xor U22621 (N_22621,N_22007,N_22350);
and U22622 (N_22622,N_22055,N_22269);
or U22623 (N_22623,N_22014,N_22473);
xor U22624 (N_22624,N_22346,N_22392);
nand U22625 (N_22625,N_22006,N_22246);
xor U22626 (N_22626,N_22058,N_22202);
and U22627 (N_22627,N_22080,N_22466);
nor U22628 (N_22628,N_22138,N_22418);
and U22629 (N_22629,N_22070,N_22128);
nor U22630 (N_22630,N_22422,N_22134);
nand U22631 (N_22631,N_22197,N_22489);
and U22632 (N_22632,N_22274,N_22012);
xnor U22633 (N_22633,N_22348,N_22458);
xor U22634 (N_22634,N_22368,N_22396);
xor U22635 (N_22635,N_22459,N_22360);
or U22636 (N_22636,N_22373,N_22369);
xor U22637 (N_22637,N_22254,N_22088);
nand U22638 (N_22638,N_22029,N_22372);
and U22639 (N_22639,N_22304,N_22344);
xor U22640 (N_22640,N_22136,N_22425);
or U22641 (N_22641,N_22352,N_22417);
or U22642 (N_22642,N_22213,N_22008);
and U22643 (N_22643,N_22212,N_22076);
or U22644 (N_22644,N_22139,N_22407);
xnor U22645 (N_22645,N_22082,N_22001);
and U22646 (N_22646,N_22364,N_22495);
nor U22647 (N_22647,N_22052,N_22268);
nand U22648 (N_22648,N_22240,N_22256);
nand U22649 (N_22649,N_22375,N_22044);
xnor U22650 (N_22650,N_22475,N_22410);
and U22651 (N_22651,N_22426,N_22061);
or U22652 (N_22652,N_22068,N_22218);
nor U22653 (N_22653,N_22314,N_22465);
nor U22654 (N_22654,N_22102,N_22067);
xor U22655 (N_22655,N_22383,N_22098);
nor U22656 (N_22656,N_22062,N_22397);
xor U22657 (N_22657,N_22419,N_22144);
xnor U22658 (N_22658,N_22374,N_22099);
and U22659 (N_22659,N_22452,N_22405);
or U22660 (N_22660,N_22227,N_22100);
or U22661 (N_22661,N_22301,N_22249);
and U22662 (N_22662,N_22191,N_22444);
nand U22663 (N_22663,N_22433,N_22491);
xor U22664 (N_22664,N_22267,N_22445);
xor U22665 (N_22665,N_22153,N_22195);
nand U22666 (N_22666,N_22343,N_22160);
nor U22667 (N_22667,N_22073,N_22140);
xor U22668 (N_22668,N_22236,N_22146);
and U22669 (N_22669,N_22395,N_22161);
nor U22670 (N_22670,N_22336,N_22137);
and U22671 (N_22671,N_22494,N_22176);
nand U22672 (N_22672,N_22184,N_22201);
nor U22673 (N_22673,N_22086,N_22315);
nand U22674 (N_22674,N_22164,N_22229);
xnor U22675 (N_22675,N_22288,N_22263);
or U22676 (N_22676,N_22449,N_22204);
or U22677 (N_22677,N_22220,N_22414);
and U22678 (N_22678,N_22172,N_22235);
and U22679 (N_22679,N_22066,N_22434);
and U22680 (N_22680,N_22110,N_22125);
xor U22681 (N_22681,N_22223,N_22041);
and U22682 (N_22682,N_22211,N_22215);
xor U22683 (N_22683,N_22030,N_22472);
nand U22684 (N_22684,N_22326,N_22341);
or U22685 (N_22685,N_22382,N_22182);
nor U22686 (N_22686,N_22059,N_22145);
nor U22687 (N_22687,N_22089,N_22015);
or U22688 (N_22688,N_22166,N_22300);
nor U22689 (N_22689,N_22285,N_22255);
and U22690 (N_22690,N_22403,N_22453);
or U22691 (N_22691,N_22331,N_22492);
nor U22692 (N_22692,N_22077,N_22293);
xnor U22693 (N_22693,N_22071,N_22056);
xor U22694 (N_22694,N_22485,N_22095);
and U22695 (N_22695,N_22400,N_22308);
nand U22696 (N_22696,N_22120,N_22388);
xnor U22697 (N_22697,N_22376,N_22154);
nand U22698 (N_22698,N_22309,N_22090);
nand U22699 (N_22699,N_22358,N_22424);
nand U22700 (N_22700,N_22296,N_22312);
and U22701 (N_22701,N_22074,N_22042);
or U22702 (N_22702,N_22408,N_22413);
nand U22703 (N_22703,N_22239,N_22038);
and U22704 (N_22704,N_22078,N_22050);
and U22705 (N_22705,N_22260,N_22157);
nor U22706 (N_22706,N_22126,N_22173);
or U22707 (N_22707,N_22390,N_22109);
or U22708 (N_22708,N_22085,N_22416);
nor U22709 (N_22709,N_22026,N_22421);
nor U22710 (N_22710,N_22342,N_22188);
nor U22711 (N_22711,N_22330,N_22318);
nor U22712 (N_22712,N_22381,N_22351);
xor U22713 (N_22713,N_22003,N_22093);
or U22714 (N_22714,N_22286,N_22428);
or U22715 (N_22715,N_22103,N_22409);
or U22716 (N_22716,N_22322,N_22337);
nand U22717 (N_22717,N_22303,N_22019);
xor U22718 (N_22718,N_22192,N_22290);
and U22719 (N_22719,N_22174,N_22438);
or U22720 (N_22720,N_22118,N_22028);
xor U22721 (N_22721,N_22432,N_22271);
xnor U22722 (N_22722,N_22210,N_22362);
nand U22723 (N_22723,N_22464,N_22439);
or U22724 (N_22724,N_22299,N_22423);
xnor U22725 (N_22725,N_22219,N_22448);
or U22726 (N_22726,N_22401,N_22178);
xor U22727 (N_22727,N_22116,N_22106);
xor U22728 (N_22728,N_22451,N_22310);
and U22729 (N_22729,N_22053,N_22371);
xnor U22730 (N_22730,N_22339,N_22363);
or U22731 (N_22731,N_22112,N_22122);
xor U22732 (N_22732,N_22377,N_22258);
and U22733 (N_22733,N_22480,N_22441);
and U22734 (N_22734,N_22253,N_22072);
xnor U22735 (N_22735,N_22436,N_22207);
nor U22736 (N_22736,N_22054,N_22132);
xnor U22737 (N_22737,N_22033,N_22018);
nor U22738 (N_22738,N_22334,N_22127);
xnor U22739 (N_22739,N_22023,N_22206);
nand U22740 (N_22740,N_22455,N_22162);
nand U22741 (N_22741,N_22484,N_22104);
or U22742 (N_22742,N_22141,N_22187);
xnor U22743 (N_22743,N_22081,N_22135);
nand U22744 (N_22744,N_22208,N_22021);
nor U22745 (N_22745,N_22032,N_22252);
nor U22746 (N_22746,N_22379,N_22005);
xor U22747 (N_22747,N_22264,N_22084);
nand U22748 (N_22748,N_22175,N_22159);
and U22749 (N_22749,N_22287,N_22149);
or U22750 (N_22750,N_22371,N_22295);
or U22751 (N_22751,N_22413,N_22080);
nor U22752 (N_22752,N_22152,N_22446);
or U22753 (N_22753,N_22268,N_22049);
xor U22754 (N_22754,N_22090,N_22103);
xnor U22755 (N_22755,N_22140,N_22184);
and U22756 (N_22756,N_22117,N_22100);
nor U22757 (N_22757,N_22450,N_22125);
xnor U22758 (N_22758,N_22092,N_22027);
or U22759 (N_22759,N_22287,N_22081);
or U22760 (N_22760,N_22326,N_22141);
xnor U22761 (N_22761,N_22494,N_22499);
xnor U22762 (N_22762,N_22304,N_22237);
or U22763 (N_22763,N_22427,N_22206);
and U22764 (N_22764,N_22379,N_22169);
and U22765 (N_22765,N_22463,N_22070);
and U22766 (N_22766,N_22230,N_22382);
and U22767 (N_22767,N_22174,N_22314);
and U22768 (N_22768,N_22067,N_22142);
nand U22769 (N_22769,N_22236,N_22474);
or U22770 (N_22770,N_22203,N_22236);
and U22771 (N_22771,N_22383,N_22408);
nor U22772 (N_22772,N_22179,N_22002);
or U22773 (N_22773,N_22492,N_22273);
nor U22774 (N_22774,N_22296,N_22089);
or U22775 (N_22775,N_22207,N_22387);
nand U22776 (N_22776,N_22171,N_22450);
xor U22777 (N_22777,N_22401,N_22472);
or U22778 (N_22778,N_22200,N_22131);
and U22779 (N_22779,N_22049,N_22017);
or U22780 (N_22780,N_22414,N_22300);
xnor U22781 (N_22781,N_22347,N_22034);
xnor U22782 (N_22782,N_22190,N_22011);
nand U22783 (N_22783,N_22305,N_22404);
nand U22784 (N_22784,N_22363,N_22443);
or U22785 (N_22785,N_22306,N_22341);
and U22786 (N_22786,N_22132,N_22319);
and U22787 (N_22787,N_22485,N_22047);
nand U22788 (N_22788,N_22334,N_22343);
nand U22789 (N_22789,N_22179,N_22137);
xor U22790 (N_22790,N_22171,N_22394);
xnor U22791 (N_22791,N_22433,N_22126);
nand U22792 (N_22792,N_22220,N_22020);
and U22793 (N_22793,N_22476,N_22463);
nor U22794 (N_22794,N_22205,N_22407);
nor U22795 (N_22795,N_22201,N_22352);
and U22796 (N_22796,N_22298,N_22155);
nand U22797 (N_22797,N_22398,N_22266);
and U22798 (N_22798,N_22318,N_22373);
nor U22799 (N_22799,N_22237,N_22267);
nand U22800 (N_22800,N_22006,N_22157);
xor U22801 (N_22801,N_22124,N_22181);
or U22802 (N_22802,N_22090,N_22480);
xnor U22803 (N_22803,N_22429,N_22205);
and U22804 (N_22804,N_22148,N_22488);
nand U22805 (N_22805,N_22023,N_22311);
or U22806 (N_22806,N_22118,N_22101);
nor U22807 (N_22807,N_22057,N_22200);
nand U22808 (N_22808,N_22285,N_22389);
xor U22809 (N_22809,N_22141,N_22484);
nand U22810 (N_22810,N_22038,N_22371);
and U22811 (N_22811,N_22459,N_22135);
or U22812 (N_22812,N_22349,N_22334);
nand U22813 (N_22813,N_22367,N_22038);
nor U22814 (N_22814,N_22433,N_22455);
nand U22815 (N_22815,N_22334,N_22398);
and U22816 (N_22816,N_22333,N_22095);
or U22817 (N_22817,N_22150,N_22246);
xnor U22818 (N_22818,N_22088,N_22189);
or U22819 (N_22819,N_22195,N_22021);
and U22820 (N_22820,N_22301,N_22205);
xnor U22821 (N_22821,N_22069,N_22385);
xor U22822 (N_22822,N_22113,N_22340);
or U22823 (N_22823,N_22183,N_22137);
xnor U22824 (N_22824,N_22093,N_22145);
and U22825 (N_22825,N_22114,N_22193);
or U22826 (N_22826,N_22490,N_22248);
or U22827 (N_22827,N_22316,N_22119);
nor U22828 (N_22828,N_22202,N_22318);
and U22829 (N_22829,N_22217,N_22211);
or U22830 (N_22830,N_22006,N_22410);
nand U22831 (N_22831,N_22132,N_22258);
and U22832 (N_22832,N_22475,N_22354);
and U22833 (N_22833,N_22115,N_22483);
and U22834 (N_22834,N_22291,N_22265);
xnor U22835 (N_22835,N_22337,N_22030);
nand U22836 (N_22836,N_22177,N_22133);
and U22837 (N_22837,N_22495,N_22137);
nand U22838 (N_22838,N_22348,N_22450);
xnor U22839 (N_22839,N_22458,N_22077);
and U22840 (N_22840,N_22246,N_22152);
or U22841 (N_22841,N_22041,N_22367);
nor U22842 (N_22842,N_22029,N_22358);
or U22843 (N_22843,N_22200,N_22000);
nor U22844 (N_22844,N_22361,N_22257);
nand U22845 (N_22845,N_22146,N_22416);
xnor U22846 (N_22846,N_22459,N_22204);
xnor U22847 (N_22847,N_22370,N_22189);
nand U22848 (N_22848,N_22008,N_22032);
xor U22849 (N_22849,N_22097,N_22094);
nor U22850 (N_22850,N_22319,N_22081);
and U22851 (N_22851,N_22380,N_22190);
or U22852 (N_22852,N_22312,N_22111);
or U22853 (N_22853,N_22084,N_22034);
nor U22854 (N_22854,N_22424,N_22299);
nand U22855 (N_22855,N_22383,N_22236);
and U22856 (N_22856,N_22217,N_22141);
nor U22857 (N_22857,N_22248,N_22051);
nor U22858 (N_22858,N_22052,N_22418);
nor U22859 (N_22859,N_22146,N_22097);
or U22860 (N_22860,N_22288,N_22154);
nor U22861 (N_22861,N_22335,N_22196);
nor U22862 (N_22862,N_22032,N_22272);
and U22863 (N_22863,N_22093,N_22265);
nor U22864 (N_22864,N_22138,N_22424);
and U22865 (N_22865,N_22142,N_22079);
or U22866 (N_22866,N_22001,N_22114);
and U22867 (N_22867,N_22102,N_22418);
nor U22868 (N_22868,N_22465,N_22478);
nor U22869 (N_22869,N_22413,N_22487);
xor U22870 (N_22870,N_22462,N_22226);
nand U22871 (N_22871,N_22466,N_22220);
nand U22872 (N_22872,N_22019,N_22135);
or U22873 (N_22873,N_22143,N_22169);
and U22874 (N_22874,N_22208,N_22419);
nand U22875 (N_22875,N_22136,N_22130);
nor U22876 (N_22876,N_22061,N_22416);
nor U22877 (N_22877,N_22123,N_22226);
or U22878 (N_22878,N_22110,N_22324);
and U22879 (N_22879,N_22051,N_22289);
xnor U22880 (N_22880,N_22167,N_22314);
or U22881 (N_22881,N_22085,N_22435);
and U22882 (N_22882,N_22466,N_22273);
nand U22883 (N_22883,N_22412,N_22394);
nand U22884 (N_22884,N_22494,N_22424);
nor U22885 (N_22885,N_22242,N_22206);
xnor U22886 (N_22886,N_22058,N_22377);
nor U22887 (N_22887,N_22479,N_22210);
nand U22888 (N_22888,N_22467,N_22261);
nor U22889 (N_22889,N_22374,N_22227);
or U22890 (N_22890,N_22329,N_22061);
nand U22891 (N_22891,N_22013,N_22086);
or U22892 (N_22892,N_22258,N_22341);
and U22893 (N_22893,N_22211,N_22334);
xor U22894 (N_22894,N_22010,N_22385);
nand U22895 (N_22895,N_22166,N_22092);
or U22896 (N_22896,N_22090,N_22370);
nor U22897 (N_22897,N_22328,N_22068);
nand U22898 (N_22898,N_22364,N_22460);
nand U22899 (N_22899,N_22019,N_22279);
xnor U22900 (N_22900,N_22407,N_22125);
and U22901 (N_22901,N_22242,N_22250);
nand U22902 (N_22902,N_22447,N_22187);
and U22903 (N_22903,N_22168,N_22286);
and U22904 (N_22904,N_22126,N_22318);
nand U22905 (N_22905,N_22315,N_22059);
nand U22906 (N_22906,N_22266,N_22354);
nand U22907 (N_22907,N_22277,N_22222);
nor U22908 (N_22908,N_22349,N_22123);
and U22909 (N_22909,N_22444,N_22264);
nor U22910 (N_22910,N_22296,N_22227);
or U22911 (N_22911,N_22399,N_22245);
xnor U22912 (N_22912,N_22366,N_22470);
or U22913 (N_22913,N_22359,N_22398);
or U22914 (N_22914,N_22109,N_22302);
and U22915 (N_22915,N_22447,N_22218);
or U22916 (N_22916,N_22022,N_22247);
nand U22917 (N_22917,N_22230,N_22142);
nand U22918 (N_22918,N_22136,N_22038);
nand U22919 (N_22919,N_22220,N_22208);
and U22920 (N_22920,N_22267,N_22366);
or U22921 (N_22921,N_22396,N_22304);
and U22922 (N_22922,N_22490,N_22292);
and U22923 (N_22923,N_22057,N_22289);
nor U22924 (N_22924,N_22287,N_22489);
or U22925 (N_22925,N_22324,N_22472);
nand U22926 (N_22926,N_22198,N_22445);
nand U22927 (N_22927,N_22343,N_22117);
nand U22928 (N_22928,N_22068,N_22298);
xnor U22929 (N_22929,N_22053,N_22138);
nand U22930 (N_22930,N_22271,N_22086);
nand U22931 (N_22931,N_22217,N_22232);
nand U22932 (N_22932,N_22312,N_22171);
xnor U22933 (N_22933,N_22438,N_22059);
xor U22934 (N_22934,N_22472,N_22053);
nand U22935 (N_22935,N_22032,N_22109);
or U22936 (N_22936,N_22285,N_22147);
or U22937 (N_22937,N_22239,N_22400);
nand U22938 (N_22938,N_22367,N_22473);
and U22939 (N_22939,N_22239,N_22348);
or U22940 (N_22940,N_22044,N_22108);
nor U22941 (N_22941,N_22476,N_22027);
nand U22942 (N_22942,N_22236,N_22283);
xnor U22943 (N_22943,N_22079,N_22032);
nand U22944 (N_22944,N_22497,N_22177);
xor U22945 (N_22945,N_22094,N_22227);
and U22946 (N_22946,N_22100,N_22478);
and U22947 (N_22947,N_22108,N_22418);
or U22948 (N_22948,N_22280,N_22371);
nand U22949 (N_22949,N_22105,N_22020);
xor U22950 (N_22950,N_22303,N_22199);
or U22951 (N_22951,N_22183,N_22396);
or U22952 (N_22952,N_22033,N_22015);
nor U22953 (N_22953,N_22012,N_22340);
nand U22954 (N_22954,N_22266,N_22128);
nor U22955 (N_22955,N_22420,N_22161);
or U22956 (N_22956,N_22479,N_22161);
xor U22957 (N_22957,N_22194,N_22057);
nand U22958 (N_22958,N_22481,N_22410);
xnor U22959 (N_22959,N_22173,N_22424);
nor U22960 (N_22960,N_22009,N_22389);
nor U22961 (N_22961,N_22025,N_22016);
nor U22962 (N_22962,N_22447,N_22114);
or U22963 (N_22963,N_22185,N_22392);
and U22964 (N_22964,N_22027,N_22186);
xnor U22965 (N_22965,N_22379,N_22406);
and U22966 (N_22966,N_22368,N_22241);
nor U22967 (N_22967,N_22122,N_22057);
xnor U22968 (N_22968,N_22023,N_22304);
and U22969 (N_22969,N_22412,N_22335);
xor U22970 (N_22970,N_22337,N_22188);
nand U22971 (N_22971,N_22164,N_22116);
nor U22972 (N_22972,N_22234,N_22272);
nand U22973 (N_22973,N_22403,N_22366);
xor U22974 (N_22974,N_22283,N_22060);
or U22975 (N_22975,N_22092,N_22288);
or U22976 (N_22976,N_22300,N_22314);
nand U22977 (N_22977,N_22383,N_22252);
and U22978 (N_22978,N_22261,N_22281);
or U22979 (N_22979,N_22158,N_22278);
nand U22980 (N_22980,N_22375,N_22083);
and U22981 (N_22981,N_22072,N_22158);
nand U22982 (N_22982,N_22084,N_22335);
and U22983 (N_22983,N_22363,N_22412);
nor U22984 (N_22984,N_22040,N_22094);
or U22985 (N_22985,N_22327,N_22358);
or U22986 (N_22986,N_22157,N_22437);
or U22987 (N_22987,N_22247,N_22015);
nor U22988 (N_22988,N_22336,N_22154);
xor U22989 (N_22989,N_22383,N_22006);
nand U22990 (N_22990,N_22235,N_22213);
or U22991 (N_22991,N_22222,N_22208);
nand U22992 (N_22992,N_22117,N_22176);
and U22993 (N_22993,N_22251,N_22206);
nand U22994 (N_22994,N_22166,N_22291);
nor U22995 (N_22995,N_22028,N_22299);
or U22996 (N_22996,N_22246,N_22327);
xor U22997 (N_22997,N_22023,N_22138);
and U22998 (N_22998,N_22062,N_22101);
xnor U22999 (N_22999,N_22171,N_22065);
or U23000 (N_23000,N_22944,N_22892);
and U23001 (N_23001,N_22950,N_22551);
and U23002 (N_23002,N_22541,N_22882);
nor U23003 (N_23003,N_22609,N_22756);
or U23004 (N_23004,N_22770,N_22643);
or U23005 (N_23005,N_22764,N_22560);
and U23006 (N_23006,N_22718,N_22947);
nand U23007 (N_23007,N_22624,N_22530);
and U23008 (N_23008,N_22837,N_22728);
or U23009 (N_23009,N_22729,N_22863);
and U23010 (N_23010,N_22675,N_22594);
nor U23011 (N_23011,N_22960,N_22716);
and U23012 (N_23012,N_22612,N_22853);
and U23013 (N_23013,N_22784,N_22719);
xor U23014 (N_23014,N_22569,N_22688);
nand U23015 (N_23015,N_22650,N_22649);
or U23016 (N_23016,N_22741,N_22606);
or U23017 (N_23017,N_22752,N_22802);
nor U23018 (N_23018,N_22740,N_22768);
or U23019 (N_23019,N_22785,N_22634);
or U23020 (N_23020,N_22655,N_22885);
nand U23021 (N_23021,N_22544,N_22769);
or U23022 (N_23022,N_22907,N_22897);
nor U23023 (N_23023,N_22818,N_22576);
nand U23024 (N_23024,N_22988,N_22889);
and U23025 (N_23025,N_22851,N_22521);
xnor U23026 (N_23026,N_22659,N_22502);
nand U23027 (N_23027,N_22873,N_22581);
nor U23028 (N_23028,N_22974,N_22758);
nor U23029 (N_23029,N_22565,N_22674);
nor U23030 (N_23030,N_22777,N_22538);
and U23031 (N_23031,N_22958,N_22680);
nand U23032 (N_23032,N_22839,N_22696);
xor U23033 (N_23033,N_22791,N_22886);
and U23034 (N_23034,N_22899,N_22671);
or U23035 (N_23035,N_22668,N_22525);
xnor U23036 (N_23036,N_22685,N_22826);
nand U23037 (N_23037,N_22898,N_22879);
xor U23038 (N_23038,N_22605,N_22985);
and U23039 (N_23039,N_22698,N_22938);
and U23040 (N_23040,N_22509,N_22996);
and U23041 (N_23041,N_22809,N_22963);
nor U23042 (N_23042,N_22788,N_22794);
and U23043 (N_23043,N_22989,N_22514);
xnor U23044 (N_23044,N_22919,N_22844);
and U23045 (N_23045,N_22939,N_22694);
xnor U23046 (N_23046,N_22547,N_22902);
xnor U23047 (N_23047,N_22692,N_22591);
and U23048 (N_23048,N_22700,N_22817);
nand U23049 (N_23049,N_22949,N_22792);
and U23050 (N_23050,N_22793,N_22747);
nand U23051 (N_23051,N_22867,N_22656);
xnor U23052 (N_23052,N_22570,N_22723);
nand U23053 (N_23053,N_22790,N_22962);
or U23054 (N_23054,N_22652,N_22568);
xor U23055 (N_23055,N_22579,N_22539);
and U23056 (N_23056,N_22614,N_22970);
and U23057 (N_23057,N_22776,N_22725);
or U23058 (N_23058,N_22517,N_22673);
and U23059 (N_23059,N_22724,N_22819);
nor U23060 (N_23060,N_22744,N_22981);
or U23061 (N_23061,N_22556,N_22992);
and U23062 (N_23062,N_22636,N_22935);
and U23063 (N_23063,N_22534,N_22778);
or U23064 (N_23064,N_22625,N_22717);
or U23065 (N_23065,N_22693,N_22558);
xnor U23066 (N_23066,N_22904,N_22987);
or U23067 (N_23067,N_22850,N_22795);
xnor U23068 (N_23068,N_22535,N_22861);
nor U23069 (N_23069,N_22948,N_22608);
xnor U23070 (N_23070,N_22805,N_22513);
or U23071 (N_23071,N_22500,N_22875);
nand U23072 (N_23072,N_22925,N_22618);
xnor U23073 (N_23073,N_22504,N_22516);
and U23074 (N_23074,N_22829,N_22707);
and U23075 (N_23075,N_22884,N_22661);
nand U23076 (N_23076,N_22737,N_22732);
and U23077 (N_23077,N_22592,N_22953);
or U23078 (N_23078,N_22520,N_22677);
and U23079 (N_23079,N_22887,N_22733);
nand U23080 (N_23080,N_22891,N_22868);
nand U23081 (N_23081,N_22531,N_22877);
xor U23082 (N_23082,N_22739,N_22993);
or U23083 (N_23083,N_22840,N_22865);
xnor U23084 (N_23084,N_22910,N_22894);
nand U23085 (N_23085,N_22751,N_22780);
or U23086 (N_23086,N_22529,N_22808);
or U23087 (N_23087,N_22982,N_22736);
nand U23088 (N_23088,N_22966,N_22611);
nand U23089 (N_23089,N_22842,N_22687);
and U23090 (N_23090,N_22603,N_22771);
or U23091 (N_23091,N_22927,N_22619);
and U23092 (N_23092,N_22772,N_22548);
and U23093 (N_23093,N_22515,N_22572);
or U23094 (N_23094,N_22590,N_22607);
nand U23095 (N_23095,N_22505,N_22943);
or U23096 (N_23096,N_22651,N_22602);
xnor U23097 (N_23097,N_22832,N_22642);
and U23098 (N_23098,N_22715,N_22601);
or U23099 (N_23099,N_22647,N_22820);
nor U23100 (N_23100,N_22749,N_22968);
nor U23101 (N_23101,N_22803,N_22691);
nor U23102 (N_23102,N_22522,N_22637);
nor U23103 (N_23103,N_22689,N_22574);
nand U23104 (N_23104,N_22980,N_22709);
or U23105 (N_23105,N_22580,N_22797);
and U23106 (N_23106,N_22566,N_22846);
xnor U23107 (N_23107,N_22893,N_22557);
and U23108 (N_23108,N_22738,N_22783);
nand U23109 (N_23109,N_22969,N_22782);
and U23110 (N_23110,N_22702,N_22774);
or U23111 (N_23111,N_22503,N_22518);
nand U23112 (N_23112,N_22930,N_22986);
xnor U23113 (N_23113,N_22816,N_22554);
nor U23114 (N_23114,N_22781,N_22633);
xor U23115 (N_23115,N_22722,N_22799);
nand U23116 (N_23116,N_22564,N_22604);
nand U23117 (N_23117,N_22712,N_22727);
nor U23118 (N_23118,N_22917,N_22562);
or U23119 (N_23119,N_22635,N_22866);
and U23120 (N_23120,N_22682,N_22951);
nor U23121 (N_23121,N_22646,N_22831);
or U23122 (N_23122,N_22654,N_22942);
nor U23123 (N_23123,N_22909,N_22613);
or U23124 (N_23124,N_22999,N_22593);
nand U23125 (N_23125,N_22552,N_22507);
and U23126 (N_23126,N_22599,N_22903);
or U23127 (N_23127,N_22825,N_22681);
and U23128 (N_23128,N_22711,N_22932);
or U23129 (N_23129,N_22561,N_22545);
nor U23130 (N_23130,N_22961,N_22888);
nor U23131 (N_23131,N_22854,N_22540);
or U23132 (N_23132,N_22860,N_22937);
nor U23133 (N_23133,N_22664,N_22676);
xor U23134 (N_23134,N_22991,N_22847);
and U23135 (N_23135,N_22838,N_22923);
nand U23136 (N_23136,N_22901,N_22775);
or U23137 (N_23137,N_22506,N_22537);
and U23138 (N_23138,N_22965,N_22559);
or U23139 (N_23139,N_22536,N_22964);
or U23140 (N_23140,N_22617,N_22952);
or U23141 (N_23141,N_22627,N_22632);
and U23142 (N_23142,N_22864,N_22742);
and U23143 (N_23143,N_22912,N_22971);
nand U23144 (N_23144,N_22929,N_22824);
and U23145 (N_23145,N_22743,N_22765);
nand U23146 (N_23146,N_22779,N_22726);
nor U23147 (N_23147,N_22998,N_22787);
and U23148 (N_23148,N_22631,N_22588);
xnor U23149 (N_23149,N_22662,N_22553);
and U23150 (N_23150,N_22928,N_22660);
or U23151 (N_23151,N_22922,N_22644);
or U23152 (N_23152,N_22849,N_22979);
nand U23153 (N_23153,N_22834,N_22527);
xor U23154 (N_23154,N_22555,N_22586);
nor U23155 (N_23155,N_22665,N_22869);
and U23156 (N_23156,N_22663,N_22757);
or U23157 (N_23157,N_22814,N_22828);
nand U23158 (N_23158,N_22683,N_22533);
and U23159 (N_23159,N_22755,N_22977);
xnor U23160 (N_23160,N_22913,N_22595);
nand U23161 (N_23161,N_22798,N_22666);
and U23162 (N_23162,N_22589,N_22622);
nor U23163 (N_23163,N_22806,N_22573);
and U23164 (N_23164,N_22512,N_22924);
nor U23165 (N_23165,N_22746,N_22669);
or U23166 (N_23166,N_22936,N_22549);
xnor U23167 (N_23167,N_22955,N_22587);
nor U23168 (N_23168,N_22759,N_22975);
nor U23169 (N_23169,N_22648,N_22994);
and U23170 (N_23170,N_22836,N_22921);
nand U23171 (N_23171,N_22653,N_22763);
nor U23172 (N_23172,N_22881,N_22670);
xnor U23173 (N_23173,N_22524,N_22896);
nor U23174 (N_23174,N_22705,N_22629);
nor U23175 (N_23175,N_22584,N_22810);
and U23176 (N_23176,N_22760,N_22915);
nor U23177 (N_23177,N_22567,N_22995);
and U23178 (N_23178,N_22597,N_22920);
or U23179 (N_23179,N_22773,N_22800);
nand U23180 (N_23180,N_22934,N_22508);
or U23181 (N_23181,N_22585,N_22857);
nor U23182 (N_23182,N_22684,N_22858);
xnor U23183 (N_23183,N_22575,N_22862);
xor U23184 (N_23184,N_22766,N_22526);
nand U23185 (N_23185,N_22628,N_22941);
nor U23186 (N_23186,N_22835,N_22621);
nor U23187 (N_23187,N_22976,N_22720);
xor U23188 (N_23188,N_22997,N_22546);
nand U23189 (N_23189,N_22911,N_22610);
nor U23190 (N_23190,N_22753,N_22890);
or U23191 (N_23191,N_22880,N_22815);
nor U23192 (N_23192,N_22657,N_22735);
nor U23193 (N_23193,N_22807,N_22871);
and U23194 (N_23194,N_22926,N_22667);
xnor U23195 (N_23195,N_22616,N_22678);
and U23196 (N_23196,N_22721,N_22931);
xnor U23197 (N_23197,N_22528,N_22914);
and U23198 (N_23198,N_22957,N_22550);
nand U23199 (N_23199,N_22672,N_22532);
and U23200 (N_23200,N_22843,N_22713);
nor U23201 (N_23201,N_22582,N_22697);
nand U23202 (N_23202,N_22543,N_22978);
or U23203 (N_23203,N_22954,N_22804);
nand U23204 (N_23204,N_22708,N_22523);
nand U23205 (N_23205,N_22600,N_22645);
and U23206 (N_23206,N_22822,N_22801);
or U23207 (N_23207,N_22821,N_22946);
or U23208 (N_23208,N_22841,N_22972);
nand U23209 (N_23209,N_22945,N_22714);
nor U23210 (N_23210,N_22542,N_22710);
nor U23211 (N_23211,N_22900,N_22827);
xnor U23212 (N_23212,N_22973,N_22870);
and U23213 (N_23213,N_22852,N_22872);
or U23214 (N_23214,N_22615,N_22990);
and U23215 (N_23215,N_22563,N_22704);
xnor U23216 (N_23216,N_22959,N_22906);
xnor U23217 (N_23217,N_22734,N_22918);
or U23218 (N_23218,N_22596,N_22811);
and U23219 (N_23219,N_22789,N_22638);
nand U23220 (N_23220,N_22577,N_22874);
xor U23221 (N_23221,N_22730,N_22883);
nor U23222 (N_23222,N_22908,N_22855);
xor U23223 (N_23223,N_22754,N_22501);
and U23224 (N_23224,N_22956,N_22511);
nand U23225 (N_23225,N_22984,N_22859);
xor U23226 (N_23226,N_22583,N_22823);
or U23227 (N_23227,N_22876,N_22750);
nor U23228 (N_23228,N_22933,N_22639);
or U23229 (N_23229,N_22571,N_22731);
nand U23230 (N_23230,N_22748,N_22690);
or U23231 (N_23231,N_22895,N_22598);
and U23232 (N_23232,N_22812,N_22916);
xor U23233 (N_23233,N_22695,N_22905);
nand U23234 (N_23234,N_22706,N_22658);
xor U23235 (N_23235,N_22767,N_22679);
nand U23236 (N_23236,N_22745,N_22786);
nand U23237 (N_23237,N_22967,N_22630);
nor U23238 (N_23238,N_22703,N_22845);
nand U23239 (N_23239,N_22699,N_22519);
and U23240 (N_23240,N_22510,N_22640);
or U23241 (N_23241,N_22856,N_22848);
or U23242 (N_23242,N_22833,N_22796);
or U23243 (N_23243,N_22620,N_22762);
xor U23244 (N_23244,N_22641,N_22761);
nor U23245 (N_23245,N_22983,N_22623);
nor U23246 (N_23246,N_22878,N_22578);
nand U23247 (N_23247,N_22686,N_22813);
nand U23248 (N_23248,N_22626,N_22830);
and U23249 (N_23249,N_22940,N_22701);
or U23250 (N_23250,N_22673,N_22769);
and U23251 (N_23251,N_22959,N_22735);
xnor U23252 (N_23252,N_22908,N_22906);
xor U23253 (N_23253,N_22918,N_22989);
or U23254 (N_23254,N_22681,N_22742);
nor U23255 (N_23255,N_22763,N_22739);
and U23256 (N_23256,N_22617,N_22714);
and U23257 (N_23257,N_22992,N_22752);
nand U23258 (N_23258,N_22683,N_22862);
or U23259 (N_23259,N_22990,N_22739);
xnor U23260 (N_23260,N_22905,N_22884);
or U23261 (N_23261,N_22928,N_22664);
nand U23262 (N_23262,N_22692,N_22548);
and U23263 (N_23263,N_22994,N_22752);
nand U23264 (N_23264,N_22734,N_22889);
and U23265 (N_23265,N_22864,N_22668);
nand U23266 (N_23266,N_22646,N_22668);
or U23267 (N_23267,N_22849,N_22611);
and U23268 (N_23268,N_22598,N_22646);
nand U23269 (N_23269,N_22511,N_22938);
or U23270 (N_23270,N_22717,N_22889);
xor U23271 (N_23271,N_22642,N_22901);
or U23272 (N_23272,N_22649,N_22623);
and U23273 (N_23273,N_22817,N_22652);
xor U23274 (N_23274,N_22983,N_22700);
nand U23275 (N_23275,N_22716,N_22725);
or U23276 (N_23276,N_22769,N_22589);
xor U23277 (N_23277,N_22993,N_22810);
xor U23278 (N_23278,N_22960,N_22503);
xor U23279 (N_23279,N_22749,N_22591);
or U23280 (N_23280,N_22739,N_22721);
and U23281 (N_23281,N_22717,N_22550);
and U23282 (N_23282,N_22890,N_22766);
and U23283 (N_23283,N_22807,N_22586);
nor U23284 (N_23284,N_22672,N_22529);
xor U23285 (N_23285,N_22702,N_22575);
nand U23286 (N_23286,N_22906,N_22533);
and U23287 (N_23287,N_22614,N_22869);
or U23288 (N_23288,N_22876,N_22868);
and U23289 (N_23289,N_22837,N_22556);
and U23290 (N_23290,N_22563,N_22744);
nand U23291 (N_23291,N_22909,N_22771);
nand U23292 (N_23292,N_22690,N_22913);
nor U23293 (N_23293,N_22787,N_22534);
or U23294 (N_23294,N_22839,N_22942);
xor U23295 (N_23295,N_22721,N_22980);
or U23296 (N_23296,N_22569,N_22864);
nor U23297 (N_23297,N_22760,N_22693);
nor U23298 (N_23298,N_22997,N_22725);
and U23299 (N_23299,N_22792,N_22899);
and U23300 (N_23300,N_22740,N_22624);
nor U23301 (N_23301,N_22510,N_22983);
and U23302 (N_23302,N_22693,N_22997);
and U23303 (N_23303,N_22971,N_22586);
and U23304 (N_23304,N_22824,N_22700);
and U23305 (N_23305,N_22687,N_22684);
and U23306 (N_23306,N_22876,N_22849);
or U23307 (N_23307,N_22703,N_22509);
nor U23308 (N_23308,N_22569,N_22887);
nand U23309 (N_23309,N_22520,N_22721);
xnor U23310 (N_23310,N_22701,N_22626);
nand U23311 (N_23311,N_22712,N_22859);
nor U23312 (N_23312,N_22975,N_22851);
and U23313 (N_23313,N_22678,N_22727);
or U23314 (N_23314,N_22548,N_22507);
nand U23315 (N_23315,N_22767,N_22964);
or U23316 (N_23316,N_22736,N_22879);
nand U23317 (N_23317,N_22715,N_22787);
nand U23318 (N_23318,N_22835,N_22921);
xor U23319 (N_23319,N_22612,N_22786);
nor U23320 (N_23320,N_22725,N_22897);
and U23321 (N_23321,N_22972,N_22653);
and U23322 (N_23322,N_22697,N_22746);
nand U23323 (N_23323,N_22753,N_22692);
or U23324 (N_23324,N_22797,N_22519);
and U23325 (N_23325,N_22555,N_22734);
nand U23326 (N_23326,N_22625,N_22615);
and U23327 (N_23327,N_22554,N_22754);
nand U23328 (N_23328,N_22851,N_22649);
nor U23329 (N_23329,N_22672,N_22633);
nand U23330 (N_23330,N_22522,N_22539);
xnor U23331 (N_23331,N_22557,N_22742);
xor U23332 (N_23332,N_22685,N_22843);
nand U23333 (N_23333,N_22607,N_22610);
nand U23334 (N_23334,N_22703,N_22856);
xnor U23335 (N_23335,N_22958,N_22649);
nand U23336 (N_23336,N_22513,N_22895);
nand U23337 (N_23337,N_22658,N_22828);
or U23338 (N_23338,N_22662,N_22780);
nor U23339 (N_23339,N_22839,N_22720);
xor U23340 (N_23340,N_22775,N_22733);
xor U23341 (N_23341,N_22519,N_22546);
or U23342 (N_23342,N_22849,N_22540);
nor U23343 (N_23343,N_22574,N_22873);
xor U23344 (N_23344,N_22682,N_22520);
nand U23345 (N_23345,N_22681,N_22650);
xor U23346 (N_23346,N_22961,N_22924);
and U23347 (N_23347,N_22918,N_22611);
nor U23348 (N_23348,N_22922,N_22955);
xnor U23349 (N_23349,N_22552,N_22630);
nor U23350 (N_23350,N_22948,N_22781);
and U23351 (N_23351,N_22841,N_22858);
xor U23352 (N_23352,N_22774,N_22693);
and U23353 (N_23353,N_22697,N_22929);
or U23354 (N_23354,N_22757,N_22631);
or U23355 (N_23355,N_22908,N_22876);
or U23356 (N_23356,N_22605,N_22793);
xor U23357 (N_23357,N_22693,N_22894);
and U23358 (N_23358,N_22646,N_22733);
xnor U23359 (N_23359,N_22982,N_22636);
and U23360 (N_23360,N_22525,N_22708);
nor U23361 (N_23361,N_22646,N_22731);
nand U23362 (N_23362,N_22859,N_22674);
xor U23363 (N_23363,N_22687,N_22771);
and U23364 (N_23364,N_22832,N_22638);
nand U23365 (N_23365,N_22538,N_22859);
nand U23366 (N_23366,N_22867,N_22915);
and U23367 (N_23367,N_22624,N_22597);
and U23368 (N_23368,N_22677,N_22591);
nand U23369 (N_23369,N_22533,N_22531);
xor U23370 (N_23370,N_22803,N_22823);
nand U23371 (N_23371,N_22898,N_22664);
and U23372 (N_23372,N_22740,N_22731);
nor U23373 (N_23373,N_22875,N_22784);
and U23374 (N_23374,N_22864,N_22796);
xnor U23375 (N_23375,N_22978,N_22692);
xnor U23376 (N_23376,N_22603,N_22720);
nor U23377 (N_23377,N_22708,N_22500);
nand U23378 (N_23378,N_22873,N_22509);
xor U23379 (N_23379,N_22957,N_22552);
or U23380 (N_23380,N_22709,N_22975);
nand U23381 (N_23381,N_22745,N_22890);
nand U23382 (N_23382,N_22668,N_22755);
nand U23383 (N_23383,N_22698,N_22944);
nand U23384 (N_23384,N_22597,N_22751);
nand U23385 (N_23385,N_22651,N_22637);
nand U23386 (N_23386,N_22577,N_22674);
nand U23387 (N_23387,N_22850,N_22595);
xor U23388 (N_23388,N_22685,N_22551);
nor U23389 (N_23389,N_22853,N_22996);
or U23390 (N_23390,N_22658,N_22588);
and U23391 (N_23391,N_22918,N_22629);
nor U23392 (N_23392,N_22917,N_22982);
xor U23393 (N_23393,N_22922,N_22536);
and U23394 (N_23394,N_22684,N_22500);
xor U23395 (N_23395,N_22806,N_22708);
nor U23396 (N_23396,N_22521,N_22863);
nor U23397 (N_23397,N_22899,N_22814);
nor U23398 (N_23398,N_22889,N_22748);
xnor U23399 (N_23399,N_22743,N_22689);
nor U23400 (N_23400,N_22688,N_22817);
nand U23401 (N_23401,N_22711,N_22716);
nor U23402 (N_23402,N_22958,N_22756);
and U23403 (N_23403,N_22789,N_22709);
nor U23404 (N_23404,N_22908,N_22810);
or U23405 (N_23405,N_22890,N_22863);
nand U23406 (N_23406,N_22724,N_22670);
or U23407 (N_23407,N_22679,N_22624);
and U23408 (N_23408,N_22553,N_22867);
nor U23409 (N_23409,N_22674,N_22701);
nand U23410 (N_23410,N_22844,N_22590);
nor U23411 (N_23411,N_22713,N_22658);
nand U23412 (N_23412,N_22921,N_22656);
and U23413 (N_23413,N_22597,N_22518);
or U23414 (N_23414,N_22943,N_22677);
nor U23415 (N_23415,N_22895,N_22625);
nor U23416 (N_23416,N_22542,N_22795);
nand U23417 (N_23417,N_22626,N_22506);
xnor U23418 (N_23418,N_22997,N_22958);
or U23419 (N_23419,N_22692,N_22524);
or U23420 (N_23420,N_22505,N_22688);
nor U23421 (N_23421,N_22632,N_22654);
nor U23422 (N_23422,N_22935,N_22672);
nand U23423 (N_23423,N_22619,N_22959);
nand U23424 (N_23424,N_22872,N_22580);
or U23425 (N_23425,N_22667,N_22863);
or U23426 (N_23426,N_22518,N_22627);
and U23427 (N_23427,N_22642,N_22772);
and U23428 (N_23428,N_22831,N_22847);
xnor U23429 (N_23429,N_22985,N_22785);
nand U23430 (N_23430,N_22536,N_22739);
and U23431 (N_23431,N_22965,N_22569);
or U23432 (N_23432,N_22747,N_22743);
nand U23433 (N_23433,N_22638,N_22767);
xnor U23434 (N_23434,N_22781,N_22520);
nor U23435 (N_23435,N_22809,N_22662);
nor U23436 (N_23436,N_22707,N_22726);
nor U23437 (N_23437,N_22866,N_22831);
xnor U23438 (N_23438,N_22694,N_22758);
xor U23439 (N_23439,N_22738,N_22786);
xor U23440 (N_23440,N_22999,N_22718);
nor U23441 (N_23441,N_22916,N_22865);
and U23442 (N_23442,N_22889,N_22875);
xor U23443 (N_23443,N_22763,N_22671);
xor U23444 (N_23444,N_22511,N_22598);
nor U23445 (N_23445,N_22520,N_22740);
nand U23446 (N_23446,N_22606,N_22610);
xnor U23447 (N_23447,N_22855,N_22617);
and U23448 (N_23448,N_22862,N_22533);
nand U23449 (N_23449,N_22890,N_22664);
nor U23450 (N_23450,N_22550,N_22642);
xor U23451 (N_23451,N_22589,N_22571);
or U23452 (N_23452,N_22556,N_22500);
xor U23453 (N_23453,N_22638,N_22596);
nor U23454 (N_23454,N_22518,N_22573);
or U23455 (N_23455,N_22757,N_22929);
or U23456 (N_23456,N_22633,N_22525);
nand U23457 (N_23457,N_22794,N_22975);
xor U23458 (N_23458,N_22636,N_22934);
and U23459 (N_23459,N_22739,N_22521);
nor U23460 (N_23460,N_22954,N_22763);
nor U23461 (N_23461,N_22543,N_22685);
and U23462 (N_23462,N_22877,N_22850);
or U23463 (N_23463,N_22772,N_22530);
nor U23464 (N_23464,N_22585,N_22988);
xor U23465 (N_23465,N_22510,N_22689);
xnor U23466 (N_23466,N_22525,N_22616);
and U23467 (N_23467,N_22523,N_22992);
nand U23468 (N_23468,N_22505,N_22729);
or U23469 (N_23469,N_22867,N_22588);
nand U23470 (N_23470,N_22504,N_22567);
nand U23471 (N_23471,N_22839,N_22902);
nor U23472 (N_23472,N_22980,N_22893);
xnor U23473 (N_23473,N_22931,N_22865);
nand U23474 (N_23474,N_22711,N_22886);
and U23475 (N_23475,N_22895,N_22572);
nand U23476 (N_23476,N_22912,N_22655);
nor U23477 (N_23477,N_22808,N_22539);
or U23478 (N_23478,N_22687,N_22948);
xor U23479 (N_23479,N_22795,N_22987);
or U23480 (N_23480,N_22677,N_22701);
or U23481 (N_23481,N_22521,N_22776);
xnor U23482 (N_23482,N_22935,N_22514);
nor U23483 (N_23483,N_22652,N_22857);
nand U23484 (N_23484,N_22798,N_22552);
nand U23485 (N_23485,N_22945,N_22502);
or U23486 (N_23486,N_22924,N_22901);
or U23487 (N_23487,N_22600,N_22602);
and U23488 (N_23488,N_22894,N_22592);
xnor U23489 (N_23489,N_22818,N_22791);
and U23490 (N_23490,N_22697,N_22728);
and U23491 (N_23491,N_22747,N_22703);
nand U23492 (N_23492,N_22875,N_22966);
and U23493 (N_23493,N_22556,N_22779);
xor U23494 (N_23494,N_22767,N_22942);
xor U23495 (N_23495,N_22642,N_22630);
and U23496 (N_23496,N_22725,N_22599);
and U23497 (N_23497,N_22996,N_22877);
and U23498 (N_23498,N_22720,N_22608);
nor U23499 (N_23499,N_22570,N_22671);
xnor U23500 (N_23500,N_23231,N_23371);
and U23501 (N_23501,N_23490,N_23002);
and U23502 (N_23502,N_23187,N_23051);
xor U23503 (N_23503,N_23112,N_23462);
xor U23504 (N_23504,N_23076,N_23131);
nor U23505 (N_23505,N_23249,N_23115);
nand U23506 (N_23506,N_23319,N_23070);
and U23507 (N_23507,N_23376,N_23454);
xor U23508 (N_23508,N_23016,N_23413);
nor U23509 (N_23509,N_23019,N_23204);
and U23510 (N_23510,N_23009,N_23244);
nor U23511 (N_23511,N_23176,N_23006);
or U23512 (N_23512,N_23260,N_23390);
or U23513 (N_23513,N_23498,N_23086);
xnor U23514 (N_23514,N_23180,N_23338);
xnor U23515 (N_23515,N_23046,N_23395);
nand U23516 (N_23516,N_23442,N_23389);
or U23517 (N_23517,N_23211,N_23484);
nor U23518 (N_23518,N_23132,N_23092);
nand U23519 (N_23519,N_23050,N_23052);
and U23520 (N_23520,N_23323,N_23202);
xnor U23521 (N_23521,N_23315,N_23440);
nand U23522 (N_23522,N_23172,N_23197);
and U23523 (N_23523,N_23380,N_23373);
nor U23524 (N_23524,N_23142,N_23174);
and U23525 (N_23525,N_23021,N_23436);
nand U23526 (N_23526,N_23038,N_23302);
nand U23527 (N_23527,N_23121,N_23457);
nand U23528 (N_23528,N_23403,N_23234);
xnor U23529 (N_23529,N_23129,N_23477);
and U23530 (N_23530,N_23497,N_23333);
and U23531 (N_23531,N_23209,N_23488);
or U23532 (N_23532,N_23257,N_23351);
nor U23533 (N_23533,N_23037,N_23201);
or U23534 (N_23534,N_23081,N_23492);
or U23535 (N_23535,N_23274,N_23054);
nand U23536 (N_23536,N_23219,N_23267);
nor U23537 (N_23537,N_23200,N_23481);
or U23538 (N_23538,N_23342,N_23383);
and U23539 (N_23539,N_23293,N_23294);
nand U23540 (N_23540,N_23183,N_23478);
nor U23541 (N_23541,N_23339,N_23365);
xnor U23542 (N_23542,N_23499,N_23025);
and U23543 (N_23543,N_23203,N_23101);
and U23544 (N_23544,N_23443,N_23362);
nor U23545 (N_23545,N_23446,N_23322);
nand U23546 (N_23546,N_23448,N_23287);
nor U23547 (N_23547,N_23066,N_23136);
xor U23548 (N_23548,N_23221,N_23075);
nand U23549 (N_23549,N_23347,N_23105);
nand U23550 (N_23550,N_23449,N_23149);
and U23551 (N_23551,N_23047,N_23337);
and U23552 (N_23552,N_23042,N_23189);
or U23553 (N_23553,N_23188,N_23169);
or U23554 (N_23554,N_23185,N_23003);
or U23555 (N_23555,N_23384,N_23001);
nor U23556 (N_23556,N_23158,N_23368);
nand U23557 (N_23557,N_23343,N_23332);
xnor U23558 (N_23558,N_23396,N_23346);
and U23559 (N_23559,N_23262,N_23080);
or U23560 (N_23560,N_23327,N_23077);
or U23561 (N_23561,N_23243,N_23217);
xor U23562 (N_23562,N_23400,N_23370);
nor U23563 (N_23563,N_23083,N_23104);
or U23564 (N_23564,N_23401,N_23297);
xnor U23565 (N_23565,N_23279,N_23458);
xnor U23566 (N_23566,N_23198,N_23005);
and U23567 (N_23567,N_23320,N_23334);
nand U23568 (N_23568,N_23124,N_23206);
and U23569 (N_23569,N_23225,N_23407);
xnor U23570 (N_23570,N_23164,N_23166);
nor U23571 (N_23571,N_23270,N_23043);
xnor U23572 (N_23572,N_23034,N_23224);
and U23573 (N_23573,N_23415,N_23153);
nor U23574 (N_23574,N_23157,N_23261);
xor U23575 (N_23575,N_23007,N_23471);
or U23576 (N_23576,N_23387,N_23058);
and U23577 (N_23577,N_23015,N_23226);
xor U23578 (N_23578,N_23160,N_23152);
xnor U23579 (N_23579,N_23283,N_23139);
and U23580 (N_23580,N_23045,N_23162);
xnor U23581 (N_23581,N_23168,N_23299);
nand U23582 (N_23582,N_23069,N_23309);
xnor U23583 (N_23583,N_23156,N_23133);
xnor U23584 (N_23584,N_23286,N_23358);
xor U23585 (N_23585,N_23350,N_23451);
and U23586 (N_23586,N_23100,N_23398);
or U23587 (N_23587,N_23487,N_23290);
or U23588 (N_23588,N_23316,N_23385);
nand U23589 (N_23589,N_23035,N_23321);
or U23590 (N_23590,N_23479,N_23404);
nor U23591 (N_23591,N_23084,N_23428);
xnor U23592 (N_23592,N_23335,N_23344);
and U23593 (N_23593,N_23113,N_23412);
nor U23594 (N_23594,N_23165,N_23378);
xor U23595 (N_23595,N_23119,N_23030);
nor U23596 (N_23596,N_23282,N_23108);
or U23597 (N_23597,N_23087,N_23388);
nand U23598 (N_23598,N_23356,N_23414);
xor U23599 (N_23599,N_23145,N_23265);
nor U23600 (N_23600,N_23360,N_23489);
and U23601 (N_23601,N_23311,N_23191);
xor U23602 (N_23602,N_23452,N_23425);
nand U23603 (N_23603,N_23272,N_23483);
xor U23604 (N_23604,N_23098,N_23430);
and U23605 (N_23605,N_23336,N_23151);
xnor U23606 (N_23606,N_23465,N_23461);
nor U23607 (N_23607,N_23127,N_23285);
nor U23608 (N_23608,N_23125,N_23017);
xnor U23609 (N_23609,N_23361,N_23111);
nor U23610 (N_23610,N_23110,N_23024);
and U23611 (N_23611,N_23314,N_23482);
xor U23612 (N_23612,N_23486,N_23055);
nand U23613 (N_23613,N_23093,N_23245);
and U23614 (N_23614,N_23215,N_23229);
nor U23615 (N_23615,N_23148,N_23057);
nand U23616 (N_23616,N_23013,N_23190);
or U23617 (N_23617,N_23372,N_23405);
nand U23618 (N_23618,N_23235,N_23438);
and U23619 (N_23619,N_23252,N_23000);
xor U23620 (N_23620,N_23277,N_23167);
nand U23621 (N_23621,N_23175,N_23212);
xnor U23622 (N_23622,N_23223,N_23422);
or U23623 (N_23623,N_23273,N_23429);
and U23624 (N_23624,N_23391,N_23324);
xnor U23625 (N_23625,N_23366,N_23144);
and U23626 (N_23626,N_23004,N_23227);
or U23627 (N_23627,N_23241,N_23210);
and U23628 (N_23628,N_23220,N_23154);
or U23629 (N_23629,N_23085,N_23467);
nor U23630 (N_23630,N_23424,N_23163);
xor U23631 (N_23631,N_23445,N_23134);
or U23632 (N_23632,N_23040,N_23096);
or U23633 (N_23633,N_23288,N_23074);
and U23634 (N_23634,N_23061,N_23318);
or U23635 (N_23635,N_23417,N_23248);
nand U23636 (N_23636,N_23247,N_23056);
xor U23637 (N_23637,N_23363,N_23008);
xor U23638 (N_23638,N_23147,N_23341);
nor U23639 (N_23639,N_23353,N_23123);
or U23640 (N_23640,N_23300,N_23444);
and U23641 (N_23641,N_23018,N_23073);
or U23642 (N_23642,N_23072,N_23060);
or U23643 (N_23643,N_23264,N_23313);
or U23644 (N_23644,N_23330,N_23431);
nand U23645 (N_23645,N_23161,N_23146);
nor U23646 (N_23646,N_23205,N_23381);
and U23647 (N_23647,N_23310,N_23182);
nand U23648 (N_23648,N_23214,N_23357);
nor U23649 (N_23649,N_23109,N_23095);
or U23650 (N_23650,N_23033,N_23432);
and U23651 (N_23651,N_23354,N_23469);
or U23652 (N_23652,N_23349,N_23485);
or U23653 (N_23653,N_23059,N_23393);
nor U23654 (N_23654,N_23213,N_23026);
nand U23655 (N_23655,N_23091,N_23420);
xnor U23656 (N_23656,N_23044,N_23359);
xor U23657 (N_23657,N_23032,N_23433);
or U23658 (N_23658,N_23418,N_23379);
and U23659 (N_23659,N_23491,N_23240);
xor U23660 (N_23660,N_23194,N_23230);
xor U23661 (N_23661,N_23308,N_23450);
and U23662 (N_23662,N_23088,N_23196);
xor U23663 (N_23663,N_23281,N_23078);
nor U23664 (N_23664,N_23495,N_23049);
xnor U23665 (N_23665,N_23325,N_23476);
or U23666 (N_23666,N_23114,N_23307);
or U23667 (N_23667,N_23468,N_23392);
nand U23668 (N_23668,N_23090,N_23303);
or U23669 (N_23669,N_23423,N_23171);
or U23670 (N_23670,N_23312,N_23455);
nand U23671 (N_23671,N_23181,N_23118);
and U23672 (N_23672,N_23386,N_23374);
and U23673 (N_23673,N_23014,N_23453);
or U23674 (N_23674,N_23269,N_23222);
or U23675 (N_23675,N_23268,N_23063);
nor U23676 (N_23676,N_23291,N_23238);
nor U23677 (N_23677,N_23232,N_23102);
or U23678 (N_23678,N_23402,N_23177);
or U23679 (N_23679,N_23421,N_23150);
nand U23680 (N_23680,N_23218,N_23305);
nor U23681 (N_23681,N_23475,N_23246);
and U23682 (N_23682,N_23460,N_23493);
or U23683 (N_23683,N_23186,N_23159);
nor U23684 (N_23684,N_23094,N_23117);
xor U23685 (N_23685,N_23340,N_23242);
or U23686 (N_23686,N_23250,N_23437);
xnor U23687 (N_23687,N_23011,N_23128);
nor U23688 (N_23688,N_23141,N_23410);
xnor U23689 (N_23689,N_23053,N_23255);
and U23690 (N_23690,N_23082,N_23416);
and U23691 (N_23691,N_23409,N_23474);
nor U23692 (N_23692,N_23280,N_23466);
nand U23693 (N_23693,N_23027,N_23237);
or U23694 (N_23694,N_23375,N_23170);
xor U23695 (N_23695,N_23199,N_23382);
nand U23696 (N_23696,N_23292,N_23048);
and U23697 (N_23697,N_23067,N_23427);
nor U23698 (N_23698,N_23022,N_23184);
and U23699 (N_23699,N_23459,N_23071);
and U23700 (N_23700,N_23331,N_23130);
xnor U23701 (N_23701,N_23369,N_23464);
xnor U23702 (N_23702,N_23065,N_23266);
or U23703 (N_23703,N_23397,N_23472);
or U23704 (N_23704,N_23263,N_23258);
nor U23705 (N_23705,N_23271,N_23289);
or U23706 (N_23706,N_23106,N_23068);
or U23707 (N_23707,N_23023,N_23317);
xor U23708 (N_23708,N_23473,N_23256);
or U23709 (N_23709,N_23195,N_23364);
or U23710 (N_23710,N_23107,N_23434);
xor U23711 (N_23711,N_23296,N_23441);
nor U23712 (N_23712,N_23216,N_23352);
nand U23713 (N_23713,N_23140,N_23377);
xor U23714 (N_23714,N_23251,N_23103);
or U23715 (N_23715,N_23079,N_23239);
xor U23716 (N_23716,N_23099,N_23259);
or U23717 (N_23717,N_23039,N_23298);
xnor U23718 (N_23718,N_23126,N_23178);
nor U23719 (N_23719,N_23143,N_23470);
xnor U23720 (N_23720,N_23276,N_23480);
nor U23721 (N_23721,N_23419,N_23345);
nand U23722 (N_23722,N_23394,N_23031);
xor U23723 (N_23723,N_23120,N_23435);
nand U23724 (N_23724,N_23399,N_23137);
and U23725 (N_23725,N_23041,N_23036);
nand U23726 (N_23726,N_23447,N_23253);
and U23727 (N_23727,N_23411,N_23228);
or U23728 (N_23728,N_23406,N_23275);
nand U23729 (N_23729,N_23028,N_23306);
nand U23730 (N_23730,N_23496,N_23193);
or U23731 (N_23731,N_23207,N_23062);
nand U23732 (N_23732,N_23064,N_23192);
nor U23733 (N_23733,N_23439,N_23329);
and U23734 (N_23734,N_23304,N_23155);
nand U23735 (N_23735,N_23233,N_23355);
nand U23736 (N_23736,N_23122,N_23138);
xnor U23737 (N_23737,N_23284,N_23089);
nor U23738 (N_23738,N_23012,N_23097);
nor U23739 (N_23739,N_23326,N_23236);
or U23740 (N_23740,N_23367,N_23010);
xor U23741 (N_23741,N_23208,N_23295);
and U23742 (N_23742,N_23348,N_23254);
nand U23743 (N_23743,N_23426,N_23328);
xor U23744 (N_23744,N_23173,N_23135);
and U23745 (N_23745,N_23278,N_23179);
and U23746 (N_23746,N_23029,N_23494);
nand U23747 (N_23747,N_23408,N_23301);
nand U23748 (N_23748,N_23020,N_23456);
and U23749 (N_23749,N_23463,N_23116);
xor U23750 (N_23750,N_23010,N_23151);
or U23751 (N_23751,N_23139,N_23192);
or U23752 (N_23752,N_23017,N_23146);
nor U23753 (N_23753,N_23378,N_23044);
nand U23754 (N_23754,N_23413,N_23278);
nand U23755 (N_23755,N_23453,N_23008);
or U23756 (N_23756,N_23228,N_23341);
or U23757 (N_23757,N_23416,N_23181);
xor U23758 (N_23758,N_23443,N_23087);
nand U23759 (N_23759,N_23482,N_23191);
or U23760 (N_23760,N_23406,N_23465);
nand U23761 (N_23761,N_23071,N_23433);
or U23762 (N_23762,N_23263,N_23119);
nand U23763 (N_23763,N_23110,N_23038);
xnor U23764 (N_23764,N_23036,N_23124);
nor U23765 (N_23765,N_23253,N_23449);
nand U23766 (N_23766,N_23410,N_23065);
nand U23767 (N_23767,N_23081,N_23376);
and U23768 (N_23768,N_23484,N_23023);
xor U23769 (N_23769,N_23079,N_23347);
and U23770 (N_23770,N_23485,N_23491);
nor U23771 (N_23771,N_23295,N_23337);
nand U23772 (N_23772,N_23224,N_23016);
nand U23773 (N_23773,N_23092,N_23264);
nor U23774 (N_23774,N_23112,N_23045);
nand U23775 (N_23775,N_23140,N_23295);
and U23776 (N_23776,N_23073,N_23017);
and U23777 (N_23777,N_23404,N_23316);
nand U23778 (N_23778,N_23170,N_23338);
and U23779 (N_23779,N_23148,N_23228);
and U23780 (N_23780,N_23479,N_23407);
nand U23781 (N_23781,N_23422,N_23430);
or U23782 (N_23782,N_23464,N_23007);
or U23783 (N_23783,N_23287,N_23008);
or U23784 (N_23784,N_23291,N_23469);
nand U23785 (N_23785,N_23127,N_23238);
and U23786 (N_23786,N_23052,N_23234);
xor U23787 (N_23787,N_23223,N_23047);
or U23788 (N_23788,N_23193,N_23308);
or U23789 (N_23789,N_23353,N_23142);
or U23790 (N_23790,N_23436,N_23015);
or U23791 (N_23791,N_23373,N_23271);
nand U23792 (N_23792,N_23179,N_23000);
or U23793 (N_23793,N_23048,N_23035);
and U23794 (N_23794,N_23447,N_23116);
xor U23795 (N_23795,N_23167,N_23034);
or U23796 (N_23796,N_23266,N_23238);
nand U23797 (N_23797,N_23109,N_23009);
and U23798 (N_23798,N_23297,N_23276);
or U23799 (N_23799,N_23344,N_23432);
and U23800 (N_23800,N_23332,N_23465);
nand U23801 (N_23801,N_23117,N_23107);
nor U23802 (N_23802,N_23248,N_23436);
or U23803 (N_23803,N_23220,N_23231);
or U23804 (N_23804,N_23402,N_23030);
nand U23805 (N_23805,N_23391,N_23408);
nand U23806 (N_23806,N_23269,N_23492);
nand U23807 (N_23807,N_23495,N_23374);
nand U23808 (N_23808,N_23026,N_23075);
nand U23809 (N_23809,N_23358,N_23162);
and U23810 (N_23810,N_23171,N_23356);
nor U23811 (N_23811,N_23186,N_23060);
nand U23812 (N_23812,N_23331,N_23273);
or U23813 (N_23813,N_23286,N_23257);
nand U23814 (N_23814,N_23460,N_23292);
or U23815 (N_23815,N_23345,N_23153);
xor U23816 (N_23816,N_23385,N_23241);
nor U23817 (N_23817,N_23352,N_23016);
and U23818 (N_23818,N_23100,N_23081);
or U23819 (N_23819,N_23426,N_23372);
and U23820 (N_23820,N_23073,N_23482);
and U23821 (N_23821,N_23488,N_23413);
nor U23822 (N_23822,N_23088,N_23095);
nor U23823 (N_23823,N_23266,N_23189);
nor U23824 (N_23824,N_23108,N_23048);
nand U23825 (N_23825,N_23238,N_23137);
xor U23826 (N_23826,N_23013,N_23299);
nor U23827 (N_23827,N_23121,N_23280);
nor U23828 (N_23828,N_23091,N_23225);
xnor U23829 (N_23829,N_23368,N_23085);
or U23830 (N_23830,N_23213,N_23053);
nand U23831 (N_23831,N_23338,N_23115);
nor U23832 (N_23832,N_23256,N_23260);
and U23833 (N_23833,N_23169,N_23180);
and U23834 (N_23834,N_23170,N_23390);
xnor U23835 (N_23835,N_23322,N_23053);
and U23836 (N_23836,N_23425,N_23033);
xor U23837 (N_23837,N_23490,N_23346);
or U23838 (N_23838,N_23119,N_23186);
nor U23839 (N_23839,N_23215,N_23075);
xnor U23840 (N_23840,N_23340,N_23400);
and U23841 (N_23841,N_23203,N_23225);
nor U23842 (N_23842,N_23133,N_23157);
xnor U23843 (N_23843,N_23260,N_23300);
nand U23844 (N_23844,N_23292,N_23423);
nor U23845 (N_23845,N_23493,N_23051);
or U23846 (N_23846,N_23112,N_23025);
nor U23847 (N_23847,N_23014,N_23170);
or U23848 (N_23848,N_23254,N_23303);
and U23849 (N_23849,N_23058,N_23174);
nand U23850 (N_23850,N_23064,N_23437);
and U23851 (N_23851,N_23249,N_23281);
xnor U23852 (N_23852,N_23176,N_23368);
and U23853 (N_23853,N_23172,N_23106);
nand U23854 (N_23854,N_23090,N_23297);
xnor U23855 (N_23855,N_23100,N_23482);
nand U23856 (N_23856,N_23177,N_23147);
and U23857 (N_23857,N_23267,N_23121);
xnor U23858 (N_23858,N_23005,N_23100);
or U23859 (N_23859,N_23484,N_23111);
xnor U23860 (N_23860,N_23358,N_23074);
nor U23861 (N_23861,N_23259,N_23094);
xnor U23862 (N_23862,N_23355,N_23186);
xor U23863 (N_23863,N_23130,N_23464);
xnor U23864 (N_23864,N_23361,N_23025);
nor U23865 (N_23865,N_23360,N_23441);
nand U23866 (N_23866,N_23410,N_23407);
or U23867 (N_23867,N_23460,N_23116);
or U23868 (N_23868,N_23371,N_23388);
nand U23869 (N_23869,N_23009,N_23097);
and U23870 (N_23870,N_23333,N_23406);
xnor U23871 (N_23871,N_23154,N_23278);
and U23872 (N_23872,N_23119,N_23079);
or U23873 (N_23873,N_23494,N_23427);
or U23874 (N_23874,N_23165,N_23478);
nand U23875 (N_23875,N_23177,N_23425);
nor U23876 (N_23876,N_23024,N_23090);
nand U23877 (N_23877,N_23316,N_23374);
or U23878 (N_23878,N_23355,N_23456);
or U23879 (N_23879,N_23356,N_23321);
xor U23880 (N_23880,N_23217,N_23215);
and U23881 (N_23881,N_23332,N_23309);
nor U23882 (N_23882,N_23367,N_23350);
nand U23883 (N_23883,N_23239,N_23033);
or U23884 (N_23884,N_23498,N_23430);
xnor U23885 (N_23885,N_23275,N_23401);
xnor U23886 (N_23886,N_23197,N_23438);
and U23887 (N_23887,N_23186,N_23346);
or U23888 (N_23888,N_23273,N_23470);
nand U23889 (N_23889,N_23025,N_23202);
nand U23890 (N_23890,N_23013,N_23462);
or U23891 (N_23891,N_23181,N_23063);
or U23892 (N_23892,N_23126,N_23115);
and U23893 (N_23893,N_23176,N_23338);
or U23894 (N_23894,N_23266,N_23152);
nor U23895 (N_23895,N_23487,N_23127);
nor U23896 (N_23896,N_23197,N_23287);
and U23897 (N_23897,N_23412,N_23028);
nand U23898 (N_23898,N_23240,N_23164);
nor U23899 (N_23899,N_23380,N_23051);
or U23900 (N_23900,N_23100,N_23383);
nand U23901 (N_23901,N_23368,N_23373);
xor U23902 (N_23902,N_23058,N_23161);
and U23903 (N_23903,N_23438,N_23297);
and U23904 (N_23904,N_23423,N_23278);
xnor U23905 (N_23905,N_23073,N_23229);
and U23906 (N_23906,N_23488,N_23486);
or U23907 (N_23907,N_23171,N_23322);
nor U23908 (N_23908,N_23388,N_23433);
or U23909 (N_23909,N_23027,N_23078);
and U23910 (N_23910,N_23470,N_23036);
or U23911 (N_23911,N_23171,N_23275);
and U23912 (N_23912,N_23126,N_23095);
xor U23913 (N_23913,N_23146,N_23029);
nor U23914 (N_23914,N_23425,N_23181);
xor U23915 (N_23915,N_23046,N_23496);
and U23916 (N_23916,N_23035,N_23339);
or U23917 (N_23917,N_23422,N_23127);
xnor U23918 (N_23918,N_23311,N_23112);
nor U23919 (N_23919,N_23146,N_23065);
nor U23920 (N_23920,N_23186,N_23191);
and U23921 (N_23921,N_23216,N_23293);
nor U23922 (N_23922,N_23005,N_23437);
or U23923 (N_23923,N_23323,N_23024);
or U23924 (N_23924,N_23332,N_23080);
nand U23925 (N_23925,N_23192,N_23244);
or U23926 (N_23926,N_23306,N_23289);
or U23927 (N_23927,N_23118,N_23455);
nand U23928 (N_23928,N_23084,N_23012);
and U23929 (N_23929,N_23387,N_23278);
nor U23930 (N_23930,N_23165,N_23452);
nand U23931 (N_23931,N_23297,N_23096);
xor U23932 (N_23932,N_23260,N_23384);
nor U23933 (N_23933,N_23082,N_23472);
nand U23934 (N_23934,N_23186,N_23298);
nor U23935 (N_23935,N_23097,N_23178);
or U23936 (N_23936,N_23182,N_23059);
nand U23937 (N_23937,N_23129,N_23051);
xnor U23938 (N_23938,N_23195,N_23071);
or U23939 (N_23939,N_23496,N_23014);
and U23940 (N_23940,N_23049,N_23154);
nor U23941 (N_23941,N_23482,N_23304);
nor U23942 (N_23942,N_23073,N_23007);
nand U23943 (N_23943,N_23021,N_23463);
nand U23944 (N_23944,N_23016,N_23466);
or U23945 (N_23945,N_23034,N_23028);
and U23946 (N_23946,N_23278,N_23137);
nand U23947 (N_23947,N_23278,N_23188);
nand U23948 (N_23948,N_23138,N_23405);
or U23949 (N_23949,N_23230,N_23444);
or U23950 (N_23950,N_23254,N_23262);
nor U23951 (N_23951,N_23456,N_23196);
or U23952 (N_23952,N_23144,N_23446);
nor U23953 (N_23953,N_23325,N_23025);
nor U23954 (N_23954,N_23477,N_23206);
or U23955 (N_23955,N_23233,N_23052);
nor U23956 (N_23956,N_23402,N_23043);
xor U23957 (N_23957,N_23144,N_23057);
or U23958 (N_23958,N_23314,N_23338);
or U23959 (N_23959,N_23463,N_23449);
and U23960 (N_23960,N_23352,N_23082);
nor U23961 (N_23961,N_23180,N_23157);
xor U23962 (N_23962,N_23349,N_23005);
nand U23963 (N_23963,N_23013,N_23369);
xor U23964 (N_23964,N_23423,N_23286);
xor U23965 (N_23965,N_23386,N_23450);
xor U23966 (N_23966,N_23112,N_23254);
xnor U23967 (N_23967,N_23165,N_23469);
or U23968 (N_23968,N_23089,N_23367);
or U23969 (N_23969,N_23045,N_23482);
nor U23970 (N_23970,N_23263,N_23247);
and U23971 (N_23971,N_23162,N_23371);
xnor U23972 (N_23972,N_23296,N_23394);
nor U23973 (N_23973,N_23208,N_23212);
and U23974 (N_23974,N_23274,N_23445);
nand U23975 (N_23975,N_23206,N_23398);
nor U23976 (N_23976,N_23278,N_23491);
and U23977 (N_23977,N_23095,N_23481);
xor U23978 (N_23978,N_23430,N_23169);
nor U23979 (N_23979,N_23221,N_23241);
and U23980 (N_23980,N_23402,N_23111);
nand U23981 (N_23981,N_23489,N_23203);
nor U23982 (N_23982,N_23452,N_23336);
nand U23983 (N_23983,N_23187,N_23258);
or U23984 (N_23984,N_23171,N_23042);
nand U23985 (N_23985,N_23104,N_23285);
and U23986 (N_23986,N_23438,N_23206);
nor U23987 (N_23987,N_23107,N_23079);
nor U23988 (N_23988,N_23232,N_23349);
nand U23989 (N_23989,N_23078,N_23394);
nor U23990 (N_23990,N_23245,N_23371);
nand U23991 (N_23991,N_23054,N_23031);
or U23992 (N_23992,N_23244,N_23334);
nor U23993 (N_23993,N_23493,N_23455);
or U23994 (N_23994,N_23051,N_23058);
and U23995 (N_23995,N_23068,N_23203);
and U23996 (N_23996,N_23084,N_23143);
nand U23997 (N_23997,N_23388,N_23448);
xor U23998 (N_23998,N_23217,N_23018);
or U23999 (N_23999,N_23191,N_23201);
xor U24000 (N_24000,N_23780,N_23746);
and U24001 (N_24001,N_23514,N_23911);
nand U24002 (N_24002,N_23633,N_23702);
and U24003 (N_24003,N_23836,N_23752);
nor U24004 (N_24004,N_23813,N_23798);
nor U24005 (N_24005,N_23992,N_23765);
xnor U24006 (N_24006,N_23951,N_23500);
xnor U24007 (N_24007,N_23907,N_23824);
nand U24008 (N_24008,N_23603,N_23677);
nor U24009 (N_24009,N_23811,N_23887);
and U24010 (N_24010,N_23738,N_23876);
nand U24011 (N_24011,N_23627,N_23850);
nor U24012 (N_24012,N_23636,N_23965);
nand U24013 (N_24013,N_23804,N_23851);
and U24014 (N_24014,N_23938,N_23833);
or U24015 (N_24015,N_23655,N_23642);
nor U24016 (N_24016,N_23674,N_23816);
or U24017 (N_24017,N_23787,N_23940);
or U24018 (N_24018,N_23873,N_23966);
xnor U24019 (N_24019,N_23689,N_23552);
nor U24020 (N_24020,N_23797,N_23519);
and U24021 (N_24021,N_23934,N_23631);
nand U24022 (N_24022,N_23678,N_23546);
nor U24023 (N_24023,N_23877,N_23892);
or U24024 (N_24024,N_23923,N_23639);
and U24025 (N_24025,N_23714,N_23721);
and U24026 (N_24026,N_23701,N_23838);
xnor U24027 (N_24027,N_23692,N_23520);
or U24028 (N_24028,N_23530,N_23592);
xor U24029 (N_24029,N_23626,N_23872);
or U24030 (N_24030,N_23572,N_23554);
nor U24031 (N_24031,N_23582,N_23645);
xor U24032 (N_24032,N_23744,N_23676);
or U24033 (N_24033,N_23600,N_23548);
or U24034 (N_24034,N_23586,N_23724);
and U24035 (N_24035,N_23613,N_23567);
xnor U24036 (N_24036,N_23644,N_23761);
nand U24037 (N_24037,N_23789,N_23704);
xor U24038 (N_24038,N_23659,N_23931);
nor U24039 (N_24039,N_23825,N_23763);
nand U24040 (N_24040,N_23890,N_23844);
or U24041 (N_24041,N_23710,N_23932);
xnor U24042 (N_24042,N_23898,N_23771);
xnor U24043 (N_24043,N_23728,N_23709);
and U24044 (N_24044,N_23889,N_23717);
nand U24045 (N_24045,N_23591,N_23802);
nor U24046 (N_24046,N_23720,N_23945);
nand U24047 (N_24047,N_23848,N_23580);
and U24048 (N_24048,N_23909,N_23980);
and U24049 (N_24049,N_23835,N_23616);
nand U24050 (N_24050,N_23896,N_23904);
nand U24051 (N_24051,N_23884,N_23905);
nor U24052 (N_24052,N_23680,N_23528);
nor U24053 (N_24053,N_23840,N_23693);
or U24054 (N_24054,N_23630,N_23681);
xnor U24055 (N_24055,N_23814,N_23682);
nor U24056 (N_24056,N_23533,N_23852);
nor U24057 (N_24057,N_23772,N_23819);
and U24058 (N_24058,N_23602,N_23999);
xnor U24059 (N_24059,N_23732,N_23641);
or U24060 (N_24060,N_23551,N_23820);
or U24061 (N_24061,N_23524,N_23886);
xnor U24062 (N_24062,N_23596,N_23975);
or U24063 (N_24063,N_23985,N_23723);
xnor U24064 (N_24064,N_23961,N_23737);
nand U24065 (N_24065,N_23978,N_23785);
nand U24066 (N_24066,N_23607,N_23529);
and U24067 (N_24067,N_23808,N_23593);
nand U24068 (N_24068,N_23537,N_23543);
xnor U24069 (N_24069,N_23866,N_23990);
xor U24070 (N_24070,N_23536,N_23733);
nor U24071 (N_24071,N_23564,N_23617);
or U24072 (N_24072,N_23656,N_23668);
nand U24073 (N_24073,N_23594,N_23981);
nor U24074 (N_24074,N_23859,N_23688);
nor U24075 (N_24075,N_23807,N_23917);
xnor U24076 (N_24076,N_23699,N_23669);
and U24077 (N_24077,N_23700,N_23918);
nor U24078 (N_24078,N_23865,N_23703);
nand U24079 (N_24079,N_23778,N_23942);
nor U24080 (N_24080,N_23657,N_23916);
nand U24081 (N_24081,N_23638,N_23827);
nand U24082 (N_24082,N_23996,N_23910);
xnor U24083 (N_24083,N_23903,N_23747);
and U24084 (N_24084,N_23513,N_23534);
or U24085 (N_24085,N_23549,N_23691);
and U24086 (N_24086,N_23518,N_23698);
xor U24087 (N_24087,N_23955,N_23768);
xnor U24088 (N_24088,N_23683,N_23870);
nor U24089 (N_24089,N_23989,N_23647);
xor U24090 (N_24090,N_23935,N_23756);
nand U24091 (N_24091,N_23803,N_23745);
or U24092 (N_24092,N_23742,N_23545);
or U24093 (N_24093,N_23949,N_23957);
nor U24094 (N_24094,N_23968,N_23502);
nand U24095 (N_24095,N_23624,N_23925);
or U24096 (N_24096,N_23954,N_23762);
and U24097 (N_24097,N_23984,N_23532);
or U24098 (N_24098,N_23615,N_23544);
nor U24099 (N_24099,N_23598,N_23505);
or U24100 (N_24100,N_23509,N_23861);
nand U24101 (N_24101,N_23900,N_23569);
nor U24102 (N_24102,N_23540,N_23766);
xnor U24103 (N_24103,N_23888,N_23716);
and U24104 (N_24104,N_23760,N_23862);
nor U24105 (N_24105,N_23727,N_23901);
or U24106 (N_24106,N_23610,N_23809);
xnor U24107 (N_24107,N_23921,N_23757);
xor U24108 (N_24108,N_23912,N_23829);
xnor U24109 (N_24109,N_23725,N_23652);
nor U24110 (N_24110,N_23628,N_23775);
xnor U24111 (N_24111,N_23566,N_23667);
or U24112 (N_24112,N_23928,N_23941);
nand U24113 (N_24113,N_23823,N_23770);
xor U24114 (N_24114,N_23690,N_23527);
or U24115 (N_24115,N_23755,N_23882);
xor U24116 (N_24116,N_23958,N_23878);
xor U24117 (N_24117,N_23854,N_23557);
or U24118 (N_24118,N_23895,N_23611);
nor U24119 (N_24119,N_23577,N_23972);
nand U24120 (N_24120,N_23541,N_23649);
nand U24121 (N_24121,N_23663,N_23601);
and U24122 (N_24122,N_23553,N_23517);
nor U24123 (N_24123,N_23585,N_23995);
and U24124 (N_24124,N_23754,N_23860);
nor U24125 (N_24125,N_23960,N_23521);
nand U24126 (N_24126,N_23563,N_23507);
nor U24127 (N_24127,N_23962,N_23672);
or U24128 (N_24128,N_23841,N_23708);
xnor U24129 (N_24129,N_23915,N_23558);
and U24130 (N_24130,N_23913,N_23881);
and U24131 (N_24131,N_23658,N_23832);
or U24132 (N_24132,N_23826,N_23830);
xnor U24133 (N_24133,N_23806,N_23774);
and U24134 (N_24134,N_23885,N_23643);
or U24135 (N_24135,N_23751,N_23654);
and U24136 (N_24136,N_23991,N_23620);
and U24137 (N_24137,N_23842,N_23512);
nand U24138 (N_24138,N_23706,N_23501);
xor U24139 (N_24139,N_23976,N_23711);
and U24140 (N_24140,N_23753,N_23697);
xnor U24141 (N_24141,N_23718,N_23587);
nand U24142 (N_24142,N_23993,N_23758);
and U24143 (N_24143,N_23969,N_23748);
xnor U24144 (N_24144,N_23719,N_23792);
nand U24145 (N_24145,N_23648,N_23695);
nor U24146 (N_24146,N_23660,N_23963);
nor U24147 (N_24147,N_23650,N_23741);
and U24148 (N_24148,N_23555,N_23570);
nor U24149 (N_24149,N_23675,N_23583);
and U24150 (N_24150,N_23967,N_23503);
or U24151 (N_24151,N_23946,N_23982);
or U24152 (N_24152,N_23791,N_23618);
nor U24153 (N_24153,N_23705,N_23696);
or U24154 (N_24154,N_23973,N_23584);
and U24155 (N_24155,N_23902,N_23855);
xnor U24156 (N_24156,N_23767,N_23879);
nor U24157 (N_24157,N_23635,N_23561);
nor U24158 (N_24158,N_23640,N_23599);
or U24159 (N_24159,N_23919,N_23783);
nand U24160 (N_24160,N_23666,N_23974);
xor U24161 (N_24161,N_23799,N_23614);
nor U24162 (N_24162,N_23927,N_23686);
nor U24163 (N_24163,N_23629,N_23531);
nand U24164 (N_24164,N_23578,N_23843);
nor U24165 (N_24165,N_23597,N_23948);
nand U24166 (N_24166,N_23573,N_23589);
nor U24167 (N_24167,N_23562,N_23550);
xor U24168 (N_24168,N_23933,N_23950);
nor U24169 (N_24169,N_23576,N_23936);
and U24170 (N_24170,N_23964,N_23883);
nand U24171 (N_24171,N_23800,N_23522);
and U24172 (N_24172,N_23930,N_23864);
and U24173 (N_24173,N_23665,N_23749);
or U24174 (N_24174,N_23997,N_23715);
xor U24175 (N_24175,N_23952,N_23712);
nor U24176 (N_24176,N_23897,N_23998);
nor U24177 (N_24177,N_23671,N_23515);
nor U24178 (N_24178,N_23739,N_23874);
and U24179 (N_24179,N_23565,N_23773);
nor U24180 (N_24180,N_23612,N_23535);
nor U24181 (N_24181,N_23730,N_23784);
or U24182 (N_24182,N_23834,N_23664);
xor U24183 (N_24183,N_23788,N_23943);
nand U24184 (N_24184,N_23619,N_23653);
or U24185 (N_24185,N_23590,N_23623);
xor U24186 (N_24186,N_23988,N_23504);
nor U24187 (N_24187,N_23894,N_23604);
nor U24188 (N_24188,N_23795,N_23729);
nor U24189 (N_24189,N_23899,N_23547);
xnor U24190 (N_24190,N_23731,N_23922);
or U24191 (N_24191,N_23891,N_23646);
nor U24192 (N_24192,N_23810,N_23818);
and U24193 (N_24193,N_23684,N_23831);
xor U24194 (N_24194,N_23822,N_23559);
nor U24195 (N_24195,N_23722,N_23673);
xor U24196 (N_24196,N_23506,N_23839);
xnor U24197 (N_24197,N_23953,N_23959);
nand U24198 (N_24198,N_23893,N_23574);
nor U24199 (N_24199,N_23581,N_23880);
or U24200 (N_24200,N_23516,N_23670);
nand U24201 (N_24201,N_23979,N_23568);
nor U24202 (N_24202,N_23863,N_23651);
nor U24203 (N_24203,N_23924,N_23853);
nand U24204 (N_24204,N_23736,N_23908);
nand U24205 (N_24205,N_23939,N_23622);
or U24206 (N_24206,N_23777,N_23871);
xor U24207 (N_24207,N_23845,N_23793);
or U24208 (N_24208,N_23595,N_23662);
nor U24209 (N_24209,N_23750,N_23634);
nand U24210 (N_24210,N_23556,N_23508);
or U24211 (N_24211,N_23782,N_23779);
xnor U24212 (N_24212,N_23511,N_23560);
xor U24213 (N_24213,N_23525,N_23867);
xor U24214 (N_24214,N_23812,N_23764);
nor U24215 (N_24215,N_23637,N_23786);
and U24216 (N_24216,N_23796,N_23875);
nor U24217 (N_24217,N_23987,N_23734);
nand U24218 (N_24218,N_23929,N_23735);
and U24219 (N_24219,N_23632,N_23856);
or U24220 (N_24220,N_23971,N_23994);
xnor U24221 (N_24221,N_23986,N_23846);
nand U24222 (N_24222,N_23801,N_23920);
xor U24223 (N_24223,N_23805,N_23970);
nor U24224 (N_24224,N_23837,N_23606);
nand U24225 (N_24225,N_23687,N_23815);
or U24226 (N_24226,N_23937,N_23707);
nor U24227 (N_24227,N_23713,N_23977);
xor U24228 (N_24228,N_23726,N_23743);
nor U24229 (N_24229,N_23588,N_23609);
and U24230 (N_24230,N_23944,N_23776);
and U24231 (N_24231,N_23625,N_23769);
and U24232 (N_24232,N_23821,N_23571);
nor U24233 (N_24233,N_23523,N_23926);
nor U24234 (N_24234,N_23621,N_23956);
nor U24235 (N_24235,N_23817,N_23510);
nand U24236 (N_24236,N_23947,N_23857);
and U24237 (N_24237,N_23526,N_23847);
and U24238 (N_24238,N_23759,N_23914);
and U24239 (N_24239,N_23538,N_23608);
xnor U24240 (N_24240,N_23661,N_23794);
or U24241 (N_24241,N_23790,N_23694);
xnor U24242 (N_24242,N_23781,N_23983);
nand U24243 (N_24243,N_23685,N_23679);
nor U24244 (N_24244,N_23858,N_23542);
or U24245 (N_24245,N_23849,N_23605);
and U24246 (N_24246,N_23579,N_23740);
nand U24247 (N_24247,N_23575,N_23868);
nand U24248 (N_24248,N_23869,N_23828);
nand U24249 (N_24249,N_23539,N_23906);
nor U24250 (N_24250,N_23970,N_23629);
nor U24251 (N_24251,N_23777,N_23764);
nand U24252 (N_24252,N_23968,N_23622);
and U24253 (N_24253,N_23807,N_23572);
or U24254 (N_24254,N_23628,N_23882);
xor U24255 (N_24255,N_23741,N_23965);
nor U24256 (N_24256,N_23600,N_23974);
nand U24257 (N_24257,N_23843,N_23678);
or U24258 (N_24258,N_23827,N_23999);
or U24259 (N_24259,N_23967,N_23871);
or U24260 (N_24260,N_23797,N_23664);
nor U24261 (N_24261,N_23514,N_23912);
nor U24262 (N_24262,N_23509,N_23873);
or U24263 (N_24263,N_23589,N_23528);
nor U24264 (N_24264,N_23680,N_23648);
and U24265 (N_24265,N_23504,N_23976);
nand U24266 (N_24266,N_23750,N_23575);
nor U24267 (N_24267,N_23923,N_23666);
or U24268 (N_24268,N_23880,N_23975);
nor U24269 (N_24269,N_23640,N_23789);
nor U24270 (N_24270,N_23623,N_23767);
nor U24271 (N_24271,N_23872,N_23967);
xnor U24272 (N_24272,N_23779,N_23873);
and U24273 (N_24273,N_23862,N_23504);
and U24274 (N_24274,N_23865,N_23560);
nor U24275 (N_24275,N_23621,N_23735);
and U24276 (N_24276,N_23543,N_23627);
nor U24277 (N_24277,N_23660,N_23740);
or U24278 (N_24278,N_23573,N_23982);
nor U24279 (N_24279,N_23947,N_23991);
or U24280 (N_24280,N_23705,N_23544);
xor U24281 (N_24281,N_23744,N_23781);
or U24282 (N_24282,N_23683,N_23785);
nand U24283 (N_24283,N_23972,N_23702);
or U24284 (N_24284,N_23543,N_23914);
nor U24285 (N_24285,N_23542,N_23854);
or U24286 (N_24286,N_23763,N_23691);
nor U24287 (N_24287,N_23532,N_23626);
xnor U24288 (N_24288,N_23923,N_23712);
xnor U24289 (N_24289,N_23578,N_23565);
nor U24290 (N_24290,N_23657,N_23810);
nor U24291 (N_24291,N_23597,N_23510);
or U24292 (N_24292,N_23767,N_23607);
xor U24293 (N_24293,N_23909,N_23579);
xnor U24294 (N_24294,N_23669,N_23936);
and U24295 (N_24295,N_23862,N_23654);
nor U24296 (N_24296,N_23721,N_23669);
xor U24297 (N_24297,N_23524,N_23755);
or U24298 (N_24298,N_23957,N_23818);
and U24299 (N_24299,N_23855,N_23847);
nand U24300 (N_24300,N_23930,N_23602);
nand U24301 (N_24301,N_23619,N_23661);
xor U24302 (N_24302,N_23680,N_23585);
or U24303 (N_24303,N_23845,N_23719);
and U24304 (N_24304,N_23571,N_23650);
and U24305 (N_24305,N_23893,N_23578);
nand U24306 (N_24306,N_23726,N_23855);
nor U24307 (N_24307,N_23735,N_23624);
xor U24308 (N_24308,N_23615,N_23754);
and U24309 (N_24309,N_23897,N_23878);
nand U24310 (N_24310,N_23920,N_23561);
nand U24311 (N_24311,N_23847,N_23867);
nor U24312 (N_24312,N_23864,N_23568);
xor U24313 (N_24313,N_23968,N_23957);
nor U24314 (N_24314,N_23775,N_23642);
nand U24315 (N_24315,N_23923,N_23613);
xor U24316 (N_24316,N_23955,N_23874);
or U24317 (N_24317,N_23780,N_23841);
xor U24318 (N_24318,N_23909,N_23536);
nand U24319 (N_24319,N_23986,N_23527);
nand U24320 (N_24320,N_23567,N_23666);
or U24321 (N_24321,N_23994,N_23591);
xor U24322 (N_24322,N_23520,N_23699);
xnor U24323 (N_24323,N_23764,N_23807);
nor U24324 (N_24324,N_23555,N_23892);
nor U24325 (N_24325,N_23696,N_23910);
nor U24326 (N_24326,N_23591,N_23617);
and U24327 (N_24327,N_23605,N_23629);
and U24328 (N_24328,N_23589,N_23970);
nand U24329 (N_24329,N_23866,N_23977);
xor U24330 (N_24330,N_23687,N_23608);
nand U24331 (N_24331,N_23731,N_23739);
nand U24332 (N_24332,N_23905,N_23679);
xnor U24333 (N_24333,N_23505,N_23818);
and U24334 (N_24334,N_23523,N_23790);
or U24335 (N_24335,N_23681,N_23570);
nor U24336 (N_24336,N_23508,N_23719);
nor U24337 (N_24337,N_23519,N_23711);
nand U24338 (N_24338,N_23875,N_23970);
or U24339 (N_24339,N_23630,N_23533);
nor U24340 (N_24340,N_23987,N_23841);
nand U24341 (N_24341,N_23574,N_23669);
nand U24342 (N_24342,N_23996,N_23693);
or U24343 (N_24343,N_23854,N_23666);
nor U24344 (N_24344,N_23506,N_23526);
xor U24345 (N_24345,N_23532,N_23517);
nor U24346 (N_24346,N_23842,N_23820);
nor U24347 (N_24347,N_23642,N_23508);
nand U24348 (N_24348,N_23756,N_23550);
or U24349 (N_24349,N_23695,N_23908);
nand U24350 (N_24350,N_23705,N_23787);
and U24351 (N_24351,N_23880,N_23731);
nand U24352 (N_24352,N_23839,N_23902);
or U24353 (N_24353,N_23512,N_23612);
or U24354 (N_24354,N_23727,N_23510);
and U24355 (N_24355,N_23745,N_23987);
xnor U24356 (N_24356,N_23779,N_23546);
and U24357 (N_24357,N_23797,N_23918);
xor U24358 (N_24358,N_23668,N_23543);
nand U24359 (N_24359,N_23991,N_23649);
xor U24360 (N_24360,N_23573,N_23832);
nand U24361 (N_24361,N_23790,N_23503);
nand U24362 (N_24362,N_23971,N_23864);
xnor U24363 (N_24363,N_23527,N_23819);
xor U24364 (N_24364,N_23773,N_23809);
or U24365 (N_24365,N_23691,N_23615);
xnor U24366 (N_24366,N_23666,N_23848);
xnor U24367 (N_24367,N_23822,N_23555);
xor U24368 (N_24368,N_23954,N_23971);
and U24369 (N_24369,N_23636,N_23717);
xnor U24370 (N_24370,N_23509,N_23592);
or U24371 (N_24371,N_23933,N_23836);
xnor U24372 (N_24372,N_23502,N_23505);
nor U24373 (N_24373,N_23804,N_23666);
nand U24374 (N_24374,N_23856,N_23879);
nand U24375 (N_24375,N_23851,N_23610);
xnor U24376 (N_24376,N_23820,N_23670);
nor U24377 (N_24377,N_23940,N_23624);
xnor U24378 (N_24378,N_23705,N_23527);
and U24379 (N_24379,N_23730,N_23796);
and U24380 (N_24380,N_23735,N_23700);
and U24381 (N_24381,N_23612,N_23711);
xor U24382 (N_24382,N_23662,N_23739);
or U24383 (N_24383,N_23864,N_23953);
nor U24384 (N_24384,N_23571,N_23674);
or U24385 (N_24385,N_23667,N_23718);
nor U24386 (N_24386,N_23971,N_23851);
xnor U24387 (N_24387,N_23887,N_23844);
nand U24388 (N_24388,N_23707,N_23682);
nor U24389 (N_24389,N_23634,N_23658);
or U24390 (N_24390,N_23972,N_23861);
xor U24391 (N_24391,N_23536,N_23746);
nor U24392 (N_24392,N_23574,N_23611);
nand U24393 (N_24393,N_23812,N_23604);
or U24394 (N_24394,N_23967,N_23615);
xor U24395 (N_24395,N_23713,N_23581);
xor U24396 (N_24396,N_23834,N_23694);
or U24397 (N_24397,N_23875,N_23727);
or U24398 (N_24398,N_23800,N_23869);
nor U24399 (N_24399,N_23971,N_23522);
or U24400 (N_24400,N_23798,N_23852);
nor U24401 (N_24401,N_23723,N_23633);
and U24402 (N_24402,N_23595,N_23917);
nand U24403 (N_24403,N_23561,N_23559);
nor U24404 (N_24404,N_23503,N_23715);
xnor U24405 (N_24405,N_23840,N_23591);
nand U24406 (N_24406,N_23562,N_23675);
nand U24407 (N_24407,N_23549,N_23539);
nand U24408 (N_24408,N_23522,N_23654);
nand U24409 (N_24409,N_23723,N_23539);
nor U24410 (N_24410,N_23698,N_23842);
and U24411 (N_24411,N_23977,N_23614);
and U24412 (N_24412,N_23629,N_23788);
and U24413 (N_24413,N_23846,N_23970);
xnor U24414 (N_24414,N_23784,N_23878);
or U24415 (N_24415,N_23913,N_23770);
nand U24416 (N_24416,N_23730,N_23648);
and U24417 (N_24417,N_23712,N_23750);
nand U24418 (N_24418,N_23665,N_23627);
nand U24419 (N_24419,N_23695,N_23878);
nor U24420 (N_24420,N_23863,N_23894);
xnor U24421 (N_24421,N_23613,N_23625);
and U24422 (N_24422,N_23505,N_23530);
xor U24423 (N_24423,N_23621,N_23680);
nand U24424 (N_24424,N_23575,N_23960);
xor U24425 (N_24425,N_23531,N_23638);
xor U24426 (N_24426,N_23787,N_23569);
nand U24427 (N_24427,N_23762,N_23504);
or U24428 (N_24428,N_23893,N_23714);
or U24429 (N_24429,N_23968,N_23836);
nand U24430 (N_24430,N_23765,N_23924);
nor U24431 (N_24431,N_23507,N_23995);
xnor U24432 (N_24432,N_23719,N_23649);
nor U24433 (N_24433,N_23551,N_23955);
and U24434 (N_24434,N_23660,N_23659);
or U24435 (N_24435,N_23656,N_23607);
nor U24436 (N_24436,N_23822,N_23656);
xnor U24437 (N_24437,N_23650,N_23902);
or U24438 (N_24438,N_23740,N_23500);
nor U24439 (N_24439,N_23535,N_23688);
or U24440 (N_24440,N_23938,N_23790);
xnor U24441 (N_24441,N_23878,N_23886);
and U24442 (N_24442,N_23932,N_23533);
nor U24443 (N_24443,N_23571,N_23942);
nor U24444 (N_24444,N_23880,N_23808);
nor U24445 (N_24445,N_23585,N_23520);
nand U24446 (N_24446,N_23565,N_23792);
or U24447 (N_24447,N_23560,N_23955);
nand U24448 (N_24448,N_23540,N_23921);
xor U24449 (N_24449,N_23630,N_23593);
nor U24450 (N_24450,N_23687,N_23787);
nor U24451 (N_24451,N_23892,N_23601);
nand U24452 (N_24452,N_23982,N_23546);
or U24453 (N_24453,N_23728,N_23577);
nor U24454 (N_24454,N_23608,N_23791);
nand U24455 (N_24455,N_23698,N_23520);
nor U24456 (N_24456,N_23696,N_23687);
nand U24457 (N_24457,N_23785,N_23869);
nor U24458 (N_24458,N_23906,N_23894);
nand U24459 (N_24459,N_23896,N_23589);
nor U24460 (N_24460,N_23673,N_23796);
xor U24461 (N_24461,N_23738,N_23960);
or U24462 (N_24462,N_23919,N_23932);
and U24463 (N_24463,N_23785,N_23952);
and U24464 (N_24464,N_23627,N_23675);
nand U24465 (N_24465,N_23688,N_23975);
nand U24466 (N_24466,N_23840,N_23603);
and U24467 (N_24467,N_23829,N_23517);
nor U24468 (N_24468,N_23884,N_23739);
or U24469 (N_24469,N_23891,N_23793);
nand U24470 (N_24470,N_23858,N_23777);
and U24471 (N_24471,N_23916,N_23576);
xnor U24472 (N_24472,N_23646,N_23752);
nor U24473 (N_24473,N_23874,N_23937);
nor U24474 (N_24474,N_23613,N_23661);
or U24475 (N_24475,N_23519,N_23902);
nand U24476 (N_24476,N_23789,N_23970);
nand U24477 (N_24477,N_23791,N_23715);
nand U24478 (N_24478,N_23556,N_23998);
nand U24479 (N_24479,N_23658,N_23803);
nand U24480 (N_24480,N_23709,N_23784);
nor U24481 (N_24481,N_23627,N_23952);
nor U24482 (N_24482,N_23912,N_23756);
xnor U24483 (N_24483,N_23523,N_23551);
xor U24484 (N_24484,N_23756,N_23762);
nor U24485 (N_24485,N_23997,N_23584);
xor U24486 (N_24486,N_23551,N_23723);
nor U24487 (N_24487,N_23701,N_23782);
xnor U24488 (N_24488,N_23888,N_23850);
nor U24489 (N_24489,N_23907,N_23650);
nor U24490 (N_24490,N_23837,N_23586);
and U24491 (N_24491,N_23780,N_23894);
or U24492 (N_24492,N_23806,N_23956);
and U24493 (N_24493,N_23762,N_23995);
and U24494 (N_24494,N_23792,N_23789);
nor U24495 (N_24495,N_23601,N_23708);
nor U24496 (N_24496,N_23559,N_23565);
and U24497 (N_24497,N_23620,N_23982);
and U24498 (N_24498,N_23564,N_23740);
and U24499 (N_24499,N_23978,N_23713);
nor U24500 (N_24500,N_24110,N_24015);
and U24501 (N_24501,N_24227,N_24012);
and U24502 (N_24502,N_24433,N_24108);
and U24503 (N_24503,N_24048,N_24182);
nand U24504 (N_24504,N_24494,N_24203);
and U24505 (N_24505,N_24323,N_24296);
xor U24506 (N_24506,N_24249,N_24345);
and U24507 (N_24507,N_24208,N_24161);
and U24508 (N_24508,N_24109,N_24214);
or U24509 (N_24509,N_24282,N_24112);
nand U24510 (N_24510,N_24097,N_24240);
nand U24511 (N_24511,N_24285,N_24280);
xnor U24512 (N_24512,N_24144,N_24247);
or U24513 (N_24513,N_24423,N_24366);
xnor U24514 (N_24514,N_24429,N_24473);
xnor U24515 (N_24515,N_24353,N_24185);
nor U24516 (N_24516,N_24337,N_24133);
nor U24517 (N_24517,N_24452,N_24238);
or U24518 (N_24518,N_24224,N_24258);
and U24519 (N_24519,N_24082,N_24043);
nand U24520 (N_24520,N_24000,N_24404);
or U24521 (N_24521,N_24402,N_24127);
or U24522 (N_24522,N_24326,N_24276);
and U24523 (N_24523,N_24167,N_24071);
and U24524 (N_24524,N_24070,N_24001);
or U24525 (N_24525,N_24287,N_24119);
and U24526 (N_24526,N_24050,N_24122);
nand U24527 (N_24527,N_24039,N_24054);
xor U24528 (N_24528,N_24221,N_24320);
nor U24529 (N_24529,N_24078,N_24014);
nor U24530 (N_24530,N_24009,N_24324);
nor U24531 (N_24531,N_24106,N_24482);
or U24532 (N_24532,N_24341,N_24389);
and U24533 (N_24533,N_24448,N_24332);
xnor U24534 (N_24534,N_24467,N_24061);
and U24535 (N_24535,N_24250,N_24201);
nor U24536 (N_24536,N_24165,N_24496);
and U24537 (N_24537,N_24321,N_24450);
nand U24538 (N_24538,N_24325,N_24126);
xor U24539 (N_24539,N_24094,N_24319);
xor U24540 (N_24540,N_24168,N_24439);
xor U24541 (N_24541,N_24408,N_24474);
and U24542 (N_24542,N_24269,N_24184);
xor U24543 (N_24543,N_24057,N_24088);
or U24544 (N_24544,N_24425,N_24053);
xnor U24545 (N_24545,N_24355,N_24362);
xnor U24546 (N_24546,N_24351,N_24415);
nor U24547 (N_24547,N_24453,N_24431);
and U24548 (N_24548,N_24260,N_24489);
xor U24549 (N_24549,N_24485,N_24446);
xor U24550 (N_24550,N_24255,N_24116);
nor U24551 (N_24551,N_24022,N_24170);
and U24552 (N_24552,N_24449,N_24079);
or U24553 (N_24553,N_24229,N_24455);
nand U24554 (N_24554,N_24157,N_24234);
nand U24555 (N_24555,N_24040,N_24062);
nand U24556 (N_24556,N_24083,N_24420);
nand U24557 (N_24557,N_24178,N_24146);
nor U24558 (N_24558,N_24365,N_24373);
or U24559 (N_24559,N_24155,N_24141);
nand U24560 (N_24560,N_24414,N_24478);
xor U24561 (N_24561,N_24120,N_24021);
and U24562 (N_24562,N_24410,N_24328);
nor U24563 (N_24563,N_24498,N_24239);
or U24564 (N_24564,N_24322,N_24372);
nor U24565 (N_24565,N_24199,N_24244);
and U24566 (N_24566,N_24186,N_24150);
xnor U24567 (N_24567,N_24388,N_24253);
xor U24568 (N_24568,N_24016,N_24215);
or U24569 (N_24569,N_24153,N_24212);
nand U24570 (N_24570,N_24367,N_24472);
and U24571 (N_24571,N_24401,N_24207);
or U24572 (N_24572,N_24095,N_24052);
nand U24573 (N_24573,N_24035,N_24192);
nand U24574 (N_24574,N_24194,N_24067);
and U24575 (N_24575,N_24063,N_24298);
xor U24576 (N_24576,N_24064,N_24486);
or U24577 (N_24577,N_24292,N_24305);
nand U24578 (N_24578,N_24069,N_24018);
or U24579 (N_24579,N_24381,N_24445);
xor U24580 (N_24580,N_24166,N_24125);
xnor U24581 (N_24581,N_24123,N_24437);
nor U24582 (N_24582,N_24087,N_24219);
and U24583 (N_24583,N_24084,N_24045);
nand U24584 (N_24584,N_24159,N_24169);
nand U24585 (N_24585,N_24363,N_24430);
nor U24586 (N_24586,N_24347,N_24010);
nor U24587 (N_24587,N_24101,N_24147);
nor U24588 (N_24588,N_24136,N_24424);
nand U24589 (N_24589,N_24469,N_24162);
nor U24590 (N_24590,N_24304,N_24435);
and U24591 (N_24591,N_24311,N_24484);
nand U24592 (N_24592,N_24349,N_24172);
or U24593 (N_24593,N_24346,N_24313);
nor U24594 (N_24594,N_24190,N_24151);
nand U24595 (N_24595,N_24198,N_24137);
xnor U24596 (N_24596,N_24275,N_24114);
xnor U24597 (N_24597,N_24444,N_24460);
nor U24598 (N_24598,N_24300,N_24216);
nand U24599 (N_24599,N_24293,N_24377);
xnor U24600 (N_24600,N_24327,N_24027);
nor U24601 (N_24601,N_24392,N_24387);
and U24602 (N_24602,N_24391,N_24447);
or U24603 (N_24603,N_24409,N_24390);
nand U24604 (N_24604,N_24130,N_24090);
nand U24605 (N_24605,N_24111,N_24038);
nor U24606 (N_24606,N_24236,N_24107);
nor U24607 (N_24607,N_24196,N_24463);
nand U24608 (N_24608,N_24128,N_24217);
and U24609 (N_24609,N_24004,N_24359);
and U24610 (N_24610,N_24330,N_24066);
nand U24611 (N_24611,N_24357,N_24003);
and U24612 (N_24612,N_24174,N_24317);
nor U24613 (N_24613,N_24295,N_24418);
and U24614 (N_24614,N_24368,N_24499);
or U24615 (N_24615,N_24013,N_24393);
xor U24616 (N_24616,N_24149,N_24289);
or U24617 (N_24617,N_24100,N_24076);
nor U24618 (N_24618,N_24413,N_24060);
nand U24619 (N_24619,N_24375,N_24102);
nand U24620 (N_24620,N_24232,N_24183);
nor U24621 (N_24621,N_24020,N_24026);
xor U24622 (N_24622,N_24302,N_24342);
xnor U24623 (N_24623,N_24451,N_24188);
xor U24624 (N_24624,N_24271,N_24117);
xnor U24625 (N_24625,N_24344,N_24092);
or U24626 (N_24626,N_24281,N_24314);
and U24627 (N_24627,N_24180,N_24462);
or U24628 (N_24628,N_24243,N_24046);
nand U24629 (N_24629,N_24458,N_24055);
or U24630 (N_24630,N_24223,N_24075);
nand U24631 (N_24631,N_24029,N_24222);
nor U24632 (N_24632,N_24378,N_24025);
nor U24633 (N_24633,N_24442,N_24051);
or U24634 (N_24634,N_24428,N_24131);
nand U24635 (N_24635,N_24471,N_24307);
xor U24636 (N_24636,N_24086,N_24242);
nor U24637 (N_24637,N_24077,N_24422);
nand U24638 (N_24638,N_24354,N_24490);
nand U24639 (N_24639,N_24384,N_24274);
or U24640 (N_24640,N_24291,N_24339);
nor U24641 (N_24641,N_24041,N_24231);
nand U24642 (N_24642,N_24383,N_24350);
nand U24643 (N_24643,N_24370,N_24220);
nor U24644 (N_24644,N_24316,N_24140);
or U24645 (N_24645,N_24403,N_24273);
and U24646 (N_24646,N_24412,N_24397);
or U24647 (N_24647,N_24461,N_24118);
or U24648 (N_24648,N_24206,N_24252);
and U24649 (N_24649,N_24139,N_24115);
or U24650 (N_24650,N_24364,N_24036);
and U24651 (N_24651,N_24358,N_24308);
nand U24652 (N_24652,N_24254,N_24121);
xnor U24653 (N_24653,N_24187,N_24481);
or U24654 (N_24654,N_24411,N_24406);
nor U24655 (N_24655,N_24209,N_24369);
nor U24656 (N_24656,N_24104,N_24310);
and U24657 (N_24657,N_24135,N_24103);
or U24658 (N_24658,N_24479,N_24177);
or U24659 (N_24659,N_24290,N_24262);
and U24660 (N_24660,N_24356,N_24303);
or U24661 (N_24661,N_24024,N_24148);
nor U24662 (N_24662,N_24343,N_24158);
xnor U24663 (N_24663,N_24030,N_24241);
xnor U24664 (N_24664,N_24438,N_24205);
xor U24665 (N_24665,N_24400,N_24268);
and U24666 (N_24666,N_24031,N_24493);
nand U24667 (N_24667,N_24007,N_24008);
or U24668 (N_24668,N_24011,N_24475);
or U24669 (N_24669,N_24338,N_24470);
xnor U24670 (N_24670,N_24204,N_24210);
and U24671 (N_24671,N_24152,N_24416);
nor U24672 (N_24672,N_24081,N_24251);
and U24673 (N_24673,N_24405,N_24432);
nand U24674 (N_24674,N_24042,N_24047);
or U24675 (N_24675,N_24417,N_24468);
and U24676 (N_24676,N_24163,N_24318);
nand U24677 (N_24677,N_24352,N_24331);
nor U24678 (N_24678,N_24002,N_24028);
nand U24679 (N_24679,N_24226,N_24213);
xnor U24680 (N_24680,N_24134,N_24235);
nor U24681 (N_24681,N_24426,N_24443);
xor U24682 (N_24682,N_24261,N_24278);
nand U24683 (N_24683,N_24477,N_24495);
nand U24684 (N_24684,N_24113,N_24465);
nand U24685 (N_24685,N_24197,N_24492);
xnor U24686 (N_24686,N_24385,N_24164);
or U24687 (N_24687,N_24309,N_24456);
xnor U24688 (N_24688,N_24267,N_24074);
nand U24689 (N_24689,N_24264,N_24091);
or U24690 (N_24690,N_24360,N_24399);
or U24691 (N_24691,N_24138,N_24124);
xnor U24692 (N_24692,N_24419,N_24072);
and U24693 (N_24693,N_24265,N_24181);
or U24694 (N_24694,N_24297,N_24259);
xnor U24695 (N_24695,N_24089,N_24301);
nand U24696 (N_24696,N_24277,N_24098);
xor U24697 (N_24697,N_24099,N_24032);
or U24698 (N_24698,N_24398,N_24476);
or U24699 (N_24699,N_24132,N_24068);
or U24700 (N_24700,N_24270,N_24440);
nor U24701 (N_24701,N_24333,N_24245);
xor U24702 (N_24702,N_24263,N_24371);
or U24703 (N_24703,N_24459,N_24160);
xor U24704 (N_24704,N_24005,N_24211);
xor U24705 (N_24705,N_24237,N_24246);
and U24706 (N_24706,N_24173,N_24033);
or U24707 (N_24707,N_24193,N_24202);
nor U24708 (N_24708,N_24142,N_24218);
or U24709 (N_24709,N_24154,N_24480);
nand U24710 (N_24710,N_24491,N_24171);
xnor U24711 (N_24711,N_24065,N_24200);
xnor U24712 (N_24712,N_24497,N_24376);
xor U24713 (N_24713,N_24315,N_24306);
and U24714 (N_24714,N_24466,N_24017);
or U24715 (N_24715,N_24457,N_24248);
or U24716 (N_24716,N_24044,N_24195);
xnor U24717 (N_24717,N_24096,N_24037);
nand U24718 (N_24718,N_24394,N_24487);
xor U24719 (N_24719,N_24230,N_24374);
and U24720 (N_24720,N_24379,N_24488);
or U24721 (N_24721,N_24034,N_24176);
and U24722 (N_24722,N_24085,N_24407);
xor U24723 (N_24723,N_24256,N_24058);
nand U24724 (N_24724,N_24329,N_24019);
nand U24725 (N_24725,N_24059,N_24340);
xnor U24726 (N_24726,N_24179,N_24434);
nor U24727 (N_24727,N_24288,N_24056);
xor U24728 (N_24728,N_24421,N_24464);
nand U24729 (N_24729,N_24380,N_24233);
nor U24730 (N_24730,N_24272,N_24454);
or U24731 (N_24731,N_24279,N_24023);
nor U24732 (N_24732,N_24294,N_24006);
xnor U24733 (N_24733,N_24143,N_24283);
or U24734 (N_24734,N_24175,N_24228);
and U24735 (N_24735,N_24436,N_24336);
nor U24736 (N_24736,N_24483,N_24284);
nand U24737 (N_24737,N_24257,N_24286);
or U24738 (N_24738,N_24189,N_24129);
and U24739 (N_24739,N_24073,N_24395);
nand U24740 (N_24740,N_24386,N_24361);
and U24741 (N_24741,N_24105,N_24335);
and U24742 (N_24742,N_24225,N_24427);
nor U24743 (N_24743,N_24093,N_24441);
nand U24744 (N_24744,N_24191,N_24080);
and U24745 (N_24745,N_24396,N_24049);
xnor U24746 (N_24746,N_24299,N_24312);
and U24747 (N_24747,N_24266,N_24145);
and U24748 (N_24748,N_24334,N_24382);
nor U24749 (N_24749,N_24156,N_24348);
nand U24750 (N_24750,N_24455,N_24210);
nand U24751 (N_24751,N_24477,N_24064);
xnor U24752 (N_24752,N_24491,N_24109);
nor U24753 (N_24753,N_24030,N_24308);
and U24754 (N_24754,N_24264,N_24282);
nor U24755 (N_24755,N_24318,N_24360);
xnor U24756 (N_24756,N_24211,N_24033);
and U24757 (N_24757,N_24201,N_24490);
xor U24758 (N_24758,N_24467,N_24480);
and U24759 (N_24759,N_24344,N_24235);
nor U24760 (N_24760,N_24245,N_24257);
nor U24761 (N_24761,N_24114,N_24052);
or U24762 (N_24762,N_24247,N_24080);
xor U24763 (N_24763,N_24398,N_24375);
or U24764 (N_24764,N_24105,N_24366);
nor U24765 (N_24765,N_24492,N_24142);
or U24766 (N_24766,N_24071,N_24125);
and U24767 (N_24767,N_24264,N_24114);
xor U24768 (N_24768,N_24175,N_24454);
nand U24769 (N_24769,N_24016,N_24293);
and U24770 (N_24770,N_24454,N_24291);
or U24771 (N_24771,N_24074,N_24072);
nor U24772 (N_24772,N_24389,N_24018);
nand U24773 (N_24773,N_24147,N_24378);
or U24774 (N_24774,N_24277,N_24181);
nor U24775 (N_24775,N_24424,N_24183);
or U24776 (N_24776,N_24167,N_24051);
or U24777 (N_24777,N_24242,N_24255);
or U24778 (N_24778,N_24012,N_24395);
or U24779 (N_24779,N_24082,N_24124);
or U24780 (N_24780,N_24394,N_24106);
xnor U24781 (N_24781,N_24360,N_24073);
nor U24782 (N_24782,N_24399,N_24120);
nor U24783 (N_24783,N_24145,N_24303);
nor U24784 (N_24784,N_24090,N_24127);
nor U24785 (N_24785,N_24258,N_24349);
nor U24786 (N_24786,N_24124,N_24449);
and U24787 (N_24787,N_24102,N_24386);
nand U24788 (N_24788,N_24424,N_24005);
nor U24789 (N_24789,N_24040,N_24385);
xor U24790 (N_24790,N_24088,N_24313);
and U24791 (N_24791,N_24227,N_24198);
or U24792 (N_24792,N_24186,N_24013);
and U24793 (N_24793,N_24427,N_24079);
xor U24794 (N_24794,N_24278,N_24236);
or U24795 (N_24795,N_24019,N_24208);
and U24796 (N_24796,N_24024,N_24022);
and U24797 (N_24797,N_24437,N_24347);
nor U24798 (N_24798,N_24359,N_24296);
nor U24799 (N_24799,N_24318,N_24219);
or U24800 (N_24800,N_24433,N_24109);
or U24801 (N_24801,N_24242,N_24112);
or U24802 (N_24802,N_24111,N_24021);
or U24803 (N_24803,N_24410,N_24384);
and U24804 (N_24804,N_24331,N_24447);
nor U24805 (N_24805,N_24396,N_24375);
xor U24806 (N_24806,N_24091,N_24468);
nor U24807 (N_24807,N_24450,N_24269);
xnor U24808 (N_24808,N_24246,N_24195);
xnor U24809 (N_24809,N_24163,N_24098);
and U24810 (N_24810,N_24085,N_24147);
or U24811 (N_24811,N_24219,N_24458);
xnor U24812 (N_24812,N_24408,N_24208);
and U24813 (N_24813,N_24113,N_24130);
nand U24814 (N_24814,N_24298,N_24132);
or U24815 (N_24815,N_24388,N_24317);
or U24816 (N_24816,N_24343,N_24277);
or U24817 (N_24817,N_24368,N_24409);
xor U24818 (N_24818,N_24198,N_24480);
xnor U24819 (N_24819,N_24497,N_24199);
nand U24820 (N_24820,N_24084,N_24042);
xor U24821 (N_24821,N_24131,N_24381);
xor U24822 (N_24822,N_24308,N_24211);
xnor U24823 (N_24823,N_24040,N_24401);
xnor U24824 (N_24824,N_24247,N_24495);
and U24825 (N_24825,N_24085,N_24349);
nand U24826 (N_24826,N_24168,N_24468);
nor U24827 (N_24827,N_24048,N_24258);
xnor U24828 (N_24828,N_24269,N_24262);
xor U24829 (N_24829,N_24219,N_24343);
nand U24830 (N_24830,N_24134,N_24115);
or U24831 (N_24831,N_24105,N_24397);
nor U24832 (N_24832,N_24155,N_24038);
nand U24833 (N_24833,N_24430,N_24082);
nor U24834 (N_24834,N_24158,N_24310);
nand U24835 (N_24835,N_24324,N_24408);
nor U24836 (N_24836,N_24379,N_24425);
nand U24837 (N_24837,N_24360,N_24412);
and U24838 (N_24838,N_24478,N_24483);
and U24839 (N_24839,N_24333,N_24372);
or U24840 (N_24840,N_24130,N_24330);
nand U24841 (N_24841,N_24377,N_24205);
or U24842 (N_24842,N_24047,N_24103);
and U24843 (N_24843,N_24259,N_24372);
and U24844 (N_24844,N_24080,N_24378);
nand U24845 (N_24845,N_24480,N_24136);
or U24846 (N_24846,N_24111,N_24254);
xnor U24847 (N_24847,N_24417,N_24448);
xnor U24848 (N_24848,N_24273,N_24465);
and U24849 (N_24849,N_24238,N_24391);
xnor U24850 (N_24850,N_24388,N_24450);
nand U24851 (N_24851,N_24111,N_24125);
xnor U24852 (N_24852,N_24301,N_24226);
nand U24853 (N_24853,N_24117,N_24144);
or U24854 (N_24854,N_24282,N_24432);
or U24855 (N_24855,N_24016,N_24108);
nand U24856 (N_24856,N_24430,N_24266);
xor U24857 (N_24857,N_24264,N_24007);
nand U24858 (N_24858,N_24002,N_24497);
nor U24859 (N_24859,N_24498,N_24320);
or U24860 (N_24860,N_24128,N_24049);
nand U24861 (N_24861,N_24467,N_24059);
or U24862 (N_24862,N_24457,N_24210);
nor U24863 (N_24863,N_24225,N_24093);
and U24864 (N_24864,N_24347,N_24072);
or U24865 (N_24865,N_24495,N_24306);
and U24866 (N_24866,N_24291,N_24351);
or U24867 (N_24867,N_24386,N_24261);
nor U24868 (N_24868,N_24382,N_24097);
or U24869 (N_24869,N_24498,N_24337);
and U24870 (N_24870,N_24102,N_24474);
nand U24871 (N_24871,N_24306,N_24054);
xor U24872 (N_24872,N_24331,N_24044);
xor U24873 (N_24873,N_24196,N_24460);
or U24874 (N_24874,N_24328,N_24251);
or U24875 (N_24875,N_24367,N_24330);
and U24876 (N_24876,N_24350,N_24274);
and U24877 (N_24877,N_24279,N_24390);
and U24878 (N_24878,N_24052,N_24149);
and U24879 (N_24879,N_24073,N_24222);
nor U24880 (N_24880,N_24078,N_24331);
and U24881 (N_24881,N_24037,N_24360);
nand U24882 (N_24882,N_24498,N_24348);
xnor U24883 (N_24883,N_24410,N_24150);
nand U24884 (N_24884,N_24097,N_24481);
and U24885 (N_24885,N_24255,N_24421);
nand U24886 (N_24886,N_24435,N_24451);
nand U24887 (N_24887,N_24306,N_24175);
xnor U24888 (N_24888,N_24481,N_24350);
or U24889 (N_24889,N_24191,N_24311);
nor U24890 (N_24890,N_24377,N_24006);
and U24891 (N_24891,N_24291,N_24213);
and U24892 (N_24892,N_24035,N_24339);
and U24893 (N_24893,N_24250,N_24040);
nand U24894 (N_24894,N_24054,N_24402);
nor U24895 (N_24895,N_24321,N_24046);
nand U24896 (N_24896,N_24233,N_24394);
and U24897 (N_24897,N_24323,N_24196);
and U24898 (N_24898,N_24196,N_24456);
xnor U24899 (N_24899,N_24348,N_24470);
nand U24900 (N_24900,N_24283,N_24296);
or U24901 (N_24901,N_24238,N_24349);
and U24902 (N_24902,N_24388,N_24351);
nor U24903 (N_24903,N_24248,N_24069);
nor U24904 (N_24904,N_24141,N_24341);
and U24905 (N_24905,N_24431,N_24310);
xnor U24906 (N_24906,N_24389,N_24195);
nand U24907 (N_24907,N_24177,N_24453);
and U24908 (N_24908,N_24042,N_24016);
and U24909 (N_24909,N_24178,N_24141);
and U24910 (N_24910,N_24190,N_24463);
and U24911 (N_24911,N_24214,N_24263);
xor U24912 (N_24912,N_24425,N_24426);
and U24913 (N_24913,N_24148,N_24191);
xnor U24914 (N_24914,N_24496,N_24057);
nand U24915 (N_24915,N_24025,N_24417);
nand U24916 (N_24916,N_24447,N_24204);
or U24917 (N_24917,N_24489,N_24424);
nor U24918 (N_24918,N_24478,N_24002);
nand U24919 (N_24919,N_24085,N_24227);
xor U24920 (N_24920,N_24174,N_24156);
xor U24921 (N_24921,N_24376,N_24410);
or U24922 (N_24922,N_24423,N_24054);
nor U24923 (N_24923,N_24054,N_24384);
and U24924 (N_24924,N_24182,N_24027);
and U24925 (N_24925,N_24273,N_24412);
or U24926 (N_24926,N_24110,N_24172);
nor U24927 (N_24927,N_24150,N_24261);
nor U24928 (N_24928,N_24012,N_24067);
or U24929 (N_24929,N_24382,N_24465);
or U24930 (N_24930,N_24286,N_24472);
nor U24931 (N_24931,N_24383,N_24483);
nand U24932 (N_24932,N_24275,N_24188);
xor U24933 (N_24933,N_24021,N_24369);
xor U24934 (N_24934,N_24193,N_24259);
nor U24935 (N_24935,N_24265,N_24080);
and U24936 (N_24936,N_24218,N_24386);
and U24937 (N_24937,N_24470,N_24214);
or U24938 (N_24938,N_24415,N_24034);
or U24939 (N_24939,N_24336,N_24195);
nor U24940 (N_24940,N_24286,N_24358);
and U24941 (N_24941,N_24382,N_24246);
xnor U24942 (N_24942,N_24367,N_24263);
nand U24943 (N_24943,N_24095,N_24069);
or U24944 (N_24944,N_24010,N_24221);
xor U24945 (N_24945,N_24080,N_24041);
xnor U24946 (N_24946,N_24351,N_24454);
and U24947 (N_24947,N_24474,N_24019);
or U24948 (N_24948,N_24179,N_24165);
nor U24949 (N_24949,N_24335,N_24072);
or U24950 (N_24950,N_24024,N_24175);
and U24951 (N_24951,N_24052,N_24384);
or U24952 (N_24952,N_24026,N_24115);
or U24953 (N_24953,N_24494,N_24282);
nor U24954 (N_24954,N_24139,N_24102);
nand U24955 (N_24955,N_24288,N_24318);
nand U24956 (N_24956,N_24441,N_24351);
and U24957 (N_24957,N_24328,N_24346);
nand U24958 (N_24958,N_24096,N_24212);
or U24959 (N_24959,N_24356,N_24182);
or U24960 (N_24960,N_24083,N_24379);
nand U24961 (N_24961,N_24077,N_24210);
xnor U24962 (N_24962,N_24066,N_24085);
nand U24963 (N_24963,N_24153,N_24154);
or U24964 (N_24964,N_24005,N_24140);
nor U24965 (N_24965,N_24456,N_24032);
xor U24966 (N_24966,N_24060,N_24393);
nor U24967 (N_24967,N_24127,N_24076);
nand U24968 (N_24968,N_24210,N_24103);
nor U24969 (N_24969,N_24316,N_24420);
xor U24970 (N_24970,N_24129,N_24139);
xnor U24971 (N_24971,N_24371,N_24447);
or U24972 (N_24972,N_24135,N_24221);
nand U24973 (N_24973,N_24032,N_24146);
xor U24974 (N_24974,N_24033,N_24189);
nor U24975 (N_24975,N_24024,N_24044);
nand U24976 (N_24976,N_24297,N_24383);
and U24977 (N_24977,N_24461,N_24062);
nand U24978 (N_24978,N_24226,N_24228);
or U24979 (N_24979,N_24331,N_24114);
and U24980 (N_24980,N_24334,N_24156);
and U24981 (N_24981,N_24204,N_24016);
or U24982 (N_24982,N_24464,N_24063);
xnor U24983 (N_24983,N_24127,N_24025);
nor U24984 (N_24984,N_24333,N_24432);
and U24985 (N_24985,N_24018,N_24287);
nor U24986 (N_24986,N_24075,N_24037);
or U24987 (N_24987,N_24163,N_24031);
and U24988 (N_24988,N_24471,N_24292);
nand U24989 (N_24989,N_24096,N_24025);
and U24990 (N_24990,N_24390,N_24254);
or U24991 (N_24991,N_24037,N_24413);
or U24992 (N_24992,N_24138,N_24295);
nand U24993 (N_24993,N_24457,N_24349);
or U24994 (N_24994,N_24194,N_24161);
nand U24995 (N_24995,N_24452,N_24033);
nand U24996 (N_24996,N_24345,N_24325);
nor U24997 (N_24997,N_24110,N_24062);
and U24998 (N_24998,N_24237,N_24222);
xnor U24999 (N_24999,N_24306,N_24052);
nor UO_0 (O_0,N_24610,N_24508);
nand UO_1 (O_1,N_24523,N_24527);
nand UO_2 (O_2,N_24712,N_24884);
and UO_3 (O_3,N_24789,N_24997);
nor UO_4 (O_4,N_24931,N_24885);
and UO_5 (O_5,N_24574,N_24830);
or UO_6 (O_6,N_24655,N_24826);
and UO_7 (O_7,N_24647,N_24595);
xnor UO_8 (O_8,N_24736,N_24987);
nand UO_9 (O_9,N_24935,N_24719);
nand UO_10 (O_10,N_24823,N_24792);
and UO_11 (O_11,N_24876,N_24594);
nand UO_12 (O_12,N_24588,N_24536);
nor UO_13 (O_13,N_24977,N_24668);
nand UO_14 (O_14,N_24533,N_24962);
and UO_15 (O_15,N_24516,N_24653);
or UO_16 (O_16,N_24846,N_24985);
and UO_17 (O_17,N_24782,N_24708);
or UO_18 (O_18,N_24517,N_24903);
and UO_19 (O_19,N_24761,N_24905);
and UO_20 (O_20,N_24552,N_24752);
xor UO_21 (O_21,N_24968,N_24917);
or UO_22 (O_22,N_24857,N_24779);
or UO_23 (O_23,N_24577,N_24642);
nand UO_24 (O_24,N_24558,N_24981);
nand UO_25 (O_25,N_24855,N_24811);
or UO_26 (O_26,N_24735,N_24866);
xnor UO_27 (O_27,N_24747,N_24518);
xnor UO_28 (O_28,N_24827,N_24899);
or UO_29 (O_29,N_24716,N_24852);
nor UO_30 (O_30,N_24908,N_24996);
xor UO_31 (O_31,N_24744,N_24812);
and UO_32 (O_32,N_24848,N_24544);
xor UO_33 (O_33,N_24785,N_24913);
nand UO_34 (O_34,N_24788,N_24822);
nor UO_35 (O_35,N_24772,N_24550);
nor UO_36 (O_36,N_24870,N_24659);
nor UO_37 (O_37,N_24839,N_24835);
nand UO_38 (O_38,N_24769,N_24941);
or UO_39 (O_39,N_24863,N_24604);
nor UO_40 (O_40,N_24947,N_24620);
xor UO_41 (O_41,N_24740,N_24990);
and UO_42 (O_42,N_24691,N_24670);
and UO_43 (O_43,N_24581,N_24810);
or UO_44 (O_44,N_24572,N_24841);
nor UO_45 (O_45,N_24618,N_24893);
nand UO_46 (O_46,N_24695,N_24502);
xnor UO_47 (O_47,N_24722,N_24948);
xor UO_48 (O_48,N_24992,N_24613);
nand UO_49 (O_49,N_24749,N_24512);
nand UO_50 (O_50,N_24748,N_24529);
or UO_51 (O_51,N_24787,N_24560);
xnor UO_52 (O_52,N_24819,N_24809);
nand UO_53 (O_53,N_24532,N_24638);
xor UO_54 (O_54,N_24955,N_24765);
nor UO_55 (O_55,N_24878,N_24715);
or UO_56 (O_56,N_24936,N_24599);
nand UO_57 (O_57,N_24578,N_24704);
xor UO_58 (O_58,N_24733,N_24692);
nor UO_59 (O_59,N_24724,N_24543);
and UO_60 (O_60,N_24808,N_24907);
and UO_61 (O_61,N_24953,N_24616);
xnor UO_62 (O_62,N_24959,N_24801);
or UO_63 (O_63,N_24622,N_24764);
or UO_64 (O_64,N_24751,N_24989);
nor UO_65 (O_65,N_24753,N_24952);
xnor UO_66 (O_66,N_24859,N_24836);
or UO_67 (O_67,N_24698,N_24979);
nor UO_68 (O_68,N_24967,N_24937);
xor UO_69 (O_69,N_24851,N_24850);
nand UO_70 (O_70,N_24661,N_24795);
or UO_71 (O_71,N_24921,N_24684);
nor UO_72 (O_72,N_24540,N_24880);
nand UO_73 (O_73,N_24958,N_24528);
or UO_74 (O_74,N_24511,N_24983);
and UO_75 (O_75,N_24793,N_24842);
xnor UO_76 (O_76,N_24549,N_24807);
or UO_77 (O_77,N_24680,N_24662);
xnor UO_78 (O_78,N_24978,N_24566);
and UO_79 (O_79,N_24521,N_24554);
nor UO_80 (O_80,N_24526,N_24825);
nor UO_81 (O_81,N_24824,N_24910);
xnor UO_82 (O_82,N_24615,N_24843);
and UO_83 (O_83,N_24929,N_24689);
nand UO_84 (O_84,N_24710,N_24833);
and UO_85 (O_85,N_24513,N_24702);
nand UO_86 (O_86,N_24760,N_24798);
and UO_87 (O_87,N_24856,N_24541);
xor UO_88 (O_88,N_24950,N_24547);
or UO_89 (O_89,N_24777,N_24865);
nand UO_90 (O_90,N_24551,N_24898);
xnor UO_91 (O_91,N_24582,N_24831);
or UO_92 (O_92,N_24963,N_24636);
and UO_93 (O_93,N_24961,N_24858);
nand UO_94 (O_94,N_24573,N_24754);
or UO_95 (O_95,N_24780,N_24840);
and UO_96 (O_96,N_24562,N_24598);
or UO_97 (O_97,N_24703,N_24862);
nor UO_98 (O_98,N_24816,N_24556);
nor UO_99 (O_99,N_24994,N_24901);
nand UO_100 (O_100,N_24944,N_24699);
xor UO_101 (O_101,N_24663,N_24970);
xnor UO_102 (O_102,N_24804,N_24732);
and UO_103 (O_103,N_24739,N_24694);
nand UO_104 (O_104,N_24927,N_24817);
nor UO_105 (O_105,N_24814,N_24806);
nand UO_106 (O_106,N_24771,N_24510);
or UO_107 (O_107,N_24626,N_24646);
xor UO_108 (O_108,N_24794,N_24845);
or UO_109 (O_109,N_24575,N_24586);
and UO_110 (O_110,N_24624,N_24776);
xor UO_111 (O_111,N_24534,N_24632);
or UO_112 (O_112,N_24949,N_24974);
nand UO_113 (O_113,N_24688,N_24922);
or UO_114 (O_114,N_24677,N_24709);
and UO_115 (O_115,N_24643,N_24943);
nor UO_116 (O_116,N_24993,N_24531);
xor UO_117 (O_117,N_24686,N_24741);
nand UO_118 (O_118,N_24768,N_24685);
nand UO_119 (O_119,N_24999,N_24998);
nor UO_120 (O_120,N_24726,N_24844);
nor UO_121 (O_121,N_24828,N_24797);
nand UO_122 (O_122,N_24660,N_24611);
nand UO_123 (O_123,N_24894,N_24627);
nand UO_124 (O_124,N_24759,N_24909);
nand UO_125 (O_125,N_24860,N_24916);
nand UO_126 (O_126,N_24890,N_24501);
xor UO_127 (O_127,N_24743,N_24886);
nand UO_128 (O_128,N_24631,N_24891);
xnor UO_129 (O_129,N_24973,N_24639);
or UO_130 (O_130,N_24939,N_24766);
nand UO_131 (O_131,N_24881,N_24567);
and UO_132 (O_132,N_24681,N_24538);
nor UO_133 (O_133,N_24569,N_24892);
and UO_134 (O_134,N_24900,N_24614);
or UO_135 (O_135,N_24606,N_24720);
and UO_136 (O_136,N_24565,N_24889);
nand UO_137 (O_137,N_24774,N_24915);
xor UO_138 (O_138,N_24644,N_24770);
or UO_139 (O_139,N_24679,N_24854);
xnor UO_140 (O_140,N_24867,N_24932);
and UO_141 (O_141,N_24803,N_24602);
and UO_142 (O_142,N_24656,N_24934);
xnor UO_143 (O_143,N_24911,N_24637);
and UO_144 (O_144,N_24737,N_24621);
xor UO_145 (O_145,N_24951,N_24729);
nand UO_146 (O_146,N_24954,N_24727);
nand UO_147 (O_147,N_24665,N_24904);
or UO_148 (O_148,N_24925,N_24589);
and UO_149 (O_149,N_24942,N_24887);
nor UO_150 (O_150,N_24995,N_24813);
nand UO_151 (O_151,N_24635,N_24832);
or UO_152 (O_152,N_24877,N_24971);
nand UO_153 (O_153,N_24930,N_24802);
nor UO_154 (O_154,N_24861,N_24649);
xor UO_155 (O_155,N_24964,N_24714);
nor UO_156 (O_156,N_24781,N_24984);
nand UO_157 (O_157,N_24975,N_24707);
xor UO_158 (O_158,N_24869,N_24555);
and UO_159 (O_159,N_24778,N_24864);
xor UO_160 (O_160,N_24587,N_24683);
nor UO_161 (O_161,N_24918,N_24608);
xnor UO_162 (O_162,N_24514,N_24628);
nand UO_163 (O_163,N_24906,N_24553);
nor UO_164 (O_164,N_24838,N_24730);
or UO_165 (O_165,N_24956,N_24799);
and UO_166 (O_166,N_24612,N_24652);
and UO_167 (O_167,N_24507,N_24522);
and UO_168 (O_168,N_24701,N_24597);
and UO_169 (O_169,N_24601,N_24821);
nor UO_170 (O_170,N_24966,N_24868);
and UO_171 (O_171,N_24731,N_24920);
xor UO_172 (O_172,N_24607,N_24596);
or UO_173 (O_173,N_24693,N_24897);
and UO_174 (O_174,N_24734,N_24982);
nand UO_175 (O_175,N_24713,N_24666);
and UO_176 (O_176,N_24658,N_24609);
and UO_177 (O_177,N_24525,N_24590);
nor UO_178 (O_178,N_24874,N_24576);
xor UO_179 (O_179,N_24758,N_24834);
nor UO_180 (O_180,N_24675,N_24928);
or UO_181 (O_181,N_24912,N_24650);
and UO_182 (O_182,N_24537,N_24746);
nor UO_183 (O_183,N_24773,N_24509);
or UO_184 (O_184,N_24548,N_24568);
nor UO_185 (O_185,N_24506,N_24672);
nor UO_186 (O_186,N_24756,N_24940);
nand UO_187 (O_187,N_24938,N_24671);
or UO_188 (O_188,N_24515,N_24657);
or UO_189 (O_189,N_24593,N_24700);
or UO_190 (O_190,N_24505,N_24718);
nand UO_191 (O_191,N_24592,N_24539);
and UO_192 (O_192,N_24853,N_24738);
nor UO_193 (O_193,N_24969,N_24728);
or UO_194 (O_194,N_24674,N_24634);
or UO_195 (O_195,N_24546,N_24872);
nand UO_196 (O_196,N_24564,N_24600);
xnor UO_197 (O_197,N_24725,N_24717);
xnor UO_198 (O_198,N_24883,N_24585);
xor UO_199 (O_199,N_24640,N_24914);
nor UO_200 (O_200,N_24757,N_24623);
nand UO_201 (O_201,N_24617,N_24545);
or UO_202 (O_202,N_24641,N_24767);
nor UO_203 (O_203,N_24775,N_24721);
nand UO_204 (O_204,N_24625,N_24705);
or UO_205 (O_205,N_24960,N_24629);
nand UO_206 (O_206,N_24619,N_24557);
and UO_207 (O_207,N_24697,N_24790);
nand UO_208 (O_208,N_24711,N_24820);
nand UO_209 (O_209,N_24815,N_24991);
nor UO_210 (O_210,N_24882,N_24957);
xor UO_211 (O_211,N_24745,N_24896);
xor UO_212 (O_212,N_24676,N_24630);
nor UO_213 (O_213,N_24669,N_24919);
xnor UO_214 (O_214,N_24933,N_24678);
xor UO_215 (O_215,N_24875,N_24603);
xnor UO_216 (O_216,N_24519,N_24879);
nor UO_217 (O_217,N_24706,N_24902);
nor UO_218 (O_218,N_24762,N_24524);
and UO_219 (O_219,N_24988,N_24980);
and UO_220 (O_220,N_24696,N_24648);
nor UO_221 (O_221,N_24924,N_24682);
nor UO_222 (O_222,N_24654,N_24645);
and UO_223 (O_223,N_24500,N_24895);
or UO_224 (O_224,N_24561,N_24796);
and UO_225 (O_225,N_24579,N_24584);
nand UO_226 (O_226,N_24535,N_24976);
and UO_227 (O_227,N_24784,N_24580);
xnor UO_228 (O_228,N_24791,N_24926);
nor UO_229 (O_229,N_24542,N_24888);
xor UO_230 (O_230,N_24965,N_24873);
xnor UO_231 (O_231,N_24829,N_24986);
and UO_232 (O_232,N_24583,N_24849);
xnor UO_233 (O_233,N_24847,N_24786);
or UO_234 (O_234,N_24520,N_24687);
and UO_235 (O_235,N_24591,N_24805);
nand UO_236 (O_236,N_24651,N_24503);
xnor UO_237 (O_237,N_24673,N_24972);
xor UO_238 (O_238,N_24763,N_24664);
nand UO_239 (O_239,N_24871,N_24818);
nand UO_240 (O_240,N_24750,N_24742);
and UO_241 (O_241,N_24633,N_24723);
nor UO_242 (O_242,N_24571,N_24504);
nor UO_243 (O_243,N_24690,N_24563);
xor UO_244 (O_244,N_24923,N_24783);
nand UO_245 (O_245,N_24945,N_24667);
xnor UO_246 (O_246,N_24570,N_24559);
and UO_247 (O_247,N_24946,N_24837);
and UO_248 (O_248,N_24755,N_24605);
nor UO_249 (O_249,N_24530,N_24800);
and UO_250 (O_250,N_24728,N_24685);
nand UO_251 (O_251,N_24700,N_24791);
nor UO_252 (O_252,N_24537,N_24699);
nand UO_253 (O_253,N_24608,N_24800);
xor UO_254 (O_254,N_24500,N_24528);
xor UO_255 (O_255,N_24586,N_24941);
nor UO_256 (O_256,N_24610,N_24801);
xnor UO_257 (O_257,N_24761,N_24823);
nor UO_258 (O_258,N_24583,N_24900);
xnor UO_259 (O_259,N_24884,N_24742);
nor UO_260 (O_260,N_24692,N_24902);
nor UO_261 (O_261,N_24883,N_24628);
and UO_262 (O_262,N_24965,N_24586);
nand UO_263 (O_263,N_24535,N_24848);
nand UO_264 (O_264,N_24857,N_24674);
nand UO_265 (O_265,N_24755,N_24545);
nand UO_266 (O_266,N_24809,N_24903);
or UO_267 (O_267,N_24633,N_24851);
nand UO_268 (O_268,N_24711,N_24636);
or UO_269 (O_269,N_24592,N_24654);
nand UO_270 (O_270,N_24666,N_24790);
xnor UO_271 (O_271,N_24519,N_24664);
nor UO_272 (O_272,N_24734,N_24933);
or UO_273 (O_273,N_24554,N_24968);
or UO_274 (O_274,N_24996,N_24679);
xor UO_275 (O_275,N_24736,N_24729);
xor UO_276 (O_276,N_24642,N_24748);
nor UO_277 (O_277,N_24781,N_24681);
xor UO_278 (O_278,N_24517,N_24994);
and UO_279 (O_279,N_24797,N_24667);
and UO_280 (O_280,N_24933,N_24993);
and UO_281 (O_281,N_24789,N_24621);
and UO_282 (O_282,N_24522,N_24550);
and UO_283 (O_283,N_24737,N_24509);
and UO_284 (O_284,N_24914,N_24843);
and UO_285 (O_285,N_24821,N_24737);
or UO_286 (O_286,N_24711,N_24623);
nand UO_287 (O_287,N_24681,N_24804);
xnor UO_288 (O_288,N_24782,N_24594);
xor UO_289 (O_289,N_24604,N_24831);
and UO_290 (O_290,N_24801,N_24797);
nor UO_291 (O_291,N_24638,N_24665);
nor UO_292 (O_292,N_24721,N_24805);
and UO_293 (O_293,N_24619,N_24646);
nor UO_294 (O_294,N_24921,N_24724);
or UO_295 (O_295,N_24574,N_24842);
nor UO_296 (O_296,N_24711,N_24602);
or UO_297 (O_297,N_24966,N_24618);
or UO_298 (O_298,N_24820,N_24707);
nor UO_299 (O_299,N_24905,N_24984);
nand UO_300 (O_300,N_24592,N_24661);
and UO_301 (O_301,N_24723,N_24830);
and UO_302 (O_302,N_24801,N_24637);
nor UO_303 (O_303,N_24985,N_24968);
or UO_304 (O_304,N_24858,N_24600);
nor UO_305 (O_305,N_24841,N_24781);
or UO_306 (O_306,N_24976,N_24882);
xnor UO_307 (O_307,N_24809,N_24642);
or UO_308 (O_308,N_24870,N_24527);
nor UO_309 (O_309,N_24862,N_24646);
and UO_310 (O_310,N_24861,N_24636);
and UO_311 (O_311,N_24687,N_24875);
or UO_312 (O_312,N_24798,N_24639);
and UO_313 (O_313,N_24737,N_24735);
and UO_314 (O_314,N_24702,N_24931);
nand UO_315 (O_315,N_24777,N_24683);
nand UO_316 (O_316,N_24730,N_24974);
or UO_317 (O_317,N_24994,N_24746);
xnor UO_318 (O_318,N_24674,N_24720);
or UO_319 (O_319,N_24625,N_24634);
nand UO_320 (O_320,N_24564,N_24508);
and UO_321 (O_321,N_24839,N_24606);
nor UO_322 (O_322,N_24986,N_24962);
xnor UO_323 (O_323,N_24631,N_24820);
nor UO_324 (O_324,N_24557,N_24991);
nand UO_325 (O_325,N_24818,N_24615);
nand UO_326 (O_326,N_24709,N_24861);
and UO_327 (O_327,N_24884,N_24730);
xnor UO_328 (O_328,N_24820,N_24685);
nand UO_329 (O_329,N_24674,N_24583);
nand UO_330 (O_330,N_24718,N_24770);
nor UO_331 (O_331,N_24791,N_24625);
xor UO_332 (O_332,N_24527,N_24789);
or UO_333 (O_333,N_24621,N_24706);
or UO_334 (O_334,N_24509,N_24642);
xor UO_335 (O_335,N_24915,N_24808);
xnor UO_336 (O_336,N_24950,N_24958);
nand UO_337 (O_337,N_24539,N_24723);
nand UO_338 (O_338,N_24689,N_24979);
nand UO_339 (O_339,N_24577,N_24809);
xor UO_340 (O_340,N_24987,N_24509);
xor UO_341 (O_341,N_24579,N_24505);
nand UO_342 (O_342,N_24696,N_24710);
nor UO_343 (O_343,N_24507,N_24624);
nor UO_344 (O_344,N_24678,N_24508);
and UO_345 (O_345,N_24864,N_24918);
nand UO_346 (O_346,N_24693,N_24559);
xor UO_347 (O_347,N_24596,N_24588);
nand UO_348 (O_348,N_24690,N_24954);
xor UO_349 (O_349,N_24588,N_24819);
nand UO_350 (O_350,N_24685,N_24916);
and UO_351 (O_351,N_24530,N_24533);
nand UO_352 (O_352,N_24778,N_24716);
and UO_353 (O_353,N_24960,N_24855);
and UO_354 (O_354,N_24916,N_24588);
or UO_355 (O_355,N_24544,N_24840);
nor UO_356 (O_356,N_24708,N_24745);
and UO_357 (O_357,N_24697,N_24654);
and UO_358 (O_358,N_24872,N_24901);
xnor UO_359 (O_359,N_24904,N_24612);
and UO_360 (O_360,N_24820,N_24558);
nor UO_361 (O_361,N_24575,N_24604);
or UO_362 (O_362,N_24929,N_24859);
nor UO_363 (O_363,N_24559,N_24624);
xnor UO_364 (O_364,N_24725,N_24619);
or UO_365 (O_365,N_24691,N_24864);
nand UO_366 (O_366,N_24875,N_24634);
or UO_367 (O_367,N_24541,N_24825);
nand UO_368 (O_368,N_24924,N_24841);
or UO_369 (O_369,N_24712,N_24584);
or UO_370 (O_370,N_24562,N_24841);
nor UO_371 (O_371,N_24664,N_24900);
or UO_372 (O_372,N_24809,N_24838);
and UO_373 (O_373,N_24649,N_24946);
or UO_374 (O_374,N_24896,N_24882);
and UO_375 (O_375,N_24844,N_24660);
nor UO_376 (O_376,N_24995,N_24987);
and UO_377 (O_377,N_24838,N_24754);
nand UO_378 (O_378,N_24799,N_24870);
or UO_379 (O_379,N_24658,N_24862);
and UO_380 (O_380,N_24703,N_24613);
or UO_381 (O_381,N_24957,N_24721);
nor UO_382 (O_382,N_24999,N_24644);
nor UO_383 (O_383,N_24598,N_24662);
or UO_384 (O_384,N_24573,N_24639);
nor UO_385 (O_385,N_24536,N_24711);
and UO_386 (O_386,N_24932,N_24907);
and UO_387 (O_387,N_24890,N_24982);
and UO_388 (O_388,N_24635,N_24649);
or UO_389 (O_389,N_24606,N_24963);
or UO_390 (O_390,N_24680,N_24924);
or UO_391 (O_391,N_24914,N_24603);
nor UO_392 (O_392,N_24884,N_24581);
xnor UO_393 (O_393,N_24913,N_24717);
xnor UO_394 (O_394,N_24900,N_24817);
and UO_395 (O_395,N_24772,N_24560);
and UO_396 (O_396,N_24606,N_24825);
and UO_397 (O_397,N_24851,N_24688);
nand UO_398 (O_398,N_24646,N_24675);
and UO_399 (O_399,N_24992,N_24939);
nand UO_400 (O_400,N_24524,N_24710);
or UO_401 (O_401,N_24942,N_24790);
and UO_402 (O_402,N_24611,N_24610);
and UO_403 (O_403,N_24891,N_24958);
or UO_404 (O_404,N_24889,N_24727);
nor UO_405 (O_405,N_24929,N_24894);
nor UO_406 (O_406,N_24840,N_24758);
and UO_407 (O_407,N_24781,N_24670);
nor UO_408 (O_408,N_24882,N_24765);
nand UO_409 (O_409,N_24796,N_24648);
nand UO_410 (O_410,N_24523,N_24799);
nand UO_411 (O_411,N_24679,N_24812);
nor UO_412 (O_412,N_24999,N_24980);
or UO_413 (O_413,N_24839,N_24814);
and UO_414 (O_414,N_24898,N_24937);
and UO_415 (O_415,N_24639,N_24783);
nor UO_416 (O_416,N_24764,N_24954);
nand UO_417 (O_417,N_24951,N_24646);
and UO_418 (O_418,N_24884,N_24905);
nor UO_419 (O_419,N_24507,N_24714);
or UO_420 (O_420,N_24686,N_24693);
xnor UO_421 (O_421,N_24770,N_24943);
nand UO_422 (O_422,N_24742,N_24971);
or UO_423 (O_423,N_24976,N_24954);
nor UO_424 (O_424,N_24683,N_24922);
or UO_425 (O_425,N_24683,N_24571);
nor UO_426 (O_426,N_24890,N_24508);
nand UO_427 (O_427,N_24525,N_24882);
nand UO_428 (O_428,N_24959,N_24636);
or UO_429 (O_429,N_24736,N_24745);
or UO_430 (O_430,N_24522,N_24627);
nor UO_431 (O_431,N_24502,N_24954);
or UO_432 (O_432,N_24891,N_24693);
nor UO_433 (O_433,N_24749,N_24907);
xnor UO_434 (O_434,N_24954,N_24745);
nor UO_435 (O_435,N_24613,N_24964);
and UO_436 (O_436,N_24837,N_24775);
nor UO_437 (O_437,N_24619,N_24832);
nor UO_438 (O_438,N_24730,N_24710);
and UO_439 (O_439,N_24934,N_24705);
and UO_440 (O_440,N_24848,N_24802);
nand UO_441 (O_441,N_24777,N_24914);
or UO_442 (O_442,N_24543,N_24512);
nor UO_443 (O_443,N_24635,N_24787);
nand UO_444 (O_444,N_24931,N_24604);
nand UO_445 (O_445,N_24606,N_24968);
xor UO_446 (O_446,N_24849,N_24665);
nor UO_447 (O_447,N_24548,N_24542);
nor UO_448 (O_448,N_24743,N_24748);
and UO_449 (O_449,N_24970,N_24693);
nor UO_450 (O_450,N_24560,N_24619);
nor UO_451 (O_451,N_24830,N_24585);
nor UO_452 (O_452,N_24629,N_24657);
xor UO_453 (O_453,N_24736,N_24726);
and UO_454 (O_454,N_24697,N_24730);
nand UO_455 (O_455,N_24619,N_24989);
and UO_456 (O_456,N_24915,N_24701);
and UO_457 (O_457,N_24932,N_24942);
nand UO_458 (O_458,N_24592,N_24972);
and UO_459 (O_459,N_24680,N_24788);
nand UO_460 (O_460,N_24627,N_24969);
nand UO_461 (O_461,N_24786,N_24591);
and UO_462 (O_462,N_24950,N_24717);
or UO_463 (O_463,N_24997,N_24823);
nor UO_464 (O_464,N_24724,N_24872);
nand UO_465 (O_465,N_24578,N_24723);
or UO_466 (O_466,N_24604,N_24912);
or UO_467 (O_467,N_24743,N_24897);
and UO_468 (O_468,N_24925,N_24809);
nor UO_469 (O_469,N_24709,N_24625);
and UO_470 (O_470,N_24932,N_24594);
nand UO_471 (O_471,N_24833,N_24842);
or UO_472 (O_472,N_24652,N_24692);
xnor UO_473 (O_473,N_24871,N_24632);
nand UO_474 (O_474,N_24859,N_24591);
nand UO_475 (O_475,N_24510,N_24961);
nor UO_476 (O_476,N_24879,N_24715);
nor UO_477 (O_477,N_24567,N_24897);
or UO_478 (O_478,N_24656,N_24797);
nor UO_479 (O_479,N_24585,N_24877);
and UO_480 (O_480,N_24623,N_24557);
or UO_481 (O_481,N_24909,N_24842);
or UO_482 (O_482,N_24561,N_24665);
and UO_483 (O_483,N_24669,N_24987);
xnor UO_484 (O_484,N_24728,N_24610);
and UO_485 (O_485,N_24778,N_24973);
xor UO_486 (O_486,N_24601,N_24830);
nor UO_487 (O_487,N_24948,N_24629);
nor UO_488 (O_488,N_24539,N_24646);
or UO_489 (O_489,N_24985,N_24593);
nand UO_490 (O_490,N_24968,N_24662);
and UO_491 (O_491,N_24638,N_24825);
nand UO_492 (O_492,N_24659,N_24920);
or UO_493 (O_493,N_24950,N_24647);
xor UO_494 (O_494,N_24920,N_24918);
xnor UO_495 (O_495,N_24543,N_24955);
xnor UO_496 (O_496,N_24628,N_24548);
and UO_497 (O_497,N_24741,N_24579);
and UO_498 (O_498,N_24754,N_24712);
nor UO_499 (O_499,N_24871,N_24748);
nand UO_500 (O_500,N_24740,N_24592);
nand UO_501 (O_501,N_24808,N_24942);
nor UO_502 (O_502,N_24780,N_24674);
nand UO_503 (O_503,N_24827,N_24523);
xor UO_504 (O_504,N_24972,N_24962);
nand UO_505 (O_505,N_24955,N_24515);
and UO_506 (O_506,N_24901,N_24568);
xor UO_507 (O_507,N_24606,N_24822);
and UO_508 (O_508,N_24649,N_24650);
nand UO_509 (O_509,N_24564,N_24840);
xor UO_510 (O_510,N_24784,N_24808);
nand UO_511 (O_511,N_24509,N_24824);
or UO_512 (O_512,N_24796,N_24779);
xnor UO_513 (O_513,N_24913,N_24730);
nand UO_514 (O_514,N_24957,N_24822);
and UO_515 (O_515,N_24739,N_24939);
xor UO_516 (O_516,N_24567,N_24628);
and UO_517 (O_517,N_24796,N_24577);
nand UO_518 (O_518,N_24705,N_24536);
xor UO_519 (O_519,N_24975,N_24743);
or UO_520 (O_520,N_24799,N_24686);
and UO_521 (O_521,N_24743,N_24761);
nor UO_522 (O_522,N_24847,N_24583);
xnor UO_523 (O_523,N_24587,N_24830);
nand UO_524 (O_524,N_24871,N_24958);
nor UO_525 (O_525,N_24567,N_24856);
and UO_526 (O_526,N_24618,N_24624);
and UO_527 (O_527,N_24679,N_24855);
nor UO_528 (O_528,N_24822,N_24758);
nand UO_529 (O_529,N_24746,N_24669);
nand UO_530 (O_530,N_24564,N_24671);
nand UO_531 (O_531,N_24679,N_24885);
xor UO_532 (O_532,N_24547,N_24523);
or UO_533 (O_533,N_24673,N_24579);
nor UO_534 (O_534,N_24641,N_24693);
xnor UO_535 (O_535,N_24813,N_24920);
nor UO_536 (O_536,N_24634,N_24550);
and UO_537 (O_537,N_24589,N_24628);
xor UO_538 (O_538,N_24873,N_24666);
and UO_539 (O_539,N_24569,N_24928);
nor UO_540 (O_540,N_24594,N_24813);
and UO_541 (O_541,N_24744,N_24749);
nor UO_542 (O_542,N_24754,N_24514);
and UO_543 (O_543,N_24576,N_24996);
or UO_544 (O_544,N_24580,N_24993);
or UO_545 (O_545,N_24984,N_24921);
xor UO_546 (O_546,N_24524,N_24711);
nand UO_547 (O_547,N_24927,N_24575);
or UO_548 (O_548,N_24608,N_24553);
xnor UO_549 (O_549,N_24927,N_24744);
and UO_550 (O_550,N_24914,N_24702);
xor UO_551 (O_551,N_24915,N_24538);
and UO_552 (O_552,N_24809,N_24785);
and UO_553 (O_553,N_24697,N_24672);
or UO_554 (O_554,N_24886,N_24593);
nand UO_555 (O_555,N_24727,N_24845);
nor UO_556 (O_556,N_24828,N_24957);
or UO_557 (O_557,N_24594,N_24652);
and UO_558 (O_558,N_24835,N_24927);
or UO_559 (O_559,N_24891,N_24836);
or UO_560 (O_560,N_24711,N_24886);
nor UO_561 (O_561,N_24657,N_24936);
xnor UO_562 (O_562,N_24826,N_24837);
xnor UO_563 (O_563,N_24593,N_24719);
and UO_564 (O_564,N_24736,N_24579);
or UO_565 (O_565,N_24957,N_24764);
xor UO_566 (O_566,N_24631,N_24626);
and UO_567 (O_567,N_24988,N_24779);
nor UO_568 (O_568,N_24864,N_24946);
or UO_569 (O_569,N_24596,N_24854);
nand UO_570 (O_570,N_24722,N_24932);
and UO_571 (O_571,N_24990,N_24634);
xor UO_572 (O_572,N_24633,N_24879);
nand UO_573 (O_573,N_24805,N_24942);
nor UO_574 (O_574,N_24949,N_24891);
or UO_575 (O_575,N_24937,N_24555);
or UO_576 (O_576,N_24849,N_24853);
and UO_577 (O_577,N_24612,N_24934);
nor UO_578 (O_578,N_24709,N_24859);
and UO_579 (O_579,N_24619,N_24687);
xnor UO_580 (O_580,N_24740,N_24973);
xnor UO_581 (O_581,N_24828,N_24776);
nor UO_582 (O_582,N_24780,N_24917);
or UO_583 (O_583,N_24514,N_24794);
and UO_584 (O_584,N_24713,N_24962);
or UO_585 (O_585,N_24675,N_24558);
or UO_586 (O_586,N_24959,N_24655);
nand UO_587 (O_587,N_24928,N_24517);
and UO_588 (O_588,N_24657,N_24610);
and UO_589 (O_589,N_24531,N_24585);
xnor UO_590 (O_590,N_24890,N_24503);
xor UO_591 (O_591,N_24548,N_24906);
xor UO_592 (O_592,N_24906,N_24910);
xnor UO_593 (O_593,N_24709,N_24564);
xor UO_594 (O_594,N_24763,N_24554);
nor UO_595 (O_595,N_24786,N_24644);
nand UO_596 (O_596,N_24958,N_24568);
and UO_597 (O_597,N_24810,N_24971);
nor UO_598 (O_598,N_24746,N_24823);
nand UO_599 (O_599,N_24603,N_24988);
nor UO_600 (O_600,N_24633,N_24615);
xor UO_601 (O_601,N_24953,N_24958);
or UO_602 (O_602,N_24908,N_24778);
nor UO_603 (O_603,N_24502,N_24806);
nand UO_604 (O_604,N_24683,N_24622);
and UO_605 (O_605,N_24797,N_24581);
or UO_606 (O_606,N_24842,N_24850);
nand UO_607 (O_607,N_24701,N_24967);
nand UO_608 (O_608,N_24895,N_24577);
nor UO_609 (O_609,N_24944,N_24746);
xnor UO_610 (O_610,N_24922,N_24740);
nor UO_611 (O_611,N_24529,N_24602);
and UO_612 (O_612,N_24966,N_24675);
and UO_613 (O_613,N_24951,N_24628);
xnor UO_614 (O_614,N_24858,N_24998);
nand UO_615 (O_615,N_24795,N_24813);
xor UO_616 (O_616,N_24734,N_24896);
nor UO_617 (O_617,N_24666,N_24573);
and UO_618 (O_618,N_24713,N_24948);
nor UO_619 (O_619,N_24501,N_24546);
nand UO_620 (O_620,N_24769,N_24999);
nand UO_621 (O_621,N_24579,N_24855);
or UO_622 (O_622,N_24924,N_24634);
nor UO_623 (O_623,N_24668,N_24874);
or UO_624 (O_624,N_24730,N_24929);
nor UO_625 (O_625,N_24932,N_24891);
nor UO_626 (O_626,N_24912,N_24930);
and UO_627 (O_627,N_24752,N_24874);
nor UO_628 (O_628,N_24610,N_24542);
and UO_629 (O_629,N_24790,N_24671);
nand UO_630 (O_630,N_24756,N_24848);
nand UO_631 (O_631,N_24501,N_24767);
xor UO_632 (O_632,N_24580,N_24999);
xnor UO_633 (O_633,N_24595,N_24525);
or UO_634 (O_634,N_24760,N_24763);
and UO_635 (O_635,N_24700,N_24571);
and UO_636 (O_636,N_24725,N_24594);
and UO_637 (O_637,N_24978,N_24641);
or UO_638 (O_638,N_24563,N_24739);
nand UO_639 (O_639,N_24912,N_24697);
nand UO_640 (O_640,N_24829,N_24892);
nor UO_641 (O_641,N_24736,N_24646);
and UO_642 (O_642,N_24591,N_24627);
or UO_643 (O_643,N_24663,N_24793);
nand UO_644 (O_644,N_24966,N_24674);
or UO_645 (O_645,N_24588,N_24580);
xnor UO_646 (O_646,N_24768,N_24959);
nand UO_647 (O_647,N_24931,N_24516);
or UO_648 (O_648,N_24698,N_24507);
and UO_649 (O_649,N_24759,N_24764);
nor UO_650 (O_650,N_24600,N_24536);
nor UO_651 (O_651,N_24583,N_24717);
nand UO_652 (O_652,N_24632,N_24526);
xor UO_653 (O_653,N_24547,N_24708);
and UO_654 (O_654,N_24727,N_24549);
or UO_655 (O_655,N_24992,N_24765);
xnor UO_656 (O_656,N_24956,N_24736);
and UO_657 (O_657,N_24612,N_24566);
and UO_658 (O_658,N_24853,N_24632);
or UO_659 (O_659,N_24905,N_24974);
and UO_660 (O_660,N_24747,N_24967);
and UO_661 (O_661,N_24879,N_24565);
or UO_662 (O_662,N_24538,N_24849);
nand UO_663 (O_663,N_24969,N_24616);
and UO_664 (O_664,N_24889,N_24790);
xor UO_665 (O_665,N_24953,N_24886);
or UO_666 (O_666,N_24943,N_24797);
and UO_667 (O_667,N_24613,N_24918);
nand UO_668 (O_668,N_24871,N_24787);
xnor UO_669 (O_669,N_24817,N_24580);
and UO_670 (O_670,N_24747,N_24547);
and UO_671 (O_671,N_24985,N_24604);
nor UO_672 (O_672,N_24946,N_24996);
nand UO_673 (O_673,N_24584,N_24969);
and UO_674 (O_674,N_24728,N_24787);
xnor UO_675 (O_675,N_24958,N_24762);
and UO_676 (O_676,N_24730,N_24703);
nand UO_677 (O_677,N_24650,N_24548);
and UO_678 (O_678,N_24597,N_24787);
or UO_679 (O_679,N_24967,N_24971);
nor UO_680 (O_680,N_24742,N_24506);
xor UO_681 (O_681,N_24851,N_24962);
and UO_682 (O_682,N_24676,N_24846);
nand UO_683 (O_683,N_24719,N_24944);
or UO_684 (O_684,N_24587,N_24704);
nand UO_685 (O_685,N_24793,N_24767);
nor UO_686 (O_686,N_24571,N_24932);
or UO_687 (O_687,N_24937,N_24743);
and UO_688 (O_688,N_24965,N_24761);
nor UO_689 (O_689,N_24868,N_24741);
nor UO_690 (O_690,N_24534,N_24797);
or UO_691 (O_691,N_24705,N_24720);
or UO_692 (O_692,N_24883,N_24713);
and UO_693 (O_693,N_24846,N_24814);
xnor UO_694 (O_694,N_24852,N_24593);
xor UO_695 (O_695,N_24911,N_24969);
xor UO_696 (O_696,N_24744,N_24563);
or UO_697 (O_697,N_24757,N_24621);
nand UO_698 (O_698,N_24941,N_24809);
or UO_699 (O_699,N_24971,N_24814);
and UO_700 (O_700,N_24531,N_24893);
nor UO_701 (O_701,N_24697,N_24752);
or UO_702 (O_702,N_24529,N_24750);
nand UO_703 (O_703,N_24960,N_24816);
or UO_704 (O_704,N_24828,N_24680);
nand UO_705 (O_705,N_24696,N_24747);
nand UO_706 (O_706,N_24534,N_24977);
xor UO_707 (O_707,N_24892,N_24645);
and UO_708 (O_708,N_24545,N_24933);
and UO_709 (O_709,N_24963,N_24625);
xnor UO_710 (O_710,N_24996,N_24600);
or UO_711 (O_711,N_24840,N_24607);
xor UO_712 (O_712,N_24562,N_24543);
and UO_713 (O_713,N_24580,N_24732);
nand UO_714 (O_714,N_24958,N_24930);
and UO_715 (O_715,N_24903,N_24989);
xnor UO_716 (O_716,N_24520,N_24707);
xor UO_717 (O_717,N_24512,N_24670);
nand UO_718 (O_718,N_24645,N_24568);
nand UO_719 (O_719,N_24935,N_24699);
nand UO_720 (O_720,N_24853,N_24942);
nor UO_721 (O_721,N_24990,N_24629);
nor UO_722 (O_722,N_24609,N_24600);
nand UO_723 (O_723,N_24732,N_24726);
xnor UO_724 (O_724,N_24690,N_24929);
xnor UO_725 (O_725,N_24757,N_24551);
nor UO_726 (O_726,N_24987,N_24881);
nor UO_727 (O_727,N_24562,N_24803);
nand UO_728 (O_728,N_24630,N_24691);
nor UO_729 (O_729,N_24942,N_24597);
or UO_730 (O_730,N_24554,N_24709);
or UO_731 (O_731,N_24880,N_24765);
xnor UO_732 (O_732,N_24860,N_24618);
or UO_733 (O_733,N_24894,N_24561);
xor UO_734 (O_734,N_24556,N_24746);
or UO_735 (O_735,N_24826,N_24704);
nand UO_736 (O_736,N_24779,N_24531);
xnor UO_737 (O_737,N_24980,N_24543);
nand UO_738 (O_738,N_24658,N_24995);
or UO_739 (O_739,N_24600,N_24748);
and UO_740 (O_740,N_24727,N_24814);
xnor UO_741 (O_741,N_24513,N_24884);
nor UO_742 (O_742,N_24677,N_24559);
nand UO_743 (O_743,N_24975,N_24812);
and UO_744 (O_744,N_24522,N_24875);
nand UO_745 (O_745,N_24642,N_24927);
or UO_746 (O_746,N_24535,N_24972);
or UO_747 (O_747,N_24664,N_24621);
nor UO_748 (O_748,N_24862,N_24734);
nor UO_749 (O_749,N_24852,N_24504);
xnor UO_750 (O_750,N_24759,N_24856);
and UO_751 (O_751,N_24927,N_24943);
xnor UO_752 (O_752,N_24907,N_24601);
nand UO_753 (O_753,N_24536,N_24551);
and UO_754 (O_754,N_24872,N_24541);
and UO_755 (O_755,N_24601,N_24974);
and UO_756 (O_756,N_24636,N_24580);
nand UO_757 (O_757,N_24676,N_24819);
xor UO_758 (O_758,N_24553,N_24745);
xnor UO_759 (O_759,N_24707,N_24910);
xor UO_760 (O_760,N_24975,N_24702);
xnor UO_761 (O_761,N_24654,N_24566);
nand UO_762 (O_762,N_24812,N_24752);
or UO_763 (O_763,N_24642,N_24703);
nor UO_764 (O_764,N_24704,N_24935);
nor UO_765 (O_765,N_24759,N_24535);
nand UO_766 (O_766,N_24891,N_24549);
nand UO_767 (O_767,N_24727,N_24972);
xnor UO_768 (O_768,N_24949,N_24518);
nor UO_769 (O_769,N_24654,N_24647);
and UO_770 (O_770,N_24681,N_24730);
xnor UO_771 (O_771,N_24508,N_24539);
and UO_772 (O_772,N_24739,N_24895);
and UO_773 (O_773,N_24919,N_24830);
nand UO_774 (O_774,N_24721,N_24923);
nand UO_775 (O_775,N_24749,N_24791);
nor UO_776 (O_776,N_24699,N_24999);
nand UO_777 (O_777,N_24914,N_24841);
nor UO_778 (O_778,N_24569,N_24505);
and UO_779 (O_779,N_24875,N_24879);
xor UO_780 (O_780,N_24941,N_24799);
xnor UO_781 (O_781,N_24687,N_24795);
and UO_782 (O_782,N_24818,N_24751);
nor UO_783 (O_783,N_24891,N_24687);
or UO_784 (O_784,N_24606,N_24820);
or UO_785 (O_785,N_24587,N_24829);
or UO_786 (O_786,N_24733,N_24746);
nand UO_787 (O_787,N_24672,N_24734);
or UO_788 (O_788,N_24734,N_24619);
or UO_789 (O_789,N_24997,N_24737);
xnor UO_790 (O_790,N_24776,N_24909);
or UO_791 (O_791,N_24533,N_24752);
or UO_792 (O_792,N_24733,N_24773);
or UO_793 (O_793,N_24600,N_24567);
nor UO_794 (O_794,N_24715,N_24616);
and UO_795 (O_795,N_24575,N_24976);
nand UO_796 (O_796,N_24898,N_24538);
and UO_797 (O_797,N_24773,N_24532);
and UO_798 (O_798,N_24943,N_24807);
nand UO_799 (O_799,N_24662,N_24984);
or UO_800 (O_800,N_24727,N_24794);
xor UO_801 (O_801,N_24988,N_24867);
xnor UO_802 (O_802,N_24719,N_24687);
xor UO_803 (O_803,N_24522,N_24667);
xor UO_804 (O_804,N_24855,N_24905);
and UO_805 (O_805,N_24913,N_24644);
nand UO_806 (O_806,N_24584,N_24763);
or UO_807 (O_807,N_24869,N_24683);
and UO_808 (O_808,N_24981,N_24667);
nor UO_809 (O_809,N_24937,N_24551);
xnor UO_810 (O_810,N_24940,N_24949);
xor UO_811 (O_811,N_24617,N_24764);
or UO_812 (O_812,N_24763,N_24548);
xnor UO_813 (O_813,N_24901,N_24910);
or UO_814 (O_814,N_24762,N_24508);
nand UO_815 (O_815,N_24661,N_24891);
or UO_816 (O_816,N_24579,N_24786);
and UO_817 (O_817,N_24617,N_24725);
xor UO_818 (O_818,N_24521,N_24792);
or UO_819 (O_819,N_24555,N_24577);
and UO_820 (O_820,N_24901,N_24917);
or UO_821 (O_821,N_24758,N_24902);
or UO_822 (O_822,N_24854,N_24945);
nand UO_823 (O_823,N_24672,N_24771);
nand UO_824 (O_824,N_24701,N_24955);
nor UO_825 (O_825,N_24561,N_24586);
or UO_826 (O_826,N_24575,N_24627);
and UO_827 (O_827,N_24658,N_24974);
and UO_828 (O_828,N_24670,N_24972);
nand UO_829 (O_829,N_24631,N_24949);
and UO_830 (O_830,N_24676,N_24901);
and UO_831 (O_831,N_24588,N_24908);
xor UO_832 (O_832,N_24609,N_24631);
nor UO_833 (O_833,N_24708,N_24638);
nor UO_834 (O_834,N_24877,N_24559);
or UO_835 (O_835,N_24712,N_24631);
and UO_836 (O_836,N_24734,N_24573);
xnor UO_837 (O_837,N_24910,N_24685);
and UO_838 (O_838,N_24539,N_24634);
or UO_839 (O_839,N_24952,N_24763);
xnor UO_840 (O_840,N_24602,N_24626);
nand UO_841 (O_841,N_24917,N_24559);
or UO_842 (O_842,N_24628,N_24600);
nand UO_843 (O_843,N_24751,N_24662);
or UO_844 (O_844,N_24701,N_24755);
xnor UO_845 (O_845,N_24733,N_24589);
nand UO_846 (O_846,N_24953,N_24977);
nand UO_847 (O_847,N_24635,N_24799);
or UO_848 (O_848,N_24712,N_24605);
and UO_849 (O_849,N_24879,N_24919);
nor UO_850 (O_850,N_24610,N_24654);
nand UO_851 (O_851,N_24961,N_24629);
nand UO_852 (O_852,N_24698,N_24885);
nand UO_853 (O_853,N_24760,N_24749);
or UO_854 (O_854,N_24978,N_24991);
nor UO_855 (O_855,N_24760,N_24907);
nand UO_856 (O_856,N_24612,N_24902);
and UO_857 (O_857,N_24895,N_24834);
xnor UO_858 (O_858,N_24600,N_24653);
xnor UO_859 (O_859,N_24586,N_24572);
and UO_860 (O_860,N_24936,N_24895);
nand UO_861 (O_861,N_24846,N_24533);
and UO_862 (O_862,N_24721,N_24870);
or UO_863 (O_863,N_24895,N_24924);
xnor UO_864 (O_864,N_24753,N_24720);
or UO_865 (O_865,N_24837,N_24922);
xor UO_866 (O_866,N_24962,N_24528);
and UO_867 (O_867,N_24971,N_24823);
xnor UO_868 (O_868,N_24571,N_24557);
xor UO_869 (O_869,N_24770,N_24648);
xor UO_870 (O_870,N_24712,N_24734);
xnor UO_871 (O_871,N_24808,N_24631);
xor UO_872 (O_872,N_24787,N_24847);
nand UO_873 (O_873,N_24751,N_24579);
nand UO_874 (O_874,N_24849,N_24962);
xnor UO_875 (O_875,N_24806,N_24527);
and UO_876 (O_876,N_24612,N_24772);
or UO_877 (O_877,N_24731,N_24591);
or UO_878 (O_878,N_24551,N_24768);
or UO_879 (O_879,N_24863,N_24753);
and UO_880 (O_880,N_24920,N_24823);
xor UO_881 (O_881,N_24730,N_24993);
nand UO_882 (O_882,N_24727,N_24772);
or UO_883 (O_883,N_24669,N_24666);
nand UO_884 (O_884,N_24802,N_24994);
xnor UO_885 (O_885,N_24518,N_24934);
nor UO_886 (O_886,N_24880,N_24754);
or UO_887 (O_887,N_24697,N_24505);
or UO_888 (O_888,N_24596,N_24663);
xnor UO_889 (O_889,N_24572,N_24850);
nand UO_890 (O_890,N_24861,N_24723);
or UO_891 (O_891,N_24792,N_24628);
xor UO_892 (O_892,N_24933,N_24675);
xor UO_893 (O_893,N_24701,N_24609);
or UO_894 (O_894,N_24762,N_24680);
xor UO_895 (O_895,N_24988,N_24906);
nand UO_896 (O_896,N_24905,N_24629);
xnor UO_897 (O_897,N_24639,N_24614);
xnor UO_898 (O_898,N_24992,N_24951);
or UO_899 (O_899,N_24624,N_24878);
xor UO_900 (O_900,N_24938,N_24720);
nand UO_901 (O_901,N_24959,N_24904);
nand UO_902 (O_902,N_24618,N_24895);
nand UO_903 (O_903,N_24553,N_24932);
nor UO_904 (O_904,N_24710,N_24538);
xnor UO_905 (O_905,N_24540,N_24700);
and UO_906 (O_906,N_24579,N_24746);
or UO_907 (O_907,N_24916,N_24824);
nand UO_908 (O_908,N_24898,N_24648);
nand UO_909 (O_909,N_24558,N_24638);
nor UO_910 (O_910,N_24779,N_24759);
and UO_911 (O_911,N_24551,N_24553);
nand UO_912 (O_912,N_24950,N_24925);
nand UO_913 (O_913,N_24552,N_24905);
nand UO_914 (O_914,N_24625,N_24556);
xor UO_915 (O_915,N_24978,N_24940);
nand UO_916 (O_916,N_24693,N_24972);
xor UO_917 (O_917,N_24829,N_24901);
and UO_918 (O_918,N_24778,N_24678);
xnor UO_919 (O_919,N_24542,N_24722);
nor UO_920 (O_920,N_24524,N_24577);
and UO_921 (O_921,N_24726,N_24879);
and UO_922 (O_922,N_24961,N_24923);
xor UO_923 (O_923,N_24520,N_24795);
nand UO_924 (O_924,N_24882,N_24998);
or UO_925 (O_925,N_24922,N_24763);
nor UO_926 (O_926,N_24730,N_24686);
or UO_927 (O_927,N_24834,N_24737);
xnor UO_928 (O_928,N_24797,N_24716);
xnor UO_929 (O_929,N_24617,N_24795);
nand UO_930 (O_930,N_24510,N_24907);
xnor UO_931 (O_931,N_24676,N_24936);
or UO_932 (O_932,N_24935,N_24529);
and UO_933 (O_933,N_24791,N_24706);
or UO_934 (O_934,N_24684,N_24729);
xnor UO_935 (O_935,N_24633,N_24919);
xnor UO_936 (O_936,N_24538,N_24574);
nand UO_937 (O_937,N_24652,N_24962);
or UO_938 (O_938,N_24928,N_24762);
nor UO_939 (O_939,N_24671,N_24699);
or UO_940 (O_940,N_24642,N_24966);
nand UO_941 (O_941,N_24769,N_24526);
and UO_942 (O_942,N_24629,N_24606);
and UO_943 (O_943,N_24591,N_24574);
xnor UO_944 (O_944,N_24782,N_24984);
xor UO_945 (O_945,N_24732,N_24877);
and UO_946 (O_946,N_24731,N_24683);
nor UO_947 (O_947,N_24660,N_24872);
xnor UO_948 (O_948,N_24539,N_24649);
or UO_949 (O_949,N_24581,N_24531);
nor UO_950 (O_950,N_24893,N_24661);
or UO_951 (O_951,N_24630,N_24900);
nand UO_952 (O_952,N_24692,N_24809);
nor UO_953 (O_953,N_24689,N_24802);
or UO_954 (O_954,N_24840,N_24583);
xnor UO_955 (O_955,N_24620,N_24734);
nand UO_956 (O_956,N_24590,N_24580);
or UO_957 (O_957,N_24811,N_24755);
xor UO_958 (O_958,N_24997,N_24954);
nand UO_959 (O_959,N_24666,N_24826);
nor UO_960 (O_960,N_24814,N_24717);
nand UO_961 (O_961,N_24587,N_24766);
or UO_962 (O_962,N_24771,N_24990);
nor UO_963 (O_963,N_24706,N_24586);
xor UO_964 (O_964,N_24938,N_24832);
nand UO_965 (O_965,N_24505,N_24957);
nor UO_966 (O_966,N_24603,N_24970);
and UO_967 (O_967,N_24695,N_24930);
nand UO_968 (O_968,N_24818,N_24600);
nor UO_969 (O_969,N_24650,N_24598);
nor UO_970 (O_970,N_24915,N_24928);
nand UO_971 (O_971,N_24976,N_24738);
xor UO_972 (O_972,N_24588,N_24841);
nand UO_973 (O_973,N_24685,N_24903);
xor UO_974 (O_974,N_24828,N_24976);
or UO_975 (O_975,N_24508,N_24609);
or UO_976 (O_976,N_24905,N_24621);
xnor UO_977 (O_977,N_24861,N_24967);
or UO_978 (O_978,N_24967,N_24581);
or UO_979 (O_979,N_24938,N_24887);
nor UO_980 (O_980,N_24906,N_24754);
and UO_981 (O_981,N_24899,N_24559);
nand UO_982 (O_982,N_24981,N_24554);
nand UO_983 (O_983,N_24646,N_24607);
nor UO_984 (O_984,N_24537,N_24863);
nor UO_985 (O_985,N_24735,N_24613);
or UO_986 (O_986,N_24706,N_24873);
nor UO_987 (O_987,N_24838,N_24567);
nor UO_988 (O_988,N_24944,N_24838);
or UO_989 (O_989,N_24922,N_24605);
nor UO_990 (O_990,N_24765,N_24730);
or UO_991 (O_991,N_24646,N_24827);
and UO_992 (O_992,N_24527,N_24940);
and UO_993 (O_993,N_24673,N_24825);
and UO_994 (O_994,N_24754,N_24666);
or UO_995 (O_995,N_24708,N_24661);
or UO_996 (O_996,N_24654,N_24637);
nor UO_997 (O_997,N_24867,N_24827);
nand UO_998 (O_998,N_24992,N_24956);
nor UO_999 (O_999,N_24734,N_24803);
or UO_1000 (O_1000,N_24963,N_24825);
xor UO_1001 (O_1001,N_24571,N_24912);
nor UO_1002 (O_1002,N_24620,N_24523);
or UO_1003 (O_1003,N_24731,N_24693);
xnor UO_1004 (O_1004,N_24667,N_24549);
xor UO_1005 (O_1005,N_24843,N_24838);
nand UO_1006 (O_1006,N_24814,N_24754);
or UO_1007 (O_1007,N_24992,N_24531);
nor UO_1008 (O_1008,N_24811,N_24972);
nand UO_1009 (O_1009,N_24940,N_24712);
nor UO_1010 (O_1010,N_24784,N_24898);
nand UO_1011 (O_1011,N_24872,N_24691);
and UO_1012 (O_1012,N_24773,N_24551);
xnor UO_1013 (O_1013,N_24719,N_24756);
xor UO_1014 (O_1014,N_24706,N_24636);
nand UO_1015 (O_1015,N_24541,N_24764);
or UO_1016 (O_1016,N_24978,N_24853);
nor UO_1017 (O_1017,N_24895,N_24542);
xnor UO_1018 (O_1018,N_24536,N_24736);
and UO_1019 (O_1019,N_24834,N_24935);
nor UO_1020 (O_1020,N_24611,N_24937);
or UO_1021 (O_1021,N_24761,N_24908);
or UO_1022 (O_1022,N_24709,N_24989);
or UO_1023 (O_1023,N_24550,N_24870);
or UO_1024 (O_1024,N_24632,N_24504);
and UO_1025 (O_1025,N_24914,N_24648);
xnor UO_1026 (O_1026,N_24589,N_24832);
or UO_1027 (O_1027,N_24950,N_24553);
nor UO_1028 (O_1028,N_24638,N_24790);
or UO_1029 (O_1029,N_24744,N_24533);
xor UO_1030 (O_1030,N_24773,N_24945);
and UO_1031 (O_1031,N_24927,N_24851);
and UO_1032 (O_1032,N_24844,N_24965);
or UO_1033 (O_1033,N_24622,N_24519);
nand UO_1034 (O_1034,N_24976,N_24905);
and UO_1035 (O_1035,N_24569,N_24907);
xor UO_1036 (O_1036,N_24774,N_24580);
nor UO_1037 (O_1037,N_24700,N_24565);
nand UO_1038 (O_1038,N_24649,N_24763);
and UO_1039 (O_1039,N_24835,N_24759);
or UO_1040 (O_1040,N_24995,N_24843);
nor UO_1041 (O_1041,N_24606,N_24984);
and UO_1042 (O_1042,N_24814,N_24988);
nand UO_1043 (O_1043,N_24579,N_24999);
nand UO_1044 (O_1044,N_24563,N_24858);
nand UO_1045 (O_1045,N_24631,N_24758);
xor UO_1046 (O_1046,N_24977,N_24777);
nand UO_1047 (O_1047,N_24727,N_24615);
or UO_1048 (O_1048,N_24841,N_24815);
xor UO_1049 (O_1049,N_24946,N_24570);
nand UO_1050 (O_1050,N_24884,N_24664);
or UO_1051 (O_1051,N_24639,N_24574);
nand UO_1052 (O_1052,N_24836,N_24504);
xnor UO_1053 (O_1053,N_24672,N_24984);
xnor UO_1054 (O_1054,N_24713,N_24961);
or UO_1055 (O_1055,N_24867,N_24568);
xor UO_1056 (O_1056,N_24704,N_24538);
nand UO_1057 (O_1057,N_24657,N_24890);
nand UO_1058 (O_1058,N_24816,N_24853);
xor UO_1059 (O_1059,N_24718,N_24942);
nand UO_1060 (O_1060,N_24859,N_24650);
nand UO_1061 (O_1061,N_24697,N_24608);
or UO_1062 (O_1062,N_24604,N_24977);
and UO_1063 (O_1063,N_24899,N_24572);
nand UO_1064 (O_1064,N_24802,N_24511);
and UO_1065 (O_1065,N_24754,N_24615);
xnor UO_1066 (O_1066,N_24872,N_24941);
or UO_1067 (O_1067,N_24641,N_24537);
nand UO_1068 (O_1068,N_24639,N_24771);
and UO_1069 (O_1069,N_24893,N_24818);
and UO_1070 (O_1070,N_24978,N_24714);
or UO_1071 (O_1071,N_24660,N_24924);
nor UO_1072 (O_1072,N_24765,N_24889);
or UO_1073 (O_1073,N_24814,N_24530);
and UO_1074 (O_1074,N_24988,N_24827);
nand UO_1075 (O_1075,N_24540,N_24871);
xnor UO_1076 (O_1076,N_24890,N_24796);
xnor UO_1077 (O_1077,N_24540,N_24628);
nor UO_1078 (O_1078,N_24900,N_24727);
xnor UO_1079 (O_1079,N_24654,N_24738);
or UO_1080 (O_1080,N_24754,N_24931);
xnor UO_1081 (O_1081,N_24580,N_24911);
nand UO_1082 (O_1082,N_24615,N_24559);
nand UO_1083 (O_1083,N_24507,N_24953);
and UO_1084 (O_1084,N_24931,N_24805);
or UO_1085 (O_1085,N_24984,N_24654);
xnor UO_1086 (O_1086,N_24552,N_24609);
nand UO_1087 (O_1087,N_24982,N_24694);
xnor UO_1088 (O_1088,N_24827,N_24987);
and UO_1089 (O_1089,N_24642,N_24886);
and UO_1090 (O_1090,N_24554,N_24744);
xnor UO_1091 (O_1091,N_24745,N_24633);
xnor UO_1092 (O_1092,N_24623,N_24534);
or UO_1093 (O_1093,N_24594,N_24854);
nand UO_1094 (O_1094,N_24757,N_24559);
nor UO_1095 (O_1095,N_24624,N_24721);
nand UO_1096 (O_1096,N_24992,N_24985);
or UO_1097 (O_1097,N_24995,N_24580);
nand UO_1098 (O_1098,N_24551,N_24589);
xnor UO_1099 (O_1099,N_24573,N_24509);
and UO_1100 (O_1100,N_24792,N_24917);
nor UO_1101 (O_1101,N_24709,N_24669);
and UO_1102 (O_1102,N_24749,N_24990);
and UO_1103 (O_1103,N_24906,N_24623);
and UO_1104 (O_1104,N_24813,N_24799);
nor UO_1105 (O_1105,N_24881,N_24819);
or UO_1106 (O_1106,N_24792,N_24957);
nand UO_1107 (O_1107,N_24934,N_24994);
and UO_1108 (O_1108,N_24559,N_24798);
xor UO_1109 (O_1109,N_24628,N_24556);
and UO_1110 (O_1110,N_24989,N_24798);
and UO_1111 (O_1111,N_24847,N_24613);
or UO_1112 (O_1112,N_24982,N_24845);
or UO_1113 (O_1113,N_24808,N_24543);
or UO_1114 (O_1114,N_24744,N_24661);
or UO_1115 (O_1115,N_24996,N_24670);
and UO_1116 (O_1116,N_24663,N_24989);
xor UO_1117 (O_1117,N_24689,N_24569);
nand UO_1118 (O_1118,N_24957,N_24922);
nor UO_1119 (O_1119,N_24579,N_24833);
nor UO_1120 (O_1120,N_24929,N_24881);
nor UO_1121 (O_1121,N_24990,N_24778);
nand UO_1122 (O_1122,N_24719,N_24982);
xor UO_1123 (O_1123,N_24947,N_24503);
and UO_1124 (O_1124,N_24923,N_24736);
nor UO_1125 (O_1125,N_24575,N_24668);
xnor UO_1126 (O_1126,N_24901,N_24911);
xor UO_1127 (O_1127,N_24835,N_24701);
and UO_1128 (O_1128,N_24840,N_24787);
or UO_1129 (O_1129,N_24529,N_24738);
xor UO_1130 (O_1130,N_24796,N_24734);
and UO_1131 (O_1131,N_24725,N_24902);
nand UO_1132 (O_1132,N_24786,N_24762);
or UO_1133 (O_1133,N_24873,N_24970);
nor UO_1134 (O_1134,N_24966,N_24921);
nand UO_1135 (O_1135,N_24611,N_24627);
xnor UO_1136 (O_1136,N_24992,N_24904);
nor UO_1137 (O_1137,N_24569,N_24795);
or UO_1138 (O_1138,N_24919,N_24533);
and UO_1139 (O_1139,N_24635,N_24692);
and UO_1140 (O_1140,N_24537,N_24995);
and UO_1141 (O_1141,N_24588,N_24718);
xnor UO_1142 (O_1142,N_24567,N_24982);
nor UO_1143 (O_1143,N_24652,N_24972);
or UO_1144 (O_1144,N_24671,N_24655);
or UO_1145 (O_1145,N_24709,N_24512);
nor UO_1146 (O_1146,N_24938,N_24953);
nand UO_1147 (O_1147,N_24929,N_24557);
xnor UO_1148 (O_1148,N_24884,N_24523);
and UO_1149 (O_1149,N_24639,N_24822);
nor UO_1150 (O_1150,N_24953,N_24717);
nand UO_1151 (O_1151,N_24885,N_24732);
and UO_1152 (O_1152,N_24803,N_24561);
nor UO_1153 (O_1153,N_24505,N_24771);
xor UO_1154 (O_1154,N_24812,N_24677);
or UO_1155 (O_1155,N_24909,N_24967);
or UO_1156 (O_1156,N_24970,N_24686);
nor UO_1157 (O_1157,N_24744,N_24951);
and UO_1158 (O_1158,N_24589,N_24795);
nor UO_1159 (O_1159,N_24931,N_24691);
and UO_1160 (O_1160,N_24586,N_24554);
nand UO_1161 (O_1161,N_24592,N_24915);
nand UO_1162 (O_1162,N_24594,N_24622);
nand UO_1163 (O_1163,N_24793,N_24617);
or UO_1164 (O_1164,N_24909,N_24625);
or UO_1165 (O_1165,N_24601,N_24618);
nand UO_1166 (O_1166,N_24901,N_24915);
nand UO_1167 (O_1167,N_24778,N_24718);
nor UO_1168 (O_1168,N_24693,N_24937);
nand UO_1169 (O_1169,N_24508,N_24506);
xnor UO_1170 (O_1170,N_24799,N_24960);
or UO_1171 (O_1171,N_24612,N_24563);
and UO_1172 (O_1172,N_24983,N_24805);
nor UO_1173 (O_1173,N_24585,N_24634);
xor UO_1174 (O_1174,N_24995,N_24723);
xor UO_1175 (O_1175,N_24835,N_24758);
xor UO_1176 (O_1176,N_24686,N_24882);
and UO_1177 (O_1177,N_24974,N_24997);
xor UO_1178 (O_1178,N_24828,N_24643);
and UO_1179 (O_1179,N_24975,N_24726);
xor UO_1180 (O_1180,N_24546,N_24512);
nor UO_1181 (O_1181,N_24659,N_24733);
or UO_1182 (O_1182,N_24651,N_24905);
nor UO_1183 (O_1183,N_24700,N_24537);
and UO_1184 (O_1184,N_24692,N_24996);
and UO_1185 (O_1185,N_24551,N_24950);
xor UO_1186 (O_1186,N_24764,N_24978);
or UO_1187 (O_1187,N_24929,N_24994);
nor UO_1188 (O_1188,N_24855,N_24745);
nor UO_1189 (O_1189,N_24851,N_24675);
nand UO_1190 (O_1190,N_24616,N_24534);
or UO_1191 (O_1191,N_24596,N_24543);
nor UO_1192 (O_1192,N_24596,N_24638);
and UO_1193 (O_1193,N_24976,N_24526);
nand UO_1194 (O_1194,N_24516,N_24784);
and UO_1195 (O_1195,N_24551,N_24640);
xnor UO_1196 (O_1196,N_24928,N_24736);
xor UO_1197 (O_1197,N_24672,N_24602);
xnor UO_1198 (O_1198,N_24761,N_24995);
and UO_1199 (O_1199,N_24515,N_24774);
xnor UO_1200 (O_1200,N_24524,N_24992);
and UO_1201 (O_1201,N_24730,N_24989);
xor UO_1202 (O_1202,N_24679,N_24857);
nor UO_1203 (O_1203,N_24556,N_24901);
or UO_1204 (O_1204,N_24504,N_24735);
nor UO_1205 (O_1205,N_24550,N_24720);
xnor UO_1206 (O_1206,N_24917,N_24775);
xnor UO_1207 (O_1207,N_24822,N_24977);
nor UO_1208 (O_1208,N_24527,N_24745);
xnor UO_1209 (O_1209,N_24651,N_24644);
and UO_1210 (O_1210,N_24745,N_24647);
or UO_1211 (O_1211,N_24594,N_24974);
and UO_1212 (O_1212,N_24574,N_24737);
xor UO_1213 (O_1213,N_24757,N_24889);
nor UO_1214 (O_1214,N_24899,N_24711);
or UO_1215 (O_1215,N_24591,N_24979);
nand UO_1216 (O_1216,N_24946,N_24505);
nand UO_1217 (O_1217,N_24707,N_24696);
xor UO_1218 (O_1218,N_24938,N_24505);
nor UO_1219 (O_1219,N_24579,N_24572);
xnor UO_1220 (O_1220,N_24805,N_24775);
xnor UO_1221 (O_1221,N_24602,N_24742);
nor UO_1222 (O_1222,N_24960,N_24599);
and UO_1223 (O_1223,N_24644,N_24614);
or UO_1224 (O_1224,N_24738,N_24828);
or UO_1225 (O_1225,N_24845,N_24752);
nor UO_1226 (O_1226,N_24805,N_24933);
nor UO_1227 (O_1227,N_24507,N_24581);
xnor UO_1228 (O_1228,N_24961,N_24694);
and UO_1229 (O_1229,N_24712,N_24722);
nor UO_1230 (O_1230,N_24527,N_24627);
nand UO_1231 (O_1231,N_24530,N_24600);
nor UO_1232 (O_1232,N_24880,N_24732);
nand UO_1233 (O_1233,N_24960,N_24710);
nor UO_1234 (O_1234,N_24886,N_24547);
and UO_1235 (O_1235,N_24851,N_24866);
or UO_1236 (O_1236,N_24690,N_24719);
xor UO_1237 (O_1237,N_24761,N_24837);
xor UO_1238 (O_1238,N_24950,N_24577);
xor UO_1239 (O_1239,N_24592,N_24941);
nand UO_1240 (O_1240,N_24842,N_24608);
and UO_1241 (O_1241,N_24931,N_24735);
nand UO_1242 (O_1242,N_24547,N_24555);
nor UO_1243 (O_1243,N_24822,N_24636);
nor UO_1244 (O_1244,N_24517,N_24726);
xnor UO_1245 (O_1245,N_24865,N_24952);
nand UO_1246 (O_1246,N_24674,N_24715);
nand UO_1247 (O_1247,N_24545,N_24743);
and UO_1248 (O_1248,N_24672,N_24634);
xor UO_1249 (O_1249,N_24552,N_24895);
and UO_1250 (O_1250,N_24529,N_24894);
nand UO_1251 (O_1251,N_24714,N_24506);
xor UO_1252 (O_1252,N_24804,N_24938);
xor UO_1253 (O_1253,N_24921,N_24754);
and UO_1254 (O_1254,N_24782,N_24615);
and UO_1255 (O_1255,N_24694,N_24880);
nand UO_1256 (O_1256,N_24540,N_24677);
nand UO_1257 (O_1257,N_24835,N_24769);
or UO_1258 (O_1258,N_24719,N_24878);
or UO_1259 (O_1259,N_24612,N_24943);
or UO_1260 (O_1260,N_24638,N_24997);
and UO_1261 (O_1261,N_24787,N_24719);
and UO_1262 (O_1262,N_24631,N_24802);
xnor UO_1263 (O_1263,N_24798,N_24911);
nand UO_1264 (O_1264,N_24531,N_24861);
or UO_1265 (O_1265,N_24553,N_24837);
xnor UO_1266 (O_1266,N_24513,N_24925);
nor UO_1267 (O_1267,N_24844,N_24767);
nand UO_1268 (O_1268,N_24517,N_24677);
and UO_1269 (O_1269,N_24718,N_24835);
or UO_1270 (O_1270,N_24961,N_24592);
xnor UO_1271 (O_1271,N_24856,N_24976);
nand UO_1272 (O_1272,N_24922,N_24977);
nand UO_1273 (O_1273,N_24535,N_24875);
and UO_1274 (O_1274,N_24513,N_24555);
or UO_1275 (O_1275,N_24955,N_24900);
or UO_1276 (O_1276,N_24741,N_24877);
or UO_1277 (O_1277,N_24782,N_24509);
xor UO_1278 (O_1278,N_24804,N_24754);
xor UO_1279 (O_1279,N_24767,N_24704);
or UO_1280 (O_1280,N_24587,N_24545);
xnor UO_1281 (O_1281,N_24985,N_24569);
and UO_1282 (O_1282,N_24525,N_24920);
nand UO_1283 (O_1283,N_24754,N_24597);
xor UO_1284 (O_1284,N_24982,N_24709);
xor UO_1285 (O_1285,N_24510,N_24642);
and UO_1286 (O_1286,N_24725,N_24948);
and UO_1287 (O_1287,N_24556,N_24897);
and UO_1288 (O_1288,N_24926,N_24798);
or UO_1289 (O_1289,N_24830,N_24580);
xor UO_1290 (O_1290,N_24510,N_24820);
and UO_1291 (O_1291,N_24704,N_24532);
or UO_1292 (O_1292,N_24798,N_24573);
xnor UO_1293 (O_1293,N_24799,N_24619);
xor UO_1294 (O_1294,N_24554,N_24857);
xor UO_1295 (O_1295,N_24777,N_24647);
nor UO_1296 (O_1296,N_24941,N_24589);
nor UO_1297 (O_1297,N_24609,N_24766);
xnor UO_1298 (O_1298,N_24685,N_24526);
or UO_1299 (O_1299,N_24698,N_24880);
nor UO_1300 (O_1300,N_24546,N_24540);
xor UO_1301 (O_1301,N_24731,N_24826);
and UO_1302 (O_1302,N_24688,N_24723);
nor UO_1303 (O_1303,N_24553,N_24670);
or UO_1304 (O_1304,N_24946,N_24734);
xnor UO_1305 (O_1305,N_24751,N_24669);
or UO_1306 (O_1306,N_24922,N_24917);
nor UO_1307 (O_1307,N_24739,N_24819);
nand UO_1308 (O_1308,N_24549,N_24618);
and UO_1309 (O_1309,N_24777,N_24826);
nor UO_1310 (O_1310,N_24521,N_24628);
nor UO_1311 (O_1311,N_24532,N_24841);
or UO_1312 (O_1312,N_24609,N_24762);
nand UO_1313 (O_1313,N_24529,N_24983);
and UO_1314 (O_1314,N_24965,N_24857);
xnor UO_1315 (O_1315,N_24700,N_24796);
nor UO_1316 (O_1316,N_24736,N_24504);
or UO_1317 (O_1317,N_24718,N_24767);
nand UO_1318 (O_1318,N_24754,N_24571);
nand UO_1319 (O_1319,N_24852,N_24963);
nor UO_1320 (O_1320,N_24719,N_24847);
nand UO_1321 (O_1321,N_24684,N_24946);
xor UO_1322 (O_1322,N_24828,N_24742);
nand UO_1323 (O_1323,N_24574,N_24535);
nor UO_1324 (O_1324,N_24851,N_24566);
or UO_1325 (O_1325,N_24720,N_24806);
nand UO_1326 (O_1326,N_24937,N_24899);
and UO_1327 (O_1327,N_24634,N_24808);
xor UO_1328 (O_1328,N_24773,N_24986);
xor UO_1329 (O_1329,N_24586,N_24781);
and UO_1330 (O_1330,N_24869,N_24908);
nor UO_1331 (O_1331,N_24695,N_24852);
nor UO_1332 (O_1332,N_24779,N_24672);
or UO_1333 (O_1333,N_24646,N_24549);
nand UO_1334 (O_1334,N_24753,N_24672);
nand UO_1335 (O_1335,N_24659,N_24924);
or UO_1336 (O_1336,N_24997,N_24666);
or UO_1337 (O_1337,N_24782,N_24864);
or UO_1338 (O_1338,N_24676,N_24930);
xor UO_1339 (O_1339,N_24773,N_24634);
and UO_1340 (O_1340,N_24622,N_24548);
nor UO_1341 (O_1341,N_24611,N_24736);
xor UO_1342 (O_1342,N_24605,N_24655);
or UO_1343 (O_1343,N_24598,N_24959);
xnor UO_1344 (O_1344,N_24622,N_24566);
and UO_1345 (O_1345,N_24526,N_24648);
nor UO_1346 (O_1346,N_24837,N_24927);
and UO_1347 (O_1347,N_24904,N_24702);
nand UO_1348 (O_1348,N_24534,N_24540);
nor UO_1349 (O_1349,N_24952,N_24790);
xor UO_1350 (O_1350,N_24959,N_24691);
or UO_1351 (O_1351,N_24808,N_24670);
and UO_1352 (O_1352,N_24598,N_24518);
xor UO_1353 (O_1353,N_24511,N_24913);
xor UO_1354 (O_1354,N_24556,N_24691);
xor UO_1355 (O_1355,N_24613,N_24818);
or UO_1356 (O_1356,N_24967,N_24989);
nor UO_1357 (O_1357,N_24529,N_24932);
nor UO_1358 (O_1358,N_24862,N_24814);
or UO_1359 (O_1359,N_24735,N_24694);
and UO_1360 (O_1360,N_24509,N_24873);
and UO_1361 (O_1361,N_24686,N_24917);
xor UO_1362 (O_1362,N_24712,N_24930);
or UO_1363 (O_1363,N_24701,N_24883);
or UO_1364 (O_1364,N_24886,N_24992);
nand UO_1365 (O_1365,N_24926,N_24685);
or UO_1366 (O_1366,N_24734,N_24889);
and UO_1367 (O_1367,N_24560,N_24752);
or UO_1368 (O_1368,N_24979,N_24738);
or UO_1369 (O_1369,N_24905,N_24666);
nand UO_1370 (O_1370,N_24793,N_24731);
nand UO_1371 (O_1371,N_24829,N_24890);
nand UO_1372 (O_1372,N_24834,N_24854);
nand UO_1373 (O_1373,N_24597,N_24860);
and UO_1374 (O_1374,N_24721,N_24847);
nor UO_1375 (O_1375,N_24611,N_24829);
and UO_1376 (O_1376,N_24767,N_24940);
xor UO_1377 (O_1377,N_24732,N_24962);
nor UO_1378 (O_1378,N_24573,N_24654);
xor UO_1379 (O_1379,N_24771,N_24582);
nand UO_1380 (O_1380,N_24901,N_24519);
or UO_1381 (O_1381,N_24808,N_24624);
xor UO_1382 (O_1382,N_24962,N_24737);
nor UO_1383 (O_1383,N_24752,N_24968);
nor UO_1384 (O_1384,N_24805,N_24787);
nand UO_1385 (O_1385,N_24922,N_24569);
or UO_1386 (O_1386,N_24762,N_24565);
and UO_1387 (O_1387,N_24549,N_24985);
xor UO_1388 (O_1388,N_24662,N_24630);
or UO_1389 (O_1389,N_24609,N_24844);
nand UO_1390 (O_1390,N_24597,N_24662);
nor UO_1391 (O_1391,N_24999,N_24677);
xnor UO_1392 (O_1392,N_24617,N_24530);
nand UO_1393 (O_1393,N_24858,N_24652);
nor UO_1394 (O_1394,N_24689,N_24935);
and UO_1395 (O_1395,N_24734,N_24794);
xnor UO_1396 (O_1396,N_24534,N_24585);
nand UO_1397 (O_1397,N_24701,N_24525);
nand UO_1398 (O_1398,N_24953,N_24793);
or UO_1399 (O_1399,N_24939,N_24949);
or UO_1400 (O_1400,N_24825,N_24788);
and UO_1401 (O_1401,N_24718,N_24892);
xor UO_1402 (O_1402,N_24582,N_24834);
or UO_1403 (O_1403,N_24713,N_24856);
xnor UO_1404 (O_1404,N_24556,N_24683);
nand UO_1405 (O_1405,N_24588,N_24583);
xnor UO_1406 (O_1406,N_24993,N_24990);
and UO_1407 (O_1407,N_24727,N_24981);
or UO_1408 (O_1408,N_24678,N_24897);
xnor UO_1409 (O_1409,N_24796,N_24767);
or UO_1410 (O_1410,N_24635,N_24877);
nand UO_1411 (O_1411,N_24684,N_24987);
nor UO_1412 (O_1412,N_24738,N_24592);
nor UO_1413 (O_1413,N_24967,N_24887);
nor UO_1414 (O_1414,N_24794,N_24685);
and UO_1415 (O_1415,N_24549,N_24888);
and UO_1416 (O_1416,N_24884,N_24853);
xnor UO_1417 (O_1417,N_24552,N_24758);
and UO_1418 (O_1418,N_24694,N_24811);
xor UO_1419 (O_1419,N_24972,N_24824);
or UO_1420 (O_1420,N_24520,N_24553);
and UO_1421 (O_1421,N_24689,N_24808);
nand UO_1422 (O_1422,N_24797,N_24809);
xnor UO_1423 (O_1423,N_24863,N_24997);
nand UO_1424 (O_1424,N_24686,N_24568);
and UO_1425 (O_1425,N_24786,N_24583);
and UO_1426 (O_1426,N_24659,N_24715);
and UO_1427 (O_1427,N_24581,N_24805);
nand UO_1428 (O_1428,N_24774,N_24793);
nor UO_1429 (O_1429,N_24998,N_24916);
and UO_1430 (O_1430,N_24539,N_24738);
and UO_1431 (O_1431,N_24841,N_24623);
nand UO_1432 (O_1432,N_24658,N_24975);
nor UO_1433 (O_1433,N_24876,N_24932);
xnor UO_1434 (O_1434,N_24959,N_24854);
xnor UO_1435 (O_1435,N_24617,N_24759);
nor UO_1436 (O_1436,N_24592,N_24630);
nor UO_1437 (O_1437,N_24654,N_24880);
or UO_1438 (O_1438,N_24861,N_24969);
or UO_1439 (O_1439,N_24569,N_24747);
nor UO_1440 (O_1440,N_24505,N_24690);
and UO_1441 (O_1441,N_24731,N_24737);
nand UO_1442 (O_1442,N_24722,N_24843);
and UO_1443 (O_1443,N_24705,N_24572);
and UO_1444 (O_1444,N_24686,N_24667);
or UO_1445 (O_1445,N_24787,N_24800);
or UO_1446 (O_1446,N_24726,N_24615);
nand UO_1447 (O_1447,N_24726,N_24511);
nand UO_1448 (O_1448,N_24551,N_24742);
nand UO_1449 (O_1449,N_24734,N_24910);
nand UO_1450 (O_1450,N_24624,N_24523);
xnor UO_1451 (O_1451,N_24756,N_24760);
xor UO_1452 (O_1452,N_24589,N_24821);
or UO_1453 (O_1453,N_24862,N_24656);
nand UO_1454 (O_1454,N_24611,N_24907);
nand UO_1455 (O_1455,N_24990,N_24909);
or UO_1456 (O_1456,N_24695,N_24771);
nand UO_1457 (O_1457,N_24564,N_24751);
nand UO_1458 (O_1458,N_24627,N_24956);
nand UO_1459 (O_1459,N_24925,N_24966);
nand UO_1460 (O_1460,N_24592,N_24984);
and UO_1461 (O_1461,N_24866,N_24653);
nor UO_1462 (O_1462,N_24927,N_24612);
nor UO_1463 (O_1463,N_24722,N_24896);
nand UO_1464 (O_1464,N_24834,N_24504);
xnor UO_1465 (O_1465,N_24709,N_24611);
nand UO_1466 (O_1466,N_24855,N_24987);
xor UO_1467 (O_1467,N_24779,N_24830);
xnor UO_1468 (O_1468,N_24762,N_24619);
xnor UO_1469 (O_1469,N_24773,N_24747);
xor UO_1470 (O_1470,N_24918,N_24720);
or UO_1471 (O_1471,N_24921,N_24544);
nand UO_1472 (O_1472,N_24841,N_24966);
nand UO_1473 (O_1473,N_24896,N_24633);
nand UO_1474 (O_1474,N_24634,N_24688);
nand UO_1475 (O_1475,N_24594,N_24635);
or UO_1476 (O_1476,N_24822,N_24815);
xnor UO_1477 (O_1477,N_24719,N_24737);
and UO_1478 (O_1478,N_24874,N_24890);
nand UO_1479 (O_1479,N_24951,N_24680);
nand UO_1480 (O_1480,N_24747,N_24643);
and UO_1481 (O_1481,N_24944,N_24602);
xor UO_1482 (O_1482,N_24651,N_24955);
or UO_1483 (O_1483,N_24541,N_24691);
nor UO_1484 (O_1484,N_24522,N_24615);
nand UO_1485 (O_1485,N_24769,N_24901);
and UO_1486 (O_1486,N_24602,N_24631);
and UO_1487 (O_1487,N_24879,N_24749);
or UO_1488 (O_1488,N_24707,N_24976);
xor UO_1489 (O_1489,N_24717,N_24631);
or UO_1490 (O_1490,N_24514,N_24898);
and UO_1491 (O_1491,N_24684,N_24739);
nor UO_1492 (O_1492,N_24873,N_24997);
xor UO_1493 (O_1493,N_24558,N_24813);
or UO_1494 (O_1494,N_24705,N_24968);
xor UO_1495 (O_1495,N_24629,N_24861);
and UO_1496 (O_1496,N_24756,N_24553);
nor UO_1497 (O_1497,N_24577,N_24988);
xor UO_1498 (O_1498,N_24505,N_24943);
xnor UO_1499 (O_1499,N_24987,N_24548);
nor UO_1500 (O_1500,N_24705,N_24784);
xor UO_1501 (O_1501,N_24519,N_24919);
or UO_1502 (O_1502,N_24544,N_24787);
nand UO_1503 (O_1503,N_24916,N_24547);
nor UO_1504 (O_1504,N_24870,N_24698);
xnor UO_1505 (O_1505,N_24523,N_24854);
nand UO_1506 (O_1506,N_24817,N_24570);
or UO_1507 (O_1507,N_24950,N_24505);
nor UO_1508 (O_1508,N_24942,N_24611);
and UO_1509 (O_1509,N_24584,N_24591);
nor UO_1510 (O_1510,N_24851,N_24808);
and UO_1511 (O_1511,N_24915,N_24822);
or UO_1512 (O_1512,N_24908,N_24824);
or UO_1513 (O_1513,N_24707,N_24955);
nor UO_1514 (O_1514,N_24717,N_24711);
nand UO_1515 (O_1515,N_24931,N_24935);
and UO_1516 (O_1516,N_24581,N_24890);
nand UO_1517 (O_1517,N_24630,N_24840);
xnor UO_1518 (O_1518,N_24922,N_24699);
nor UO_1519 (O_1519,N_24929,N_24707);
or UO_1520 (O_1520,N_24964,N_24935);
and UO_1521 (O_1521,N_24506,N_24861);
nand UO_1522 (O_1522,N_24774,N_24966);
nand UO_1523 (O_1523,N_24517,N_24552);
xnor UO_1524 (O_1524,N_24906,N_24775);
nor UO_1525 (O_1525,N_24645,N_24512);
or UO_1526 (O_1526,N_24664,N_24501);
and UO_1527 (O_1527,N_24938,N_24713);
or UO_1528 (O_1528,N_24575,N_24583);
and UO_1529 (O_1529,N_24744,N_24540);
nor UO_1530 (O_1530,N_24529,N_24885);
and UO_1531 (O_1531,N_24842,N_24765);
nor UO_1532 (O_1532,N_24956,N_24910);
and UO_1533 (O_1533,N_24680,N_24639);
nor UO_1534 (O_1534,N_24881,N_24619);
nand UO_1535 (O_1535,N_24675,N_24804);
and UO_1536 (O_1536,N_24727,N_24761);
nand UO_1537 (O_1537,N_24617,N_24923);
nand UO_1538 (O_1538,N_24507,N_24692);
nor UO_1539 (O_1539,N_24821,N_24847);
and UO_1540 (O_1540,N_24897,N_24744);
nand UO_1541 (O_1541,N_24662,N_24804);
nand UO_1542 (O_1542,N_24547,N_24904);
xnor UO_1543 (O_1543,N_24730,N_24772);
or UO_1544 (O_1544,N_24877,N_24887);
and UO_1545 (O_1545,N_24652,N_24904);
nor UO_1546 (O_1546,N_24849,N_24602);
and UO_1547 (O_1547,N_24876,N_24549);
xnor UO_1548 (O_1548,N_24771,N_24872);
and UO_1549 (O_1549,N_24987,N_24638);
and UO_1550 (O_1550,N_24531,N_24856);
nor UO_1551 (O_1551,N_24808,N_24599);
nor UO_1552 (O_1552,N_24941,N_24846);
nor UO_1553 (O_1553,N_24710,N_24908);
nor UO_1554 (O_1554,N_24793,N_24981);
nand UO_1555 (O_1555,N_24888,N_24689);
nand UO_1556 (O_1556,N_24673,N_24831);
nor UO_1557 (O_1557,N_24842,N_24668);
xnor UO_1558 (O_1558,N_24900,N_24972);
nor UO_1559 (O_1559,N_24764,N_24763);
nor UO_1560 (O_1560,N_24552,N_24907);
nor UO_1561 (O_1561,N_24659,N_24602);
nor UO_1562 (O_1562,N_24670,N_24532);
or UO_1563 (O_1563,N_24854,N_24831);
xor UO_1564 (O_1564,N_24834,N_24565);
xor UO_1565 (O_1565,N_24933,N_24708);
xor UO_1566 (O_1566,N_24847,N_24805);
or UO_1567 (O_1567,N_24612,N_24968);
or UO_1568 (O_1568,N_24839,N_24509);
nand UO_1569 (O_1569,N_24667,N_24847);
nor UO_1570 (O_1570,N_24788,N_24855);
xnor UO_1571 (O_1571,N_24878,N_24984);
and UO_1572 (O_1572,N_24898,N_24776);
or UO_1573 (O_1573,N_24533,N_24572);
nor UO_1574 (O_1574,N_24534,N_24563);
or UO_1575 (O_1575,N_24550,N_24578);
and UO_1576 (O_1576,N_24578,N_24535);
xnor UO_1577 (O_1577,N_24858,N_24871);
and UO_1578 (O_1578,N_24521,N_24866);
or UO_1579 (O_1579,N_24500,N_24812);
or UO_1580 (O_1580,N_24547,N_24943);
and UO_1581 (O_1581,N_24605,N_24504);
nor UO_1582 (O_1582,N_24996,N_24757);
or UO_1583 (O_1583,N_24754,N_24933);
or UO_1584 (O_1584,N_24789,N_24626);
or UO_1585 (O_1585,N_24995,N_24781);
nand UO_1586 (O_1586,N_24865,N_24614);
or UO_1587 (O_1587,N_24999,N_24986);
nor UO_1588 (O_1588,N_24791,N_24788);
xor UO_1589 (O_1589,N_24759,N_24509);
and UO_1590 (O_1590,N_24883,N_24501);
nand UO_1591 (O_1591,N_24693,N_24663);
nand UO_1592 (O_1592,N_24833,N_24558);
and UO_1593 (O_1593,N_24788,N_24836);
nand UO_1594 (O_1594,N_24755,N_24542);
and UO_1595 (O_1595,N_24983,N_24702);
xor UO_1596 (O_1596,N_24674,N_24890);
xor UO_1597 (O_1597,N_24632,N_24950);
and UO_1598 (O_1598,N_24549,N_24935);
and UO_1599 (O_1599,N_24899,N_24862);
or UO_1600 (O_1600,N_24990,N_24551);
nor UO_1601 (O_1601,N_24541,N_24756);
nor UO_1602 (O_1602,N_24523,N_24889);
nor UO_1603 (O_1603,N_24787,N_24517);
nor UO_1604 (O_1604,N_24738,N_24845);
or UO_1605 (O_1605,N_24971,N_24748);
or UO_1606 (O_1606,N_24868,N_24866);
or UO_1607 (O_1607,N_24646,N_24703);
nor UO_1608 (O_1608,N_24779,N_24556);
or UO_1609 (O_1609,N_24764,N_24709);
nand UO_1610 (O_1610,N_24804,N_24875);
and UO_1611 (O_1611,N_24790,N_24686);
or UO_1612 (O_1612,N_24517,N_24549);
nand UO_1613 (O_1613,N_24914,N_24753);
and UO_1614 (O_1614,N_24617,N_24542);
xnor UO_1615 (O_1615,N_24878,N_24733);
nand UO_1616 (O_1616,N_24862,N_24638);
nand UO_1617 (O_1617,N_24942,N_24882);
or UO_1618 (O_1618,N_24652,N_24999);
xnor UO_1619 (O_1619,N_24767,N_24609);
and UO_1620 (O_1620,N_24557,N_24847);
nor UO_1621 (O_1621,N_24643,N_24574);
nor UO_1622 (O_1622,N_24877,N_24876);
nor UO_1623 (O_1623,N_24885,N_24810);
nor UO_1624 (O_1624,N_24504,N_24613);
xnor UO_1625 (O_1625,N_24872,N_24565);
or UO_1626 (O_1626,N_24777,N_24999);
nand UO_1627 (O_1627,N_24839,N_24644);
nand UO_1628 (O_1628,N_24668,N_24753);
nor UO_1629 (O_1629,N_24978,N_24659);
or UO_1630 (O_1630,N_24577,N_24757);
and UO_1631 (O_1631,N_24878,N_24597);
and UO_1632 (O_1632,N_24958,N_24664);
and UO_1633 (O_1633,N_24752,N_24772);
or UO_1634 (O_1634,N_24716,N_24924);
or UO_1635 (O_1635,N_24627,N_24941);
or UO_1636 (O_1636,N_24961,N_24969);
nor UO_1637 (O_1637,N_24672,N_24785);
or UO_1638 (O_1638,N_24585,N_24724);
and UO_1639 (O_1639,N_24800,N_24715);
and UO_1640 (O_1640,N_24944,N_24546);
nand UO_1641 (O_1641,N_24828,N_24589);
xor UO_1642 (O_1642,N_24933,N_24800);
nor UO_1643 (O_1643,N_24540,N_24562);
nor UO_1644 (O_1644,N_24978,N_24870);
or UO_1645 (O_1645,N_24619,N_24606);
or UO_1646 (O_1646,N_24880,N_24534);
xnor UO_1647 (O_1647,N_24687,N_24915);
nor UO_1648 (O_1648,N_24898,N_24772);
nor UO_1649 (O_1649,N_24990,N_24668);
nand UO_1650 (O_1650,N_24536,N_24518);
nor UO_1651 (O_1651,N_24969,N_24999);
and UO_1652 (O_1652,N_24805,N_24728);
xnor UO_1653 (O_1653,N_24915,N_24819);
and UO_1654 (O_1654,N_24932,N_24656);
nor UO_1655 (O_1655,N_24575,N_24725);
or UO_1656 (O_1656,N_24548,N_24826);
nor UO_1657 (O_1657,N_24725,N_24632);
or UO_1658 (O_1658,N_24880,N_24961);
nand UO_1659 (O_1659,N_24970,N_24907);
nand UO_1660 (O_1660,N_24730,N_24779);
xnor UO_1661 (O_1661,N_24727,N_24585);
or UO_1662 (O_1662,N_24660,N_24860);
and UO_1663 (O_1663,N_24990,N_24722);
nor UO_1664 (O_1664,N_24784,N_24586);
and UO_1665 (O_1665,N_24530,N_24888);
nor UO_1666 (O_1666,N_24810,N_24572);
or UO_1667 (O_1667,N_24793,N_24662);
and UO_1668 (O_1668,N_24682,N_24652);
nand UO_1669 (O_1669,N_24529,N_24899);
and UO_1670 (O_1670,N_24887,N_24832);
nand UO_1671 (O_1671,N_24656,N_24639);
nand UO_1672 (O_1672,N_24791,N_24765);
and UO_1673 (O_1673,N_24586,N_24975);
and UO_1674 (O_1674,N_24717,N_24895);
xnor UO_1675 (O_1675,N_24516,N_24589);
and UO_1676 (O_1676,N_24928,N_24965);
xor UO_1677 (O_1677,N_24859,N_24551);
nor UO_1678 (O_1678,N_24543,N_24959);
nor UO_1679 (O_1679,N_24961,N_24716);
nor UO_1680 (O_1680,N_24927,N_24561);
or UO_1681 (O_1681,N_24648,N_24511);
nand UO_1682 (O_1682,N_24738,N_24589);
nand UO_1683 (O_1683,N_24833,N_24680);
nand UO_1684 (O_1684,N_24542,N_24869);
or UO_1685 (O_1685,N_24650,N_24640);
nand UO_1686 (O_1686,N_24849,N_24842);
nor UO_1687 (O_1687,N_24857,N_24596);
or UO_1688 (O_1688,N_24796,N_24631);
or UO_1689 (O_1689,N_24852,N_24666);
and UO_1690 (O_1690,N_24666,N_24936);
nand UO_1691 (O_1691,N_24706,N_24896);
nand UO_1692 (O_1692,N_24734,N_24890);
xor UO_1693 (O_1693,N_24672,N_24844);
nand UO_1694 (O_1694,N_24899,N_24835);
xnor UO_1695 (O_1695,N_24858,N_24695);
xor UO_1696 (O_1696,N_24526,N_24752);
nand UO_1697 (O_1697,N_24603,N_24653);
xnor UO_1698 (O_1698,N_24907,N_24950);
and UO_1699 (O_1699,N_24717,N_24841);
nor UO_1700 (O_1700,N_24525,N_24835);
nand UO_1701 (O_1701,N_24610,N_24843);
nand UO_1702 (O_1702,N_24874,N_24905);
or UO_1703 (O_1703,N_24571,N_24878);
and UO_1704 (O_1704,N_24543,N_24850);
nor UO_1705 (O_1705,N_24602,N_24798);
nor UO_1706 (O_1706,N_24532,N_24640);
or UO_1707 (O_1707,N_24872,N_24938);
or UO_1708 (O_1708,N_24982,N_24897);
and UO_1709 (O_1709,N_24525,N_24987);
xnor UO_1710 (O_1710,N_24840,N_24654);
and UO_1711 (O_1711,N_24803,N_24585);
and UO_1712 (O_1712,N_24930,N_24917);
and UO_1713 (O_1713,N_24730,N_24961);
and UO_1714 (O_1714,N_24722,N_24508);
or UO_1715 (O_1715,N_24906,N_24570);
or UO_1716 (O_1716,N_24817,N_24815);
nor UO_1717 (O_1717,N_24742,N_24787);
xnor UO_1718 (O_1718,N_24844,N_24552);
nor UO_1719 (O_1719,N_24996,N_24770);
or UO_1720 (O_1720,N_24751,N_24761);
and UO_1721 (O_1721,N_24919,N_24804);
and UO_1722 (O_1722,N_24870,N_24832);
nand UO_1723 (O_1723,N_24994,N_24768);
xor UO_1724 (O_1724,N_24879,N_24980);
nor UO_1725 (O_1725,N_24804,N_24702);
or UO_1726 (O_1726,N_24523,N_24910);
or UO_1727 (O_1727,N_24793,N_24886);
xnor UO_1728 (O_1728,N_24657,N_24573);
xnor UO_1729 (O_1729,N_24744,N_24697);
or UO_1730 (O_1730,N_24572,N_24715);
or UO_1731 (O_1731,N_24906,N_24855);
nor UO_1732 (O_1732,N_24617,N_24933);
and UO_1733 (O_1733,N_24739,N_24770);
or UO_1734 (O_1734,N_24892,N_24795);
and UO_1735 (O_1735,N_24885,N_24700);
or UO_1736 (O_1736,N_24788,N_24893);
xnor UO_1737 (O_1737,N_24957,N_24918);
and UO_1738 (O_1738,N_24849,N_24987);
nand UO_1739 (O_1739,N_24679,N_24723);
xor UO_1740 (O_1740,N_24520,N_24898);
and UO_1741 (O_1741,N_24529,N_24671);
or UO_1742 (O_1742,N_24957,N_24591);
nand UO_1743 (O_1743,N_24940,N_24873);
or UO_1744 (O_1744,N_24606,N_24639);
and UO_1745 (O_1745,N_24989,N_24923);
nor UO_1746 (O_1746,N_24629,N_24889);
nor UO_1747 (O_1747,N_24838,N_24798);
nand UO_1748 (O_1748,N_24947,N_24527);
xnor UO_1749 (O_1749,N_24664,N_24864);
nand UO_1750 (O_1750,N_24919,N_24732);
xor UO_1751 (O_1751,N_24543,N_24922);
and UO_1752 (O_1752,N_24683,N_24723);
nand UO_1753 (O_1753,N_24886,N_24929);
xnor UO_1754 (O_1754,N_24606,N_24798);
and UO_1755 (O_1755,N_24657,N_24903);
or UO_1756 (O_1756,N_24810,N_24721);
nand UO_1757 (O_1757,N_24659,N_24834);
and UO_1758 (O_1758,N_24629,N_24823);
xnor UO_1759 (O_1759,N_24968,N_24953);
or UO_1760 (O_1760,N_24856,N_24858);
nor UO_1761 (O_1761,N_24700,N_24877);
or UO_1762 (O_1762,N_24872,N_24716);
nand UO_1763 (O_1763,N_24928,N_24523);
and UO_1764 (O_1764,N_24944,N_24881);
or UO_1765 (O_1765,N_24579,N_24589);
nand UO_1766 (O_1766,N_24997,N_24508);
or UO_1767 (O_1767,N_24980,N_24857);
and UO_1768 (O_1768,N_24666,N_24711);
nand UO_1769 (O_1769,N_24677,N_24769);
and UO_1770 (O_1770,N_24965,N_24848);
or UO_1771 (O_1771,N_24875,N_24661);
and UO_1772 (O_1772,N_24790,N_24542);
nand UO_1773 (O_1773,N_24926,N_24731);
or UO_1774 (O_1774,N_24679,N_24770);
or UO_1775 (O_1775,N_24836,N_24964);
nand UO_1776 (O_1776,N_24733,N_24717);
or UO_1777 (O_1777,N_24534,N_24817);
xnor UO_1778 (O_1778,N_24750,N_24555);
nand UO_1779 (O_1779,N_24790,N_24881);
xor UO_1780 (O_1780,N_24813,N_24610);
nor UO_1781 (O_1781,N_24779,N_24729);
nand UO_1782 (O_1782,N_24773,N_24850);
and UO_1783 (O_1783,N_24608,N_24836);
xnor UO_1784 (O_1784,N_24994,N_24864);
xor UO_1785 (O_1785,N_24807,N_24622);
nor UO_1786 (O_1786,N_24842,N_24696);
or UO_1787 (O_1787,N_24810,N_24752);
nor UO_1788 (O_1788,N_24689,N_24583);
nand UO_1789 (O_1789,N_24810,N_24604);
nor UO_1790 (O_1790,N_24986,N_24993);
and UO_1791 (O_1791,N_24933,N_24514);
nand UO_1792 (O_1792,N_24705,N_24722);
nand UO_1793 (O_1793,N_24793,N_24889);
xnor UO_1794 (O_1794,N_24646,N_24627);
or UO_1795 (O_1795,N_24855,N_24509);
nor UO_1796 (O_1796,N_24935,N_24639);
nand UO_1797 (O_1797,N_24898,N_24698);
or UO_1798 (O_1798,N_24995,N_24992);
nor UO_1799 (O_1799,N_24835,N_24559);
nor UO_1800 (O_1800,N_24701,N_24650);
and UO_1801 (O_1801,N_24694,N_24973);
nand UO_1802 (O_1802,N_24564,N_24527);
xor UO_1803 (O_1803,N_24864,N_24631);
or UO_1804 (O_1804,N_24731,N_24974);
nand UO_1805 (O_1805,N_24781,N_24886);
and UO_1806 (O_1806,N_24699,N_24928);
nor UO_1807 (O_1807,N_24977,N_24544);
nand UO_1808 (O_1808,N_24536,N_24710);
and UO_1809 (O_1809,N_24583,N_24896);
xor UO_1810 (O_1810,N_24989,N_24586);
and UO_1811 (O_1811,N_24539,N_24889);
and UO_1812 (O_1812,N_24698,N_24751);
nand UO_1813 (O_1813,N_24513,N_24549);
nor UO_1814 (O_1814,N_24978,N_24555);
and UO_1815 (O_1815,N_24717,N_24747);
or UO_1816 (O_1816,N_24586,N_24621);
nor UO_1817 (O_1817,N_24737,N_24682);
nor UO_1818 (O_1818,N_24632,N_24960);
and UO_1819 (O_1819,N_24718,N_24538);
and UO_1820 (O_1820,N_24768,N_24813);
xor UO_1821 (O_1821,N_24568,N_24646);
nor UO_1822 (O_1822,N_24698,N_24939);
and UO_1823 (O_1823,N_24565,N_24570);
nor UO_1824 (O_1824,N_24636,N_24615);
and UO_1825 (O_1825,N_24588,N_24712);
xnor UO_1826 (O_1826,N_24857,N_24858);
and UO_1827 (O_1827,N_24810,N_24505);
xor UO_1828 (O_1828,N_24821,N_24776);
nand UO_1829 (O_1829,N_24567,N_24502);
xnor UO_1830 (O_1830,N_24605,N_24785);
xnor UO_1831 (O_1831,N_24533,N_24786);
xor UO_1832 (O_1832,N_24770,N_24902);
nor UO_1833 (O_1833,N_24868,N_24925);
nand UO_1834 (O_1834,N_24924,N_24526);
nand UO_1835 (O_1835,N_24615,N_24619);
or UO_1836 (O_1836,N_24582,N_24844);
or UO_1837 (O_1837,N_24913,N_24955);
or UO_1838 (O_1838,N_24841,N_24571);
and UO_1839 (O_1839,N_24633,N_24736);
xnor UO_1840 (O_1840,N_24865,N_24670);
xor UO_1841 (O_1841,N_24744,N_24888);
nand UO_1842 (O_1842,N_24751,N_24987);
nand UO_1843 (O_1843,N_24593,N_24995);
or UO_1844 (O_1844,N_24684,N_24888);
or UO_1845 (O_1845,N_24811,N_24625);
xor UO_1846 (O_1846,N_24709,N_24624);
nand UO_1847 (O_1847,N_24714,N_24896);
nor UO_1848 (O_1848,N_24730,N_24950);
and UO_1849 (O_1849,N_24779,N_24891);
or UO_1850 (O_1850,N_24665,N_24512);
xor UO_1851 (O_1851,N_24936,N_24799);
and UO_1852 (O_1852,N_24575,N_24710);
nand UO_1853 (O_1853,N_24843,N_24906);
nand UO_1854 (O_1854,N_24639,N_24678);
or UO_1855 (O_1855,N_24986,N_24757);
and UO_1856 (O_1856,N_24660,N_24812);
nor UO_1857 (O_1857,N_24863,N_24920);
nand UO_1858 (O_1858,N_24849,N_24941);
and UO_1859 (O_1859,N_24506,N_24782);
or UO_1860 (O_1860,N_24644,N_24587);
or UO_1861 (O_1861,N_24505,N_24606);
xnor UO_1862 (O_1862,N_24556,N_24777);
nand UO_1863 (O_1863,N_24835,N_24727);
or UO_1864 (O_1864,N_24842,N_24596);
xnor UO_1865 (O_1865,N_24830,N_24731);
or UO_1866 (O_1866,N_24772,N_24903);
nor UO_1867 (O_1867,N_24929,N_24538);
and UO_1868 (O_1868,N_24784,N_24950);
nor UO_1869 (O_1869,N_24676,N_24909);
xnor UO_1870 (O_1870,N_24857,N_24789);
nand UO_1871 (O_1871,N_24981,N_24998);
and UO_1872 (O_1872,N_24712,N_24993);
xor UO_1873 (O_1873,N_24620,N_24951);
nand UO_1874 (O_1874,N_24866,N_24977);
xor UO_1875 (O_1875,N_24836,N_24941);
nand UO_1876 (O_1876,N_24821,N_24792);
xor UO_1877 (O_1877,N_24531,N_24685);
nor UO_1878 (O_1878,N_24911,N_24547);
or UO_1879 (O_1879,N_24829,N_24865);
nor UO_1880 (O_1880,N_24655,N_24511);
xor UO_1881 (O_1881,N_24732,N_24718);
xnor UO_1882 (O_1882,N_24887,N_24997);
xnor UO_1883 (O_1883,N_24527,N_24902);
nand UO_1884 (O_1884,N_24824,N_24825);
or UO_1885 (O_1885,N_24731,N_24610);
and UO_1886 (O_1886,N_24531,N_24865);
or UO_1887 (O_1887,N_24750,N_24979);
nand UO_1888 (O_1888,N_24840,N_24682);
nor UO_1889 (O_1889,N_24658,N_24690);
nor UO_1890 (O_1890,N_24532,N_24899);
nor UO_1891 (O_1891,N_24996,N_24574);
nor UO_1892 (O_1892,N_24794,N_24859);
or UO_1893 (O_1893,N_24624,N_24567);
or UO_1894 (O_1894,N_24911,N_24764);
or UO_1895 (O_1895,N_24636,N_24764);
and UO_1896 (O_1896,N_24528,N_24617);
xor UO_1897 (O_1897,N_24768,N_24608);
xnor UO_1898 (O_1898,N_24963,N_24942);
xor UO_1899 (O_1899,N_24842,N_24758);
nor UO_1900 (O_1900,N_24755,N_24572);
nand UO_1901 (O_1901,N_24611,N_24751);
or UO_1902 (O_1902,N_24511,N_24950);
or UO_1903 (O_1903,N_24745,N_24878);
or UO_1904 (O_1904,N_24539,N_24633);
xnor UO_1905 (O_1905,N_24795,N_24807);
or UO_1906 (O_1906,N_24706,N_24821);
nor UO_1907 (O_1907,N_24709,N_24850);
and UO_1908 (O_1908,N_24831,N_24562);
and UO_1909 (O_1909,N_24938,N_24912);
nor UO_1910 (O_1910,N_24852,N_24717);
or UO_1911 (O_1911,N_24907,N_24902);
nor UO_1912 (O_1912,N_24687,N_24607);
xor UO_1913 (O_1913,N_24736,N_24600);
xor UO_1914 (O_1914,N_24659,N_24536);
xnor UO_1915 (O_1915,N_24988,N_24816);
xor UO_1916 (O_1916,N_24850,N_24918);
or UO_1917 (O_1917,N_24525,N_24646);
xnor UO_1918 (O_1918,N_24862,N_24600);
nand UO_1919 (O_1919,N_24805,N_24643);
nor UO_1920 (O_1920,N_24841,N_24775);
nand UO_1921 (O_1921,N_24600,N_24659);
xor UO_1922 (O_1922,N_24598,N_24634);
or UO_1923 (O_1923,N_24955,N_24941);
xor UO_1924 (O_1924,N_24738,N_24827);
or UO_1925 (O_1925,N_24876,N_24639);
or UO_1926 (O_1926,N_24644,N_24547);
nand UO_1927 (O_1927,N_24864,N_24608);
and UO_1928 (O_1928,N_24810,N_24875);
xor UO_1929 (O_1929,N_24606,N_24795);
or UO_1930 (O_1930,N_24808,N_24987);
and UO_1931 (O_1931,N_24688,N_24507);
xor UO_1932 (O_1932,N_24638,N_24876);
and UO_1933 (O_1933,N_24659,N_24930);
or UO_1934 (O_1934,N_24510,N_24852);
nand UO_1935 (O_1935,N_24733,N_24512);
or UO_1936 (O_1936,N_24801,N_24717);
nor UO_1937 (O_1937,N_24735,N_24506);
and UO_1938 (O_1938,N_24931,N_24684);
nand UO_1939 (O_1939,N_24798,N_24717);
nand UO_1940 (O_1940,N_24810,N_24995);
nand UO_1941 (O_1941,N_24834,N_24866);
nor UO_1942 (O_1942,N_24840,N_24597);
xnor UO_1943 (O_1943,N_24677,N_24939);
nand UO_1944 (O_1944,N_24857,N_24711);
xor UO_1945 (O_1945,N_24832,N_24954);
nor UO_1946 (O_1946,N_24689,N_24589);
nor UO_1947 (O_1947,N_24537,N_24730);
and UO_1948 (O_1948,N_24689,N_24648);
and UO_1949 (O_1949,N_24667,N_24539);
nor UO_1950 (O_1950,N_24845,N_24579);
nand UO_1951 (O_1951,N_24586,N_24796);
and UO_1952 (O_1952,N_24635,N_24562);
or UO_1953 (O_1953,N_24852,N_24625);
nor UO_1954 (O_1954,N_24510,N_24712);
and UO_1955 (O_1955,N_24664,N_24727);
or UO_1956 (O_1956,N_24812,N_24737);
and UO_1957 (O_1957,N_24538,N_24772);
xor UO_1958 (O_1958,N_24794,N_24830);
or UO_1959 (O_1959,N_24737,N_24538);
nand UO_1960 (O_1960,N_24691,N_24921);
nand UO_1961 (O_1961,N_24870,N_24699);
or UO_1962 (O_1962,N_24924,N_24685);
nor UO_1963 (O_1963,N_24631,N_24896);
or UO_1964 (O_1964,N_24843,N_24523);
and UO_1965 (O_1965,N_24886,N_24819);
or UO_1966 (O_1966,N_24531,N_24976);
nor UO_1967 (O_1967,N_24574,N_24884);
nand UO_1968 (O_1968,N_24871,N_24795);
xor UO_1969 (O_1969,N_24821,N_24717);
nor UO_1970 (O_1970,N_24959,N_24675);
or UO_1971 (O_1971,N_24957,N_24528);
nor UO_1972 (O_1972,N_24792,N_24971);
and UO_1973 (O_1973,N_24984,N_24730);
nor UO_1974 (O_1974,N_24918,N_24715);
nand UO_1975 (O_1975,N_24525,N_24527);
nor UO_1976 (O_1976,N_24632,N_24880);
nand UO_1977 (O_1977,N_24633,N_24609);
nor UO_1978 (O_1978,N_24992,N_24744);
and UO_1979 (O_1979,N_24947,N_24612);
and UO_1980 (O_1980,N_24936,N_24559);
or UO_1981 (O_1981,N_24649,N_24690);
nor UO_1982 (O_1982,N_24686,N_24605);
and UO_1983 (O_1983,N_24995,N_24551);
nor UO_1984 (O_1984,N_24563,N_24908);
nand UO_1985 (O_1985,N_24941,N_24818);
and UO_1986 (O_1986,N_24788,N_24562);
nor UO_1987 (O_1987,N_24990,N_24843);
nand UO_1988 (O_1988,N_24855,N_24569);
nand UO_1989 (O_1989,N_24907,N_24837);
nor UO_1990 (O_1990,N_24977,N_24734);
xnor UO_1991 (O_1991,N_24940,N_24880);
nor UO_1992 (O_1992,N_24794,N_24674);
and UO_1993 (O_1993,N_24815,N_24832);
or UO_1994 (O_1994,N_24701,N_24907);
xor UO_1995 (O_1995,N_24567,N_24683);
or UO_1996 (O_1996,N_24830,N_24898);
nor UO_1997 (O_1997,N_24894,N_24879);
nand UO_1998 (O_1998,N_24995,N_24918);
nand UO_1999 (O_1999,N_24596,N_24513);
or UO_2000 (O_2000,N_24551,N_24712);
nand UO_2001 (O_2001,N_24696,N_24608);
nor UO_2002 (O_2002,N_24956,N_24618);
nand UO_2003 (O_2003,N_24921,N_24672);
and UO_2004 (O_2004,N_24509,N_24844);
nor UO_2005 (O_2005,N_24560,N_24508);
xnor UO_2006 (O_2006,N_24840,N_24850);
xnor UO_2007 (O_2007,N_24827,N_24875);
or UO_2008 (O_2008,N_24568,N_24632);
and UO_2009 (O_2009,N_24653,N_24820);
nand UO_2010 (O_2010,N_24961,N_24632);
or UO_2011 (O_2011,N_24724,N_24536);
xor UO_2012 (O_2012,N_24520,N_24820);
xor UO_2013 (O_2013,N_24861,N_24878);
nor UO_2014 (O_2014,N_24995,N_24538);
and UO_2015 (O_2015,N_24762,N_24624);
or UO_2016 (O_2016,N_24613,N_24950);
xnor UO_2017 (O_2017,N_24731,N_24979);
and UO_2018 (O_2018,N_24765,N_24531);
or UO_2019 (O_2019,N_24562,N_24865);
or UO_2020 (O_2020,N_24716,N_24828);
and UO_2021 (O_2021,N_24544,N_24742);
and UO_2022 (O_2022,N_24717,N_24517);
or UO_2023 (O_2023,N_24589,N_24600);
or UO_2024 (O_2024,N_24959,N_24742);
xnor UO_2025 (O_2025,N_24722,N_24903);
and UO_2026 (O_2026,N_24519,N_24791);
nand UO_2027 (O_2027,N_24922,N_24606);
or UO_2028 (O_2028,N_24868,N_24666);
nand UO_2029 (O_2029,N_24789,N_24939);
or UO_2030 (O_2030,N_24714,N_24882);
xnor UO_2031 (O_2031,N_24970,N_24935);
nand UO_2032 (O_2032,N_24567,N_24821);
or UO_2033 (O_2033,N_24504,N_24942);
xor UO_2034 (O_2034,N_24941,N_24647);
and UO_2035 (O_2035,N_24768,N_24615);
or UO_2036 (O_2036,N_24541,N_24724);
and UO_2037 (O_2037,N_24544,N_24644);
and UO_2038 (O_2038,N_24632,N_24537);
nand UO_2039 (O_2039,N_24993,N_24922);
xor UO_2040 (O_2040,N_24820,N_24768);
nor UO_2041 (O_2041,N_24757,N_24936);
nand UO_2042 (O_2042,N_24504,N_24597);
nor UO_2043 (O_2043,N_24737,N_24588);
nor UO_2044 (O_2044,N_24618,N_24681);
or UO_2045 (O_2045,N_24921,N_24920);
nor UO_2046 (O_2046,N_24599,N_24973);
or UO_2047 (O_2047,N_24560,N_24688);
or UO_2048 (O_2048,N_24579,N_24784);
xor UO_2049 (O_2049,N_24630,N_24901);
or UO_2050 (O_2050,N_24566,N_24817);
and UO_2051 (O_2051,N_24606,N_24599);
or UO_2052 (O_2052,N_24697,N_24686);
xor UO_2053 (O_2053,N_24968,N_24764);
and UO_2054 (O_2054,N_24906,N_24589);
nand UO_2055 (O_2055,N_24579,N_24737);
nand UO_2056 (O_2056,N_24618,N_24854);
and UO_2057 (O_2057,N_24917,N_24570);
nor UO_2058 (O_2058,N_24955,N_24739);
and UO_2059 (O_2059,N_24871,N_24561);
or UO_2060 (O_2060,N_24580,N_24900);
xnor UO_2061 (O_2061,N_24858,N_24949);
nand UO_2062 (O_2062,N_24549,N_24706);
and UO_2063 (O_2063,N_24626,N_24562);
nand UO_2064 (O_2064,N_24730,N_24670);
xnor UO_2065 (O_2065,N_24708,N_24646);
and UO_2066 (O_2066,N_24839,N_24996);
nor UO_2067 (O_2067,N_24945,N_24944);
and UO_2068 (O_2068,N_24722,N_24639);
and UO_2069 (O_2069,N_24930,N_24947);
xor UO_2070 (O_2070,N_24755,N_24883);
xor UO_2071 (O_2071,N_24558,N_24535);
nor UO_2072 (O_2072,N_24977,N_24998);
nor UO_2073 (O_2073,N_24508,N_24824);
or UO_2074 (O_2074,N_24861,N_24782);
xnor UO_2075 (O_2075,N_24749,N_24790);
nor UO_2076 (O_2076,N_24699,N_24552);
nor UO_2077 (O_2077,N_24629,N_24862);
or UO_2078 (O_2078,N_24936,N_24616);
nand UO_2079 (O_2079,N_24581,N_24670);
nand UO_2080 (O_2080,N_24980,N_24856);
or UO_2081 (O_2081,N_24618,N_24756);
nor UO_2082 (O_2082,N_24812,N_24599);
nand UO_2083 (O_2083,N_24849,N_24565);
nor UO_2084 (O_2084,N_24939,N_24881);
nand UO_2085 (O_2085,N_24696,N_24569);
nor UO_2086 (O_2086,N_24785,N_24714);
or UO_2087 (O_2087,N_24974,N_24665);
xor UO_2088 (O_2088,N_24598,N_24895);
nand UO_2089 (O_2089,N_24762,N_24647);
and UO_2090 (O_2090,N_24781,N_24527);
nand UO_2091 (O_2091,N_24643,N_24521);
nor UO_2092 (O_2092,N_24535,N_24832);
nor UO_2093 (O_2093,N_24998,N_24779);
nor UO_2094 (O_2094,N_24579,N_24724);
nor UO_2095 (O_2095,N_24853,N_24868);
xnor UO_2096 (O_2096,N_24529,N_24956);
nand UO_2097 (O_2097,N_24533,N_24807);
nand UO_2098 (O_2098,N_24630,N_24604);
nor UO_2099 (O_2099,N_24534,N_24661);
or UO_2100 (O_2100,N_24925,N_24597);
xnor UO_2101 (O_2101,N_24528,N_24688);
nor UO_2102 (O_2102,N_24950,N_24913);
nor UO_2103 (O_2103,N_24951,N_24515);
and UO_2104 (O_2104,N_24901,N_24712);
xnor UO_2105 (O_2105,N_24525,N_24593);
or UO_2106 (O_2106,N_24615,N_24548);
xnor UO_2107 (O_2107,N_24950,N_24900);
or UO_2108 (O_2108,N_24988,N_24964);
nand UO_2109 (O_2109,N_24647,N_24575);
xnor UO_2110 (O_2110,N_24964,N_24721);
or UO_2111 (O_2111,N_24619,N_24838);
and UO_2112 (O_2112,N_24579,N_24641);
nor UO_2113 (O_2113,N_24786,N_24925);
xor UO_2114 (O_2114,N_24847,N_24526);
and UO_2115 (O_2115,N_24516,N_24693);
and UO_2116 (O_2116,N_24567,N_24546);
xor UO_2117 (O_2117,N_24624,N_24509);
nand UO_2118 (O_2118,N_24985,N_24966);
or UO_2119 (O_2119,N_24685,N_24575);
xnor UO_2120 (O_2120,N_24904,N_24945);
and UO_2121 (O_2121,N_24607,N_24979);
xnor UO_2122 (O_2122,N_24888,N_24852);
nor UO_2123 (O_2123,N_24747,N_24949);
xor UO_2124 (O_2124,N_24909,N_24681);
xnor UO_2125 (O_2125,N_24937,N_24581);
xor UO_2126 (O_2126,N_24872,N_24777);
nand UO_2127 (O_2127,N_24609,N_24861);
nand UO_2128 (O_2128,N_24643,N_24777);
and UO_2129 (O_2129,N_24559,N_24676);
or UO_2130 (O_2130,N_24927,N_24608);
nor UO_2131 (O_2131,N_24999,N_24595);
and UO_2132 (O_2132,N_24951,N_24818);
xnor UO_2133 (O_2133,N_24879,N_24804);
or UO_2134 (O_2134,N_24878,N_24754);
and UO_2135 (O_2135,N_24975,N_24649);
nand UO_2136 (O_2136,N_24831,N_24511);
nand UO_2137 (O_2137,N_24772,N_24598);
nand UO_2138 (O_2138,N_24950,N_24848);
xnor UO_2139 (O_2139,N_24500,N_24767);
nand UO_2140 (O_2140,N_24638,N_24939);
xor UO_2141 (O_2141,N_24900,N_24681);
nand UO_2142 (O_2142,N_24993,N_24930);
nor UO_2143 (O_2143,N_24593,N_24942);
or UO_2144 (O_2144,N_24856,N_24714);
xnor UO_2145 (O_2145,N_24901,N_24553);
nand UO_2146 (O_2146,N_24998,N_24564);
and UO_2147 (O_2147,N_24666,N_24654);
nand UO_2148 (O_2148,N_24588,N_24549);
and UO_2149 (O_2149,N_24545,N_24702);
xor UO_2150 (O_2150,N_24655,N_24646);
nand UO_2151 (O_2151,N_24778,N_24673);
xor UO_2152 (O_2152,N_24885,N_24832);
nand UO_2153 (O_2153,N_24900,N_24946);
nand UO_2154 (O_2154,N_24921,N_24519);
and UO_2155 (O_2155,N_24802,N_24537);
and UO_2156 (O_2156,N_24729,N_24773);
nand UO_2157 (O_2157,N_24815,N_24876);
and UO_2158 (O_2158,N_24843,N_24841);
and UO_2159 (O_2159,N_24608,N_24884);
nand UO_2160 (O_2160,N_24855,N_24739);
or UO_2161 (O_2161,N_24862,N_24533);
xnor UO_2162 (O_2162,N_24616,N_24566);
or UO_2163 (O_2163,N_24988,N_24649);
nor UO_2164 (O_2164,N_24950,N_24793);
or UO_2165 (O_2165,N_24666,N_24623);
and UO_2166 (O_2166,N_24818,N_24998);
nor UO_2167 (O_2167,N_24805,N_24772);
xor UO_2168 (O_2168,N_24814,N_24925);
nand UO_2169 (O_2169,N_24717,N_24524);
and UO_2170 (O_2170,N_24617,N_24551);
nand UO_2171 (O_2171,N_24714,N_24759);
or UO_2172 (O_2172,N_24770,N_24820);
nor UO_2173 (O_2173,N_24737,N_24985);
and UO_2174 (O_2174,N_24537,N_24690);
and UO_2175 (O_2175,N_24761,N_24563);
xnor UO_2176 (O_2176,N_24862,N_24964);
nand UO_2177 (O_2177,N_24598,N_24809);
or UO_2178 (O_2178,N_24822,N_24972);
nor UO_2179 (O_2179,N_24758,N_24738);
nand UO_2180 (O_2180,N_24880,N_24860);
or UO_2181 (O_2181,N_24823,N_24510);
nor UO_2182 (O_2182,N_24987,N_24554);
nand UO_2183 (O_2183,N_24836,N_24906);
xnor UO_2184 (O_2184,N_24605,N_24847);
nor UO_2185 (O_2185,N_24898,N_24959);
nor UO_2186 (O_2186,N_24672,N_24998);
nand UO_2187 (O_2187,N_24932,N_24921);
and UO_2188 (O_2188,N_24997,N_24996);
nor UO_2189 (O_2189,N_24886,N_24947);
and UO_2190 (O_2190,N_24850,N_24547);
xnor UO_2191 (O_2191,N_24549,N_24827);
xor UO_2192 (O_2192,N_24553,N_24693);
xnor UO_2193 (O_2193,N_24868,N_24775);
xnor UO_2194 (O_2194,N_24637,N_24828);
nand UO_2195 (O_2195,N_24973,N_24531);
and UO_2196 (O_2196,N_24829,N_24889);
nand UO_2197 (O_2197,N_24966,N_24892);
and UO_2198 (O_2198,N_24664,N_24667);
and UO_2199 (O_2199,N_24719,N_24594);
and UO_2200 (O_2200,N_24604,N_24694);
xnor UO_2201 (O_2201,N_24779,N_24763);
and UO_2202 (O_2202,N_24563,N_24792);
xor UO_2203 (O_2203,N_24587,N_24677);
and UO_2204 (O_2204,N_24821,N_24903);
nor UO_2205 (O_2205,N_24793,N_24760);
or UO_2206 (O_2206,N_24754,N_24703);
nand UO_2207 (O_2207,N_24579,N_24533);
xnor UO_2208 (O_2208,N_24695,N_24635);
or UO_2209 (O_2209,N_24750,N_24881);
xnor UO_2210 (O_2210,N_24790,N_24634);
and UO_2211 (O_2211,N_24584,N_24859);
nor UO_2212 (O_2212,N_24572,N_24996);
or UO_2213 (O_2213,N_24570,N_24611);
xor UO_2214 (O_2214,N_24861,N_24786);
and UO_2215 (O_2215,N_24564,N_24755);
nand UO_2216 (O_2216,N_24695,N_24733);
nand UO_2217 (O_2217,N_24569,N_24647);
nand UO_2218 (O_2218,N_24540,N_24618);
or UO_2219 (O_2219,N_24838,N_24695);
nand UO_2220 (O_2220,N_24722,N_24757);
and UO_2221 (O_2221,N_24576,N_24821);
and UO_2222 (O_2222,N_24846,N_24914);
or UO_2223 (O_2223,N_24545,N_24765);
nand UO_2224 (O_2224,N_24952,N_24617);
and UO_2225 (O_2225,N_24572,N_24634);
nor UO_2226 (O_2226,N_24821,N_24725);
and UO_2227 (O_2227,N_24900,N_24963);
xnor UO_2228 (O_2228,N_24541,N_24864);
xor UO_2229 (O_2229,N_24837,N_24855);
or UO_2230 (O_2230,N_24921,N_24956);
and UO_2231 (O_2231,N_24577,N_24824);
or UO_2232 (O_2232,N_24626,N_24913);
or UO_2233 (O_2233,N_24918,N_24855);
xor UO_2234 (O_2234,N_24845,N_24690);
or UO_2235 (O_2235,N_24818,N_24549);
nor UO_2236 (O_2236,N_24919,N_24974);
nand UO_2237 (O_2237,N_24594,N_24562);
and UO_2238 (O_2238,N_24771,N_24939);
or UO_2239 (O_2239,N_24905,N_24642);
nor UO_2240 (O_2240,N_24855,N_24511);
nand UO_2241 (O_2241,N_24727,N_24630);
or UO_2242 (O_2242,N_24869,N_24508);
nand UO_2243 (O_2243,N_24856,N_24764);
and UO_2244 (O_2244,N_24840,N_24795);
or UO_2245 (O_2245,N_24898,N_24941);
xor UO_2246 (O_2246,N_24728,N_24860);
xor UO_2247 (O_2247,N_24657,N_24730);
xor UO_2248 (O_2248,N_24771,N_24878);
nand UO_2249 (O_2249,N_24860,N_24631);
nand UO_2250 (O_2250,N_24722,N_24636);
nor UO_2251 (O_2251,N_24935,N_24914);
nand UO_2252 (O_2252,N_24847,N_24832);
nand UO_2253 (O_2253,N_24926,N_24552);
nor UO_2254 (O_2254,N_24747,N_24783);
xnor UO_2255 (O_2255,N_24602,N_24977);
nor UO_2256 (O_2256,N_24696,N_24604);
or UO_2257 (O_2257,N_24835,N_24760);
xor UO_2258 (O_2258,N_24910,N_24513);
and UO_2259 (O_2259,N_24853,N_24572);
xnor UO_2260 (O_2260,N_24568,N_24868);
and UO_2261 (O_2261,N_24821,N_24935);
and UO_2262 (O_2262,N_24616,N_24535);
xor UO_2263 (O_2263,N_24831,N_24556);
and UO_2264 (O_2264,N_24839,N_24668);
and UO_2265 (O_2265,N_24795,N_24738);
and UO_2266 (O_2266,N_24724,N_24875);
nand UO_2267 (O_2267,N_24699,N_24924);
xnor UO_2268 (O_2268,N_24648,N_24715);
nor UO_2269 (O_2269,N_24681,N_24753);
or UO_2270 (O_2270,N_24949,N_24667);
xor UO_2271 (O_2271,N_24648,N_24664);
nor UO_2272 (O_2272,N_24744,N_24687);
nor UO_2273 (O_2273,N_24922,N_24849);
and UO_2274 (O_2274,N_24828,N_24806);
and UO_2275 (O_2275,N_24783,N_24931);
xor UO_2276 (O_2276,N_24889,N_24769);
xor UO_2277 (O_2277,N_24732,N_24900);
or UO_2278 (O_2278,N_24931,N_24894);
xnor UO_2279 (O_2279,N_24544,N_24788);
xnor UO_2280 (O_2280,N_24705,N_24920);
or UO_2281 (O_2281,N_24615,N_24996);
nand UO_2282 (O_2282,N_24855,N_24785);
or UO_2283 (O_2283,N_24747,N_24805);
nand UO_2284 (O_2284,N_24767,N_24635);
nor UO_2285 (O_2285,N_24868,N_24769);
nor UO_2286 (O_2286,N_24569,N_24594);
xnor UO_2287 (O_2287,N_24760,N_24938);
nand UO_2288 (O_2288,N_24688,N_24573);
xnor UO_2289 (O_2289,N_24895,N_24660);
and UO_2290 (O_2290,N_24664,N_24696);
xnor UO_2291 (O_2291,N_24732,N_24666);
nor UO_2292 (O_2292,N_24948,N_24745);
and UO_2293 (O_2293,N_24618,N_24726);
and UO_2294 (O_2294,N_24985,N_24756);
xor UO_2295 (O_2295,N_24723,N_24514);
and UO_2296 (O_2296,N_24601,N_24861);
or UO_2297 (O_2297,N_24939,N_24653);
nor UO_2298 (O_2298,N_24956,N_24609);
xnor UO_2299 (O_2299,N_24884,N_24804);
nand UO_2300 (O_2300,N_24745,N_24741);
nor UO_2301 (O_2301,N_24561,N_24929);
xnor UO_2302 (O_2302,N_24639,N_24979);
nand UO_2303 (O_2303,N_24994,N_24933);
nor UO_2304 (O_2304,N_24719,N_24609);
nor UO_2305 (O_2305,N_24904,N_24827);
and UO_2306 (O_2306,N_24759,N_24652);
nand UO_2307 (O_2307,N_24742,N_24992);
nand UO_2308 (O_2308,N_24592,N_24875);
or UO_2309 (O_2309,N_24578,N_24606);
xor UO_2310 (O_2310,N_24617,N_24942);
or UO_2311 (O_2311,N_24992,N_24771);
nor UO_2312 (O_2312,N_24704,N_24853);
or UO_2313 (O_2313,N_24811,N_24691);
nor UO_2314 (O_2314,N_24913,N_24696);
xor UO_2315 (O_2315,N_24677,N_24849);
nand UO_2316 (O_2316,N_24871,N_24520);
nand UO_2317 (O_2317,N_24875,N_24871);
or UO_2318 (O_2318,N_24893,N_24705);
nor UO_2319 (O_2319,N_24501,N_24809);
or UO_2320 (O_2320,N_24694,N_24778);
xnor UO_2321 (O_2321,N_24998,N_24621);
xnor UO_2322 (O_2322,N_24802,N_24536);
nor UO_2323 (O_2323,N_24924,N_24985);
and UO_2324 (O_2324,N_24578,N_24791);
xor UO_2325 (O_2325,N_24730,N_24956);
and UO_2326 (O_2326,N_24618,N_24587);
nor UO_2327 (O_2327,N_24878,N_24579);
nor UO_2328 (O_2328,N_24616,N_24652);
or UO_2329 (O_2329,N_24899,N_24665);
nor UO_2330 (O_2330,N_24994,N_24774);
nand UO_2331 (O_2331,N_24891,N_24833);
and UO_2332 (O_2332,N_24925,N_24900);
or UO_2333 (O_2333,N_24640,N_24511);
xor UO_2334 (O_2334,N_24879,N_24939);
xnor UO_2335 (O_2335,N_24619,N_24792);
nand UO_2336 (O_2336,N_24611,N_24592);
nor UO_2337 (O_2337,N_24521,N_24637);
nand UO_2338 (O_2338,N_24589,N_24848);
nor UO_2339 (O_2339,N_24817,N_24637);
or UO_2340 (O_2340,N_24940,N_24699);
xnor UO_2341 (O_2341,N_24981,N_24634);
nand UO_2342 (O_2342,N_24861,N_24953);
or UO_2343 (O_2343,N_24530,N_24575);
nand UO_2344 (O_2344,N_24708,N_24675);
nand UO_2345 (O_2345,N_24838,N_24692);
and UO_2346 (O_2346,N_24918,N_24624);
nand UO_2347 (O_2347,N_24629,N_24938);
and UO_2348 (O_2348,N_24574,N_24995);
xnor UO_2349 (O_2349,N_24835,N_24504);
nand UO_2350 (O_2350,N_24597,N_24586);
nand UO_2351 (O_2351,N_24568,N_24597);
or UO_2352 (O_2352,N_24924,N_24988);
and UO_2353 (O_2353,N_24996,N_24976);
nand UO_2354 (O_2354,N_24504,N_24689);
nor UO_2355 (O_2355,N_24572,N_24856);
nand UO_2356 (O_2356,N_24516,N_24845);
xnor UO_2357 (O_2357,N_24802,N_24696);
xor UO_2358 (O_2358,N_24751,N_24778);
xnor UO_2359 (O_2359,N_24673,N_24711);
and UO_2360 (O_2360,N_24918,N_24785);
or UO_2361 (O_2361,N_24592,N_24739);
nor UO_2362 (O_2362,N_24531,N_24688);
nor UO_2363 (O_2363,N_24532,N_24771);
and UO_2364 (O_2364,N_24981,N_24984);
nor UO_2365 (O_2365,N_24772,N_24955);
nor UO_2366 (O_2366,N_24801,N_24694);
and UO_2367 (O_2367,N_24995,N_24531);
nand UO_2368 (O_2368,N_24910,N_24588);
nand UO_2369 (O_2369,N_24606,N_24837);
and UO_2370 (O_2370,N_24753,N_24501);
xnor UO_2371 (O_2371,N_24538,N_24913);
and UO_2372 (O_2372,N_24719,N_24871);
or UO_2373 (O_2373,N_24569,N_24547);
nor UO_2374 (O_2374,N_24750,N_24894);
nand UO_2375 (O_2375,N_24761,N_24779);
nor UO_2376 (O_2376,N_24909,N_24779);
nand UO_2377 (O_2377,N_24606,N_24570);
nand UO_2378 (O_2378,N_24901,N_24672);
or UO_2379 (O_2379,N_24539,N_24605);
nand UO_2380 (O_2380,N_24824,N_24955);
nor UO_2381 (O_2381,N_24949,N_24828);
and UO_2382 (O_2382,N_24651,N_24980);
nand UO_2383 (O_2383,N_24681,N_24997);
nand UO_2384 (O_2384,N_24623,N_24756);
and UO_2385 (O_2385,N_24790,N_24503);
and UO_2386 (O_2386,N_24621,N_24699);
and UO_2387 (O_2387,N_24765,N_24973);
nor UO_2388 (O_2388,N_24514,N_24610);
nor UO_2389 (O_2389,N_24653,N_24919);
or UO_2390 (O_2390,N_24633,N_24890);
and UO_2391 (O_2391,N_24842,N_24698);
xor UO_2392 (O_2392,N_24746,N_24651);
nor UO_2393 (O_2393,N_24580,N_24996);
xnor UO_2394 (O_2394,N_24921,N_24668);
and UO_2395 (O_2395,N_24716,N_24690);
nor UO_2396 (O_2396,N_24742,N_24706);
or UO_2397 (O_2397,N_24530,N_24591);
and UO_2398 (O_2398,N_24600,N_24940);
nor UO_2399 (O_2399,N_24597,N_24538);
xor UO_2400 (O_2400,N_24747,N_24848);
and UO_2401 (O_2401,N_24502,N_24651);
or UO_2402 (O_2402,N_24974,N_24543);
xnor UO_2403 (O_2403,N_24986,N_24729);
or UO_2404 (O_2404,N_24893,N_24780);
and UO_2405 (O_2405,N_24885,N_24807);
and UO_2406 (O_2406,N_24736,N_24889);
xor UO_2407 (O_2407,N_24588,N_24710);
xnor UO_2408 (O_2408,N_24663,N_24655);
xnor UO_2409 (O_2409,N_24610,N_24798);
or UO_2410 (O_2410,N_24808,N_24986);
nor UO_2411 (O_2411,N_24715,N_24733);
xor UO_2412 (O_2412,N_24652,N_24922);
or UO_2413 (O_2413,N_24772,N_24913);
nand UO_2414 (O_2414,N_24719,N_24641);
or UO_2415 (O_2415,N_24633,N_24906);
nand UO_2416 (O_2416,N_24740,N_24783);
nand UO_2417 (O_2417,N_24844,N_24945);
nand UO_2418 (O_2418,N_24621,N_24632);
nand UO_2419 (O_2419,N_24916,N_24802);
nor UO_2420 (O_2420,N_24882,N_24771);
xor UO_2421 (O_2421,N_24684,N_24659);
nand UO_2422 (O_2422,N_24629,N_24846);
and UO_2423 (O_2423,N_24696,N_24716);
and UO_2424 (O_2424,N_24537,N_24900);
nand UO_2425 (O_2425,N_24656,N_24757);
nor UO_2426 (O_2426,N_24805,N_24845);
nand UO_2427 (O_2427,N_24594,N_24948);
nor UO_2428 (O_2428,N_24854,N_24976);
and UO_2429 (O_2429,N_24594,N_24840);
or UO_2430 (O_2430,N_24913,N_24878);
or UO_2431 (O_2431,N_24686,N_24652);
xnor UO_2432 (O_2432,N_24918,N_24767);
xor UO_2433 (O_2433,N_24962,N_24571);
nand UO_2434 (O_2434,N_24758,N_24500);
or UO_2435 (O_2435,N_24584,N_24963);
nand UO_2436 (O_2436,N_24958,N_24689);
and UO_2437 (O_2437,N_24935,N_24636);
or UO_2438 (O_2438,N_24504,N_24842);
xnor UO_2439 (O_2439,N_24653,N_24895);
nor UO_2440 (O_2440,N_24830,N_24903);
and UO_2441 (O_2441,N_24798,N_24566);
xor UO_2442 (O_2442,N_24559,N_24716);
and UO_2443 (O_2443,N_24504,N_24525);
nand UO_2444 (O_2444,N_24968,N_24667);
xor UO_2445 (O_2445,N_24970,N_24808);
nand UO_2446 (O_2446,N_24665,N_24600);
nor UO_2447 (O_2447,N_24607,N_24540);
or UO_2448 (O_2448,N_24791,N_24736);
or UO_2449 (O_2449,N_24681,N_24565);
xor UO_2450 (O_2450,N_24885,N_24988);
nor UO_2451 (O_2451,N_24688,N_24877);
nor UO_2452 (O_2452,N_24691,N_24536);
and UO_2453 (O_2453,N_24695,N_24823);
or UO_2454 (O_2454,N_24872,N_24680);
nor UO_2455 (O_2455,N_24726,N_24635);
and UO_2456 (O_2456,N_24700,N_24646);
xnor UO_2457 (O_2457,N_24904,N_24978);
or UO_2458 (O_2458,N_24973,N_24925);
nand UO_2459 (O_2459,N_24781,N_24744);
or UO_2460 (O_2460,N_24865,N_24656);
xor UO_2461 (O_2461,N_24669,N_24543);
and UO_2462 (O_2462,N_24580,N_24738);
or UO_2463 (O_2463,N_24728,N_24797);
nand UO_2464 (O_2464,N_24680,N_24732);
nor UO_2465 (O_2465,N_24630,N_24920);
nor UO_2466 (O_2466,N_24754,N_24564);
and UO_2467 (O_2467,N_24673,N_24921);
nor UO_2468 (O_2468,N_24511,N_24734);
or UO_2469 (O_2469,N_24918,N_24562);
nand UO_2470 (O_2470,N_24636,N_24676);
xor UO_2471 (O_2471,N_24721,N_24564);
nand UO_2472 (O_2472,N_24716,N_24779);
xnor UO_2473 (O_2473,N_24549,N_24663);
and UO_2474 (O_2474,N_24791,N_24815);
nand UO_2475 (O_2475,N_24724,N_24618);
nand UO_2476 (O_2476,N_24522,N_24611);
or UO_2477 (O_2477,N_24702,N_24712);
and UO_2478 (O_2478,N_24600,N_24829);
nor UO_2479 (O_2479,N_24593,N_24620);
nand UO_2480 (O_2480,N_24957,N_24559);
and UO_2481 (O_2481,N_24676,N_24690);
nand UO_2482 (O_2482,N_24749,N_24525);
xor UO_2483 (O_2483,N_24544,N_24531);
nand UO_2484 (O_2484,N_24788,N_24531);
nor UO_2485 (O_2485,N_24720,N_24798);
xor UO_2486 (O_2486,N_24791,N_24667);
nor UO_2487 (O_2487,N_24592,N_24952);
nor UO_2488 (O_2488,N_24847,N_24997);
xnor UO_2489 (O_2489,N_24548,N_24913);
xnor UO_2490 (O_2490,N_24821,N_24951);
or UO_2491 (O_2491,N_24576,N_24854);
xor UO_2492 (O_2492,N_24831,N_24600);
or UO_2493 (O_2493,N_24561,N_24584);
nor UO_2494 (O_2494,N_24972,N_24757);
nor UO_2495 (O_2495,N_24686,N_24922);
or UO_2496 (O_2496,N_24549,N_24789);
and UO_2497 (O_2497,N_24650,N_24681);
nand UO_2498 (O_2498,N_24827,N_24562);
or UO_2499 (O_2499,N_24868,N_24918);
nor UO_2500 (O_2500,N_24809,N_24904);
and UO_2501 (O_2501,N_24598,N_24566);
xor UO_2502 (O_2502,N_24606,N_24870);
and UO_2503 (O_2503,N_24800,N_24518);
nor UO_2504 (O_2504,N_24819,N_24564);
nor UO_2505 (O_2505,N_24617,N_24618);
nand UO_2506 (O_2506,N_24800,N_24808);
or UO_2507 (O_2507,N_24663,N_24934);
nor UO_2508 (O_2508,N_24854,N_24652);
or UO_2509 (O_2509,N_24505,N_24749);
nand UO_2510 (O_2510,N_24524,N_24630);
nor UO_2511 (O_2511,N_24952,N_24821);
nor UO_2512 (O_2512,N_24639,N_24609);
xor UO_2513 (O_2513,N_24724,N_24500);
xnor UO_2514 (O_2514,N_24633,N_24874);
xor UO_2515 (O_2515,N_24593,N_24750);
nor UO_2516 (O_2516,N_24715,N_24758);
nand UO_2517 (O_2517,N_24571,N_24540);
and UO_2518 (O_2518,N_24665,N_24588);
nor UO_2519 (O_2519,N_24950,N_24986);
nor UO_2520 (O_2520,N_24704,N_24785);
xor UO_2521 (O_2521,N_24697,N_24700);
and UO_2522 (O_2522,N_24823,N_24755);
or UO_2523 (O_2523,N_24752,N_24850);
and UO_2524 (O_2524,N_24784,N_24625);
nand UO_2525 (O_2525,N_24656,N_24615);
and UO_2526 (O_2526,N_24569,N_24621);
nand UO_2527 (O_2527,N_24757,N_24863);
nand UO_2528 (O_2528,N_24568,N_24662);
or UO_2529 (O_2529,N_24560,N_24816);
xor UO_2530 (O_2530,N_24818,N_24813);
nand UO_2531 (O_2531,N_24741,N_24610);
xor UO_2532 (O_2532,N_24762,N_24787);
nand UO_2533 (O_2533,N_24996,N_24571);
and UO_2534 (O_2534,N_24612,N_24734);
nor UO_2535 (O_2535,N_24556,N_24611);
nor UO_2536 (O_2536,N_24887,N_24514);
nand UO_2537 (O_2537,N_24721,N_24686);
and UO_2538 (O_2538,N_24611,N_24793);
and UO_2539 (O_2539,N_24803,N_24885);
and UO_2540 (O_2540,N_24772,N_24616);
nor UO_2541 (O_2541,N_24643,N_24875);
or UO_2542 (O_2542,N_24779,N_24747);
nand UO_2543 (O_2543,N_24518,N_24822);
nand UO_2544 (O_2544,N_24902,N_24883);
nor UO_2545 (O_2545,N_24707,N_24739);
and UO_2546 (O_2546,N_24536,N_24953);
xnor UO_2547 (O_2547,N_24894,N_24775);
nand UO_2548 (O_2548,N_24884,N_24650);
xnor UO_2549 (O_2549,N_24802,N_24892);
or UO_2550 (O_2550,N_24535,N_24544);
or UO_2551 (O_2551,N_24823,N_24562);
nand UO_2552 (O_2552,N_24769,N_24794);
nor UO_2553 (O_2553,N_24752,N_24863);
or UO_2554 (O_2554,N_24680,N_24637);
nor UO_2555 (O_2555,N_24905,N_24910);
nor UO_2556 (O_2556,N_24928,N_24624);
and UO_2557 (O_2557,N_24743,N_24874);
nand UO_2558 (O_2558,N_24961,N_24966);
and UO_2559 (O_2559,N_24535,N_24715);
or UO_2560 (O_2560,N_24549,N_24500);
xor UO_2561 (O_2561,N_24590,N_24671);
and UO_2562 (O_2562,N_24969,N_24831);
or UO_2563 (O_2563,N_24941,N_24978);
and UO_2564 (O_2564,N_24746,N_24905);
xnor UO_2565 (O_2565,N_24607,N_24807);
and UO_2566 (O_2566,N_24728,N_24522);
and UO_2567 (O_2567,N_24501,N_24592);
nand UO_2568 (O_2568,N_24964,N_24976);
and UO_2569 (O_2569,N_24888,N_24874);
and UO_2570 (O_2570,N_24693,N_24584);
xnor UO_2571 (O_2571,N_24670,N_24891);
nor UO_2572 (O_2572,N_24643,N_24966);
and UO_2573 (O_2573,N_24599,N_24876);
and UO_2574 (O_2574,N_24783,N_24833);
and UO_2575 (O_2575,N_24885,N_24627);
nand UO_2576 (O_2576,N_24596,N_24952);
or UO_2577 (O_2577,N_24962,N_24556);
and UO_2578 (O_2578,N_24889,N_24961);
and UO_2579 (O_2579,N_24511,N_24711);
xnor UO_2580 (O_2580,N_24625,N_24991);
and UO_2581 (O_2581,N_24594,N_24770);
or UO_2582 (O_2582,N_24650,N_24933);
or UO_2583 (O_2583,N_24815,N_24689);
and UO_2584 (O_2584,N_24653,N_24643);
or UO_2585 (O_2585,N_24895,N_24576);
or UO_2586 (O_2586,N_24854,N_24977);
xor UO_2587 (O_2587,N_24879,N_24775);
xor UO_2588 (O_2588,N_24628,N_24838);
nor UO_2589 (O_2589,N_24974,N_24923);
and UO_2590 (O_2590,N_24811,N_24701);
xor UO_2591 (O_2591,N_24827,N_24567);
xnor UO_2592 (O_2592,N_24848,N_24803);
or UO_2593 (O_2593,N_24820,N_24538);
and UO_2594 (O_2594,N_24601,N_24983);
or UO_2595 (O_2595,N_24646,N_24753);
nand UO_2596 (O_2596,N_24668,N_24516);
nor UO_2597 (O_2597,N_24506,N_24615);
nor UO_2598 (O_2598,N_24532,N_24573);
and UO_2599 (O_2599,N_24949,N_24961);
nor UO_2600 (O_2600,N_24907,N_24927);
nand UO_2601 (O_2601,N_24718,N_24605);
nand UO_2602 (O_2602,N_24715,N_24948);
or UO_2603 (O_2603,N_24729,N_24576);
nand UO_2604 (O_2604,N_24767,N_24569);
or UO_2605 (O_2605,N_24578,N_24913);
nor UO_2606 (O_2606,N_24681,N_24920);
and UO_2607 (O_2607,N_24934,N_24803);
or UO_2608 (O_2608,N_24712,N_24726);
or UO_2609 (O_2609,N_24516,N_24873);
or UO_2610 (O_2610,N_24500,N_24508);
or UO_2611 (O_2611,N_24702,N_24923);
xnor UO_2612 (O_2612,N_24723,N_24758);
and UO_2613 (O_2613,N_24656,N_24566);
and UO_2614 (O_2614,N_24793,N_24993);
nand UO_2615 (O_2615,N_24865,N_24998);
or UO_2616 (O_2616,N_24522,N_24960);
nor UO_2617 (O_2617,N_24790,N_24804);
xor UO_2618 (O_2618,N_24707,N_24549);
nor UO_2619 (O_2619,N_24804,N_24827);
and UO_2620 (O_2620,N_24897,N_24870);
nand UO_2621 (O_2621,N_24970,N_24839);
nor UO_2622 (O_2622,N_24988,N_24716);
nor UO_2623 (O_2623,N_24928,N_24588);
nor UO_2624 (O_2624,N_24889,N_24767);
and UO_2625 (O_2625,N_24966,N_24731);
and UO_2626 (O_2626,N_24954,N_24863);
or UO_2627 (O_2627,N_24598,N_24867);
nor UO_2628 (O_2628,N_24503,N_24652);
xnor UO_2629 (O_2629,N_24784,N_24738);
xnor UO_2630 (O_2630,N_24592,N_24979);
nand UO_2631 (O_2631,N_24813,N_24893);
and UO_2632 (O_2632,N_24770,N_24986);
nor UO_2633 (O_2633,N_24568,N_24806);
nand UO_2634 (O_2634,N_24992,N_24555);
and UO_2635 (O_2635,N_24682,N_24746);
nor UO_2636 (O_2636,N_24507,N_24885);
nor UO_2637 (O_2637,N_24786,N_24830);
nand UO_2638 (O_2638,N_24504,N_24881);
or UO_2639 (O_2639,N_24536,N_24793);
xor UO_2640 (O_2640,N_24995,N_24929);
nor UO_2641 (O_2641,N_24563,N_24784);
nand UO_2642 (O_2642,N_24857,N_24951);
or UO_2643 (O_2643,N_24784,N_24897);
or UO_2644 (O_2644,N_24616,N_24866);
or UO_2645 (O_2645,N_24766,N_24692);
nor UO_2646 (O_2646,N_24527,N_24681);
nand UO_2647 (O_2647,N_24594,N_24867);
nor UO_2648 (O_2648,N_24662,N_24895);
and UO_2649 (O_2649,N_24925,N_24828);
nor UO_2650 (O_2650,N_24635,N_24983);
nand UO_2651 (O_2651,N_24978,N_24849);
nand UO_2652 (O_2652,N_24598,N_24731);
xor UO_2653 (O_2653,N_24697,N_24702);
or UO_2654 (O_2654,N_24562,N_24815);
and UO_2655 (O_2655,N_24953,N_24939);
nand UO_2656 (O_2656,N_24820,N_24851);
nand UO_2657 (O_2657,N_24809,N_24603);
nor UO_2658 (O_2658,N_24573,N_24809);
nand UO_2659 (O_2659,N_24586,N_24678);
xnor UO_2660 (O_2660,N_24541,N_24534);
nor UO_2661 (O_2661,N_24577,N_24714);
nand UO_2662 (O_2662,N_24620,N_24597);
nand UO_2663 (O_2663,N_24537,N_24984);
nor UO_2664 (O_2664,N_24562,N_24694);
nand UO_2665 (O_2665,N_24736,N_24840);
xor UO_2666 (O_2666,N_24645,N_24933);
and UO_2667 (O_2667,N_24549,N_24969);
xnor UO_2668 (O_2668,N_24626,N_24541);
xor UO_2669 (O_2669,N_24645,N_24841);
and UO_2670 (O_2670,N_24575,N_24722);
xnor UO_2671 (O_2671,N_24512,N_24805);
xnor UO_2672 (O_2672,N_24981,N_24770);
nor UO_2673 (O_2673,N_24977,N_24630);
or UO_2674 (O_2674,N_24638,N_24883);
nand UO_2675 (O_2675,N_24741,N_24925);
or UO_2676 (O_2676,N_24918,N_24847);
xor UO_2677 (O_2677,N_24871,N_24816);
nand UO_2678 (O_2678,N_24880,N_24962);
or UO_2679 (O_2679,N_24991,N_24760);
xor UO_2680 (O_2680,N_24629,N_24683);
and UO_2681 (O_2681,N_24665,N_24502);
and UO_2682 (O_2682,N_24942,N_24529);
or UO_2683 (O_2683,N_24925,N_24578);
xor UO_2684 (O_2684,N_24903,N_24607);
or UO_2685 (O_2685,N_24579,N_24954);
nand UO_2686 (O_2686,N_24604,N_24990);
and UO_2687 (O_2687,N_24951,N_24614);
and UO_2688 (O_2688,N_24935,N_24999);
nand UO_2689 (O_2689,N_24644,N_24706);
xnor UO_2690 (O_2690,N_24925,N_24818);
xnor UO_2691 (O_2691,N_24778,N_24765);
xnor UO_2692 (O_2692,N_24557,N_24909);
or UO_2693 (O_2693,N_24766,N_24987);
and UO_2694 (O_2694,N_24562,N_24507);
nand UO_2695 (O_2695,N_24797,N_24884);
or UO_2696 (O_2696,N_24703,N_24969);
xnor UO_2697 (O_2697,N_24983,N_24896);
nand UO_2698 (O_2698,N_24551,N_24766);
nor UO_2699 (O_2699,N_24670,N_24727);
nand UO_2700 (O_2700,N_24634,N_24703);
nor UO_2701 (O_2701,N_24959,N_24714);
or UO_2702 (O_2702,N_24818,N_24913);
or UO_2703 (O_2703,N_24700,N_24723);
nor UO_2704 (O_2704,N_24838,N_24539);
and UO_2705 (O_2705,N_24804,N_24930);
and UO_2706 (O_2706,N_24555,N_24526);
nand UO_2707 (O_2707,N_24983,N_24653);
nand UO_2708 (O_2708,N_24821,N_24545);
nand UO_2709 (O_2709,N_24977,N_24646);
or UO_2710 (O_2710,N_24735,N_24980);
xnor UO_2711 (O_2711,N_24693,N_24682);
nand UO_2712 (O_2712,N_24860,N_24707);
xnor UO_2713 (O_2713,N_24712,N_24864);
nand UO_2714 (O_2714,N_24584,N_24562);
nand UO_2715 (O_2715,N_24502,N_24887);
xor UO_2716 (O_2716,N_24814,N_24981);
nand UO_2717 (O_2717,N_24966,N_24671);
nand UO_2718 (O_2718,N_24902,N_24983);
and UO_2719 (O_2719,N_24909,N_24826);
nand UO_2720 (O_2720,N_24640,N_24536);
xor UO_2721 (O_2721,N_24787,N_24727);
nand UO_2722 (O_2722,N_24969,N_24940);
nor UO_2723 (O_2723,N_24741,N_24561);
nor UO_2724 (O_2724,N_24740,N_24898);
nor UO_2725 (O_2725,N_24840,N_24963);
xor UO_2726 (O_2726,N_24557,N_24704);
nand UO_2727 (O_2727,N_24904,N_24980);
nand UO_2728 (O_2728,N_24583,N_24610);
and UO_2729 (O_2729,N_24762,N_24742);
and UO_2730 (O_2730,N_24756,N_24731);
and UO_2731 (O_2731,N_24869,N_24714);
nand UO_2732 (O_2732,N_24688,N_24529);
xor UO_2733 (O_2733,N_24792,N_24709);
and UO_2734 (O_2734,N_24630,N_24693);
or UO_2735 (O_2735,N_24905,N_24682);
xor UO_2736 (O_2736,N_24862,N_24745);
and UO_2737 (O_2737,N_24908,N_24911);
and UO_2738 (O_2738,N_24665,N_24530);
xor UO_2739 (O_2739,N_24894,N_24661);
or UO_2740 (O_2740,N_24937,N_24907);
and UO_2741 (O_2741,N_24832,N_24719);
nor UO_2742 (O_2742,N_24506,N_24652);
nor UO_2743 (O_2743,N_24646,N_24711);
nor UO_2744 (O_2744,N_24649,N_24881);
or UO_2745 (O_2745,N_24549,N_24681);
and UO_2746 (O_2746,N_24855,N_24902);
or UO_2747 (O_2747,N_24524,N_24511);
or UO_2748 (O_2748,N_24848,N_24641);
nand UO_2749 (O_2749,N_24901,N_24921);
and UO_2750 (O_2750,N_24763,N_24772);
and UO_2751 (O_2751,N_24966,N_24621);
nor UO_2752 (O_2752,N_24626,N_24531);
or UO_2753 (O_2753,N_24627,N_24910);
xnor UO_2754 (O_2754,N_24731,N_24647);
or UO_2755 (O_2755,N_24938,N_24520);
or UO_2756 (O_2756,N_24832,N_24656);
nor UO_2757 (O_2757,N_24685,N_24889);
or UO_2758 (O_2758,N_24878,N_24656);
xor UO_2759 (O_2759,N_24861,N_24637);
xnor UO_2760 (O_2760,N_24930,N_24852);
xor UO_2761 (O_2761,N_24865,N_24681);
and UO_2762 (O_2762,N_24607,N_24638);
nand UO_2763 (O_2763,N_24752,N_24503);
and UO_2764 (O_2764,N_24686,N_24920);
xor UO_2765 (O_2765,N_24662,N_24889);
nor UO_2766 (O_2766,N_24847,N_24534);
nor UO_2767 (O_2767,N_24900,N_24574);
or UO_2768 (O_2768,N_24719,N_24696);
or UO_2769 (O_2769,N_24885,N_24600);
or UO_2770 (O_2770,N_24567,N_24920);
and UO_2771 (O_2771,N_24671,N_24974);
nand UO_2772 (O_2772,N_24943,N_24656);
and UO_2773 (O_2773,N_24696,N_24506);
nand UO_2774 (O_2774,N_24979,N_24605);
and UO_2775 (O_2775,N_24832,N_24863);
or UO_2776 (O_2776,N_24500,N_24624);
nand UO_2777 (O_2777,N_24616,N_24778);
or UO_2778 (O_2778,N_24638,N_24683);
xnor UO_2779 (O_2779,N_24836,N_24802);
nor UO_2780 (O_2780,N_24898,N_24986);
xnor UO_2781 (O_2781,N_24722,N_24934);
or UO_2782 (O_2782,N_24753,N_24663);
or UO_2783 (O_2783,N_24665,N_24802);
and UO_2784 (O_2784,N_24769,N_24581);
nand UO_2785 (O_2785,N_24517,N_24504);
or UO_2786 (O_2786,N_24569,N_24912);
xor UO_2787 (O_2787,N_24802,N_24876);
and UO_2788 (O_2788,N_24989,N_24787);
xor UO_2789 (O_2789,N_24889,N_24839);
and UO_2790 (O_2790,N_24910,N_24947);
xor UO_2791 (O_2791,N_24943,N_24850);
nor UO_2792 (O_2792,N_24596,N_24966);
xnor UO_2793 (O_2793,N_24824,N_24840);
nor UO_2794 (O_2794,N_24900,N_24965);
and UO_2795 (O_2795,N_24939,N_24598);
nor UO_2796 (O_2796,N_24932,N_24973);
nand UO_2797 (O_2797,N_24888,N_24681);
nor UO_2798 (O_2798,N_24929,N_24725);
nor UO_2799 (O_2799,N_24724,N_24854);
and UO_2800 (O_2800,N_24880,N_24848);
nor UO_2801 (O_2801,N_24915,N_24831);
or UO_2802 (O_2802,N_24586,N_24961);
xnor UO_2803 (O_2803,N_24939,N_24599);
nand UO_2804 (O_2804,N_24816,N_24516);
or UO_2805 (O_2805,N_24638,N_24934);
or UO_2806 (O_2806,N_24765,N_24508);
nor UO_2807 (O_2807,N_24518,N_24577);
or UO_2808 (O_2808,N_24720,N_24863);
or UO_2809 (O_2809,N_24915,N_24666);
and UO_2810 (O_2810,N_24567,N_24977);
xor UO_2811 (O_2811,N_24707,N_24709);
nor UO_2812 (O_2812,N_24837,N_24684);
nand UO_2813 (O_2813,N_24605,N_24699);
nor UO_2814 (O_2814,N_24860,N_24671);
nand UO_2815 (O_2815,N_24752,N_24800);
nor UO_2816 (O_2816,N_24884,N_24943);
nand UO_2817 (O_2817,N_24564,N_24964);
and UO_2818 (O_2818,N_24844,N_24522);
nor UO_2819 (O_2819,N_24702,N_24662);
or UO_2820 (O_2820,N_24726,N_24599);
or UO_2821 (O_2821,N_24889,N_24927);
and UO_2822 (O_2822,N_24760,N_24540);
nand UO_2823 (O_2823,N_24904,N_24553);
or UO_2824 (O_2824,N_24739,N_24818);
nor UO_2825 (O_2825,N_24805,N_24624);
or UO_2826 (O_2826,N_24936,N_24819);
xnor UO_2827 (O_2827,N_24639,N_24992);
and UO_2828 (O_2828,N_24906,N_24823);
xor UO_2829 (O_2829,N_24819,N_24616);
and UO_2830 (O_2830,N_24588,N_24561);
and UO_2831 (O_2831,N_24909,N_24704);
xnor UO_2832 (O_2832,N_24678,N_24990);
xnor UO_2833 (O_2833,N_24794,N_24645);
nor UO_2834 (O_2834,N_24591,N_24589);
nor UO_2835 (O_2835,N_24603,N_24698);
xor UO_2836 (O_2836,N_24527,N_24996);
xor UO_2837 (O_2837,N_24803,N_24909);
or UO_2838 (O_2838,N_24662,N_24713);
nor UO_2839 (O_2839,N_24531,N_24760);
nand UO_2840 (O_2840,N_24716,N_24665);
or UO_2841 (O_2841,N_24520,N_24550);
or UO_2842 (O_2842,N_24676,N_24788);
and UO_2843 (O_2843,N_24995,N_24874);
nand UO_2844 (O_2844,N_24900,N_24621);
or UO_2845 (O_2845,N_24867,N_24733);
or UO_2846 (O_2846,N_24744,N_24602);
xnor UO_2847 (O_2847,N_24675,N_24727);
nor UO_2848 (O_2848,N_24876,N_24937);
or UO_2849 (O_2849,N_24732,N_24831);
xor UO_2850 (O_2850,N_24667,N_24662);
nor UO_2851 (O_2851,N_24973,N_24965);
nand UO_2852 (O_2852,N_24625,N_24574);
nand UO_2853 (O_2853,N_24853,N_24918);
or UO_2854 (O_2854,N_24653,N_24929);
nand UO_2855 (O_2855,N_24509,N_24962);
nor UO_2856 (O_2856,N_24967,N_24790);
or UO_2857 (O_2857,N_24914,N_24515);
and UO_2858 (O_2858,N_24695,N_24664);
or UO_2859 (O_2859,N_24946,N_24627);
and UO_2860 (O_2860,N_24592,N_24510);
or UO_2861 (O_2861,N_24702,N_24619);
and UO_2862 (O_2862,N_24738,N_24999);
xor UO_2863 (O_2863,N_24829,N_24848);
and UO_2864 (O_2864,N_24935,N_24942);
xor UO_2865 (O_2865,N_24954,N_24870);
xnor UO_2866 (O_2866,N_24814,N_24995);
xnor UO_2867 (O_2867,N_24883,N_24583);
nand UO_2868 (O_2868,N_24704,N_24943);
or UO_2869 (O_2869,N_24865,N_24516);
and UO_2870 (O_2870,N_24752,N_24546);
or UO_2871 (O_2871,N_24846,N_24874);
nand UO_2872 (O_2872,N_24880,N_24647);
or UO_2873 (O_2873,N_24955,N_24850);
nor UO_2874 (O_2874,N_24508,N_24995);
nand UO_2875 (O_2875,N_24640,N_24624);
nor UO_2876 (O_2876,N_24822,N_24721);
nand UO_2877 (O_2877,N_24985,N_24583);
and UO_2878 (O_2878,N_24501,N_24778);
nand UO_2879 (O_2879,N_24798,N_24558);
or UO_2880 (O_2880,N_24862,N_24821);
xnor UO_2881 (O_2881,N_24890,N_24901);
and UO_2882 (O_2882,N_24629,N_24977);
nand UO_2883 (O_2883,N_24564,N_24983);
and UO_2884 (O_2884,N_24541,N_24639);
nand UO_2885 (O_2885,N_24883,N_24554);
nor UO_2886 (O_2886,N_24887,N_24716);
nor UO_2887 (O_2887,N_24555,N_24544);
nand UO_2888 (O_2888,N_24654,N_24581);
or UO_2889 (O_2889,N_24970,N_24567);
nor UO_2890 (O_2890,N_24858,N_24791);
or UO_2891 (O_2891,N_24513,N_24674);
nand UO_2892 (O_2892,N_24625,N_24577);
nand UO_2893 (O_2893,N_24687,N_24769);
or UO_2894 (O_2894,N_24832,N_24813);
and UO_2895 (O_2895,N_24505,N_24740);
nor UO_2896 (O_2896,N_24773,N_24809);
nand UO_2897 (O_2897,N_24545,N_24715);
nor UO_2898 (O_2898,N_24644,N_24564);
and UO_2899 (O_2899,N_24916,N_24987);
nor UO_2900 (O_2900,N_24659,N_24609);
xor UO_2901 (O_2901,N_24968,N_24575);
xnor UO_2902 (O_2902,N_24897,N_24620);
and UO_2903 (O_2903,N_24741,N_24716);
and UO_2904 (O_2904,N_24639,N_24802);
and UO_2905 (O_2905,N_24864,N_24733);
and UO_2906 (O_2906,N_24881,N_24604);
and UO_2907 (O_2907,N_24773,N_24508);
or UO_2908 (O_2908,N_24550,N_24986);
nor UO_2909 (O_2909,N_24876,N_24765);
nand UO_2910 (O_2910,N_24960,N_24655);
xor UO_2911 (O_2911,N_24769,N_24744);
or UO_2912 (O_2912,N_24682,N_24725);
or UO_2913 (O_2913,N_24861,N_24965);
or UO_2914 (O_2914,N_24957,N_24926);
or UO_2915 (O_2915,N_24868,N_24710);
nand UO_2916 (O_2916,N_24676,N_24625);
xor UO_2917 (O_2917,N_24803,N_24586);
xor UO_2918 (O_2918,N_24878,N_24981);
and UO_2919 (O_2919,N_24759,N_24519);
nor UO_2920 (O_2920,N_24813,N_24922);
nor UO_2921 (O_2921,N_24897,N_24747);
xor UO_2922 (O_2922,N_24654,N_24963);
or UO_2923 (O_2923,N_24840,N_24951);
xor UO_2924 (O_2924,N_24663,N_24571);
and UO_2925 (O_2925,N_24614,N_24682);
and UO_2926 (O_2926,N_24547,N_24703);
nor UO_2927 (O_2927,N_24948,N_24984);
nor UO_2928 (O_2928,N_24696,N_24895);
nand UO_2929 (O_2929,N_24950,N_24965);
xnor UO_2930 (O_2930,N_24641,N_24861);
or UO_2931 (O_2931,N_24986,N_24984);
nor UO_2932 (O_2932,N_24555,N_24697);
xnor UO_2933 (O_2933,N_24782,N_24639);
or UO_2934 (O_2934,N_24754,N_24579);
nor UO_2935 (O_2935,N_24740,N_24813);
nor UO_2936 (O_2936,N_24671,N_24777);
and UO_2937 (O_2937,N_24934,N_24608);
nor UO_2938 (O_2938,N_24670,N_24795);
or UO_2939 (O_2939,N_24719,N_24674);
nor UO_2940 (O_2940,N_24678,N_24527);
or UO_2941 (O_2941,N_24972,N_24781);
or UO_2942 (O_2942,N_24652,N_24855);
or UO_2943 (O_2943,N_24801,N_24774);
nand UO_2944 (O_2944,N_24780,N_24501);
or UO_2945 (O_2945,N_24955,N_24677);
or UO_2946 (O_2946,N_24760,N_24810);
nand UO_2947 (O_2947,N_24518,N_24787);
xnor UO_2948 (O_2948,N_24981,N_24657);
and UO_2949 (O_2949,N_24652,N_24721);
or UO_2950 (O_2950,N_24516,N_24876);
and UO_2951 (O_2951,N_24843,N_24575);
xnor UO_2952 (O_2952,N_24704,N_24820);
or UO_2953 (O_2953,N_24899,N_24570);
and UO_2954 (O_2954,N_24975,N_24787);
nor UO_2955 (O_2955,N_24821,N_24942);
and UO_2956 (O_2956,N_24558,N_24789);
and UO_2957 (O_2957,N_24642,N_24620);
or UO_2958 (O_2958,N_24560,N_24742);
nand UO_2959 (O_2959,N_24865,N_24877);
and UO_2960 (O_2960,N_24754,N_24787);
and UO_2961 (O_2961,N_24567,N_24919);
nand UO_2962 (O_2962,N_24692,N_24612);
nand UO_2963 (O_2963,N_24782,N_24686);
nor UO_2964 (O_2964,N_24635,N_24708);
nand UO_2965 (O_2965,N_24644,N_24746);
nor UO_2966 (O_2966,N_24897,N_24625);
nor UO_2967 (O_2967,N_24632,N_24753);
nor UO_2968 (O_2968,N_24851,N_24711);
and UO_2969 (O_2969,N_24612,N_24610);
and UO_2970 (O_2970,N_24755,N_24534);
xnor UO_2971 (O_2971,N_24933,N_24568);
nor UO_2972 (O_2972,N_24595,N_24892);
nor UO_2973 (O_2973,N_24917,N_24727);
nand UO_2974 (O_2974,N_24573,N_24818);
nand UO_2975 (O_2975,N_24975,N_24617);
xor UO_2976 (O_2976,N_24572,N_24782);
and UO_2977 (O_2977,N_24668,N_24902);
nand UO_2978 (O_2978,N_24813,N_24604);
nand UO_2979 (O_2979,N_24557,N_24779);
or UO_2980 (O_2980,N_24573,N_24801);
nand UO_2981 (O_2981,N_24514,N_24592);
or UO_2982 (O_2982,N_24934,N_24502);
nand UO_2983 (O_2983,N_24505,N_24828);
nand UO_2984 (O_2984,N_24993,N_24653);
or UO_2985 (O_2985,N_24792,N_24950);
xnor UO_2986 (O_2986,N_24587,N_24679);
or UO_2987 (O_2987,N_24658,N_24768);
or UO_2988 (O_2988,N_24679,N_24872);
nor UO_2989 (O_2989,N_24576,N_24583);
nand UO_2990 (O_2990,N_24926,N_24670);
xnor UO_2991 (O_2991,N_24570,N_24682);
nor UO_2992 (O_2992,N_24561,N_24565);
or UO_2993 (O_2993,N_24842,N_24810);
and UO_2994 (O_2994,N_24940,N_24686);
xnor UO_2995 (O_2995,N_24593,N_24753);
and UO_2996 (O_2996,N_24581,N_24708);
or UO_2997 (O_2997,N_24755,N_24870);
or UO_2998 (O_2998,N_24973,N_24824);
xor UO_2999 (O_2999,N_24883,N_24742);
endmodule