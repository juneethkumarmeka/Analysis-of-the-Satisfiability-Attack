module basic_1000_10000_1500_10_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
xnor U0 (N_0,In_502,In_152);
nor U1 (N_1,In_325,In_508);
or U2 (N_2,In_206,In_440);
nand U3 (N_3,In_839,In_824);
nor U4 (N_4,In_357,In_285);
nand U5 (N_5,In_434,In_735);
xor U6 (N_6,In_992,In_775);
nor U7 (N_7,In_204,In_500);
nor U8 (N_8,In_111,In_305);
nand U9 (N_9,In_197,In_956);
nor U10 (N_10,In_23,In_6);
nand U11 (N_11,In_699,In_378);
and U12 (N_12,In_898,In_495);
and U13 (N_13,In_39,In_670);
nand U14 (N_14,In_84,In_424);
xnor U15 (N_15,In_104,In_696);
and U16 (N_16,In_350,In_468);
nor U17 (N_17,In_634,In_487);
nand U18 (N_18,In_202,In_90);
nand U19 (N_19,In_109,In_740);
or U20 (N_20,In_118,In_342);
and U21 (N_21,In_368,In_801);
nand U22 (N_22,In_506,In_601);
and U23 (N_23,In_580,In_287);
or U24 (N_24,In_96,In_836);
and U25 (N_25,In_609,In_834);
nor U26 (N_26,In_460,In_29);
and U27 (N_27,In_223,In_681);
or U28 (N_28,In_449,In_192);
nand U29 (N_29,In_522,In_222);
or U30 (N_30,In_174,In_71);
xor U31 (N_31,In_910,In_555);
or U32 (N_32,In_635,In_312);
xnor U33 (N_33,In_383,In_143);
nand U34 (N_34,In_727,In_885);
nor U35 (N_35,In_913,In_893);
nand U36 (N_36,In_139,In_11);
xnor U37 (N_37,In_124,In_878);
and U38 (N_38,In_238,In_266);
xnor U39 (N_39,In_429,In_618);
or U40 (N_40,In_716,In_320);
xnor U41 (N_41,In_796,In_289);
nand U42 (N_42,In_113,In_827);
and U43 (N_43,In_328,In_911);
and U44 (N_44,In_133,In_67);
xor U45 (N_45,In_515,In_20);
or U46 (N_46,In_448,In_486);
nor U47 (N_47,In_229,In_87);
nand U48 (N_48,In_12,In_848);
nand U49 (N_49,In_709,In_822);
xnor U50 (N_50,In_711,In_5);
or U51 (N_51,In_554,In_509);
and U52 (N_52,In_676,In_231);
nand U53 (N_53,In_852,In_311);
or U54 (N_54,In_729,In_776);
nand U55 (N_55,In_470,In_388);
nand U56 (N_56,In_200,In_184);
nand U57 (N_57,In_217,In_54);
xnor U58 (N_58,In_373,In_177);
and U59 (N_59,In_584,In_213);
or U60 (N_60,In_546,In_792);
or U61 (N_61,In_674,In_472);
nor U62 (N_62,In_410,In_921);
nor U63 (N_63,In_928,In_105);
or U64 (N_64,In_561,In_786);
and U65 (N_65,In_948,In_58);
and U66 (N_66,In_163,In_809);
nor U67 (N_67,In_704,In_171);
nor U68 (N_68,In_813,In_541);
nor U69 (N_69,In_220,In_647);
nor U70 (N_70,In_692,In_773);
or U71 (N_71,In_236,In_52);
nand U72 (N_72,In_671,In_563);
nand U73 (N_73,In_95,In_940);
nand U74 (N_74,In_130,In_833);
or U75 (N_75,In_384,In_724);
nor U76 (N_76,In_430,In_151);
xnor U77 (N_77,In_534,In_664);
nand U78 (N_78,In_450,In_596);
nor U79 (N_79,In_247,In_597);
nand U80 (N_80,In_503,In_490);
nor U81 (N_81,In_492,In_234);
nor U82 (N_82,In_544,In_351);
or U83 (N_83,In_10,In_690);
nor U84 (N_84,In_923,In_805);
xnor U85 (N_85,In_94,In_160);
or U86 (N_86,In_625,In_933);
xor U87 (N_87,In_537,In_34);
and U88 (N_88,In_708,In_167);
and U89 (N_89,In_321,In_138);
xnor U90 (N_90,In_760,In_176);
and U91 (N_91,In_154,In_722);
and U92 (N_92,In_372,In_327);
nand U93 (N_93,In_274,In_624);
or U94 (N_94,In_525,In_838);
and U95 (N_95,In_489,In_977);
or U96 (N_96,In_874,In_349);
and U97 (N_97,In_803,In_912);
or U98 (N_98,In_987,In_759);
nor U99 (N_99,In_296,In_396);
or U100 (N_100,In_299,In_628);
and U101 (N_101,In_876,In_966);
nand U102 (N_102,In_499,In_98);
nand U103 (N_103,In_294,In_998);
nand U104 (N_104,In_286,In_248);
xnor U105 (N_105,In_78,In_80);
nor U106 (N_106,In_455,In_538);
xor U107 (N_107,In_386,In_302);
nand U108 (N_108,In_497,In_527);
nor U109 (N_109,In_602,In_25);
xor U110 (N_110,In_929,In_938);
nand U111 (N_111,In_92,In_230);
nor U112 (N_112,In_203,In_245);
xnor U113 (N_113,In_33,In_185);
nor U114 (N_114,In_984,In_445);
and U115 (N_115,In_648,In_412);
and U116 (N_116,In_811,In_605);
nand U117 (N_117,In_968,In_645);
or U118 (N_118,In_369,In_770);
nor U119 (N_119,In_844,In_919);
and U120 (N_120,In_677,In_479);
and U121 (N_121,In_790,In_707);
or U122 (N_122,In_417,In_401);
or U123 (N_123,In_267,In_530);
xnor U124 (N_124,In_24,In_239);
xor U125 (N_125,In_902,In_900);
xor U126 (N_126,In_505,In_744);
and U127 (N_127,In_140,In_436);
nand U128 (N_128,In_57,In_399);
xor U129 (N_129,In_221,In_56);
or U130 (N_130,In_93,In_841);
xor U131 (N_131,In_79,In_753);
and U132 (N_132,In_421,In_346);
nand U133 (N_133,In_157,In_632);
and U134 (N_134,In_849,In_381);
and U135 (N_135,In_661,In_477);
nand U136 (N_136,In_535,In_644);
nand U137 (N_137,In_627,In_443);
nand U138 (N_138,In_757,In_188);
xor U139 (N_139,In_817,In_164);
or U140 (N_140,In_687,In_607);
or U141 (N_141,In_678,In_99);
nand U142 (N_142,In_100,In_411);
nand U143 (N_143,In_53,In_309);
nor U144 (N_144,In_345,In_864);
and U145 (N_145,In_685,In_225);
xor U146 (N_146,In_818,In_300);
nand U147 (N_147,In_387,In_227);
or U148 (N_148,In_832,In_651);
nand U149 (N_149,In_768,In_646);
xor U150 (N_150,In_49,In_592);
xor U151 (N_151,In_623,In_179);
nand U152 (N_152,In_144,In_339);
xnor U153 (N_153,In_533,In_280);
nor U154 (N_154,In_859,In_380);
and U155 (N_155,In_319,In_0);
nand U156 (N_156,In_74,In_715);
xnor U157 (N_157,In_123,In_214);
nand U158 (N_158,In_61,In_719);
nand U159 (N_159,In_442,In_993);
nor U160 (N_160,In_21,In_615);
nand U161 (N_161,In_64,In_804);
and U162 (N_162,In_110,In_51);
or U163 (N_163,In_957,In_665);
xor U164 (N_164,In_301,In_598);
xnor U165 (N_165,In_293,In_662);
nor U166 (N_166,In_918,In_166);
nand U167 (N_167,In_467,In_212);
xor U168 (N_168,In_942,In_720);
and U169 (N_169,In_344,In_954);
and U170 (N_170,In_393,In_684);
and U171 (N_171,In_920,In_193);
nand U172 (N_172,In_959,In_857);
nand U173 (N_173,In_137,In_636);
nor U174 (N_174,In_262,In_173);
or U175 (N_175,In_556,In_19);
nand U176 (N_176,In_103,In_447);
nand U177 (N_177,In_44,In_960);
and U178 (N_178,In_785,In_358);
and U179 (N_179,In_802,In_35);
nor U180 (N_180,In_772,In_643);
xor U181 (N_181,In_807,In_191);
nor U182 (N_182,In_897,In_433);
nor U183 (N_183,In_374,In_997);
and U184 (N_184,In_85,In_691);
and U185 (N_185,In_367,In_738);
and U186 (N_186,In_480,In_867);
xor U187 (N_187,In_149,In_577);
or U188 (N_188,In_30,In_831);
nor U189 (N_189,In_816,In_181);
or U190 (N_190,In_899,In_250);
xor U191 (N_191,In_746,In_553);
xnor U192 (N_192,In_710,In_81);
or U193 (N_193,In_279,In_540);
nand U194 (N_194,In_270,In_228);
nand U195 (N_195,In_806,In_583);
or U196 (N_196,In_531,In_416);
and U197 (N_197,In_117,In_917);
and U198 (N_198,In_516,In_963);
nand U199 (N_199,In_178,In_656);
xor U200 (N_200,In_712,In_941);
nor U201 (N_201,In_481,In_475);
and U202 (N_202,In_879,In_595);
nor U203 (N_203,In_86,In_689);
nand U204 (N_204,In_575,In_400);
nor U205 (N_205,In_43,In_850);
or U206 (N_206,In_253,In_778);
nand U207 (N_207,In_364,In_721);
or U208 (N_208,In_573,In_175);
and U209 (N_209,In_895,In_903);
nor U210 (N_210,In_780,In_557);
or U211 (N_211,In_69,In_937);
and U212 (N_212,In_745,In_265);
or U213 (N_213,In_322,In_18);
nor U214 (N_214,In_638,In_465);
nor U215 (N_215,In_953,In_258);
xor U216 (N_216,In_952,In_565);
and U217 (N_217,In_574,In_697);
xnor U218 (N_218,In_996,In_593);
or U219 (N_219,In_949,In_908);
and U220 (N_220,In_862,In_454);
nor U221 (N_221,In_307,In_600);
or U222 (N_222,In_868,In_518);
and U223 (N_223,In_112,In_855);
nand U224 (N_224,In_965,In_717);
nand U225 (N_225,In_652,In_990);
nand U226 (N_226,In_281,In_980);
xnor U227 (N_227,In_201,In_491);
or U228 (N_228,In_414,In_156);
and U229 (N_229,In_754,In_141);
nor U230 (N_230,In_612,In_385);
and U231 (N_231,In_9,In_298);
and U232 (N_232,In_370,In_962);
xor U233 (N_233,In_675,In_914);
or U234 (N_234,In_389,In_260);
and U235 (N_235,In_283,In_458);
or U236 (N_236,In_331,In_362);
nor U237 (N_237,In_762,In_264);
nand U238 (N_238,In_925,In_734);
and U239 (N_239,In_889,In_865);
xnor U240 (N_240,In_669,In_249);
nand U241 (N_241,In_860,In_316);
nor U242 (N_242,In_31,In_617);
nor U243 (N_243,In_891,In_934);
xor U244 (N_244,In_438,In_730);
or U245 (N_245,In_916,In_91);
nand U246 (N_246,In_484,In_413);
xor U247 (N_247,In_616,In_935);
nand U248 (N_248,In_944,In_861);
and U249 (N_249,In_218,In_254);
nor U250 (N_250,In_457,In_409);
or U251 (N_251,In_115,In_306);
nor U252 (N_252,In_659,In_1);
nand U253 (N_253,In_545,In_750);
nor U254 (N_254,In_579,In_295);
nor U255 (N_255,In_732,In_971);
xor U256 (N_256,In_701,In_27);
or U257 (N_257,In_986,In_453);
xnor U258 (N_258,In_682,In_277);
and U259 (N_259,In_524,In_14);
nor U260 (N_260,In_107,In_189);
and U261 (N_261,In_564,In_927);
and U262 (N_262,In_604,In_382);
and U263 (N_263,In_884,In_359);
nor U264 (N_264,In_145,In_165);
or U265 (N_265,In_147,In_572);
xor U266 (N_266,In_828,In_131);
nand U267 (N_267,In_415,In_748);
xor U268 (N_268,In_931,In_869);
nor U269 (N_269,In_974,In_581);
or U270 (N_270,In_733,In_569);
nor U271 (N_271,In_886,In_106);
nor U272 (N_272,In_257,In_566);
or U273 (N_273,In_32,In_585);
nand U274 (N_274,In_526,In_303);
or U275 (N_275,In_964,In_45);
and U276 (N_276,In_207,In_232);
or U277 (N_277,In_168,In_972);
or U278 (N_278,In_840,In_808);
nor U279 (N_279,In_820,In_683);
or U280 (N_280,In_875,In_698);
xor U281 (N_281,In_469,In_680);
xnor U282 (N_282,In_404,In_586);
nor U283 (N_283,In_788,In_242);
and U284 (N_284,In_854,In_55);
nor U285 (N_285,In_226,In_452);
nor U286 (N_286,In_660,In_501);
nor U287 (N_287,In_706,In_969);
and U288 (N_288,In_407,In_153);
and U289 (N_289,In_883,In_425);
xor U290 (N_290,In_28,In_48);
nand U291 (N_291,In_356,In_282);
nand U292 (N_292,In_4,In_946);
xnor U293 (N_293,In_743,In_766);
and U294 (N_294,In_695,In_126);
nand U295 (N_295,In_473,In_391);
nand U296 (N_296,In_765,In_471);
or U297 (N_297,In_858,In_244);
nand U298 (N_298,In_405,In_62);
xor U299 (N_299,In_507,In_630);
nor U300 (N_300,In_323,In_939);
and U301 (N_301,In_756,In_890);
nor U302 (N_302,In_403,In_552);
nor U303 (N_303,In_985,In_582);
xor U304 (N_304,In_463,In_65);
nand U305 (N_305,In_116,In_485);
or U306 (N_306,In_343,In_406);
or U307 (N_307,In_922,In_132);
nand U308 (N_308,In_190,In_390);
nand U309 (N_309,In_958,In_764);
or U310 (N_310,In_394,In_774);
nor U311 (N_311,In_290,In_975);
and U312 (N_312,In_246,In_863);
xor U313 (N_313,In_633,In_315);
xnor U314 (N_314,In_686,In_983);
or U315 (N_315,In_40,In_700);
xnor U316 (N_316,In_261,In_881);
nor U317 (N_317,In_46,In_650);
nor U318 (N_318,In_208,In_7);
xnor U319 (N_319,In_135,In_233);
nand U320 (N_320,In_134,In_608);
nand U321 (N_321,In_787,In_829);
xor U322 (N_322,In_63,In_16);
nand U323 (N_323,In_512,In_657);
xnor U324 (N_324,In_845,In_637);
and U325 (N_325,In_128,In_375);
nand U326 (N_326,In_119,In_2);
or U327 (N_327,In_894,In_548);
xor U328 (N_328,In_211,In_395);
and U329 (N_329,In_38,In_308);
nor U330 (N_330,In_866,In_13);
or U331 (N_331,In_930,In_210);
or U332 (N_332,In_640,In_631);
or U333 (N_333,In_755,In_483);
xor U334 (N_334,In_613,In_324);
nor U335 (N_335,In_408,In_142);
or U336 (N_336,In_767,In_560);
nor U337 (N_337,In_679,In_310);
nor U338 (N_338,In_620,In_273);
xor U339 (N_339,In_694,In_714);
xnor U340 (N_340,In_906,In_705);
xnor U341 (N_341,In_591,In_498);
or U342 (N_342,In_125,In_550);
and U343 (N_343,In_752,In_422);
and U344 (N_344,In_547,In_37);
or U345 (N_345,In_588,In_418);
nor U346 (N_346,In_170,In_474);
nand U347 (N_347,In_276,In_114);
and U348 (N_348,In_318,In_673);
or U349 (N_349,In_68,In_8);
nor U350 (N_350,In_420,In_590);
xor U351 (N_351,In_314,In_431);
or U352 (N_352,In_194,In_291);
or U353 (N_353,In_549,In_688);
or U354 (N_354,In_991,In_761);
or U355 (N_355,In_519,In_901);
xor U356 (N_356,In_797,In_847);
nand U357 (N_357,In_464,In_379);
and U358 (N_358,In_26,In_663);
or U359 (N_359,In_870,In_363);
xnor U360 (N_360,In_837,In_17);
nor U361 (N_361,In_256,In_317);
or U362 (N_362,In_587,In_146);
nor U363 (N_363,In_955,In_215);
nor U364 (N_364,In_713,In_741);
nor U365 (N_365,In_887,In_880);
xor U366 (N_366,In_819,In_288);
xor U367 (N_367,In_60,In_578);
or U368 (N_368,In_970,In_747);
nor U369 (N_369,In_441,In_195);
and U370 (N_370,In_779,In_313);
and U371 (N_371,In_523,In_932);
and U372 (N_372,In_877,In_159);
and U373 (N_373,In_799,In_108);
xnor U374 (N_374,In_341,In_558);
xor U375 (N_375,In_494,In_89);
xor U376 (N_376,In_329,In_621);
xnor U377 (N_377,In_158,In_205);
xor U378 (N_378,In_798,In_428);
nor U379 (N_379,In_278,In_888);
xor U380 (N_380,In_842,In_334);
or U381 (N_381,In_655,In_493);
nor U382 (N_382,In_186,In_567);
xor U383 (N_383,In_129,In_488);
xnor U384 (N_384,In_476,In_397);
nand U385 (N_385,In_551,In_800);
or U386 (N_386,In_872,In_843);
or U387 (N_387,In_543,In_76);
nand U388 (N_388,In_402,In_703);
or U389 (N_389,In_726,In_513);
nor U390 (N_390,In_326,In_209);
nor U391 (N_391,In_853,In_528);
nand U392 (N_392,In_514,In_529);
nor U393 (N_393,In_482,In_275);
nand U394 (N_394,In_951,In_347);
xor U395 (N_395,In_924,In_243);
xor U396 (N_396,In_994,In_668);
and U397 (N_397,In_943,In_871);
and U398 (N_398,In_196,In_366);
and U399 (N_399,In_36,In_532);
xor U400 (N_400,In_162,In_371);
xnor U401 (N_401,In_999,In_905);
nor U402 (N_402,In_102,In_255);
and U403 (N_403,In_961,In_791);
nor U404 (N_404,In_622,In_172);
xnor U405 (N_405,In_340,In_432);
and U406 (N_406,In_466,In_771);
and U407 (N_407,In_536,In_439);
nor U408 (N_408,In_459,In_169);
nor U409 (N_409,In_610,In_603);
or U410 (N_410,In_693,In_784);
xnor U411 (N_411,In_148,In_121);
xor U412 (N_412,In_520,In_731);
and U413 (N_413,In_224,In_377);
or U414 (N_414,In_702,In_654);
nor U415 (N_415,In_967,In_199);
xnor U416 (N_416,In_161,In_570);
or U417 (N_417,In_97,In_241);
and U418 (N_418,In_562,In_444);
nand U419 (N_419,In_728,In_446);
nand U420 (N_420,In_462,In_376);
xnor U421 (N_421,In_873,In_978);
nor U422 (N_422,In_136,In_435);
nand U423 (N_423,In_672,In_269);
or U424 (N_424,In_988,In_437);
xor U425 (N_425,In_611,In_973);
nand U426 (N_426,In_830,In_47);
or U427 (N_427,In_120,In_263);
or U428 (N_428,In_510,In_777);
nor U429 (N_429,In_271,In_907);
nor U430 (N_430,In_751,In_355);
or U431 (N_431,In_904,In_216);
nor U432 (N_432,In_22,In_235);
xnor U433 (N_433,In_915,In_789);
nand U434 (N_434,In_649,In_348);
or U435 (N_435,In_122,In_268);
xnor U436 (N_436,In_629,In_769);
nor U437 (N_437,In_338,In_252);
nand U438 (N_438,In_653,In_187);
or U439 (N_439,In_180,In_825);
nand U440 (N_440,In_667,In_979);
and U441 (N_441,In_846,In_150);
nand U442 (N_442,In_66,In_3);
or U443 (N_443,In_737,In_423);
nor U444 (N_444,In_511,In_182);
nor U445 (N_445,In_976,In_272);
and U446 (N_446,In_542,In_936);
xor U447 (N_447,In_75,In_82);
nor U448 (N_448,In_101,In_795);
nor U449 (N_449,In_426,In_821);
or U450 (N_450,In_815,In_571);
xor U451 (N_451,In_599,In_183);
nand U452 (N_452,In_398,In_360);
or U453 (N_453,In_723,In_892);
nand U454 (N_454,In_606,In_292);
and U455 (N_455,In_259,In_427);
and U456 (N_456,In_77,In_826);
xnor U457 (N_457,In_337,In_725);
and U458 (N_458,In_794,In_198);
or U459 (N_459,In_83,In_823);
xnor U460 (N_460,In_330,In_219);
or U461 (N_461,In_926,In_718);
or U462 (N_462,In_856,In_361);
or U463 (N_463,In_642,In_461);
xnor U464 (N_464,In_882,In_782);
or U465 (N_465,In_127,In_559);
or U466 (N_466,In_909,In_981);
and U467 (N_467,In_240,In_504);
nor U468 (N_468,In_88,In_50);
nand U469 (N_469,In_521,In_950);
xor U470 (N_470,In_626,In_812);
nor U471 (N_471,In_352,In_666);
and U472 (N_472,In_851,In_658);
nand U473 (N_473,In_781,In_42);
nand U474 (N_474,In_835,In_594);
and U475 (N_475,In_72,In_619);
xnor U476 (N_476,In_284,In_758);
xnor U477 (N_477,In_763,In_451);
nor U478 (N_478,In_392,In_641);
and U479 (N_479,In_810,In_15);
and U480 (N_480,In_736,In_517);
or U481 (N_481,In_783,In_332);
and U482 (N_482,In_70,In_478);
and U483 (N_483,In_742,In_945);
xor U484 (N_484,In_251,In_639);
or U485 (N_485,In_237,In_539);
or U486 (N_486,In_41,In_793);
nor U487 (N_487,In_568,In_896);
nand U488 (N_488,In_335,In_496);
xor U489 (N_489,In_989,In_749);
or U490 (N_490,In_304,In_333);
xnor U491 (N_491,In_995,In_59);
or U492 (N_492,In_947,In_456);
or U493 (N_493,In_365,In_814);
nor U494 (N_494,In_576,In_419);
nand U495 (N_495,In_589,In_614);
or U496 (N_496,In_353,In_336);
and U497 (N_497,In_982,In_739);
nand U498 (N_498,In_297,In_155);
xor U499 (N_499,In_354,In_73);
or U500 (N_500,In_525,In_708);
nand U501 (N_501,In_533,In_205);
nand U502 (N_502,In_946,In_326);
xor U503 (N_503,In_309,In_76);
nor U504 (N_504,In_950,In_54);
nor U505 (N_505,In_24,In_523);
nand U506 (N_506,In_421,In_120);
and U507 (N_507,In_906,In_372);
and U508 (N_508,In_461,In_995);
xor U509 (N_509,In_231,In_667);
nand U510 (N_510,In_352,In_803);
or U511 (N_511,In_105,In_519);
nand U512 (N_512,In_876,In_592);
xor U513 (N_513,In_805,In_835);
and U514 (N_514,In_251,In_984);
xor U515 (N_515,In_167,In_920);
nand U516 (N_516,In_541,In_692);
and U517 (N_517,In_58,In_993);
or U518 (N_518,In_112,In_766);
nor U519 (N_519,In_512,In_248);
and U520 (N_520,In_344,In_735);
nor U521 (N_521,In_344,In_978);
and U522 (N_522,In_709,In_677);
or U523 (N_523,In_67,In_644);
nand U524 (N_524,In_295,In_898);
xor U525 (N_525,In_661,In_140);
and U526 (N_526,In_706,In_471);
xnor U527 (N_527,In_342,In_616);
nor U528 (N_528,In_994,In_106);
and U529 (N_529,In_667,In_682);
xor U530 (N_530,In_979,In_85);
nand U531 (N_531,In_563,In_689);
xor U532 (N_532,In_631,In_350);
and U533 (N_533,In_600,In_785);
xnor U534 (N_534,In_810,In_581);
xnor U535 (N_535,In_545,In_282);
and U536 (N_536,In_623,In_894);
nand U537 (N_537,In_991,In_526);
nand U538 (N_538,In_605,In_449);
nor U539 (N_539,In_577,In_660);
or U540 (N_540,In_712,In_36);
and U541 (N_541,In_989,In_661);
or U542 (N_542,In_479,In_426);
nor U543 (N_543,In_381,In_855);
or U544 (N_544,In_494,In_722);
xnor U545 (N_545,In_997,In_991);
and U546 (N_546,In_192,In_573);
and U547 (N_547,In_169,In_406);
nand U548 (N_548,In_879,In_309);
and U549 (N_549,In_766,In_213);
xor U550 (N_550,In_975,In_160);
nor U551 (N_551,In_563,In_838);
nor U552 (N_552,In_940,In_46);
xor U553 (N_553,In_257,In_518);
or U554 (N_554,In_46,In_686);
and U555 (N_555,In_829,In_201);
and U556 (N_556,In_465,In_239);
nand U557 (N_557,In_947,In_540);
nor U558 (N_558,In_75,In_323);
or U559 (N_559,In_921,In_445);
nand U560 (N_560,In_186,In_865);
nor U561 (N_561,In_939,In_369);
nand U562 (N_562,In_384,In_292);
or U563 (N_563,In_933,In_179);
and U564 (N_564,In_475,In_173);
xnor U565 (N_565,In_287,In_707);
and U566 (N_566,In_758,In_840);
or U567 (N_567,In_131,In_794);
nor U568 (N_568,In_326,In_180);
nand U569 (N_569,In_345,In_876);
or U570 (N_570,In_565,In_782);
or U571 (N_571,In_845,In_512);
and U572 (N_572,In_104,In_389);
or U573 (N_573,In_405,In_973);
and U574 (N_574,In_449,In_328);
and U575 (N_575,In_803,In_705);
nor U576 (N_576,In_394,In_775);
xnor U577 (N_577,In_349,In_634);
xor U578 (N_578,In_540,In_125);
xor U579 (N_579,In_811,In_352);
xnor U580 (N_580,In_327,In_354);
nand U581 (N_581,In_896,In_86);
nor U582 (N_582,In_140,In_535);
xor U583 (N_583,In_213,In_225);
xor U584 (N_584,In_304,In_374);
nand U585 (N_585,In_682,In_352);
nor U586 (N_586,In_652,In_829);
nor U587 (N_587,In_676,In_531);
or U588 (N_588,In_402,In_840);
and U589 (N_589,In_944,In_466);
nor U590 (N_590,In_761,In_49);
nor U591 (N_591,In_654,In_503);
xor U592 (N_592,In_336,In_53);
and U593 (N_593,In_646,In_722);
xor U594 (N_594,In_955,In_536);
nor U595 (N_595,In_850,In_303);
nor U596 (N_596,In_914,In_275);
nand U597 (N_597,In_228,In_258);
and U598 (N_598,In_915,In_124);
nor U599 (N_599,In_641,In_47);
xor U600 (N_600,In_100,In_154);
nor U601 (N_601,In_159,In_145);
nand U602 (N_602,In_874,In_312);
or U603 (N_603,In_950,In_132);
nor U604 (N_604,In_180,In_999);
nand U605 (N_605,In_219,In_773);
or U606 (N_606,In_646,In_346);
and U607 (N_607,In_23,In_596);
nor U608 (N_608,In_424,In_159);
and U609 (N_609,In_829,In_456);
and U610 (N_610,In_969,In_995);
nor U611 (N_611,In_814,In_16);
or U612 (N_612,In_535,In_488);
and U613 (N_613,In_308,In_598);
nand U614 (N_614,In_566,In_689);
and U615 (N_615,In_251,In_894);
or U616 (N_616,In_382,In_126);
or U617 (N_617,In_907,In_273);
or U618 (N_618,In_159,In_901);
nand U619 (N_619,In_318,In_937);
xnor U620 (N_620,In_7,In_849);
or U621 (N_621,In_270,In_358);
and U622 (N_622,In_0,In_847);
nand U623 (N_623,In_734,In_997);
and U624 (N_624,In_899,In_207);
xnor U625 (N_625,In_706,In_259);
nand U626 (N_626,In_538,In_570);
or U627 (N_627,In_333,In_557);
and U628 (N_628,In_425,In_918);
and U629 (N_629,In_357,In_892);
nand U630 (N_630,In_633,In_946);
or U631 (N_631,In_114,In_210);
xor U632 (N_632,In_435,In_203);
nand U633 (N_633,In_557,In_45);
nand U634 (N_634,In_247,In_747);
xnor U635 (N_635,In_534,In_820);
xor U636 (N_636,In_368,In_231);
nor U637 (N_637,In_390,In_660);
and U638 (N_638,In_114,In_121);
xnor U639 (N_639,In_127,In_890);
xor U640 (N_640,In_120,In_11);
nand U641 (N_641,In_366,In_348);
nand U642 (N_642,In_520,In_213);
or U643 (N_643,In_42,In_944);
and U644 (N_644,In_230,In_344);
and U645 (N_645,In_876,In_539);
or U646 (N_646,In_537,In_604);
and U647 (N_647,In_160,In_959);
or U648 (N_648,In_559,In_876);
or U649 (N_649,In_181,In_876);
nand U650 (N_650,In_440,In_787);
and U651 (N_651,In_286,In_970);
and U652 (N_652,In_983,In_742);
xnor U653 (N_653,In_948,In_403);
xnor U654 (N_654,In_11,In_521);
or U655 (N_655,In_288,In_766);
nor U656 (N_656,In_299,In_681);
nand U657 (N_657,In_865,In_917);
and U658 (N_658,In_277,In_817);
xor U659 (N_659,In_490,In_304);
and U660 (N_660,In_492,In_403);
xor U661 (N_661,In_927,In_733);
nand U662 (N_662,In_342,In_921);
nor U663 (N_663,In_599,In_963);
xnor U664 (N_664,In_963,In_21);
xor U665 (N_665,In_67,In_989);
xnor U666 (N_666,In_113,In_675);
nand U667 (N_667,In_437,In_506);
or U668 (N_668,In_740,In_785);
nand U669 (N_669,In_149,In_583);
nand U670 (N_670,In_390,In_666);
and U671 (N_671,In_940,In_715);
and U672 (N_672,In_807,In_769);
nand U673 (N_673,In_449,In_647);
or U674 (N_674,In_354,In_41);
or U675 (N_675,In_205,In_841);
nor U676 (N_676,In_891,In_959);
or U677 (N_677,In_576,In_325);
nor U678 (N_678,In_523,In_680);
nor U679 (N_679,In_832,In_886);
or U680 (N_680,In_327,In_454);
and U681 (N_681,In_589,In_221);
or U682 (N_682,In_605,In_568);
and U683 (N_683,In_729,In_972);
xnor U684 (N_684,In_857,In_615);
and U685 (N_685,In_745,In_222);
nor U686 (N_686,In_122,In_92);
and U687 (N_687,In_416,In_480);
xnor U688 (N_688,In_245,In_567);
nand U689 (N_689,In_788,In_99);
nor U690 (N_690,In_426,In_263);
nor U691 (N_691,In_395,In_975);
nand U692 (N_692,In_448,In_788);
nor U693 (N_693,In_368,In_46);
nand U694 (N_694,In_878,In_650);
nand U695 (N_695,In_820,In_656);
nand U696 (N_696,In_3,In_34);
nand U697 (N_697,In_616,In_165);
xnor U698 (N_698,In_60,In_751);
and U699 (N_699,In_344,In_654);
or U700 (N_700,In_799,In_81);
xnor U701 (N_701,In_300,In_60);
xor U702 (N_702,In_271,In_253);
and U703 (N_703,In_445,In_204);
and U704 (N_704,In_738,In_739);
xor U705 (N_705,In_274,In_118);
nor U706 (N_706,In_871,In_274);
nand U707 (N_707,In_299,In_613);
nor U708 (N_708,In_683,In_110);
or U709 (N_709,In_93,In_11);
nand U710 (N_710,In_515,In_397);
nand U711 (N_711,In_71,In_790);
and U712 (N_712,In_980,In_847);
and U713 (N_713,In_60,In_123);
xnor U714 (N_714,In_529,In_528);
or U715 (N_715,In_774,In_616);
xor U716 (N_716,In_283,In_54);
xnor U717 (N_717,In_706,In_501);
or U718 (N_718,In_544,In_642);
and U719 (N_719,In_323,In_203);
nand U720 (N_720,In_344,In_938);
xor U721 (N_721,In_53,In_117);
nor U722 (N_722,In_360,In_97);
nand U723 (N_723,In_994,In_985);
nand U724 (N_724,In_831,In_171);
nor U725 (N_725,In_145,In_517);
or U726 (N_726,In_857,In_403);
nor U727 (N_727,In_625,In_243);
xnor U728 (N_728,In_306,In_190);
nand U729 (N_729,In_365,In_869);
and U730 (N_730,In_804,In_987);
and U731 (N_731,In_246,In_173);
or U732 (N_732,In_275,In_678);
or U733 (N_733,In_544,In_199);
or U734 (N_734,In_292,In_420);
or U735 (N_735,In_173,In_331);
xnor U736 (N_736,In_397,In_51);
nand U737 (N_737,In_19,In_84);
nand U738 (N_738,In_343,In_746);
xor U739 (N_739,In_368,In_110);
and U740 (N_740,In_208,In_888);
or U741 (N_741,In_212,In_953);
nor U742 (N_742,In_629,In_960);
xor U743 (N_743,In_319,In_118);
nor U744 (N_744,In_971,In_404);
xnor U745 (N_745,In_308,In_663);
nor U746 (N_746,In_202,In_649);
xnor U747 (N_747,In_648,In_690);
or U748 (N_748,In_880,In_240);
xor U749 (N_749,In_798,In_100);
nor U750 (N_750,In_112,In_590);
xor U751 (N_751,In_768,In_541);
nor U752 (N_752,In_876,In_487);
nand U753 (N_753,In_163,In_587);
nand U754 (N_754,In_954,In_256);
nand U755 (N_755,In_407,In_279);
or U756 (N_756,In_467,In_38);
or U757 (N_757,In_111,In_657);
nand U758 (N_758,In_761,In_9);
nand U759 (N_759,In_839,In_610);
or U760 (N_760,In_532,In_291);
xnor U761 (N_761,In_467,In_749);
xor U762 (N_762,In_639,In_424);
or U763 (N_763,In_961,In_99);
and U764 (N_764,In_314,In_604);
and U765 (N_765,In_874,In_889);
nor U766 (N_766,In_695,In_775);
xor U767 (N_767,In_421,In_98);
nor U768 (N_768,In_446,In_729);
xor U769 (N_769,In_579,In_831);
and U770 (N_770,In_169,In_323);
and U771 (N_771,In_486,In_810);
or U772 (N_772,In_750,In_938);
or U773 (N_773,In_117,In_677);
nand U774 (N_774,In_879,In_329);
and U775 (N_775,In_902,In_388);
nand U776 (N_776,In_1,In_730);
nor U777 (N_777,In_551,In_110);
nor U778 (N_778,In_209,In_152);
and U779 (N_779,In_735,In_763);
nand U780 (N_780,In_477,In_776);
nor U781 (N_781,In_502,In_874);
nor U782 (N_782,In_895,In_680);
or U783 (N_783,In_691,In_140);
or U784 (N_784,In_924,In_167);
or U785 (N_785,In_545,In_710);
and U786 (N_786,In_803,In_684);
or U787 (N_787,In_865,In_715);
xor U788 (N_788,In_679,In_613);
or U789 (N_789,In_587,In_551);
nor U790 (N_790,In_544,In_630);
nand U791 (N_791,In_776,In_210);
nor U792 (N_792,In_786,In_961);
xor U793 (N_793,In_319,In_145);
xnor U794 (N_794,In_157,In_549);
nor U795 (N_795,In_700,In_709);
and U796 (N_796,In_744,In_710);
and U797 (N_797,In_632,In_298);
nor U798 (N_798,In_800,In_192);
nand U799 (N_799,In_548,In_74);
and U800 (N_800,In_370,In_808);
nor U801 (N_801,In_862,In_450);
nor U802 (N_802,In_53,In_115);
nor U803 (N_803,In_177,In_278);
and U804 (N_804,In_249,In_931);
and U805 (N_805,In_265,In_891);
or U806 (N_806,In_770,In_787);
nor U807 (N_807,In_42,In_320);
or U808 (N_808,In_29,In_608);
nand U809 (N_809,In_42,In_355);
or U810 (N_810,In_511,In_691);
or U811 (N_811,In_972,In_418);
nor U812 (N_812,In_443,In_388);
and U813 (N_813,In_788,In_163);
nand U814 (N_814,In_775,In_169);
or U815 (N_815,In_621,In_438);
xor U816 (N_816,In_122,In_322);
and U817 (N_817,In_937,In_640);
and U818 (N_818,In_198,In_531);
nand U819 (N_819,In_457,In_581);
or U820 (N_820,In_877,In_152);
nor U821 (N_821,In_640,In_831);
xnor U822 (N_822,In_474,In_248);
xnor U823 (N_823,In_125,In_982);
or U824 (N_824,In_713,In_633);
nor U825 (N_825,In_766,In_325);
xor U826 (N_826,In_484,In_268);
or U827 (N_827,In_349,In_514);
xnor U828 (N_828,In_460,In_964);
and U829 (N_829,In_127,In_117);
or U830 (N_830,In_23,In_545);
nor U831 (N_831,In_900,In_435);
or U832 (N_832,In_592,In_879);
or U833 (N_833,In_96,In_926);
and U834 (N_834,In_553,In_632);
nor U835 (N_835,In_186,In_970);
nor U836 (N_836,In_319,In_521);
and U837 (N_837,In_229,In_499);
xor U838 (N_838,In_413,In_595);
or U839 (N_839,In_835,In_762);
and U840 (N_840,In_572,In_217);
xnor U841 (N_841,In_168,In_83);
or U842 (N_842,In_953,In_490);
nor U843 (N_843,In_522,In_363);
xor U844 (N_844,In_722,In_446);
nand U845 (N_845,In_368,In_929);
or U846 (N_846,In_992,In_811);
or U847 (N_847,In_144,In_970);
nand U848 (N_848,In_686,In_241);
xnor U849 (N_849,In_917,In_672);
or U850 (N_850,In_517,In_714);
nand U851 (N_851,In_379,In_791);
nand U852 (N_852,In_709,In_637);
nand U853 (N_853,In_692,In_174);
or U854 (N_854,In_635,In_249);
and U855 (N_855,In_717,In_972);
or U856 (N_856,In_339,In_44);
nand U857 (N_857,In_602,In_178);
xnor U858 (N_858,In_511,In_898);
and U859 (N_859,In_151,In_504);
and U860 (N_860,In_758,In_527);
nand U861 (N_861,In_532,In_846);
nand U862 (N_862,In_302,In_811);
or U863 (N_863,In_91,In_935);
nand U864 (N_864,In_877,In_200);
xnor U865 (N_865,In_395,In_807);
and U866 (N_866,In_102,In_56);
and U867 (N_867,In_977,In_372);
nand U868 (N_868,In_632,In_631);
xor U869 (N_869,In_146,In_169);
xnor U870 (N_870,In_975,In_712);
or U871 (N_871,In_991,In_330);
and U872 (N_872,In_190,In_206);
nand U873 (N_873,In_818,In_972);
or U874 (N_874,In_875,In_337);
nand U875 (N_875,In_236,In_622);
nand U876 (N_876,In_748,In_570);
xor U877 (N_877,In_546,In_833);
nand U878 (N_878,In_955,In_592);
nand U879 (N_879,In_937,In_23);
or U880 (N_880,In_263,In_683);
or U881 (N_881,In_876,In_228);
nand U882 (N_882,In_264,In_103);
and U883 (N_883,In_697,In_893);
nand U884 (N_884,In_616,In_981);
nand U885 (N_885,In_917,In_317);
and U886 (N_886,In_722,In_802);
nor U887 (N_887,In_977,In_798);
nand U888 (N_888,In_183,In_469);
nand U889 (N_889,In_831,In_938);
and U890 (N_890,In_132,In_942);
nand U891 (N_891,In_878,In_652);
and U892 (N_892,In_596,In_178);
xor U893 (N_893,In_537,In_845);
nor U894 (N_894,In_107,In_62);
and U895 (N_895,In_169,In_490);
nor U896 (N_896,In_193,In_956);
and U897 (N_897,In_982,In_664);
nor U898 (N_898,In_228,In_801);
nand U899 (N_899,In_887,In_632);
and U900 (N_900,In_618,In_760);
nor U901 (N_901,In_210,In_350);
nand U902 (N_902,In_81,In_166);
or U903 (N_903,In_204,In_386);
and U904 (N_904,In_827,In_127);
and U905 (N_905,In_51,In_470);
nand U906 (N_906,In_33,In_416);
xor U907 (N_907,In_902,In_986);
xor U908 (N_908,In_17,In_782);
and U909 (N_909,In_78,In_648);
xnor U910 (N_910,In_187,In_733);
and U911 (N_911,In_10,In_205);
nand U912 (N_912,In_379,In_863);
xnor U913 (N_913,In_323,In_266);
or U914 (N_914,In_673,In_107);
and U915 (N_915,In_183,In_767);
nand U916 (N_916,In_232,In_692);
and U917 (N_917,In_112,In_44);
nor U918 (N_918,In_744,In_898);
xnor U919 (N_919,In_94,In_857);
or U920 (N_920,In_80,In_21);
nor U921 (N_921,In_712,In_16);
or U922 (N_922,In_689,In_46);
nor U923 (N_923,In_760,In_824);
and U924 (N_924,In_745,In_623);
nor U925 (N_925,In_857,In_68);
or U926 (N_926,In_138,In_955);
or U927 (N_927,In_27,In_549);
or U928 (N_928,In_4,In_59);
and U929 (N_929,In_243,In_576);
or U930 (N_930,In_803,In_469);
xor U931 (N_931,In_515,In_171);
nor U932 (N_932,In_614,In_224);
and U933 (N_933,In_84,In_856);
nand U934 (N_934,In_142,In_544);
or U935 (N_935,In_659,In_125);
nand U936 (N_936,In_833,In_289);
and U937 (N_937,In_167,In_815);
nand U938 (N_938,In_75,In_456);
nand U939 (N_939,In_898,In_958);
nor U940 (N_940,In_335,In_798);
and U941 (N_941,In_421,In_614);
nand U942 (N_942,In_224,In_604);
nor U943 (N_943,In_649,In_692);
or U944 (N_944,In_719,In_505);
xor U945 (N_945,In_516,In_314);
nand U946 (N_946,In_943,In_352);
xnor U947 (N_947,In_706,In_251);
and U948 (N_948,In_307,In_506);
xnor U949 (N_949,In_980,In_942);
nand U950 (N_950,In_524,In_55);
nand U951 (N_951,In_293,In_600);
nor U952 (N_952,In_84,In_215);
and U953 (N_953,In_199,In_757);
nor U954 (N_954,In_793,In_8);
and U955 (N_955,In_70,In_744);
xnor U956 (N_956,In_409,In_177);
and U957 (N_957,In_650,In_979);
nand U958 (N_958,In_268,In_976);
and U959 (N_959,In_498,In_631);
nor U960 (N_960,In_719,In_818);
nand U961 (N_961,In_416,In_311);
and U962 (N_962,In_36,In_576);
or U963 (N_963,In_429,In_323);
and U964 (N_964,In_868,In_841);
and U965 (N_965,In_556,In_314);
xor U966 (N_966,In_564,In_667);
or U967 (N_967,In_488,In_536);
xnor U968 (N_968,In_853,In_358);
xnor U969 (N_969,In_107,In_369);
xnor U970 (N_970,In_52,In_133);
xor U971 (N_971,In_878,In_572);
xor U972 (N_972,In_608,In_562);
nand U973 (N_973,In_490,In_256);
nand U974 (N_974,In_86,In_484);
nor U975 (N_975,In_601,In_732);
nand U976 (N_976,In_12,In_959);
xor U977 (N_977,In_55,In_122);
xnor U978 (N_978,In_993,In_335);
xor U979 (N_979,In_1,In_333);
and U980 (N_980,In_907,In_567);
or U981 (N_981,In_212,In_140);
and U982 (N_982,In_716,In_502);
nor U983 (N_983,In_627,In_634);
and U984 (N_984,In_202,In_612);
and U985 (N_985,In_292,In_184);
xor U986 (N_986,In_36,In_221);
xor U987 (N_987,In_623,In_106);
or U988 (N_988,In_831,In_336);
and U989 (N_989,In_519,In_882);
and U990 (N_990,In_976,In_628);
or U991 (N_991,In_185,In_855);
or U992 (N_992,In_605,In_104);
xor U993 (N_993,In_265,In_18);
xnor U994 (N_994,In_2,In_292);
nor U995 (N_995,In_726,In_326);
nor U996 (N_996,In_105,In_245);
nor U997 (N_997,In_803,In_492);
nor U998 (N_998,In_931,In_935);
xor U999 (N_999,In_551,In_266);
and U1000 (N_1000,N_614,N_647);
or U1001 (N_1001,N_923,N_936);
nand U1002 (N_1002,N_15,N_251);
or U1003 (N_1003,N_120,N_9);
xor U1004 (N_1004,N_659,N_868);
and U1005 (N_1005,N_947,N_856);
xor U1006 (N_1006,N_830,N_842);
and U1007 (N_1007,N_416,N_701);
xnor U1008 (N_1008,N_841,N_152);
nor U1009 (N_1009,N_697,N_446);
xor U1010 (N_1010,N_543,N_845);
nor U1011 (N_1011,N_121,N_21);
nor U1012 (N_1012,N_79,N_784);
nand U1013 (N_1013,N_698,N_816);
xor U1014 (N_1014,N_849,N_450);
or U1015 (N_1015,N_768,N_459);
xnor U1016 (N_1016,N_866,N_872);
nor U1017 (N_1017,N_430,N_186);
and U1018 (N_1018,N_387,N_775);
xnor U1019 (N_1019,N_809,N_794);
nand U1020 (N_1020,N_798,N_192);
and U1021 (N_1021,N_577,N_759);
xor U1022 (N_1022,N_435,N_392);
nor U1023 (N_1023,N_293,N_709);
or U1024 (N_1024,N_945,N_238);
nor U1025 (N_1025,N_632,N_780);
or U1026 (N_1026,N_68,N_307);
nand U1027 (N_1027,N_425,N_541);
xor U1028 (N_1028,N_937,N_593);
nand U1029 (N_1029,N_276,N_189);
xnor U1030 (N_1030,N_523,N_566);
and U1031 (N_1031,N_822,N_742);
xor U1032 (N_1032,N_438,N_175);
or U1033 (N_1033,N_404,N_542);
xor U1034 (N_1034,N_448,N_288);
xor U1035 (N_1035,N_454,N_990);
and U1036 (N_1036,N_88,N_20);
or U1037 (N_1037,N_887,N_801);
nand U1038 (N_1038,N_820,N_624);
and U1039 (N_1039,N_789,N_442);
nand U1040 (N_1040,N_8,N_386);
nor U1041 (N_1041,N_876,N_568);
and U1042 (N_1042,N_907,N_229);
xor U1043 (N_1043,N_117,N_639);
or U1044 (N_1044,N_359,N_787);
nor U1045 (N_1045,N_244,N_802);
nor U1046 (N_1046,N_729,N_908);
or U1047 (N_1047,N_146,N_714);
or U1048 (N_1048,N_751,N_839);
and U1049 (N_1049,N_656,N_417);
and U1050 (N_1050,N_153,N_981);
and U1051 (N_1051,N_38,N_418);
or U1052 (N_1052,N_264,N_389);
xnor U1053 (N_1053,N_89,N_920);
and U1054 (N_1054,N_69,N_185);
nand U1055 (N_1055,N_808,N_865);
or U1056 (N_1056,N_473,N_154);
nand U1057 (N_1057,N_444,N_852);
nand U1058 (N_1058,N_375,N_504);
nor U1059 (N_1059,N_556,N_319);
and U1060 (N_1060,N_664,N_427);
xor U1061 (N_1061,N_327,N_573);
nor U1062 (N_1062,N_525,N_447);
or U1063 (N_1063,N_661,N_467);
nor U1064 (N_1064,N_901,N_226);
nand U1065 (N_1065,N_772,N_626);
nand U1066 (N_1066,N_518,N_61);
or U1067 (N_1067,N_341,N_619);
xor U1068 (N_1068,N_259,N_892);
and U1069 (N_1069,N_900,N_562);
nand U1070 (N_1070,N_674,N_301);
nor U1071 (N_1071,N_403,N_95);
xnor U1072 (N_1072,N_660,N_917);
and U1073 (N_1073,N_815,N_893);
or U1074 (N_1074,N_456,N_198);
or U1075 (N_1075,N_972,N_196);
and U1076 (N_1076,N_671,N_851);
and U1077 (N_1077,N_648,N_123);
nand U1078 (N_1078,N_883,N_17);
nand U1079 (N_1079,N_247,N_401);
nor U1080 (N_1080,N_296,N_678);
nor U1081 (N_1081,N_212,N_685);
nand U1082 (N_1082,N_505,N_126);
or U1083 (N_1083,N_576,N_382);
or U1084 (N_1084,N_623,N_788);
nand U1085 (N_1085,N_457,N_135);
nor U1086 (N_1086,N_93,N_383);
or U1087 (N_1087,N_724,N_493);
nor U1088 (N_1088,N_30,N_928);
nor U1089 (N_1089,N_687,N_326);
nand U1090 (N_1090,N_155,N_33);
and U1091 (N_1091,N_988,N_168);
or U1092 (N_1092,N_80,N_517);
xnor U1093 (N_1093,N_708,N_285);
nand U1094 (N_1094,N_220,N_646);
nor U1095 (N_1095,N_743,N_354);
nor U1096 (N_1096,N_421,N_76);
nor U1097 (N_1097,N_846,N_799);
or U1098 (N_1098,N_333,N_254);
or U1099 (N_1099,N_863,N_510);
xnor U1100 (N_1100,N_462,N_796);
or U1101 (N_1101,N_358,N_591);
and U1102 (N_1102,N_635,N_443);
xor U1103 (N_1103,N_987,N_282);
or U1104 (N_1104,N_162,N_311);
and U1105 (N_1105,N_379,N_419);
nor U1106 (N_1106,N_193,N_173);
or U1107 (N_1107,N_1,N_546);
nand U1108 (N_1108,N_12,N_859);
nand U1109 (N_1109,N_368,N_848);
xnor U1110 (N_1110,N_754,N_817);
or U1111 (N_1111,N_262,N_658);
and U1112 (N_1112,N_39,N_715);
nor U1113 (N_1113,N_575,N_873);
or U1114 (N_1114,N_677,N_284);
xnor U1115 (N_1115,N_233,N_51);
nor U1116 (N_1116,N_400,N_879);
or U1117 (N_1117,N_654,N_234);
nand U1118 (N_1118,N_180,N_738);
and U1119 (N_1119,N_686,N_101);
xor U1120 (N_1120,N_871,N_533);
nor U1121 (N_1121,N_104,N_663);
xor U1122 (N_1122,N_766,N_156);
xor U1123 (N_1123,N_862,N_115);
or U1124 (N_1124,N_271,N_971);
nand U1125 (N_1125,N_265,N_74);
nor U1126 (N_1126,N_627,N_719);
xor U1127 (N_1127,N_370,N_538);
and U1128 (N_1128,N_585,N_471);
nand U1129 (N_1129,N_158,N_867);
or U1130 (N_1130,N_753,N_277);
xor U1131 (N_1131,N_581,N_445);
nand U1132 (N_1132,N_339,N_548);
nand U1133 (N_1133,N_116,N_726);
and U1134 (N_1134,N_463,N_71);
or U1135 (N_1135,N_100,N_975);
nor U1136 (N_1136,N_433,N_394);
xnor U1137 (N_1137,N_765,N_390);
and U1138 (N_1138,N_377,N_520);
xor U1139 (N_1139,N_353,N_622);
and U1140 (N_1140,N_838,N_615);
nand U1141 (N_1141,N_300,N_309);
and U1142 (N_1142,N_771,N_391);
xnor U1143 (N_1143,N_369,N_323);
xor U1144 (N_1144,N_63,N_953);
nand U1145 (N_1145,N_710,N_306);
nand U1146 (N_1146,N_823,N_910);
nor U1147 (N_1147,N_365,N_964);
or U1148 (N_1148,N_746,N_672);
nor U1149 (N_1149,N_48,N_338);
nor U1150 (N_1150,N_269,N_636);
xnor U1151 (N_1151,N_167,N_439);
xor U1152 (N_1152,N_536,N_275);
nor U1153 (N_1153,N_62,N_938);
or U1154 (N_1154,N_436,N_980);
nor U1155 (N_1155,N_372,N_332);
nand U1156 (N_1156,N_501,N_385);
nand U1157 (N_1157,N_376,N_878);
and U1158 (N_1158,N_885,N_346);
nand U1159 (N_1159,N_652,N_415);
nor U1160 (N_1160,N_764,N_472);
nor U1161 (N_1161,N_611,N_992);
xor U1162 (N_1162,N_408,N_916);
or U1163 (N_1163,N_800,N_197);
or U1164 (N_1164,N_747,N_940);
and U1165 (N_1165,N_166,N_625);
or U1166 (N_1166,N_485,N_720);
or U1167 (N_1167,N_924,N_513);
nor U1168 (N_1168,N_606,N_983);
or U1169 (N_1169,N_412,N_289);
nor U1170 (N_1170,N_861,N_807);
or U1171 (N_1171,N_644,N_200);
and U1172 (N_1172,N_590,N_592);
nand U1173 (N_1173,N_605,N_218);
xnor U1174 (N_1174,N_294,N_381);
nand U1175 (N_1175,N_734,N_7);
nor U1176 (N_1176,N_287,N_31);
and U1177 (N_1177,N_767,N_854);
or U1178 (N_1178,N_0,N_290);
or U1179 (N_1179,N_92,N_597);
nand U1180 (N_1180,N_570,N_302);
nor U1181 (N_1181,N_763,N_578);
and U1182 (N_1182,N_237,N_349);
and U1183 (N_1183,N_178,N_215);
or U1184 (N_1184,N_559,N_99);
xnor U1185 (N_1185,N_305,N_986);
or U1186 (N_1186,N_616,N_736);
and U1187 (N_1187,N_491,N_109);
and U1188 (N_1188,N_213,N_966);
and U1189 (N_1189,N_222,N_34);
or U1190 (N_1190,N_880,N_728);
nor U1191 (N_1191,N_963,N_752);
and U1192 (N_1192,N_835,N_308);
and U1193 (N_1193,N_558,N_257);
nor U1194 (N_1194,N_703,N_179);
and U1195 (N_1195,N_814,N_779);
or U1196 (N_1196,N_669,N_718);
xor U1197 (N_1197,N_49,N_778);
nor U1198 (N_1198,N_310,N_514);
or U1199 (N_1199,N_844,N_500);
nand U1200 (N_1200,N_151,N_610);
or U1201 (N_1201,N_40,N_557);
nand U1202 (N_1202,N_364,N_994);
nand U1203 (N_1203,N_933,N_827);
or U1204 (N_1204,N_409,N_930);
and U1205 (N_1205,N_563,N_201);
and U1206 (N_1206,N_477,N_492);
nand U1207 (N_1207,N_261,N_604);
xor U1208 (N_1208,N_607,N_97);
and U1209 (N_1209,N_423,N_165);
xor U1210 (N_1210,N_706,N_342);
and U1211 (N_1211,N_414,N_723);
or U1212 (N_1212,N_206,N_942);
or U1213 (N_1213,N_344,N_329);
nor U1214 (N_1214,N_857,N_114);
xnor U1215 (N_1215,N_111,N_191);
xor U1216 (N_1216,N_793,N_203);
or U1217 (N_1217,N_13,N_52);
nor U1218 (N_1218,N_470,N_108);
xor U1219 (N_1219,N_941,N_733);
xor U1220 (N_1220,N_997,N_598);
xnor U1221 (N_1221,N_758,N_509);
or U1222 (N_1222,N_690,N_795);
xnor U1223 (N_1223,N_974,N_850);
and U1224 (N_1224,N_662,N_5);
xor U1225 (N_1225,N_449,N_670);
or U1226 (N_1226,N_934,N_223);
xnor U1227 (N_1227,N_324,N_561);
and U1228 (N_1228,N_896,N_781);
or U1229 (N_1229,N_374,N_487);
xor U1230 (N_1230,N_818,N_322);
xnor U1231 (N_1231,N_172,N_965);
and U1232 (N_1232,N_995,N_833);
nand U1233 (N_1233,N_441,N_594);
nor U1234 (N_1234,N_534,N_949);
and U1235 (N_1235,N_628,N_83);
nand U1236 (N_1236,N_834,N_482);
nand U1237 (N_1237,N_829,N_84);
or U1238 (N_1238,N_174,N_516);
xnor U1239 (N_1239,N_739,N_805);
and U1240 (N_1240,N_927,N_47);
and U1241 (N_1241,N_66,N_321);
xnor U1242 (N_1242,N_999,N_479);
nor U1243 (N_1243,N_147,N_657);
and U1244 (N_1244,N_434,N_161);
nand U1245 (N_1245,N_864,N_774);
nand U1246 (N_1246,N_511,N_320);
nor U1247 (N_1247,N_260,N_355);
and U1248 (N_1248,N_406,N_127);
and U1249 (N_1249,N_216,N_843);
and U1250 (N_1250,N_948,N_612);
and U1251 (N_1251,N_828,N_551);
xor U1252 (N_1252,N_130,N_977);
nor U1253 (N_1253,N_325,N_884);
and U1254 (N_1254,N_967,N_199);
nor U1255 (N_1255,N_554,N_26);
nor U1256 (N_1256,N_73,N_569);
or U1257 (N_1257,N_14,N_451);
or U1258 (N_1258,N_515,N_803);
and U1259 (N_1259,N_190,N_388);
and U1260 (N_1260,N_731,N_340);
and U1261 (N_1261,N_684,N_314);
and U1262 (N_1262,N_366,N_889);
nor U1263 (N_1263,N_812,N_757);
and U1264 (N_1264,N_717,N_481);
xor U1265 (N_1265,N_335,N_673);
xnor U1266 (N_1266,N_177,N_960);
or U1267 (N_1267,N_455,N_134);
nor U1268 (N_1268,N_783,N_735);
nor U1269 (N_1269,N_280,N_537);
nand U1270 (N_1270,N_224,N_527);
xnor U1271 (N_1271,N_693,N_2);
or U1272 (N_1272,N_499,N_617);
nor U1273 (N_1273,N_860,N_211);
nor U1274 (N_1274,N_621,N_904);
xnor U1275 (N_1275,N_776,N_711);
nand U1276 (N_1276,N_603,N_642);
nor U1277 (N_1277,N_60,N_564);
xor U1278 (N_1278,N_330,N_630);
or U1279 (N_1279,N_384,N_651);
or U1280 (N_1280,N_702,N_207);
nand U1281 (N_1281,N_897,N_431);
or U1282 (N_1282,N_291,N_985);
nand U1283 (N_1283,N_745,N_295);
nor U1284 (N_1284,N_53,N_968);
nor U1285 (N_1285,N_125,N_643);
nor U1286 (N_1286,N_11,N_777);
and U1287 (N_1287,N_331,N_649);
nand U1288 (N_1288,N_242,N_373);
or U1289 (N_1289,N_955,N_19);
xor U1290 (N_1290,N_722,N_890);
and U1291 (N_1291,N_484,N_954);
or U1292 (N_1292,N_131,N_221);
or U1293 (N_1293,N_973,N_958);
nor U1294 (N_1294,N_810,N_847);
nand U1295 (N_1295,N_716,N_918);
nor U1296 (N_1296,N_836,N_502);
nor U1297 (N_1297,N_540,N_490);
nand U1298 (N_1298,N_503,N_970);
nand U1299 (N_1299,N_371,N_351);
or U1300 (N_1300,N_498,N_397);
or U1301 (N_1301,N_993,N_468);
and U1302 (N_1302,N_24,N_931);
and U1303 (N_1303,N_398,N_464);
xnor U1304 (N_1304,N_352,N_667);
and U1305 (N_1305,N_813,N_613);
xor U1306 (N_1306,N_730,N_411);
xnor U1307 (N_1307,N_749,N_547);
or U1308 (N_1308,N_105,N_692);
and U1309 (N_1309,N_959,N_27);
nand U1310 (N_1310,N_507,N_725);
nor U1311 (N_1311,N_478,N_826);
or U1312 (N_1312,N_316,N_225);
and U1313 (N_1313,N_476,N_420);
xnor U1314 (N_1314,N_204,N_22);
nand U1315 (N_1315,N_645,N_696);
and U1316 (N_1316,N_469,N_691);
xnor U1317 (N_1317,N_205,N_28);
and U1318 (N_1318,N_665,N_41);
or U1319 (N_1319,N_655,N_453);
or U1320 (N_1320,N_832,N_582);
nand U1321 (N_1321,N_303,N_951);
xor U1322 (N_1322,N_486,N_571);
and U1323 (N_1323,N_962,N_106);
and U1324 (N_1324,N_919,N_32);
and U1325 (N_1325,N_681,N_825);
or U1326 (N_1326,N_258,N_524);
nand U1327 (N_1327,N_946,N_922);
xor U1328 (N_1328,N_292,N_188);
and U1329 (N_1329,N_526,N_694);
or U1330 (N_1330,N_148,N_782);
and U1331 (N_1331,N_508,N_72);
and U1332 (N_1332,N_160,N_584);
nor U1333 (N_1333,N_903,N_81);
or U1334 (N_1334,N_236,N_94);
xnor U1335 (N_1335,N_35,N_898);
and U1336 (N_1336,N_54,N_957);
or U1337 (N_1337,N_773,N_638);
nand U1338 (N_1338,N_539,N_96);
and U1339 (N_1339,N_666,N_361);
xor U1340 (N_1340,N_700,N_304);
nand U1341 (N_1341,N_998,N_629);
nand U1342 (N_1342,N_182,N_187);
xor U1343 (N_1343,N_894,N_680);
nor U1344 (N_1344,N_235,N_550);
nand U1345 (N_1345,N_797,N_82);
nor U1346 (N_1346,N_43,N_65);
and U1347 (N_1347,N_183,N_343);
and U1348 (N_1348,N_682,N_202);
and U1349 (N_1349,N_334,N_925);
nor U1350 (N_1350,N_653,N_877);
xor U1351 (N_1351,N_580,N_618);
and U1352 (N_1352,N_978,N_858);
and U1353 (N_1353,N_452,N_256);
and U1354 (N_1354,N_29,N_679);
nor U1355 (N_1355,N_939,N_113);
xnor U1356 (N_1356,N_55,N_926);
xor U1357 (N_1357,N_437,N_110);
and U1358 (N_1358,N_668,N_219);
and U1359 (N_1359,N_164,N_488);
nor U1360 (N_1360,N_602,N_675);
xor U1361 (N_1361,N_112,N_145);
xor U1362 (N_1362,N_75,N_159);
nor U1363 (N_1363,N_519,N_982);
nand U1364 (N_1364,N_313,N_270);
xor U1365 (N_1365,N_209,N_579);
xnor U1366 (N_1366,N_750,N_348);
and U1367 (N_1367,N_552,N_138);
or U1368 (N_1368,N_283,N_588);
or U1369 (N_1369,N_976,N_683);
xnor U1370 (N_1370,N_140,N_86);
nand U1371 (N_1371,N_461,N_497);
and U1372 (N_1372,N_90,N_150);
and U1373 (N_1373,N_704,N_87);
xnor U1374 (N_1374,N_357,N_405);
and U1375 (N_1375,N_956,N_422);
xor U1376 (N_1376,N_128,N_785);
xnor U1377 (N_1377,N_227,N_59);
nand U1378 (N_1378,N_929,N_297);
and U1379 (N_1379,N_124,N_531);
xor U1380 (N_1380,N_882,N_133);
nor U1381 (N_1381,N_979,N_278);
xor U1382 (N_1382,N_239,N_495);
nor U1383 (N_1383,N_18,N_921);
and U1384 (N_1384,N_157,N_424);
nand U1385 (N_1385,N_744,N_45);
nand U1386 (N_1386,N_760,N_641);
and U1387 (N_1387,N_909,N_16);
nor U1388 (N_1388,N_494,N_712);
and U1389 (N_1389,N_572,N_267);
or U1390 (N_1390,N_824,N_347);
and U1391 (N_1391,N_853,N_249);
xnor U1392 (N_1392,N_608,N_312);
xnor U1393 (N_1393,N_380,N_360);
nor U1394 (N_1394,N_184,N_6);
and U1395 (N_1395,N_631,N_240);
and U1396 (N_1396,N_194,N_132);
or U1397 (N_1397,N_740,N_46);
nand U1398 (N_1398,N_840,N_410);
xnor U1399 (N_1399,N_522,N_231);
and U1400 (N_1400,N_466,N_791);
nor U1401 (N_1401,N_741,N_44);
and U1402 (N_1402,N_77,N_600);
and U1403 (N_1403,N_119,N_640);
nand U1404 (N_1404,N_350,N_393);
xnor U1405 (N_1405,N_230,N_961);
or U1406 (N_1406,N_756,N_574);
and U1407 (N_1407,N_804,N_328);
and U1408 (N_1408,N_943,N_620);
or U1409 (N_1409,N_298,N_819);
xnor U1410 (N_1410,N_902,N_881);
nor U1411 (N_1411,N_143,N_914);
and U1412 (N_1412,N_378,N_888);
nand U1413 (N_1413,N_549,N_855);
or U1414 (N_1414,N_699,N_214);
nand U1415 (N_1415,N_944,N_169);
xnor U1416 (N_1416,N_869,N_886);
and U1417 (N_1417,N_601,N_413);
and U1418 (N_1418,N_689,N_506);
nand U1419 (N_1419,N_426,N_208);
nand U1420 (N_1420,N_475,N_250);
xnor U1421 (N_1421,N_634,N_952);
or U1422 (N_1422,N_905,N_609);
and U1423 (N_1423,N_336,N_695);
nor U1424 (N_1424,N_118,N_279);
nor U1425 (N_1425,N_195,N_37);
and U1426 (N_1426,N_458,N_589);
nor U1427 (N_1427,N_255,N_565);
or U1428 (N_1428,N_268,N_595);
nand U1429 (N_1429,N_483,N_560);
and U1430 (N_1430,N_489,N_243);
nand U1431 (N_1431,N_4,N_122);
or U1432 (N_1432,N_732,N_367);
xnor U1433 (N_1433,N_899,N_637);
xnor U1434 (N_1434,N_395,N_103);
nor U1435 (N_1435,N_67,N_318);
or U1436 (N_1436,N_586,N_769);
and U1437 (N_1437,N_78,N_228);
nand U1438 (N_1438,N_363,N_465);
xnor U1439 (N_1439,N_529,N_432);
xor U1440 (N_1440,N_407,N_761);
xor U1441 (N_1441,N_567,N_3);
nand U1442 (N_1442,N_428,N_599);
and U1443 (N_1443,N_528,N_286);
nor U1444 (N_1444,N_210,N_50);
or U1445 (N_1445,N_480,N_831);
or U1446 (N_1446,N_274,N_107);
xnor U1447 (N_1447,N_163,N_912);
nor U1448 (N_1448,N_521,N_544);
nand U1449 (N_1449,N_906,N_142);
and U1450 (N_1450,N_460,N_266);
nor U1451 (N_1451,N_317,N_932);
nor U1452 (N_1452,N_633,N_786);
nor U1453 (N_1453,N_440,N_396);
or U1454 (N_1454,N_790,N_530);
nor U1455 (N_1455,N_770,N_356);
nor U1456 (N_1456,N_402,N_102);
nand U1457 (N_1457,N_545,N_707);
xnor U1458 (N_1458,N_950,N_915);
and U1459 (N_1459,N_874,N_36);
nand U1460 (N_1460,N_56,N_676);
and U1461 (N_1461,N_245,N_149);
or U1462 (N_1462,N_806,N_253);
xor U1463 (N_1463,N_913,N_837);
and U1464 (N_1464,N_64,N_58);
xnor U1465 (N_1465,N_984,N_875);
and U1466 (N_1466,N_70,N_399);
nand U1467 (N_1467,N_232,N_248);
nand U1468 (N_1468,N_792,N_429);
or U1469 (N_1469,N_553,N_713);
and U1470 (N_1470,N_144,N_587);
nor U1471 (N_1471,N_171,N_345);
and U1472 (N_1472,N_755,N_246);
nand U1473 (N_1473,N_217,N_737);
or U1474 (N_1474,N_721,N_10);
nor U1475 (N_1475,N_762,N_811);
or U1476 (N_1476,N_727,N_98);
and U1477 (N_1477,N_989,N_252);
xnor U1478 (N_1478,N_991,N_136);
or U1479 (N_1479,N_650,N_85);
nand U1480 (N_1480,N_532,N_748);
or U1481 (N_1481,N_911,N_137);
nor U1482 (N_1482,N_895,N_935);
nand U1483 (N_1483,N_362,N_496);
nand U1484 (N_1484,N_870,N_170);
or U1485 (N_1485,N_583,N_969);
nand U1486 (N_1486,N_596,N_57);
nand U1487 (N_1487,N_315,N_181);
and U1488 (N_1488,N_23,N_555);
or U1489 (N_1489,N_141,N_129);
nor U1490 (N_1490,N_337,N_281);
xnor U1491 (N_1491,N_535,N_705);
or U1492 (N_1492,N_91,N_25);
nor U1493 (N_1493,N_42,N_263);
xor U1494 (N_1494,N_176,N_996);
or U1495 (N_1495,N_474,N_821);
nor U1496 (N_1496,N_688,N_891);
and U1497 (N_1497,N_512,N_272);
nor U1498 (N_1498,N_241,N_273);
nor U1499 (N_1499,N_139,N_299);
or U1500 (N_1500,N_346,N_531);
nand U1501 (N_1501,N_428,N_16);
or U1502 (N_1502,N_66,N_981);
nor U1503 (N_1503,N_124,N_958);
or U1504 (N_1504,N_245,N_235);
or U1505 (N_1505,N_852,N_730);
or U1506 (N_1506,N_625,N_87);
xor U1507 (N_1507,N_580,N_658);
nor U1508 (N_1508,N_533,N_869);
and U1509 (N_1509,N_461,N_22);
nor U1510 (N_1510,N_193,N_847);
nand U1511 (N_1511,N_734,N_491);
xor U1512 (N_1512,N_842,N_485);
nand U1513 (N_1513,N_547,N_650);
xnor U1514 (N_1514,N_275,N_128);
nor U1515 (N_1515,N_305,N_241);
nor U1516 (N_1516,N_304,N_495);
nor U1517 (N_1517,N_965,N_622);
nor U1518 (N_1518,N_15,N_889);
nor U1519 (N_1519,N_390,N_264);
nor U1520 (N_1520,N_514,N_583);
or U1521 (N_1521,N_801,N_879);
or U1522 (N_1522,N_746,N_347);
nand U1523 (N_1523,N_283,N_266);
nand U1524 (N_1524,N_765,N_620);
nand U1525 (N_1525,N_518,N_91);
or U1526 (N_1526,N_265,N_231);
or U1527 (N_1527,N_628,N_895);
or U1528 (N_1528,N_624,N_774);
xnor U1529 (N_1529,N_32,N_326);
nor U1530 (N_1530,N_420,N_446);
and U1531 (N_1531,N_15,N_579);
xnor U1532 (N_1532,N_958,N_190);
or U1533 (N_1533,N_642,N_526);
nor U1534 (N_1534,N_94,N_550);
xnor U1535 (N_1535,N_991,N_643);
nand U1536 (N_1536,N_179,N_266);
nor U1537 (N_1537,N_112,N_292);
or U1538 (N_1538,N_244,N_699);
or U1539 (N_1539,N_257,N_655);
nand U1540 (N_1540,N_9,N_398);
or U1541 (N_1541,N_741,N_132);
or U1542 (N_1542,N_446,N_406);
xnor U1543 (N_1543,N_480,N_762);
nand U1544 (N_1544,N_765,N_937);
nor U1545 (N_1545,N_642,N_548);
and U1546 (N_1546,N_484,N_155);
nor U1547 (N_1547,N_703,N_561);
nand U1548 (N_1548,N_702,N_22);
xor U1549 (N_1549,N_303,N_919);
or U1550 (N_1550,N_783,N_414);
or U1551 (N_1551,N_231,N_717);
xor U1552 (N_1552,N_222,N_375);
nand U1553 (N_1553,N_691,N_871);
xor U1554 (N_1554,N_730,N_601);
xnor U1555 (N_1555,N_685,N_779);
and U1556 (N_1556,N_769,N_763);
nand U1557 (N_1557,N_3,N_699);
xnor U1558 (N_1558,N_621,N_550);
and U1559 (N_1559,N_133,N_377);
nor U1560 (N_1560,N_601,N_652);
or U1561 (N_1561,N_693,N_794);
and U1562 (N_1562,N_169,N_843);
and U1563 (N_1563,N_1,N_813);
nor U1564 (N_1564,N_978,N_557);
and U1565 (N_1565,N_194,N_514);
nor U1566 (N_1566,N_686,N_409);
xnor U1567 (N_1567,N_504,N_917);
or U1568 (N_1568,N_90,N_937);
xnor U1569 (N_1569,N_27,N_53);
nor U1570 (N_1570,N_526,N_992);
nor U1571 (N_1571,N_343,N_565);
nor U1572 (N_1572,N_463,N_611);
and U1573 (N_1573,N_136,N_551);
and U1574 (N_1574,N_897,N_332);
nor U1575 (N_1575,N_508,N_402);
xor U1576 (N_1576,N_300,N_791);
xor U1577 (N_1577,N_797,N_98);
xnor U1578 (N_1578,N_308,N_606);
nand U1579 (N_1579,N_122,N_512);
or U1580 (N_1580,N_590,N_611);
nand U1581 (N_1581,N_681,N_777);
nor U1582 (N_1582,N_117,N_643);
and U1583 (N_1583,N_799,N_211);
xnor U1584 (N_1584,N_526,N_788);
or U1585 (N_1585,N_739,N_938);
nor U1586 (N_1586,N_971,N_320);
nor U1587 (N_1587,N_172,N_342);
or U1588 (N_1588,N_120,N_456);
nand U1589 (N_1589,N_727,N_37);
nand U1590 (N_1590,N_437,N_744);
nand U1591 (N_1591,N_849,N_379);
or U1592 (N_1592,N_645,N_625);
nor U1593 (N_1593,N_650,N_388);
nand U1594 (N_1594,N_192,N_254);
xor U1595 (N_1595,N_316,N_377);
nor U1596 (N_1596,N_362,N_147);
or U1597 (N_1597,N_310,N_89);
nand U1598 (N_1598,N_401,N_838);
nor U1599 (N_1599,N_634,N_754);
or U1600 (N_1600,N_863,N_188);
or U1601 (N_1601,N_602,N_137);
xnor U1602 (N_1602,N_379,N_142);
nand U1603 (N_1603,N_456,N_604);
nor U1604 (N_1604,N_289,N_449);
xnor U1605 (N_1605,N_195,N_311);
xnor U1606 (N_1606,N_103,N_418);
xnor U1607 (N_1607,N_844,N_204);
and U1608 (N_1608,N_869,N_625);
and U1609 (N_1609,N_153,N_705);
nand U1610 (N_1610,N_698,N_366);
nand U1611 (N_1611,N_986,N_120);
nand U1612 (N_1612,N_677,N_214);
nand U1613 (N_1613,N_537,N_112);
and U1614 (N_1614,N_954,N_926);
and U1615 (N_1615,N_441,N_415);
nand U1616 (N_1616,N_660,N_817);
and U1617 (N_1617,N_340,N_53);
or U1618 (N_1618,N_142,N_674);
xnor U1619 (N_1619,N_702,N_109);
nand U1620 (N_1620,N_730,N_614);
nor U1621 (N_1621,N_228,N_251);
nor U1622 (N_1622,N_241,N_715);
nand U1623 (N_1623,N_231,N_581);
xor U1624 (N_1624,N_792,N_467);
xor U1625 (N_1625,N_898,N_62);
xnor U1626 (N_1626,N_574,N_339);
and U1627 (N_1627,N_0,N_344);
and U1628 (N_1628,N_432,N_907);
or U1629 (N_1629,N_857,N_286);
or U1630 (N_1630,N_944,N_587);
and U1631 (N_1631,N_320,N_649);
xnor U1632 (N_1632,N_573,N_591);
nor U1633 (N_1633,N_896,N_94);
nor U1634 (N_1634,N_912,N_723);
xnor U1635 (N_1635,N_267,N_963);
or U1636 (N_1636,N_127,N_956);
nor U1637 (N_1637,N_931,N_751);
xor U1638 (N_1638,N_335,N_283);
nor U1639 (N_1639,N_666,N_944);
nor U1640 (N_1640,N_249,N_361);
nand U1641 (N_1641,N_966,N_866);
and U1642 (N_1642,N_875,N_995);
nand U1643 (N_1643,N_983,N_921);
nor U1644 (N_1644,N_379,N_910);
xnor U1645 (N_1645,N_141,N_991);
nand U1646 (N_1646,N_136,N_831);
xor U1647 (N_1647,N_387,N_515);
xor U1648 (N_1648,N_925,N_867);
nand U1649 (N_1649,N_456,N_133);
nand U1650 (N_1650,N_852,N_258);
or U1651 (N_1651,N_148,N_171);
xor U1652 (N_1652,N_530,N_906);
and U1653 (N_1653,N_486,N_156);
or U1654 (N_1654,N_689,N_135);
nand U1655 (N_1655,N_954,N_550);
and U1656 (N_1656,N_407,N_116);
nor U1657 (N_1657,N_85,N_217);
nor U1658 (N_1658,N_249,N_625);
xor U1659 (N_1659,N_695,N_424);
nand U1660 (N_1660,N_587,N_371);
nand U1661 (N_1661,N_709,N_788);
and U1662 (N_1662,N_208,N_686);
xnor U1663 (N_1663,N_551,N_494);
xnor U1664 (N_1664,N_875,N_362);
or U1665 (N_1665,N_629,N_589);
nand U1666 (N_1666,N_963,N_610);
xor U1667 (N_1667,N_251,N_528);
nand U1668 (N_1668,N_235,N_964);
nand U1669 (N_1669,N_252,N_546);
nor U1670 (N_1670,N_784,N_21);
nand U1671 (N_1671,N_24,N_417);
xnor U1672 (N_1672,N_949,N_88);
nor U1673 (N_1673,N_369,N_618);
nand U1674 (N_1674,N_407,N_510);
nand U1675 (N_1675,N_629,N_65);
xnor U1676 (N_1676,N_87,N_86);
or U1677 (N_1677,N_778,N_869);
nand U1678 (N_1678,N_192,N_997);
and U1679 (N_1679,N_946,N_745);
nand U1680 (N_1680,N_50,N_679);
nand U1681 (N_1681,N_783,N_790);
xnor U1682 (N_1682,N_961,N_42);
and U1683 (N_1683,N_708,N_404);
xor U1684 (N_1684,N_184,N_367);
nor U1685 (N_1685,N_544,N_480);
or U1686 (N_1686,N_74,N_757);
and U1687 (N_1687,N_356,N_312);
or U1688 (N_1688,N_269,N_822);
nand U1689 (N_1689,N_47,N_538);
nand U1690 (N_1690,N_144,N_309);
and U1691 (N_1691,N_370,N_399);
xor U1692 (N_1692,N_612,N_820);
or U1693 (N_1693,N_230,N_530);
nand U1694 (N_1694,N_123,N_161);
and U1695 (N_1695,N_476,N_174);
and U1696 (N_1696,N_466,N_464);
and U1697 (N_1697,N_258,N_182);
and U1698 (N_1698,N_857,N_552);
nor U1699 (N_1699,N_478,N_614);
and U1700 (N_1700,N_667,N_278);
and U1701 (N_1701,N_334,N_951);
and U1702 (N_1702,N_340,N_212);
nor U1703 (N_1703,N_99,N_778);
and U1704 (N_1704,N_287,N_239);
nor U1705 (N_1705,N_39,N_189);
or U1706 (N_1706,N_240,N_433);
xnor U1707 (N_1707,N_706,N_881);
or U1708 (N_1708,N_941,N_97);
or U1709 (N_1709,N_491,N_406);
nand U1710 (N_1710,N_341,N_665);
and U1711 (N_1711,N_760,N_560);
xor U1712 (N_1712,N_351,N_763);
and U1713 (N_1713,N_153,N_839);
nand U1714 (N_1714,N_860,N_698);
and U1715 (N_1715,N_483,N_172);
nand U1716 (N_1716,N_551,N_45);
and U1717 (N_1717,N_411,N_690);
or U1718 (N_1718,N_924,N_256);
nand U1719 (N_1719,N_71,N_301);
nor U1720 (N_1720,N_859,N_968);
or U1721 (N_1721,N_806,N_759);
nor U1722 (N_1722,N_941,N_259);
or U1723 (N_1723,N_517,N_496);
or U1724 (N_1724,N_207,N_288);
or U1725 (N_1725,N_99,N_354);
xor U1726 (N_1726,N_372,N_187);
xnor U1727 (N_1727,N_269,N_735);
nand U1728 (N_1728,N_503,N_483);
nor U1729 (N_1729,N_256,N_98);
or U1730 (N_1730,N_940,N_296);
xor U1731 (N_1731,N_726,N_308);
nor U1732 (N_1732,N_26,N_680);
or U1733 (N_1733,N_588,N_178);
nor U1734 (N_1734,N_321,N_670);
or U1735 (N_1735,N_38,N_837);
or U1736 (N_1736,N_729,N_962);
xnor U1737 (N_1737,N_641,N_887);
nand U1738 (N_1738,N_520,N_239);
nor U1739 (N_1739,N_318,N_192);
xor U1740 (N_1740,N_333,N_939);
xnor U1741 (N_1741,N_259,N_615);
nand U1742 (N_1742,N_834,N_264);
xnor U1743 (N_1743,N_409,N_164);
or U1744 (N_1744,N_140,N_369);
nand U1745 (N_1745,N_135,N_261);
or U1746 (N_1746,N_692,N_562);
and U1747 (N_1747,N_486,N_344);
xnor U1748 (N_1748,N_43,N_604);
and U1749 (N_1749,N_81,N_920);
nor U1750 (N_1750,N_183,N_299);
nor U1751 (N_1751,N_264,N_103);
nand U1752 (N_1752,N_381,N_606);
xor U1753 (N_1753,N_260,N_876);
or U1754 (N_1754,N_493,N_271);
xor U1755 (N_1755,N_477,N_909);
and U1756 (N_1756,N_65,N_544);
nand U1757 (N_1757,N_297,N_976);
or U1758 (N_1758,N_295,N_764);
or U1759 (N_1759,N_531,N_623);
xor U1760 (N_1760,N_923,N_778);
or U1761 (N_1761,N_625,N_886);
nand U1762 (N_1762,N_753,N_362);
nor U1763 (N_1763,N_26,N_96);
nor U1764 (N_1764,N_845,N_338);
xor U1765 (N_1765,N_273,N_166);
and U1766 (N_1766,N_260,N_99);
nand U1767 (N_1767,N_268,N_888);
and U1768 (N_1768,N_982,N_463);
nand U1769 (N_1769,N_99,N_556);
nand U1770 (N_1770,N_673,N_580);
nor U1771 (N_1771,N_85,N_75);
or U1772 (N_1772,N_737,N_512);
or U1773 (N_1773,N_44,N_84);
or U1774 (N_1774,N_800,N_909);
nand U1775 (N_1775,N_960,N_429);
xor U1776 (N_1776,N_39,N_696);
nand U1777 (N_1777,N_194,N_817);
and U1778 (N_1778,N_377,N_930);
or U1779 (N_1779,N_738,N_619);
nand U1780 (N_1780,N_660,N_963);
xnor U1781 (N_1781,N_173,N_941);
nor U1782 (N_1782,N_983,N_276);
and U1783 (N_1783,N_115,N_522);
xnor U1784 (N_1784,N_938,N_944);
and U1785 (N_1785,N_88,N_509);
xor U1786 (N_1786,N_881,N_302);
xnor U1787 (N_1787,N_994,N_246);
nand U1788 (N_1788,N_284,N_506);
nor U1789 (N_1789,N_575,N_384);
or U1790 (N_1790,N_411,N_56);
nand U1791 (N_1791,N_616,N_497);
and U1792 (N_1792,N_756,N_55);
nand U1793 (N_1793,N_285,N_990);
nand U1794 (N_1794,N_740,N_656);
nand U1795 (N_1795,N_493,N_521);
and U1796 (N_1796,N_547,N_797);
xor U1797 (N_1797,N_751,N_281);
nand U1798 (N_1798,N_654,N_470);
and U1799 (N_1799,N_311,N_879);
xnor U1800 (N_1800,N_790,N_670);
and U1801 (N_1801,N_944,N_755);
and U1802 (N_1802,N_155,N_24);
nand U1803 (N_1803,N_358,N_101);
xnor U1804 (N_1804,N_165,N_56);
xor U1805 (N_1805,N_883,N_534);
or U1806 (N_1806,N_704,N_967);
nand U1807 (N_1807,N_428,N_358);
or U1808 (N_1808,N_447,N_963);
nand U1809 (N_1809,N_746,N_663);
or U1810 (N_1810,N_172,N_484);
nor U1811 (N_1811,N_757,N_404);
xnor U1812 (N_1812,N_724,N_738);
xor U1813 (N_1813,N_692,N_366);
nand U1814 (N_1814,N_732,N_182);
nor U1815 (N_1815,N_864,N_998);
nor U1816 (N_1816,N_665,N_462);
nand U1817 (N_1817,N_748,N_120);
xor U1818 (N_1818,N_216,N_757);
and U1819 (N_1819,N_349,N_467);
and U1820 (N_1820,N_903,N_961);
and U1821 (N_1821,N_20,N_967);
and U1822 (N_1822,N_408,N_92);
nor U1823 (N_1823,N_662,N_726);
nor U1824 (N_1824,N_990,N_774);
xor U1825 (N_1825,N_527,N_72);
or U1826 (N_1826,N_609,N_542);
or U1827 (N_1827,N_160,N_765);
nand U1828 (N_1828,N_944,N_789);
nand U1829 (N_1829,N_995,N_885);
xnor U1830 (N_1830,N_670,N_11);
and U1831 (N_1831,N_706,N_846);
or U1832 (N_1832,N_197,N_55);
xnor U1833 (N_1833,N_856,N_406);
nor U1834 (N_1834,N_284,N_627);
xnor U1835 (N_1835,N_978,N_654);
nand U1836 (N_1836,N_433,N_188);
xor U1837 (N_1837,N_958,N_596);
and U1838 (N_1838,N_991,N_873);
nand U1839 (N_1839,N_957,N_113);
nand U1840 (N_1840,N_862,N_81);
xor U1841 (N_1841,N_278,N_595);
or U1842 (N_1842,N_211,N_339);
nor U1843 (N_1843,N_434,N_914);
or U1844 (N_1844,N_578,N_286);
or U1845 (N_1845,N_314,N_120);
xnor U1846 (N_1846,N_888,N_641);
nand U1847 (N_1847,N_90,N_137);
and U1848 (N_1848,N_30,N_477);
or U1849 (N_1849,N_291,N_774);
and U1850 (N_1850,N_648,N_337);
nor U1851 (N_1851,N_280,N_759);
and U1852 (N_1852,N_40,N_147);
xor U1853 (N_1853,N_109,N_874);
or U1854 (N_1854,N_400,N_602);
and U1855 (N_1855,N_953,N_797);
or U1856 (N_1856,N_898,N_713);
or U1857 (N_1857,N_443,N_988);
or U1858 (N_1858,N_754,N_941);
or U1859 (N_1859,N_173,N_391);
or U1860 (N_1860,N_707,N_198);
nand U1861 (N_1861,N_99,N_500);
and U1862 (N_1862,N_834,N_675);
and U1863 (N_1863,N_264,N_23);
nor U1864 (N_1864,N_175,N_703);
and U1865 (N_1865,N_490,N_211);
nor U1866 (N_1866,N_642,N_338);
or U1867 (N_1867,N_288,N_212);
xor U1868 (N_1868,N_9,N_527);
nor U1869 (N_1869,N_412,N_339);
or U1870 (N_1870,N_568,N_6);
or U1871 (N_1871,N_878,N_349);
and U1872 (N_1872,N_323,N_221);
and U1873 (N_1873,N_759,N_422);
and U1874 (N_1874,N_787,N_251);
and U1875 (N_1875,N_748,N_150);
xor U1876 (N_1876,N_891,N_585);
xor U1877 (N_1877,N_991,N_964);
or U1878 (N_1878,N_147,N_508);
and U1879 (N_1879,N_755,N_502);
and U1880 (N_1880,N_60,N_409);
nor U1881 (N_1881,N_30,N_523);
or U1882 (N_1882,N_676,N_243);
xor U1883 (N_1883,N_796,N_220);
or U1884 (N_1884,N_442,N_88);
nand U1885 (N_1885,N_238,N_164);
nand U1886 (N_1886,N_988,N_931);
and U1887 (N_1887,N_40,N_784);
and U1888 (N_1888,N_912,N_477);
nand U1889 (N_1889,N_997,N_726);
and U1890 (N_1890,N_630,N_979);
nand U1891 (N_1891,N_615,N_388);
and U1892 (N_1892,N_74,N_357);
xor U1893 (N_1893,N_179,N_507);
or U1894 (N_1894,N_108,N_344);
and U1895 (N_1895,N_809,N_509);
xor U1896 (N_1896,N_109,N_439);
nor U1897 (N_1897,N_933,N_993);
nor U1898 (N_1898,N_197,N_461);
nand U1899 (N_1899,N_906,N_588);
nand U1900 (N_1900,N_637,N_935);
nor U1901 (N_1901,N_212,N_146);
xor U1902 (N_1902,N_29,N_725);
xnor U1903 (N_1903,N_901,N_725);
nand U1904 (N_1904,N_327,N_559);
nand U1905 (N_1905,N_282,N_497);
and U1906 (N_1906,N_409,N_380);
nand U1907 (N_1907,N_190,N_91);
or U1908 (N_1908,N_987,N_538);
or U1909 (N_1909,N_890,N_59);
nand U1910 (N_1910,N_917,N_711);
or U1911 (N_1911,N_570,N_852);
nand U1912 (N_1912,N_935,N_640);
nor U1913 (N_1913,N_563,N_773);
xor U1914 (N_1914,N_104,N_907);
or U1915 (N_1915,N_447,N_625);
xnor U1916 (N_1916,N_32,N_18);
or U1917 (N_1917,N_643,N_835);
and U1918 (N_1918,N_149,N_126);
and U1919 (N_1919,N_111,N_4);
nor U1920 (N_1920,N_863,N_279);
nand U1921 (N_1921,N_576,N_710);
and U1922 (N_1922,N_74,N_341);
or U1923 (N_1923,N_575,N_519);
nand U1924 (N_1924,N_184,N_60);
or U1925 (N_1925,N_800,N_347);
nor U1926 (N_1926,N_942,N_484);
and U1927 (N_1927,N_689,N_88);
or U1928 (N_1928,N_275,N_761);
or U1929 (N_1929,N_404,N_833);
nand U1930 (N_1930,N_742,N_768);
xor U1931 (N_1931,N_918,N_277);
and U1932 (N_1932,N_759,N_203);
nand U1933 (N_1933,N_923,N_422);
nor U1934 (N_1934,N_895,N_530);
nor U1935 (N_1935,N_644,N_798);
xor U1936 (N_1936,N_983,N_33);
nand U1937 (N_1937,N_672,N_836);
or U1938 (N_1938,N_594,N_193);
and U1939 (N_1939,N_695,N_822);
xor U1940 (N_1940,N_569,N_805);
and U1941 (N_1941,N_638,N_873);
nand U1942 (N_1942,N_31,N_792);
xor U1943 (N_1943,N_75,N_506);
and U1944 (N_1944,N_88,N_931);
and U1945 (N_1945,N_175,N_32);
nor U1946 (N_1946,N_344,N_917);
xor U1947 (N_1947,N_829,N_720);
xor U1948 (N_1948,N_38,N_785);
or U1949 (N_1949,N_569,N_292);
nand U1950 (N_1950,N_163,N_940);
nor U1951 (N_1951,N_496,N_225);
nor U1952 (N_1952,N_144,N_292);
or U1953 (N_1953,N_343,N_650);
or U1954 (N_1954,N_890,N_485);
or U1955 (N_1955,N_676,N_53);
nor U1956 (N_1956,N_520,N_533);
xnor U1957 (N_1957,N_648,N_404);
nand U1958 (N_1958,N_256,N_353);
nor U1959 (N_1959,N_918,N_486);
nor U1960 (N_1960,N_646,N_149);
or U1961 (N_1961,N_804,N_431);
nor U1962 (N_1962,N_407,N_462);
or U1963 (N_1963,N_393,N_867);
nor U1964 (N_1964,N_534,N_952);
xor U1965 (N_1965,N_136,N_855);
nor U1966 (N_1966,N_683,N_765);
nand U1967 (N_1967,N_462,N_721);
nand U1968 (N_1968,N_433,N_832);
and U1969 (N_1969,N_10,N_75);
and U1970 (N_1970,N_648,N_465);
xor U1971 (N_1971,N_531,N_52);
and U1972 (N_1972,N_539,N_621);
and U1973 (N_1973,N_735,N_198);
and U1974 (N_1974,N_782,N_637);
xor U1975 (N_1975,N_546,N_92);
xnor U1976 (N_1976,N_462,N_366);
nor U1977 (N_1977,N_954,N_907);
nand U1978 (N_1978,N_786,N_386);
or U1979 (N_1979,N_522,N_12);
xor U1980 (N_1980,N_971,N_608);
nor U1981 (N_1981,N_764,N_884);
nand U1982 (N_1982,N_639,N_740);
and U1983 (N_1983,N_903,N_157);
xor U1984 (N_1984,N_689,N_892);
nand U1985 (N_1985,N_59,N_85);
and U1986 (N_1986,N_22,N_462);
and U1987 (N_1987,N_283,N_343);
and U1988 (N_1988,N_120,N_368);
nor U1989 (N_1989,N_241,N_563);
or U1990 (N_1990,N_843,N_936);
xnor U1991 (N_1991,N_351,N_67);
or U1992 (N_1992,N_825,N_4);
and U1993 (N_1993,N_973,N_933);
xor U1994 (N_1994,N_526,N_754);
or U1995 (N_1995,N_938,N_894);
nor U1996 (N_1996,N_274,N_830);
and U1997 (N_1997,N_141,N_701);
xor U1998 (N_1998,N_70,N_339);
xor U1999 (N_1999,N_381,N_342);
xor U2000 (N_2000,N_1579,N_1504);
nand U2001 (N_2001,N_1490,N_1422);
or U2002 (N_2002,N_1054,N_1330);
nand U2003 (N_2003,N_1898,N_1272);
xor U2004 (N_2004,N_1952,N_1282);
and U2005 (N_2005,N_1912,N_1210);
and U2006 (N_2006,N_1373,N_1318);
nor U2007 (N_2007,N_1388,N_1602);
nor U2008 (N_2008,N_1804,N_1917);
and U2009 (N_2009,N_1637,N_1578);
or U2010 (N_2010,N_1135,N_1420);
nand U2011 (N_2011,N_1093,N_1699);
xor U2012 (N_2012,N_1295,N_1499);
or U2013 (N_2013,N_1261,N_1718);
nand U2014 (N_2014,N_1211,N_1307);
nand U2015 (N_2015,N_1344,N_1667);
and U2016 (N_2016,N_1893,N_1516);
nand U2017 (N_2017,N_1111,N_1956);
nand U2018 (N_2018,N_1584,N_1438);
xor U2019 (N_2019,N_1421,N_1145);
nor U2020 (N_2020,N_1765,N_1216);
or U2021 (N_2021,N_1920,N_1041);
nor U2022 (N_2022,N_1990,N_1911);
xnor U2023 (N_2023,N_1779,N_1062);
nand U2024 (N_2024,N_1725,N_1037);
or U2025 (N_2025,N_1019,N_1632);
nand U2026 (N_2026,N_1970,N_1255);
or U2027 (N_2027,N_1554,N_1189);
nand U2028 (N_2028,N_1839,N_1007);
or U2029 (N_2029,N_1716,N_1266);
xor U2030 (N_2030,N_1885,N_1121);
or U2031 (N_2031,N_1994,N_1565);
and U2032 (N_2032,N_1739,N_1158);
nor U2033 (N_2033,N_1692,N_1751);
and U2034 (N_2034,N_1620,N_1348);
nand U2035 (N_2035,N_1673,N_1288);
nor U2036 (N_2036,N_1112,N_1088);
nor U2037 (N_2037,N_1810,N_1290);
nor U2038 (N_2038,N_1657,N_1817);
nor U2039 (N_2039,N_1557,N_1709);
xor U2040 (N_2040,N_1489,N_1091);
xnor U2041 (N_2041,N_1863,N_1649);
or U2042 (N_2042,N_1205,N_1841);
xor U2043 (N_2043,N_1476,N_1232);
and U2044 (N_2044,N_1224,N_1221);
nand U2045 (N_2045,N_1212,N_1249);
or U2046 (N_2046,N_1443,N_1464);
or U2047 (N_2047,N_1943,N_1909);
xor U2048 (N_2048,N_1460,N_1923);
or U2049 (N_2049,N_1387,N_1745);
and U2050 (N_2050,N_1555,N_1774);
or U2051 (N_2051,N_1461,N_1381);
or U2052 (N_2052,N_1500,N_1071);
nor U2053 (N_2053,N_1764,N_1333);
nand U2054 (N_2054,N_1069,N_1389);
or U2055 (N_2055,N_1619,N_1030);
xor U2056 (N_2056,N_1763,N_1177);
nor U2057 (N_2057,N_1941,N_1454);
or U2058 (N_2058,N_1782,N_1197);
nand U2059 (N_2059,N_1060,N_1860);
xor U2060 (N_2060,N_1983,N_1222);
xor U2061 (N_2061,N_1978,N_1524);
and U2062 (N_2062,N_1077,N_1834);
and U2063 (N_2063,N_1679,N_1016);
nor U2064 (N_2064,N_1188,N_1332);
xnor U2065 (N_2065,N_1882,N_1690);
xor U2066 (N_2066,N_1129,N_1564);
xor U2067 (N_2067,N_1992,N_1090);
or U2068 (N_2068,N_1998,N_1240);
and U2069 (N_2069,N_1595,N_1850);
nor U2070 (N_2070,N_1650,N_1004);
xor U2071 (N_2071,N_1870,N_1130);
and U2072 (N_2072,N_1410,N_1270);
nor U2073 (N_2073,N_1230,N_1819);
nor U2074 (N_2074,N_1024,N_1651);
nand U2075 (N_2075,N_1588,N_1097);
and U2076 (N_2076,N_1648,N_1049);
nor U2077 (N_2077,N_1456,N_1823);
and U2078 (N_2078,N_1302,N_1052);
and U2079 (N_2079,N_1572,N_1323);
nor U2080 (N_2080,N_1877,N_1937);
nor U2081 (N_2081,N_1191,N_1193);
or U2082 (N_2082,N_1787,N_1689);
and U2083 (N_2083,N_1283,N_1018);
nor U2084 (N_2084,N_1328,N_1467);
xor U2085 (N_2085,N_1811,N_1873);
or U2086 (N_2086,N_1644,N_1525);
xnor U2087 (N_2087,N_1192,N_1435);
nor U2088 (N_2088,N_1708,N_1631);
or U2089 (N_2089,N_1748,N_1675);
xnor U2090 (N_2090,N_1510,N_1587);
nand U2091 (N_2091,N_1600,N_1700);
nor U2092 (N_2092,N_1124,N_1132);
nand U2093 (N_2093,N_1895,N_1790);
xnor U2094 (N_2094,N_1605,N_1022);
nand U2095 (N_2095,N_1768,N_1393);
and U2096 (N_2096,N_1292,N_1173);
nand U2097 (N_2097,N_1369,N_1806);
nor U2098 (N_2098,N_1026,N_1519);
and U2099 (N_2099,N_1082,N_1084);
nor U2100 (N_2100,N_1465,N_1663);
or U2101 (N_2101,N_1549,N_1902);
or U2102 (N_2102,N_1820,N_1728);
nor U2103 (N_2103,N_1246,N_1714);
nand U2104 (N_2104,N_1967,N_1710);
nand U2105 (N_2105,N_1220,N_1000);
and U2106 (N_2106,N_1131,N_1206);
nor U2107 (N_2107,N_1845,N_1691);
or U2108 (N_2108,N_1033,N_1469);
and U2109 (N_2109,N_1342,N_1159);
or U2110 (N_2110,N_1652,N_1080);
xnor U2111 (N_2111,N_1753,N_1532);
and U2112 (N_2112,N_1788,N_1264);
nand U2113 (N_2113,N_1375,N_1696);
nand U2114 (N_2114,N_1045,N_1259);
or U2115 (N_2115,N_1048,N_1304);
xor U2116 (N_2116,N_1281,N_1448);
nor U2117 (N_2117,N_1223,N_1854);
nor U2118 (N_2118,N_1756,N_1309);
nor U2119 (N_2119,N_1544,N_1047);
or U2120 (N_2120,N_1357,N_1042);
xor U2121 (N_2121,N_1953,N_1615);
and U2122 (N_2122,N_1875,N_1398);
nor U2123 (N_2123,N_1451,N_1163);
nand U2124 (N_2124,N_1546,N_1248);
nand U2125 (N_2125,N_1827,N_1997);
and U2126 (N_2126,N_1301,N_1027);
nor U2127 (N_2127,N_1948,N_1066);
xor U2128 (N_2128,N_1833,N_1053);
and U2129 (N_2129,N_1161,N_1686);
xor U2130 (N_2130,N_1889,N_1012);
nand U2131 (N_2131,N_1432,N_1701);
and U2132 (N_2132,N_1401,N_1390);
or U2133 (N_2133,N_1878,N_1798);
and U2134 (N_2134,N_1263,N_1128);
xnor U2135 (N_2135,N_1236,N_1299);
and U2136 (N_2136,N_1791,N_1829);
and U2137 (N_2137,N_1972,N_1168);
nand U2138 (N_2138,N_1868,N_1317);
and U2139 (N_2139,N_1008,N_1979);
and U2140 (N_2140,N_1147,N_1591);
nor U2141 (N_2141,N_1784,N_1757);
xor U2142 (N_2142,N_1645,N_1310);
xor U2143 (N_2143,N_1403,N_1512);
nor U2144 (N_2144,N_1092,N_1639);
and U2145 (N_2145,N_1103,N_1471);
xnor U2146 (N_2146,N_1174,N_1086);
xor U2147 (N_2147,N_1431,N_1297);
xor U2148 (N_2148,N_1859,N_1562);
or U2149 (N_2149,N_1133,N_1795);
nor U2150 (N_2150,N_1630,N_1102);
nand U2151 (N_2151,N_1537,N_1356);
and U2152 (N_2152,N_1918,N_1237);
nand U2153 (N_2153,N_1640,N_1148);
nand U2154 (N_2154,N_1606,N_1761);
xor U2155 (N_2155,N_1813,N_1522);
nor U2156 (N_2156,N_1190,N_1569);
and U2157 (N_2157,N_1940,N_1906);
nand U2158 (N_2158,N_1105,N_1151);
or U2159 (N_2159,N_1265,N_1382);
or U2160 (N_2160,N_1711,N_1296);
and U2161 (N_2161,N_1869,N_1169);
nand U2162 (N_2162,N_1995,N_1267);
xnor U2163 (N_2163,N_1553,N_1526);
xnor U2164 (N_2164,N_1647,N_1786);
nor U2165 (N_2165,N_1364,N_1427);
nand U2166 (N_2166,N_1225,N_1021);
xor U2167 (N_2167,N_1036,N_1634);
or U2168 (N_2168,N_1530,N_1609);
nand U2169 (N_2169,N_1843,N_1586);
or U2170 (N_2170,N_1039,N_1963);
xor U2171 (N_2171,N_1046,N_1442);
nor U2172 (N_2172,N_1853,N_1621);
or U2173 (N_2173,N_1440,N_1029);
and U2174 (N_2174,N_1737,N_1271);
or U2175 (N_2175,N_1372,N_1095);
or U2176 (N_2176,N_1417,N_1959);
xnor U2177 (N_2177,N_1340,N_1981);
or U2178 (N_2178,N_1862,N_1883);
or U2179 (N_2179,N_1073,N_1646);
nand U2180 (N_2180,N_1423,N_1034);
nand U2181 (N_2181,N_1391,N_1472);
xnor U2182 (N_2182,N_1167,N_1762);
and U2183 (N_2183,N_1365,N_1180);
nand U2184 (N_2184,N_1684,N_1613);
nand U2185 (N_2185,N_1919,N_1104);
xnor U2186 (N_2186,N_1478,N_1927);
xor U2187 (N_2187,N_1463,N_1153);
and U2188 (N_2188,N_1485,N_1933);
nor U2189 (N_2189,N_1628,N_1611);
nor U2190 (N_2190,N_1429,N_1867);
nor U2191 (N_2191,N_1426,N_1346);
or U2192 (N_2192,N_1723,N_1141);
nor U2193 (N_2193,N_1334,N_1107);
xor U2194 (N_2194,N_1503,N_1961);
xor U2195 (N_2195,N_1496,N_1368);
xnor U2196 (N_2196,N_1257,N_1155);
or U2197 (N_2197,N_1558,N_1406);
xnor U2198 (N_2198,N_1362,N_1314);
xor U2199 (N_2199,N_1685,N_1734);
nor U2200 (N_2200,N_1229,N_1234);
or U2201 (N_2201,N_1541,N_1379);
or U2202 (N_2202,N_1597,N_1468);
and U2203 (N_2203,N_1766,N_1688);
nand U2204 (N_2204,N_1152,N_1962);
or U2205 (N_2205,N_1306,N_1198);
or U2206 (N_2206,N_1925,N_1089);
xnor U2207 (N_2207,N_1003,N_1740);
xor U2208 (N_2208,N_1020,N_1542);
and U2209 (N_2209,N_1010,N_1146);
nand U2210 (N_2210,N_1035,N_1109);
and U2211 (N_2211,N_1023,N_1722);
nand U2212 (N_2212,N_1642,N_1445);
nand U2213 (N_2213,N_1217,N_1808);
nand U2214 (N_2214,N_1358,N_1079);
xor U2215 (N_2215,N_1293,N_1098);
xor U2216 (N_2216,N_1258,N_1444);
and U2217 (N_2217,N_1363,N_1319);
or U2218 (N_2218,N_1057,N_1832);
nor U2219 (N_2219,N_1209,N_1985);
and U2220 (N_2220,N_1497,N_1437);
nor U2221 (N_2221,N_1245,N_1777);
nand U2222 (N_2222,N_1987,N_1337);
and U2223 (N_2223,N_1074,N_1395);
xor U2224 (N_2224,N_1719,N_1625);
or U2225 (N_2225,N_1849,N_1114);
nand U2226 (N_2226,N_1352,N_1502);
or U2227 (N_2227,N_1311,N_1575);
or U2228 (N_2228,N_1947,N_1848);
nand U2229 (N_2229,N_1374,N_1446);
and U2230 (N_2230,N_1687,N_1670);
xnor U2231 (N_2231,N_1165,N_1831);
or U2232 (N_2232,N_1252,N_1612);
or U2233 (N_2233,N_1694,N_1922);
or U2234 (N_2234,N_1697,N_1498);
and U2235 (N_2235,N_1596,N_1874);
nand U2236 (N_2236,N_1488,N_1371);
xnor U2237 (N_2237,N_1759,N_1861);
nand U2238 (N_2238,N_1935,N_1123);
xor U2239 (N_2239,N_1247,N_1428);
nand U2240 (N_2240,N_1812,N_1207);
and U2241 (N_2241,N_1715,N_1244);
nand U2242 (N_2242,N_1325,N_1914);
nor U2243 (N_2243,N_1884,N_1286);
xnor U2244 (N_2244,N_1936,N_1682);
nand U2245 (N_2245,N_1561,N_1031);
xnor U2246 (N_2246,N_1603,N_1964);
or U2247 (N_2247,N_1775,N_1164);
nand U2248 (N_2248,N_1618,N_1083);
nand U2249 (N_2249,N_1322,N_1744);
nand U2250 (N_2250,N_1338,N_1495);
xnor U2251 (N_2251,N_1559,N_1355);
or U2252 (N_2252,N_1085,N_1926);
xnor U2253 (N_2253,N_1359,N_1666);
or U2254 (N_2254,N_1608,N_1622);
or U2255 (N_2255,N_1858,N_1780);
and U2256 (N_2256,N_1397,N_1094);
nand U2257 (N_2257,N_1533,N_1106);
or U2258 (N_2258,N_1730,N_1186);
xor U2259 (N_2259,N_1857,N_1514);
and U2260 (N_2260,N_1156,N_1733);
and U2261 (N_2261,N_1396,N_1743);
xnor U2262 (N_2262,N_1616,N_1453);
or U2263 (N_2263,N_1957,N_1816);
or U2264 (N_2264,N_1269,N_1966);
nand U2265 (N_2265,N_1360,N_1814);
xor U2266 (N_2266,N_1415,N_1385);
nand U2267 (N_2267,N_1096,N_1900);
and U2268 (N_2268,N_1001,N_1942);
xnor U2269 (N_2269,N_1720,N_1916);
or U2270 (N_2270,N_1032,N_1413);
nand U2271 (N_2271,N_1695,N_1162);
or U2272 (N_2272,N_1305,N_1050);
and U2273 (N_2273,N_1969,N_1243);
or U2274 (N_2274,N_1386,N_1517);
or U2275 (N_2275,N_1507,N_1005);
xor U2276 (N_2276,N_1072,N_1181);
nand U2277 (N_2277,N_1932,N_1002);
and U2278 (N_2278,N_1626,N_1674);
or U2279 (N_2279,N_1518,N_1137);
and U2280 (N_2280,N_1452,N_1480);
nand U2281 (N_2281,N_1576,N_1044);
and U2282 (N_2282,N_1303,N_1930);
and U2283 (N_2283,N_1108,N_1924);
nor U2284 (N_2284,N_1436,N_1607);
or U2285 (N_2285,N_1971,N_1989);
or U2286 (N_2286,N_1614,N_1231);
or U2287 (N_2287,N_1797,N_1081);
nand U2288 (N_2288,N_1552,N_1056);
and U2289 (N_2289,N_1199,N_1599);
or U2290 (N_2290,N_1732,N_1439);
nand U2291 (N_2291,N_1624,N_1891);
nand U2292 (N_2292,N_1219,N_1545);
and U2293 (N_2293,N_1425,N_1126);
xor U2294 (N_2294,N_1384,N_1075);
and U2295 (N_2295,N_1704,N_1218);
and U2296 (N_2296,N_1771,N_1345);
nand U2297 (N_2297,N_1999,N_1892);
or U2298 (N_2298,N_1662,N_1101);
and U2299 (N_2299,N_1043,N_1313);
or U2300 (N_2300,N_1897,N_1122);
and U2301 (N_2301,N_1855,N_1538);
nand U2302 (N_2302,N_1598,N_1176);
nand U2303 (N_2303,N_1915,N_1268);
xnor U2304 (N_2304,N_1949,N_1536);
nor U2305 (N_2305,N_1459,N_1376);
nand U2306 (N_2306,N_1982,N_1581);
and U2307 (N_2307,N_1776,N_1157);
and U2308 (N_2308,N_1531,N_1273);
or U2309 (N_2309,N_1278,N_1287);
nand U2310 (N_2310,N_1991,N_1566);
nand U2311 (N_2311,N_1567,N_1896);
or U2312 (N_2312,N_1713,N_1803);
nand U2313 (N_2313,N_1547,N_1825);
xnor U2314 (N_2314,N_1411,N_1871);
nor U2315 (N_2315,N_1513,N_1887);
or U2316 (N_2316,N_1593,N_1326);
or U2317 (N_2317,N_1370,N_1773);
nor U2318 (N_2318,N_1589,N_1905);
and U2319 (N_2319,N_1668,N_1457);
or U2320 (N_2320,N_1543,N_1521);
nor U2321 (N_2321,N_1754,N_1215);
and U2322 (N_2322,N_1473,N_1506);
xor U2323 (N_2323,N_1341,N_1316);
nand U2324 (N_2324,N_1527,N_1353);
and U2325 (N_2325,N_1681,N_1462);
nor U2326 (N_2326,N_1412,N_1481);
nand U2327 (N_2327,N_1767,N_1907);
or U2328 (N_2328,N_1928,N_1138);
nor U2329 (N_2329,N_1494,N_1866);
or U2330 (N_2330,N_1227,N_1339);
and U2331 (N_2331,N_1847,N_1913);
xnor U2332 (N_2332,N_1592,N_1134);
nor U2333 (N_2333,N_1635,N_1349);
or U2334 (N_2334,N_1419,N_1993);
or U2335 (N_2335,N_1150,N_1945);
nand U2336 (N_2336,N_1946,N_1028);
nand U2337 (N_2337,N_1683,N_1178);
nor U2338 (N_2338,N_1805,N_1087);
nor U2339 (N_2339,N_1366,N_1377);
or U2340 (N_2340,N_1470,N_1856);
nor U2341 (N_2341,N_1321,N_1785);
and U2342 (N_2342,N_1880,N_1846);
or U2343 (N_2343,N_1617,N_1793);
nand U2344 (N_2344,N_1404,N_1051);
xnor U2345 (N_2345,N_1799,N_1807);
and U2346 (N_2346,N_1721,N_1013);
nor U2347 (N_2347,N_1772,N_1204);
nand U2348 (N_2348,N_1291,N_1336);
and U2349 (N_2349,N_1818,N_1678);
or U2350 (N_2350,N_1741,N_1166);
nor U2351 (N_2351,N_1367,N_1483);
and U2352 (N_2352,N_1703,N_1707);
nor U2353 (N_2353,N_1399,N_1408);
nor U2354 (N_2354,N_1233,N_1254);
nand U2355 (N_2355,N_1560,N_1511);
nor U2356 (N_2356,N_1822,N_1815);
xnor U2357 (N_2357,N_1573,N_1633);
nand U2358 (N_2358,N_1886,N_1934);
nand U2359 (N_2359,N_1837,N_1059);
or U2360 (N_2360,N_1801,N_1890);
nand U2361 (N_2361,N_1604,N_1235);
or U2362 (N_2362,N_1430,N_1656);
nor U2363 (N_2363,N_1119,N_1014);
xnor U2364 (N_2364,N_1750,N_1838);
and U2365 (N_2365,N_1735,N_1580);
or U2366 (N_2366,N_1571,N_1182);
nand U2367 (N_2367,N_1724,N_1142);
nor U2368 (N_2368,N_1331,N_1712);
nor U2369 (N_2369,N_1653,N_1185);
and U2370 (N_2370,N_1154,N_1975);
xnor U2371 (N_2371,N_1954,N_1241);
xor U2372 (N_2372,N_1594,N_1183);
xor U2373 (N_2373,N_1623,N_1570);
and U2374 (N_2374,N_1015,N_1872);
xor U2375 (N_2375,N_1455,N_1213);
xor U2376 (N_2376,N_1195,N_1486);
nor U2377 (N_2377,N_1800,N_1040);
xor U2378 (N_2378,N_1300,N_1262);
or U2379 (N_2379,N_1851,N_1556);
nand U2380 (N_2380,N_1706,N_1601);
xor U2381 (N_2381,N_1038,N_1747);
and U2382 (N_2382,N_1654,N_1354);
xor U2383 (N_2383,N_1529,N_1076);
nand U2384 (N_2384,N_1583,N_1064);
nand U2385 (N_2385,N_1574,N_1852);
nor U2386 (N_2386,N_1110,N_1789);
nor U2387 (N_2387,N_1414,N_1778);
nor U2388 (N_2388,N_1065,N_1988);
xnor U2389 (N_2389,N_1061,N_1659);
nor U2390 (N_2390,N_1260,N_1226);
xnor U2391 (N_2391,N_1548,N_1285);
or U2392 (N_2392,N_1738,N_1996);
and U2393 (N_2393,N_1202,N_1921);
or U2394 (N_2394,N_1680,N_1493);
and U2395 (N_2395,N_1025,N_1184);
or U2396 (N_2396,N_1239,N_1824);
xor U2397 (N_2397,N_1017,N_1441);
and U2398 (N_2398,N_1171,N_1758);
nand U2399 (N_2399,N_1253,N_1641);
xnor U2400 (N_2400,N_1350,N_1068);
nand U2401 (N_2401,N_1770,N_1908);
nand U2402 (N_2402,N_1899,N_1402);
or U2403 (N_2403,N_1705,N_1796);
xnor U2404 (N_2404,N_1727,N_1693);
nand U2405 (N_2405,N_1347,N_1528);
xnor U2406 (N_2406,N_1378,N_1127);
and U2407 (N_2407,N_1351,N_1534);
nand U2408 (N_2408,N_1279,N_1729);
nor U2409 (N_2409,N_1939,N_1894);
xor U2410 (N_2410,N_1479,N_1901);
nand U2411 (N_2411,N_1055,N_1380);
and U2412 (N_2412,N_1783,N_1876);
nand U2413 (N_2413,N_1830,N_1835);
or U2414 (N_2414,N_1904,N_1515);
and U2415 (N_2415,N_1676,N_1327);
or U2416 (N_2416,N_1214,N_1658);
or U2417 (N_2417,N_1958,N_1120);
and U2418 (N_2418,N_1117,N_1903);
xnor U2419 (N_2419,N_1280,N_1187);
or U2420 (N_2420,N_1143,N_1407);
nand U2421 (N_2421,N_1755,N_1736);
xor U2422 (N_2422,N_1879,N_1492);
or U2423 (N_2423,N_1746,N_1568);
nand U2424 (N_2424,N_1477,N_1011);
and U2425 (N_2425,N_1067,N_1242);
xnor U2426 (N_2426,N_1540,N_1535);
nor U2427 (N_2427,N_1434,N_1208);
nand U2428 (N_2428,N_1298,N_1636);
and U2429 (N_2429,N_1201,N_1200);
or U2430 (N_2430,N_1394,N_1329);
nand U2431 (N_2431,N_1888,N_1424);
nand U2432 (N_2432,N_1172,N_1335);
nand U2433 (N_2433,N_1383,N_1509);
nor U2434 (N_2434,N_1475,N_1842);
xnor U2435 (N_2435,N_1433,N_1125);
and U2436 (N_2436,N_1006,N_1099);
nand U2437 (N_2437,N_1965,N_1760);
and U2438 (N_2438,N_1643,N_1238);
nor U2439 (N_2439,N_1742,N_1487);
xor U2440 (N_2440,N_1505,N_1113);
and U2441 (N_2441,N_1661,N_1361);
nand U2442 (N_2442,N_1416,N_1009);
nand U2443 (N_2443,N_1638,N_1610);
and U2444 (N_2444,N_1929,N_1931);
nor U2445 (N_2445,N_1160,N_1315);
and U2446 (N_2446,N_1140,N_1840);
or U2447 (N_2447,N_1449,N_1501);
xnor U2448 (N_2448,N_1070,N_1660);
xnor U2449 (N_2449,N_1203,N_1276);
nor U2450 (N_2450,N_1251,N_1312);
nor U2451 (N_2451,N_1175,N_1582);
and U2452 (N_2452,N_1275,N_1228);
nand U2453 (N_2453,N_1447,N_1466);
nor U2454 (N_2454,N_1629,N_1960);
nand U2455 (N_2455,N_1551,N_1977);
nand U2456 (N_2456,N_1577,N_1450);
and U2457 (N_2457,N_1274,N_1726);
nand U2458 (N_2458,N_1474,N_1974);
and U2459 (N_2459,N_1702,N_1523);
or U2460 (N_2460,N_1520,N_1149);
nor U2461 (N_2461,N_1698,N_1256);
xor U2462 (N_2462,N_1405,N_1627);
or U2463 (N_2463,N_1938,N_1491);
nor U2464 (N_2464,N_1116,N_1968);
and U2465 (N_2465,N_1664,N_1655);
or U2466 (N_2466,N_1585,N_1194);
or U2467 (N_2467,N_1950,N_1955);
xor U2468 (N_2468,N_1343,N_1324);
nand U2469 (N_2469,N_1769,N_1749);
nor U2470 (N_2470,N_1731,N_1836);
nand U2471 (N_2471,N_1802,N_1951);
nand U2472 (N_2472,N_1482,N_1539);
and U2473 (N_2473,N_1910,N_1115);
nand U2474 (N_2474,N_1118,N_1973);
xnor U2475 (N_2475,N_1136,N_1308);
xnor U2476 (N_2476,N_1250,N_1677);
nor U2477 (N_2477,N_1717,N_1508);
nor U2478 (N_2478,N_1139,N_1828);
or U2479 (N_2479,N_1409,N_1984);
and U2480 (N_2480,N_1864,N_1078);
nor U2481 (N_2481,N_1672,N_1392);
and U2482 (N_2482,N_1986,N_1809);
or U2483 (N_2483,N_1484,N_1058);
xor U2484 (N_2484,N_1294,N_1458);
or U2485 (N_2485,N_1980,N_1144);
or U2486 (N_2486,N_1320,N_1196);
or U2487 (N_2487,N_1794,N_1277);
nor U2488 (N_2488,N_1170,N_1669);
or U2489 (N_2489,N_1550,N_1400);
nand U2490 (N_2490,N_1781,N_1289);
nand U2491 (N_2491,N_1944,N_1671);
nor U2492 (N_2492,N_1826,N_1792);
nand U2493 (N_2493,N_1418,N_1063);
xor U2494 (N_2494,N_1665,N_1590);
and U2495 (N_2495,N_1821,N_1563);
nor U2496 (N_2496,N_1100,N_1976);
xnor U2497 (N_2497,N_1179,N_1284);
or U2498 (N_2498,N_1752,N_1844);
xnor U2499 (N_2499,N_1881,N_1865);
nand U2500 (N_2500,N_1008,N_1365);
or U2501 (N_2501,N_1929,N_1584);
nor U2502 (N_2502,N_1938,N_1948);
nor U2503 (N_2503,N_1638,N_1607);
nor U2504 (N_2504,N_1633,N_1034);
or U2505 (N_2505,N_1843,N_1663);
xnor U2506 (N_2506,N_1722,N_1623);
xor U2507 (N_2507,N_1046,N_1616);
xnor U2508 (N_2508,N_1552,N_1958);
and U2509 (N_2509,N_1933,N_1213);
xor U2510 (N_2510,N_1770,N_1947);
nor U2511 (N_2511,N_1423,N_1728);
xor U2512 (N_2512,N_1238,N_1151);
and U2513 (N_2513,N_1845,N_1718);
xor U2514 (N_2514,N_1017,N_1478);
and U2515 (N_2515,N_1395,N_1849);
nand U2516 (N_2516,N_1875,N_1719);
xor U2517 (N_2517,N_1900,N_1360);
xor U2518 (N_2518,N_1585,N_1092);
and U2519 (N_2519,N_1045,N_1048);
nand U2520 (N_2520,N_1393,N_1425);
or U2521 (N_2521,N_1258,N_1105);
and U2522 (N_2522,N_1001,N_1963);
xnor U2523 (N_2523,N_1786,N_1395);
and U2524 (N_2524,N_1641,N_1194);
xnor U2525 (N_2525,N_1240,N_1027);
xnor U2526 (N_2526,N_1429,N_1481);
or U2527 (N_2527,N_1550,N_1719);
and U2528 (N_2528,N_1702,N_1313);
nor U2529 (N_2529,N_1259,N_1806);
nand U2530 (N_2530,N_1573,N_1542);
nor U2531 (N_2531,N_1523,N_1698);
nor U2532 (N_2532,N_1546,N_1394);
xnor U2533 (N_2533,N_1163,N_1609);
nor U2534 (N_2534,N_1885,N_1162);
or U2535 (N_2535,N_1022,N_1696);
and U2536 (N_2536,N_1525,N_1794);
or U2537 (N_2537,N_1656,N_1369);
nand U2538 (N_2538,N_1438,N_1098);
nor U2539 (N_2539,N_1127,N_1979);
nand U2540 (N_2540,N_1515,N_1741);
nor U2541 (N_2541,N_1710,N_1887);
nand U2542 (N_2542,N_1665,N_1935);
xnor U2543 (N_2543,N_1261,N_1578);
or U2544 (N_2544,N_1024,N_1157);
nand U2545 (N_2545,N_1145,N_1497);
nor U2546 (N_2546,N_1383,N_1145);
xor U2547 (N_2547,N_1620,N_1308);
nor U2548 (N_2548,N_1324,N_1239);
or U2549 (N_2549,N_1833,N_1163);
xor U2550 (N_2550,N_1867,N_1765);
xor U2551 (N_2551,N_1148,N_1057);
nand U2552 (N_2552,N_1240,N_1910);
xor U2553 (N_2553,N_1655,N_1377);
nor U2554 (N_2554,N_1950,N_1322);
nor U2555 (N_2555,N_1575,N_1588);
nor U2556 (N_2556,N_1739,N_1674);
nor U2557 (N_2557,N_1593,N_1492);
nor U2558 (N_2558,N_1419,N_1366);
and U2559 (N_2559,N_1628,N_1972);
xor U2560 (N_2560,N_1031,N_1322);
or U2561 (N_2561,N_1297,N_1032);
nand U2562 (N_2562,N_1391,N_1640);
or U2563 (N_2563,N_1641,N_1735);
nor U2564 (N_2564,N_1614,N_1560);
nand U2565 (N_2565,N_1040,N_1638);
nor U2566 (N_2566,N_1252,N_1605);
or U2567 (N_2567,N_1110,N_1400);
nand U2568 (N_2568,N_1756,N_1111);
nor U2569 (N_2569,N_1198,N_1338);
or U2570 (N_2570,N_1659,N_1448);
nand U2571 (N_2571,N_1669,N_1495);
nor U2572 (N_2572,N_1093,N_1805);
and U2573 (N_2573,N_1962,N_1169);
and U2574 (N_2574,N_1345,N_1763);
and U2575 (N_2575,N_1140,N_1477);
nand U2576 (N_2576,N_1935,N_1640);
nand U2577 (N_2577,N_1907,N_1899);
or U2578 (N_2578,N_1217,N_1743);
or U2579 (N_2579,N_1949,N_1385);
xnor U2580 (N_2580,N_1620,N_1285);
and U2581 (N_2581,N_1603,N_1893);
or U2582 (N_2582,N_1386,N_1073);
and U2583 (N_2583,N_1161,N_1360);
and U2584 (N_2584,N_1440,N_1066);
or U2585 (N_2585,N_1560,N_1218);
nor U2586 (N_2586,N_1238,N_1147);
nand U2587 (N_2587,N_1178,N_1433);
nand U2588 (N_2588,N_1203,N_1637);
and U2589 (N_2589,N_1990,N_1041);
or U2590 (N_2590,N_1601,N_1320);
xor U2591 (N_2591,N_1877,N_1871);
or U2592 (N_2592,N_1070,N_1254);
nor U2593 (N_2593,N_1240,N_1185);
or U2594 (N_2594,N_1613,N_1629);
nor U2595 (N_2595,N_1701,N_1097);
nand U2596 (N_2596,N_1244,N_1875);
and U2597 (N_2597,N_1627,N_1674);
nand U2598 (N_2598,N_1664,N_1649);
nand U2599 (N_2599,N_1849,N_1365);
nor U2600 (N_2600,N_1311,N_1110);
xnor U2601 (N_2601,N_1084,N_1351);
xnor U2602 (N_2602,N_1718,N_1395);
nor U2603 (N_2603,N_1935,N_1195);
nor U2604 (N_2604,N_1740,N_1542);
and U2605 (N_2605,N_1946,N_1436);
and U2606 (N_2606,N_1215,N_1506);
xnor U2607 (N_2607,N_1583,N_1984);
or U2608 (N_2608,N_1265,N_1985);
xnor U2609 (N_2609,N_1451,N_1746);
and U2610 (N_2610,N_1441,N_1572);
and U2611 (N_2611,N_1091,N_1341);
and U2612 (N_2612,N_1111,N_1401);
xor U2613 (N_2613,N_1716,N_1095);
and U2614 (N_2614,N_1817,N_1922);
or U2615 (N_2615,N_1780,N_1779);
nand U2616 (N_2616,N_1105,N_1359);
nand U2617 (N_2617,N_1517,N_1335);
xor U2618 (N_2618,N_1568,N_1935);
or U2619 (N_2619,N_1715,N_1403);
nor U2620 (N_2620,N_1865,N_1541);
nand U2621 (N_2621,N_1072,N_1710);
xnor U2622 (N_2622,N_1547,N_1065);
xnor U2623 (N_2623,N_1464,N_1582);
and U2624 (N_2624,N_1410,N_1520);
or U2625 (N_2625,N_1219,N_1757);
nand U2626 (N_2626,N_1376,N_1400);
xor U2627 (N_2627,N_1468,N_1302);
nor U2628 (N_2628,N_1210,N_1625);
xnor U2629 (N_2629,N_1945,N_1051);
xnor U2630 (N_2630,N_1518,N_1029);
xnor U2631 (N_2631,N_1598,N_1923);
nor U2632 (N_2632,N_1477,N_1082);
xor U2633 (N_2633,N_1629,N_1029);
xnor U2634 (N_2634,N_1136,N_1245);
nand U2635 (N_2635,N_1400,N_1042);
nor U2636 (N_2636,N_1718,N_1531);
and U2637 (N_2637,N_1582,N_1390);
nor U2638 (N_2638,N_1190,N_1586);
nand U2639 (N_2639,N_1156,N_1723);
nand U2640 (N_2640,N_1058,N_1468);
nand U2641 (N_2641,N_1430,N_1648);
xor U2642 (N_2642,N_1131,N_1838);
xnor U2643 (N_2643,N_1294,N_1197);
nor U2644 (N_2644,N_1234,N_1297);
or U2645 (N_2645,N_1288,N_1323);
and U2646 (N_2646,N_1323,N_1339);
or U2647 (N_2647,N_1052,N_1939);
nand U2648 (N_2648,N_1033,N_1506);
and U2649 (N_2649,N_1838,N_1674);
xor U2650 (N_2650,N_1186,N_1077);
nor U2651 (N_2651,N_1177,N_1067);
and U2652 (N_2652,N_1174,N_1444);
xor U2653 (N_2653,N_1887,N_1118);
nor U2654 (N_2654,N_1668,N_1311);
nor U2655 (N_2655,N_1602,N_1296);
nor U2656 (N_2656,N_1337,N_1435);
and U2657 (N_2657,N_1878,N_1100);
or U2658 (N_2658,N_1093,N_1185);
or U2659 (N_2659,N_1326,N_1972);
nor U2660 (N_2660,N_1569,N_1296);
nor U2661 (N_2661,N_1072,N_1830);
nand U2662 (N_2662,N_1201,N_1298);
or U2663 (N_2663,N_1000,N_1013);
nand U2664 (N_2664,N_1479,N_1578);
or U2665 (N_2665,N_1874,N_1295);
nand U2666 (N_2666,N_1024,N_1272);
nand U2667 (N_2667,N_1894,N_1918);
or U2668 (N_2668,N_1491,N_1840);
xor U2669 (N_2669,N_1293,N_1614);
xnor U2670 (N_2670,N_1557,N_1380);
and U2671 (N_2671,N_1050,N_1021);
or U2672 (N_2672,N_1384,N_1186);
or U2673 (N_2673,N_1944,N_1877);
and U2674 (N_2674,N_1410,N_1015);
nand U2675 (N_2675,N_1718,N_1191);
xor U2676 (N_2676,N_1631,N_1531);
xor U2677 (N_2677,N_1968,N_1807);
nand U2678 (N_2678,N_1594,N_1510);
nor U2679 (N_2679,N_1297,N_1394);
nand U2680 (N_2680,N_1884,N_1471);
nand U2681 (N_2681,N_1601,N_1764);
nor U2682 (N_2682,N_1003,N_1009);
nand U2683 (N_2683,N_1314,N_1794);
xnor U2684 (N_2684,N_1915,N_1187);
nor U2685 (N_2685,N_1520,N_1236);
xor U2686 (N_2686,N_1357,N_1836);
xnor U2687 (N_2687,N_1624,N_1501);
xnor U2688 (N_2688,N_1066,N_1766);
xor U2689 (N_2689,N_1434,N_1972);
and U2690 (N_2690,N_1025,N_1345);
xor U2691 (N_2691,N_1007,N_1607);
and U2692 (N_2692,N_1050,N_1789);
xnor U2693 (N_2693,N_1286,N_1498);
nand U2694 (N_2694,N_1128,N_1746);
or U2695 (N_2695,N_1110,N_1198);
and U2696 (N_2696,N_1515,N_1791);
xor U2697 (N_2697,N_1217,N_1588);
and U2698 (N_2698,N_1369,N_1723);
nand U2699 (N_2699,N_1208,N_1731);
xor U2700 (N_2700,N_1142,N_1095);
xnor U2701 (N_2701,N_1429,N_1890);
and U2702 (N_2702,N_1425,N_1810);
xnor U2703 (N_2703,N_1428,N_1106);
and U2704 (N_2704,N_1336,N_1016);
xor U2705 (N_2705,N_1623,N_1717);
nand U2706 (N_2706,N_1197,N_1366);
and U2707 (N_2707,N_1704,N_1418);
or U2708 (N_2708,N_1345,N_1097);
and U2709 (N_2709,N_1426,N_1409);
xor U2710 (N_2710,N_1769,N_1730);
nor U2711 (N_2711,N_1850,N_1287);
and U2712 (N_2712,N_1737,N_1689);
nor U2713 (N_2713,N_1892,N_1219);
nand U2714 (N_2714,N_1634,N_1875);
or U2715 (N_2715,N_1318,N_1363);
or U2716 (N_2716,N_1019,N_1813);
xor U2717 (N_2717,N_1766,N_1820);
nor U2718 (N_2718,N_1151,N_1380);
nor U2719 (N_2719,N_1582,N_1627);
or U2720 (N_2720,N_1311,N_1930);
and U2721 (N_2721,N_1075,N_1828);
xnor U2722 (N_2722,N_1443,N_1800);
nand U2723 (N_2723,N_1058,N_1443);
nand U2724 (N_2724,N_1280,N_1408);
nor U2725 (N_2725,N_1877,N_1979);
xnor U2726 (N_2726,N_1913,N_1356);
and U2727 (N_2727,N_1666,N_1099);
nand U2728 (N_2728,N_1506,N_1245);
xor U2729 (N_2729,N_1116,N_1085);
and U2730 (N_2730,N_1756,N_1449);
xor U2731 (N_2731,N_1917,N_1806);
nand U2732 (N_2732,N_1485,N_1087);
or U2733 (N_2733,N_1813,N_1614);
nand U2734 (N_2734,N_1620,N_1877);
and U2735 (N_2735,N_1467,N_1846);
xnor U2736 (N_2736,N_1636,N_1389);
nor U2737 (N_2737,N_1265,N_1850);
xnor U2738 (N_2738,N_1632,N_1340);
xor U2739 (N_2739,N_1144,N_1360);
nor U2740 (N_2740,N_1535,N_1215);
nor U2741 (N_2741,N_1177,N_1476);
nand U2742 (N_2742,N_1217,N_1079);
xor U2743 (N_2743,N_1932,N_1017);
and U2744 (N_2744,N_1285,N_1254);
xnor U2745 (N_2745,N_1224,N_1334);
nor U2746 (N_2746,N_1720,N_1987);
xnor U2747 (N_2747,N_1177,N_1520);
and U2748 (N_2748,N_1946,N_1601);
xnor U2749 (N_2749,N_1014,N_1938);
nor U2750 (N_2750,N_1733,N_1891);
xnor U2751 (N_2751,N_1524,N_1036);
and U2752 (N_2752,N_1335,N_1898);
xnor U2753 (N_2753,N_1268,N_1991);
nor U2754 (N_2754,N_1049,N_1829);
and U2755 (N_2755,N_1326,N_1513);
nor U2756 (N_2756,N_1697,N_1189);
or U2757 (N_2757,N_1926,N_1064);
and U2758 (N_2758,N_1027,N_1270);
nand U2759 (N_2759,N_1482,N_1584);
xor U2760 (N_2760,N_1357,N_1707);
xnor U2761 (N_2761,N_1861,N_1378);
xnor U2762 (N_2762,N_1997,N_1497);
and U2763 (N_2763,N_1726,N_1470);
nor U2764 (N_2764,N_1118,N_1134);
nand U2765 (N_2765,N_1618,N_1057);
xnor U2766 (N_2766,N_1031,N_1658);
or U2767 (N_2767,N_1279,N_1252);
or U2768 (N_2768,N_1883,N_1815);
nand U2769 (N_2769,N_1630,N_1503);
nor U2770 (N_2770,N_1785,N_1986);
xnor U2771 (N_2771,N_1789,N_1735);
nor U2772 (N_2772,N_1055,N_1585);
nand U2773 (N_2773,N_1865,N_1803);
xor U2774 (N_2774,N_1528,N_1376);
xnor U2775 (N_2775,N_1811,N_1453);
and U2776 (N_2776,N_1579,N_1419);
nand U2777 (N_2777,N_1282,N_1484);
nor U2778 (N_2778,N_1713,N_1489);
nor U2779 (N_2779,N_1430,N_1493);
xnor U2780 (N_2780,N_1501,N_1253);
nand U2781 (N_2781,N_1695,N_1509);
and U2782 (N_2782,N_1571,N_1712);
nor U2783 (N_2783,N_1686,N_1512);
or U2784 (N_2784,N_1050,N_1076);
nor U2785 (N_2785,N_1808,N_1850);
and U2786 (N_2786,N_1066,N_1505);
xnor U2787 (N_2787,N_1336,N_1320);
nor U2788 (N_2788,N_1879,N_1826);
or U2789 (N_2789,N_1694,N_1193);
or U2790 (N_2790,N_1932,N_1919);
nand U2791 (N_2791,N_1944,N_1855);
or U2792 (N_2792,N_1952,N_1117);
and U2793 (N_2793,N_1760,N_1715);
xor U2794 (N_2794,N_1842,N_1894);
nand U2795 (N_2795,N_1362,N_1934);
xnor U2796 (N_2796,N_1074,N_1016);
xor U2797 (N_2797,N_1549,N_1699);
xnor U2798 (N_2798,N_1919,N_1245);
nor U2799 (N_2799,N_1089,N_1270);
or U2800 (N_2800,N_1406,N_1086);
xor U2801 (N_2801,N_1563,N_1829);
nand U2802 (N_2802,N_1284,N_1787);
nand U2803 (N_2803,N_1553,N_1755);
nor U2804 (N_2804,N_1098,N_1626);
xor U2805 (N_2805,N_1393,N_1033);
xor U2806 (N_2806,N_1238,N_1919);
or U2807 (N_2807,N_1409,N_1016);
nand U2808 (N_2808,N_1860,N_1362);
nand U2809 (N_2809,N_1182,N_1673);
nand U2810 (N_2810,N_1136,N_1602);
nor U2811 (N_2811,N_1905,N_1472);
nand U2812 (N_2812,N_1836,N_1749);
nand U2813 (N_2813,N_1290,N_1012);
or U2814 (N_2814,N_1493,N_1066);
or U2815 (N_2815,N_1996,N_1074);
and U2816 (N_2816,N_1369,N_1547);
xor U2817 (N_2817,N_1608,N_1805);
and U2818 (N_2818,N_1993,N_1258);
nor U2819 (N_2819,N_1996,N_1545);
and U2820 (N_2820,N_1259,N_1998);
xnor U2821 (N_2821,N_1803,N_1816);
or U2822 (N_2822,N_1642,N_1621);
or U2823 (N_2823,N_1953,N_1013);
or U2824 (N_2824,N_1795,N_1563);
nor U2825 (N_2825,N_1542,N_1719);
or U2826 (N_2826,N_1964,N_1619);
nand U2827 (N_2827,N_1849,N_1699);
and U2828 (N_2828,N_1936,N_1194);
nor U2829 (N_2829,N_1516,N_1773);
and U2830 (N_2830,N_1582,N_1973);
nand U2831 (N_2831,N_1521,N_1297);
nand U2832 (N_2832,N_1380,N_1372);
xor U2833 (N_2833,N_1623,N_1134);
and U2834 (N_2834,N_1944,N_1218);
and U2835 (N_2835,N_1083,N_1667);
nor U2836 (N_2836,N_1784,N_1808);
or U2837 (N_2837,N_1990,N_1410);
or U2838 (N_2838,N_1708,N_1042);
nand U2839 (N_2839,N_1367,N_1030);
xnor U2840 (N_2840,N_1958,N_1103);
and U2841 (N_2841,N_1875,N_1960);
nor U2842 (N_2842,N_1333,N_1470);
nand U2843 (N_2843,N_1177,N_1293);
nand U2844 (N_2844,N_1302,N_1836);
xnor U2845 (N_2845,N_1871,N_1047);
or U2846 (N_2846,N_1011,N_1049);
nand U2847 (N_2847,N_1559,N_1187);
or U2848 (N_2848,N_1681,N_1828);
or U2849 (N_2849,N_1562,N_1696);
and U2850 (N_2850,N_1148,N_1549);
and U2851 (N_2851,N_1546,N_1516);
nand U2852 (N_2852,N_1941,N_1160);
xnor U2853 (N_2853,N_1700,N_1581);
nor U2854 (N_2854,N_1578,N_1951);
and U2855 (N_2855,N_1950,N_1181);
nand U2856 (N_2856,N_1037,N_1473);
nand U2857 (N_2857,N_1346,N_1003);
xor U2858 (N_2858,N_1495,N_1433);
or U2859 (N_2859,N_1312,N_1726);
nor U2860 (N_2860,N_1643,N_1333);
nand U2861 (N_2861,N_1372,N_1277);
or U2862 (N_2862,N_1572,N_1946);
xor U2863 (N_2863,N_1450,N_1293);
nor U2864 (N_2864,N_1517,N_1519);
and U2865 (N_2865,N_1369,N_1349);
or U2866 (N_2866,N_1684,N_1250);
nor U2867 (N_2867,N_1388,N_1683);
or U2868 (N_2868,N_1158,N_1363);
nand U2869 (N_2869,N_1644,N_1076);
xnor U2870 (N_2870,N_1897,N_1530);
or U2871 (N_2871,N_1790,N_1481);
and U2872 (N_2872,N_1417,N_1361);
nor U2873 (N_2873,N_1827,N_1001);
nor U2874 (N_2874,N_1969,N_1725);
nand U2875 (N_2875,N_1954,N_1681);
nand U2876 (N_2876,N_1611,N_1243);
and U2877 (N_2877,N_1670,N_1804);
nand U2878 (N_2878,N_1649,N_1932);
xor U2879 (N_2879,N_1047,N_1605);
xnor U2880 (N_2880,N_1637,N_1466);
xor U2881 (N_2881,N_1585,N_1175);
nor U2882 (N_2882,N_1016,N_1230);
nor U2883 (N_2883,N_1948,N_1687);
or U2884 (N_2884,N_1851,N_1452);
nand U2885 (N_2885,N_1336,N_1844);
or U2886 (N_2886,N_1408,N_1387);
nand U2887 (N_2887,N_1334,N_1011);
xnor U2888 (N_2888,N_1356,N_1393);
xnor U2889 (N_2889,N_1183,N_1314);
and U2890 (N_2890,N_1743,N_1434);
and U2891 (N_2891,N_1047,N_1761);
or U2892 (N_2892,N_1709,N_1578);
and U2893 (N_2893,N_1350,N_1648);
xnor U2894 (N_2894,N_1078,N_1715);
nand U2895 (N_2895,N_1088,N_1372);
or U2896 (N_2896,N_1419,N_1094);
xor U2897 (N_2897,N_1122,N_1412);
and U2898 (N_2898,N_1881,N_1366);
nor U2899 (N_2899,N_1692,N_1985);
nand U2900 (N_2900,N_1240,N_1671);
or U2901 (N_2901,N_1336,N_1279);
nand U2902 (N_2902,N_1835,N_1038);
nor U2903 (N_2903,N_1814,N_1714);
nand U2904 (N_2904,N_1760,N_1311);
xor U2905 (N_2905,N_1732,N_1195);
or U2906 (N_2906,N_1590,N_1821);
and U2907 (N_2907,N_1190,N_1899);
or U2908 (N_2908,N_1736,N_1023);
and U2909 (N_2909,N_1810,N_1305);
or U2910 (N_2910,N_1225,N_1464);
nor U2911 (N_2911,N_1806,N_1196);
xor U2912 (N_2912,N_1107,N_1055);
nor U2913 (N_2913,N_1018,N_1046);
xor U2914 (N_2914,N_1447,N_1362);
xor U2915 (N_2915,N_1733,N_1605);
xor U2916 (N_2916,N_1032,N_1053);
and U2917 (N_2917,N_1851,N_1615);
nor U2918 (N_2918,N_1390,N_1126);
or U2919 (N_2919,N_1563,N_1186);
or U2920 (N_2920,N_1657,N_1117);
or U2921 (N_2921,N_1435,N_1096);
nor U2922 (N_2922,N_1872,N_1833);
nand U2923 (N_2923,N_1011,N_1439);
or U2924 (N_2924,N_1529,N_1446);
xnor U2925 (N_2925,N_1342,N_1456);
nor U2926 (N_2926,N_1902,N_1840);
and U2927 (N_2927,N_1514,N_1873);
nand U2928 (N_2928,N_1119,N_1430);
nand U2929 (N_2929,N_1387,N_1497);
xor U2930 (N_2930,N_1105,N_1248);
and U2931 (N_2931,N_1651,N_1317);
nand U2932 (N_2932,N_1628,N_1858);
xor U2933 (N_2933,N_1539,N_1383);
and U2934 (N_2934,N_1437,N_1831);
nand U2935 (N_2935,N_1877,N_1748);
nor U2936 (N_2936,N_1876,N_1808);
xnor U2937 (N_2937,N_1350,N_1304);
nor U2938 (N_2938,N_1910,N_1981);
nor U2939 (N_2939,N_1928,N_1383);
and U2940 (N_2940,N_1033,N_1585);
nand U2941 (N_2941,N_1240,N_1664);
xnor U2942 (N_2942,N_1548,N_1237);
and U2943 (N_2943,N_1070,N_1037);
nand U2944 (N_2944,N_1403,N_1630);
or U2945 (N_2945,N_1608,N_1466);
xnor U2946 (N_2946,N_1483,N_1311);
or U2947 (N_2947,N_1580,N_1238);
nand U2948 (N_2948,N_1214,N_1487);
nand U2949 (N_2949,N_1331,N_1467);
nor U2950 (N_2950,N_1408,N_1237);
nor U2951 (N_2951,N_1526,N_1947);
nor U2952 (N_2952,N_1740,N_1951);
nand U2953 (N_2953,N_1179,N_1865);
nand U2954 (N_2954,N_1774,N_1461);
or U2955 (N_2955,N_1970,N_1949);
or U2956 (N_2956,N_1218,N_1166);
nor U2957 (N_2957,N_1552,N_1345);
xor U2958 (N_2958,N_1812,N_1021);
nor U2959 (N_2959,N_1202,N_1701);
or U2960 (N_2960,N_1430,N_1440);
xnor U2961 (N_2961,N_1679,N_1048);
xnor U2962 (N_2962,N_1847,N_1932);
and U2963 (N_2963,N_1872,N_1032);
or U2964 (N_2964,N_1339,N_1855);
or U2965 (N_2965,N_1418,N_1327);
or U2966 (N_2966,N_1645,N_1411);
xor U2967 (N_2967,N_1895,N_1047);
and U2968 (N_2968,N_1294,N_1887);
nand U2969 (N_2969,N_1477,N_1986);
nor U2970 (N_2970,N_1237,N_1323);
and U2971 (N_2971,N_1566,N_1709);
nand U2972 (N_2972,N_1728,N_1780);
nor U2973 (N_2973,N_1906,N_1972);
nor U2974 (N_2974,N_1611,N_1499);
nand U2975 (N_2975,N_1835,N_1455);
and U2976 (N_2976,N_1644,N_1757);
xnor U2977 (N_2977,N_1602,N_1093);
and U2978 (N_2978,N_1313,N_1620);
nand U2979 (N_2979,N_1241,N_1352);
nor U2980 (N_2980,N_1400,N_1187);
nor U2981 (N_2981,N_1424,N_1573);
and U2982 (N_2982,N_1296,N_1836);
and U2983 (N_2983,N_1766,N_1366);
nand U2984 (N_2984,N_1412,N_1917);
or U2985 (N_2985,N_1592,N_1049);
nand U2986 (N_2986,N_1665,N_1999);
or U2987 (N_2987,N_1674,N_1437);
nor U2988 (N_2988,N_1540,N_1497);
and U2989 (N_2989,N_1137,N_1840);
nor U2990 (N_2990,N_1752,N_1026);
xor U2991 (N_2991,N_1488,N_1895);
and U2992 (N_2992,N_1590,N_1208);
or U2993 (N_2993,N_1296,N_1604);
nand U2994 (N_2994,N_1006,N_1804);
or U2995 (N_2995,N_1856,N_1504);
nor U2996 (N_2996,N_1149,N_1682);
or U2997 (N_2997,N_1863,N_1035);
xnor U2998 (N_2998,N_1838,N_1417);
xnor U2999 (N_2999,N_1336,N_1248);
nand U3000 (N_3000,N_2533,N_2945);
or U3001 (N_3001,N_2279,N_2290);
or U3002 (N_3002,N_2361,N_2814);
and U3003 (N_3003,N_2088,N_2657);
nor U3004 (N_3004,N_2900,N_2033);
nand U3005 (N_3005,N_2451,N_2539);
nor U3006 (N_3006,N_2655,N_2261);
xor U3007 (N_3007,N_2395,N_2706);
nor U3008 (N_3008,N_2422,N_2469);
xor U3009 (N_3009,N_2083,N_2488);
and U3010 (N_3010,N_2891,N_2623);
and U3011 (N_3011,N_2330,N_2888);
and U3012 (N_3012,N_2136,N_2140);
nand U3013 (N_3013,N_2271,N_2311);
xnor U3014 (N_3014,N_2421,N_2711);
or U3015 (N_3015,N_2478,N_2955);
nand U3016 (N_3016,N_2739,N_2508);
and U3017 (N_3017,N_2748,N_2081);
or U3018 (N_3018,N_2281,N_2807);
xnor U3019 (N_3019,N_2825,N_2021);
or U3020 (N_3020,N_2650,N_2602);
nor U3021 (N_3021,N_2198,N_2565);
nor U3022 (N_3022,N_2201,N_2598);
or U3023 (N_3023,N_2845,N_2354);
or U3024 (N_3024,N_2284,N_2642);
or U3025 (N_3025,N_2546,N_2663);
xor U3026 (N_3026,N_2087,N_2892);
or U3027 (N_3027,N_2819,N_2157);
xnor U3028 (N_3028,N_2893,N_2069);
xor U3029 (N_3029,N_2728,N_2673);
and U3030 (N_3030,N_2034,N_2832);
nor U3031 (N_3031,N_2454,N_2437);
or U3032 (N_3032,N_2118,N_2744);
and U3033 (N_3033,N_2780,N_2821);
or U3034 (N_3034,N_2643,N_2371);
nand U3035 (N_3035,N_2159,N_2741);
nand U3036 (N_3036,N_2818,N_2192);
or U3037 (N_3037,N_2876,N_2370);
nor U3038 (N_3038,N_2759,N_2023);
nand U3039 (N_3039,N_2869,N_2073);
and U3040 (N_3040,N_2029,N_2683);
or U3041 (N_3041,N_2638,N_2849);
nand U3042 (N_3042,N_2324,N_2144);
or U3043 (N_3043,N_2003,N_2779);
xor U3044 (N_3044,N_2368,N_2274);
and U3045 (N_3045,N_2336,N_2342);
nor U3046 (N_3046,N_2439,N_2054);
or U3047 (N_3047,N_2122,N_2015);
nor U3048 (N_3048,N_2458,N_2681);
xor U3049 (N_3049,N_2002,N_2344);
xor U3050 (N_3050,N_2335,N_2889);
and U3051 (N_3051,N_2640,N_2147);
xnor U3052 (N_3052,N_2108,N_2383);
and U3053 (N_3053,N_2872,N_2696);
xnor U3054 (N_3054,N_2875,N_2751);
nand U3055 (N_3055,N_2106,N_2094);
nor U3056 (N_3056,N_2247,N_2403);
xor U3057 (N_3057,N_2625,N_2090);
nand U3058 (N_3058,N_2408,N_2927);
or U3059 (N_3059,N_2510,N_2704);
and U3060 (N_3060,N_2651,N_2117);
xnor U3061 (N_3061,N_2263,N_2440);
or U3062 (N_3062,N_2115,N_2661);
or U3063 (N_3063,N_2690,N_2841);
nor U3064 (N_3064,N_2262,N_2323);
or U3065 (N_3065,N_2039,N_2639);
and U3066 (N_3066,N_2961,N_2092);
nor U3067 (N_3067,N_2360,N_2205);
nand U3068 (N_3068,N_2647,N_2575);
nor U3069 (N_3069,N_2166,N_2550);
nand U3070 (N_3070,N_2404,N_2163);
and U3071 (N_3071,N_2967,N_2237);
xor U3072 (N_3072,N_2133,N_2098);
nand U3073 (N_3073,N_2297,N_2309);
nor U3074 (N_3074,N_2534,N_2597);
nor U3075 (N_3075,N_2227,N_2037);
and U3076 (N_3076,N_2203,N_2848);
and U3077 (N_3077,N_2386,N_2871);
or U3078 (N_3078,N_2479,N_2540);
nor U3079 (N_3079,N_2399,N_2170);
nor U3080 (N_3080,N_2600,N_2664);
nand U3081 (N_3081,N_2703,N_2836);
and U3082 (N_3082,N_2905,N_2014);
and U3083 (N_3083,N_2606,N_2242);
or U3084 (N_3084,N_2061,N_2005);
nand U3085 (N_3085,N_2352,N_2523);
nand U3086 (N_3086,N_2969,N_2246);
xor U3087 (N_3087,N_2908,N_2200);
nor U3088 (N_3088,N_2020,N_2180);
nand U3089 (N_3089,N_2992,N_2617);
xor U3090 (N_3090,N_2936,N_2607);
xor U3091 (N_3091,N_2929,N_2331);
nor U3092 (N_3092,N_2438,N_2957);
nand U3093 (N_3093,N_2152,N_2394);
and U3094 (N_3094,N_2350,N_2027);
nor U3095 (N_3095,N_2175,N_2940);
xor U3096 (N_3096,N_2149,N_2334);
nor U3097 (N_3097,N_2485,N_2169);
or U3098 (N_3098,N_2858,N_2199);
nand U3099 (N_3099,N_2025,N_2302);
nor U3100 (N_3100,N_2911,N_2578);
nor U3101 (N_3101,N_2505,N_2435);
xor U3102 (N_3102,N_2058,N_2702);
and U3103 (N_3103,N_2884,N_2393);
nor U3104 (N_3104,N_2031,N_2009);
or U3105 (N_3105,N_2328,N_2926);
nand U3106 (N_3106,N_2616,N_2495);
and U3107 (N_3107,N_2068,N_2656);
nor U3108 (N_3108,N_2093,N_2786);
xnor U3109 (N_3109,N_2299,N_2490);
nand U3110 (N_3110,N_2110,N_2229);
nand U3111 (N_3111,N_2486,N_2794);
xnor U3112 (N_3112,N_2298,N_2254);
and U3113 (N_3113,N_2189,N_2579);
and U3114 (N_3114,N_2053,N_2839);
and U3115 (N_3115,N_2462,N_2145);
or U3116 (N_3116,N_2428,N_2275);
nor U3117 (N_3117,N_2179,N_2862);
nand U3118 (N_3118,N_2958,N_2672);
xor U3119 (N_3119,N_2358,N_2436);
xnor U3120 (N_3120,N_2621,N_2007);
nor U3121 (N_3121,N_2662,N_2820);
nor U3122 (N_3122,N_2844,N_2288);
or U3123 (N_3123,N_2494,N_2959);
or U3124 (N_3124,N_2287,N_2218);
or U3125 (N_3125,N_2266,N_2613);
nor U3126 (N_3126,N_2215,N_2563);
nand U3127 (N_3127,N_2585,N_2783);
xnor U3128 (N_3128,N_2817,N_2195);
nand U3129 (N_3129,N_2943,N_2286);
xnor U3130 (N_3130,N_2951,N_2402);
xor U3131 (N_3131,N_2989,N_2172);
xnor U3132 (N_3132,N_2749,N_2592);
or U3133 (N_3133,N_2325,N_2852);
nor U3134 (N_3134,N_2504,N_2968);
xor U3135 (N_3135,N_2292,N_2134);
nor U3136 (N_3136,N_2351,N_2496);
nor U3137 (N_3137,N_2729,N_2156);
or U3138 (N_3138,N_2979,N_2720);
nor U3139 (N_3139,N_2762,N_2396);
or U3140 (N_3140,N_2097,N_2500);
nor U3141 (N_3141,N_2787,N_2191);
nand U3142 (N_3142,N_2670,N_2167);
xnor U3143 (N_3143,N_2448,N_2388);
nor U3144 (N_3144,N_2249,N_2129);
and U3145 (N_3145,N_2080,N_2830);
and U3146 (N_3146,N_2569,N_2318);
nand U3147 (N_3147,N_2173,N_2502);
nor U3148 (N_3148,N_2446,N_2919);
xnor U3149 (N_3149,N_2503,N_2828);
nor U3150 (N_3150,N_2684,N_2853);
nand U3151 (N_3151,N_2686,N_2558);
xnor U3152 (N_3152,N_2411,N_2082);
nor U3153 (N_3153,N_2216,N_2410);
and U3154 (N_3154,N_2840,N_2444);
nand U3155 (N_3155,N_2085,N_2303);
xnor U3156 (N_3156,N_2709,N_2329);
and U3157 (N_3157,N_2378,N_2582);
nand U3158 (N_3158,N_2461,N_2362);
nand U3159 (N_3159,N_2793,N_2296);
xor U3160 (N_3160,N_2909,N_2813);
nand U3161 (N_3161,N_2635,N_2024);
or U3162 (N_3162,N_2238,N_2482);
nor U3163 (N_3163,N_2590,N_2712);
nand U3164 (N_3164,N_2036,N_2019);
nor U3165 (N_3165,N_2863,N_2948);
or U3166 (N_3166,N_2320,N_2030);
or U3167 (N_3167,N_2987,N_2594);
or U3168 (N_3168,N_2018,N_2895);
or U3169 (N_3169,N_2123,N_2774);
xor U3170 (N_3170,N_2996,N_2956);
and U3171 (N_3171,N_2944,N_2012);
nor U3172 (N_3172,N_2628,N_2521);
and U3173 (N_3173,N_2834,N_2622);
or U3174 (N_3174,N_2481,N_2074);
nand U3175 (N_3175,N_2798,N_2797);
or U3176 (N_3176,N_2509,N_2079);
nor U3177 (N_3177,N_2861,N_2804);
nor U3178 (N_3178,N_2356,N_2102);
xor U3179 (N_3179,N_2537,N_2308);
xnor U3180 (N_3180,N_2599,N_2051);
or U3181 (N_3181,N_2000,N_2788);
or U3182 (N_3182,N_2515,N_2235);
xor U3183 (N_3183,N_2040,N_2928);
nor U3184 (N_3184,N_2520,N_2885);
and U3185 (N_3185,N_2187,N_2213);
or U3186 (N_3186,N_2796,N_2507);
xor U3187 (N_3187,N_2910,N_2326);
or U3188 (N_3188,N_2443,N_2682);
and U3189 (N_3189,N_2120,N_2269);
xnor U3190 (N_3190,N_2781,N_2758);
nor U3191 (N_3191,N_2829,N_2161);
xnor U3192 (N_3192,N_2631,N_2332);
xor U3193 (N_3193,N_2747,N_2066);
nand U3194 (N_3194,N_2208,N_2210);
and U3195 (N_3195,N_2155,N_2468);
nor U3196 (N_3196,N_2963,N_2746);
and U3197 (N_3197,N_2931,N_2822);
or U3198 (N_3198,N_2973,N_2001);
nor U3199 (N_3199,N_2491,N_2312);
or U3200 (N_3200,N_2214,N_2418);
nand U3201 (N_3201,N_2010,N_2391);
and U3202 (N_3202,N_2131,N_2886);
and U3203 (N_3203,N_2552,N_2904);
and U3204 (N_3204,N_2775,N_2990);
nand U3205 (N_3205,N_2737,N_2165);
or U3206 (N_3206,N_2896,N_2970);
nand U3207 (N_3207,N_2267,N_2251);
xnor U3208 (N_3208,N_2319,N_2517);
xor U3209 (N_3209,N_2412,N_2933);
xor U3210 (N_3210,N_2755,N_2450);
or U3211 (N_3211,N_2935,N_2004);
and U3212 (N_3212,N_2555,N_2233);
nor U3213 (N_3213,N_2525,N_2044);
and U3214 (N_3214,N_2276,N_2812);
nor U3215 (N_3215,N_2974,N_2392);
nor U3216 (N_3216,N_2567,N_2826);
nand U3217 (N_3217,N_2988,N_2679);
and U3218 (N_3218,N_2801,N_2314);
xor U3219 (N_3219,N_2802,N_2135);
xor U3220 (N_3220,N_2950,N_2501);
nor U3221 (N_3221,N_2553,N_2736);
or U3222 (N_3222,N_2576,N_2649);
and U3223 (N_3223,N_2917,N_2070);
nand U3224 (N_3224,N_2560,N_2295);
or U3225 (N_3225,N_2032,N_2574);
xor U3226 (N_3226,N_2048,N_2595);
xor U3227 (N_3227,N_2777,N_2049);
or U3228 (N_3228,N_2441,N_2381);
nand U3229 (N_3229,N_2960,N_2277);
nand U3230 (N_3230,N_2072,N_2865);
xor U3231 (N_3231,N_2902,N_2268);
xor U3232 (N_3232,N_2250,N_2062);
or U3233 (N_3233,N_2202,N_2678);
xnor U3234 (N_3234,N_2089,N_2528);
and U3235 (N_3235,N_2805,N_2060);
nor U3236 (N_3236,N_2160,N_2285);
and U3237 (N_3237,N_2084,N_2924);
or U3238 (N_3238,N_2473,N_2897);
nor U3239 (N_3239,N_2516,N_2513);
nor U3240 (N_3240,N_2369,N_2116);
nand U3241 (N_3241,N_2126,N_2442);
nand U3242 (N_3242,N_2573,N_2204);
or U3243 (N_3243,N_2773,N_2301);
and U3244 (N_3244,N_2417,N_2333);
and U3245 (N_3245,N_2273,N_2692);
or U3246 (N_3246,N_2374,N_2965);
and U3247 (N_3247,N_2006,N_2986);
or U3248 (N_3248,N_2976,N_2077);
and U3249 (N_3249,N_2721,N_2300);
xor U3250 (N_3250,N_2549,N_2874);
or U3251 (N_3251,N_2447,N_2244);
or U3252 (N_3252,N_2168,N_2224);
nand U3253 (N_3253,N_2547,N_2816);
or U3254 (N_3254,N_2419,N_2132);
xnor U3255 (N_3255,N_2708,N_2824);
nor U3256 (N_3256,N_2873,N_2536);
xnor U3257 (N_3257,N_2499,N_2256);
or U3258 (N_3258,N_2305,N_2859);
and U3259 (N_3259,N_2677,N_2942);
or U3260 (N_3260,N_2150,N_2280);
nor U3261 (N_3261,N_2075,N_2338);
and U3262 (N_3262,N_2860,N_2236);
nor U3263 (N_3263,N_2511,N_2810);
or U3264 (N_3264,N_2367,N_2178);
or U3265 (N_3265,N_2733,N_2207);
and U3266 (N_3266,N_2761,N_2130);
or U3267 (N_3267,N_2121,N_2601);
nand U3268 (N_3268,N_2270,N_2671);
nand U3269 (N_3269,N_2645,N_2467);
nand U3270 (N_3270,N_2630,N_2581);
xor U3271 (N_3271,N_2633,N_2105);
nor U3272 (N_3272,N_2743,N_2637);
nor U3273 (N_3273,N_2838,N_2222);
nand U3274 (N_3274,N_2206,N_2699);
nand U3275 (N_3275,N_2890,N_2980);
or U3276 (N_3276,N_2609,N_2903);
and U3277 (N_3277,N_2415,N_2545);
nor U3278 (N_3278,N_2566,N_2915);
or U3279 (N_3279,N_2694,N_2212);
nand U3280 (N_3280,N_2526,N_2346);
nor U3281 (N_3281,N_2837,N_2676);
xor U3282 (N_3282,N_2453,N_2390);
or U3283 (N_3283,N_2939,N_2197);
nand U3284 (N_3284,N_2128,N_2659);
nand U3285 (N_3285,N_2991,N_2753);
xor U3286 (N_3286,N_2688,N_2137);
nor U3287 (N_3287,N_2055,N_2142);
nand U3288 (N_3288,N_2241,N_2518);
or U3289 (N_3289,N_2634,N_2008);
xor U3290 (N_3290,N_2345,N_2067);
xor U3291 (N_3291,N_2416,N_2669);
xnor U3292 (N_3292,N_2522,N_2475);
nand U3293 (N_3293,N_2022,N_2349);
nand U3294 (N_3294,N_2561,N_2855);
nand U3295 (N_3295,N_2717,N_2757);
and U3296 (N_3296,N_2259,N_2385);
xnor U3297 (N_3297,N_2177,N_2947);
xor U3298 (N_3298,N_2770,N_2376);
and U3299 (N_3299,N_2867,N_2593);
or U3300 (N_3300,N_2257,N_2405);
nor U3301 (N_3301,N_2282,N_2190);
xnor U3302 (N_3302,N_2498,N_2785);
nand U3303 (N_3303,N_2589,N_2099);
nand U3304 (N_3304,N_2745,N_2457);
and U3305 (N_3305,N_2146,N_2543);
nor U3306 (N_3306,N_2174,N_2975);
xnor U3307 (N_3307,N_2994,N_2719);
or U3308 (N_3308,N_2618,N_2815);
nor U3309 (N_3309,N_2898,N_2493);
or U3310 (N_3310,N_2343,N_2811);
or U3311 (N_3311,N_2687,N_2716);
nor U3312 (N_3312,N_2047,N_2680);
nand U3313 (N_3313,N_2586,N_2045);
xor U3314 (N_3314,N_2771,N_2772);
or U3315 (N_3315,N_2401,N_2791);
and U3316 (N_3316,N_2766,N_2432);
nand U3317 (N_3317,N_2359,N_2026);
nand U3318 (N_3318,N_2164,N_2985);
or U3319 (N_3319,N_2138,N_2742);
and U3320 (N_3320,N_2624,N_2689);
xor U3321 (N_3321,N_2530,N_2866);
xor U3322 (N_3322,N_2763,N_2400);
nand U3323 (N_3323,N_2377,N_2397);
xor U3324 (N_3324,N_2472,N_2551);
xnor U3325 (N_3325,N_2426,N_2809);
and U3326 (N_3326,N_2907,N_2660);
or U3327 (N_3327,N_2615,N_2760);
nand U3328 (N_3328,N_2953,N_2219);
xnor U3329 (N_3329,N_2078,N_2713);
or U3330 (N_3330,N_2559,N_2313);
nor U3331 (N_3331,N_2248,N_2307);
nor U3332 (N_3332,N_2291,N_2456);
nor U3333 (N_3333,N_2756,N_2459);
nor U3334 (N_3334,N_2252,N_2949);
nand U3335 (N_3335,N_2398,N_2532);
nand U3336 (N_3336,N_2932,N_2920);
nand U3337 (N_3337,N_2572,N_2856);
and U3338 (N_3338,N_2220,N_2583);
nor U3339 (N_3339,N_2423,N_2347);
and U3340 (N_3340,N_2487,N_2148);
and U3341 (N_3341,N_2341,N_2535);
nor U3342 (N_3342,N_2221,N_2225);
nand U3343 (N_3343,N_2715,N_2186);
and U3344 (N_3344,N_2043,N_2476);
nand U3345 (N_3345,N_2188,N_2596);
nand U3346 (N_3346,N_2614,N_2310);
xor U3347 (N_3347,N_2880,N_2827);
nor U3348 (N_3348,N_2112,N_2557);
nor U3349 (N_3349,N_2228,N_2611);
nand U3350 (N_3350,N_2240,N_2730);
nor U3351 (N_3351,N_2407,N_2529);
and U3352 (N_3352,N_2666,N_2769);
nor U3353 (N_3353,N_2750,N_2675);
or U3354 (N_3354,N_2209,N_2153);
or U3355 (N_3355,N_2258,N_2854);
nand U3356 (N_3356,N_2612,N_2833);
nand U3357 (N_3357,N_2104,N_2564);
nor U3358 (N_3358,N_2835,N_2922);
xor U3359 (N_3359,N_2652,N_2591);
nor U3360 (N_3360,N_2548,N_2823);
nand U3361 (N_3361,N_2223,N_2355);
and U3362 (N_3362,N_2430,N_2452);
nand U3363 (N_3363,N_2971,N_2851);
or U3364 (N_3364,N_2648,N_2264);
nor U3365 (N_3365,N_2512,N_2489);
and U3366 (N_3366,N_2455,N_2778);
or U3367 (N_3367,N_2941,N_2883);
nor U3368 (N_3368,N_2619,N_2293);
and U3369 (N_3369,N_2705,N_2668);
nand U3370 (N_3370,N_2348,N_2665);
or U3371 (N_3371,N_2464,N_2767);
xnor U3372 (N_3372,N_2086,N_2765);
or U3373 (N_3373,N_2913,N_2918);
xnor U3374 (N_3374,N_2923,N_2556);
nor U3375 (N_3375,N_2519,N_2124);
nand U3376 (N_3376,N_2253,N_2114);
xnor U3377 (N_3377,N_2226,N_2231);
nor U3378 (N_3378,N_2171,N_2752);
nand U3379 (N_3379,N_2095,N_2843);
and U3380 (N_3380,N_2340,N_2185);
nand U3381 (N_3381,N_2064,N_2899);
and U3382 (N_3382,N_2982,N_2966);
nand U3383 (N_3383,N_2808,N_2691);
nand U3384 (N_3384,N_2806,N_2406);
nand U3385 (N_3385,N_2842,N_2109);
and U3386 (N_3386,N_2790,N_2125);
and U3387 (N_3387,N_2445,N_2373);
nand U3388 (N_3388,N_2995,N_2930);
nor U3389 (N_3389,N_2580,N_2707);
nor U3390 (N_3390,N_2998,N_2554);
xnor U3391 (N_3391,N_2984,N_2868);
and U3392 (N_3392,N_2646,N_2604);
and U3393 (N_3393,N_2725,N_2141);
and U3394 (N_3394,N_2050,N_2731);
xor U3395 (N_3395,N_2046,N_2799);
nand U3396 (N_3396,N_2337,N_2568);
nand U3397 (N_3397,N_2847,N_2471);
nor U3398 (N_3398,N_2658,N_2339);
and U3399 (N_3399,N_2632,N_2570);
nor U3400 (N_3400,N_2413,N_2409);
xnor U3401 (N_3401,N_2764,N_2038);
nor U3402 (N_3402,N_2700,N_2420);
nor U3403 (N_3403,N_2740,N_2096);
and U3404 (N_3404,N_2531,N_2784);
nor U3405 (N_3405,N_2366,N_2071);
and U3406 (N_3406,N_2977,N_2372);
and U3407 (N_3407,N_2541,N_2584);
xor U3408 (N_3408,N_2260,N_2571);
nor U3409 (N_3409,N_2964,N_2914);
xor U3410 (N_3410,N_2857,N_2674);
nand U3411 (N_3411,N_2514,N_2232);
and U3412 (N_3412,N_2107,N_2434);
and U3413 (N_3413,N_2724,N_2162);
and U3414 (N_3414,N_2063,N_2184);
nor U3415 (N_3415,N_2727,N_2474);
and U3416 (N_3416,N_2925,N_2641);
nand U3417 (N_3417,N_2732,N_2954);
or U3418 (N_3418,N_2685,N_2894);
and U3419 (N_3419,N_2483,N_2091);
and U3420 (N_3420,N_2879,N_2538);
xnor U3421 (N_3421,N_2542,N_2978);
nand U3422 (N_3422,N_2937,N_2608);
or U3423 (N_3423,N_2588,N_2993);
and U3424 (N_3424,N_2387,N_2353);
xor U3425 (N_3425,N_2906,N_2938);
and U3426 (N_3426,N_2357,N_2056);
and U3427 (N_3427,N_2620,N_2052);
and U3428 (N_3428,N_2317,N_2997);
xnor U3429 (N_3429,N_2850,N_2484);
or U3430 (N_3430,N_2272,N_2389);
nor U3431 (N_3431,N_2734,N_2878);
xnor U3432 (N_3432,N_2524,N_2100);
nand U3433 (N_3433,N_2754,N_2304);
or U3434 (N_3434,N_2243,N_2718);
xor U3435 (N_3435,N_2921,N_2946);
and U3436 (N_3436,N_2429,N_2076);
or U3437 (N_3437,N_2544,N_2846);
nand U3438 (N_3438,N_2375,N_2463);
and U3439 (N_3439,N_2782,N_2603);
xor U3440 (N_3440,N_2013,N_2972);
nor U3441 (N_3441,N_2042,N_2431);
and U3442 (N_3442,N_2211,N_2113);
or U3443 (N_3443,N_2726,N_2433);
nor U3444 (N_3444,N_2644,N_2363);
xnor U3445 (N_3445,N_2887,N_2882);
and U3446 (N_3446,N_2427,N_2028);
nor U3447 (N_3447,N_2017,N_2952);
or U3448 (N_3448,N_2610,N_2800);
and U3449 (N_3449,N_2239,N_2695);
xnor U3450 (N_3450,N_2492,N_2315);
nand U3451 (N_3451,N_2414,N_2470);
nor U3452 (N_3452,N_2181,N_2831);
or U3453 (N_3453,N_2035,N_2194);
or U3454 (N_3454,N_2710,N_2527);
xor U3455 (N_3455,N_2654,N_2183);
nor U3456 (N_3456,N_2101,N_2425);
or U3457 (N_3457,N_2999,N_2154);
nor U3458 (N_3458,N_2577,N_2011);
or U3459 (N_3459,N_2016,N_2497);
and U3460 (N_3460,N_2723,N_2289);
or U3461 (N_3461,N_2294,N_2449);
or U3462 (N_3462,N_2041,N_2127);
nand U3463 (N_3463,N_2701,N_2693);
nand U3464 (N_3464,N_2424,N_2182);
xnor U3465 (N_3465,N_2480,N_2803);
xor U3466 (N_3466,N_2234,N_2278);
xor U3467 (N_3467,N_2176,N_2962);
nand U3468 (N_3468,N_2626,N_2714);
nor U3469 (N_3469,N_2864,N_2667);
and U3470 (N_3470,N_2697,N_2629);
nor U3471 (N_3471,N_2143,N_2139);
nand U3472 (N_3472,N_2916,N_2103);
or U3473 (N_3473,N_2877,N_2158);
nor U3474 (N_3474,N_2477,N_2698);
xnor U3475 (N_3475,N_2065,N_2983);
xnor U3476 (N_3476,N_2379,N_2306);
xor U3477 (N_3477,N_2057,N_2722);
xor U3478 (N_3478,N_2870,N_2627);
xnor U3479 (N_3479,N_2912,N_2193);
nor U3480 (N_3480,N_2382,N_2789);
nor U3481 (N_3481,N_2283,N_2327);
or U3482 (N_3482,N_2230,N_2119);
xnor U3483 (N_3483,N_2321,N_2265);
or U3484 (N_3484,N_2466,N_2653);
nor U3485 (N_3485,N_2506,N_2380);
or U3486 (N_3486,N_2981,N_2196);
and U3487 (N_3487,N_2587,N_2735);
nand U3488 (N_3488,N_2636,N_2151);
nor U3489 (N_3489,N_2881,N_2365);
and U3490 (N_3490,N_2460,N_2901);
and U3491 (N_3491,N_2934,N_2364);
xor U3492 (N_3492,N_2245,N_2465);
nand U3493 (N_3493,N_2059,N_2795);
nand U3494 (N_3494,N_2384,N_2738);
nand U3495 (N_3495,N_2322,N_2792);
nor U3496 (N_3496,N_2316,N_2776);
nor U3497 (N_3497,N_2217,N_2255);
nand U3498 (N_3498,N_2111,N_2768);
or U3499 (N_3499,N_2562,N_2605);
or U3500 (N_3500,N_2012,N_2428);
nand U3501 (N_3501,N_2108,N_2058);
and U3502 (N_3502,N_2466,N_2555);
nand U3503 (N_3503,N_2079,N_2959);
and U3504 (N_3504,N_2614,N_2354);
and U3505 (N_3505,N_2019,N_2677);
or U3506 (N_3506,N_2023,N_2172);
nor U3507 (N_3507,N_2749,N_2697);
or U3508 (N_3508,N_2015,N_2691);
nor U3509 (N_3509,N_2899,N_2276);
and U3510 (N_3510,N_2466,N_2030);
nor U3511 (N_3511,N_2595,N_2059);
xnor U3512 (N_3512,N_2386,N_2085);
and U3513 (N_3513,N_2981,N_2356);
nand U3514 (N_3514,N_2783,N_2149);
or U3515 (N_3515,N_2780,N_2978);
and U3516 (N_3516,N_2332,N_2472);
or U3517 (N_3517,N_2558,N_2680);
xor U3518 (N_3518,N_2470,N_2797);
nor U3519 (N_3519,N_2928,N_2310);
xnor U3520 (N_3520,N_2257,N_2999);
xor U3521 (N_3521,N_2832,N_2081);
and U3522 (N_3522,N_2525,N_2289);
or U3523 (N_3523,N_2807,N_2355);
nor U3524 (N_3524,N_2427,N_2722);
and U3525 (N_3525,N_2779,N_2338);
xor U3526 (N_3526,N_2657,N_2228);
nand U3527 (N_3527,N_2797,N_2564);
xor U3528 (N_3528,N_2442,N_2570);
and U3529 (N_3529,N_2956,N_2216);
or U3530 (N_3530,N_2515,N_2069);
nand U3531 (N_3531,N_2023,N_2272);
or U3532 (N_3532,N_2402,N_2368);
xnor U3533 (N_3533,N_2168,N_2170);
nor U3534 (N_3534,N_2560,N_2440);
xor U3535 (N_3535,N_2121,N_2974);
nor U3536 (N_3536,N_2916,N_2527);
nand U3537 (N_3537,N_2042,N_2732);
xnor U3538 (N_3538,N_2849,N_2229);
or U3539 (N_3539,N_2643,N_2334);
nand U3540 (N_3540,N_2976,N_2186);
nand U3541 (N_3541,N_2202,N_2368);
nor U3542 (N_3542,N_2281,N_2066);
nand U3543 (N_3543,N_2004,N_2052);
and U3544 (N_3544,N_2822,N_2311);
and U3545 (N_3545,N_2333,N_2811);
nor U3546 (N_3546,N_2304,N_2641);
nand U3547 (N_3547,N_2210,N_2979);
nor U3548 (N_3548,N_2387,N_2059);
nand U3549 (N_3549,N_2508,N_2429);
or U3550 (N_3550,N_2169,N_2314);
or U3551 (N_3551,N_2711,N_2697);
xor U3552 (N_3552,N_2185,N_2167);
and U3553 (N_3553,N_2632,N_2635);
nor U3554 (N_3554,N_2025,N_2805);
and U3555 (N_3555,N_2438,N_2220);
and U3556 (N_3556,N_2227,N_2426);
or U3557 (N_3557,N_2513,N_2751);
nor U3558 (N_3558,N_2994,N_2378);
nor U3559 (N_3559,N_2886,N_2779);
nor U3560 (N_3560,N_2614,N_2181);
nor U3561 (N_3561,N_2534,N_2283);
nand U3562 (N_3562,N_2499,N_2987);
nand U3563 (N_3563,N_2445,N_2196);
nor U3564 (N_3564,N_2384,N_2306);
nand U3565 (N_3565,N_2574,N_2916);
nand U3566 (N_3566,N_2131,N_2208);
xnor U3567 (N_3567,N_2356,N_2213);
or U3568 (N_3568,N_2857,N_2921);
nor U3569 (N_3569,N_2901,N_2547);
or U3570 (N_3570,N_2443,N_2064);
nor U3571 (N_3571,N_2876,N_2858);
xnor U3572 (N_3572,N_2444,N_2019);
and U3573 (N_3573,N_2632,N_2380);
and U3574 (N_3574,N_2032,N_2628);
or U3575 (N_3575,N_2817,N_2289);
xor U3576 (N_3576,N_2203,N_2163);
or U3577 (N_3577,N_2248,N_2110);
or U3578 (N_3578,N_2225,N_2927);
or U3579 (N_3579,N_2617,N_2503);
nand U3580 (N_3580,N_2784,N_2931);
xnor U3581 (N_3581,N_2284,N_2601);
xor U3582 (N_3582,N_2222,N_2680);
xor U3583 (N_3583,N_2621,N_2781);
nor U3584 (N_3584,N_2627,N_2291);
nor U3585 (N_3585,N_2383,N_2692);
and U3586 (N_3586,N_2347,N_2861);
and U3587 (N_3587,N_2808,N_2029);
and U3588 (N_3588,N_2816,N_2857);
nand U3589 (N_3589,N_2085,N_2543);
and U3590 (N_3590,N_2369,N_2589);
and U3591 (N_3591,N_2029,N_2374);
nand U3592 (N_3592,N_2729,N_2868);
nand U3593 (N_3593,N_2412,N_2195);
xnor U3594 (N_3594,N_2646,N_2841);
and U3595 (N_3595,N_2869,N_2429);
and U3596 (N_3596,N_2533,N_2024);
or U3597 (N_3597,N_2230,N_2953);
and U3598 (N_3598,N_2160,N_2219);
nand U3599 (N_3599,N_2716,N_2604);
and U3600 (N_3600,N_2432,N_2618);
nor U3601 (N_3601,N_2148,N_2047);
xnor U3602 (N_3602,N_2005,N_2685);
or U3603 (N_3603,N_2758,N_2691);
xnor U3604 (N_3604,N_2480,N_2455);
or U3605 (N_3605,N_2747,N_2608);
or U3606 (N_3606,N_2515,N_2281);
nor U3607 (N_3607,N_2264,N_2409);
xor U3608 (N_3608,N_2730,N_2188);
nand U3609 (N_3609,N_2893,N_2191);
and U3610 (N_3610,N_2726,N_2454);
nor U3611 (N_3611,N_2660,N_2062);
or U3612 (N_3612,N_2679,N_2387);
nand U3613 (N_3613,N_2576,N_2316);
nand U3614 (N_3614,N_2984,N_2325);
and U3615 (N_3615,N_2849,N_2111);
or U3616 (N_3616,N_2313,N_2340);
nor U3617 (N_3617,N_2397,N_2731);
and U3618 (N_3618,N_2941,N_2256);
nand U3619 (N_3619,N_2817,N_2241);
nor U3620 (N_3620,N_2387,N_2899);
and U3621 (N_3621,N_2882,N_2916);
nand U3622 (N_3622,N_2619,N_2383);
xnor U3623 (N_3623,N_2551,N_2124);
nor U3624 (N_3624,N_2792,N_2299);
or U3625 (N_3625,N_2314,N_2981);
xor U3626 (N_3626,N_2384,N_2431);
nor U3627 (N_3627,N_2813,N_2699);
and U3628 (N_3628,N_2345,N_2037);
and U3629 (N_3629,N_2039,N_2196);
nand U3630 (N_3630,N_2096,N_2365);
nand U3631 (N_3631,N_2147,N_2574);
nand U3632 (N_3632,N_2820,N_2795);
or U3633 (N_3633,N_2138,N_2372);
or U3634 (N_3634,N_2998,N_2182);
xnor U3635 (N_3635,N_2558,N_2400);
xor U3636 (N_3636,N_2523,N_2682);
or U3637 (N_3637,N_2602,N_2767);
and U3638 (N_3638,N_2142,N_2920);
and U3639 (N_3639,N_2558,N_2084);
and U3640 (N_3640,N_2238,N_2940);
xor U3641 (N_3641,N_2425,N_2085);
nor U3642 (N_3642,N_2834,N_2933);
nor U3643 (N_3643,N_2320,N_2701);
xnor U3644 (N_3644,N_2191,N_2550);
nand U3645 (N_3645,N_2450,N_2018);
xor U3646 (N_3646,N_2360,N_2118);
nand U3647 (N_3647,N_2112,N_2715);
nor U3648 (N_3648,N_2590,N_2747);
nor U3649 (N_3649,N_2136,N_2909);
nor U3650 (N_3650,N_2869,N_2039);
or U3651 (N_3651,N_2751,N_2156);
xor U3652 (N_3652,N_2339,N_2200);
nand U3653 (N_3653,N_2928,N_2879);
or U3654 (N_3654,N_2302,N_2529);
xnor U3655 (N_3655,N_2435,N_2624);
or U3656 (N_3656,N_2792,N_2722);
and U3657 (N_3657,N_2630,N_2652);
nor U3658 (N_3658,N_2481,N_2759);
nand U3659 (N_3659,N_2915,N_2982);
or U3660 (N_3660,N_2388,N_2488);
nor U3661 (N_3661,N_2700,N_2843);
nor U3662 (N_3662,N_2330,N_2700);
nand U3663 (N_3663,N_2428,N_2571);
xor U3664 (N_3664,N_2193,N_2270);
or U3665 (N_3665,N_2447,N_2552);
nand U3666 (N_3666,N_2747,N_2973);
and U3667 (N_3667,N_2444,N_2746);
nand U3668 (N_3668,N_2390,N_2789);
xnor U3669 (N_3669,N_2766,N_2721);
or U3670 (N_3670,N_2231,N_2450);
xor U3671 (N_3671,N_2258,N_2248);
or U3672 (N_3672,N_2673,N_2357);
and U3673 (N_3673,N_2015,N_2270);
or U3674 (N_3674,N_2555,N_2526);
xor U3675 (N_3675,N_2062,N_2421);
and U3676 (N_3676,N_2653,N_2674);
nor U3677 (N_3677,N_2160,N_2794);
nand U3678 (N_3678,N_2074,N_2106);
nand U3679 (N_3679,N_2257,N_2080);
or U3680 (N_3680,N_2422,N_2622);
nor U3681 (N_3681,N_2773,N_2536);
nand U3682 (N_3682,N_2922,N_2865);
nand U3683 (N_3683,N_2284,N_2065);
xor U3684 (N_3684,N_2945,N_2147);
nor U3685 (N_3685,N_2464,N_2191);
or U3686 (N_3686,N_2433,N_2815);
nor U3687 (N_3687,N_2596,N_2762);
and U3688 (N_3688,N_2492,N_2924);
and U3689 (N_3689,N_2348,N_2352);
nor U3690 (N_3690,N_2849,N_2616);
and U3691 (N_3691,N_2027,N_2505);
nand U3692 (N_3692,N_2305,N_2944);
nand U3693 (N_3693,N_2135,N_2475);
xnor U3694 (N_3694,N_2041,N_2510);
nand U3695 (N_3695,N_2216,N_2883);
nand U3696 (N_3696,N_2283,N_2261);
or U3697 (N_3697,N_2573,N_2610);
and U3698 (N_3698,N_2948,N_2169);
and U3699 (N_3699,N_2661,N_2739);
nor U3700 (N_3700,N_2329,N_2916);
xor U3701 (N_3701,N_2326,N_2597);
and U3702 (N_3702,N_2844,N_2441);
or U3703 (N_3703,N_2409,N_2992);
or U3704 (N_3704,N_2339,N_2348);
xor U3705 (N_3705,N_2962,N_2761);
nand U3706 (N_3706,N_2972,N_2186);
or U3707 (N_3707,N_2905,N_2663);
xnor U3708 (N_3708,N_2800,N_2355);
and U3709 (N_3709,N_2202,N_2126);
nand U3710 (N_3710,N_2278,N_2366);
and U3711 (N_3711,N_2817,N_2757);
xor U3712 (N_3712,N_2210,N_2768);
or U3713 (N_3713,N_2750,N_2865);
and U3714 (N_3714,N_2124,N_2186);
nand U3715 (N_3715,N_2594,N_2224);
xor U3716 (N_3716,N_2777,N_2435);
or U3717 (N_3717,N_2501,N_2537);
nor U3718 (N_3718,N_2139,N_2897);
xnor U3719 (N_3719,N_2777,N_2788);
nand U3720 (N_3720,N_2559,N_2632);
or U3721 (N_3721,N_2039,N_2978);
and U3722 (N_3722,N_2306,N_2654);
xor U3723 (N_3723,N_2397,N_2141);
nor U3724 (N_3724,N_2166,N_2012);
xor U3725 (N_3725,N_2275,N_2014);
or U3726 (N_3726,N_2729,N_2329);
or U3727 (N_3727,N_2163,N_2513);
xnor U3728 (N_3728,N_2833,N_2062);
nand U3729 (N_3729,N_2436,N_2902);
xnor U3730 (N_3730,N_2001,N_2046);
nor U3731 (N_3731,N_2547,N_2866);
nand U3732 (N_3732,N_2446,N_2623);
nor U3733 (N_3733,N_2433,N_2841);
or U3734 (N_3734,N_2801,N_2842);
nand U3735 (N_3735,N_2295,N_2038);
xor U3736 (N_3736,N_2384,N_2138);
nor U3737 (N_3737,N_2091,N_2439);
xnor U3738 (N_3738,N_2944,N_2702);
nand U3739 (N_3739,N_2083,N_2486);
nor U3740 (N_3740,N_2945,N_2672);
and U3741 (N_3741,N_2690,N_2851);
and U3742 (N_3742,N_2399,N_2648);
xor U3743 (N_3743,N_2251,N_2040);
or U3744 (N_3744,N_2992,N_2593);
nand U3745 (N_3745,N_2672,N_2572);
nor U3746 (N_3746,N_2994,N_2221);
nand U3747 (N_3747,N_2099,N_2281);
nand U3748 (N_3748,N_2316,N_2812);
xnor U3749 (N_3749,N_2773,N_2154);
and U3750 (N_3750,N_2831,N_2808);
nor U3751 (N_3751,N_2280,N_2679);
and U3752 (N_3752,N_2794,N_2000);
nand U3753 (N_3753,N_2478,N_2793);
nand U3754 (N_3754,N_2247,N_2487);
nand U3755 (N_3755,N_2154,N_2004);
nand U3756 (N_3756,N_2013,N_2637);
xor U3757 (N_3757,N_2142,N_2563);
or U3758 (N_3758,N_2031,N_2425);
xor U3759 (N_3759,N_2527,N_2226);
nand U3760 (N_3760,N_2956,N_2997);
or U3761 (N_3761,N_2013,N_2608);
and U3762 (N_3762,N_2114,N_2652);
xnor U3763 (N_3763,N_2411,N_2620);
xnor U3764 (N_3764,N_2828,N_2002);
nor U3765 (N_3765,N_2925,N_2837);
or U3766 (N_3766,N_2903,N_2496);
and U3767 (N_3767,N_2921,N_2557);
xor U3768 (N_3768,N_2658,N_2347);
nand U3769 (N_3769,N_2921,N_2229);
or U3770 (N_3770,N_2735,N_2898);
nand U3771 (N_3771,N_2719,N_2027);
and U3772 (N_3772,N_2534,N_2795);
xnor U3773 (N_3773,N_2866,N_2809);
xor U3774 (N_3774,N_2921,N_2479);
nor U3775 (N_3775,N_2687,N_2001);
nand U3776 (N_3776,N_2953,N_2373);
or U3777 (N_3777,N_2365,N_2291);
xor U3778 (N_3778,N_2847,N_2698);
nor U3779 (N_3779,N_2689,N_2920);
nand U3780 (N_3780,N_2199,N_2716);
nand U3781 (N_3781,N_2919,N_2662);
and U3782 (N_3782,N_2391,N_2511);
and U3783 (N_3783,N_2427,N_2656);
nand U3784 (N_3784,N_2157,N_2669);
or U3785 (N_3785,N_2567,N_2726);
and U3786 (N_3786,N_2940,N_2929);
xor U3787 (N_3787,N_2995,N_2256);
nor U3788 (N_3788,N_2398,N_2448);
nand U3789 (N_3789,N_2895,N_2541);
or U3790 (N_3790,N_2774,N_2932);
nand U3791 (N_3791,N_2168,N_2744);
or U3792 (N_3792,N_2480,N_2412);
nand U3793 (N_3793,N_2750,N_2699);
nor U3794 (N_3794,N_2237,N_2153);
and U3795 (N_3795,N_2626,N_2338);
nand U3796 (N_3796,N_2707,N_2885);
and U3797 (N_3797,N_2488,N_2457);
xor U3798 (N_3798,N_2735,N_2450);
or U3799 (N_3799,N_2107,N_2536);
or U3800 (N_3800,N_2593,N_2667);
or U3801 (N_3801,N_2516,N_2759);
or U3802 (N_3802,N_2434,N_2168);
and U3803 (N_3803,N_2653,N_2597);
nand U3804 (N_3804,N_2895,N_2132);
nor U3805 (N_3805,N_2819,N_2309);
or U3806 (N_3806,N_2938,N_2781);
nand U3807 (N_3807,N_2988,N_2655);
nand U3808 (N_3808,N_2464,N_2612);
or U3809 (N_3809,N_2839,N_2020);
xor U3810 (N_3810,N_2556,N_2273);
and U3811 (N_3811,N_2931,N_2794);
nor U3812 (N_3812,N_2321,N_2437);
and U3813 (N_3813,N_2818,N_2534);
xor U3814 (N_3814,N_2276,N_2931);
or U3815 (N_3815,N_2611,N_2562);
or U3816 (N_3816,N_2730,N_2513);
and U3817 (N_3817,N_2563,N_2938);
xor U3818 (N_3818,N_2425,N_2537);
nand U3819 (N_3819,N_2947,N_2493);
xor U3820 (N_3820,N_2117,N_2670);
or U3821 (N_3821,N_2902,N_2962);
nor U3822 (N_3822,N_2142,N_2829);
and U3823 (N_3823,N_2054,N_2193);
and U3824 (N_3824,N_2805,N_2114);
or U3825 (N_3825,N_2479,N_2927);
or U3826 (N_3826,N_2285,N_2447);
and U3827 (N_3827,N_2380,N_2820);
nand U3828 (N_3828,N_2542,N_2583);
nand U3829 (N_3829,N_2931,N_2271);
and U3830 (N_3830,N_2806,N_2205);
and U3831 (N_3831,N_2428,N_2489);
nor U3832 (N_3832,N_2521,N_2382);
nor U3833 (N_3833,N_2696,N_2635);
nand U3834 (N_3834,N_2513,N_2615);
or U3835 (N_3835,N_2554,N_2114);
or U3836 (N_3836,N_2690,N_2914);
xor U3837 (N_3837,N_2684,N_2632);
nor U3838 (N_3838,N_2315,N_2569);
and U3839 (N_3839,N_2727,N_2940);
and U3840 (N_3840,N_2028,N_2685);
nand U3841 (N_3841,N_2453,N_2054);
and U3842 (N_3842,N_2980,N_2808);
nor U3843 (N_3843,N_2256,N_2998);
nor U3844 (N_3844,N_2014,N_2731);
xor U3845 (N_3845,N_2501,N_2068);
nand U3846 (N_3846,N_2317,N_2657);
nand U3847 (N_3847,N_2123,N_2984);
nor U3848 (N_3848,N_2439,N_2765);
nor U3849 (N_3849,N_2565,N_2308);
or U3850 (N_3850,N_2867,N_2012);
xnor U3851 (N_3851,N_2702,N_2453);
or U3852 (N_3852,N_2295,N_2197);
nand U3853 (N_3853,N_2343,N_2883);
and U3854 (N_3854,N_2450,N_2861);
nand U3855 (N_3855,N_2151,N_2908);
and U3856 (N_3856,N_2695,N_2279);
or U3857 (N_3857,N_2425,N_2842);
xnor U3858 (N_3858,N_2535,N_2930);
xnor U3859 (N_3859,N_2883,N_2870);
nor U3860 (N_3860,N_2500,N_2609);
or U3861 (N_3861,N_2427,N_2649);
xor U3862 (N_3862,N_2043,N_2755);
xor U3863 (N_3863,N_2715,N_2573);
xnor U3864 (N_3864,N_2440,N_2783);
and U3865 (N_3865,N_2874,N_2512);
xor U3866 (N_3866,N_2085,N_2289);
nor U3867 (N_3867,N_2113,N_2311);
xnor U3868 (N_3868,N_2194,N_2447);
or U3869 (N_3869,N_2016,N_2322);
nor U3870 (N_3870,N_2992,N_2188);
nor U3871 (N_3871,N_2926,N_2119);
xnor U3872 (N_3872,N_2379,N_2202);
and U3873 (N_3873,N_2225,N_2483);
xnor U3874 (N_3874,N_2813,N_2664);
nor U3875 (N_3875,N_2494,N_2011);
or U3876 (N_3876,N_2750,N_2541);
and U3877 (N_3877,N_2535,N_2602);
nand U3878 (N_3878,N_2753,N_2648);
and U3879 (N_3879,N_2476,N_2233);
or U3880 (N_3880,N_2640,N_2964);
or U3881 (N_3881,N_2227,N_2255);
nand U3882 (N_3882,N_2263,N_2743);
and U3883 (N_3883,N_2991,N_2491);
nor U3884 (N_3884,N_2158,N_2452);
nor U3885 (N_3885,N_2587,N_2866);
nor U3886 (N_3886,N_2375,N_2322);
xor U3887 (N_3887,N_2434,N_2447);
and U3888 (N_3888,N_2810,N_2405);
nor U3889 (N_3889,N_2984,N_2268);
or U3890 (N_3890,N_2254,N_2139);
nand U3891 (N_3891,N_2171,N_2534);
xor U3892 (N_3892,N_2396,N_2560);
nand U3893 (N_3893,N_2772,N_2449);
and U3894 (N_3894,N_2137,N_2544);
xnor U3895 (N_3895,N_2842,N_2671);
nand U3896 (N_3896,N_2816,N_2092);
nand U3897 (N_3897,N_2842,N_2686);
nor U3898 (N_3898,N_2240,N_2580);
or U3899 (N_3899,N_2311,N_2933);
nand U3900 (N_3900,N_2203,N_2589);
and U3901 (N_3901,N_2481,N_2657);
or U3902 (N_3902,N_2522,N_2864);
and U3903 (N_3903,N_2392,N_2419);
or U3904 (N_3904,N_2989,N_2943);
nand U3905 (N_3905,N_2348,N_2668);
nand U3906 (N_3906,N_2504,N_2633);
or U3907 (N_3907,N_2235,N_2276);
nor U3908 (N_3908,N_2313,N_2481);
or U3909 (N_3909,N_2850,N_2240);
or U3910 (N_3910,N_2033,N_2839);
or U3911 (N_3911,N_2413,N_2048);
or U3912 (N_3912,N_2955,N_2568);
xor U3913 (N_3913,N_2778,N_2033);
nand U3914 (N_3914,N_2692,N_2670);
xnor U3915 (N_3915,N_2993,N_2973);
nand U3916 (N_3916,N_2386,N_2234);
and U3917 (N_3917,N_2084,N_2478);
nor U3918 (N_3918,N_2604,N_2011);
nand U3919 (N_3919,N_2418,N_2118);
xnor U3920 (N_3920,N_2018,N_2419);
nor U3921 (N_3921,N_2590,N_2142);
and U3922 (N_3922,N_2387,N_2811);
xnor U3923 (N_3923,N_2413,N_2622);
nor U3924 (N_3924,N_2864,N_2372);
nor U3925 (N_3925,N_2155,N_2962);
nor U3926 (N_3926,N_2611,N_2034);
nand U3927 (N_3927,N_2632,N_2547);
or U3928 (N_3928,N_2802,N_2510);
xnor U3929 (N_3929,N_2632,N_2251);
xor U3930 (N_3930,N_2157,N_2426);
nand U3931 (N_3931,N_2006,N_2240);
nand U3932 (N_3932,N_2105,N_2959);
xnor U3933 (N_3933,N_2679,N_2095);
xor U3934 (N_3934,N_2987,N_2138);
and U3935 (N_3935,N_2050,N_2084);
or U3936 (N_3936,N_2076,N_2319);
and U3937 (N_3937,N_2896,N_2254);
nand U3938 (N_3938,N_2805,N_2945);
or U3939 (N_3939,N_2741,N_2614);
or U3940 (N_3940,N_2383,N_2326);
nand U3941 (N_3941,N_2091,N_2356);
nand U3942 (N_3942,N_2093,N_2328);
nand U3943 (N_3943,N_2182,N_2633);
or U3944 (N_3944,N_2340,N_2090);
xnor U3945 (N_3945,N_2566,N_2393);
or U3946 (N_3946,N_2067,N_2408);
or U3947 (N_3947,N_2030,N_2776);
nor U3948 (N_3948,N_2309,N_2963);
xor U3949 (N_3949,N_2197,N_2058);
nand U3950 (N_3950,N_2334,N_2296);
and U3951 (N_3951,N_2172,N_2101);
or U3952 (N_3952,N_2599,N_2490);
xnor U3953 (N_3953,N_2747,N_2922);
nand U3954 (N_3954,N_2276,N_2525);
and U3955 (N_3955,N_2541,N_2628);
xnor U3956 (N_3956,N_2899,N_2486);
xnor U3957 (N_3957,N_2550,N_2086);
nor U3958 (N_3958,N_2649,N_2671);
nand U3959 (N_3959,N_2971,N_2341);
or U3960 (N_3960,N_2465,N_2491);
nor U3961 (N_3961,N_2154,N_2390);
nor U3962 (N_3962,N_2984,N_2440);
or U3963 (N_3963,N_2664,N_2527);
and U3964 (N_3964,N_2170,N_2158);
nor U3965 (N_3965,N_2386,N_2732);
nand U3966 (N_3966,N_2216,N_2714);
nor U3967 (N_3967,N_2584,N_2340);
nand U3968 (N_3968,N_2704,N_2347);
nor U3969 (N_3969,N_2116,N_2198);
and U3970 (N_3970,N_2421,N_2965);
or U3971 (N_3971,N_2462,N_2090);
or U3972 (N_3972,N_2428,N_2688);
nand U3973 (N_3973,N_2277,N_2204);
nand U3974 (N_3974,N_2090,N_2817);
nand U3975 (N_3975,N_2014,N_2091);
nor U3976 (N_3976,N_2949,N_2797);
and U3977 (N_3977,N_2069,N_2895);
xor U3978 (N_3978,N_2797,N_2836);
and U3979 (N_3979,N_2288,N_2687);
or U3980 (N_3980,N_2161,N_2419);
or U3981 (N_3981,N_2706,N_2317);
xor U3982 (N_3982,N_2467,N_2477);
or U3983 (N_3983,N_2309,N_2750);
nor U3984 (N_3984,N_2653,N_2520);
or U3985 (N_3985,N_2538,N_2948);
xnor U3986 (N_3986,N_2676,N_2736);
nor U3987 (N_3987,N_2568,N_2771);
or U3988 (N_3988,N_2652,N_2298);
xor U3989 (N_3989,N_2513,N_2437);
or U3990 (N_3990,N_2084,N_2582);
nand U3991 (N_3991,N_2293,N_2607);
xor U3992 (N_3992,N_2849,N_2935);
and U3993 (N_3993,N_2021,N_2860);
xor U3994 (N_3994,N_2804,N_2859);
and U3995 (N_3995,N_2481,N_2720);
and U3996 (N_3996,N_2594,N_2418);
nand U3997 (N_3997,N_2705,N_2212);
xnor U3998 (N_3998,N_2439,N_2339);
and U3999 (N_3999,N_2209,N_2770);
and U4000 (N_4000,N_3879,N_3032);
or U4001 (N_4001,N_3489,N_3491);
xor U4002 (N_4002,N_3782,N_3091);
nand U4003 (N_4003,N_3533,N_3043);
or U4004 (N_4004,N_3900,N_3812);
xor U4005 (N_4005,N_3632,N_3529);
nand U4006 (N_4006,N_3102,N_3270);
nor U4007 (N_4007,N_3579,N_3029);
nor U4008 (N_4008,N_3890,N_3444);
or U4009 (N_4009,N_3758,N_3098);
nor U4010 (N_4010,N_3395,N_3714);
or U4011 (N_4011,N_3025,N_3298);
nand U4012 (N_4012,N_3122,N_3016);
and U4013 (N_4013,N_3795,N_3327);
or U4014 (N_4014,N_3921,N_3435);
or U4015 (N_4015,N_3648,N_3980);
or U4016 (N_4016,N_3168,N_3328);
and U4017 (N_4017,N_3382,N_3239);
or U4018 (N_4018,N_3911,N_3715);
xnor U4019 (N_4019,N_3377,N_3257);
nor U4020 (N_4020,N_3344,N_3740);
and U4021 (N_4021,N_3062,N_3502);
nand U4022 (N_4022,N_3272,N_3710);
or U4023 (N_4023,N_3954,N_3373);
xnor U4024 (N_4024,N_3517,N_3238);
and U4025 (N_4025,N_3880,N_3527);
xnor U4026 (N_4026,N_3528,N_3744);
and U4027 (N_4027,N_3903,N_3179);
nor U4028 (N_4028,N_3623,N_3271);
nor U4029 (N_4029,N_3110,N_3277);
nor U4030 (N_4030,N_3158,N_3638);
or U4031 (N_4031,N_3470,N_3707);
xnor U4032 (N_4032,N_3881,N_3213);
or U4033 (N_4033,N_3316,N_3627);
nor U4034 (N_4034,N_3588,N_3676);
nand U4035 (N_4035,N_3525,N_3495);
xnor U4036 (N_4036,N_3336,N_3656);
nor U4037 (N_4037,N_3645,N_3150);
nor U4038 (N_4038,N_3636,N_3640);
or U4039 (N_4039,N_3516,N_3453);
xor U4040 (N_4040,N_3927,N_3193);
nand U4041 (N_4041,N_3695,N_3190);
xor U4042 (N_4042,N_3819,N_3905);
nor U4043 (N_4043,N_3657,N_3616);
xnor U4044 (N_4044,N_3538,N_3133);
and U4045 (N_4045,N_3273,N_3294);
nand U4046 (N_4046,N_3814,N_3412);
and U4047 (N_4047,N_3910,N_3075);
or U4048 (N_4048,N_3416,N_3708);
nand U4049 (N_4049,N_3622,N_3671);
nor U4050 (N_4050,N_3868,N_3368);
nor U4051 (N_4051,N_3406,N_3821);
nand U4052 (N_4052,N_3978,N_3496);
xnor U4053 (N_4053,N_3914,N_3262);
xor U4054 (N_4054,N_3558,N_3006);
nand U4055 (N_4055,N_3767,N_3665);
nand U4056 (N_4056,N_3305,N_3400);
nand U4057 (N_4057,N_3263,N_3584);
nor U4058 (N_4058,N_3765,N_3661);
xor U4059 (N_4059,N_3786,N_3574);
nor U4060 (N_4060,N_3358,N_3154);
or U4061 (N_4061,N_3349,N_3654);
xor U4062 (N_4062,N_3866,N_3861);
and U4063 (N_4063,N_3383,N_3843);
nor U4064 (N_4064,N_3693,N_3136);
nand U4065 (N_4065,N_3557,N_3074);
xnor U4066 (N_4066,N_3668,N_3600);
nand U4067 (N_4067,N_3863,N_3601);
nor U4068 (N_4068,N_3899,N_3148);
nor U4069 (N_4069,N_3514,N_3418);
or U4070 (N_4070,N_3434,N_3571);
nand U4071 (N_4071,N_3176,N_3526);
nand U4072 (N_4072,N_3287,N_3051);
and U4073 (N_4073,N_3070,N_3609);
nor U4074 (N_4074,N_3572,N_3724);
xnor U4075 (N_4075,N_3066,N_3482);
nor U4076 (N_4076,N_3918,N_3149);
nand U4077 (N_4077,N_3152,N_3776);
or U4078 (N_4078,N_3332,N_3773);
or U4079 (N_4079,N_3974,N_3893);
xnor U4080 (N_4080,N_3072,N_3145);
and U4081 (N_4081,N_3803,N_3207);
nand U4082 (N_4082,N_3224,N_3991);
nand U4083 (N_4083,N_3854,N_3564);
xor U4084 (N_4084,N_3713,N_3894);
nor U4085 (N_4085,N_3490,N_3721);
nand U4086 (N_4086,N_3460,N_3583);
and U4087 (N_4087,N_3194,N_3251);
nand U4088 (N_4088,N_3858,N_3889);
and U4089 (N_4089,N_3080,N_3994);
xor U4090 (N_4090,N_3586,N_3030);
xnor U4091 (N_4091,N_3322,N_3988);
and U4092 (N_4092,N_3913,N_3604);
nand U4093 (N_4093,N_3424,N_3350);
nor U4094 (N_4094,N_3591,N_3013);
nand U4095 (N_4095,N_3473,N_3365);
or U4096 (N_4096,N_3997,N_3709);
xnor U4097 (N_4097,N_3965,N_3628);
or U4098 (N_4098,N_3275,N_3670);
nand U4099 (N_4099,N_3875,N_3679);
nor U4100 (N_4100,N_3372,N_3963);
and U4101 (N_4101,N_3820,N_3120);
nand U4102 (N_4102,N_3907,N_3521);
nor U4103 (N_4103,N_3682,N_3888);
nor U4104 (N_4104,N_3909,N_3141);
nand U4105 (N_4105,N_3433,N_3643);
or U4106 (N_4106,N_3589,N_3602);
nor U4107 (N_4107,N_3872,N_3408);
or U4108 (N_4108,N_3342,N_3220);
and U4109 (N_4109,N_3664,N_3293);
nor U4110 (N_4110,N_3598,N_3218);
or U4111 (N_4111,N_3596,N_3401);
xnor U4112 (N_4112,N_3204,N_3123);
and U4113 (N_4113,N_3097,N_3252);
xor U4114 (N_4114,N_3042,N_3303);
nand U4115 (N_4115,N_3165,N_3518);
nor U4116 (N_4116,N_3329,N_3835);
and U4117 (N_4117,N_3582,N_3335);
nor U4118 (N_4118,N_3174,N_3639);
nor U4119 (N_4119,N_3551,N_3069);
nand U4120 (N_4120,N_3736,N_3493);
or U4121 (N_4121,N_3947,N_3700);
and U4122 (N_4122,N_3107,N_3157);
nand U4123 (N_4123,N_3685,N_3807);
nor U4124 (N_4124,N_3594,N_3292);
and U4125 (N_4125,N_3090,N_3612);
nor U4126 (N_4126,N_3989,N_3983);
or U4127 (N_4127,N_3520,N_3508);
or U4128 (N_4128,N_3926,N_3092);
xor U4129 (N_4129,N_3361,N_3902);
nand U4130 (N_4130,N_3816,N_3050);
and U4131 (N_4131,N_3901,N_3403);
xor U4132 (N_4132,N_3290,N_3236);
and U4133 (N_4133,N_3569,N_3577);
xor U4134 (N_4134,N_3461,N_3229);
xor U4135 (N_4135,N_3541,N_3870);
nand U4136 (N_4136,N_3487,N_3950);
and U4137 (N_4137,N_3105,N_3924);
xor U4138 (N_4138,N_3456,N_3626);
nand U4139 (N_4139,N_3119,N_3908);
nor U4140 (N_4140,N_3146,N_3004);
and U4141 (N_4141,N_3394,N_3501);
and U4142 (N_4142,N_3333,N_3917);
nand U4143 (N_4143,N_3234,N_3512);
nor U4144 (N_4144,N_3652,N_3308);
and U4145 (N_4145,N_3566,N_3916);
or U4146 (N_4146,N_3155,N_3537);
nand U4147 (N_4147,N_3367,N_3221);
or U4148 (N_4148,N_3673,N_3667);
nor U4149 (N_4149,N_3000,N_3706);
nand U4150 (N_4150,N_3973,N_3028);
nand U4151 (N_4151,N_3937,N_3254);
xor U4152 (N_4152,N_3341,N_3912);
xnor U4153 (N_4153,N_3241,N_3100);
nand U4154 (N_4154,N_3940,N_3956);
or U4155 (N_4155,N_3620,N_3641);
or U4156 (N_4156,N_3427,N_3633);
nor U4157 (N_4157,N_3935,N_3946);
nor U4158 (N_4158,N_3180,N_3389);
xnor U4159 (N_4159,N_3058,N_3513);
nor U4160 (N_4160,N_3302,N_3167);
xnor U4161 (N_4161,N_3283,N_3892);
nand U4162 (N_4162,N_3530,N_3992);
and U4163 (N_4163,N_3445,N_3048);
xor U4164 (N_4164,N_3245,N_3339);
xnor U4165 (N_4165,N_3730,N_3701);
xor U4166 (N_4166,N_3568,N_3544);
nor U4167 (N_4167,N_3307,N_3542);
or U4168 (N_4168,N_3555,N_3166);
nor U4169 (N_4169,N_3472,N_3178);
and U4170 (N_4170,N_3304,N_3338);
and U4171 (N_4171,N_3056,N_3337);
xor U4172 (N_4172,N_3686,N_3018);
and U4173 (N_4173,N_3188,N_3015);
nor U4174 (N_4174,N_3354,N_3446);
xnor U4175 (N_4175,N_3692,N_3347);
or U4176 (N_4176,N_3126,N_3014);
or U4177 (N_4177,N_3206,N_3993);
and U4178 (N_4178,N_3431,N_3356);
nand U4179 (N_4179,N_3635,N_3702);
xnor U4180 (N_4180,N_3871,N_3480);
and U4181 (N_4181,N_3757,N_3109);
and U4182 (N_4182,N_3545,N_3198);
xnor U4183 (N_4183,N_3929,N_3862);
and U4184 (N_4184,N_3759,N_3792);
and U4185 (N_4185,N_3041,N_3053);
and U4186 (N_4186,N_3413,N_3727);
and U4187 (N_4187,N_3611,N_3524);
nand U4188 (N_4188,N_3233,N_3195);
nor U4189 (N_4189,N_3143,N_3297);
nand U4190 (N_4190,N_3306,N_3184);
nor U4191 (N_4191,N_3462,N_3312);
nor U4192 (N_4192,N_3256,N_3644);
and U4193 (N_4193,N_3440,N_3442);
and U4194 (N_4194,N_3173,N_3390);
and U4195 (N_4195,N_3982,N_3849);
and U4196 (N_4196,N_3827,N_3002);
or U4197 (N_4197,N_3138,N_3007);
xor U4198 (N_4198,N_3450,N_3919);
nor U4199 (N_4199,N_3115,N_3603);
nand U4200 (N_4200,N_3559,N_3033);
and U4201 (N_4201,N_3824,N_3887);
nand U4202 (N_4202,N_3311,N_3563);
nand U4203 (N_4203,N_3108,N_3183);
xor U4204 (N_4204,N_3610,N_3592);
or U4205 (N_4205,N_3121,N_3210);
nor U4206 (N_4206,N_3960,N_3240);
or U4207 (N_4207,N_3651,N_3464);
xnor U4208 (N_4208,N_3286,N_3718);
nor U4209 (N_4209,N_3082,N_3265);
nand U4210 (N_4210,N_3781,N_3246);
nand U4211 (N_4211,N_3959,N_3078);
xor U4212 (N_4212,N_3546,N_3852);
xnor U4213 (N_4213,N_3024,N_3019);
xor U4214 (N_4214,N_3300,N_3647);
nor U4215 (N_4215,N_3222,N_3509);
xor U4216 (N_4216,N_3877,N_3289);
or U4217 (N_4217,N_3398,N_3362);
or U4218 (N_4218,N_3585,N_3345);
or U4219 (N_4219,N_3649,N_3742);
and U4220 (N_4220,N_3248,N_3753);
xor U4221 (N_4221,N_3818,N_3500);
and U4222 (N_4222,N_3118,N_3215);
nor U4223 (N_4223,N_3379,N_3772);
or U4224 (N_4224,N_3452,N_3415);
nand U4225 (N_4225,N_3479,N_3031);
xnor U4226 (N_4226,N_3244,N_3247);
nand U4227 (N_4227,N_3185,N_3986);
nor U4228 (N_4228,N_3750,N_3055);
xor U4229 (N_4229,N_3005,N_3561);
and U4230 (N_4230,N_3192,N_3723);
nand U4231 (N_4231,N_3751,N_3429);
nand U4232 (N_4232,N_3884,N_3719);
or U4233 (N_4233,N_3079,N_3798);
and U4234 (N_4234,N_3111,N_3969);
xor U4235 (N_4235,N_3340,N_3876);
nor U4236 (N_4236,N_3567,N_3475);
or U4237 (N_4237,N_3878,N_3743);
xnor U4238 (N_4238,N_3330,N_3712);
xnor U4239 (N_4239,N_3953,N_3027);
or U4240 (N_4240,N_3681,N_3481);
or U4241 (N_4241,N_3729,N_3853);
and U4242 (N_4242,N_3531,N_3556);
xor U4243 (N_4243,N_3288,N_3381);
or U4244 (N_4244,N_3003,N_3597);
or U4245 (N_4245,N_3939,N_3351);
nor U4246 (N_4246,N_3762,N_3189);
nor U4247 (N_4247,N_3523,N_3384);
nor U4248 (N_4248,N_3883,N_3483);
xor U4249 (N_4249,N_3425,N_3313);
and U4250 (N_4250,N_3134,N_3411);
nor U4251 (N_4251,N_3223,N_3432);
xnor U4252 (N_4252,N_3933,N_3949);
or U4253 (N_4253,N_3857,N_3507);
and U4254 (N_4254,N_3366,N_3590);
or U4255 (N_4255,N_3299,N_3923);
and U4256 (N_4256,N_3739,N_3570);
nand U4257 (N_4257,N_3318,N_3216);
or U4258 (N_4258,N_3182,N_3457);
nand U4259 (N_4259,N_3404,N_3360);
xnor U4260 (N_4260,N_3067,N_3151);
or U4261 (N_4261,N_3488,N_3124);
nor U4262 (N_4262,N_3804,N_3725);
or U4263 (N_4263,N_3874,N_3439);
or U4264 (N_4264,N_3506,N_3060);
nand U4265 (N_4265,N_3310,N_3618);
nand U4266 (N_4266,N_3576,N_3607);
and U4267 (N_4267,N_3650,N_3552);
nor U4268 (N_4268,N_3451,N_3769);
or U4269 (N_4269,N_3720,N_3448);
xnor U4270 (N_4270,N_3274,N_3637);
or U4271 (N_4271,N_3137,N_3437);
nor U4272 (N_4272,N_3784,N_3698);
and U4273 (N_4273,N_3052,N_3231);
nor U4274 (N_4274,N_3282,N_3235);
nor U4275 (N_4275,N_3979,N_3915);
nand U4276 (N_4276,N_3426,N_3430);
nand U4277 (N_4277,N_3696,N_3276);
and U4278 (N_4278,N_3955,N_3653);
and U4279 (N_4279,N_3565,N_3187);
xor U4280 (N_4280,N_3793,N_3331);
and U4281 (N_4281,N_3012,N_3791);
nor U4282 (N_4282,N_3129,N_3458);
xor U4283 (N_4283,N_3175,N_3093);
nand U4284 (N_4284,N_3886,N_3226);
nand U4285 (N_4285,N_3388,N_3497);
or U4286 (N_4286,N_3117,N_3735);
nor U4287 (N_4287,N_3811,N_3957);
nand U4288 (N_4288,N_3968,N_3057);
and U4289 (N_4289,N_3353,N_3455);
or U4290 (N_4290,N_3951,N_3621);
or U4291 (N_4291,N_3212,N_3396);
or U4292 (N_4292,N_3943,N_3897);
and U4293 (N_4293,N_3799,N_3694);
nand U4294 (N_4294,N_3838,N_3970);
nor U4295 (N_4295,N_3630,N_3699);
nor U4296 (N_4296,N_3967,N_3573);
or U4297 (N_4297,N_3595,N_3071);
and U4298 (N_4298,N_3380,N_3634);
nand U4299 (N_4299,N_3617,N_3447);
nor U4300 (N_4300,N_3112,N_3385);
or U4301 (N_4301,N_3324,N_3746);
nand U4302 (N_4302,N_3454,N_3554);
xor U4303 (N_4303,N_3766,N_3466);
xor U4304 (N_4304,N_3284,N_3840);
nand U4305 (N_4305,N_3205,N_3815);
nand U4306 (N_4306,N_3785,N_3441);
xnor U4307 (N_4307,N_3089,N_3680);
nand U4308 (N_4308,N_3044,N_3443);
and U4309 (N_4309,N_3153,N_3201);
nor U4310 (N_4310,N_3140,N_3690);
nand U4311 (N_4311,N_3976,N_3219);
nor U4312 (N_4312,N_3064,N_3995);
and U4313 (N_4313,N_3659,N_3810);
and U4314 (N_4314,N_3845,N_3580);
xnor U4315 (N_4315,N_3159,N_3486);
nor U4316 (N_4316,N_3505,N_3320);
nand U4317 (N_4317,N_3186,N_3787);
nand U4318 (N_4318,N_3629,N_3823);
and U4319 (N_4319,N_3436,N_3998);
nand U4320 (N_4320,N_3761,N_3672);
nor U4321 (N_4321,N_3017,N_3774);
and U4322 (N_4322,N_3428,N_3829);
nand U4323 (N_4323,N_3510,N_3142);
or U4324 (N_4324,N_3160,N_3625);
and U4325 (N_4325,N_3386,N_3741);
and U4326 (N_4326,N_3532,N_3864);
nand U4327 (N_4327,N_3906,N_3987);
and U4328 (N_4328,N_3737,N_3608);
and U4329 (N_4329,N_3675,N_3088);
xor U4330 (N_4330,N_3036,N_3484);
and U4331 (N_4331,N_3225,N_3267);
nor U4332 (N_4332,N_3397,N_3999);
nor U4333 (N_4333,N_3749,N_3836);
nand U4334 (N_4334,N_3981,N_3095);
and U4335 (N_4335,N_3499,N_3200);
xor U4336 (N_4336,N_3208,N_3944);
nand U4337 (N_4337,N_3261,N_3731);
nand U4338 (N_4338,N_3841,N_3139);
xor U4339 (N_4339,N_3800,N_3278);
xnor U4340 (N_4340,N_3471,N_3966);
or U4341 (N_4341,N_3837,N_3717);
nand U4342 (N_4342,N_3961,N_3073);
xor U4343 (N_4343,N_3756,N_3034);
nor U4344 (N_4344,N_3021,N_3850);
nor U4345 (N_4345,N_3783,N_3230);
and U4346 (N_4346,N_3063,N_3535);
or U4347 (N_4347,N_3931,N_3655);
nand U4348 (N_4348,N_3106,N_3099);
and U4349 (N_4349,N_3407,N_3678);
and U4350 (N_4350,N_3202,N_3593);
nor U4351 (N_4351,N_3801,N_3144);
or U4352 (N_4352,N_3562,N_3511);
nand U4353 (N_4353,N_3777,N_3203);
nand U4354 (N_4354,N_3449,N_3116);
xor U4355 (N_4355,N_3260,N_3237);
nor U4356 (N_4356,N_3387,N_3920);
and U4357 (N_4357,N_3494,N_3975);
nand U4358 (N_4358,N_3227,N_3171);
xor U4359 (N_4359,N_3391,N_3291);
nor U4360 (N_4360,N_3001,N_3164);
or U4361 (N_4361,N_3355,N_3035);
xnor U4362 (N_4362,N_3778,N_3172);
or U4363 (N_4363,N_3964,N_3054);
nor U4364 (N_4364,N_3898,N_3059);
xor U4365 (N_4365,N_3832,N_3217);
xnor U4366 (N_4366,N_3962,N_3156);
nand U4367 (N_4367,N_3420,N_3677);
xor U4368 (N_4368,N_3614,N_3922);
or U4369 (N_4369,N_3972,N_3985);
and U4370 (N_4370,N_3469,N_3253);
or U4371 (N_4371,N_3323,N_3352);
and U4372 (N_4372,N_3409,N_3515);
nand U4373 (N_4373,N_3477,N_3711);
nor U4374 (N_4374,N_3476,N_3705);
xnor U4375 (N_4375,N_3605,N_3285);
and U4376 (N_4376,N_3996,N_3642);
xor U4377 (N_4377,N_3860,N_3697);
nor U4378 (N_4378,N_3045,N_3846);
nand U4379 (N_4379,N_3938,N_3301);
nor U4380 (N_4380,N_3125,N_3734);
nand U4381 (N_4381,N_3942,N_3049);
xor U4382 (N_4382,N_3687,N_3789);
nor U4383 (N_4383,N_3147,N_3296);
xor U4384 (N_4384,N_3211,N_3357);
xnor U4385 (N_4385,N_3733,N_3891);
and U4386 (N_4386,N_3728,N_3945);
nor U4387 (N_4387,N_3314,N_3258);
xor U4388 (N_4388,N_3334,N_3770);
xor U4389 (N_4389,N_3806,N_3726);
or U4390 (N_4390,N_3468,N_3393);
and U4391 (N_4391,N_3809,N_3405);
nand U4392 (N_4392,N_3348,N_3813);
or U4393 (N_4393,N_3833,N_3103);
and U4394 (N_4394,N_3410,N_3378);
and U4395 (N_4395,N_3790,N_3936);
or U4396 (N_4396,N_3259,N_3930);
and U4397 (N_4397,N_3704,N_3228);
or U4398 (N_4398,N_3805,N_3536);
nand U4399 (N_4399,N_3780,N_3309);
nand U4400 (N_4400,N_3519,N_3904);
nand U4401 (N_4401,N_3076,N_3232);
xnor U4402 (N_4402,N_3161,N_3086);
nor U4403 (N_4403,N_3022,N_3885);
or U4404 (N_4404,N_3419,N_3747);
nand U4405 (N_4405,N_3127,N_3842);
xnor U4406 (N_4406,N_3660,N_3011);
nor U4407 (N_4407,N_3703,N_3752);
nor U4408 (N_4408,N_3094,N_3825);
xor U4409 (N_4409,N_3763,N_3169);
nand U4410 (N_4410,N_3038,N_3279);
and U4411 (N_4411,N_3925,N_3748);
nand U4412 (N_4412,N_3859,N_3896);
nor U4413 (N_4413,N_3851,N_3077);
and U4414 (N_4414,N_3280,N_3374);
and U4415 (N_4415,N_3392,N_3738);
nand U4416 (N_4416,N_3130,N_3855);
and U4417 (N_4417,N_3873,N_3065);
nor U4418 (N_4418,N_3485,N_3463);
and U4419 (N_4419,N_3421,N_3587);
xnor U4420 (N_4420,N_3008,N_3465);
nand U4421 (N_4421,N_3423,N_3266);
xnor U4422 (N_4422,N_3839,N_3826);
xnor U4423 (N_4423,N_3068,N_3243);
nand U4424 (N_4424,N_3163,N_3895);
and U4425 (N_4425,N_3135,N_3177);
xnor U4426 (N_4426,N_3321,N_3376);
xor U4427 (N_4427,N_3666,N_3856);
nor U4428 (N_4428,N_3199,N_3547);
nand U4429 (N_4429,N_3295,N_3689);
and U4430 (N_4430,N_3788,N_3534);
or U4431 (N_4431,N_3503,N_3847);
and U4432 (N_4432,N_3663,N_3369);
and U4433 (N_4433,N_3319,N_3414);
or U4434 (N_4434,N_3662,N_3869);
nor U4435 (N_4435,N_3802,N_3264);
nor U4436 (N_4436,N_3315,N_3317);
nor U4437 (N_4437,N_3540,N_3478);
nor U4438 (N_4438,N_3459,N_3834);
or U4439 (N_4439,N_3948,N_3504);
nor U4440 (N_4440,N_3615,N_3581);
nand U4441 (N_4441,N_3755,N_3669);
or U4442 (N_4442,N_3249,N_3754);
nor U4443 (N_4443,N_3745,N_3364);
or U4444 (N_4444,N_3422,N_3242);
and U4445 (N_4445,N_3732,N_3771);
or U4446 (N_4446,N_3326,N_3359);
and U4447 (N_4447,N_3467,N_3114);
nor U4448 (N_4448,N_3363,N_3191);
xor U4449 (N_4449,N_3269,N_3087);
nand U4450 (N_4450,N_3658,N_3085);
xnor U4451 (N_4451,N_3081,N_3325);
xor U4452 (N_4452,N_3683,N_3402);
nand U4453 (N_4453,N_3399,N_3197);
nand U4454 (N_4454,N_3848,N_3631);
or U4455 (N_4455,N_3096,N_3560);
or U4456 (N_4456,N_3684,N_3128);
xnor U4457 (N_4457,N_3779,N_3474);
nor U4458 (N_4458,N_3214,N_3047);
nor U4459 (N_4459,N_3831,N_3844);
xor U4460 (N_4460,N_3599,N_3250);
and U4461 (N_4461,N_3984,N_3797);
or U4462 (N_4462,N_3830,N_3775);
nor U4463 (N_4463,N_3343,N_3865);
nor U4464 (N_4464,N_3764,N_3104);
nand U4465 (N_4465,N_3162,N_3255);
or U4466 (N_4466,N_3822,N_3674);
nand U4467 (N_4467,N_3794,N_3020);
nand U4468 (N_4468,N_3928,N_3934);
nand U4469 (N_4469,N_3281,N_3131);
nand U4470 (N_4470,N_3613,N_3026);
nand U4471 (N_4471,N_3796,N_3539);
nand U4472 (N_4472,N_3417,N_3646);
nand U4473 (N_4473,N_3543,N_3619);
nor U4474 (N_4474,N_3578,N_3941);
nand U4475 (N_4475,N_3688,N_3932);
nor U4476 (N_4476,N_3023,N_3375);
xnor U4477 (N_4477,N_3952,N_3196);
xor U4478 (N_4478,N_3716,N_3037);
nand U4479 (N_4479,N_3808,N_3209);
nand U4480 (N_4480,N_3882,N_3575);
and U4481 (N_4481,N_3977,N_3817);
xnor U4482 (N_4482,N_3268,N_3550);
nor U4483 (N_4483,N_3522,N_3548);
or U4484 (N_4484,N_3760,N_3132);
nor U4485 (N_4485,N_3039,N_3867);
nor U4486 (N_4486,N_3009,N_3606);
nor U4487 (N_4487,N_3553,N_3370);
and U4488 (N_4488,N_3371,N_3346);
and U4489 (N_4489,N_3101,N_3768);
nor U4490 (N_4490,N_3498,N_3549);
or U4491 (N_4491,N_3958,N_3438);
xnor U4492 (N_4492,N_3170,N_3061);
nand U4493 (N_4493,N_3624,N_3971);
xnor U4494 (N_4494,N_3040,N_3691);
or U4495 (N_4495,N_3083,N_3084);
or U4496 (N_4496,N_3990,N_3181);
nand U4497 (N_4497,N_3492,N_3113);
or U4498 (N_4498,N_3046,N_3828);
xor U4499 (N_4499,N_3010,N_3722);
xnor U4500 (N_4500,N_3231,N_3288);
nor U4501 (N_4501,N_3305,N_3013);
and U4502 (N_4502,N_3525,N_3739);
xnor U4503 (N_4503,N_3807,N_3106);
or U4504 (N_4504,N_3359,N_3392);
and U4505 (N_4505,N_3150,N_3201);
and U4506 (N_4506,N_3833,N_3429);
or U4507 (N_4507,N_3144,N_3737);
nor U4508 (N_4508,N_3095,N_3723);
nand U4509 (N_4509,N_3827,N_3077);
and U4510 (N_4510,N_3465,N_3637);
nor U4511 (N_4511,N_3865,N_3335);
xnor U4512 (N_4512,N_3682,N_3118);
nand U4513 (N_4513,N_3358,N_3921);
nand U4514 (N_4514,N_3738,N_3370);
nor U4515 (N_4515,N_3833,N_3524);
and U4516 (N_4516,N_3041,N_3917);
nand U4517 (N_4517,N_3173,N_3300);
xnor U4518 (N_4518,N_3514,N_3634);
or U4519 (N_4519,N_3543,N_3024);
or U4520 (N_4520,N_3984,N_3625);
or U4521 (N_4521,N_3855,N_3599);
or U4522 (N_4522,N_3947,N_3955);
nand U4523 (N_4523,N_3774,N_3657);
xnor U4524 (N_4524,N_3532,N_3596);
xor U4525 (N_4525,N_3289,N_3385);
or U4526 (N_4526,N_3352,N_3375);
nor U4527 (N_4527,N_3522,N_3153);
and U4528 (N_4528,N_3607,N_3562);
or U4529 (N_4529,N_3437,N_3431);
nand U4530 (N_4530,N_3882,N_3414);
and U4531 (N_4531,N_3047,N_3846);
nand U4532 (N_4532,N_3937,N_3282);
or U4533 (N_4533,N_3622,N_3039);
xnor U4534 (N_4534,N_3463,N_3381);
nand U4535 (N_4535,N_3435,N_3501);
and U4536 (N_4536,N_3252,N_3583);
or U4537 (N_4537,N_3911,N_3792);
nand U4538 (N_4538,N_3145,N_3050);
and U4539 (N_4539,N_3746,N_3058);
nor U4540 (N_4540,N_3667,N_3171);
xnor U4541 (N_4541,N_3329,N_3247);
nor U4542 (N_4542,N_3550,N_3304);
nor U4543 (N_4543,N_3943,N_3937);
nor U4544 (N_4544,N_3917,N_3278);
and U4545 (N_4545,N_3998,N_3431);
nand U4546 (N_4546,N_3972,N_3173);
nand U4547 (N_4547,N_3183,N_3079);
xnor U4548 (N_4548,N_3033,N_3318);
nor U4549 (N_4549,N_3324,N_3847);
and U4550 (N_4550,N_3635,N_3129);
xnor U4551 (N_4551,N_3153,N_3550);
nand U4552 (N_4552,N_3023,N_3395);
and U4553 (N_4553,N_3583,N_3110);
xnor U4554 (N_4554,N_3655,N_3039);
and U4555 (N_4555,N_3678,N_3450);
xor U4556 (N_4556,N_3392,N_3689);
nor U4557 (N_4557,N_3008,N_3109);
and U4558 (N_4558,N_3051,N_3144);
and U4559 (N_4559,N_3923,N_3859);
or U4560 (N_4560,N_3988,N_3074);
and U4561 (N_4561,N_3498,N_3187);
nor U4562 (N_4562,N_3373,N_3145);
nor U4563 (N_4563,N_3344,N_3978);
nor U4564 (N_4564,N_3710,N_3192);
nand U4565 (N_4565,N_3321,N_3476);
and U4566 (N_4566,N_3969,N_3029);
nand U4567 (N_4567,N_3372,N_3855);
xor U4568 (N_4568,N_3766,N_3027);
and U4569 (N_4569,N_3097,N_3424);
xnor U4570 (N_4570,N_3218,N_3440);
or U4571 (N_4571,N_3387,N_3645);
nor U4572 (N_4572,N_3937,N_3620);
or U4573 (N_4573,N_3168,N_3265);
or U4574 (N_4574,N_3933,N_3002);
nor U4575 (N_4575,N_3317,N_3147);
nand U4576 (N_4576,N_3335,N_3666);
xnor U4577 (N_4577,N_3304,N_3788);
nor U4578 (N_4578,N_3654,N_3195);
nand U4579 (N_4579,N_3540,N_3406);
nand U4580 (N_4580,N_3347,N_3037);
and U4581 (N_4581,N_3497,N_3164);
xor U4582 (N_4582,N_3706,N_3215);
and U4583 (N_4583,N_3871,N_3730);
or U4584 (N_4584,N_3807,N_3654);
xnor U4585 (N_4585,N_3544,N_3580);
nand U4586 (N_4586,N_3694,N_3753);
or U4587 (N_4587,N_3875,N_3267);
nand U4588 (N_4588,N_3031,N_3976);
xor U4589 (N_4589,N_3287,N_3105);
and U4590 (N_4590,N_3184,N_3584);
nor U4591 (N_4591,N_3127,N_3848);
xnor U4592 (N_4592,N_3111,N_3965);
xor U4593 (N_4593,N_3018,N_3795);
xor U4594 (N_4594,N_3976,N_3142);
or U4595 (N_4595,N_3488,N_3173);
nor U4596 (N_4596,N_3411,N_3329);
and U4597 (N_4597,N_3783,N_3499);
xnor U4598 (N_4598,N_3267,N_3107);
xnor U4599 (N_4599,N_3259,N_3372);
and U4600 (N_4600,N_3263,N_3300);
nand U4601 (N_4601,N_3428,N_3540);
and U4602 (N_4602,N_3294,N_3123);
and U4603 (N_4603,N_3005,N_3765);
nand U4604 (N_4604,N_3111,N_3944);
or U4605 (N_4605,N_3431,N_3017);
and U4606 (N_4606,N_3403,N_3678);
or U4607 (N_4607,N_3413,N_3790);
xor U4608 (N_4608,N_3207,N_3254);
or U4609 (N_4609,N_3499,N_3279);
nand U4610 (N_4610,N_3093,N_3996);
and U4611 (N_4611,N_3488,N_3327);
xor U4612 (N_4612,N_3113,N_3782);
nor U4613 (N_4613,N_3052,N_3900);
nand U4614 (N_4614,N_3256,N_3835);
nor U4615 (N_4615,N_3475,N_3396);
and U4616 (N_4616,N_3266,N_3765);
or U4617 (N_4617,N_3411,N_3734);
nand U4618 (N_4618,N_3576,N_3109);
and U4619 (N_4619,N_3441,N_3311);
or U4620 (N_4620,N_3449,N_3408);
nor U4621 (N_4621,N_3917,N_3484);
and U4622 (N_4622,N_3915,N_3552);
xnor U4623 (N_4623,N_3765,N_3712);
nor U4624 (N_4624,N_3203,N_3667);
xnor U4625 (N_4625,N_3063,N_3696);
nor U4626 (N_4626,N_3444,N_3802);
and U4627 (N_4627,N_3273,N_3572);
xor U4628 (N_4628,N_3141,N_3226);
nor U4629 (N_4629,N_3106,N_3589);
or U4630 (N_4630,N_3912,N_3600);
or U4631 (N_4631,N_3511,N_3053);
nand U4632 (N_4632,N_3816,N_3789);
or U4633 (N_4633,N_3743,N_3919);
or U4634 (N_4634,N_3370,N_3118);
nand U4635 (N_4635,N_3551,N_3400);
xnor U4636 (N_4636,N_3322,N_3636);
nor U4637 (N_4637,N_3618,N_3997);
nor U4638 (N_4638,N_3601,N_3814);
or U4639 (N_4639,N_3655,N_3331);
nand U4640 (N_4640,N_3818,N_3534);
or U4641 (N_4641,N_3634,N_3490);
and U4642 (N_4642,N_3863,N_3600);
or U4643 (N_4643,N_3583,N_3461);
nand U4644 (N_4644,N_3598,N_3713);
nand U4645 (N_4645,N_3153,N_3423);
or U4646 (N_4646,N_3385,N_3708);
nor U4647 (N_4647,N_3226,N_3299);
nand U4648 (N_4648,N_3383,N_3836);
or U4649 (N_4649,N_3481,N_3541);
nand U4650 (N_4650,N_3895,N_3396);
nand U4651 (N_4651,N_3856,N_3836);
or U4652 (N_4652,N_3031,N_3442);
nand U4653 (N_4653,N_3111,N_3268);
and U4654 (N_4654,N_3647,N_3417);
and U4655 (N_4655,N_3581,N_3844);
nor U4656 (N_4656,N_3257,N_3867);
nor U4657 (N_4657,N_3246,N_3791);
xor U4658 (N_4658,N_3415,N_3331);
and U4659 (N_4659,N_3353,N_3140);
or U4660 (N_4660,N_3394,N_3667);
nand U4661 (N_4661,N_3936,N_3317);
xor U4662 (N_4662,N_3159,N_3899);
or U4663 (N_4663,N_3834,N_3098);
xnor U4664 (N_4664,N_3988,N_3851);
and U4665 (N_4665,N_3329,N_3449);
nor U4666 (N_4666,N_3557,N_3853);
nor U4667 (N_4667,N_3862,N_3335);
xor U4668 (N_4668,N_3059,N_3372);
nand U4669 (N_4669,N_3589,N_3235);
or U4670 (N_4670,N_3256,N_3794);
nor U4671 (N_4671,N_3109,N_3754);
nand U4672 (N_4672,N_3768,N_3994);
nor U4673 (N_4673,N_3698,N_3427);
nand U4674 (N_4674,N_3645,N_3794);
or U4675 (N_4675,N_3060,N_3092);
and U4676 (N_4676,N_3282,N_3828);
nor U4677 (N_4677,N_3566,N_3336);
nand U4678 (N_4678,N_3835,N_3593);
nand U4679 (N_4679,N_3249,N_3950);
or U4680 (N_4680,N_3796,N_3789);
nor U4681 (N_4681,N_3740,N_3287);
nand U4682 (N_4682,N_3239,N_3887);
or U4683 (N_4683,N_3999,N_3468);
nand U4684 (N_4684,N_3713,N_3859);
xnor U4685 (N_4685,N_3826,N_3833);
or U4686 (N_4686,N_3238,N_3056);
nor U4687 (N_4687,N_3673,N_3630);
xnor U4688 (N_4688,N_3618,N_3911);
nor U4689 (N_4689,N_3919,N_3011);
nand U4690 (N_4690,N_3533,N_3834);
xnor U4691 (N_4691,N_3189,N_3396);
xor U4692 (N_4692,N_3324,N_3977);
nor U4693 (N_4693,N_3408,N_3885);
xor U4694 (N_4694,N_3020,N_3624);
and U4695 (N_4695,N_3080,N_3509);
nand U4696 (N_4696,N_3639,N_3328);
xnor U4697 (N_4697,N_3807,N_3354);
nor U4698 (N_4698,N_3146,N_3768);
xor U4699 (N_4699,N_3996,N_3934);
nand U4700 (N_4700,N_3515,N_3084);
xor U4701 (N_4701,N_3134,N_3974);
nor U4702 (N_4702,N_3860,N_3951);
nand U4703 (N_4703,N_3327,N_3421);
nand U4704 (N_4704,N_3593,N_3664);
nor U4705 (N_4705,N_3292,N_3647);
and U4706 (N_4706,N_3066,N_3774);
xor U4707 (N_4707,N_3231,N_3805);
xnor U4708 (N_4708,N_3317,N_3507);
or U4709 (N_4709,N_3327,N_3110);
nand U4710 (N_4710,N_3812,N_3452);
or U4711 (N_4711,N_3670,N_3841);
nand U4712 (N_4712,N_3380,N_3009);
or U4713 (N_4713,N_3499,N_3739);
nand U4714 (N_4714,N_3028,N_3866);
nor U4715 (N_4715,N_3313,N_3874);
and U4716 (N_4716,N_3485,N_3293);
nor U4717 (N_4717,N_3341,N_3956);
nor U4718 (N_4718,N_3408,N_3078);
and U4719 (N_4719,N_3088,N_3862);
or U4720 (N_4720,N_3243,N_3806);
or U4721 (N_4721,N_3776,N_3813);
or U4722 (N_4722,N_3859,N_3864);
xor U4723 (N_4723,N_3667,N_3619);
nand U4724 (N_4724,N_3776,N_3506);
xor U4725 (N_4725,N_3414,N_3160);
nor U4726 (N_4726,N_3573,N_3511);
and U4727 (N_4727,N_3068,N_3973);
or U4728 (N_4728,N_3400,N_3333);
xor U4729 (N_4729,N_3241,N_3842);
and U4730 (N_4730,N_3977,N_3630);
nor U4731 (N_4731,N_3922,N_3871);
nand U4732 (N_4732,N_3187,N_3033);
xnor U4733 (N_4733,N_3810,N_3164);
nor U4734 (N_4734,N_3379,N_3344);
nor U4735 (N_4735,N_3918,N_3625);
nand U4736 (N_4736,N_3251,N_3025);
or U4737 (N_4737,N_3463,N_3740);
or U4738 (N_4738,N_3844,N_3975);
and U4739 (N_4739,N_3613,N_3286);
nand U4740 (N_4740,N_3924,N_3705);
xnor U4741 (N_4741,N_3294,N_3660);
xor U4742 (N_4742,N_3094,N_3594);
or U4743 (N_4743,N_3554,N_3489);
xor U4744 (N_4744,N_3563,N_3395);
xnor U4745 (N_4745,N_3938,N_3957);
and U4746 (N_4746,N_3562,N_3661);
nand U4747 (N_4747,N_3376,N_3827);
xor U4748 (N_4748,N_3335,N_3942);
or U4749 (N_4749,N_3558,N_3923);
or U4750 (N_4750,N_3599,N_3141);
and U4751 (N_4751,N_3350,N_3221);
xor U4752 (N_4752,N_3595,N_3913);
nand U4753 (N_4753,N_3235,N_3542);
nand U4754 (N_4754,N_3947,N_3697);
or U4755 (N_4755,N_3656,N_3031);
nor U4756 (N_4756,N_3263,N_3742);
nand U4757 (N_4757,N_3758,N_3734);
nand U4758 (N_4758,N_3800,N_3810);
or U4759 (N_4759,N_3152,N_3411);
xor U4760 (N_4760,N_3261,N_3896);
xnor U4761 (N_4761,N_3472,N_3789);
nor U4762 (N_4762,N_3296,N_3346);
nand U4763 (N_4763,N_3240,N_3733);
xnor U4764 (N_4764,N_3245,N_3702);
nand U4765 (N_4765,N_3728,N_3423);
nor U4766 (N_4766,N_3091,N_3698);
nand U4767 (N_4767,N_3003,N_3043);
or U4768 (N_4768,N_3170,N_3096);
and U4769 (N_4769,N_3071,N_3092);
and U4770 (N_4770,N_3836,N_3361);
xor U4771 (N_4771,N_3447,N_3651);
nand U4772 (N_4772,N_3862,N_3767);
and U4773 (N_4773,N_3688,N_3568);
nor U4774 (N_4774,N_3598,N_3627);
xor U4775 (N_4775,N_3807,N_3213);
nand U4776 (N_4776,N_3705,N_3411);
xnor U4777 (N_4777,N_3304,N_3571);
and U4778 (N_4778,N_3098,N_3061);
and U4779 (N_4779,N_3483,N_3779);
nand U4780 (N_4780,N_3397,N_3146);
xor U4781 (N_4781,N_3463,N_3304);
and U4782 (N_4782,N_3287,N_3229);
xnor U4783 (N_4783,N_3242,N_3774);
nand U4784 (N_4784,N_3453,N_3851);
nor U4785 (N_4785,N_3392,N_3448);
and U4786 (N_4786,N_3373,N_3987);
nor U4787 (N_4787,N_3321,N_3962);
nand U4788 (N_4788,N_3944,N_3823);
nand U4789 (N_4789,N_3028,N_3987);
nand U4790 (N_4790,N_3275,N_3168);
or U4791 (N_4791,N_3274,N_3668);
or U4792 (N_4792,N_3943,N_3892);
xor U4793 (N_4793,N_3611,N_3735);
nand U4794 (N_4794,N_3156,N_3815);
xor U4795 (N_4795,N_3645,N_3876);
and U4796 (N_4796,N_3790,N_3024);
and U4797 (N_4797,N_3447,N_3256);
nand U4798 (N_4798,N_3656,N_3172);
xnor U4799 (N_4799,N_3104,N_3077);
nand U4800 (N_4800,N_3753,N_3261);
xnor U4801 (N_4801,N_3179,N_3316);
nor U4802 (N_4802,N_3243,N_3905);
and U4803 (N_4803,N_3048,N_3486);
xnor U4804 (N_4804,N_3991,N_3968);
xor U4805 (N_4805,N_3847,N_3273);
nand U4806 (N_4806,N_3183,N_3642);
nand U4807 (N_4807,N_3607,N_3849);
nor U4808 (N_4808,N_3665,N_3446);
nor U4809 (N_4809,N_3484,N_3062);
nand U4810 (N_4810,N_3027,N_3694);
xor U4811 (N_4811,N_3949,N_3499);
or U4812 (N_4812,N_3903,N_3784);
or U4813 (N_4813,N_3840,N_3499);
nor U4814 (N_4814,N_3523,N_3705);
nand U4815 (N_4815,N_3551,N_3604);
nand U4816 (N_4816,N_3986,N_3806);
nor U4817 (N_4817,N_3590,N_3510);
nand U4818 (N_4818,N_3359,N_3595);
xor U4819 (N_4819,N_3225,N_3736);
xor U4820 (N_4820,N_3979,N_3277);
xnor U4821 (N_4821,N_3675,N_3702);
and U4822 (N_4822,N_3427,N_3347);
and U4823 (N_4823,N_3404,N_3720);
or U4824 (N_4824,N_3960,N_3309);
and U4825 (N_4825,N_3183,N_3798);
xnor U4826 (N_4826,N_3869,N_3041);
and U4827 (N_4827,N_3497,N_3883);
nor U4828 (N_4828,N_3076,N_3793);
and U4829 (N_4829,N_3070,N_3227);
xor U4830 (N_4830,N_3119,N_3257);
nor U4831 (N_4831,N_3975,N_3819);
nand U4832 (N_4832,N_3583,N_3637);
and U4833 (N_4833,N_3786,N_3121);
xnor U4834 (N_4834,N_3238,N_3906);
or U4835 (N_4835,N_3935,N_3693);
or U4836 (N_4836,N_3403,N_3914);
and U4837 (N_4837,N_3443,N_3039);
xor U4838 (N_4838,N_3872,N_3509);
nor U4839 (N_4839,N_3212,N_3138);
nand U4840 (N_4840,N_3321,N_3697);
xnor U4841 (N_4841,N_3962,N_3417);
nor U4842 (N_4842,N_3736,N_3035);
xnor U4843 (N_4843,N_3398,N_3468);
or U4844 (N_4844,N_3897,N_3076);
nand U4845 (N_4845,N_3653,N_3952);
and U4846 (N_4846,N_3321,N_3199);
xnor U4847 (N_4847,N_3203,N_3551);
nand U4848 (N_4848,N_3218,N_3236);
xnor U4849 (N_4849,N_3787,N_3655);
or U4850 (N_4850,N_3068,N_3169);
xnor U4851 (N_4851,N_3118,N_3319);
or U4852 (N_4852,N_3936,N_3333);
and U4853 (N_4853,N_3346,N_3513);
and U4854 (N_4854,N_3650,N_3769);
nand U4855 (N_4855,N_3437,N_3846);
nor U4856 (N_4856,N_3573,N_3118);
nor U4857 (N_4857,N_3476,N_3377);
and U4858 (N_4858,N_3084,N_3661);
nor U4859 (N_4859,N_3342,N_3742);
and U4860 (N_4860,N_3948,N_3560);
xnor U4861 (N_4861,N_3469,N_3626);
xnor U4862 (N_4862,N_3075,N_3941);
xnor U4863 (N_4863,N_3884,N_3158);
or U4864 (N_4864,N_3329,N_3435);
nor U4865 (N_4865,N_3121,N_3003);
xnor U4866 (N_4866,N_3803,N_3809);
and U4867 (N_4867,N_3474,N_3369);
nor U4868 (N_4868,N_3373,N_3111);
nand U4869 (N_4869,N_3445,N_3346);
nor U4870 (N_4870,N_3404,N_3811);
xnor U4871 (N_4871,N_3591,N_3990);
nand U4872 (N_4872,N_3386,N_3578);
xnor U4873 (N_4873,N_3316,N_3169);
or U4874 (N_4874,N_3097,N_3178);
or U4875 (N_4875,N_3001,N_3419);
and U4876 (N_4876,N_3688,N_3705);
nand U4877 (N_4877,N_3590,N_3732);
nand U4878 (N_4878,N_3972,N_3268);
nand U4879 (N_4879,N_3066,N_3471);
and U4880 (N_4880,N_3021,N_3926);
and U4881 (N_4881,N_3393,N_3382);
xor U4882 (N_4882,N_3976,N_3133);
nand U4883 (N_4883,N_3595,N_3596);
and U4884 (N_4884,N_3010,N_3862);
or U4885 (N_4885,N_3538,N_3280);
or U4886 (N_4886,N_3358,N_3981);
xnor U4887 (N_4887,N_3618,N_3759);
xnor U4888 (N_4888,N_3544,N_3368);
or U4889 (N_4889,N_3983,N_3606);
or U4890 (N_4890,N_3585,N_3701);
and U4891 (N_4891,N_3062,N_3305);
or U4892 (N_4892,N_3213,N_3560);
and U4893 (N_4893,N_3919,N_3147);
xor U4894 (N_4894,N_3009,N_3865);
xnor U4895 (N_4895,N_3196,N_3293);
nand U4896 (N_4896,N_3220,N_3932);
nor U4897 (N_4897,N_3327,N_3906);
nand U4898 (N_4898,N_3543,N_3341);
xor U4899 (N_4899,N_3567,N_3823);
or U4900 (N_4900,N_3499,N_3882);
and U4901 (N_4901,N_3657,N_3328);
nor U4902 (N_4902,N_3946,N_3374);
xnor U4903 (N_4903,N_3337,N_3373);
and U4904 (N_4904,N_3489,N_3648);
and U4905 (N_4905,N_3013,N_3923);
and U4906 (N_4906,N_3043,N_3517);
and U4907 (N_4907,N_3329,N_3512);
nand U4908 (N_4908,N_3604,N_3275);
and U4909 (N_4909,N_3902,N_3724);
or U4910 (N_4910,N_3950,N_3952);
nand U4911 (N_4911,N_3602,N_3960);
or U4912 (N_4912,N_3292,N_3692);
xor U4913 (N_4913,N_3258,N_3584);
nor U4914 (N_4914,N_3027,N_3330);
nor U4915 (N_4915,N_3230,N_3347);
xnor U4916 (N_4916,N_3007,N_3869);
xor U4917 (N_4917,N_3397,N_3995);
or U4918 (N_4918,N_3252,N_3668);
or U4919 (N_4919,N_3455,N_3848);
xor U4920 (N_4920,N_3474,N_3468);
xnor U4921 (N_4921,N_3678,N_3864);
xnor U4922 (N_4922,N_3703,N_3705);
or U4923 (N_4923,N_3304,N_3720);
xor U4924 (N_4924,N_3737,N_3790);
or U4925 (N_4925,N_3767,N_3921);
xor U4926 (N_4926,N_3839,N_3001);
or U4927 (N_4927,N_3284,N_3735);
and U4928 (N_4928,N_3163,N_3362);
xnor U4929 (N_4929,N_3217,N_3116);
or U4930 (N_4930,N_3915,N_3211);
nand U4931 (N_4931,N_3790,N_3180);
or U4932 (N_4932,N_3459,N_3743);
nor U4933 (N_4933,N_3617,N_3101);
and U4934 (N_4934,N_3909,N_3847);
xor U4935 (N_4935,N_3976,N_3660);
nand U4936 (N_4936,N_3582,N_3317);
nor U4937 (N_4937,N_3227,N_3441);
nor U4938 (N_4938,N_3918,N_3638);
xnor U4939 (N_4939,N_3025,N_3333);
nand U4940 (N_4940,N_3877,N_3148);
and U4941 (N_4941,N_3264,N_3968);
and U4942 (N_4942,N_3736,N_3566);
or U4943 (N_4943,N_3810,N_3049);
or U4944 (N_4944,N_3093,N_3839);
nand U4945 (N_4945,N_3980,N_3613);
or U4946 (N_4946,N_3392,N_3938);
and U4947 (N_4947,N_3128,N_3962);
and U4948 (N_4948,N_3607,N_3808);
and U4949 (N_4949,N_3984,N_3590);
nand U4950 (N_4950,N_3865,N_3090);
and U4951 (N_4951,N_3393,N_3580);
xor U4952 (N_4952,N_3405,N_3401);
nor U4953 (N_4953,N_3422,N_3555);
and U4954 (N_4954,N_3099,N_3713);
xnor U4955 (N_4955,N_3641,N_3434);
nand U4956 (N_4956,N_3104,N_3134);
or U4957 (N_4957,N_3029,N_3815);
or U4958 (N_4958,N_3602,N_3887);
or U4959 (N_4959,N_3888,N_3742);
nor U4960 (N_4960,N_3375,N_3956);
nor U4961 (N_4961,N_3948,N_3751);
nor U4962 (N_4962,N_3040,N_3983);
xnor U4963 (N_4963,N_3263,N_3298);
and U4964 (N_4964,N_3653,N_3826);
or U4965 (N_4965,N_3971,N_3161);
or U4966 (N_4966,N_3893,N_3664);
nand U4967 (N_4967,N_3118,N_3911);
or U4968 (N_4968,N_3963,N_3080);
nand U4969 (N_4969,N_3065,N_3182);
or U4970 (N_4970,N_3072,N_3925);
xor U4971 (N_4971,N_3751,N_3248);
nand U4972 (N_4972,N_3106,N_3300);
or U4973 (N_4973,N_3980,N_3404);
or U4974 (N_4974,N_3516,N_3502);
or U4975 (N_4975,N_3106,N_3431);
or U4976 (N_4976,N_3035,N_3409);
xnor U4977 (N_4977,N_3578,N_3032);
nor U4978 (N_4978,N_3696,N_3839);
nand U4979 (N_4979,N_3025,N_3232);
and U4980 (N_4980,N_3411,N_3075);
nor U4981 (N_4981,N_3235,N_3221);
nand U4982 (N_4982,N_3669,N_3364);
and U4983 (N_4983,N_3314,N_3517);
and U4984 (N_4984,N_3403,N_3844);
nand U4985 (N_4985,N_3836,N_3520);
and U4986 (N_4986,N_3251,N_3057);
and U4987 (N_4987,N_3597,N_3810);
nand U4988 (N_4988,N_3612,N_3171);
nand U4989 (N_4989,N_3593,N_3974);
nor U4990 (N_4990,N_3645,N_3489);
and U4991 (N_4991,N_3757,N_3283);
nor U4992 (N_4992,N_3125,N_3356);
or U4993 (N_4993,N_3821,N_3379);
or U4994 (N_4994,N_3565,N_3620);
xnor U4995 (N_4995,N_3629,N_3575);
nand U4996 (N_4996,N_3545,N_3351);
nor U4997 (N_4997,N_3646,N_3328);
xor U4998 (N_4998,N_3567,N_3269);
and U4999 (N_4999,N_3226,N_3276);
or U5000 (N_5000,N_4356,N_4735);
nor U5001 (N_5001,N_4746,N_4681);
or U5002 (N_5002,N_4352,N_4239);
or U5003 (N_5003,N_4864,N_4678);
xnor U5004 (N_5004,N_4748,N_4092);
or U5005 (N_5005,N_4299,N_4667);
xnor U5006 (N_5006,N_4599,N_4258);
and U5007 (N_5007,N_4710,N_4884);
and U5008 (N_5008,N_4097,N_4665);
and U5009 (N_5009,N_4605,N_4608);
and U5010 (N_5010,N_4272,N_4777);
and U5011 (N_5011,N_4377,N_4195);
and U5012 (N_5012,N_4270,N_4187);
nand U5013 (N_5013,N_4213,N_4883);
nand U5014 (N_5014,N_4370,N_4996);
or U5015 (N_5015,N_4703,N_4968);
nand U5016 (N_5016,N_4277,N_4330);
and U5017 (N_5017,N_4516,N_4953);
or U5018 (N_5018,N_4985,N_4829);
or U5019 (N_5019,N_4128,N_4569);
xor U5020 (N_5020,N_4933,N_4276);
and U5021 (N_5021,N_4631,N_4344);
and U5022 (N_5022,N_4408,N_4707);
nor U5023 (N_5023,N_4298,N_4168);
nand U5024 (N_5024,N_4124,N_4300);
or U5025 (N_5025,N_4692,N_4436);
nand U5026 (N_5026,N_4753,N_4926);
and U5027 (N_5027,N_4882,N_4487);
and U5028 (N_5028,N_4222,N_4910);
and U5029 (N_5029,N_4798,N_4456);
xor U5030 (N_5030,N_4254,N_4016);
or U5031 (N_5031,N_4020,N_4078);
and U5032 (N_5032,N_4334,N_4028);
or U5033 (N_5033,N_4257,N_4190);
xnor U5034 (N_5034,N_4642,N_4717);
xnor U5035 (N_5035,N_4267,N_4034);
nand U5036 (N_5036,N_4694,N_4649);
nor U5037 (N_5037,N_4853,N_4689);
xnor U5038 (N_5038,N_4747,N_4768);
nand U5039 (N_5039,N_4009,N_4443);
xor U5040 (N_5040,N_4363,N_4463);
nor U5041 (N_5041,N_4205,N_4314);
and U5042 (N_5042,N_4739,N_4137);
nor U5043 (N_5043,N_4148,N_4900);
nand U5044 (N_5044,N_4297,N_4350);
nand U5045 (N_5045,N_4003,N_4947);
xor U5046 (N_5046,N_4627,N_4194);
and U5047 (N_5047,N_4042,N_4146);
xor U5048 (N_5048,N_4371,N_4030);
xnor U5049 (N_5049,N_4616,N_4368);
or U5050 (N_5050,N_4155,N_4952);
or U5051 (N_5051,N_4074,N_4278);
xor U5052 (N_5052,N_4850,N_4779);
or U5053 (N_5053,N_4607,N_4970);
and U5054 (N_5054,N_4211,N_4560);
xor U5055 (N_5055,N_4957,N_4000);
or U5056 (N_5056,N_4865,N_4388);
or U5057 (N_5057,N_4564,N_4675);
nor U5058 (N_5058,N_4134,N_4818);
or U5059 (N_5059,N_4058,N_4801);
and U5060 (N_5060,N_4082,N_4696);
nand U5061 (N_5061,N_4365,N_4986);
or U5062 (N_5062,N_4790,N_4342);
and U5063 (N_5063,N_4907,N_4328);
nor U5064 (N_5064,N_4052,N_4458);
xor U5065 (N_5065,N_4118,N_4320);
xnor U5066 (N_5066,N_4781,N_4589);
or U5067 (N_5067,N_4555,N_4012);
and U5068 (N_5068,N_4131,N_4121);
and U5069 (N_5069,N_4789,N_4571);
and U5070 (N_5070,N_4231,N_4077);
xnor U5071 (N_5071,N_4975,N_4863);
and U5072 (N_5072,N_4142,N_4899);
nor U5073 (N_5073,N_4946,N_4089);
nand U5074 (N_5074,N_4086,N_4604);
and U5075 (N_5075,N_4307,N_4473);
xor U5076 (N_5076,N_4111,N_4039);
nor U5077 (N_5077,N_4888,N_4002);
or U5078 (N_5078,N_4448,N_4215);
nor U5079 (N_5079,N_4308,N_4679);
xor U5080 (N_5080,N_4057,N_4859);
and U5081 (N_5081,N_4592,N_4819);
and U5082 (N_5082,N_4524,N_4218);
nor U5083 (N_5083,N_4745,N_4999);
or U5084 (N_5084,N_4858,N_4432);
nor U5085 (N_5085,N_4886,N_4561);
or U5086 (N_5086,N_4241,N_4136);
nand U5087 (N_5087,N_4714,N_4378);
and U5088 (N_5088,N_4598,N_4705);
and U5089 (N_5089,N_4274,N_4655);
nand U5090 (N_5090,N_4848,N_4005);
nand U5091 (N_5091,N_4201,N_4430);
or U5092 (N_5092,N_4491,N_4527);
nor U5093 (N_5093,N_4243,N_4935);
nor U5094 (N_5094,N_4816,N_4806);
and U5095 (N_5095,N_4855,N_4475);
xnor U5096 (N_5096,N_4618,N_4664);
nor U5097 (N_5097,N_4398,N_4785);
xnor U5098 (N_5098,N_4204,N_4088);
nand U5099 (N_5099,N_4949,N_4619);
nand U5100 (N_5100,N_4327,N_4446);
xor U5101 (N_5101,N_4465,N_4425);
and U5102 (N_5102,N_4026,N_4301);
nor U5103 (N_5103,N_4706,N_4911);
nor U5104 (N_5104,N_4860,N_4565);
nor U5105 (N_5105,N_4479,N_4893);
nor U5106 (N_5106,N_4586,N_4245);
nor U5107 (N_5107,N_4400,N_4867);
or U5108 (N_5108,N_4355,N_4185);
xnor U5109 (N_5109,N_4927,N_4252);
and U5110 (N_5110,N_4715,N_4658);
nand U5111 (N_5111,N_4915,N_4332);
xor U5112 (N_5112,N_4529,N_4251);
nor U5113 (N_5113,N_4288,N_4490);
nand U5114 (N_5114,N_4493,N_4442);
or U5115 (N_5115,N_4362,N_4059);
nor U5116 (N_5116,N_4771,N_4866);
nand U5117 (N_5117,N_4499,N_4075);
xnor U5118 (N_5118,N_4094,N_4849);
xor U5119 (N_5119,N_4551,N_4581);
nor U5120 (N_5120,N_4541,N_4438);
and U5121 (N_5121,N_4421,N_4595);
or U5122 (N_5122,N_4025,N_4263);
nor U5123 (N_5123,N_4722,N_4208);
or U5124 (N_5124,N_4410,N_4343);
and U5125 (N_5125,N_4196,N_4316);
and U5126 (N_5126,N_4138,N_4462);
xor U5127 (N_5127,N_4593,N_4125);
or U5128 (N_5128,N_4729,N_4763);
or U5129 (N_5129,N_4740,N_4702);
and U5130 (N_5130,N_4047,N_4104);
xnor U5131 (N_5131,N_4046,N_4407);
nand U5132 (N_5132,N_4804,N_4772);
xor U5133 (N_5133,N_4109,N_4956);
nand U5134 (N_5134,N_4548,N_4285);
nand U5135 (N_5135,N_4672,N_4787);
nor U5136 (N_5136,N_4240,N_4445);
nor U5137 (N_5137,N_4008,N_4021);
or U5138 (N_5138,N_4776,N_4471);
xnor U5139 (N_5139,N_4147,N_4158);
nor U5140 (N_5140,N_4289,N_4048);
and U5141 (N_5141,N_4885,N_4067);
xor U5142 (N_5142,N_4498,N_4965);
nor U5143 (N_5143,N_4038,N_4625);
or U5144 (N_5144,N_4071,N_4180);
xnor U5145 (N_5145,N_4698,N_4731);
or U5146 (N_5146,N_4451,N_4684);
nand U5147 (N_5147,N_4096,N_4010);
nand U5148 (N_5148,N_4594,N_4271);
nand U5149 (N_5149,N_4721,N_4757);
nor U5150 (N_5150,N_4405,N_4178);
xor U5151 (N_5151,N_4765,N_4478);
nand U5152 (N_5152,N_4359,N_4466);
or U5153 (N_5153,N_4526,N_4113);
xnor U5154 (N_5154,N_4384,N_4961);
xor U5155 (N_5155,N_4152,N_4967);
xor U5156 (N_5156,N_4457,N_4032);
nand U5157 (N_5157,N_4073,N_4114);
xor U5158 (N_5158,N_4105,N_4165);
or U5159 (N_5159,N_4756,N_4439);
and U5160 (N_5160,N_4264,N_4351);
nand U5161 (N_5161,N_4317,N_4216);
or U5162 (N_5162,N_4648,N_4651);
and U5163 (N_5163,N_4390,N_4022);
and U5164 (N_5164,N_4523,N_4993);
xor U5165 (N_5165,N_4719,N_4662);
xnor U5166 (N_5166,N_4634,N_4287);
xor U5167 (N_5167,N_4991,N_4857);
nor U5168 (N_5168,N_4794,N_4821);
xnor U5169 (N_5169,N_4381,N_4921);
xor U5170 (N_5170,N_4982,N_4040);
nor U5171 (N_5171,N_4902,N_4934);
nor U5172 (N_5172,N_4494,N_4574);
xor U5173 (N_5173,N_4331,N_4076);
nand U5174 (N_5174,N_4606,N_4875);
xnor U5175 (N_5175,N_4467,N_4019);
nor U5176 (N_5176,N_4006,N_4955);
nand U5177 (N_5177,N_4530,N_4512);
xor U5178 (N_5178,N_4936,N_4718);
nor U5179 (N_5179,N_4637,N_4657);
xor U5180 (N_5180,N_4203,N_4292);
and U5181 (N_5181,N_4509,N_4108);
and U5182 (N_5182,N_4418,N_4214);
or U5183 (N_5183,N_4909,N_4830);
and U5184 (N_5184,N_4923,N_4533);
and U5185 (N_5185,N_4353,N_4966);
nand U5186 (N_5186,N_4697,N_4575);
nor U5187 (N_5187,N_4741,N_4504);
xor U5188 (N_5188,N_4597,N_4962);
or U5189 (N_5189,N_4179,N_4358);
xor U5190 (N_5190,N_4227,N_4820);
xor U5191 (N_5191,N_4157,N_4199);
or U5192 (N_5192,N_4751,N_4474);
nand U5193 (N_5193,N_4519,N_4452);
nor U5194 (N_5194,N_4145,N_4782);
xor U5195 (N_5195,N_4470,N_4960);
xor U5196 (N_5196,N_4338,N_4995);
nand U5197 (N_5197,N_4141,N_4401);
xnor U5198 (N_5198,N_4416,N_4303);
or U5199 (N_5199,N_4389,N_4001);
xnor U5200 (N_5200,N_4337,N_4126);
nor U5201 (N_5201,N_4554,N_4450);
xor U5202 (N_5202,N_4024,N_4412);
nand U5203 (N_5203,N_4060,N_4708);
or U5204 (N_5204,N_4322,N_4209);
nor U5205 (N_5205,N_4954,N_4500);
and U5206 (N_5206,N_4318,N_4730);
nand U5207 (N_5207,N_4674,N_4248);
nor U5208 (N_5208,N_4815,N_4544);
or U5209 (N_5209,N_4424,N_4382);
xnor U5210 (N_5210,N_4319,N_4603);
nor U5211 (N_5211,N_4576,N_4894);
and U5212 (N_5212,N_4916,N_4366);
nor U5213 (N_5213,N_4834,N_4015);
and U5214 (N_5214,N_4069,N_4472);
and U5215 (N_5215,N_4054,N_4172);
or U5216 (N_5216,N_4117,N_4221);
nor U5217 (N_5217,N_4827,N_4100);
xor U5218 (N_5218,N_4345,N_4904);
or U5219 (N_5219,N_4877,N_4045);
and U5220 (N_5220,N_4266,N_4811);
nor U5221 (N_5221,N_4486,N_4079);
or U5222 (N_5222,N_4433,N_4626);
or U5223 (N_5223,N_4656,N_4053);
or U5224 (N_5224,N_4453,N_4406);
xor U5225 (N_5225,N_4990,N_4693);
nor U5226 (N_5226,N_4531,N_4206);
and U5227 (N_5227,N_4628,N_4572);
nor U5228 (N_5228,N_4070,N_4984);
or U5229 (N_5229,N_4154,N_4403);
or U5230 (N_5230,N_4455,N_4315);
nor U5231 (N_5231,N_4396,N_4978);
and U5232 (N_5232,N_4153,N_4485);
or U5233 (N_5233,N_4612,N_4423);
nand U5234 (N_5234,N_4583,N_4164);
and U5235 (N_5235,N_4163,N_4321);
and U5236 (N_5236,N_4035,N_4732);
or U5237 (N_5237,N_4766,N_4435);
nor U5238 (N_5238,N_4856,N_4895);
nand U5239 (N_5239,N_4103,N_4828);
and U5240 (N_5240,N_4232,N_4226);
or U5241 (N_5241,N_4686,N_4711);
nand U5242 (N_5242,N_4582,N_4809);
nor U5243 (N_5243,N_4036,N_4210);
or U5244 (N_5244,N_4461,N_4795);
or U5245 (N_5245,N_4380,N_4284);
xnor U5246 (N_5246,N_4712,N_4197);
nand U5247 (N_5247,N_4652,N_4633);
nand U5248 (N_5248,N_4511,N_4584);
or U5249 (N_5249,N_4552,N_4106);
or U5250 (N_5250,N_4842,N_4268);
nor U5251 (N_5251,N_4228,N_4023);
and U5252 (N_5252,N_4728,N_4269);
nor U5253 (N_5253,N_4041,N_4229);
and U5254 (N_5254,N_4341,N_4691);
nor U5255 (N_5255,N_4528,N_4309);
nor U5256 (N_5256,N_4115,N_4087);
or U5257 (N_5257,N_4399,N_4460);
xor U5258 (N_5258,N_4476,N_4862);
or U5259 (N_5259,N_4579,N_4174);
nor U5260 (N_5260,N_4761,N_4505);
nor U5261 (N_5261,N_4778,N_4083);
nor U5262 (N_5262,N_4558,N_4013);
and U5263 (N_5263,N_4814,N_4373);
and U5264 (N_5264,N_4437,N_4379);
or U5265 (N_5265,N_4037,N_4736);
nand U5266 (N_5266,N_4852,N_4890);
xnor U5267 (N_5267,N_4081,N_4621);
nand U5268 (N_5268,N_4235,N_4930);
nand U5269 (N_5269,N_4127,N_4906);
nand U5270 (N_5270,N_4896,N_4585);
xnor U5271 (N_5271,N_4831,N_4149);
and U5272 (N_5272,N_4979,N_4754);
nor U5273 (N_5273,N_4653,N_4539);
nor U5274 (N_5274,N_4496,N_4540);
xor U5275 (N_5275,N_4004,N_4974);
nor U5276 (N_5276,N_4912,N_4690);
xor U5277 (N_5277,N_4903,N_4800);
nand U5278 (N_5278,N_4347,N_4207);
and U5279 (N_5279,N_4791,N_4639);
nand U5280 (N_5280,N_4293,N_4596);
or U5281 (N_5281,N_4843,N_4361);
and U5282 (N_5282,N_4976,N_4826);
nor U5283 (N_5283,N_4159,N_4783);
nor U5284 (N_5284,N_4176,N_4668);
xor U5285 (N_5285,N_4660,N_4914);
nand U5286 (N_5286,N_4255,N_4411);
and U5287 (N_5287,N_4223,N_4063);
nand U5288 (N_5288,N_4644,N_4464);
nand U5289 (N_5289,N_4562,N_4357);
or U5290 (N_5290,N_4622,N_4901);
nand U5291 (N_5291,N_4868,N_4329);
or U5292 (N_5292,N_4680,N_4503);
nor U5293 (N_5293,N_4397,N_4259);
and U5294 (N_5294,N_4913,N_4426);
nand U5295 (N_5295,N_4051,N_4685);
xnor U5296 (N_5296,N_4310,N_4727);
and U5297 (N_5297,N_4260,N_4119);
or U5298 (N_5298,N_4845,N_4969);
nor U5299 (N_5299,N_4056,N_4265);
nand U5300 (N_5300,N_4281,N_4250);
and U5301 (N_5301,N_4769,N_4247);
nor U5302 (N_5302,N_4977,N_4107);
nor U5303 (N_5303,N_4542,N_4261);
xnor U5304 (N_5304,N_4171,N_4510);
nand U5305 (N_5305,N_4173,N_4892);
or U5306 (N_5306,N_4534,N_4973);
nand U5307 (N_5307,N_4546,N_4017);
nor U5308 (N_5308,N_4374,N_4792);
nand U5309 (N_5309,N_4093,N_4162);
nand U5310 (N_5310,N_4609,N_4387);
or U5311 (N_5311,N_4212,N_4198);
xor U5312 (N_5312,N_4872,N_4733);
or U5313 (N_5313,N_4532,N_4773);
xor U5314 (N_5314,N_4713,N_4553);
nand U5315 (N_5315,N_4099,N_4312);
nor U5316 (N_5316,N_4803,N_4988);
xnor U5317 (N_5317,N_4784,N_4755);
nor U5318 (N_5318,N_4588,N_4233);
nand U5319 (N_5319,N_4573,N_4280);
and U5320 (N_5320,N_4525,N_4360);
nor U5321 (N_5321,N_4924,N_4372);
nor U5322 (N_5322,N_4156,N_4066);
xor U5323 (N_5323,N_4839,N_4624);
nor U5324 (N_5324,N_4177,N_4919);
xnor U5325 (N_5325,N_4749,N_4671);
xor U5326 (N_5326,N_4029,N_4482);
xnor U5327 (N_5327,N_4072,N_4797);
xor U5328 (N_5328,N_4630,N_4502);
nand U5329 (N_5329,N_4182,N_4659);
nor U5330 (N_5330,N_4286,N_4760);
xnor U5331 (N_5331,N_4150,N_4349);
xnor U5332 (N_5332,N_4987,N_4447);
or U5333 (N_5333,N_4796,N_4964);
xor U5334 (N_5334,N_4011,N_4014);
nor U5335 (N_5335,N_4963,N_4774);
nand U5336 (N_5336,N_4567,N_4018);
and U5337 (N_5337,N_4234,N_4682);
and U5338 (N_5338,N_4033,N_4663);
or U5339 (N_5339,N_4441,N_4997);
and U5340 (N_5340,N_4333,N_4454);
xnor U5341 (N_5341,N_4770,N_4563);
and U5342 (N_5342,N_4880,N_4143);
or U5343 (N_5343,N_4189,N_4538);
and U5344 (N_5344,N_4807,N_4217);
xnor U5345 (N_5345,N_4940,N_4413);
and U5346 (N_5346,N_4495,N_4549);
nor U5347 (N_5347,N_4305,N_4402);
nor U5348 (N_5348,N_4869,N_4767);
or U5349 (N_5349,N_4151,N_4972);
or U5350 (N_5350,N_4238,N_4611);
or U5351 (N_5351,N_4780,N_4578);
and U5352 (N_5352,N_4091,N_4700);
xnor U5353 (N_5353,N_4677,N_4687);
xor U5354 (N_5354,N_4175,N_4296);
nand U5355 (N_5355,N_4556,N_4937);
nand U5356 (N_5356,N_4044,N_4220);
and U5357 (N_5357,N_4459,N_4422);
nor U5358 (N_5358,N_4701,N_4295);
nor U5359 (N_5359,N_4734,N_4339);
nor U5360 (N_5360,N_4090,N_4429);
nor U5361 (N_5361,N_4537,N_4920);
nor U5362 (N_5362,N_4181,N_4874);
xor U5363 (N_5363,N_4517,N_4031);
xnor U5364 (N_5364,N_4550,N_4282);
nand U5365 (N_5365,N_4810,N_4647);
nor U5366 (N_5366,N_4545,N_4992);
nand U5367 (N_5367,N_4098,N_4870);
or U5368 (N_5368,N_4068,N_4536);
nor U5369 (N_5369,N_4050,N_4654);
or U5370 (N_5370,N_4983,N_4354);
nor U5371 (N_5371,N_4580,N_4738);
nor U5372 (N_5372,N_4835,N_4417);
nand U5373 (N_5373,N_4393,N_4161);
or U5374 (N_5374,N_4294,N_4188);
or U5375 (N_5375,N_4489,N_4879);
or U5376 (N_5376,N_4887,N_4521);
or U5377 (N_5377,N_4786,N_4805);
nand U5378 (N_5378,N_4587,N_4950);
and U5379 (N_5379,N_4394,N_4184);
nor U5380 (N_5380,N_4385,N_4939);
nand U5381 (N_5381,N_4507,N_4420);
xor U5382 (N_5382,N_4336,N_4431);
or U5383 (N_5383,N_4646,N_4193);
xor U5384 (N_5384,N_4323,N_4833);
nor U5385 (N_5385,N_4237,N_4602);
nor U5386 (N_5386,N_4958,N_4951);
nor U5387 (N_5387,N_4645,N_4610);
and U5388 (N_5388,N_4673,N_4291);
and U5389 (N_5389,N_4824,N_4905);
and U5390 (N_5390,N_4386,N_4948);
and U5391 (N_5391,N_4167,N_4304);
or U5392 (N_5392,N_4515,N_4891);
and U5393 (N_5393,N_4752,N_4670);
nor U5394 (N_5394,N_4275,N_4825);
and U5395 (N_5395,N_4832,N_4166);
or U5396 (N_5396,N_4808,N_4742);
nor U5397 (N_5397,N_4847,N_4183);
xnor U5398 (N_5398,N_4615,N_4709);
or U5399 (N_5399,N_4623,N_4262);
nand U5400 (N_5400,N_4844,N_4364);
or U5401 (N_5401,N_4737,N_4169);
nor U5402 (N_5402,N_4346,N_4650);
or U5403 (N_5403,N_4929,N_4139);
xnor U5404 (N_5404,N_4302,N_4557);
nor U5405 (N_5405,N_4129,N_4120);
nand U5406 (N_5406,N_4219,N_4007);
nor U5407 (N_5407,N_4468,N_4084);
xnor U5408 (N_5408,N_4632,N_4027);
xnor U5409 (N_5409,N_4917,N_4812);
or U5410 (N_5410,N_4348,N_4409);
xnor U5411 (N_5411,N_4311,N_4080);
and U5412 (N_5412,N_4723,N_4484);
nand U5413 (N_5413,N_4871,N_4192);
nor U5414 (N_5414,N_4376,N_4959);
nand U5415 (N_5415,N_4375,N_4942);
nand U5416 (N_5416,N_4873,N_4635);
or U5417 (N_5417,N_4989,N_4876);
nor U5418 (N_5418,N_4501,N_4392);
or U5419 (N_5419,N_4764,N_4547);
nor U5420 (N_5420,N_4061,N_4617);
nand U5421 (N_5421,N_4908,N_4383);
xor U5422 (N_5422,N_4492,N_4638);
nor U5423 (N_5423,N_4676,N_4591);
xor U5424 (N_5424,N_4508,N_4123);
xor U5425 (N_5425,N_4799,N_4759);
nand U5426 (N_5426,N_4506,N_4922);
nor U5427 (N_5427,N_4724,N_4716);
nand U5428 (N_5428,N_4559,N_4725);
or U5429 (N_5429,N_4140,N_4613);
xor U5430 (N_5430,N_4112,N_4481);
nor U5431 (N_5431,N_4434,N_4324);
and U5432 (N_5432,N_4981,N_4202);
or U5433 (N_5433,N_4590,N_4941);
nor U5434 (N_5434,N_4980,N_4273);
nor U5435 (N_5435,N_4750,N_4878);
or U5436 (N_5436,N_4062,N_4513);
xor U5437 (N_5437,N_4971,N_4699);
and U5438 (N_5438,N_4244,N_4191);
xor U5439 (N_5439,N_4846,N_4225);
or U5440 (N_5440,N_4683,N_4444);
xor U5441 (N_5441,N_4775,N_4943);
or U5442 (N_5442,N_4522,N_4535);
and U5443 (N_5443,N_4427,N_4838);
xor U5444 (N_5444,N_4313,N_4279);
nor U5445 (N_5445,N_4395,N_4897);
nand U5446 (N_5446,N_4095,N_4793);
xor U5447 (N_5447,N_4283,N_4854);
nor U5448 (N_5448,N_4695,N_4998);
or U5449 (N_5449,N_4325,N_4116);
nand U5450 (N_5450,N_4837,N_4823);
nor U5451 (N_5451,N_4132,N_4469);
xor U5452 (N_5452,N_4110,N_4130);
nand U5453 (N_5453,N_4520,N_4881);
or U5454 (N_5454,N_4851,N_4600);
and U5455 (N_5455,N_4813,N_4160);
or U5456 (N_5456,N_4928,N_4643);
or U5457 (N_5457,N_4568,N_4641);
nand U5458 (N_5458,N_4601,N_4788);
or U5459 (N_5459,N_4661,N_4440);
or U5460 (N_5460,N_4744,N_4367);
nor U5461 (N_5461,N_4629,N_4122);
nand U5462 (N_5462,N_4415,N_4514);
xnor U5463 (N_5463,N_4817,N_4326);
or U5464 (N_5464,N_4841,N_4931);
nand U5465 (N_5465,N_4570,N_4135);
nor U5466 (N_5466,N_4428,N_4566);
nor U5467 (N_5467,N_4840,N_4861);
and U5468 (N_5468,N_4994,N_4055);
nand U5469 (N_5469,N_4704,N_4144);
nor U5470 (N_5470,N_4497,N_4449);
nor U5471 (N_5471,N_4688,N_4918);
or U5472 (N_5472,N_4932,N_4085);
nor U5473 (N_5473,N_4836,N_4404);
xor U5474 (N_5474,N_4743,N_4669);
nand U5475 (N_5475,N_4043,N_4577);
and U5476 (N_5476,N_4480,N_4101);
nand U5477 (N_5477,N_4726,N_4065);
nor U5478 (N_5478,N_4200,N_4306);
or U5479 (N_5479,N_4614,N_4249);
nand U5480 (N_5480,N_4369,N_4518);
and U5481 (N_5481,N_4335,N_4340);
and U5482 (N_5482,N_4483,N_4666);
nand U5483 (N_5483,N_4944,N_4477);
or U5484 (N_5484,N_4898,N_4640);
and U5485 (N_5485,N_4543,N_4758);
or U5486 (N_5486,N_4186,N_4419);
or U5487 (N_5487,N_4242,N_4236);
nand U5488 (N_5488,N_4720,N_4925);
xor U5489 (N_5489,N_4391,N_4636);
xor U5490 (N_5490,N_4224,N_4762);
and U5491 (N_5491,N_4246,N_4938);
and U5492 (N_5492,N_4620,N_4290);
nor U5493 (N_5493,N_4102,N_4064);
xor U5494 (N_5494,N_4049,N_4256);
and U5495 (N_5495,N_4414,N_4170);
nor U5496 (N_5496,N_4253,N_4133);
and U5497 (N_5497,N_4889,N_4230);
or U5498 (N_5498,N_4488,N_4802);
nor U5499 (N_5499,N_4822,N_4945);
and U5500 (N_5500,N_4565,N_4731);
and U5501 (N_5501,N_4822,N_4400);
xor U5502 (N_5502,N_4995,N_4580);
nand U5503 (N_5503,N_4011,N_4746);
or U5504 (N_5504,N_4896,N_4377);
xor U5505 (N_5505,N_4651,N_4513);
and U5506 (N_5506,N_4855,N_4503);
nor U5507 (N_5507,N_4067,N_4056);
xor U5508 (N_5508,N_4187,N_4707);
or U5509 (N_5509,N_4947,N_4562);
and U5510 (N_5510,N_4466,N_4997);
nand U5511 (N_5511,N_4103,N_4042);
xnor U5512 (N_5512,N_4997,N_4564);
or U5513 (N_5513,N_4220,N_4066);
and U5514 (N_5514,N_4129,N_4414);
nor U5515 (N_5515,N_4962,N_4954);
and U5516 (N_5516,N_4418,N_4772);
nand U5517 (N_5517,N_4499,N_4399);
xor U5518 (N_5518,N_4069,N_4823);
or U5519 (N_5519,N_4135,N_4281);
or U5520 (N_5520,N_4099,N_4143);
nor U5521 (N_5521,N_4879,N_4600);
nand U5522 (N_5522,N_4590,N_4400);
and U5523 (N_5523,N_4853,N_4321);
xor U5524 (N_5524,N_4972,N_4748);
xor U5525 (N_5525,N_4930,N_4366);
nand U5526 (N_5526,N_4971,N_4347);
nor U5527 (N_5527,N_4967,N_4787);
nand U5528 (N_5528,N_4021,N_4539);
and U5529 (N_5529,N_4177,N_4860);
xor U5530 (N_5530,N_4562,N_4557);
nand U5531 (N_5531,N_4597,N_4633);
nand U5532 (N_5532,N_4157,N_4540);
or U5533 (N_5533,N_4145,N_4550);
and U5534 (N_5534,N_4134,N_4425);
and U5535 (N_5535,N_4108,N_4125);
or U5536 (N_5536,N_4054,N_4524);
and U5537 (N_5537,N_4147,N_4374);
nor U5538 (N_5538,N_4061,N_4024);
nor U5539 (N_5539,N_4547,N_4573);
or U5540 (N_5540,N_4681,N_4618);
or U5541 (N_5541,N_4271,N_4925);
or U5542 (N_5542,N_4937,N_4545);
and U5543 (N_5543,N_4930,N_4863);
nor U5544 (N_5544,N_4781,N_4012);
and U5545 (N_5545,N_4989,N_4601);
and U5546 (N_5546,N_4082,N_4675);
nor U5547 (N_5547,N_4670,N_4346);
or U5548 (N_5548,N_4076,N_4812);
or U5549 (N_5549,N_4231,N_4100);
or U5550 (N_5550,N_4026,N_4086);
nand U5551 (N_5551,N_4942,N_4115);
and U5552 (N_5552,N_4060,N_4835);
nor U5553 (N_5553,N_4965,N_4102);
nor U5554 (N_5554,N_4030,N_4409);
and U5555 (N_5555,N_4916,N_4199);
nor U5556 (N_5556,N_4529,N_4631);
xnor U5557 (N_5557,N_4594,N_4258);
nand U5558 (N_5558,N_4823,N_4575);
or U5559 (N_5559,N_4749,N_4336);
nor U5560 (N_5560,N_4523,N_4888);
xor U5561 (N_5561,N_4019,N_4624);
xor U5562 (N_5562,N_4262,N_4986);
xnor U5563 (N_5563,N_4168,N_4847);
nand U5564 (N_5564,N_4542,N_4320);
nor U5565 (N_5565,N_4613,N_4163);
nor U5566 (N_5566,N_4901,N_4018);
nor U5567 (N_5567,N_4220,N_4646);
xnor U5568 (N_5568,N_4274,N_4716);
and U5569 (N_5569,N_4868,N_4982);
and U5570 (N_5570,N_4710,N_4059);
or U5571 (N_5571,N_4918,N_4566);
or U5572 (N_5572,N_4755,N_4815);
nand U5573 (N_5573,N_4708,N_4795);
nor U5574 (N_5574,N_4931,N_4978);
nor U5575 (N_5575,N_4560,N_4141);
and U5576 (N_5576,N_4277,N_4236);
nor U5577 (N_5577,N_4227,N_4074);
and U5578 (N_5578,N_4423,N_4425);
or U5579 (N_5579,N_4600,N_4745);
nand U5580 (N_5580,N_4935,N_4582);
or U5581 (N_5581,N_4809,N_4850);
nor U5582 (N_5582,N_4981,N_4910);
nor U5583 (N_5583,N_4394,N_4964);
and U5584 (N_5584,N_4625,N_4670);
and U5585 (N_5585,N_4617,N_4442);
nand U5586 (N_5586,N_4663,N_4163);
or U5587 (N_5587,N_4745,N_4545);
or U5588 (N_5588,N_4883,N_4728);
or U5589 (N_5589,N_4888,N_4471);
or U5590 (N_5590,N_4531,N_4333);
xnor U5591 (N_5591,N_4145,N_4279);
and U5592 (N_5592,N_4988,N_4309);
xor U5593 (N_5593,N_4077,N_4254);
nor U5594 (N_5594,N_4746,N_4409);
xnor U5595 (N_5595,N_4912,N_4589);
xor U5596 (N_5596,N_4596,N_4466);
xnor U5597 (N_5597,N_4234,N_4629);
or U5598 (N_5598,N_4514,N_4134);
xnor U5599 (N_5599,N_4735,N_4469);
nand U5600 (N_5600,N_4837,N_4347);
nor U5601 (N_5601,N_4961,N_4940);
xnor U5602 (N_5602,N_4441,N_4748);
nand U5603 (N_5603,N_4144,N_4213);
nor U5604 (N_5604,N_4712,N_4299);
nor U5605 (N_5605,N_4917,N_4701);
or U5606 (N_5606,N_4711,N_4505);
nand U5607 (N_5607,N_4688,N_4641);
nor U5608 (N_5608,N_4263,N_4660);
xor U5609 (N_5609,N_4265,N_4257);
xnor U5610 (N_5610,N_4308,N_4373);
or U5611 (N_5611,N_4788,N_4113);
or U5612 (N_5612,N_4276,N_4374);
and U5613 (N_5613,N_4609,N_4856);
nand U5614 (N_5614,N_4903,N_4223);
nor U5615 (N_5615,N_4292,N_4719);
and U5616 (N_5616,N_4729,N_4565);
nor U5617 (N_5617,N_4590,N_4104);
nor U5618 (N_5618,N_4269,N_4025);
or U5619 (N_5619,N_4819,N_4611);
and U5620 (N_5620,N_4363,N_4859);
xor U5621 (N_5621,N_4458,N_4981);
and U5622 (N_5622,N_4693,N_4875);
xor U5623 (N_5623,N_4830,N_4393);
or U5624 (N_5624,N_4630,N_4202);
nand U5625 (N_5625,N_4662,N_4273);
xnor U5626 (N_5626,N_4560,N_4452);
and U5627 (N_5627,N_4360,N_4984);
and U5628 (N_5628,N_4574,N_4493);
or U5629 (N_5629,N_4950,N_4797);
xor U5630 (N_5630,N_4755,N_4645);
xnor U5631 (N_5631,N_4923,N_4244);
nand U5632 (N_5632,N_4458,N_4684);
xor U5633 (N_5633,N_4533,N_4643);
nand U5634 (N_5634,N_4696,N_4217);
xor U5635 (N_5635,N_4027,N_4480);
xnor U5636 (N_5636,N_4171,N_4308);
xor U5637 (N_5637,N_4367,N_4560);
or U5638 (N_5638,N_4533,N_4502);
nor U5639 (N_5639,N_4222,N_4594);
and U5640 (N_5640,N_4773,N_4321);
xnor U5641 (N_5641,N_4456,N_4552);
xor U5642 (N_5642,N_4383,N_4145);
xor U5643 (N_5643,N_4758,N_4609);
or U5644 (N_5644,N_4040,N_4776);
nor U5645 (N_5645,N_4883,N_4081);
and U5646 (N_5646,N_4085,N_4450);
or U5647 (N_5647,N_4332,N_4079);
xnor U5648 (N_5648,N_4721,N_4057);
and U5649 (N_5649,N_4753,N_4875);
nor U5650 (N_5650,N_4056,N_4661);
and U5651 (N_5651,N_4218,N_4076);
nand U5652 (N_5652,N_4308,N_4183);
or U5653 (N_5653,N_4707,N_4492);
nand U5654 (N_5654,N_4050,N_4916);
and U5655 (N_5655,N_4865,N_4787);
nand U5656 (N_5656,N_4725,N_4798);
nor U5657 (N_5657,N_4899,N_4190);
xor U5658 (N_5658,N_4848,N_4011);
and U5659 (N_5659,N_4914,N_4099);
or U5660 (N_5660,N_4515,N_4460);
and U5661 (N_5661,N_4302,N_4153);
or U5662 (N_5662,N_4811,N_4351);
nand U5663 (N_5663,N_4417,N_4178);
xnor U5664 (N_5664,N_4993,N_4642);
and U5665 (N_5665,N_4829,N_4152);
nor U5666 (N_5666,N_4709,N_4935);
or U5667 (N_5667,N_4284,N_4538);
nor U5668 (N_5668,N_4873,N_4703);
and U5669 (N_5669,N_4407,N_4691);
xor U5670 (N_5670,N_4431,N_4737);
nor U5671 (N_5671,N_4830,N_4305);
nand U5672 (N_5672,N_4736,N_4739);
xor U5673 (N_5673,N_4298,N_4162);
nand U5674 (N_5674,N_4024,N_4467);
and U5675 (N_5675,N_4603,N_4394);
nand U5676 (N_5676,N_4125,N_4491);
nor U5677 (N_5677,N_4423,N_4979);
and U5678 (N_5678,N_4931,N_4057);
nor U5679 (N_5679,N_4260,N_4564);
and U5680 (N_5680,N_4450,N_4305);
xor U5681 (N_5681,N_4919,N_4861);
xnor U5682 (N_5682,N_4406,N_4412);
nand U5683 (N_5683,N_4272,N_4065);
nand U5684 (N_5684,N_4700,N_4861);
nor U5685 (N_5685,N_4651,N_4094);
or U5686 (N_5686,N_4162,N_4064);
xnor U5687 (N_5687,N_4140,N_4300);
nor U5688 (N_5688,N_4177,N_4695);
xnor U5689 (N_5689,N_4679,N_4798);
and U5690 (N_5690,N_4736,N_4777);
xor U5691 (N_5691,N_4112,N_4746);
nor U5692 (N_5692,N_4429,N_4156);
xnor U5693 (N_5693,N_4984,N_4875);
nor U5694 (N_5694,N_4727,N_4006);
or U5695 (N_5695,N_4394,N_4498);
and U5696 (N_5696,N_4497,N_4213);
xor U5697 (N_5697,N_4534,N_4037);
nand U5698 (N_5698,N_4080,N_4376);
or U5699 (N_5699,N_4979,N_4536);
xnor U5700 (N_5700,N_4710,N_4493);
and U5701 (N_5701,N_4746,N_4962);
or U5702 (N_5702,N_4490,N_4954);
nand U5703 (N_5703,N_4732,N_4936);
nand U5704 (N_5704,N_4181,N_4638);
or U5705 (N_5705,N_4750,N_4830);
and U5706 (N_5706,N_4064,N_4935);
or U5707 (N_5707,N_4833,N_4953);
xor U5708 (N_5708,N_4098,N_4071);
and U5709 (N_5709,N_4620,N_4726);
and U5710 (N_5710,N_4984,N_4503);
and U5711 (N_5711,N_4964,N_4921);
xnor U5712 (N_5712,N_4894,N_4621);
nor U5713 (N_5713,N_4448,N_4919);
nor U5714 (N_5714,N_4405,N_4105);
nor U5715 (N_5715,N_4777,N_4307);
xor U5716 (N_5716,N_4474,N_4033);
nor U5717 (N_5717,N_4274,N_4583);
nand U5718 (N_5718,N_4756,N_4648);
nand U5719 (N_5719,N_4145,N_4275);
or U5720 (N_5720,N_4592,N_4467);
xor U5721 (N_5721,N_4949,N_4966);
nand U5722 (N_5722,N_4555,N_4273);
and U5723 (N_5723,N_4339,N_4030);
nand U5724 (N_5724,N_4463,N_4090);
nand U5725 (N_5725,N_4200,N_4375);
nand U5726 (N_5726,N_4303,N_4968);
and U5727 (N_5727,N_4519,N_4896);
nor U5728 (N_5728,N_4010,N_4637);
xnor U5729 (N_5729,N_4013,N_4347);
nor U5730 (N_5730,N_4038,N_4258);
or U5731 (N_5731,N_4813,N_4540);
and U5732 (N_5732,N_4337,N_4678);
nor U5733 (N_5733,N_4781,N_4351);
and U5734 (N_5734,N_4686,N_4308);
nor U5735 (N_5735,N_4911,N_4821);
or U5736 (N_5736,N_4014,N_4518);
xor U5737 (N_5737,N_4417,N_4908);
nand U5738 (N_5738,N_4506,N_4159);
nand U5739 (N_5739,N_4649,N_4280);
or U5740 (N_5740,N_4293,N_4484);
and U5741 (N_5741,N_4104,N_4602);
nor U5742 (N_5742,N_4911,N_4754);
or U5743 (N_5743,N_4128,N_4604);
and U5744 (N_5744,N_4743,N_4977);
nor U5745 (N_5745,N_4468,N_4933);
nor U5746 (N_5746,N_4183,N_4495);
nand U5747 (N_5747,N_4181,N_4500);
or U5748 (N_5748,N_4784,N_4201);
xor U5749 (N_5749,N_4319,N_4062);
or U5750 (N_5750,N_4414,N_4734);
and U5751 (N_5751,N_4953,N_4272);
nand U5752 (N_5752,N_4908,N_4891);
or U5753 (N_5753,N_4221,N_4368);
and U5754 (N_5754,N_4584,N_4242);
and U5755 (N_5755,N_4577,N_4222);
nand U5756 (N_5756,N_4404,N_4620);
and U5757 (N_5757,N_4296,N_4793);
and U5758 (N_5758,N_4034,N_4664);
and U5759 (N_5759,N_4784,N_4068);
xnor U5760 (N_5760,N_4559,N_4999);
nor U5761 (N_5761,N_4704,N_4693);
nor U5762 (N_5762,N_4933,N_4866);
nor U5763 (N_5763,N_4990,N_4405);
nand U5764 (N_5764,N_4872,N_4932);
nand U5765 (N_5765,N_4892,N_4290);
or U5766 (N_5766,N_4575,N_4098);
nand U5767 (N_5767,N_4044,N_4532);
and U5768 (N_5768,N_4737,N_4141);
and U5769 (N_5769,N_4404,N_4313);
xor U5770 (N_5770,N_4688,N_4197);
xnor U5771 (N_5771,N_4343,N_4980);
and U5772 (N_5772,N_4977,N_4693);
nand U5773 (N_5773,N_4677,N_4905);
xor U5774 (N_5774,N_4464,N_4899);
xor U5775 (N_5775,N_4995,N_4541);
nand U5776 (N_5776,N_4727,N_4092);
xor U5777 (N_5777,N_4465,N_4131);
and U5778 (N_5778,N_4043,N_4139);
nand U5779 (N_5779,N_4310,N_4151);
xor U5780 (N_5780,N_4678,N_4861);
nand U5781 (N_5781,N_4969,N_4426);
or U5782 (N_5782,N_4770,N_4519);
nand U5783 (N_5783,N_4968,N_4708);
nor U5784 (N_5784,N_4648,N_4044);
or U5785 (N_5785,N_4435,N_4448);
nor U5786 (N_5786,N_4932,N_4742);
xor U5787 (N_5787,N_4936,N_4282);
xnor U5788 (N_5788,N_4093,N_4030);
xor U5789 (N_5789,N_4297,N_4026);
xor U5790 (N_5790,N_4031,N_4683);
xnor U5791 (N_5791,N_4075,N_4071);
and U5792 (N_5792,N_4893,N_4175);
and U5793 (N_5793,N_4568,N_4827);
nor U5794 (N_5794,N_4326,N_4168);
xor U5795 (N_5795,N_4400,N_4791);
or U5796 (N_5796,N_4329,N_4192);
or U5797 (N_5797,N_4589,N_4128);
or U5798 (N_5798,N_4823,N_4410);
nand U5799 (N_5799,N_4405,N_4311);
xnor U5800 (N_5800,N_4682,N_4363);
or U5801 (N_5801,N_4592,N_4230);
and U5802 (N_5802,N_4119,N_4933);
nor U5803 (N_5803,N_4514,N_4964);
or U5804 (N_5804,N_4337,N_4052);
or U5805 (N_5805,N_4716,N_4072);
nor U5806 (N_5806,N_4496,N_4382);
and U5807 (N_5807,N_4108,N_4433);
nand U5808 (N_5808,N_4936,N_4211);
nand U5809 (N_5809,N_4036,N_4227);
nand U5810 (N_5810,N_4435,N_4242);
or U5811 (N_5811,N_4584,N_4889);
xnor U5812 (N_5812,N_4422,N_4237);
xnor U5813 (N_5813,N_4725,N_4466);
nor U5814 (N_5814,N_4943,N_4994);
and U5815 (N_5815,N_4618,N_4892);
or U5816 (N_5816,N_4834,N_4872);
and U5817 (N_5817,N_4848,N_4792);
nor U5818 (N_5818,N_4121,N_4125);
xor U5819 (N_5819,N_4761,N_4815);
or U5820 (N_5820,N_4953,N_4486);
nand U5821 (N_5821,N_4811,N_4114);
and U5822 (N_5822,N_4727,N_4251);
and U5823 (N_5823,N_4002,N_4465);
xnor U5824 (N_5824,N_4415,N_4245);
xor U5825 (N_5825,N_4283,N_4007);
xor U5826 (N_5826,N_4129,N_4043);
xor U5827 (N_5827,N_4269,N_4848);
and U5828 (N_5828,N_4011,N_4326);
nand U5829 (N_5829,N_4502,N_4074);
or U5830 (N_5830,N_4983,N_4932);
nand U5831 (N_5831,N_4474,N_4973);
or U5832 (N_5832,N_4766,N_4673);
xor U5833 (N_5833,N_4697,N_4052);
and U5834 (N_5834,N_4242,N_4915);
nor U5835 (N_5835,N_4957,N_4215);
nor U5836 (N_5836,N_4323,N_4418);
nand U5837 (N_5837,N_4131,N_4593);
nor U5838 (N_5838,N_4469,N_4864);
nand U5839 (N_5839,N_4480,N_4831);
nand U5840 (N_5840,N_4283,N_4835);
nor U5841 (N_5841,N_4502,N_4324);
nand U5842 (N_5842,N_4166,N_4519);
nor U5843 (N_5843,N_4423,N_4743);
and U5844 (N_5844,N_4729,N_4890);
nor U5845 (N_5845,N_4088,N_4550);
and U5846 (N_5846,N_4327,N_4630);
nor U5847 (N_5847,N_4701,N_4993);
nand U5848 (N_5848,N_4611,N_4410);
nand U5849 (N_5849,N_4152,N_4343);
xnor U5850 (N_5850,N_4632,N_4035);
or U5851 (N_5851,N_4993,N_4650);
or U5852 (N_5852,N_4372,N_4144);
nand U5853 (N_5853,N_4041,N_4154);
xor U5854 (N_5854,N_4840,N_4558);
or U5855 (N_5855,N_4833,N_4094);
nor U5856 (N_5856,N_4946,N_4657);
xnor U5857 (N_5857,N_4834,N_4478);
nor U5858 (N_5858,N_4723,N_4860);
and U5859 (N_5859,N_4914,N_4782);
nor U5860 (N_5860,N_4773,N_4406);
nand U5861 (N_5861,N_4480,N_4596);
xnor U5862 (N_5862,N_4385,N_4330);
nor U5863 (N_5863,N_4391,N_4733);
nor U5864 (N_5864,N_4276,N_4229);
and U5865 (N_5865,N_4728,N_4971);
or U5866 (N_5866,N_4753,N_4829);
xnor U5867 (N_5867,N_4130,N_4596);
and U5868 (N_5868,N_4240,N_4702);
or U5869 (N_5869,N_4395,N_4108);
nor U5870 (N_5870,N_4863,N_4431);
nand U5871 (N_5871,N_4914,N_4104);
or U5872 (N_5872,N_4687,N_4601);
nor U5873 (N_5873,N_4788,N_4581);
nor U5874 (N_5874,N_4591,N_4625);
xnor U5875 (N_5875,N_4492,N_4252);
or U5876 (N_5876,N_4682,N_4357);
nand U5877 (N_5877,N_4873,N_4821);
nand U5878 (N_5878,N_4114,N_4334);
or U5879 (N_5879,N_4466,N_4935);
nor U5880 (N_5880,N_4611,N_4961);
or U5881 (N_5881,N_4808,N_4010);
nor U5882 (N_5882,N_4577,N_4400);
and U5883 (N_5883,N_4423,N_4868);
nand U5884 (N_5884,N_4705,N_4446);
nor U5885 (N_5885,N_4946,N_4486);
and U5886 (N_5886,N_4307,N_4355);
and U5887 (N_5887,N_4091,N_4409);
or U5888 (N_5888,N_4291,N_4415);
or U5889 (N_5889,N_4453,N_4546);
xnor U5890 (N_5890,N_4879,N_4093);
or U5891 (N_5891,N_4042,N_4668);
nand U5892 (N_5892,N_4582,N_4599);
or U5893 (N_5893,N_4977,N_4850);
or U5894 (N_5894,N_4907,N_4946);
and U5895 (N_5895,N_4093,N_4863);
and U5896 (N_5896,N_4636,N_4399);
or U5897 (N_5897,N_4710,N_4480);
and U5898 (N_5898,N_4461,N_4241);
nand U5899 (N_5899,N_4150,N_4013);
nor U5900 (N_5900,N_4267,N_4826);
nor U5901 (N_5901,N_4504,N_4061);
xnor U5902 (N_5902,N_4158,N_4772);
xor U5903 (N_5903,N_4756,N_4496);
nand U5904 (N_5904,N_4978,N_4715);
nor U5905 (N_5905,N_4806,N_4486);
nand U5906 (N_5906,N_4552,N_4976);
or U5907 (N_5907,N_4334,N_4049);
or U5908 (N_5908,N_4822,N_4251);
xnor U5909 (N_5909,N_4591,N_4353);
or U5910 (N_5910,N_4712,N_4051);
xnor U5911 (N_5911,N_4766,N_4247);
xor U5912 (N_5912,N_4548,N_4675);
or U5913 (N_5913,N_4355,N_4592);
nand U5914 (N_5914,N_4389,N_4611);
and U5915 (N_5915,N_4674,N_4258);
or U5916 (N_5916,N_4961,N_4771);
and U5917 (N_5917,N_4944,N_4563);
or U5918 (N_5918,N_4999,N_4752);
or U5919 (N_5919,N_4788,N_4115);
xnor U5920 (N_5920,N_4161,N_4322);
nand U5921 (N_5921,N_4109,N_4254);
xor U5922 (N_5922,N_4781,N_4971);
xor U5923 (N_5923,N_4977,N_4520);
nand U5924 (N_5924,N_4521,N_4419);
and U5925 (N_5925,N_4355,N_4629);
or U5926 (N_5926,N_4245,N_4532);
and U5927 (N_5927,N_4152,N_4555);
nor U5928 (N_5928,N_4195,N_4557);
and U5929 (N_5929,N_4209,N_4749);
nand U5930 (N_5930,N_4559,N_4569);
nor U5931 (N_5931,N_4560,N_4756);
or U5932 (N_5932,N_4193,N_4253);
or U5933 (N_5933,N_4033,N_4378);
nor U5934 (N_5934,N_4043,N_4599);
nand U5935 (N_5935,N_4665,N_4141);
nand U5936 (N_5936,N_4013,N_4384);
nand U5937 (N_5937,N_4876,N_4146);
xor U5938 (N_5938,N_4446,N_4295);
and U5939 (N_5939,N_4600,N_4639);
and U5940 (N_5940,N_4136,N_4592);
nor U5941 (N_5941,N_4807,N_4134);
and U5942 (N_5942,N_4269,N_4927);
and U5943 (N_5943,N_4954,N_4138);
nor U5944 (N_5944,N_4380,N_4099);
xor U5945 (N_5945,N_4332,N_4580);
nand U5946 (N_5946,N_4947,N_4365);
or U5947 (N_5947,N_4134,N_4364);
nand U5948 (N_5948,N_4237,N_4014);
nor U5949 (N_5949,N_4282,N_4442);
nor U5950 (N_5950,N_4441,N_4599);
nor U5951 (N_5951,N_4470,N_4527);
nor U5952 (N_5952,N_4084,N_4092);
nor U5953 (N_5953,N_4827,N_4025);
nand U5954 (N_5954,N_4203,N_4533);
nor U5955 (N_5955,N_4676,N_4374);
nand U5956 (N_5956,N_4540,N_4762);
and U5957 (N_5957,N_4489,N_4917);
or U5958 (N_5958,N_4462,N_4168);
or U5959 (N_5959,N_4183,N_4676);
nand U5960 (N_5960,N_4340,N_4974);
nor U5961 (N_5961,N_4466,N_4900);
and U5962 (N_5962,N_4471,N_4793);
nor U5963 (N_5963,N_4187,N_4720);
and U5964 (N_5964,N_4260,N_4659);
nor U5965 (N_5965,N_4833,N_4907);
xor U5966 (N_5966,N_4232,N_4973);
nor U5967 (N_5967,N_4256,N_4705);
xor U5968 (N_5968,N_4168,N_4425);
nand U5969 (N_5969,N_4541,N_4088);
nor U5970 (N_5970,N_4664,N_4011);
or U5971 (N_5971,N_4410,N_4318);
and U5972 (N_5972,N_4836,N_4165);
xnor U5973 (N_5973,N_4475,N_4629);
xnor U5974 (N_5974,N_4695,N_4437);
nand U5975 (N_5975,N_4719,N_4269);
nand U5976 (N_5976,N_4166,N_4480);
nor U5977 (N_5977,N_4457,N_4776);
or U5978 (N_5978,N_4784,N_4132);
and U5979 (N_5979,N_4494,N_4784);
nand U5980 (N_5980,N_4794,N_4085);
nand U5981 (N_5981,N_4535,N_4776);
and U5982 (N_5982,N_4023,N_4854);
xnor U5983 (N_5983,N_4319,N_4584);
nor U5984 (N_5984,N_4776,N_4665);
or U5985 (N_5985,N_4011,N_4876);
nor U5986 (N_5986,N_4961,N_4496);
nand U5987 (N_5987,N_4199,N_4060);
and U5988 (N_5988,N_4999,N_4594);
nor U5989 (N_5989,N_4466,N_4213);
nor U5990 (N_5990,N_4754,N_4958);
nand U5991 (N_5991,N_4877,N_4821);
nor U5992 (N_5992,N_4798,N_4092);
and U5993 (N_5993,N_4547,N_4761);
nor U5994 (N_5994,N_4181,N_4084);
xor U5995 (N_5995,N_4690,N_4610);
nand U5996 (N_5996,N_4679,N_4231);
nor U5997 (N_5997,N_4255,N_4642);
and U5998 (N_5998,N_4328,N_4858);
nand U5999 (N_5999,N_4761,N_4877);
or U6000 (N_6000,N_5025,N_5213);
and U6001 (N_6001,N_5968,N_5194);
and U6002 (N_6002,N_5529,N_5693);
nand U6003 (N_6003,N_5954,N_5270);
nor U6004 (N_6004,N_5915,N_5625);
nor U6005 (N_6005,N_5227,N_5958);
or U6006 (N_6006,N_5516,N_5598);
xnor U6007 (N_6007,N_5171,N_5990);
xor U6008 (N_6008,N_5081,N_5276);
nor U6009 (N_6009,N_5736,N_5433);
nor U6010 (N_6010,N_5146,N_5112);
xor U6011 (N_6011,N_5997,N_5315);
xnor U6012 (N_6012,N_5196,N_5104);
and U6013 (N_6013,N_5463,N_5048);
nand U6014 (N_6014,N_5881,N_5240);
and U6015 (N_6015,N_5897,N_5019);
or U6016 (N_6016,N_5861,N_5153);
nand U6017 (N_6017,N_5623,N_5280);
and U6018 (N_6018,N_5775,N_5924);
nor U6019 (N_6019,N_5036,N_5945);
nand U6020 (N_6020,N_5841,N_5498);
or U6021 (N_6021,N_5798,N_5829);
nor U6022 (N_6022,N_5416,N_5307);
nand U6023 (N_6023,N_5940,N_5778);
xor U6024 (N_6024,N_5965,N_5192);
nor U6025 (N_6025,N_5344,N_5957);
nand U6026 (N_6026,N_5197,N_5089);
and U6027 (N_6027,N_5577,N_5052);
or U6028 (N_6028,N_5278,N_5855);
nor U6029 (N_6029,N_5319,N_5637);
nand U6030 (N_6030,N_5900,N_5215);
nand U6031 (N_6031,N_5604,N_5730);
and U6032 (N_6032,N_5642,N_5528);
and U6033 (N_6033,N_5804,N_5523);
xor U6034 (N_6034,N_5888,N_5842);
and U6035 (N_6035,N_5147,N_5876);
and U6036 (N_6036,N_5088,N_5993);
nor U6037 (N_6037,N_5282,N_5752);
or U6038 (N_6038,N_5672,N_5445);
nor U6039 (N_6039,N_5012,N_5426);
xor U6040 (N_6040,N_5667,N_5558);
or U6041 (N_6041,N_5039,N_5718);
nor U6042 (N_6042,N_5294,N_5066);
and U6043 (N_6043,N_5184,N_5468);
nor U6044 (N_6044,N_5093,N_5480);
nor U6045 (N_6045,N_5476,N_5305);
nand U6046 (N_6046,N_5053,N_5844);
and U6047 (N_6047,N_5273,N_5700);
xor U6048 (N_6048,N_5148,N_5072);
or U6049 (N_6049,N_5701,N_5359);
or U6050 (N_6050,N_5601,N_5919);
nand U6051 (N_6051,N_5521,N_5921);
or U6052 (N_6052,N_5596,N_5208);
nand U6053 (N_6053,N_5210,N_5483);
nand U6054 (N_6054,N_5682,N_5152);
nand U6055 (N_6055,N_5602,N_5226);
nand U6056 (N_6056,N_5974,N_5744);
and U6057 (N_6057,N_5246,N_5203);
xor U6058 (N_6058,N_5544,N_5615);
and U6059 (N_6059,N_5982,N_5326);
and U6060 (N_6060,N_5320,N_5794);
and U6061 (N_6061,N_5253,N_5686);
nor U6062 (N_6062,N_5046,N_5892);
nand U6063 (N_6063,N_5934,N_5875);
xnor U6064 (N_6064,N_5448,N_5149);
xor U6065 (N_6065,N_5885,N_5230);
nor U6066 (N_6066,N_5398,N_5159);
nand U6067 (N_6067,N_5809,N_5662);
nand U6068 (N_6068,N_5348,N_5256);
nand U6069 (N_6069,N_5008,N_5435);
or U6070 (N_6070,N_5456,N_5741);
nand U6071 (N_6071,N_5204,N_5591);
or U6072 (N_6072,N_5179,N_5639);
nand U6073 (N_6073,N_5317,N_5296);
nor U6074 (N_6074,N_5034,N_5430);
nand U6075 (N_6075,N_5125,N_5368);
or U6076 (N_6076,N_5078,N_5947);
or U6077 (N_6077,N_5422,N_5525);
xnor U6078 (N_6078,N_5813,N_5816);
and U6079 (N_6079,N_5927,N_5151);
nor U6080 (N_6080,N_5929,N_5189);
or U6081 (N_6081,N_5057,N_5572);
and U6082 (N_6082,N_5477,N_5669);
nor U6083 (N_6083,N_5366,N_5561);
or U6084 (N_6084,N_5201,N_5956);
nand U6085 (N_6085,N_5935,N_5966);
xnor U6086 (N_6086,N_5894,N_5026);
xnor U6087 (N_6087,N_5407,N_5489);
and U6088 (N_6088,N_5652,N_5583);
or U6089 (N_6089,N_5461,N_5136);
and U6090 (N_6090,N_5117,N_5796);
nand U6091 (N_6091,N_5560,N_5097);
nand U6092 (N_6092,N_5524,N_5410);
nor U6093 (N_6093,N_5336,N_5910);
nand U6094 (N_6094,N_5427,N_5989);
nor U6095 (N_6095,N_5724,N_5338);
nand U6096 (N_6096,N_5379,N_5312);
xnor U6097 (N_6097,N_5756,N_5099);
and U6098 (N_6098,N_5570,N_5621);
and U6099 (N_6099,N_5354,N_5092);
or U6100 (N_6100,N_5534,N_5386);
or U6101 (N_6101,N_5697,N_5631);
nor U6102 (N_6102,N_5007,N_5383);
nor U6103 (N_6103,N_5364,N_5167);
xnor U6104 (N_6104,N_5976,N_5423);
and U6105 (N_6105,N_5339,N_5978);
nor U6106 (N_6106,N_5872,N_5771);
xor U6107 (N_6107,N_5992,N_5102);
and U6108 (N_6108,N_5851,N_5987);
nand U6109 (N_6109,N_5031,N_5825);
nor U6110 (N_6110,N_5399,N_5458);
nor U6111 (N_6111,N_5882,N_5030);
xnor U6112 (N_6112,N_5634,N_5706);
xnor U6113 (N_6113,N_5404,N_5389);
or U6114 (N_6114,N_5231,N_5506);
nand U6115 (N_6115,N_5460,N_5758);
nor U6116 (N_6116,N_5126,N_5396);
or U6117 (N_6117,N_5916,N_5713);
and U6118 (N_6118,N_5447,N_5831);
xor U6119 (N_6119,N_5879,N_5562);
or U6120 (N_6120,N_5703,N_5109);
and U6121 (N_6121,N_5302,N_5580);
xor U6122 (N_6122,N_5076,N_5856);
and U6123 (N_6123,N_5245,N_5905);
and U6124 (N_6124,N_5229,N_5907);
and U6125 (N_6125,N_5363,N_5691);
nand U6126 (N_6126,N_5219,N_5252);
or U6127 (N_6127,N_5135,N_5536);
xor U6128 (N_6128,N_5020,N_5384);
xor U6129 (N_6129,N_5556,N_5217);
xnor U6130 (N_6130,N_5335,N_5763);
nand U6131 (N_6131,N_5134,N_5047);
or U6132 (N_6132,N_5058,N_5510);
nand U6133 (N_6133,N_5795,N_5564);
nand U6134 (N_6134,N_5801,N_5285);
nand U6135 (N_6135,N_5808,N_5522);
nand U6136 (N_6136,N_5378,N_5472);
nor U6137 (N_6137,N_5453,N_5158);
nand U6138 (N_6138,N_5838,N_5926);
nor U6139 (N_6139,N_5206,N_5819);
and U6140 (N_6140,N_5455,N_5610);
nand U6141 (N_6141,N_5543,N_5963);
nand U6142 (N_6142,N_5083,N_5177);
and U6143 (N_6143,N_5566,N_5883);
nand U6144 (N_6144,N_5501,N_5180);
and U6145 (N_6145,N_5818,N_5663);
nand U6146 (N_6146,N_5715,N_5131);
xor U6147 (N_6147,N_5859,N_5822);
nand U6148 (N_6148,N_5100,N_5984);
nand U6149 (N_6149,N_5866,N_5133);
and U6150 (N_6150,N_5620,N_5614);
nand U6151 (N_6151,N_5917,N_5001);
and U6152 (N_6152,N_5494,N_5165);
and U6153 (N_6153,N_5434,N_5174);
nand U6154 (N_6154,N_5199,N_5714);
xnor U6155 (N_6155,N_5860,N_5027);
nor U6156 (N_6156,N_5138,N_5640);
xnor U6157 (N_6157,N_5537,N_5836);
xnor U6158 (N_6158,N_5854,N_5792);
xor U6159 (N_6159,N_5038,N_5509);
and U6160 (N_6160,N_5635,N_5503);
or U6161 (N_6161,N_5225,N_5616);
nand U6162 (N_6162,N_5130,N_5708);
or U6163 (N_6163,N_5606,N_5327);
nand U6164 (N_6164,N_5920,N_5360);
xnor U6165 (N_6165,N_5720,N_5450);
nand U6166 (N_6166,N_5732,N_5937);
or U6167 (N_6167,N_5840,N_5666);
nor U6168 (N_6168,N_5906,N_5518);
nand U6169 (N_6169,N_5768,N_5548);
xnor U6170 (N_6170,N_5600,N_5791);
nand U6171 (N_6171,N_5555,N_5938);
nand U6172 (N_6172,N_5181,N_5943);
xor U6173 (N_6173,N_5952,N_5559);
nor U6174 (N_6174,N_5833,N_5579);
or U6175 (N_6175,N_5857,N_5535);
xnor U6176 (N_6176,N_5397,N_5214);
nand U6177 (N_6177,N_5847,N_5195);
xor U6178 (N_6178,N_5550,N_5696);
or U6179 (N_6179,N_5520,N_5357);
nand U6180 (N_6180,N_5006,N_5323);
or U6181 (N_6181,N_5250,N_5306);
or U6182 (N_6182,N_5584,N_5124);
xnor U6183 (N_6183,N_5022,N_5603);
nor U6184 (N_6184,N_5291,N_5050);
nor U6185 (N_6185,N_5557,N_5878);
nand U6186 (N_6186,N_5617,N_5582);
nand U6187 (N_6187,N_5998,N_5727);
xnor U6188 (N_6188,N_5161,N_5488);
xor U6189 (N_6189,N_5111,N_5193);
xnor U6190 (N_6190,N_5408,N_5690);
xor U6191 (N_6191,N_5168,N_5912);
nand U6192 (N_6192,N_5372,N_5340);
xnor U6193 (N_6193,N_5395,N_5182);
nand U6194 (N_6194,N_5400,N_5699);
or U6195 (N_6195,N_5266,N_5547);
nor U6196 (N_6196,N_5734,N_5154);
xor U6197 (N_6197,N_5757,N_5624);
or U6198 (N_6198,N_5655,N_5079);
xnor U6199 (N_6199,N_5769,N_5032);
nand U6200 (N_6200,N_5073,N_5781);
nor U6201 (N_6201,N_5457,N_5973);
xnor U6202 (N_6202,N_5542,N_5028);
or U6203 (N_6203,N_5514,N_5971);
nand U6204 (N_6204,N_5689,N_5183);
nand U6205 (N_6205,N_5721,N_5733);
or U6206 (N_6206,N_5321,N_5874);
nand U6207 (N_6207,N_5928,N_5401);
nand U6208 (N_6208,N_5292,N_5352);
xnor U6209 (N_6209,N_5411,N_5793);
nor U6210 (N_6210,N_5800,N_5356);
and U6211 (N_6211,N_5259,N_5517);
nand U6212 (N_6212,N_5261,N_5465);
xor U6213 (N_6213,N_5018,N_5108);
and U6214 (N_6214,N_5964,N_5473);
nand U6215 (N_6215,N_5970,N_5257);
and U6216 (N_6216,N_5139,N_5061);
nand U6217 (N_6217,N_5644,N_5554);
nor U6218 (N_6218,N_5123,N_5590);
and U6219 (N_6219,N_5674,N_5478);
xnor U6220 (N_6220,N_5205,N_5593);
xnor U6221 (N_6221,N_5661,N_5739);
or U6222 (N_6222,N_5750,N_5242);
xor U6223 (N_6223,N_5827,N_5037);
or U6224 (N_6224,N_5486,N_5063);
xor U6225 (N_6225,N_5980,N_5527);
or U6226 (N_6226,N_5649,N_5519);
nor U6227 (N_6227,N_5005,N_5533);
nor U6228 (N_6228,N_5909,N_5746);
nor U6229 (N_6229,N_5896,N_5283);
nand U6230 (N_6230,N_5986,N_5082);
nor U6231 (N_6231,N_5029,N_5675);
xor U6232 (N_6232,N_5611,N_5086);
nor U6233 (N_6233,N_5254,N_5490);
nand U6234 (N_6234,N_5173,N_5380);
nor U6235 (N_6235,N_5545,N_5420);
xnor U6236 (N_6236,N_5981,N_5500);
xor U6237 (N_6237,N_5913,N_5754);
and U6238 (N_6238,N_5576,N_5419);
or U6239 (N_6239,N_5688,N_5931);
nor U6240 (N_6240,N_5513,N_5495);
xor U6241 (N_6241,N_5071,N_5780);
xnor U6242 (N_6242,N_5526,N_5889);
xnor U6243 (N_6243,N_5824,N_5755);
nand U6244 (N_6244,N_5497,N_5232);
or U6245 (N_6245,N_5479,N_5678);
or U6246 (N_6246,N_5712,N_5350);
nor U6247 (N_6247,N_5122,N_5898);
xor U6248 (N_6248,N_5627,N_5160);
and U6249 (N_6249,N_5328,N_5729);
nand U6250 (N_6250,N_5351,N_5286);
xnor U6251 (N_6251,N_5392,N_5373);
nor U6252 (N_6252,N_5507,N_5143);
and U6253 (N_6253,N_5128,N_5299);
nand U6254 (N_6254,N_5070,N_5091);
and U6255 (N_6255,N_5272,N_5355);
or U6256 (N_6256,N_5806,N_5316);
and U6257 (N_6257,N_5784,N_5132);
or U6258 (N_6258,N_5726,N_5760);
nand U6259 (N_6259,N_5475,N_5995);
nor U6260 (N_6260,N_5651,N_5238);
xnor U6261 (N_6261,N_5051,N_5975);
xnor U6262 (N_6262,N_5650,N_5951);
and U6263 (N_6263,N_5633,N_5207);
nand U6264 (N_6264,N_5432,N_5942);
and U6265 (N_6265,N_5466,N_5187);
or U6266 (N_6266,N_5474,N_5228);
and U6267 (N_6267,N_5504,N_5248);
nor U6268 (N_6268,N_5394,N_5334);
xnor U6269 (N_6269,N_5835,N_5428);
nor U6270 (N_6270,N_5087,N_5630);
nand U6271 (N_6271,N_5371,N_5540);
and U6272 (N_6272,N_5711,N_5443);
xor U6273 (N_6273,N_5587,N_5777);
and U6274 (N_6274,N_5431,N_5459);
xor U6275 (N_6275,N_5991,N_5369);
nor U6276 (N_6276,N_5834,N_5439);
and U6277 (N_6277,N_5594,N_5056);
nand U6278 (N_6278,N_5839,N_5810);
xnor U6279 (N_6279,N_5679,N_5994);
or U6280 (N_6280,N_5065,N_5962);
or U6281 (N_6281,N_5698,N_5553);
nor U6282 (N_6282,N_5090,N_5023);
xnor U6283 (N_6283,N_5176,N_5300);
xor U6284 (N_6284,N_5737,N_5178);
nor U6285 (N_6285,N_5449,N_5345);
and U6286 (N_6286,N_5293,N_5367);
or U6287 (N_6287,N_5852,N_5060);
and U6288 (N_6288,N_5609,N_5681);
nand U6289 (N_6289,N_5766,N_5901);
xnor U6290 (N_6290,N_5508,N_5880);
or U6291 (N_6291,N_5551,N_5843);
nand U6292 (N_6292,N_5961,N_5324);
and U6293 (N_6293,N_5121,N_5251);
xor U6294 (N_6294,N_5709,N_5493);
nor U6295 (N_6295,N_5484,N_5045);
and U6296 (N_6296,N_5502,N_5865);
xor U6297 (N_6297,N_5370,N_5331);
nand U6298 (N_6298,N_5972,N_5764);
or U6299 (N_6299,N_5573,N_5314);
nor U6300 (N_6300,N_5753,N_5802);
nand U6301 (N_6301,N_5923,N_5884);
and U6302 (N_6302,N_5377,N_5773);
xor U6303 (N_6303,N_5164,N_5264);
nor U6304 (N_6304,N_5024,N_5789);
or U6305 (N_6305,N_5805,N_5779);
nand U6306 (N_6306,N_5094,N_5983);
or U6307 (N_6307,N_5871,N_5096);
nand U6308 (N_6308,N_5823,N_5237);
nor U6309 (N_6309,N_5003,N_5288);
or U6310 (N_6310,N_5608,N_5011);
xnor U6311 (N_6311,N_5599,N_5393);
or U6312 (N_6312,N_5767,N_5255);
xor U6313 (N_6313,N_5429,N_5743);
nor U6314 (N_6314,N_5597,N_5999);
nand U6315 (N_6315,N_5749,N_5683);
nor U6316 (N_6316,N_5645,N_5902);
or U6317 (N_6317,N_5832,N_5062);
or U6318 (N_6318,N_5731,N_5702);
and U6319 (N_6319,N_5191,N_5589);
nand U6320 (N_6320,N_5303,N_5939);
and U6321 (N_6321,N_5960,N_5166);
nand U6322 (N_6322,N_5632,N_5342);
xnor U6323 (N_6323,N_5774,N_5770);
nand U6324 (N_6324,N_5638,N_5850);
or U6325 (N_6325,N_5365,N_5004);
and U6326 (N_6326,N_5586,N_5095);
and U6327 (N_6327,N_5425,N_5641);
xnor U6328 (N_6328,N_5469,N_5175);
xnor U6329 (N_6329,N_5233,N_5725);
nand U6330 (N_6330,N_5863,N_5381);
xor U6331 (N_6331,N_5665,N_5619);
and U6332 (N_6332,N_5362,N_5200);
xnor U6333 (N_6333,N_5988,N_5908);
xor U6334 (N_6334,N_5142,N_5115);
or U6335 (N_6335,N_5765,N_5969);
and U6336 (N_6336,N_5119,N_5471);
nor U6337 (N_6337,N_5155,N_5812);
or U6338 (N_6338,N_5783,N_5499);
nor U6339 (N_6339,N_5330,N_5849);
nand U6340 (N_6340,N_5612,N_5436);
nand U6341 (N_6341,N_5613,N_5761);
nor U6342 (N_6342,N_5343,N_5156);
nand U6343 (N_6343,N_5922,N_5297);
and U6344 (N_6344,N_5748,N_5899);
and U6345 (N_6345,N_5241,N_5332);
nor U6346 (N_6346,N_5414,N_5275);
nor U6347 (N_6347,N_5269,N_5388);
nand U6348 (N_6348,N_5745,N_5157);
xnor U6349 (N_6349,N_5224,N_5064);
or U6350 (N_6350,N_5141,N_5347);
nand U6351 (N_6351,N_5218,N_5762);
nand U6352 (N_6352,N_5271,N_5044);
nor U6353 (N_6353,N_5914,N_5626);
nand U6354 (N_6354,N_5129,N_5444);
nand U6355 (N_6355,N_5442,N_5869);
and U6356 (N_6356,N_5904,N_5040);
nand U6357 (N_6357,N_5830,N_5605);
xor U6358 (N_6358,N_5585,N_5120);
xor U6359 (N_6359,N_5895,N_5387);
and U6360 (N_6360,N_5873,N_5890);
and U6361 (N_6361,N_5150,N_5185);
xor U6362 (N_6362,N_5325,N_5837);
xor U6363 (N_6363,N_5546,N_5452);
xor U6364 (N_6364,N_5670,N_5629);
and U6365 (N_6365,N_5304,N_5864);
nor U6366 (N_6366,N_5281,N_5440);
nor U6367 (N_6367,N_5870,N_5977);
nand U6368 (N_6368,N_5482,N_5657);
and U6369 (N_6369,N_5144,N_5877);
nor U6370 (N_6370,N_5563,N_5035);
xor U6371 (N_6371,N_5933,N_5704);
and U6372 (N_6372,N_5467,N_5375);
or U6373 (N_6373,N_5803,N_5487);
nand U6374 (N_6374,N_5009,N_5868);
nor U6375 (N_6375,N_5318,N_5979);
xor U6376 (N_6376,N_5680,N_5886);
xnor U6377 (N_6377,N_5595,N_5786);
and U6378 (N_6378,N_5772,N_5887);
xor U6379 (N_6379,N_5235,N_5417);
xnor U6380 (N_6380,N_5322,N_5298);
xnor U6381 (N_6381,N_5636,N_5013);
xnor U6382 (N_6382,N_5049,N_5660);
xor U6383 (N_6383,N_5391,N_5249);
nand U6384 (N_6384,N_5267,N_5575);
xor U6385 (N_6385,N_5170,N_5017);
and U6386 (N_6386,N_5221,N_5274);
or U6387 (N_6387,N_5127,N_5692);
and U6388 (N_6388,N_5668,N_5828);
and U6389 (N_6389,N_5376,N_5239);
xnor U6390 (N_6390,N_5069,N_5646);
nor U6391 (N_6391,N_5891,N_5068);
nand U6392 (N_6392,N_5740,N_5911);
or U6393 (N_6393,N_5787,N_5511);
and U6394 (N_6394,N_5216,N_5137);
nor U6395 (N_6395,N_5930,N_5140);
or U6396 (N_6396,N_5985,N_5287);
or U6397 (N_6397,N_5742,N_5084);
nand U6398 (N_6398,N_5247,N_5080);
and U6399 (N_6399,N_5222,N_5485);
nor U6400 (N_6400,N_5492,N_5571);
nand U6401 (N_6401,N_5313,N_5234);
nor U6402 (N_6402,N_5932,N_5628);
and U6403 (N_6403,N_5853,N_5867);
and U6404 (N_6404,N_5588,N_5530);
and U6405 (N_6405,N_5390,N_5446);
nor U6406 (N_6406,N_5268,N_5042);
and U6407 (N_6407,N_5212,N_5759);
nor U6408 (N_6408,N_5067,N_5103);
nor U6409 (N_6409,N_5413,N_5110);
and U6410 (N_6410,N_5858,N_5574);
or U6411 (N_6411,N_5654,N_5202);
nor U6412 (N_6412,N_5685,N_5244);
xnor U6413 (N_6413,N_5105,N_5451);
nand U6414 (N_6414,N_5015,N_5936);
xnor U6415 (N_6415,N_5815,N_5162);
xor U6416 (N_6416,N_5967,N_5925);
or U6417 (N_6417,N_5265,N_5710);
nand U6418 (N_6418,N_5659,N_5747);
xnor U6419 (N_6419,N_5918,N_5811);
nand U6420 (N_6420,N_5728,N_5054);
nand U6421 (N_6421,N_5211,N_5705);
or U6422 (N_6422,N_5113,N_5016);
xor U6423 (N_6423,N_5941,N_5186);
nor U6424 (N_6424,N_5262,N_5707);
or U6425 (N_6425,N_5671,N_5209);
xor U6426 (N_6426,N_5021,N_5043);
nor U6427 (N_6427,N_5505,N_5041);
xnor U6428 (N_6428,N_5223,N_5532);
or U6429 (N_6429,N_5098,N_5569);
nand U6430 (N_6430,N_5751,N_5101);
nand U6431 (N_6431,N_5955,N_5673);
nand U6432 (N_6432,N_5512,N_5694);
nand U6433 (N_6433,N_5950,N_5676);
and U6434 (N_6434,N_5409,N_5953);
or U6435 (N_6435,N_5776,N_5567);
nand U6436 (N_6436,N_5308,N_5311);
xor U6437 (N_6437,N_5785,N_5277);
nand U6438 (N_6438,N_5799,N_5059);
nand U6439 (N_6439,N_5491,N_5341);
or U6440 (N_6440,N_5418,N_5814);
nor U6441 (N_6441,N_5648,N_5944);
xnor U6442 (N_6442,N_5719,N_5656);
and U6443 (N_6443,N_5353,N_5116);
nand U6444 (N_6444,N_5415,N_5807);
nand U6445 (N_6445,N_5470,N_5496);
nand U6446 (N_6446,N_5684,N_5075);
nand U6447 (N_6447,N_5552,N_5301);
or U6448 (N_6448,N_5515,N_5826);
or U6449 (N_6449,N_5258,N_5438);
and U6450 (N_6450,N_5289,N_5437);
nand U6451 (N_6451,N_5658,N_5310);
or U6452 (N_6452,N_5948,N_5664);
and U6453 (N_6453,N_5647,N_5163);
or U6454 (N_6454,N_5592,N_5169);
and U6455 (N_6455,N_5722,N_5188);
nand U6456 (N_6456,N_5622,N_5329);
nand U6457 (N_6457,N_5541,N_5687);
and U6458 (N_6458,N_5996,N_5959);
or U6459 (N_6459,N_5821,N_5424);
nor U6460 (N_6460,N_5565,N_5903);
nor U6461 (N_6461,N_5581,N_5074);
xor U6462 (N_6462,N_5531,N_5385);
or U6463 (N_6463,N_5464,N_5114);
nor U6464 (N_6464,N_5279,N_5361);
and U6465 (N_6465,N_5643,N_5788);
or U6466 (N_6466,N_5441,N_5695);
and U6467 (N_6467,N_5735,N_5893);
nor U6468 (N_6468,N_5949,N_5817);
xor U6469 (N_6469,N_5106,N_5260);
or U6470 (N_6470,N_5014,N_5421);
xor U6471 (N_6471,N_5405,N_5402);
xnor U6472 (N_6472,N_5145,N_5118);
or U6473 (N_6473,N_5846,N_5607);
and U6474 (N_6474,N_5010,N_5454);
xnor U6475 (N_6475,N_5716,N_5033);
nor U6476 (N_6476,N_5462,N_5481);
or U6477 (N_6477,N_5295,N_5374);
nand U6478 (N_6478,N_5000,N_5077);
or U6479 (N_6479,N_5797,N_5406);
nor U6480 (N_6480,N_5848,N_5220);
xor U6481 (N_6481,N_5538,N_5333);
nand U6482 (N_6482,N_5677,N_5568);
or U6483 (N_6483,N_5236,N_5172);
nor U6484 (N_6484,N_5198,N_5578);
nor U6485 (N_6485,N_5717,N_5085);
nand U6486 (N_6486,N_5539,N_5403);
or U6487 (N_6487,N_5738,N_5055);
or U6488 (N_6488,N_5382,N_5862);
nor U6489 (N_6489,N_5790,N_5349);
xnor U6490 (N_6490,N_5243,N_5346);
nor U6491 (N_6491,N_5845,N_5263);
xnor U6492 (N_6492,N_5309,N_5107);
nand U6493 (N_6493,N_5284,N_5002);
or U6494 (N_6494,N_5337,N_5723);
or U6495 (N_6495,N_5290,N_5820);
nand U6496 (N_6496,N_5358,N_5618);
and U6497 (N_6497,N_5412,N_5653);
nand U6498 (N_6498,N_5190,N_5549);
or U6499 (N_6499,N_5946,N_5782);
nor U6500 (N_6500,N_5655,N_5974);
nand U6501 (N_6501,N_5264,N_5868);
or U6502 (N_6502,N_5283,N_5985);
xor U6503 (N_6503,N_5247,N_5942);
nor U6504 (N_6504,N_5796,N_5160);
xnor U6505 (N_6505,N_5918,N_5651);
and U6506 (N_6506,N_5912,N_5906);
nor U6507 (N_6507,N_5060,N_5442);
nand U6508 (N_6508,N_5020,N_5693);
and U6509 (N_6509,N_5603,N_5591);
and U6510 (N_6510,N_5435,N_5399);
xor U6511 (N_6511,N_5570,N_5693);
xor U6512 (N_6512,N_5940,N_5597);
xor U6513 (N_6513,N_5060,N_5999);
xnor U6514 (N_6514,N_5226,N_5874);
or U6515 (N_6515,N_5095,N_5057);
and U6516 (N_6516,N_5221,N_5494);
nand U6517 (N_6517,N_5363,N_5897);
nor U6518 (N_6518,N_5314,N_5927);
or U6519 (N_6519,N_5649,N_5532);
or U6520 (N_6520,N_5213,N_5955);
nand U6521 (N_6521,N_5257,N_5540);
xnor U6522 (N_6522,N_5799,N_5427);
or U6523 (N_6523,N_5331,N_5131);
nand U6524 (N_6524,N_5959,N_5932);
nand U6525 (N_6525,N_5537,N_5427);
nand U6526 (N_6526,N_5094,N_5457);
nand U6527 (N_6527,N_5432,N_5539);
nand U6528 (N_6528,N_5984,N_5263);
or U6529 (N_6529,N_5661,N_5844);
and U6530 (N_6530,N_5599,N_5561);
or U6531 (N_6531,N_5386,N_5445);
and U6532 (N_6532,N_5199,N_5554);
or U6533 (N_6533,N_5927,N_5958);
and U6534 (N_6534,N_5085,N_5819);
and U6535 (N_6535,N_5256,N_5197);
nor U6536 (N_6536,N_5328,N_5182);
and U6537 (N_6537,N_5302,N_5069);
nand U6538 (N_6538,N_5990,N_5801);
nor U6539 (N_6539,N_5248,N_5059);
and U6540 (N_6540,N_5682,N_5971);
nor U6541 (N_6541,N_5293,N_5674);
nor U6542 (N_6542,N_5954,N_5022);
or U6543 (N_6543,N_5045,N_5275);
or U6544 (N_6544,N_5968,N_5645);
and U6545 (N_6545,N_5207,N_5968);
and U6546 (N_6546,N_5495,N_5259);
xor U6547 (N_6547,N_5378,N_5381);
or U6548 (N_6548,N_5345,N_5885);
or U6549 (N_6549,N_5518,N_5502);
xnor U6550 (N_6550,N_5362,N_5529);
xor U6551 (N_6551,N_5941,N_5477);
nand U6552 (N_6552,N_5927,N_5759);
and U6553 (N_6553,N_5592,N_5837);
nor U6554 (N_6554,N_5804,N_5728);
and U6555 (N_6555,N_5158,N_5499);
nor U6556 (N_6556,N_5113,N_5706);
or U6557 (N_6557,N_5790,N_5911);
and U6558 (N_6558,N_5816,N_5716);
xor U6559 (N_6559,N_5468,N_5745);
nor U6560 (N_6560,N_5948,N_5682);
xor U6561 (N_6561,N_5066,N_5559);
nand U6562 (N_6562,N_5823,N_5665);
or U6563 (N_6563,N_5914,N_5441);
or U6564 (N_6564,N_5064,N_5836);
nand U6565 (N_6565,N_5935,N_5331);
nor U6566 (N_6566,N_5577,N_5765);
nand U6567 (N_6567,N_5019,N_5494);
nor U6568 (N_6568,N_5428,N_5914);
or U6569 (N_6569,N_5174,N_5474);
nor U6570 (N_6570,N_5343,N_5362);
nor U6571 (N_6571,N_5958,N_5398);
nor U6572 (N_6572,N_5210,N_5402);
nor U6573 (N_6573,N_5830,N_5115);
xor U6574 (N_6574,N_5397,N_5003);
xor U6575 (N_6575,N_5358,N_5694);
nand U6576 (N_6576,N_5283,N_5560);
or U6577 (N_6577,N_5071,N_5498);
xor U6578 (N_6578,N_5762,N_5874);
xor U6579 (N_6579,N_5001,N_5353);
xnor U6580 (N_6580,N_5789,N_5219);
nand U6581 (N_6581,N_5679,N_5816);
or U6582 (N_6582,N_5473,N_5919);
nand U6583 (N_6583,N_5887,N_5901);
nor U6584 (N_6584,N_5806,N_5391);
nor U6585 (N_6585,N_5611,N_5847);
nand U6586 (N_6586,N_5247,N_5811);
or U6587 (N_6587,N_5954,N_5518);
nor U6588 (N_6588,N_5674,N_5935);
and U6589 (N_6589,N_5424,N_5976);
nor U6590 (N_6590,N_5381,N_5851);
and U6591 (N_6591,N_5897,N_5319);
and U6592 (N_6592,N_5096,N_5490);
nor U6593 (N_6593,N_5093,N_5646);
and U6594 (N_6594,N_5834,N_5876);
nand U6595 (N_6595,N_5198,N_5421);
nor U6596 (N_6596,N_5879,N_5161);
xnor U6597 (N_6597,N_5995,N_5963);
nand U6598 (N_6598,N_5229,N_5821);
xor U6599 (N_6599,N_5193,N_5849);
nor U6600 (N_6600,N_5497,N_5946);
nand U6601 (N_6601,N_5645,N_5858);
or U6602 (N_6602,N_5255,N_5986);
and U6603 (N_6603,N_5124,N_5468);
and U6604 (N_6604,N_5051,N_5390);
or U6605 (N_6605,N_5700,N_5211);
and U6606 (N_6606,N_5563,N_5355);
nand U6607 (N_6607,N_5921,N_5472);
nor U6608 (N_6608,N_5569,N_5249);
and U6609 (N_6609,N_5065,N_5524);
and U6610 (N_6610,N_5838,N_5962);
and U6611 (N_6611,N_5632,N_5726);
or U6612 (N_6612,N_5326,N_5529);
and U6613 (N_6613,N_5824,N_5750);
xor U6614 (N_6614,N_5533,N_5334);
nand U6615 (N_6615,N_5082,N_5601);
xor U6616 (N_6616,N_5058,N_5633);
or U6617 (N_6617,N_5972,N_5514);
xnor U6618 (N_6618,N_5685,N_5609);
nor U6619 (N_6619,N_5202,N_5240);
nand U6620 (N_6620,N_5551,N_5612);
and U6621 (N_6621,N_5978,N_5940);
nor U6622 (N_6622,N_5458,N_5952);
xor U6623 (N_6623,N_5627,N_5813);
and U6624 (N_6624,N_5109,N_5104);
and U6625 (N_6625,N_5150,N_5983);
and U6626 (N_6626,N_5233,N_5736);
nor U6627 (N_6627,N_5209,N_5082);
or U6628 (N_6628,N_5372,N_5891);
xor U6629 (N_6629,N_5681,N_5782);
and U6630 (N_6630,N_5641,N_5568);
nand U6631 (N_6631,N_5122,N_5969);
nor U6632 (N_6632,N_5149,N_5796);
and U6633 (N_6633,N_5785,N_5678);
or U6634 (N_6634,N_5117,N_5820);
xor U6635 (N_6635,N_5244,N_5963);
nor U6636 (N_6636,N_5624,N_5282);
nor U6637 (N_6637,N_5026,N_5394);
and U6638 (N_6638,N_5263,N_5344);
and U6639 (N_6639,N_5550,N_5775);
and U6640 (N_6640,N_5181,N_5752);
and U6641 (N_6641,N_5236,N_5138);
xor U6642 (N_6642,N_5374,N_5973);
nor U6643 (N_6643,N_5265,N_5248);
or U6644 (N_6644,N_5448,N_5335);
and U6645 (N_6645,N_5383,N_5810);
or U6646 (N_6646,N_5428,N_5596);
nand U6647 (N_6647,N_5776,N_5518);
xor U6648 (N_6648,N_5693,N_5092);
or U6649 (N_6649,N_5412,N_5027);
and U6650 (N_6650,N_5830,N_5175);
nor U6651 (N_6651,N_5547,N_5263);
or U6652 (N_6652,N_5418,N_5825);
or U6653 (N_6653,N_5637,N_5215);
nand U6654 (N_6654,N_5180,N_5960);
and U6655 (N_6655,N_5194,N_5793);
xor U6656 (N_6656,N_5802,N_5856);
xor U6657 (N_6657,N_5070,N_5811);
nor U6658 (N_6658,N_5434,N_5621);
xor U6659 (N_6659,N_5705,N_5346);
and U6660 (N_6660,N_5937,N_5557);
xnor U6661 (N_6661,N_5914,N_5764);
nor U6662 (N_6662,N_5881,N_5337);
nand U6663 (N_6663,N_5089,N_5457);
nand U6664 (N_6664,N_5928,N_5596);
and U6665 (N_6665,N_5677,N_5742);
or U6666 (N_6666,N_5163,N_5791);
and U6667 (N_6667,N_5999,N_5719);
and U6668 (N_6668,N_5543,N_5626);
and U6669 (N_6669,N_5308,N_5741);
xnor U6670 (N_6670,N_5814,N_5178);
xnor U6671 (N_6671,N_5756,N_5354);
nor U6672 (N_6672,N_5325,N_5662);
and U6673 (N_6673,N_5857,N_5272);
nand U6674 (N_6674,N_5613,N_5605);
nand U6675 (N_6675,N_5650,N_5731);
nor U6676 (N_6676,N_5048,N_5351);
or U6677 (N_6677,N_5275,N_5947);
nand U6678 (N_6678,N_5278,N_5703);
xnor U6679 (N_6679,N_5797,N_5001);
nand U6680 (N_6680,N_5971,N_5681);
and U6681 (N_6681,N_5386,N_5791);
nor U6682 (N_6682,N_5682,N_5336);
xor U6683 (N_6683,N_5247,N_5344);
nor U6684 (N_6684,N_5291,N_5999);
xor U6685 (N_6685,N_5894,N_5589);
or U6686 (N_6686,N_5749,N_5069);
xor U6687 (N_6687,N_5604,N_5188);
and U6688 (N_6688,N_5768,N_5083);
or U6689 (N_6689,N_5575,N_5198);
and U6690 (N_6690,N_5732,N_5617);
nor U6691 (N_6691,N_5132,N_5100);
nor U6692 (N_6692,N_5115,N_5971);
nor U6693 (N_6693,N_5998,N_5889);
and U6694 (N_6694,N_5972,N_5558);
and U6695 (N_6695,N_5691,N_5410);
xnor U6696 (N_6696,N_5143,N_5791);
xor U6697 (N_6697,N_5371,N_5446);
or U6698 (N_6698,N_5839,N_5375);
nand U6699 (N_6699,N_5595,N_5544);
and U6700 (N_6700,N_5410,N_5004);
and U6701 (N_6701,N_5308,N_5733);
nor U6702 (N_6702,N_5519,N_5175);
xnor U6703 (N_6703,N_5289,N_5751);
xnor U6704 (N_6704,N_5829,N_5384);
xnor U6705 (N_6705,N_5982,N_5381);
nor U6706 (N_6706,N_5945,N_5976);
and U6707 (N_6707,N_5586,N_5954);
nor U6708 (N_6708,N_5258,N_5671);
xnor U6709 (N_6709,N_5624,N_5174);
or U6710 (N_6710,N_5230,N_5565);
nand U6711 (N_6711,N_5043,N_5568);
xnor U6712 (N_6712,N_5780,N_5376);
xnor U6713 (N_6713,N_5712,N_5981);
or U6714 (N_6714,N_5699,N_5519);
nand U6715 (N_6715,N_5777,N_5067);
or U6716 (N_6716,N_5670,N_5271);
xnor U6717 (N_6717,N_5221,N_5043);
nor U6718 (N_6718,N_5242,N_5156);
and U6719 (N_6719,N_5538,N_5952);
and U6720 (N_6720,N_5427,N_5321);
nor U6721 (N_6721,N_5817,N_5699);
or U6722 (N_6722,N_5603,N_5007);
or U6723 (N_6723,N_5894,N_5188);
xnor U6724 (N_6724,N_5109,N_5294);
nand U6725 (N_6725,N_5242,N_5996);
xnor U6726 (N_6726,N_5917,N_5190);
nor U6727 (N_6727,N_5571,N_5180);
and U6728 (N_6728,N_5037,N_5306);
and U6729 (N_6729,N_5156,N_5227);
or U6730 (N_6730,N_5635,N_5992);
and U6731 (N_6731,N_5149,N_5942);
or U6732 (N_6732,N_5732,N_5188);
and U6733 (N_6733,N_5032,N_5671);
and U6734 (N_6734,N_5067,N_5849);
or U6735 (N_6735,N_5012,N_5049);
xnor U6736 (N_6736,N_5337,N_5296);
xor U6737 (N_6737,N_5605,N_5657);
xor U6738 (N_6738,N_5496,N_5563);
nand U6739 (N_6739,N_5366,N_5472);
or U6740 (N_6740,N_5958,N_5544);
nand U6741 (N_6741,N_5736,N_5696);
or U6742 (N_6742,N_5784,N_5959);
or U6743 (N_6743,N_5704,N_5074);
and U6744 (N_6744,N_5322,N_5496);
nor U6745 (N_6745,N_5598,N_5188);
nand U6746 (N_6746,N_5336,N_5898);
and U6747 (N_6747,N_5818,N_5099);
xnor U6748 (N_6748,N_5321,N_5359);
nand U6749 (N_6749,N_5512,N_5156);
xor U6750 (N_6750,N_5956,N_5284);
or U6751 (N_6751,N_5377,N_5825);
and U6752 (N_6752,N_5924,N_5939);
nand U6753 (N_6753,N_5009,N_5993);
nand U6754 (N_6754,N_5394,N_5949);
and U6755 (N_6755,N_5815,N_5266);
and U6756 (N_6756,N_5251,N_5285);
and U6757 (N_6757,N_5362,N_5036);
or U6758 (N_6758,N_5113,N_5609);
or U6759 (N_6759,N_5116,N_5279);
nand U6760 (N_6760,N_5108,N_5542);
nand U6761 (N_6761,N_5474,N_5553);
nor U6762 (N_6762,N_5536,N_5388);
and U6763 (N_6763,N_5498,N_5490);
xnor U6764 (N_6764,N_5820,N_5849);
nand U6765 (N_6765,N_5854,N_5393);
and U6766 (N_6766,N_5315,N_5578);
nand U6767 (N_6767,N_5870,N_5988);
and U6768 (N_6768,N_5804,N_5602);
nand U6769 (N_6769,N_5257,N_5711);
xnor U6770 (N_6770,N_5056,N_5934);
nor U6771 (N_6771,N_5248,N_5899);
xor U6772 (N_6772,N_5856,N_5836);
and U6773 (N_6773,N_5243,N_5535);
xnor U6774 (N_6774,N_5624,N_5432);
xnor U6775 (N_6775,N_5922,N_5363);
or U6776 (N_6776,N_5073,N_5384);
and U6777 (N_6777,N_5438,N_5992);
xor U6778 (N_6778,N_5675,N_5072);
nand U6779 (N_6779,N_5108,N_5515);
and U6780 (N_6780,N_5805,N_5449);
xnor U6781 (N_6781,N_5178,N_5700);
nand U6782 (N_6782,N_5319,N_5850);
nor U6783 (N_6783,N_5592,N_5734);
nand U6784 (N_6784,N_5150,N_5008);
and U6785 (N_6785,N_5220,N_5230);
and U6786 (N_6786,N_5479,N_5081);
nor U6787 (N_6787,N_5061,N_5870);
xor U6788 (N_6788,N_5366,N_5771);
xnor U6789 (N_6789,N_5251,N_5258);
nand U6790 (N_6790,N_5985,N_5479);
or U6791 (N_6791,N_5173,N_5662);
nand U6792 (N_6792,N_5713,N_5746);
nor U6793 (N_6793,N_5409,N_5047);
and U6794 (N_6794,N_5668,N_5401);
xnor U6795 (N_6795,N_5430,N_5839);
xor U6796 (N_6796,N_5307,N_5058);
nand U6797 (N_6797,N_5004,N_5013);
nand U6798 (N_6798,N_5170,N_5668);
nand U6799 (N_6799,N_5153,N_5045);
and U6800 (N_6800,N_5643,N_5974);
nand U6801 (N_6801,N_5041,N_5630);
and U6802 (N_6802,N_5568,N_5117);
nand U6803 (N_6803,N_5908,N_5372);
xnor U6804 (N_6804,N_5616,N_5982);
and U6805 (N_6805,N_5302,N_5674);
nand U6806 (N_6806,N_5773,N_5925);
xor U6807 (N_6807,N_5266,N_5942);
xnor U6808 (N_6808,N_5130,N_5515);
xor U6809 (N_6809,N_5435,N_5136);
nand U6810 (N_6810,N_5551,N_5913);
xor U6811 (N_6811,N_5005,N_5048);
and U6812 (N_6812,N_5311,N_5667);
nor U6813 (N_6813,N_5920,N_5531);
nor U6814 (N_6814,N_5954,N_5883);
and U6815 (N_6815,N_5153,N_5062);
xor U6816 (N_6816,N_5383,N_5138);
or U6817 (N_6817,N_5618,N_5995);
nor U6818 (N_6818,N_5839,N_5777);
nand U6819 (N_6819,N_5559,N_5278);
nand U6820 (N_6820,N_5376,N_5571);
or U6821 (N_6821,N_5804,N_5827);
nand U6822 (N_6822,N_5775,N_5814);
nand U6823 (N_6823,N_5729,N_5964);
nor U6824 (N_6824,N_5562,N_5926);
xor U6825 (N_6825,N_5079,N_5155);
xor U6826 (N_6826,N_5371,N_5763);
or U6827 (N_6827,N_5007,N_5554);
nand U6828 (N_6828,N_5728,N_5317);
xnor U6829 (N_6829,N_5464,N_5533);
nor U6830 (N_6830,N_5299,N_5443);
nor U6831 (N_6831,N_5246,N_5265);
nor U6832 (N_6832,N_5407,N_5365);
and U6833 (N_6833,N_5160,N_5474);
nand U6834 (N_6834,N_5326,N_5149);
nand U6835 (N_6835,N_5340,N_5656);
nand U6836 (N_6836,N_5874,N_5006);
or U6837 (N_6837,N_5146,N_5636);
xor U6838 (N_6838,N_5316,N_5451);
or U6839 (N_6839,N_5127,N_5634);
or U6840 (N_6840,N_5700,N_5162);
nand U6841 (N_6841,N_5897,N_5033);
and U6842 (N_6842,N_5419,N_5646);
xnor U6843 (N_6843,N_5968,N_5960);
nor U6844 (N_6844,N_5529,N_5120);
nand U6845 (N_6845,N_5618,N_5547);
or U6846 (N_6846,N_5553,N_5390);
nor U6847 (N_6847,N_5754,N_5743);
xnor U6848 (N_6848,N_5766,N_5445);
xor U6849 (N_6849,N_5026,N_5996);
nor U6850 (N_6850,N_5036,N_5465);
or U6851 (N_6851,N_5238,N_5710);
and U6852 (N_6852,N_5349,N_5639);
nand U6853 (N_6853,N_5404,N_5973);
xor U6854 (N_6854,N_5374,N_5892);
xor U6855 (N_6855,N_5857,N_5436);
and U6856 (N_6856,N_5795,N_5405);
nand U6857 (N_6857,N_5891,N_5877);
nand U6858 (N_6858,N_5114,N_5016);
and U6859 (N_6859,N_5698,N_5193);
nand U6860 (N_6860,N_5294,N_5473);
nor U6861 (N_6861,N_5551,N_5641);
nand U6862 (N_6862,N_5106,N_5730);
and U6863 (N_6863,N_5456,N_5919);
nand U6864 (N_6864,N_5325,N_5112);
or U6865 (N_6865,N_5963,N_5648);
and U6866 (N_6866,N_5946,N_5467);
xor U6867 (N_6867,N_5141,N_5172);
or U6868 (N_6868,N_5413,N_5927);
or U6869 (N_6869,N_5210,N_5760);
nor U6870 (N_6870,N_5941,N_5778);
or U6871 (N_6871,N_5586,N_5447);
or U6872 (N_6872,N_5433,N_5667);
nor U6873 (N_6873,N_5659,N_5390);
nand U6874 (N_6874,N_5288,N_5956);
or U6875 (N_6875,N_5902,N_5017);
nor U6876 (N_6876,N_5017,N_5837);
or U6877 (N_6877,N_5671,N_5233);
or U6878 (N_6878,N_5717,N_5023);
and U6879 (N_6879,N_5888,N_5849);
xnor U6880 (N_6880,N_5721,N_5797);
or U6881 (N_6881,N_5423,N_5711);
or U6882 (N_6882,N_5452,N_5295);
or U6883 (N_6883,N_5983,N_5065);
and U6884 (N_6884,N_5066,N_5016);
or U6885 (N_6885,N_5060,N_5217);
nand U6886 (N_6886,N_5093,N_5805);
nor U6887 (N_6887,N_5947,N_5301);
or U6888 (N_6888,N_5022,N_5731);
or U6889 (N_6889,N_5493,N_5944);
nor U6890 (N_6890,N_5884,N_5990);
xor U6891 (N_6891,N_5900,N_5804);
nand U6892 (N_6892,N_5561,N_5139);
and U6893 (N_6893,N_5876,N_5808);
and U6894 (N_6894,N_5017,N_5298);
and U6895 (N_6895,N_5287,N_5218);
nand U6896 (N_6896,N_5915,N_5766);
nand U6897 (N_6897,N_5263,N_5203);
or U6898 (N_6898,N_5165,N_5155);
and U6899 (N_6899,N_5307,N_5042);
nor U6900 (N_6900,N_5375,N_5588);
xnor U6901 (N_6901,N_5219,N_5917);
and U6902 (N_6902,N_5096,N_5562);
or U6903 (N_6903,N_5362,N_5396);
and U6904 (N_6904,N_5584,N_5143);
nand U6905 (N_6905,N_5269,N_5205);
nand U6906 (N_6906,N_5610,N_5205);
and U6907 (N_6907,N_5290,N_5666);
or U6908 (N_6908,N_5267,N_5531);
or U6909 (N_6909,N_5488,N_5290);
xor U6910 (N_6910,N_5276,N_5123);
nor U6911 (N_6911,N_5604,N_5015);
nor U6912 (N_6912,N_5515,N_5866);
or U6913 (N_6913,N_5619,N_5839);
nand U6914 (N_6914,N_5918,N_5389);
nor U6915 (N_6915,N_5683,N_5271);
and U6916 (N_6916,N_5063,N_5483);
nor U6917 (N_6917,N_5115,N_5503);
nand U6918 (N_6918,N_5422,N_5094);
xnor U6919 (N_6919,N_5955,N_5142);
and U6920 (N_6920,N_5630,N_5515);
or U6921 (N_6921,N_5841,N_5421);
or U6922 (N_6922,N_5299,N_5596);
xor U6923 (N_6923,N_5838,N_5361);
xor U6924 (N_6924,N_5658,N_5735);
nand U6925 (N_6925,N_5965,N_5009);
nand U6926 (N_6926,N_5994,N_5294);
and U6927 (N_6927,N_5220,N_5722);
nor U6928 (N_6928,N_5387,N_5231);
nand U6929 (N_6929,N_5980,N_5024);
nor U6930 (N_6930,N_5309,N_5434);
nand U6931 (N_6931,N_5528,N_5603);
nor U6932 (N_6932,N_5022,N_5721);
and U6933 (N_6933,N_5837,N_5632);
nand U6934 (N_6934,N_5754,N_5452);
xor U6935 (N_6935,N_5791,N_5221);
or U6936 (N_6936,N_5059,N_5640);
and U6937 (N_6937,N_5868,N_5373);
nand U6938 (N_6938,N_5050,N_5299);
nor U6939 (N_6939,N_5027,N_5450);
and U6940 (N_6940,N_5173,N_5492);
xor U6941 (N_6941,N_5609,N_5978);
or U6942 (N_6942,N_5227,N_5426);
nor U6943 (N_6943,N_5722,N_5709);
or U6944 (N_6944,N_5512,N_5378);
nor U6945 (N_6945,N_5755,N_5267);
nor U6946 (N_6946,N_5450,N_5894);
nand U6947 (N_6947,N_5393,N_5201);
nor U6948 (N_6948,N_5817,N_5082);
xnor U6949 (N_6949,N_5632,N_5580);
nand U6950 (N_6950,N_5242,N_5466);
xor U6951 (N_6951,N_5724,N_5583);
nor U6952 (N_6952,N_5342,N_5109);
nor U6953 (N_6953,N_5458,N_5420);
nor U6954 (N_6954,N_5661,N_5967);
or U6955 (N_6955,N_5046,N_5841);
xor U6956 (N_6956,N_5611,N_5570);
nor U6957 (N_6957,N_5366,N_5680);
or U6958 (N_6958,N_5637,N_5889);
xor U6959 (N_6959,N_5798,N_5989);
or U6960 (N_6960,N_5783,N_5893);
nand U6961 (N_6961,N_5863,N_5906);
nor U6962 (N_6962,N_5907,N_5591);
nand U6963 (N_6963,N_5400,N_5940);
nor U6964 (N_6964,N_5132,N_5997);
nor U6965 (N_6965,N_5621,N_5144);
and U6966 (N_6966,N_5725,N_5315);
or U6967 (N_6967,N_5089,N_5162);
xor U6968 (N_6968,N_5697,N_5144);
and U6969 (N_6969,N_5829,N_5537);
nand U6970 (N_6970,N_5452,N_5154);
and U6971 (N_6971,N_5877,N_5811);
and U6972 (N_6972,N_5501,N_5733);
nor U6973 (N_6973,N_5520,N_5921);
xor U6974 (N_6974,N_5997,N_5759);
or U6975 (N_6975,N_5307,N_5370);
nand U6976 (N_6976,N_5072,N_5025);
nand U6977 (N_6977,N_5400,N_5771);
xnor U6978 (N_6978,N_5162,N_5764);
and U6979 (N_6979,N_5125,N_5647);
nand U6980 (N_6980,N_5531,N_5386);
nor U6981 (N_6981,N_5656,N_5302);
nand U6982 (N_6982,N_5876,N_5192);
xor U6983 (N_6983,N_5124,N_5611);
xnor U6984 (N_6984,N_5930,N_5293);
xor U6985 (N_6985,N_5240,N_5844);
or U6986 (N_6986,N_5613,N_5082);
nand U6987 (N_6987,N_5449,N_5819);
nor U6988 (N_6988,N_5791,N_5167);
nand U6989 (N_6989,N_5848,N_5315);
xor U6990 (N_6990,N_5656,N_5459);
xnor U6991 (N_6991,N_5738,N_5028);
nor U6992 (N_6992,N_5672,N_5545);
or U6993 (N_6993,N_5680,N_5552);
or U6994 (N_6994,N_5901,N_5872);
and U6995 (N_6995,N_5656,N_5146);
nand U6996 (N_6996,N_5523,N_5941);
xnor U6997 (N_6997,N_5063,N_5552);
or U6998 (N_6998,N_5270,N_5642);
nand U6999 (N_6999,N_5858,N_5138);
nand U7000 (N_7000,N_6738,N_6274);
and U7001 (N_7001,N_6138,N_6090);
nand U7002 (N_7002,N_6316,N_6523);
and U7003 (N_7003,N_6172,N_6204);
nor U7004 (N_7004,N_6192,N_6552);
or U7005 (N_7005,N_6355,N_6254);
and U7006 (N_7006,N_6685,N_6174);
or U7007 (N_7007,N_6111,N_6021);
nor U7008 (N_7008,N_6703,N_6640);
nor U7009 (N_7009,N_6647,N_6811);
or U7010 (N_7010,N_6026,N_6371);
or U7011 (N_7011,N_6938,N_6345);
or U7012 (N_7012,N_6566,N_6203);
or U7013 (N_7013,N_6067,N_6814);
or U7014 (N_7014,N_6144,N_6844);
nor U7015 (N_7015,N_6549,N_6619);
nand U7016 (N_7016,N_6957,N_6550);
xnor U7017 (N_7017,N_6396,N_6408);
and U7018 (N_7018,N_6893,N_6568);
nor U7019 (N_7019,N_6229,N_6792);
and U7020 (N_7020,N_6770,N_6939);
nand U7021 (N_7021,N_6728,N_6098);
nand U7022 (N_7022,N_6522,N_6638);
nand U7023 (N_7023,N_6535,N_6635);
nand U7024 (N_7024,N_6029,N_6722);
xor U7025 (N_7025,N_6973,N_6841);
or U7026 (N_7026,N_6056,N_6520);
nor U7027 (N_7027,N_6285,N_6187);
nand U7028 (N_7028,N_6199,N_6795);
nand U7029 (N_7029,N_6305,N_6912);
nand U7030 (N_7030,N_6579,N_6014);
nand U7031 (N_7031,N_6166,N_6981);
nor U7032 (N_7032,N_6262,N_6495);
or U7033 (N_7033,N_6244,N_6452);
nand U7034 (N_7034,N_6626,N_6235);
nand U7035 (N_7035,N_6819,N_6857);
and U7036 (N_7036,N_6466,N_6931);
nor U7037 (N_7037,N_6242,N_6188);
or U7038 (N_7038,N_6175,N_6654);
or U7039 (N_7039,N_6443,N_6010);
nor U7040 (N_7040,N_6313,N_6221);
xnor U7041 (N_7041,N_6460,N_6983);
or U7042 (N_7042,N_6093,N_6817);
or U7043 (N_7043,N_6249,N_6212);
xor U7044 (N_7044,N_6965,N_6444);
nor U7045 (N_7045,N_6789,N_6941);
or U7046 (N_7046,N_6489,N_6168);
xor U7047 (N_7047,N_6480,N_6830);
nand U7048 (N_7048,N_6483,N_6406);
nor U7049 (N_7049,N_6195,N_6031);
nor U7050 (N_7050,N_6639,N_6704);
or U7051 (N_7051,N_6159,N_6349);
or U7052 (N_7052,N_6757,N_6446);
and U7053 (N_7053,N_6864,N_6760);
nor U7054 (N_7054,N_6504,N_6456);
nor U7055 (N_7055,N_6266,N_6820);
nor U7056 (N_7056,N_6362,N_6911);
or U7057 (N_7057,N_6851,N_6954);
nand U7058 (N_7058,N_6512,N_6106);
and U7059 (N_7059,N_6945,N_6694);
xor U7060 (N_7060,N_6332,N_6592);
nand U7061 (N_7061,N_6241,N_6643);
or U7062 (N_7062,N_6538,N_6384);
and U7063 (N_7063,N_6264,N_6899);
nand U7064 (N_7064,N_6440,N_6590);
and U7065 (N_7065,N_6875,N_6907);
nand U7066 (N_7066,N_6220,N_6367);
and U7067 (N_7067,N_6651,N_6263);
nor U7068 (N_7068,N_6824,N_6223);
xor U7069 (N_7069,N_6877,N_6622);
xnor U7070 (N_7070,N_6471,N_6633);
xor U7071 (N_7071,N_6149,N_6683);
nand U7072 (N_7072,N_6324,N_6730);
or U7073 (N_7073,N_6154,N_6702);
or U7074 (N_7074,N_6729,N_6066);
nand U7075 (N_7075,N_6200,N_6075);
xnor U7076 (N_7076,N_6255,N_6748);
and U7077 (N_7077,N_6381,N_6074);
xor U7078 (N_7078,N_6554,N_6339);
xnor U7079 (N_7079,N_6663,N_6755);
or U7080 (N_7080,N_6561,N_6602);
and U7081 (N_7081,N_6900,N_6562);
nor U7082 (N_7082,N_6445,N_6454);
or U7083 (N_7083,N_6859,N_6065);
and U7084 (N_7084,N_6534,N_6777);
or U7085 (N_7085,N_6427,N_6231);
and U7086 (N_7086,N_6846,N_6426);
nand U7087 (N_7087,N_6048,N_6832);
and U7088 (N_7088,N_6948,N_6675);
nand U7089 (N_7089,N_6542,N_6351);
nor U7090 (N_7090,N_6723,N_6013);
nor U7091 (N_7091,N_6419,N_6287);
or U7092 (N_7092,N_6118,N_6334);
xnor U7093 (N_7093,N_6247,N_6173);
nor U7094 (N_7094,N_6314,N_6799);
nand U7095 (N_7095,N_6767,N_6039);
nor U7096 (N_7096,N_6448,N_6320);
or U7097 (N_7097,N_6769,N_6024);
xnor U7098 (N_7098,N_6887,N_6046);
nor U7099 (N_7099,N_6020,N_6055);
nand U7100 (N_7100,N_6493,N_6879);
nor U7101 (N_7101,N_6881,N_6089);
nand U7102 (N_7102,N_6398,N_6658);
xor U7103 (N_7103,N_6906,N_6257);
nand U7104 (N_7104,N_6671,N_6781);
or U7105 (N_7105,N_6719,N_6956);
nor U7106 (N_7106,N_6894,N_6077);
and U7107 (N_7107,N_6563,N_6272);
nand U7108 (N_7108,N_6226,N_6688);
nor U7109 (N_7109,N_6838,N_6937);
xor U7110 (N_7110,N_6128,N_6068);
or U7111 (N_7111,N_6153,N_6517);
and U7112 (N_7112,N_6301,N_6585);
nand U7113 (N_7113,N_6428,N_6499);
or U7114 (N_7114,N_6315,N_6978);
and U7115 (N_7115,N_6214,N_6528);
xnor U7116 (N_7116,N_6696,N_6509);
nor U7117 (N_7117,N_6155,N_6027);
and U7118 (N_7118,N_6752,N_6125);
nand U7119 (N_7119,N_6677,N_6641);
xor U7120 (N_7120,N_6136,N_6481);
xnor U7121 (N_7121,N_6082,N_6016);
xor U7122 (N_7122,N_6399,N_6225);
or U7123 (N_7123,N_6925,N_6525);
or U7124 (N_7124,N_6331,N_6724);
or U7125 (N_7125,N_6656,N_6710);
xor U7126 (N_7126,N_6474,N_6270);
or U7127 (N_7127,N_6599,N_6356);
or U7128 (N_7128,N_6197,N_6596);
and U7129 (N_7129,N_6835,N_6179);
and U7130 (N_7130,N_6213,N_6459);
nor U7131 (N_7131,N_6700,N_6547);
and U7132 (N_7132,N_6492,N_6400);
or U7133 (N_7133,N_6104,N_6442);
and U7134 (N_7134,N_6533,N_6441);
or U7135 (N_7135,N_6556,N_6980);
xor U7136 (N_7136,N_6224,N_6142);
xor U7137 (N_7137,N_6623,N_6910);
nand U7138 (N_7138,N_6580,N_6327);
and U7139 (N_7139,N_6787,N_6583);
xnor U7140 (N_7140,N_6934,N_6524);
nor U7141 (N_7141,N_6734,N_6006);
nor U7142 (N_7142,N_6123,N_6207);
nand U7143 (N_7143,N_6275,N_6030);
or U7144 (N_7144,N_6008,N_6145);
nor U7145 (N_7145,N_6099,N_6127);
or U7146 (N_7146,N_6932,N_6854);
nor U7147 (N_7147,N_6108,N_6572);
or U7148 (N_7148,N_6347,N_6727);
or U7149 (N_7149,N_6397,N_6189);
xor U7150 (N_7150,N_6181,N_6880);
xnor U7151 (N_7151,N_6836,N_6253);
xor U7152 (N_7152,N_6490,N_6037);
or U7153 (N_7153,N_6823,N_6196);
or U7154 (N_7154,N_6482,N_6372);
xor U7155 (N_7155,N_6968,N_6236);
and U7156 (N_7156,N_6141,N_6182);
or U7157 (N_7157,N_6551,N_6309);
xnor U7158 (N_7158,N_6791,N_6160);
nand U7159 (N_7159,N_6126,N_6896);
xnor U7160 (N_7160,N_6348,N_6260);
nand U7161 (N_7161,N_6465,N_6299);
nor U7162 (N_7162,N_6903,N_6344);
xnor U7163 (N_7163,N_6855,N_6637);
or U7164 (N_7164,N_6432,N_6073);
nand U7165 (N_7165,N_6989,N_6165);
nor U7166 (N_7166,N_6712,N_6373);
nand U7167 (N_7167,N_6059,N_6438);
nand U7168 (N_7168,N_6582,N_6737);
and U7169 (N_7169,N_6018,N_6005);
or U7170 (N_7170,N_6361,N_6497);
or U7171 (N_7171,N_6624,N_6537);
xor U7172 (N_7172,N_6988,N_6668);
xor U7173 (N_7173,N_6079,N_6813);
and U7174 (N_7174,N_6674,N_6962);
or U7175 (N_7175,N_6087,N_6085);
and U7176 (N_7176,N_6918,N_6601);
nand U7177 (N_7177,N_6574,N_6237);
xor U7178 (N_7178,N_6276,N_6783);
or U7179 (N_7179,N_6714,N_6377);
nor U7180 (N_7180,N_6358,N_6570);
or U7181 (N_7181,N_6246,N_6084);
and U7182 (N_7182,N_6395,N_6913);
or U7183 (N_7183,N_6464,N_6022);
xor U7184 (N_7184,N_6183,N_6115);
nand U7185 (N_7185,N_6457,N_6659);
and U7186 (N_7186,N_6884,N_6972);
and U7187 (N_7187,N_6686,N_6749);
or U7188 (N_7188,N_6888,N_6232);
and U7189 (N_7189,N_6975,N_6088);
or U7190 (N_7190,N_6271,N_6340);
or U7191 (N_7191,N_6634,N_6889);
or U7192 (N_7192,N_6215,N_6424);
nor U7193 (N_7193,N_6869,N_6023);
nor U7194 (N_7194,N_6532,N_6914);
nand U7195 (N_7195,N_6387,N_6919);
xor U7196 (N_7196,N_6451,N_6019);
nand U7197 (N_7197,N_6655,N_6506);
and U7198 (N_7198,N_6773,N_6935);
and U7199 (N_7199,N_6721,N_6076);
and U7200 (N_7200,N_6336,N_6302);
and U7201 (N_7201,N_6664,N_6167);
and U7202 (N_7202,N_6286,N_6025);
or U7203 (N_7203,N_6430,N_6343);
xnor U7204 (N_7204,N_6810,N_6614);
or U7205 (N_7205,N_6709,N_6708);
xnor U7206 (N_7206,N_6186,N_6051);
xor U7207 (N_7207,N_6868,N_6007);
nand U7208 (N_7208,N_6389,N_6184);
nor U7209 (N_7209,N_6961,N_6540);
or U7210 (N_7210,N_6856,N_6742);
nand U7211 (N_7211,N_6958,N_6776);
nor U7212 (N_7212,N_6329,N_6682);
and U7213 (N_7213,N_6133,N_6094);
or U7214 (N_7214,N_6064,N_6629);
nor U7215 (N_7215,N_6543,N_6248);
or U7216 (N_7216,N_6002,N_6421);
nand U7217 (N_7217,N_6797,N_6758);
nor U7218 (N_7218,N_6891,N_6964);
or U7219 (N_7219,N_6494,N_6303);
xor U7220 (N_7220,N_6132,N_6233);
nand U7221 (N_7221,N_6735,N_6843);
nand U7222 (N_7222,N_6822,N_6625);
and U7223 (N_7223,N_6711,N_6297);
or U7224 (N_7224,N_6407,N_6670);
and U7225 (N_7225,N_6743,N_6342);
nand U7226 (N_7226,N_6805,N_6564);
or U7227 (N_7227,N_6417,N_6439);
or U7228 (N_7228,N_6134,N_6825);
or U7229 (N_7229,N_6121,N_6762);
nand U7230 (N_7230,N_6850,N_6852);
nand U7231 (N_7231,N_6839,N_6295);
nand U7232 (N_7232,N_6573,N_6279);
or U7233 (N_7233,N_6505,N_6586);
and U7234 (N_7234,N_6120,N_6541);
and U7235 (N_7235,N_6992,N_6650);
nand U7236 (N_7236,N_6565,N_6611);
xor U7237 (N_7237,N_6933,N_6359);
nor U7238 (N_7238,N_6597,N_6994);
nand U7239 (N_7239,N_6034,N_6593);
xnor U7240 (N_7240,N_6536,N_6618);
nor U7241 (N_7241,N_6282,N_6936);
or U7242 (N_7242,N_6256,N_6208);
nand U7243 (N_7243,N_6831,N_6669);
nand U7244 (N_7244,N_6058,N_6865);
or U7245 (N_7245,N_6458,N_6273);
nand U7246 (N_7246,N_6943,N_6673);
xor U7247 (N_7247,N_6812,N_6576);
nor U7248 (N_7248,N_6969,N_6882);
nand U7249 (N_7249,N_6692,N_6672);
and U7250 (N_7250,N_6162,N_6388);
nand U7251 (N_7251,N_6240,N_6152);
nand U7252 (N_7252,N_6405,N_6291);
nor U7253 (N_7253,N_6050,N_6069);
or U7254 (N_7254,N_6953,N_6928);
xnor U7255 (N_7255,N_6418,N_6578);
xor U7256 (N_7256,N_6326,N_6904);
nor U7257 (N_7257,N_6521,N_6927);
nor U7258 (N_7258,N_6690,N_6415);
or U7259 (N_7259,N_6995,N_6527);
or U7260 (N_7260,N_6569,N_6720);
nand U7261 (N_7261,N_6496,N_6425);
nor U7262 (N_7262,N_6170,N_6277);
and U7263 (N_7263,N_6804,N_6778);
or U7264 (N_7264,N_6951,N_6739);
and U7265 (N_7265,N_6837,N_6821);
and U7266 (N_7266,N_6292,N_6060);
and U7267 (N_7267,N_6860,N_6131);
nor U7268 (N_7268,N_6849,N_6258);
xor U7269 (N_7269,N_6678,N_6621);
nand U7270 (N_7270,N_6984,N_6510);
nand U7271 (N_7271,N_6000,N_6293);
xor U7272 (N_7272,N_6594,N_6756);
or U7273 (N_7273,N_6402,N_6967);
nor U7274 (N_7274,N_6947,N_6311);
nor U7275 (N_7275,N_6986,N_6103);
and U7276 (N_7276,N_6699,N_6798);
nor U7277 (N_7277,N_6871,N_6976);
nand U7278 (N_7278,N_6015,N_6436);
nor U7279 (N_7279,N_6977,N_6139);
nor U7280 (N_7280,N_6267,N_6507);
nand U7281 (N_7281,N_6487,N_6210);
or U7282 (N_7282,N_6095,N_6401);
or U7283 (N_7283,N_6230,N_6319);
nor U7284 (N_7284,N_6486,N_6895);
nor U7285 (N_7285,N_6243,N_6431);
nand U7286 (N_7286,N_6705,N_6876);
and U7287 (N_7287,N_6449,N_6265);
xnor U7288 (N_7288,N_6807,N_6475);
nor U7289 (N_7289,N_6478,N_6312);
nor U7290 (N_7290,N_6909,N_6940);
xnor U7291 (N_7291,N_6886,N_6999);
or U7292 (N_7292,N_6330,N_6216);
nand U7293 (N_7293,N_6294,N_6238);
and U7294 (N_7294,N_6740,N_6392);
and U7295 (N_7295,N_6222,N_6963);
xor U7296 (N_7296,N_6930,N_6413);
xnor U7297 (N_7297,N_6818,N_6245);
nor U7298 (N_7298,N_6269,N_6515);
nor U7299 (N_7299,N_6915,N_6502);
nor U7300 (N_7300,N_6130,N_6544);
or U7301 (N_7301,N_6679,N_6878);
xnor U7302 (N_7302,N_6078,N_6178);
xnor U7303 (N_7303,N_6529,N_6600);
or U7304 (N_7304,N_6001,N_6357);
nand U7305 (N_7305,N_6109,N_6768);
or U7306 (N_7306,N_6902,N_6143);
nand U7307 (N_7307,N_6375,N_6217);
nor U7308 (N_7308,N_6318,N_6982);
xnor U7309 (N_7309,N_6741,N_6605);
nand U7310 (N_7310,N_6463,N_6146);
nand U7311 (N_7311,N_6433,N_6530);
nor U7312 (N_7312,N_6288,N_6322);
nor U7313 (N_7313,N_6630,N_6416);
nor U7314 (N_7314,N_6300,N_6386);
and U7315 (N_7315,N_6393,N_6833);
nor U7316 (N_7316,N_6110,N_6800);
xnor U7317 (N_7317,N_6991,N_6648);
nand U7318 (N_7318,N_6205,N_6555);
xor U7319 (N_7319,N_6861,N_6194);
nor U7320 (N_7320,N_6575,N_6137);
nand U7321 (N_7321,N_6571,N_6717);
nand U7322 (N_7322,N_6017,N_6979);
xnor U7323 (N_7323,N_6866,N_6012);
or U7324 (N_7324,N_6996,N_6041);
nor U7325 (N_7325,N_6676,N_6353);
or U7326 (N_7326,N_6853,N_6140);
xnor U7327 (N_7327,N_6598,N_6628);
or U7328 (N_7328,N_6049,N_6774);
nor U7329 (N_7329,N_6645,N_6086);
or U7330 (N_7330,N_6863,N_6306);
and U7331 (N_7331,N_6100,N_6746);
xor U7332 (N_7332,N_6870,N_6113);
xnor U7333 (N_7333,N_6105,N_6751);
xnor U7334 (N_7334,N_6701,N_6054);
nor U7335 (N_7335,N_6011,N_6158);
nand U7336 (N_7336,N_6698,N_6403);
or U7337 (N_7337,N_6045,N_6202);
nand U7338 (N_7338,N_6198,N_6206);
or U7339 (N_7339,N_6642,N_6560);
and U7340 (N_7340,N_6040,N_6595);
xnor U7341 (N_7341,N_6503,N_6558);
and U7342 (N_7342,N_6063,N_6157);
and U7343 (N_7343,N_6009,N_6514);
and U7344 (N_7344,N_6666,N_6083);
or U7345 (N_7345,N_6747,N_6809);
nor U7346 (N_7346,N_6364,N_6298);
nor U7347 (N_7347,N_6112,N_6061);
nor U7348 (N_7348,N_6290,N_6376);
xnor U7349 (N_7349,N_6379,N_6107);
and U7350 (N_7350,N_6693,N_6135);
or U7351 (N_7351,N_6070,N_6352);
or U7352 (N_7352,N_6097,N_6610);
xor U7353 (N_7353,N_6374,N_6631);
nor U7354 (N_7354,N_6434,N_6488);
nand U7355 (N_7355,N_6885,N_6122);
nor U7356 (N_7356,N_6032,N_6924);
xor U7357 (N_7357,N_6259,N_6296);
nand U7358 (N_7358,N_6508,N_6250);
or U7359 (N_7359,N_6588,N_6950);
nand U7360 (N_7360,N_6239,N_6763);
nor U7361 (N_7361,N_6307,N_6794);
or U7362 (N_7362,N_6462,N_6905);
and U7363 (N_7363,N_6604,N_6472);
and U7364 (N_7364,N_6808,N_6848);
nand U7365 (N_7365,N_6518,N_6929);
nand U7366 (N_7366,N_6971,N_6081);
nand U7367 (N_7367,N_6476,N_6771);
nor U7368 (N_7368,N_6917,N_6354);
nor U7369 (N_7369,N_6412,N_6053);
xnor U7370 (N_7370,N_6796,N_6447);
nor U7371 (N_7371,N_6491,N_6453);
nor U7372 (N_7372,N_6661,N_6479);
nor U7373 (N_7373,N_6072,N_6323);
xnor U7374 (N_7374,N_6959,N_6657);
or U7375 (N_7375,N_6176,N_6338);
nor U7376 (N_7376,N_6816,N_6680);
nand U7377 (N_7377,N_6922,N_6567);
xnor U7378 (N_7378,N_6872,N_6681);
or U7379 (N_7379,N_6461,N_6890);
and U7380 (N_7380,N_6731,N_6511);
nor U7381 (N_7381,N_6501,N_6341);
xor U7382 (N_7382,N_6469,N_6684);
xnor U7383 (N_7383,N_6845,N_6589);
and U7384 (N_7384,N_6378,N_6036);
nor U7385 (N_7385,N_6620,N_6328);
and U7386 (N_7386,N_6304,N_6793);
nor U7387 (N_7387,N_6840,N_6662);
xor U7388 (N_7388,N_6193,N_6513);
or U7389 (N_7389,N_6759,N_6119);
nor U7390 (N_7390,N_6500,N_6190);
nor U7391 (N_7391,N_6163,N_6960);
and U7392 (N_7392,N_6761,N_6004);
nor U7393 (N_7393,N_6993,N_6591);
and U7394 (N_7394,N_6057,N_6219);
nand U7395 (N_7395,N_6033,N_6707);
or U7396 (N_7396,N_6689,N_6784);
nand U7397 (N_7397,N_6873,N_6897);
and U7398 (N_7398,N_6091,N_6766);
nor U7399 (N_7399,N_6390,N_6827);
and U7400 (N_7400,N_6780,N_6468);
and U7401 (N_7401,N_6251,N_6252);
nor U7402 (N_7402,N_6786,N_6923);
nor U7403 (N_7403,N_6382,N_6608);
xor U7404 (N_7404,N_6612,N_6764);
or U7405 (N_7405,N_6990,N_6736);
nand U7406 (N_7406,N_6926,N_6636);
nor U7407 (N_7407,N_6801,N_6834);
nor U7408 (N_7408,N_6559,N_6949);
nor U7409 (N_7409,N_6955,N_6409);
nand U7410 (N_7410,N_6733,N_6035);
xnor U7411 (N_7411,N_6952,N_6627);
nor U7412 (N_7412,N_6394,N_6695);
and U7413 (N_7413,N_6970,N_6516);
or U7414 (N_7414,N_6450,N_6557);
nand U7415 (N_7415,N_6467,N_6308);
nor U7416 (N_7416,N_6102,N_6519);
nor U7417 (N_7417,N_6363,N_6209);
and U7418 (N_7418,N_6718,N_6360);
and U7419 (N_7419,N_6539,N_6148);
or U7420 (N_7420,N_6346,N_6646);
xor U7421 (N_7421,N_6171,N_6268);
nor U7422 (N_7422,N_6667,N_6003);
or U7423 (N_7423,N_6715,N_6691);
and U7424 (N_7424,N_6043,N_6716);
xnor U7425 (N_7425,N_6147,N_6211);
and U7426 (N_7426,N_6985,N_6803);
xor U7427 (N_7427,N_6942,N_6603);
nor U7428 (N_7428,N_6609,N_6584);
or U7429 (N_7429,N_6788,N_6410);
and U7430 (N_7430,N_6191,N_6745);
xor U7431 (N_7431,N_6124,N_6826);
and U7432 (N_7432,N_6096,N_6321);
nand U7433 (N_7433,N_6725,N_6867);
nor U7434 (N_7434,N_6847,N_6435);
or U7435 (N_7435,N_6802,N_6874);
or U7436 (N_7436,N_6422,N_6484);
or U7437 (N_7437,N_6317,N_6546);
xor U7438 (N_7438,N_6042,N_6782);
nor U7439 (N_7439,N_6883,N_6908);
nand U7440 (N_7440,N_6713,N_6790);
nand U7441 (N_7441,N_6744,N_6653);
and U7442 (N_7442,N_6587,N_6470);
nor U7443 (N_7443,N_6779,N_6151);
nand U7444 (N_7444,N_6177,N_6862);
and U7445 (N_7445,N_6335,N_6665);
nand U7446 (N_7446,N_6581,N_6129);
xnor U7447 (N_7447,N_6278,N_6946);
nor U7448 (N_7448,N_6649,N_6333);
xor U7449 (N_7449,N_6828,N_6898);
nor U7450 (N_7450,N_6485,N_6369);
and U7451 (N_7451,N_6772,N_6169);
nand U7452 (N_7452,N_6380,N_6892);
or U7453 (N_7453,N_6101,N_6944);
or U7454 (N_7454,N_6732,N_6185);
and U7455 (N_7455,N_6350,N_6545);
and U7456 (N_7456,N_6901,N_6644);
xnor U7457 (N_7457,N_6383,N_6385);
nor U7458 (N_7458,N_6161,N_6785);
xnor U7459 (N_7459,N_6281,N_6473);
nand U7460 (N_7460,N_6829,N_6365);
nor U7461 (N_7461,N_6310,N_6553);
nor U7462 (N_7462,N_6047,N_6150);
nor U7463 (N_7463,N_6411,N_6606);
and U7464 (N_7464,N_6815,N_6201);
nor U7465 (N_7465,N_6337,N_6164);
nor U7466 (N_7466,N_6726,N_6080);
nor U7467 (N_7467,N_6753,N_6404);
and U7468 (N_7468,N_6998,N_6156);
or U7469 (N_7469,N_6616,N_6613);
nor U7470 (N_7470,N_6577,N_6607);
nand U7471 (N_7471,N_6498,N_6754);
and U7472 (N_7472,N_6391,N_6966);
nand U7473 (N_7473,N_6234,N_6062);
nor U7474 (N_7474,N_6765,N_6660);
nor U7475 (N_7475,N_6280,N_6916);
xnor U7476 (N_7476,N_6044,N_6180);
nand U7477 (N_7477,N_6368,N_6052);
nand U7478 (N_7478,N_6218,N_6806);
nor U7479 (N_7479,N_6414,N_6261);
xor U7480 (N_7480,N_6289,N_6858);
xor U7481 (N_7481,N_6071,N_6437);
nor U7482 (N_7482,N_6632,N_6974);
or U7483 (N_7483,N_6548,N_6775);
nand U7484 (N_7484,N_6423,N_6652);
nand U7485 (N_7485,N_6227,N_6366);
or U7486 (N_7486,N_6092,N_6706);
xnor U7487 (N_7487,N_6750,N_6531);
nor U7488 (N_7488,N_6429,N_6325);
nor U7489 (N_7489,N_6028,N_6116);
and U7490 (N_7490,N_6687,N_6526);
nand U7491 (N_7491,N_6114,N_6117);
nand U7492 (N_7492,N_6842,N_6697);
and U7493 (N_7493,N_6997,N_6921);
and U7494 (N_7494,N_6370,N_6284);
and U7495 (N_7495,N_6617,N_6987);
and U7496 (N_7496,N_6038,N_6228);
and U7497 (N_7497,N_6477,N_6283);
and U7498 (N_7498,N_6615,N_6455);
nor U7499 (N_7499,N_6420,N_6920);
xnor U7500 (N_7500,N_6838,N_6080);
or U7501 (N_7501,N_6941,N_6801);
and U7502 (N_7502,N_6166,N_6372);
nand U7503 (N_7503,N_6385,N_6155);
xor U7504 (N_7504,N_6113,N_6381);
xor U7505 (N_7505,N_6811,N_6723);
xor U7506 (N_7506,N_6267,N_6757);
and U7507 (N_7507,N_6381,N_6030);
nand U7508 (N_7508,N_6349,N_6330);
and U7509 (N_7509,N_6949,N_6837);
nand U7510 (N_7510,N_6922,N_6069);
nor U7511 (N_7511,N_6320,N_6079);
or U7512 (N_7512,N_6402,N_6529);
nand U7513 (N_7513,N_6105,N_6461);
and U7514 (N_7514,N_6412,N_6761);
nand U7515 (N_7515,N_6897,N_6366);
nor U7516 (N_7516,N_6146,N_6290);
xor U7517 (N_7517,N_6451,N_6982);
nor U7518 (N_7518,N_6370,N_6552);
nor U7519 (N_7519,N_6922,N_6101);
and U7520 (N_7520,N_6956,N_6705);
or U7521 (N_7521,N_6133,N_6773);
nor U7522 (N_7522,N_6394,N_6469);
and U7523 (N_7523,N_6675,N_6150);
nand U7524 (N_7524,N_6681,N_6529);
xnor U7525 (N_7525,N_6840,N_6093);
or U7526 (N_7526,N_6810,N_6491);
nand U7527 (N_7527,N_6136,N_6538);
nor U7528 (N_7528,N_6529,N_6541);
nor U7529 (N_7529,N_6670,N_6695);
and U7530 (N_7530,N_6463,N_6440);
and U7531 (N_7531,N_6228,N_6913);
or U7532 (N_7532,N_6592,N_6112);
xnor U7533 (N_7533,N_6436,N_6988);
nor U7534 (N_7534,N_6007,N_6357);
or U7535 (N_7535,N_6534,N_6591);
xor U7536 (N_7536,N_6635,N_6092);
or U7537 (N_7537,N_6688,N_6967);
and U7538 (N_7538,N_6164,N_6166);
nand U7539 (N_7539,N_6612,N_6976);
and U7540 (N_7540,N_6496,N_6566);
xnor U7541 (N_7541,N_6439,N_6286);
nor U7542 (N_7542,N_6975,N_6056);
or U7543 (N_7543,N_6682,N_6930);
nand U7544 (N_7544,N_6483,N_6009);
or U7545 (N_7545,N_6212,N_6539);
or U7546 (N_7546,N_6104,N_6630);
or U7547 (N_7547,N_6484,N_6664);
xor U7548 (N_7548,N_6146,N_6232);
nor U7549 (N_7549,N_6833,N_6361);
or U7550 (N_7550,N_6797,N_6649);
or U7551 (N_7551,N_6783,N_6441);
nor U7552 (N_7552,N_6553,N_6924);
nand U7553 (N_7553,N_6863,N_6938);
nor U7554 (N_7554,N_6050,N_6857);
or U7555 (N_7555,N_6658,N_6104);
or U7556 (N_7556,N_6579,N_6979);
xor U7557 (N_7557,N_6213,N_6498);
or U7558 (N_7558,N_6450,N_6266);
nor U7559 (N_7559,N_6481,N_6355);
or U7560 (N_7560,N_6317,N_6195);
or U7561 (N_7561,N_6909,N_6359);
nor U7562 (N_7562,N_6773,N_6367);
or U7563 (N_7563,N_6716,N_6817);
nor U7564 (N_7564,N_6076,N_6712);
xnor U7565 (N_7565,N_6529,N_6771);
nor U7566 (N_7566,N_6904,N_6148);
or U7567 (N_7567,N_6226,N_6386);
or U7568 (N_7568,N_6886,N_6795);
xor U7569 (N_7569,N_6272,N_6334);
xor U7570 (N_7570,N_6877,N_6779);
nor U7571 (N_7571,N_6833,N_6548);
and U7572 (N_7572,N_6840,N_6561);
nand U7573 (N_7573,N_6774,N_6986);
or U7574 (N_7574,N_6342,N_6628);
nor U7575 (N_7575,N_6641,N_6369);
nand U7576 (N_7576,N_6145,N_6120);
nor U7577 (N_7577,N_6763,N_6076);
or U7578 (N_7578,N_6974,N_6888);
nor U7579 (N_7579,N_6017,N_6170);
nor U7580 (N_7580,N_6245,N_6516);
or U7581 (N_7581,N_6857,N_6840);
nor U7582 (N_7582,N_6383,N_6495);
or U7583 (N_7583,N_6476,N_6647);
xnor U7584 (N_7584,N_6792,N_6159);
xor U7585 (N_7585,N_6735,N_6123);
or U7586 (N_7586,N_6633,N_6934);
nor U7587 (N_7587,N_6251,N_6150);
and U7588 (N_7588,N_6556,N_6503);
or U7589 (N_7589,N_6994,N_6422);
and U7590 (N_7590,N_6987,N_6296);
and U7591 (N_7591,N_6137,N_6428);
and U7592 (N_7592,N_6592,N_6039);
or U7593 (N_7593,N_6866,N_6981);
xor U7594 (N_7594,N_6628,N_6900);
nand U7595 (N_7595,N_6869,N_6484);
xnor U7596 (N_7596,N_6588,N_6016);
nand U7597 (N_7597,N_6286,N_6376);
and U7598 (N_7598,N_6380,N_6047);
xnor U7599 (N_7599,N_6484,N_6001);
and U7600 (N_7600,N_6881,N_6680);
or U7601 (N_7601,N_6530,N_6010);
nor U7602 (N_7602,N_6906,N_6747);
nor U7603 (N_7603,N_6849,N_6282);
nor U7604 (N_7604,N_6817,N_6196);
and U7605 (N_7605,N_6726,N_6816);
or U7606 (N_7606,N_6265,N_6588);
or U7607 (N_7607,N_6666,N_6301);
and U7608 (N_7608,N_6786,N_6828);
nand U7609 (N_7609,N_6890,N_6388);
nand U7610 (N_7610,N_6645,N_6363);
nor U7611 (N_7611,N_6086,N_6466);
nor U7612 (N_7612,N_6619,N_6477);
xnor U7613 (N_7613,N_6130,N_6899);
xnor U7614 (N_7614,N_6401,N_6806);
or U7615 (N_7615,N_6669,N_6438);
nor U7616 (N_7616,N_6371,N_6714);
and U7617 (N_7617,N_6632,N_6729);
nand U7618 (N_7618,N_6043,N_6618);
or U7619 (N_7619,N_6143,N_6701);
nor U7620 (N_7620,N_6199,N_6904);
and U7621 (N_7621,N_6507,N_6099);
xor U7622 (N_7622,N_6541,N_6478);
or U7623 (N_7623,N_6316,N_6804);
nor U7624 (N_7624,N_6224,N_6031);
and U7625 (N_7625,N_6268,N_6936);
or U7626 (N_7626,N_6894,N_6091);
and U7627 (N_7627,N_6937,N_6490);
xnor U7628 (N_7628,N_6402,N_6835);
xnor U7629 (N_7629,N_6658,N_6056);
or U7630 (N_7630,N_6569,N_6606);
and U7631 (N_7631,N_6211,N_6322);
and U7632 (N_7632,N_6972,N_6332);
or U7633 (N_7633,N_6662,N_6465);
nand U7634 (N_7634,N_6377,N_6057);
nand U7635 (N_7635,N_6450,N_6563);
nor U7636 (N_7636,N_6267,N_6599);
xor U7637 (N_7637,N_6622,N_6526);
or U7638 (N_7638,N_6248,N_6542);
or U7639 (N_7639,N_6609,N_6305);
nand U7640 (N_7640,N_6637,N_6117);
or U7641 (N_7641,N_6167,N_6721);
nand U7642 (N_7642,N_6911,N_6904);
nand U7643 (N_7643,N_6297,N_6284);
and U7644 (N_7644,N_6688,N_6333);
xnor U7645 (N_7645,N_6083,N_6703);
nand U7646 (N_7646,N_6513,N_6248);
nor U7647 (N_7647,N_6645,N_6470);
and U7648 (N_7648,N_6575,N_6207);
xnor U7649 (N_7649,N_6003,N_6053);
or U7650 (N_7650,N_6078,N_6779);
nor U7651 (N_7651,N_6672,N_6224);
nor U7652 (N_7652,N_6837,N_6261);
xnor U7653 (N_7653,N_6501,N_6683);
nand U7654 (N_7654,N_6071,N_6760);
nor U7655 (N_7655,N_6668,N_6746);
and U7656 (N_7656,N_6283,N_6063);
and U7657 (N_7657,N_6116,N_6520);
or U7658 (N_7658,N_6396,N_6031);
xnor U7659 (N_7659,N_6059,N_6443);
and U7660 (N_7660,N_6299,N_6757);
or U7661 (N_7661,N_6529,N_6483);
nand U7662 (N_7662,N_6345,N_6868);
or U7663 (N_7663,N_6292,N_6121);
or U7664 (N_7664,N_6316,N_6958);
xor U7665 (N_7665,N_6766,N_6460);
nand U7666 (N_7666,N_6312,N_6790);
xnor U7667 (N_7667,N_6607,N_6902);
nor U7668 (N_7668,N_6295,N_6694);
and U7669 (N_7669,N_6148,N_6134);
nor U7670 (N_7670,N_6736,N_6583);
or U7671 (N_7671,N_6231,N_6880);
nor U7672 (N_7672,N_6898,N_6637);
and U7673 (N_7673,N_6871,N_6102);
xnor U7674 (N_7674,N_6782,N_6652);
nor U7675 (N_7675,N_6789,N_6807);
and U7676 (N_7676,N_6163,N_6265);
nand U7677 (N_7677,N_6369,N_6002);
nand U7678 (N_7678,N_6481,N_6822);
and U7679 (N_7679,N_6845,N_6286);
and U7680 (N_7680,N_6367,N_6248);
nor U7681 (N_7681,N_6886,N_6979);
xor U7682 (N_7682,N_6299,N_6053);
xor U7683 (N_7683,N_6623,N_6861);
and U7684 (N_7684,N_6765,N_6320);
nand U7685 (N_7685,N_6216,N_6156);
xnor U7686 (N_7686,N_6177,N_6024);
or U7687 (N_7687,N_6866,N_6129);
or U7688 (N_7688,N_6141,N_6970);
nand U7689 (N_7689,N_6926,N_6630);
xor U7690 (N_7690,N_6124,N_6298);
and U7691 (N_7691,N_6176,N_6179);
nor U7692 (N_7692,N_6787,N_6392);
and U7693 (N_7693,N_6019,N_6086);
nor U7694 (N_7694,N_6429,N_6232);
or U7695 (N_7695,N_6160,N_6789);
xor U7696 (N_7696,N_6431,N_6498);
and U7697 (N_7697,N_6008,N_6398);
xnor U7698 (N_7698,N_6629,N_6613);
nand U7699 (N_7699,N_6458,N_6812);
or U7700 (N_7700,N_6471,N_6222);
or U7701 (N_7701,N_6990,N_6711);
nor U7702 (N_7702,N_6875,N_6612);
or U7703 (N_7703,N_6208,N_6438);
xnor U7704 (N_7704,N_6290,N_6680);
or U7705 (N_7705,N_6689,N_6375);
nor U7706 (N_7706,N_6386,N_6304);
xor U7707 (N_7707,N_6777,N_6753);
or U7708 (N_7708,N_6882,N_6442);
xnor U7709 (N_7709,N_6073,N_6566);
nor U7710 (N_7710,N_6487,N_6301);
nor U7711 (N_7711,N_6237,N_6354);
nor U7712 (N_7712,N_6935,N_6739);
nand U7713 (N_7713,N_6752,N_6568);
xnor U7714 (N_7714,N_6578,N_6180);
nor U7715 (N_7715,N_6581,N_6394);
and U7716 (N_7716,N_6149,N_6182);
nand U7717 (N_7717,N_6992,N_6360);
and U7718 (N_7718,N_6446,N_6782);
xor U7719 (N_7719,N_6249,N_6986);
and U7720 (N_7720,N_6519,N_6845);
xnor U7721 (N_7721,N_6856,N_6863);
and U7722 (N_7722,N_6512,N_6480);
nand U7723 (N_7723,N_6993,N_6077);
and U7724 (N_7724,N_6989,N_6939);
nor U7725 (N_7725,N_6873,N_6194);
xnor U7726 (N_7726,N_6850,N_6483);
nor U7727 (N_7727,N_6804,N_6631);
xnor U7728 (N_7728,N_6371,N_6891);
or U7729 (N_7729,N_6010,N_6277);
nor U7730 (N_7730,N_6014,N_6959);
or U7731 (N_7731,N_6221,N_6584);
xor U7732 (N_7732,N_6891,N_6467);
and U7733 (N_7733,N_6776,N_6610);
or U7734 (N_7734,N_6822,N_6679);
or U7735 (N_7735,N_6719,N_6414);
nand U7736 (N_7736,N_6507,N_6310);
nand U7737 (N_7737,N_6750,N_6644);
nor U7738 (N_7738,N_6028,N_6258);
nor U7739 (N_7739,N_6527,N_6970);
xnor U7740 (N_7740,N_6818,N_6375);
nand U7741 (N_7741,N_6084,N_6591);
nand U7742 (N_7742,N_6174,N_6192);
nand U7743 (N_7743,N_6114,N_6128);
and U7744 (N_7744,N_6062,N_6378);
or U7745 (N_7745,N_6004,N_6765);
or U7746 (N_7746,N_6206,N_6390);
xor U7747 (N_7747,N_6941,N_6293);
or U7748 (N_7748,N_6504,N_6111);
nand U7749 (N_7749,N_6070,N_6019);
and U7750 (N_7750,N_6802,N_6073);
or U7751 (N_7751,N_6549,N_6586);
nand U7752 (N_7752,N_6230,N_6336);
xor U7753 (N_7753,N_6776,N_6104);
nand U7754 (N_7754,N_6428,N_6127);
and U7755 (N_7755,N_6767,N_6022);
xnor U7756 (N_7756,N_6326,N_6339);
or U7757 (N_7757,N_6306,N_6552);
and U7758 (N_7758,N_6080,N_6277);
nand U7759 (N_7759,N_6483,N_6729);
nor U7760 (N_7760,N_6433,N_6289);
and U7761 (N_7761,N_6480,N_6280);
or U7762 (N_7762,N_6305,N_6667);
or U7763 (N_7763,N_6530,N_6979);
nand U7764 (N_7764,N_6912,N_6913);
nand U7765 (N_7765,N_6820,N_6236);
nand U7766 (N_7766,N_6434,N_6184);
nand U7767 (N_7767,N_6829,N_6029);
nor U7768 (N_7768,N_6555,N_6417);
nor U7769 (N_7769,N_6093,N_6189);
or U7770 (N_7770,N_6500,N_6736);
nor U7771 (N_7771,N_6231,N_6615);
nor U7772 (N_7772,N_6796,N_6840);
or U7773 (N_7773,N_6005,N_6028);
and U7774 (N_7774,N_6153,N_6333);
nor U7775 (N_7775,N_6269,N_6134);
xnor U7776 (N_7776,N_6278,N_6765);
and U7777 (N_7777,N_6670,N_6333);
xor U7778 (N_7778,N_6698,N_6521);
and U7779 (N_7779,N_6122,N_6250);
and U7780 (N_7780,N_6525,N_6848);
nand U7781 (N_7781,N_6057,N_6889);
or U7782 (N_7782,N_6294,N_6907);
and U7783 (N_7783,N_6262,N_6451);
nor U7784 (N_7784,N_6574,N_6948);
xor U7785 (N_7785,N_6950,N_6434);
nand U7786 (N_7786,N_6476,N_6561);
or U7787 (N_7787,N_6218,N_6196);
nand U7788 (N_7788,N_6176,N_6844);
nand U7789 (N_7789,N_6470,N_6859);
or U7790 (N_7790,N_6237,N_6780);
nand U7791 (N_7791,N_6231,N_6540);
or U7792 (N_7792,N_6516,N_6369);
xnor U7793 (N_7793,N_6903,N_6206);
nor U7794 (N_7794,N_6594,N_6507);
and U7795 (N_7795,N_6353,N_6115);
xnor U7796 (N_7796,N_6387,N_6717);
and U7797 (N_7797,N_6390,N_6744);
xor U7798 (N_7798,N_6581,N_6563);
or U7799 (N_7799,N_6426,N_6382);
or U7800 (N_7800,N_6741,N_6286);
and U7801 (N_7801,N_6463,N_6459);
or U7802 (N_7802,N_6891,N_6177);
nor U7803 (N_7803,N_6210,N_6749);
xor U7804 (N_7804,N_6848,N_6225);
or U7805 (N_7805,N_6150,N_6789);
nor U7806 (N_7806,N_6218,N_6922);
or U7807 (N_7807,N_6845,N_6488);
or U7808 (N_7808,N_6155,N_6619);
and U7809 (N_7809,N_6396,N_6180);
or U7810 (N_7810,N_6304,N_6296);
or U7811 (N_7811,N_6985,N_6412);
xnor U7812 (N_7812,N_6191,N_6305);
nand U7813 (N_7813,N_6557,N_6246);
or U7814 (N_7814,N_6194,N_6781);
or U7815 (N_7815,N_6068,N_6906);
nand U7816 (N_7816,N_6435,N_6084);
nor U7817 (N_7817,N_6702,N_6583);
and U7818 (N_7818,N_6557,N_6385);
or U7819 (N_7819,N_6497,N_6864);
and U7820 (N_7820,N_6437,N_6662);
nand U7821 (N_7821,N_6786,N_6216);
nor U7822 (N_7822,N_6568,N_6955);
nand U7823 (N_7823,N_6781,N_6892);
nor U7824 (N_7824,N_6587,N_6334);
nand U7825 (N_7825,N_6761,N_6087);
nor U7826 (N_7826,N_6237,N_6494);
or U7827 (N_7827,N_6470,N_6056);
or U7828 (N_7828,N_6291,N_6011);
nand U7829 (N_7829,N_6835,N_6532);
or U7830 (N_7830,N_6493,N_6946);
xnor U7831 (N_7831,N_6709,N_6618);
nor U7832 (N_7832,N_6449,N_6459);
xor U7833 (N_7833,N_6341,N_6553);
nor U7834 (N_7834,N_6405,N_6848);
or U7835 (N_7835,N_6079,N_6143);
nand U7836 (N_7836,N_6716,N_6275);
nand U7837 (N_7837,N_6891,N_6897);
and U7838 (N_7838,N_6613,N_6324);
or U7839 (N_7839,N_6327,N_6154);
xor U7840 (N_7840,N_6226,N_6371);
xnor U7841 (N_7841,N_6307,N_6929);
nor U7842 (N_7842,N_6207,N_6372);
or U7843 (N_7843,N_6494,N_6351);
xor U7844 (N_7844,N_6703,N_6078);
or U7845 (N_7845,N_6314,N_6838);
or U7846 (N_7846,N_6025,N_6296);
nand U7847 (N_7847,N_6967,N_6766);
nand U7848 (N_7848,N_6703,N_6921);
or U7849 (N_7849,N_6305,N_6640);
or U7850 (N_7850,N_6541,N_6139);
xnor U7851 (N_7851,N_6070,N_6102);
nand U7852 (N_7852,N_6052,N_6791);
nor U7853 (N_7853,N_6880,N_6796);
nor U7854 (N_7854,N_6165,N_6592);
or U7855 (N_7855,N_6820,N_6847);
nand U7856 (N_7856,N_6232,N_6991);
and U7857 (N_7857,N_6182,N_6727);
nor U7858 (N_7858,N_6248,N_6577);
or U7859 (N_7859,N_6846,N_6576);
and U7860 (N_7860,N_6088,N_6307);
or U7861 (N_7861,N_6710,N_6387);
and U7862 (N_7862,N_6009,N_6473);
or U7863 (N_7863,N_6469,N_6319);
xnor U7864 (N_7864,N_6877,N_6149);
and U7865 (N_7865,N_6682,N_6271);
or U7866 (N_7866,N_6915,N_6520);
nor U7867 (N_7867,N_6445,N_6183);
or U7868 (N_7868,N_6714,N_6334);
nor U7869 (N_7869,N_6920,N_6520);
nor U7870 (N_7870,N_6957,N_6253);
nand U7871 (N_7871,N_6114,N_6943);
or U7872 (N_7872,N_6464,N_6770);
nand U7873 (N_7873,N_6008,N_6112);
or U7874 (N_7874,N_6717,N_6006);
xnor U7875 (N_7875,N_6806,N_6297);
xor U7876 (N_7876,N_6785,N_6808);
and U7877 (N_7877,N_6146,N_6476);
and U7878 (N_7878,N_6234,N_6422);
nand U7879 (N_7879,N_6431,N_6679);
xor U7880 (N_7880,N_6460,N_6690);
xor U7881 (N_7881,N_6533,N_6033);
nor U7882 (N_7882,N_6262,N_6321);
xnor U7883 (N_7883,N_6074,N_6434);
xnor U7884 (N_7884,N_6943,N_6583);
or U7885 (N_7885,N_6827,N_6124);
and U7886 (N_7886,N_6539,N_6193);
xor U7887 (N_7887,N_6265,N_6986);
xor U7888 (N_7888,N_6174,N_6680);
nand U7889 (N_7889,N_6957,N_6752);
and U7890 (N_7890,N_6521,N_6714);
or U7891 (N_7891,N_6146,N_6224);
xnor U7892 (N_7892,N_6649,N_6379);
nor U7893 (N_7893,N_6729,N_6623);
xor U7894 (N_7894,N_6231,N_6600);
xor U7895 (N_7895,N_6402,N_6314);
xnor U7896 (N_7896,N_6937,N_6085);
nor U7897 (N_7897,N_6150,N_6590);
and U7898 (N_7898,N_6748,N_6070);
xor U7899 (N_7899,N_6150,N_6331);
nand U7900 (N_7900,N_6311,N_6778);
or U7901 (N_7901,N_6703,N_6305);
and U7902 (N_7902,N_6740,N_6851);
and U7903 (N_7903,N_6415,N_6441);
xor U7904 (N_7904,N_6363,N_6056);
nor U7905 (N_7905,N_6808,N_6925);
nand U7906 (N_7906,N_6269,N_6165);
nor U7907 (N_7907,N_6214,N_6795);
and U7908 (N_7908,N_6924,N_6707);
and U7909 (N_7909,N_6698,N_6852);
nor U7910 (N_7910,N_6240,N_6416);
nand U7911 (N_7911,N_6284,N_6028);
and U7912 (N_7912,N_6255,N_6910);
xnor U7913 (N_7913,N_6530,N_6565);
or U7914 (N_7914,N_6521,N_6702);
and U7915 (N_7915,N_6932,N_6408);
or U7916 (N_7916,N_6065,N_6268);
nand U7917 (N_7917,N_6197,N_6100);
nand U7918 (N_7918,N_6228,N_6935);
or U7919 (N_7919,N_6129,N_6640);
xnor U7920 (N_7920,N_6166,N_6992);
nand U7921 (N_7921,N_6962,N_6509);
and U7922 (N_7922,N_6131,N_6395);
nand U7923 (N_7923,N_6575,N_6952);
or U7924 (N_7924,N_6887,N_6142);
nand U7925 (N_7925,N_6920,N_6822);
and U7926 (N_7926,N_6016,N_6180);
nor U7927 (N_7927,N_6333,N_6855);
nand U7928 (N_7928,N_6102,N_6729);
and U7929 (N_7929,N_6176,N_6489);
and U7930 (N_7930,N_6285,N_6997);
and U7931 (N_7931,N_6494,N_6657);
nor U7932 (N_7932,N_6010,N_6391);
nor U7933 (N_7933,N_6708,N_6198);
nand U7934 (N_7934,N_6588,N_6151);
or U7935 (N_7935,N_6766,N_6186);
or U7936 (N_7936,N_6679,N_6101);
nor U7937 (N_7937,N_6289,N_6287);
nor U7938 (N_7938,N_6798,N_6371);
or U7939 (N_7939,N_6845,N_6989);
or U7940 (N_7940,N_6270,N_6959);
nand U7941 (N_7941,N_6469,N_6785);
nand U7942 (N_7942,N_6033,N_6473);
or U7943 (N_7943,N_6516,N_6739);
nand U7944 (N_7944,N_6471,N_6256);
and U7945 (N_7945,N_6941,N_6772);
and U7946 (N_7946,N_6510,N_6212);
xnor U7947 (N_7947,N_6907,N_6278);
or U7948 (N_7948,N_6105,N_6189);
or U7949 (N_7949,N_6267,N_6544);
nand U7950 (N_7950,N_6574,N_6324);
or U7951 (N_7951,N_6489,N_6118);
or U7952 (N_7952,N_6214,N_6264);
nor U7953 (N_7953,N_6146,N_6821);
and U7954 (N_7954,N_6079,N_6005);
and U7955 (N_7955,N_6225,N_6568);
xnor U7956 (N_7956,N_6552,N_6502);
nand U7957 (N_7957,N_6254,N_6398);
nor U7958 (N_7958,N_6545,N_6929);
xnor U7959 (N_7959,N_6599,N_6008);
and U7960 (N_7960,N_6928,N_6423);
xnor U7961 (N_7961,N_6250,N_6307);
and U7962 (N_7962,N_6161,N_6535);
nor U7963 (N_7963,N_6397,N_6674);
or U7964 (N_7964,N_6219,N_6980);
nand U7965 (N_7965,N_6470,N_6272);
xnor U7966 (N_7966,N_6464,N_6766);
or U7967 (N_7967,N_6103,N_6502);
nor U7968 (N_7968,N_6423,N_6750);
and U7969 (N_7969,N_6526,N_6868);
nor U7970 (N_7970,N_6606,N_6152);
nor U7971 (N_7971,N_6050,N_6550);
nor U7972 (N_7972,N_6350,N_6600);
nor U7973 (N_7973,N_6565,N_6434);
nand U7974 (N_7974,N_6973,N_6430);
xor U7975 (N_7975,N_6684,N_6259);
or U7976 (N_7976,N_6403,N_6798);
or U7977 (N_7977,N_6926,N_6191);
or U7978 (N_7978,N_6595,N_6893);
and U7979 (N_7979,N_6136,N_6568);
or U7980 (N_7980,N_6086,N_6148);
xor U7981 (N_7981,N_6793,N_6651);
xnor U7982 (N_7982,N_6343,N_6934);
nand U7983 (N_7983,N_6843,N_6145);
or U7984 (N_7984,N_6338,N_6242);
nor U7985 (N_7985,N_6967,N_6755);
or U7986 (N_7986,N_6421,N_6780);
or U7987 (N_7987,N_6179,N_6884);
and U7988 (N_7988,N_6487,N_6641);
and U7989 (N_7989,N_6219,N_6340);
nand U7990 (N_7990,N_6950,N_6526);
and U7991 (N_7991,N_6973,N_6659);
or U7992 (N_7992,N_6036,N_6484);
nor U7993 (N_7993,N_6269,N_6585);
nand U7994 (N_7994,N_6717,N_6611);
and U7995 (N_7995,N_6709,N_6484);
and U7996 (N_7996,N_6808,N_6772);
nor U7997 (N_7997,N_6326,N_6062);
or U7998 (N_7998,N_6373,N_6729);
nor U7999 (N_7999,N_6890,N_6834);
xnor U8000 (N_8000,N_7347,N_7868);
and U8001 (N_8001,N_7070,N_7394);
and U8002 (N_8002,N_7950,N_7917);
or U8003 (N_8003,N_7874,N_7283);
or U8004 (N_8004,N_7136,N_7991);
xor U8005 (N_8005,N_7530,N_7822);
or U8006 (N_8006,N_7816,N_7527);
xnor U8007 (N_8007,N_7463,N_7230);
nor U8008 (N_8008,N_7037,N_7248);
xnor U8009 (N_8009,N_7867,N_7449);
and U8010 (N_8010,N_7190,N_7340);
nand U8011 (N_8011,N_7054,N_7817);
nor U8012 (N_8012,N_7495,N_7351);
xnor U8013 (N_8013,N_7523,N_7643);
or U8014 (N_8014,N_7303,N_7943);
and U8015 (N_8015,N_7119,N_7003);
and U8016 (N_8016,N_7737,N_7494);
nor U8017 (N_8017,N_7490,N_7338);
and U8018 (N_8018,N_7468,N_7242);
nor U8019 (N_8019,N_7424,N_7327);
and U8020 (N_8020,N_7906,N_7751);
nand U8021 (N_8021,N_7672,N_7369);
nand U8022 (N_8022,N_7216,N_7529);
nand U8023 (N_8023,N_7464,N_7202);
or U8024 (N_8024,N_7035,N_7728);
or U8025 (N_8025,N_7115,N_7844);
xor U8026 (N_8026,N_7189,N_7050);
or U8027 (N_8027,N_7741,N_7573);
nand U8028 (N_8028,N_7286,N_7325);
nor U8029 (N_8029,N_7184,N_7368);
nand U8030 (N_8030,N_7264,N_7241);
or U8031 (N_8031,N_7379,N_7632);
or U8032 (N_8032,N_7461,N_7767);
or U8033 (N_8033,N_7235,N_7363);
or U8034 (N_8034,N_7251,N_7642);
xor U8035 (N_8035,N_7063,N_7373);
xor U8036 (N_8036,N_7160,N_7743);
xnor U8037 (N_8037,N_7467,N_7598);
and U8038 (N_8038,N_7181,N_7945);
nand U8039 (N_8039,N_7295,N_7634);
nand U8040 (N_8040,N_7317,N_7278);
xnor U8041 (N_8041,N_7339,N_7756);
xnor U8042 (N_8042,N_7196,N_7687);
nor U8043 (N_8043,N_7900,N_7214);
xor U8044 (N_8044,N_7707,N_7504);
nor U8045 (N_8045,N_7668,N_7094);
or U8046 (N_8046,N_7191,N_7567);
nor U8047 (N_8047,N_7179,N_7122);
or U8048 (N_8048,N_7093,N_7055);
xnor U8049 (N_8049,N_7139,N_7383);
or U8050 (N_8050,N_7371,N_7857);
nand U8051 (N_8051,N_7064,N_7477);
nor U8052 (N_8052,N_7350,N_7971);
xnor U8053 (N_8053,N_7987,N_7306);
nor U8054 (N_8054,N_7636,N_7689);
nor U8055 (N_8055,N_7272,N_7135);
and U8056 (N_8056,N_7103,N_7676);
nand U8057 (N_8057,N_7096,N_7946);
xnor U8058 (N_8058,N_7503,N_7526);
xor U8059 (N_8059,N_7076,N_7755);
xnor U8060 (N_8060,N_7141,N_7630);
or U8061 (N_8061,N_7296,N_7675);
nand U8062 (N_8062,N_7980,N_7718);
nand U8063 (N_8063,N_7903,N_7257);
and U8064 (N_8064,N_7388,N_7428);
nand U8065 (N_8065,N_7968,N_7914);
nand U8066 (N_8066,N_7405,N_7892);
xor U8067 (N_8067,N_7701,N_7051);
or U8068 (N_8068,N_7800,N_7229);
xnor U8069 (N_8069,N_7832,N_7033);
nand U8070 (N_8070,N_7966,N_7533);
nor U8071 (N_8071,N_7261,N_7481);
and U8072 (N_8072,N_7474,N_7250);
nor U8073 (N_8073,N_7397,N_7806);
xnor U8074 (N_8074,N_7854,N_7731);
xnor U8075 (N_8075,N_7435,N_7084);
or U8076 (N_8076,N_7426,N_7622);
xor U8077 (N_8077,N_7548,N_7356);
xnor U8078 (N_8078,N_7492,N_7357);
and U8079 (N_8079,N_7819,N_7409);
and U8080 (N_8080,N_7036,N_7572);
and U8081 (N_8081,N_7195,N_7606);
or U8082 (N_8082,N_7341,N_7437);
or U8083 (N_8083,N_7015,N_7006);
xor U8084 (N_8084,N_7042,N_7244);
xor U8085 (N_8085,N_7352,N_7847);
or U8086 (N_8086,N_7535,N_7765);
nand U8087 (N_8087,N_7721,N_7043);
nor U8088 (N_8088,N_7575,N_7650);
or U8089 (N_8089,N_7175,N_7716);
or U8090 (N_8090,N_7846,N_7276);
nor U8091 (N_8091,N_7863,N_7274);
nand U8092 (N_8092,N_7612,N_7071);
xor U8093 (N_8093,N_7029,N_7030);
xor U8094 (N_8094,N_7508,N_7838);
nor U8095 (N_8095,N_7955,N_7666);
and U8096 (N_8096,N_7910,N_7805);
nand U8097 (N_8097,N_7670,N_7332);
or U8098 (N_8098,N_7079,N_7709);
nor U8099 (N_8099,N_7434,N_7802);
or U8100 (N_8100,N_7140,N_7759);
nor U8101 (N_8101,N_7986,N_7167);
nand U8102 (N_8102,N_7528,N_7501);
or U8103 (N_8103,N_7952,N_7515);
or U8104 (N_8104,N_7281,N_7101);
xnor U8105 (N_8105,N_7011,N_7932);
nor U8106 (N_8106,N_7112,N_7331);
xnor U8107 (N_8107,N_7957,N_7629);
and U8108 (N_8108,N_7279,N_7496);
or U8109 (N_8109,N_7764,N_7912);
or U8110 (N_8110,N_7542,N_7605);
or U8111 (N_8111,N_7761,N_7640);
xnor U8112 (N_8112,N_7811,N_7156);
nor U8113 (N_8113,N_7110,N_7406);
nand U8114 (N_8114,N_7165,N_7859);
nand U8115 (N_8115,N_7180,N_7192);
xnor U8116 (N_8116,N_7482,N_7786);
or U8117 (N_8117,N_7750,N_7164);
or U8118 (N_8118,N_7412,N_7944);
nand U8119 (N_8119,N_7182,N_7221);
or U8120 (N_8120,N_7473,N_7713);
or U8121 (N_8121,N_7516,N_7861);
nor U8122 (N_8122,N_7403,N_7194);
and U8123 (N_8123,N_7308,N_7413);
nand U8124 (N_8124,N_7977,N_7088);
nor U8125 (N_8125,N_7326,N_7137);
and U8126 (N_8126,N_7858,N_7022);
nand U8127 (N_8127,N_7671,N_7291);
xnor U8128 (N_8128,N_7730,N_7563);
or U8129 (N_8129,N_7399,N_7999);
xnor U8130 (N_8130,N_7995,N_7807);
nor U8131 (N_8131,N_7734,N_7316);
nor U8132 (N_8132,N_7348,N_7599);
nand U8133 (N_8133,N_7465,N_7284);
nand U8134 (N_8134,N_7753,N_7420);
xor U8135 (N_8135,N_7688,N_7089);
nand U8136 (N_8136,N_7522,N_7908);
xor U8137 (N_8137,N_7448,N_7615);
nor U8138 (N_8138,N_7566,N_7451);
or U8139 (N_8139,N_7983,N_7581);
nor U8140 (N_8140,N_7480,N_7085);
nor U8141 (N_8141,N_7183,N_7068);
and U8142 (N_8142,N_7659,N_7519);
nand U8143 (N_8143,N_7875,N_7290);
xor U8144 (N_8144,N_7158,N_7964);
nor U8145 (N_8145,N_7213,N_7540);
nand U8146 (N_8146,N_7518,N_7849);
and U8147 (N_8147,N_7418,N_7500);
xor U8148 (N_8148,N_7323,N_7610);
or U8149 (N_8149,N_7002,N_7578);
and U8150 (N_8150,N_7813,N_7635);
or U8151 (N_8151,N_7942,N_7851);
nor U8152 (N_8152,N_7470,N_7733);
nand U8153 (N_8153,N_7381,N_7186);
nand U8154 (N_8154,N_7704,N_7395);
nor U8155 (N_8155,N_7255,N_7355);
nor U8156 (N_8156,N_7661,N_7834);
and U8157 (N_8157,N_7887,N_7869);
nand U8158 (N_8158,N_7021,N_7722);
xnor U8159 (N_8159,N_7346,N_7611);
nand U8160 (N_8160,N_7928,N_7719);
and U8161 (N_8161,N_7387,N_7065);
xor U8162 (N_8162,N_7218,N_7052);
or U8163 (N_8163,N_7300,N_7010);
xnor U8164 (N_8164,N_7146,N_7442);
xnor U8165 (N_8165,N_7389,N_7994);
xor U8166 (N_8166,N_7618,N_7365);
or U8167 (N_8167,N_7328,N_7142);
or U8168 (N_8168,N_7393,N_7826);
or U8169 (N_8169,N_7249,N_7027);
nand U8170 (N_8170,N_7174,N_7072);
or U8171 (N_8171,N_7729,N_7120);
and U8172 (N_8172,N_7770,N_7993);
and U8173 (N_8173,N_7711,N_7493);
or U8174 (N_8174,N_7873,N_7265);
xnor U8175 (N_8175,N_7697,N_7367);
and U8176 (N_8176,N_7792,N_7114);
nand U8177 (N_8177,N_7524,N_7775);
xnor U8178 (N_8178,N_7109,N_7954);
or U8179 (N_8179,N_7538,N_7602);
xnor U8180 (N_8180,N_7656,N_7419);
xnor U8181 (N_8181,N_7440,N_7400);
or U8182 (N_8182,N_7374,N_7947);
and U8183 (N_8183,N_7648,N_7510);
nand U8184 (N_8184,N_7886,N_7329);
nor U8185 (N_8185,N_7517,N_7057);
nand U8186 (N_8186,N_7143,N_7880);
nand U8187 (N_8187,N_7879,N_7016);
xor U8188 (N_8188,N_7209,N_7941);
or U8189 (N_8189,N_7271,N_7568);
nor U8190 (N_8190,N_7360,N_7876);
nand U8191 (N_8191,N_7099,N_7511);
xor U8192 (N_8192,N_7008,N_7998);
and U8193 (N_8193,N_7842,N_7318);
xnor U8194 (N_8194,N_7708,N_7665);
nor U8195 (N_8195,N_7282,N_7092);
xnor U8196 (N_8196,N_7322,N_7692);
xnor U8197 (N_8197,N_7131,N_7226);
xnor U8198 (N_8198,N_7684,N_7227);
nor U8199 (N_8199,N_7937,N_7929);
nor U8200 (N_8200,N_7445,N_7580);
nor U8201 (N_8201,N_7965,N_7049);
or U8202 (N_8202,N_7233,N_7651);
nor U8203 (N_8203,N_7550,N_7746);
nor U8204 (N_8204,N_7150,N_7979);
xor U8205 (N_8205,N_7956,N_7774);
xor U8206 (N_8206,N_7658,N_7162);
nand U8207 (N_8207,N_7311,N_7380);
and U8208 (N_8208,N_7973,N_7116);
or U8209 (N_8209,N_7415,N_7628);
nor U8210 (N_8210,N_7211,N_7410);
or U8211 (N_8211,N_7877,N_7349);
nand U8212 (N_8212,N_7555,N_7169);
or U8213 (N_8213,N_7913,N_7940);
nor U8214 (N_8214,N_7781,N_7577);
nand U8215 (N_8215,N_7171,N_7818);
or U8216 (N_8216,N_7031,N_7292);
and U8217 (N_8217,N_7458,N_7416);
nor U8218 (N_8218,N_7990,N_7924);
and U8219 (N_8219,N_7803,N_7588);
and U8220 (N_8220,N_7696,N_7794);
nor U8221 (N_8221,N_7004,N_7304);
nor U8222 (N_8222,N_7881,N_7507);
nor U8223 (N_8223,N_7660,N_7337);
nor U8224 (N_8224,N_7314,N_7173);
xnor U8225 (N_8225,N_7830,N_7982);
or U8226 (N_8226,N_7153,N_7690);
nand U8227 (N_8227,N_7839,N_7275);
nor U8228 (N_8228,N_7040,N_7958);
xor U8229 (N_8229,N_7444,N_7038);
or U8230 (N_8230,N_7425,N_7238);
xnor U8231 (N_8231,N_7831,N_7354);
and U8232 (N_8232,N_7564,N_7923);
or U8233 (N_8233,N_7200,N_7256);
and U8234 (N_8234,N_7569,N_7613);
and U8235 (N_8235,N_7080,N_7607);
nor U8236 (N_8236,N_7320,N_7185);
or U8237 (N_8237,N_7432,N_7752);
nor U8238 (N_8238,N_7654,N_7897);
nor U8239 (N_8239,N_7309,N_7682);
nand U8240 (N_8240,N_7013,N_7960);
and U8241 (N_8241,N_7260,N_7152);
nand U8242 (N_8242,N_7107,N_7223);
or U8243 (N_8243,N_7307,N_7975);
xor U8244 (N_8244,N_7460,N_7835);
xnor U8245 (N_8245,N_7144,N_7885);
nor U8246 (N_8246,N_7203,N_7047);
and U8247 (N_8247,N_7336,N_7375);
or U8248 (N_8248,N_7561,N_7310);
nand U8249 (N_8249,N_7560,N_7889);
nand U8250 (N_8250,N_7126,N_7591);
and U8251 (N_8251,N_7520,N_7453);
nand U8252 (N_8252,N_7936,N_7121);
xor U8253 (N_8253,N_7901,N_7188);
nor U8254 (N_8254,N_7554,N_7837);
nand U8255 (N_8255,N_7760,N_7537);
nor U8256 (N_8256,N_7582,N_7514);
xor U8257 (N_8257,N_7549,N_7075);
nand U8258 (N_8258,N_7231,N_7335);
xor U8259 (N_8259,N_7667,N_7976);
or U8260 (N_8260,N_7366,N_7804);
xnor U8261 (N_8261,N_7681,N_7170);
nand U8262 (N_8262,N_7565,N_7780);
and U8263 (N_8263,N_7254,N_7083);
nor U8264 (N_8264,N_7732,N_7299);
xor U8265 (N_8265,N_7408,N_7757);
and U8266 (N_8266,N_7270,N_7091);
and U8267 (N_8267,N_7872,N_7758);
nand U8268 (N_8268,N_7237,N_7893);
nand U8269 (N_8269,N_7625,N_7724);
nand U8270 (N_8270,N_7649,N_7498);
nand U8271 (N_8271,N_7154,N_7475);
and U8272 (N_8272,N_7225,N_7117);
xnor U8273 (N_8273,N_7601,N_7044);
nor U8274 (N_8274,N_7815,N_7978);
or U8275 (N_8275,N_7509,N_7870);
xor U8276 (N_8276,N_7372,N_7269);
and U8277 (N_8277,N_7710,N_7603);
and U8278 (N_8278,N_7172,N_7106);
xor U8279 (N_8279,N_7521,N_7104);
and U8280 (N_8280,N_7609,N_7032);
nor U8281 (N_8281,N_7014,N_7862);
xor U8282 (N_8282,N_7129,N_7438);
or U8283 (N_8283,N_7178,N_7204);
nand U8284 (N_8284,N_7793,N_7334);
xor U8285 (N_8285,N_7860,N_7919);
nor U8286 (N_8286,N_7723,N_7997);
xnor U8287 (N_8287,N_7809,N_7902);
and U8288 (N_8288,N_7621,N_7012);
nor U8289 (N_8289,N_7895,N_7552);
nor U8290 (N_8290,N_7985,N_7486);
xnor U8291 (N_8291,N_7878,N_7090);
or U8292 (N_8292,N_7545,N_7882);
nand U8293 (N_8293,N_7224,N_7487);
and U8294 (N_8294,N_7078,N_7285);
or U8295 (N_8295,N_7703,N_7077);
and U8296 (N_8296,N_7187,N_7715);
nor U8297 (N_8297,N_7996,N_7574);
nand U8298 (N_8298,N_7396,N_7201);
or U8299 (N_8299,N_7417,N_7392);
and U8300 (N_8300,N_7735,N_7151);
nor U8301 (N_8301,N_7132,N_7048);
and U8302 (N_8302,N_7583,N_7546);
xnor U8303 (N_8303,N_7447,N_7268);
and U8304 (N_8304,N_7108,N_7820);
or U8305 (N_8305,N_7801,N_7896);
nor U8306 (N_8306,N_7871,N_7828);
or U8307 (N_8307,N_7930,N_7313);
or U8308 (N_8308,N_7747,N_7390);
or U8309 (N_8309,N_7045,N_7280);
xor U8310 (N_8310,N_7236,N_7647);
nor U8311 (N_8311,N_7208,N_7544);
nand U8312 (N_8312,N_7215,N_7148);
and U8313 (N_8313,N_7594,N_7812);
and U8314 (N_8314,N_7641,N_7992);
xnor U8315 (N_8315,N_7614,N_7386);
nor U8316 (N_8316,N_7541,N_7138);
xor U8317 (N_8317,N_7097,N_7769);
nand U8318 (N_8318,N_7364,N_7430);
xnor U8319 (N_8319,N_7422,N_7543);
xnor U8320 (N_8320,N_7198,N_7748);
and U8321 (N_8321,N_7778,N_7497);
nor U8322 (N_8322,N_7926,N_7845);
and U8323 (N_8323,N_7698,N_7127);
or U8324 (N_8324,N_7305,N_7789);
nand U8325 (N_8325,N_7825,N_7294);
or U8326 (N_8326,N_7534,N_7981);
nand U8327 (N_8327,N_7590,N_7843);
xor U8328 (N_8328,N_7691,N_7633);
nand U8329 (N_8329,N_7934,N_7680);
nand U8330 (N_8330,N_7865,N_7974);
nand U8331 (N_8331,N_7663,N_7478);
or U8332 (N_8332,N_7333,N_7246);
nand U8333 (N_8333,N_7061,N_7678);
or U8334 (N_8334,N_7505,N_7799);
or U8335 (N_8335,N_7370,N_7252);
xnor U8336 (N_8336,N_7777,N_7967);
nor U8337 (N_8337,N_7714,N_7134);
nand U8338 (N_8338,N_7531,N_7489);
or U8339 (N_8339,N_7571,N_7645);
xor U8340 (N_8340,N_7073,N_7962);
nor U8341 (N_8341,N_7069,N_7087);
nor U8342 (N_8342,N_7939,N_7407);
xnor U8343 (N_8343,N_7784,N_7771);
xor U8344 (N_8344,N_7124,N_7557);
nor U8345 (N_8345,N_7066,N_7788);
nor U8346 (N_8346,N_7626,N_7970);
and U8347 (N_8347,N_7228,N_7576);
nor U8348 (N_8348,N_7797,N_7988);
nor U8349 (N_8349,N_7450,N_7953);
xnor U8350 (N_8350,N_7920,N_7024);
or U8351 (N_8351,N_7884,N_7827);
nand U8352 (N_8352,N_7657,N_7456);
or U8353 (N_8353,N_7377,N_7210);
nor U8354 (N_8354,N_7028,N_7699);
nor U8355 (N_8355,N_7536,N_7829);
nor U8356 (N_8356,N_7017,N_7664);
and U8357 (N_8357,N_7653,N_7959);
nor U8358 (N_8358,N_7197,N_7585);
nand U8359 (N_8359,N_7586,N_7620);
nor U8360 (N_8360,N_7499,N_7060);
nand U8361 (N_8361,N_7039,N_7289);
nand U8362 (N_8362,N_7814,N_7302);
nand U8363 (N_8363,N_7627,N_7677);
nand U8364 (N_8364,N_7020,N_7362);
and U8365 (N_8365,N_7398,N_7824);
and U8366 (N_8366,N_7921,N_7702);
nand U8367 (N_8367,N_7726,N_7401);
or U8368 (N_8368,N_7159,N_7287);
and U8369 (N_8369,N_7744,N_7712);
nor U8370 (N_8370,N_7506,N_7059);
nor U8371 (N_8371,N_7023,N_7853);
nand U8372 (N_8372,N_7742,N_7911);
nor U8373 (N_8373,N_7111,N_7081);
and U8374 (N_8374,N_7841,N_7795);
nor U8375 (N_8375,N_7457,N_7624);
nor U8376 (N_8376,N_7277,N_7909);
nand U8377 (N_8377,N_7925,N_7247);
nor U8378 (N_8378,N_7446,N_7695);
and U8379 (N_8379,N_7161,N_7219);
nor U8380 (N_8380,N_7113,N_7798);
or U8381 (N_8381,N_7513,N_7596);
xnor U8382 (N_8382,N_7562,N_7471);
xnor U8383 (N_8383,N_7391,N_7086);
nor U8384 (N_8384,N_7850,N_7705);
nand U8385 (N_8385,N_7273,N_7969);
nand U8386 (N_8386,N_7423,N_7644);
nand U8387 (N_8387,N_7205,N_7915);
nand U8388 (N_8388,N_7483,N_7963);
and U8389 (N_8389,N_7199,N_7429);
xnor U8390 (N_8390,N_7848,N_7258);
xor U8391 (N_8391,N_7894,N_7454);
nor U8392 (N_8392,N_7810,N_7253);
and U8393 (N_8393,N_7669,N_7787);
or U8394 (N_8394,N_7009,N_7123);
xnor U8395 (N_8395,N_7149,N_7790);
and U8396 (N_8396,N_7864,N_7342);
nand U8397 (N_8397,N_7559,N_7376);
or U8398 (N_8398,N_7100,N_7046);
nor U8399 (N_8399,N_7931,N_7888);
xor U8400 (N_8400,N_7821,N_7679);
or U8401 (N_8401,N_7935,N_7808);
nor U8402 (N_8402,N_7345,N_7866);
and U8403 (N_8403,N_7319,N_7469);
or U8404 (N_8404,N_7321,N_7344);
xnor U8405 (N_8405,N_7856,N_7539);
nor U8406 (N_8406,N_7502,N_7662);
nor U8407 (N_8407,N_7776,N_7617);
xor U8408 (N_8408,N_7382,N_7836);
nand U8409 (N_8409,N_7163,N_7763);
and U8410 (N_8410,N_7700,N_7619);
nand U8411 (N_8411,N_7479,N_7720);
or U8412 (N_8412,N_7484,N_7899);
nand U8413 (N_8413,N_7476,N_7315);
nand U8414 (N_8414,N_7402,N_7595);
or U8415 (N_8415,N_7949,N_7532);
nand U8416 (N_8416,N_7018,N_7683);
nor U8417 (N_8417,N_7783,N_7485);
xor U8418 (N_8418,N_7234,N_7655);
and U8419 (N_8419,N_7358,N_7587);
nand U8420 (N_8420,N_7074,N_7938);
or U8421 (N_8421,N_7176,N_7785);
and U8422 (N_8422,N_7616,N_7740);
xor U8423 (N_8423,N_7082,N_7001);
and U8424 (N_8424,N_7951,N_7948);
and U8425 (N_8425,N_7833,N_7907);
or U8426 (N_8426,N_7491,N_7007);
xnor U8427 (N_8427,N_7570,N_7421);
nand U8428 (N_8428,N_7916,N_7608);
nand U8429 (N_8429,N_7062,N_7589);
nand U8430 (N_8430,N_7593,N_7462);
nor U8431 (N_8431,N_7439,N_7259);
nor U8432 (N_8432,N_7168,N_7472);
nor U8433 (N_8433,N_7989,N_7972);
nor U8434 (N_8434,N_7488,N_7220);
nor U8435 (N_8435,N_7768,N_7905);
or U8436 (N_8436,N_7005,N_7239);
nand U8437 (N_8437,N_7312,N_7556);
xor U8438 (N_8438,N_7041,N_7772);
nand U8439 (N_8439,N_7034,N_7243);
and U8440 (N_8440,N_7361,N_7693);
xor U8441 (N_8441,N_7433,N_7782);
nand U8442 (N_8442,N_7706,N_7293);
nand U8443 (N_8443,N_7694,N_7353);
or U8444 (N_8444,N_7686,N_7431);
and U8445 (N_8445,N_7193,N_7455);
or U8446 (N_8446,N_7717,N_7918);
nand U8447 (N_8447,N_7206,N_7597);
xnor U8448 (N_8448,N_7118,N_7891);
nand U8449 (N_8449,N_7459,N_7000);
xor U8450 (N_8450,N_7301,N_7102);
xor U8451 (N_8451,N_7145,N_7378);
xor U8452 (N_8452,N_7166,N_7553);
nand U8453 (N_8453,N_7098,N_7262);
xnor U8454 (N_8454,N_7933,N_7823);
nor U8455 (N_8455,N_7922,N_7266);
nand U8456 (N_8456,N_7898,N_7385);
and U8457 (N_8457,N_7674,N_7147);
or U8458 (N_8458,N_7288,N_7592);
nand U8459 (N_8459,N_7427,N_7298);
nand U8460 (N_8460,N_7762,N_7324);
nor U8461 (N_8461,N_7773,N_7212);
xnor U8462 (N_8462,N_7411,N_7095);
xnor U8463 (N_8463,N_7652,N_7840);
xnor U8464 (N_8464,N_7155,N_7125);
or U8465 (N_8465,N_7738,N_7754);
nand U8466 (N_8466,N_7359,N_7558);
nand U8467 (N_8467,N_7736,N_7441);
or U8468 (N_8468,N_7404,N_7791);
nand U8469 (N_8469,N_7384,N_7638);
xnor U8470 (N_8470,N_7058,N_7623);
and U8471 (N_8471,N_7157,N_7512);
nor U8472 (N_8472,N_7207,N_7739);
nor U8473 (N_8473,N_7105,N_7240);
nor U8474 (N_8474,N_7796,N_7579);
xor U8475 (N_8475,N_7984,N_7904);
and U8476 (N_8476,N_7436,N_7646);
xnor U8477 (N_8477,N_7452,N_7547);
nand U8478 (N_8478,N_7749,N_7673);
nand U8479 (N_8479,N_7631,N_7727);
xnor U8480 (N_8480,N_7053,N_7177);
nand U8481 (N_8481,N_7961,N_7056);
or U8482 (N_8482,N_7130,N_7855);
xor U8483 (N_8483,N_7222,N_7551);
nor U8484 (N_8484,N_7128,N_7343);
and U8485 (N_8485,N_7019,N_7600);
nand U8486 (N_8486,N_7330,N_7685);
and U8487 (N_8487,N_7883,N_7890);
xnor U8488 (N_8488,N_7414,N_7639);
nand U8489 (N_8489,N_7025,N_7637);
or U8490 (N_8490,N_7267,N_7745);
xnor U8491 (N_8491,N_7026,N_7245);
or U8492 (N_8492,N_7297,N_7604);
nand U8493 (N_8493,N_7927,N_7067);
or U8494 (N_8494,N_7584,N_7217);
nand U8495 (N_8495,N_7443,N_7779);
nor U8496 (N_8496,N_7766,N_7232);
nor U8497 (N_8497,N_7525,N_7466);
and U8498 (N_8498,N_7133,N_7725);
and U8499 (N_8499,N_7263,N_7852);
nand U8500 (N_8500,N_7283,N_7976);
nand U8501 (N_8501,N_7217,N_7288);
and U8502 (N_8502,N_7362,N_7987);
xor U8503 (N_8503,N_7236,N_7208);
or U8504 (N_8504,N_7219,N_7014);
or U8505 (N_8505,N_7189,N_7709);
or U8506 (N_8506,N_7662,N_7536);
xor U8507 (N_8507,N_7360,N_7020);
nand U8508 (N_8508,N_7104,N_7967);
and U8509 (N_8509,N_7851,N_7830);
nand U8510 (N_8510,N_7340,N_7145);
xor U8511 (N_8511,N_7696,N_7949);
nor U8512 (N_8512,N_7228,N_7747);
or U8513 (N_8513,N_7612,N_7505);
xor U8514 (N_8514,N_7540,N_7394);
xnor U8515 (N_8515,N_7934,N_7964);
xnor U8516 (N_8516,N_7369,N_7425);
or U8517 (N_8517,N_7664,N_7072);
or U8518 (N_8518,N_7856,N_7562);
and U8519 (N_8519,N_7488,N_7140);
xor U8520 (N_8520,N_7468,N_7365);
xnor U8521 (N_8521,N_7355,N_7558);
and U8522 (N_8522,N_7499,N_7866);
and U8523 (N_8523,N_7905,N_7073);
nand U8524 (N_8524,N_7612,N_7919);
nor U8525 (N_8525,N_7763,N_7809);
nand U8526 (N_8526,N_7050,N_7988);
or U8527 (N_8527,N_7011,N_7353);
xnor U8528 (N_8528,N_7181,N_7563);
xnor U8529 (N_8529,N_7203,N_7537);
nand U8530 (N_8530,N_7854,N_7683);
or U8531 (N_8531,N_7401,N_7182);
or U8532 (N_8532,N_7442,N_7215);
and U8533 (N_8533,N_7869,N_7344);
nand U8534 (N_8534,N_7372,N_7040);
or U8535 (N_8535,N_7185,N_7870);
and U8536 (N_8536,N_7688,N_7272);
nand U8537 (N_8537,N_7545,N_7014);
nand U8538 (N_8538,N_7877,N_7975);
and U8539 (N_8539,N_7896,N_7459);
nor U8540 (N_8540,N_7485,N_7704);
nand U8541 (N_8541,N_7259,N_7252);
nand U8542 (N_8542,N_7724,N_7088);
and U8543 (N_8543,N_7582,N_7161);
nor U8544 (N_8544,N_7360,N_7586);
nand U8545 (N_8545,N_7789,N_7893);
and U8546 (N_8546,N_7135,N_7718);
xnor U8547 (N_8547,N_7088,N_7252);
nand U8548 (N_8548,N_7937,N_7413);
xor U8549 (N_8549,N_7045,N_7060);
xor U8550 (N_8550,N_7197,N_7517);
xnor U8551 (N_8551,N_7333,N_7632);
or U8552 (N_8552,N_7442,N_7278);
xnor U8553 (N_8553,N_7702,N_7845);
or U8554 (N_8554,N_7578,N_7744);
nor U8555 (N_8555,N_7583,N_7225);
and U8556 (N_8556,N_7068,N_7666);
and U8557 (N_8557,N_7991,N_7719);
or U8558 (N_8558,N_7754,N_7430);
nor U8559 (N_8559,N_7631,N_7451);
nor U8560 (N_8560,N_7672,N_7535);
nand U8561 (N_8561,N_7165,N_7432);
or U8562 (N_8562,N_7511,N_7414);
and U8563 (N_8563,N_7600,N_7399);
or U8564 (N_8564,N_7808,N_7931);
and U8565 (N_8565,N_7190,N_7775);
xor U8566 (N_8566,N_7596,N_7316);
nand U8567 (N_8567,N_7027,N_7419);
and U8568 (N_8568,N_7540,N_7399);
and U8569 (N_8569,N_7418,N_7676);
and U8570 (N_8570,N_7440,N_7196);
or U8571 (N_8571,N_7787,N_7878);
or U8572 (N_8572,N_7245,N_7395);
and U8573 (N_8573,N_7592,N_7139);
xor U8574 (N_8574,N_7947,N_7003);
nand U8575 (N_8575,N_7963,N_7373);
or U8576 (N_8576,N_7085,N_7623);
or U8577 (N_8577,N_7355,N_7464);
nand U8578 (N_8578,N_7216,N_7923);
and U8579 (N_8579,N_7207,N_7070);
nor U8580 (N_8580,N_7621,N_7338);
nand U8581 (N_8581,N_7324,N_7071);
xor U8582 (N_8582,N_7817,N_7546);
and U8583 (N_8583,N_7632,N_7694);
or U8584 (N_8584,N_7413,N_7747);
nand U8585 (N_8585,N_7095,N_7660);
or U8586 (N_8586,N_7027,N_7947);
and U8587 (N_8587,N_7261,N_7079);
and U8588 (N_8588,N_7050,N_7544);
or U8589 (N_8589,N_7666,N_7637);
xnor U8590 (N_8590,N_7375,N_7069);
or U8591 (N_8591,N_7520,N_7070);
nor U8592 (N_8592,N_7635,N_7025);
or U8593 (N_8593,N_7471,N_7313);
nand U8594 (N_8594,N_7769,N_7056);
or U8595 (N_8595,N_7441,N_7816);
nor U8596 (N_8596,N_7998,N_7185);
nand U8597 (N_8597,N_7548,N_7680);
or U8598 (N_8598,N_7198,N_7140);
and U8599 (N_8599,N_7584,N_7727);
nor U8600 (N_8600,N_7081,N_7739);
nor U8601 (N_8601,N_7948,N_7271);
nor U8602 (N_8602,N_7035,N_7016);
nor U8603 (N_8603,N_7955,N_7858);
and U8604 (N_8604,N_7755,N_7090);
and U8605 (N_8605,N_7198,N_7529);
or U8606 (N_8606,N_7365,N_7123);
and U8607 (N_8607,N_7412,N_7342);
xnor U8608 (N_8608,N_7787,N_7645);
or U8609 (N_8609,N_7646,N_7428);
nor U8610 (N_8610,N_7366,N_7445);
nand U8611 (N_8611,N_7797,N_7069);
nand U8612 (N_8612,N_7742,N_7146);
and U8613 (N_8613,N_7088,N_7723);
xor U8614 (N_8614,N_7090,N_7347);
nand U8615 (N_8615,N_7271,N_7172);
or U8616 (N_8616,N_7996,N_7666);
or U8617 (N_8617,N_7418,N_7982);
xnor U8618 (N_8618,N_7747,N_7052);
nand U8619 (N_8619,N_7554,N_7564);
nand U8620 (N_8620,N_7131,N_7665);
nor U8621 (N_8621,N_7293,N_7250);
nor U8622 (N_8622,N_7320,N_7495);
nor U8623 (N_8623,N_7897,N_7458);
xnor U8624 (N_8624,N_7809,N_7511);
or U8625 (N_8625,N_7574,N_7268);
nand U8626 (N_8626,N_7249,N_7276);
or U8627 (N_8627,N_7269,N_7924);
xnor U8628 (N_8628,N_7805,N_7828);
and U8629 (N_8629,N_7694,N_7517);
or U8630 (N_8630,N_7346,N_7417);
nor U8631 (N_8631,N_7341,N_7220);
and U8632 (N_8632,N_7931,N_7285);
or U8633 (N_8633,N_7142,N_7528);
nand U8634 (N_8634,N_7417,N_7137);
or U8635 (N_8635,N_7870,N_7144);
and U8636 (N_8636,N_7058,N_7294);
nor U8637 (N_8637,N_7842,N_7605);
and U8638 (N_8638,N_7912,N_7862);
xnor U8639 (N_8639,N_7286,N_7370);
nand U8640 (N_8640,N_7328,N_7293);
or U8641 (N_8641,N_7220,N_7590);
or U8642 (N_8642,N_7368,N_7620);
or U8643 (N_8643,N_7170,N_7378);
nor U8644 (N_8644,N_7269,N_7870);
nand U8645 (N_8645,N_7712,N_7185);
or U8646 (N_8646,N_7087,N_7393);
nor U8647 (N_8647,N_7403,N_7294);
xor U8648 (N_8648,N_7931,N_7608);
nand U8649 (N_8649,N_7803,N_7857);
nor U8650 (N_8650,N_7724,N_7392);
nand U8651 (N_8651,N_7141,N_7916);
xor U8652 (N_8652,N_7310,N_7749);
and U8653 (N_8653,N_7370,N_7593);
and U8654 (N_8654,N_7995,N_7608);
nand U8655 (N_8655,N_7360,N_7499);
xnor U8656 (N_8656,N_7171,N_7175);
or U8657 (N_8657,N_7095,N_7240);
and U8658 (N_8658,N_7054,N_7478);
nand U8659 (N_8659,N_7882,N_7135);
and U8660 (N_8660,N_7504,N_7057);
nor U8661 (N_8661,N_7927,N_7490);
nand U8662 (N_8662,N_7150,N_7085);
nand U8663 (N_8663,N_7960,N_7167);
and U8664 (N_8664,N_7511,N_7698);
and U8665 (N_8665,N_7785,N_7354);
nand U8666 (N_8666,N_7193,N_7437);
nor U8667 (N_8667,N_7345,N_7688);
nand U8668 (N_8668,N_7197,N_7072);
xor U8669 (N_8669,N_7871,N_7518);
or U8670 (N_8670,N_7097,N_7849);
nand U8671 (N_8671,N_7137,N_7426);
xor U8672 (N_8672,N_7601,N_7640);
or U8673 (N_8673,N_7458,N_7864);
nand U8674 (N_8674,N_7455,N_7328);
nor U8675 (N_8675,N_7694,N_7037);
nand U8676 (N_8676,N_7758,N_7924);
nand U8677 (N_8677,N_7050,N_7750);
nand U8678 (N_8678,N_7445,N_7284);
nor U8679 (N_8679,N_7664,N_7133);
or U8680 (N_8680,N_7080,N_7834);
nor U8681 (N_8681,N_7397,N_7582);
and U8682 (N_8682,N_7064,N_7795);
and U8683 (N_8683,N_7939,N_7955);
and U8684 (N_8684,N_7329,N_7589);
nand U8685 (N_8685,N_7023,N_7199);
or U8686 (N_8686,N_7634,N_7918);
and U8687 (N_8687,N_7369,N_7443);
nor U8688 (N_8688,N_7999,N_7366);
nand U8689 (N_8689,N_7935,N_7270);
nand U8690 (N_8690,N_7338,N_7827);
or U8691 (N_8691,N_7595,N_7780);
or U8692 (N_8692,N_7801,N_7758);
and U8693 (N_8693,N_7716,N_7579);
or U8694 (N_8694,N_7866,N_7689);
or U8695 (N_8695,N_7233,N_7466);
nor U8696 (N_8696,N_7865,N_7829);
and U8697 (N_8697,N_7235,N_7481);
xor U8698 (N_8698,N_7768,N_7140);
nand U8699 (N_8699,N_7302,N_7470);
nor U8700 (N_8700,N_7452,N_7543);
and U8701 (N_8701,N_7500,N_7344);
and U8702 (N_8702,N_7535,N_7007);
or U8703 (N_8703,N_7914,N_7181);
nor U8704 (N_8704,N_7155,N_7781);
or U8705 (N_8705,N_7493,N_7799);
or U8706 (N_8706,N_7988,N_7975);
nand U8707 (N_8707,N_7914,N_7419);
nand U8708 (N_8708,N_7024,N_7413);
nor U8709 (N_8709,N_7934,N_7751);
xnor U8710 (N_8710,N_7168,N_7549);
and U8711 (N_8711,N_7645,N_7319);
nor U8712 (N_8712,N_7895,N_7905);
xor U8713 (N_8713,N_7174,N_7678);
and U8714 (N_8714,N_7009,N_7816);
or U8715 (N_8715,N_7305,N_7921);
nor U8716 (N_8716,N_7418,N_7353);
and U8717 (N_8717,N_7704,N_7170);
nor U8718 (N_8718,N_7257,N_7692);
nand U8719 (N_8719,N_7934,N_7890);
nand U8720 (N_8720,N_7606,N_7726);
or U8721 (N_8721,N_7599,N_7540);
and U8722 (N_8722,N_7312,N_7045);
nor U8723 (N_8723,N_7802,N_7411);
or U8724 (N_8724,N_7346,N_7680);
or U8725 (N_8725,N_7196,N_7623);
and U8726 (N_8726,N_7007,N_7506);
or U8727 (N_8727,N_7485,N_7403);
or U8728 (N_8728,N_7418,N_7478);
or U8729 (N_8729,N_7609,N_7197);
or U8730 (N_8730,N_7835,N_7355);
xnor U8731 (N_8731,N_7409,N_7429);
nand U8732 (N_8732,N_7666,N_7974);
or U8733 (N_8733,N_7396,N_7807);
or U8734 (N_8734,N_7307,N_7047);
nand U8735 (N_8735,N_7119,N_7664);
and U8736 (N_8736,N_7626,N_7000);
nand U8737 (N_8737,N_7963,N_7803);
and U8738 (N_8738,N_7376,N_7429);
and U8739 (N_8739,N_7595,N_7787);
or U8740 (N_8740,N_7073,N_7576);
nor U8741 (N_8741,N_7300,N_7343);
and U8742 (N_8742,N_7145,N_7458);
xor U8743 (N_8743,N_7349,N_7818);
nand U8744 (N_8744,N_7930,N_7632);
or U8745 (N_8745,N_7257,N_7281);
or U8746 (N_8746,N_7536,N_7467);
nor U8747 (N_8747,N_7127,N_7122);
nand U8748 (N_8748,N_7225,N_7954);
and U8749 (N_8749,N_7858,N_7659);
nor U8750 (N_8750,N_7411,N_7678);
xor U8751 (N_8751,N_7988,N_7167);
or U8752 (N_8752,N_7678,N_7945);
nor U8753 (N_8753,N_7213,N_7178);
or U8754 (N_8754,N_7590,N_7465);
xnor U8755 (N_8755,N_7809,N_7546);
xnor U8756 (N_8756,N_7513,N_7730);
and U8757 (N_8757,N_7827,N_7342);
or U8758 (N_8758,N_7559,N_7828);
or U8759 (N_8759,N_7931,N_7343);
nand U8760 (N_8760,N_7473,N_7867);
xnor U8761 (N_8761,N_7560,N_7380);
nand U8762 (N_8762,N_7463,N_7948);
nand U8763 (N_8763,N_7621,N_7246);
and U8764 (N_8764,N_7988,N_7960);
xor U8765 (N_8765,N_7515,N_7336);
and U8766 (N_8766,N_7576,N_7708);
nand U8767 (N_8767,N_7415,N_7525);
nand U8768 (N_8768,N_7494,N_7865);
xnor U8769 (N_8769,N_7914,N_7477);
and U8770 (N_8770,N_7989,N_7026);
nand U8771 (N_8771,N_7292,N_7158);
and U8772 (N_8772,N_7146,N_7401);
nor U8773 (N_8773,N_7926,N_7606);
or U8774 (N_8774,N_7370,N_7208);
or U8775 (N_8775,N_7991,N_7638);
nand U8776 (N_8776,N_7198,N_7063);
nor U8777 (N_8777,N_7071,N_7955);
nor U8778 (N_8778,N_7080,N_7454);
nor U8779 (N_8779,N_7119,N_7879);
or U8780 (N_8780,N_7982,N_7550);
and U8781 (N_8781,N_7069,N_7202);
nor U8782 (N_8782,N_7067,N_7557);
xor U8783 (N_8783,N_7416,N_7522);
nand U8784 (N_8784,N_7338,N_7840);
nor U8785 (N_8785,N_7983,N_7440);
nand U8786 (N_8786,N_7354,N_7489);
nor U8787 (N_8787,N_7205,N_7021);
nand U8788 (N_8788,N_7470,N_7999);
nor U8789 (N_8789,N_7606,N_7521);
and U8790 (N_8790,N_7630,N_7577);
nand U8791 (N_8791,N_7418,N_7149);
xnor U8792 (N_8792,N_7400,N_7740);
and U8793 (N_8793,N_7269,N_7880);
or U8794 (N_8794,N_7933,N_7564);
xor U8795 (N_8795,N_7862,N_7449);
or U8796 (N_8796,N_7544,N_7410);
or U8797 (N_8797,N_7910,N_7148);
xnor U8798 (N_8798,N_7684,N_7065);
and U8799 (N_8799,N_7836,N_7147);
nand U8800 (N_8800,N_7743,N_7944);
nor U8801 (N_8801,N_7079,N_7911);
and U8802 (N_8802,N_7289,N_7561);
and U8803 (N_8803,N_7423,N_7509);
and U8804 (N_8804,N_7460,N_7795);
xor U8805 (N_8805,N_7902,N_7484);
nand U8806 (N_8806,N_7958,N_7582);
nand U8807 (N_8807,N_7466,N_7482);
nor U8808 (N_8808,N_7740,N_7792);
nand U8809 (N_8809,N_7858,N_7037);
nand U8810 (N_8810,N_7224,N_7373);
nor U8811 (N_8811,N_7576,N_7310);
nand U8812 (N_8812,N_7596,N_7266);
nor U8813 (N_8813,N_7061,N_7147);
or U8814 (N_8814,N_7386,N_7132);
nor U8815 (N_8815,N_7593,N_7868);
and U8816 (N_8816,N_7253,N_7478);
xnor U8817 (N_8817,N_7071,N_7309);
and U8818 (N_8818,N_7281,N_7365);
or U8819 (N_8819,N_7181,N_7028);
xnor U8820 (N_8820,N_7020,N_7282);
or U8821 (N_8821,N_7899,N_7739);
or U8822 (N_8822,N_7512,N_7708);
nand U8823 (N_8823,N_7944,N_7485);
nor U8824 (N_8824,N_7122,N_7721);
and U8825 (N_8825,N_7394,N_7907);
or U8826 (N_8826,N_7156,N_7998);
nor U8827 (N_8827,N_7786,N_7363);
xor U8828 (N_8828,N_7559,N_7728);
nand U8829 (N_8829,N_7351,N_7987);
nor U8830 (N_8830,N_7915,N_7334);
xor U8831 (N_8831,N_7318,N_7055);
nand U8832 (N_8832,N_7676,N_7301);
nand U8833 (N_8833,N_7208,N_7484);
nor U8834 (N_8834,N_7264,N_7489);
xor U8835 (N_8835,N_7913,N_7127);
nand U8836 (N_8836,N_7711,N_7235);
xor U8837 (N_8837,N_7179,N_7603);
or U8838 (N_8838,N_7239,N_7993);
nand U8839 (N_8839,N_7595,N_7815);
xor U8840 (N_8840,N_7865,N_7299);
and U8841 (N_8841,N_7518,N_7434);
and U8842 (N_8842,N_7125,N_7691);
nor U8843 (N_8843,N_7314,N_7635);
xor U8844 (N_8844,N_7492,N_7154);
xor U8845 (N_8845,N_7928,N_7778);
nand U8846 (N_8846,N_7983,N_7547);
nor U8847 (N_8847,N_7265,N_7692);
or U8848 (N_8848,N_7196,N_7734);
or U8849 (N_8849,N_7771,N_7883);
xor U8850 (N_8850,N_7367,N_7278);
or U8851 (N_8851,N_7686,N_7007);
and U8852 (N_8852,N_7686,N_7081);
nand U8853 (N_8853,N_7665,N_7080);
nand U8854 (N_8854,N_7227,N_7037);
or U8855 (N_8855,N_7790,N_7906);
xnor U8856 (N_8856,N_7676,N_7918);
and U8857 (N_8857,N_7480,N_7321);
nand U8858 (N_8858,N_7531,N_7914);
or U8859 (N_8859,N_7513,N_7741);
nand U8860 (N_8860,N_7583,N_7138);
and U8861 (N_8861,N_7345,N_7787);
nor U8862 (N_8862,N_7920,N_7803);
xnor U8863 (N_8863,N_7741,N_7616);
xor U8864 (N_8864,N_7900,N_7466);
and U8865 (N_8865,N_7818,N_7580);
or U8866 (N_8866,N_7153,N_7834);
nand U8867 (N_8867,N_7900,N_7180);
and U8868 (N_8868,N_7517,N_7004);
nor U8869 (N_8869,N_7322,N_7848);
and U8870 (N_8870,N_7873,N_7239);
nor U8871 (N_8871,N_7532,N_7313);
nand U8872 (N_8872,N_7627,N_7731);
or U8873 (N_8873,N_7672,N_7262);
nor U8874 (N_8874,N_7747,N_7106);
nor U8875 (N_8875,N_7609,N_7987);
xnor U8876 (N_8876,N_7815,N_7793);
nand U8877 (N_8877,N_7927,N_7306);
or U8878 (N_8878,N_7006,N_7948);
or U8879 (N_8879,N_7433,N_7998);
nand U8880 (N_8880,N_7893,N_7610);
nand U8881 (N_8881,N_7624,N_7630);
nor U8882 (N_8882,N_7094,N_7172);
and U8883 (N_8883,N_7682,N_7603);
or U8884 (N_8884,N_7153,N_7547);
nor U8885 (N_8885,N_7260,N_7726);
or U8886 (N_8886,N_7638,N_7110);
nor U8887 (N_8887,N_7258,N_7914);
xor U8888 (N_8888,N_7123,N_7754);
or U8889 (N_8889,N_7048,N_7189);
xor U8890 (N_8890,N_7520,N_7165);
and U8891 (N_8891,N_7375,N_7771);
or U8892 (N_8892,N_7632,N_7846);
or U8893 (N_8893,N_7760,N_7568);
nand U8894 (N_8894,N_7029,N_7708);
and U8895 (N_8895,N_7910,N_7817);
nand U8896 (N_8896,N_7973,N_7477);
and U8897 (N_8897,N_7915,N_7254);
xor U8898 (N_8898,N_7567,N_7052);
xor U8899 (N_8899,N_7247,N_7026);
nor U8900 (N_8900,N_7087,N_7941);
nor U8901 (N_8901,N_7682,N_7776);
or U8902 (N_8902,N_7132,N_7448);
and U8903 (N_8903,N_7076,N_7793);
and U8904 (N_8904,N_7743,N_7462);
or U8905 (N_8905,N_7208,N_7984);
xor U8906 (N_8906,N_7328,N_7695);
or U8907 (N_8907,N_7813,N_7224);
nand U8908 (N_8908,N_7706,N_7959);
nor U8909 (N_8909,N_7869,N_7635);
xor U8910 (N_8910,N_7550,N_7803);
and U8911 (N_8911,N_7249,N_7661);
or U8912 (N_8912,N_7417,N_7618);
nand U8913 (N_8913,N_7545,N_7846);
nand U8914 (N_8914,N_7675,N_7739);
or U8915 (N_8915,N_7352,N_7989);
nor U8916 (N_8916,N_7261,N_7379);
nand U8917 (N_8917,N_7164,N_7417);
or U8918 (N_8918,N_7777,N_7445);
or U8919 (N_8919,N_7806,N_7801);
and U8920 (N_8920,N_7443,N_7670);
or U8921 (N_8921,N_7819,N_7828);
nand U8922 (N_8922,N_7253,N_7623);
nand U8923 (N_8923,N_7488,N_7631);
nand U8924 (N_8924,N_7281,N_7350);
and U8925 (N_8925,N_7322,N_7680);
nand U8926 (N_8926,N_7428,N_7253);
nor U8927 (N_8927,N_7907,N_7914);
nand U8928 (N_8928,N_7771,N_7541);
xor U8929 (N_8929,N_7834,N_7693);
xor U8930 (N_8930,N_7611,N_7569);
or U8931 (N_8931,N_7242,N_7338);
or U8932 (N_8932,N_7862,N_7482);
and U8933 (N_8933,N_7832,N_7346);
or U8934 (N_8934,N_7589,N_7339);
nor U8935 (N_8935,N_7307,N_7214);
or U8936 (N_8936,N_7914,N_7527);
or U8937 (N_8937,N_7893,N_7315);
or U8938 (N_8938,N_7390,N_7127);
or U8939 (N_8939,N_7695,N_7475);
nand U8940 (N_8940,N_7275,N_7331);
nor U8941 (N_8941,N_7849,N_7182);
or U8942 (N_8942,N_7756,N_7908);
or U8943 (N_8943,N_7499,N_7125);
and U8944 (N_8944,N_7038,N_7950);
and U8945 (N_8945,N_7247,N_7943);
and U8946 (N_8946,N_7070,N_7456);
xnor U8947 (N_8947,N_7643,N_7618);
nor U8948 (N_8948,N_7376,N_7443);
or U8949 (N_8949,N_7375,N_7649);
and U8950 (N_8950,N_7065,N_7373);
nor U8951 (N_8951,N_7509,N_7979);
or U8952 (N_8952,N_7536,N_7917);
nor U8953 (N_8953,N_7752,N_7926);
and U8954 (N_8954,N_7252,N_7215);
nor U8955 (N_8955,N_7879,N_7924);
xor U8956 (N_8956,N_7099,N_7664);
nor U8957 (N_8957,N_7269,N_7186);
nor U8958 (N_8958,N_7016,N_7394);
nand U8959 (N_8959,N_7257,N_7173);
or U8960 (N_8960,N_7825,N_7850);
nor U8961 (N_8961,N_7500,N_7040);
and U8962 (N_8962,N_7556,N_7107);
xnor U8963 (N_8963,N_7821,N_7828);
xnor U8964 (N_8964,N_7663,N_7967);
nor U8965 (N_8965,N_7664,N_7077);
xor U8966 (N_8966,N_7081,N_7607);
nor U8967 (N_8967,N_7594,N_7229);
or U8968 (N_8968,N_7676,N_7093);
nand U8969 (N_8969,N_7698,N_7359);
or U8970 (N_8970,N_7854,N_7668);
xnor U8971 (N_8971,N_7775,N_7055);
and U8972 (N_8972,N_7401,N_7433);
or U8973 (N_8973,N_7880,N_7331);
and U8974 (N_8974,N_7778,N_7828);
or U8975 (N_8975,N_7918,N_7387);
xor U8976 (N_8976,N_7534,N_7409);
xnor U8977 (N_8977,N_7192,N_7126);
and U8978 (N_8978,N_7147,N_7287);
nand U8979 (N_8979,N_7936,N_7732);
xor U8980 (N_8980,N_7050,N_7464);
nor U8981 (N_8981,N_7316,N_7222);
or U8982 (N_8982,N_7564,N_7719);
xnor U8983 (N_8983,N_7061,N_7017);
nand U8984 (N_8984,N_7449,N_7761);
xnor U8985 (N_8985,N_7580,N_7389);
xnor U8986 (N_8986,N_7797,N_7284);
nand U8987 (N_8987,N_7625,N_7897);
or U8988 (N_8988,N_7710,N_7833);
or U8989 (N_8989,N_7277,N_7327);
xnor U8990 (N_8990,N_7029,N_7021);
and U8991 (N_8991,N_7685,N_7903);
and U8992 (N_8992,N_7268,N_7354);
or U8993 (N_8993,N_7773,N_7060);
xnor U8994 (N_8994,N_7135,N_7739);
nand U8995 (N_8995,N_7182,N_7170);
or U8996 (N_8996,N_7678,N_7169);
xnor U8997 (N_8997,N_7626,N_7880);
xor U8998 (N_8998,N_7746,N_7903);
and U8999 (N_8999,N_7380,N_7941);
and U9000 (N_9000,N_8046,N_8359);
and U9001 (N_9001,N_8710,N_8714);
or U9002 (N_9002,N_8537,N_8028);
or U9003 (N_9003,N_8368,N_8733);
nand U9004 (N_9004,N_8533,N_8044);
nor U9005 (N_9005,N_8116,N_8174);
and U9006 (N_9006,N_8437,N_8936);
nand U9007 (N_9007,N_8867,N_8752);
xor U9008 (N_9008,N_8755,N_8062);
nor U9009 (N_9009,N_8324,N_8056);
and U9010 (N_9010,N_8943,N_8011);
or U9011 (N_9011,N_8541,N_8959);
nor U9012 (N_9012,N_8346,N_8038);
nor U9013 (N_9013,N_8683,N_8754);
xor U9014 (N_9014,N_8309,N_8431);
nand U9015 (N_9015,N_8965,N_8492);
nor U9016 (N_9016,N_8204,N_8886);
xnor U9017 (N_9017,N_8709,N_8920);
and U9018 (N_9018,N_8022,N_8110);
and U9019 (N_9019,N_8612,N_8254);
nor U9020 (N_9020,N_8523,N_8386);
and U9021 (N_9021,N_8640,N_8184);
nand U9022 (N_9022,N_8701,N_8181);
nand U9023 (N_9023,N_8360,N_8272);
nor U9024 (N_9024,N_8105,N_8750);
nor U9025 (N_9025,N_8190,N_8076);
nand U9026 (N_9026,N_8529,N_8252);
and U9027 (N_9027,N_8978,N_8852);
or U9028 (N_9028,N_8747,N_8446);
and U9029 (N_9029,N_8824,N_8927);
or U9030 (N_9030,N_8840,N_8939);
nor U9031 (N_9031,N_8343,N_8394);
and U9032 (N_9032,N_8687,N_8909);
and U9033 (N_9033,N_8719,N_8525);
nor U9034 (N_9034,N_8361,N_8816);
or U9035 (N_9035,N_8877,N_8844);
or U9036 (N_9036,N_8785,N_8057);
nand U9037 (N_9037,N_8042,N_8260);
and U9038 (N_9038,N_8398,N_8273);
xnor U9039 (N_9039,N_8863,N_8600);
or U9040 (N_9040,N_8702,N_8085);
nand U9041 (N_9041,N_8677,N_8552);
xnor U9042 (N_9042,N_8622,N_8783);
and U9043 (N_9043,N_8207,N_8591);
nand U9044 (N_9044,N_8756,N_8746);
xnor U9045 (N_9045,N_8822,N_8292);
nand U9046 (N_9046,N_8545,N_8151);
xnor U9047 (N_9047,N_8299,N_8019);
nor U9048 (N_9048,N_8325,N_8045);
and U9049 (N_9049,N_8013,N_8145);
nand U9050 (N_9050,N_8220,N_8811);
xor U9051 (N_9051,N_8761,N_8699);
nand U9052 (N_9052,N_8407,N_8499);
and U9053 (N_9053,N_8109,N_8584);
xor U9054 (N_9054,N_8333,N_8708);
or U9055 (N_9055,N_8937,N_8037);
and U9056 (N_9056,N_8704,N_8946);
or U9057 (N_9057,N_8594,N_8808);
and U9058 (N_9058,N_8675,N_8486);
xnor U9059 (N_9059,N_8510,N_8236);
nor U9060 (N_9060,N_8757,N_8203);
xnor U9061 (N_9061,N_8847,N_8362);
xor U9062 (N_9062,N_8912,N_8268);
xor U9063 (N_9063,N_8957,N_8505);
xor U9064 (N_9064,N_8770,N_8030);
nor U9065 (N_9065,N_8794,N_8083);
nor U9066 (N_9066,N_8147,N_8780);
or U9067 (N_9067,N_8370,N_8348);
nand U9068 (N_9068,N_8763,N_8450);
xor U9069 (N_9069,N_8508,N_8357);
nor U9070 (N_9070,N_8933,N_8715);
xnor U9071 (N_9071,N_8396,N_8742);
nand U9072 (N_9072,N_8137,N_8784);
nor U9073 (N_9073,N_8623,N_8717);
and U9074 (N_9074,N_8438,N_8532);
nor U9075 (N_9075,N_8389,N_8314);
or U9076 (N_9076,N_8131,N_8981);
xor U9077 (N_9077,N_8405,N_8269);
nand U9078 (N_9078,N_8373,N_8259);
nand U9079 (N_9079,N_8164,N_8601);
or U9080 (N_9080,N_8494,N_8255);
xnor U9081 (N_9081,N_8974,N_8010);
nand U9082 (N_9082,N_8725,N_8179);
nor U9083 (N_9083,N_8634,N_8311);
nand U9084 (N_9084,N_8191,N_8614);
and U9085 (N_9085,N_8300,N_8200);
and U9086 (N_9086,N_8583,N_8691);
and U9087 (N_9087,N_8999,N_8310);
nor U9088 (N_9088,N_8592,N_8341);
or U9089 (N_9089,N_8960,N_8342);
nand U9090 (N_9090,N_8466,N_8654);
or U9091 (N_9091,N_8941,N_8376);
nor U9092 (N_9092,N_8703,N_8734);
or U9093 (N_9093,N_8293,N_8246);
xnor U9094 (N_9094,N_8497,N_8551);
nand U9095 (N_9095,N_8048,N_8970);
nand U9096 (N_9096,N_8520,N_8651);
or U9097 (N_9097,N_8738,N_8740);
nand U9098 (N_9098,N_8227,N_8706);
or U9099 (N_9099,N_8379,N_8673);
and U9100 (N_9100,N_8888,N_8091);
or U9101 (N_9101,N_8507,N_8636);
and U9102 (N_9102,N_8629,N_8152);
and U9103 (N_9103,N_8558,N_8180);
nand U9104 (N_9104,N_8445,N_8410);
nor U9105 (N_9105,N_8667,N_8657);
or U9106 (N_9106,N_8830,N_8873);
xnor U9107 (N_9107,N_8225,N_8842);
or U9108 (N_9108,N_8457,N_8149);
or U9109 (N_9109,N_8531,N_8158);
xor U9110 (N_9110,N_8161,N_8895);
nand U9111 (N_9111,N_8915,N_8890);
xnor U9112 (N_9112,N_8728,N_8201);
nand U9113 (N_9113,N_8579,N_8328);
and U9114 (N_9114,N_8274,N_8114);
xnor U9115 (N_9115,N_8662,N_8278);
or U9116 (N_9116,N_8332,N_8550);
nand U9117 (N_9117,N_8097,N_8723);
and U9118 (N_9118,N_8698,N_8034);
or U9119 (N_9119,N_8340,N_8012);
nand U9120 (N_9120,N_8779,N_8823);
or U9121 (N_9121,N_8819,N_8232);
or U9122 (N_9122,N_8365,N_8925);
xnor U9123 (N_9123,N_8914,N_8670);
and U9124 (N_9124,N_8366,N_8994);
nor U9125 (N_9125,N_8512,N_8442);
nand U9126 (N_9126,N_8380,N_8918);
and U9127 (N_9127,N_8422,N_8337);
or U9128 (N_9128,N_8081,N_8369);
and U9129 (N_9129,N_8305,N_8390);
or U9130 (N_9130,N_8408,N_8615);
nor U9131 (N_9131,N_8838,N_8006);
xnor U9132 (N_9132,N_8522,N_8788);
xnor U9133 (N_9133,N_8899,N_8007);
xnor U9134 (N_9134,N_8344,N_8904);
and U9135 (N_9135,N_8289,N_8118);
nand U9136 (N_9136,N_8774,N_8125);
nor U9137 (N_9137,N_8572,N_8940);
xor U9138 (N_9138,N_8047,N_8850);
nor U9139 (N_9139,N_8251,N_8593);
xor U9140 (N_9140,N_8606,N_8582);
xnor U9141 (N_9141,N_8475,N_8972);
nor U9142 (N_9142,N_8697,N_8597);
or U9143 (N_9143,N_8176,N_8777);
xnor U9144 (N_9144,N_8595,N_8247);
nand U9145 (N_9145,N_8477,N_8224);
nor U9146 (N_9146,N_8133,N_8991);
nand U9147 (N_9147,N_8711,N_8024);
nor U9148 (N_9148,N_8156,N_8196);
or U9149 (N_9149,N_8094,N_8542);
xor U9150 (N_9150,N_8077,N_8737);
nand U9151 (N_9151,N_8833,N_8067);
or U9152 (N_9152,N_8679,N_8144);
xor U9153 (N_9153,N_8182,N_8501);
or U9154 (N_9154,N_8996,N_8907);
nor U9155 (N_9155,N_8868,N_8172);
nand U9156 (N_9156,N_8900,N_8686);
xor U9157 (N_9157,N_8079,N_8568);
nand U9158 (N_9158,N_8910,N_8096);
xor U9159 (N_9159,N_8949,N_8120);
or U9160 (N_9160,N_8417,N_8605);
nor U9161 (N_9161,N_8767,N_8950);
nand U9162 (N_9162,N_8456,N_8535);
xor U9163 (N_9163,N_8163,N_8841);
and U9164 (N_9164,N_8620,N_8319);
nor U9165 (N_9165,N_8923,N_8626);
and U9166 (N_9166,N_8294,N_8449);
nand U9167 (N_9167,N_8813,N_8467);
nor U9168 (N_9168,N_8917,N_8547);
nand U9169 (N_9169,N_8906,N_8855);
and U9170 (N_9170,N_8088,N_8213);
nor U9171 (N_9171,N_8801,N_8335);
nor U9172 (N_9172,N_8036,N_8393);
nand U9173 (N_9173,N_8485,N_8800);
nand U9174 (N_9174,N_8652,N_8188);
or U9175 (N_9175,N_8284,N_8948);
nand U9176 (N_9176,N_8881,N_8316);
nor U9177 (N_9177,N_8643,N_8569);
nand U9178 (N_9178,N_8329,N_8303);
xnor U9179 (N_9179,N_8173,N_8954);
or U9180 (N_9180,N_8166,N_8549);
or U9181 (N_9181,N_8185,N_8039);
or U9182 (N_9182,N_8193,N_8372);
nand U9183 (N_9183,N_8488,N_8140);
or U9184 (N_9184,N_8425,N_8222);
and U9185 (N_9185,N_8321,N_8101);
and U9186 (N_9186,N_8753,N_8049);
nand U9187 (N_9187,N_8973,N_8645);
nor U9188 (N_9188,N_8435,N_8980);
nor U9189 (N_9189,N_8472,N_8257);
or U9190 (N_9190,N_8170,N_8155);
xnor U9191 (N_9191,N_8502,N_8413);
nor U9192 (N_9192,N_8587,N_8474);
and U9193 (N_9193,N_8384,N_8644);
nor U9194 (N_9194,N_8664,N_8471);
or U9195 (N_9195,N_8264,N_8689);
nand U9196 (N_9196,N_8235,N_8460);
nor U9197 (N_9197,N_8302,N_8849);
or U9198 (N_9198,N_8290,N_8955);
nor U9199 (N_9199,N_8952,N_8588);
and U9200 (N_9200,N_8573,N_8596);
or U9201 (N_9201,N_8866,N_8197);
xnor U9202 (N_9202,N_8397,N_8616);
and U9203 (N_9203,N_8848,N_8356);
nor U9204 (N_9204,N_8436,N_8967);
xor U9205 (N_9205,N_8861,N_8392);
xor U9206 (N_9206,N_8810,N_8355);
nand U9207 (N_9207,N_8619,N_8560);
xnor U9208 (N_9208,N_8743,N_8998);
nand U9209 (N_9209,N_8879,N_8003);
xor U9210 (N_9210,N_8404,N_8987);
nand U9211 (N_9211,N_8060,N_8237);
and U9212 (N_9212,N_8598,N_8997);
nor U9213 (N_9213,N_8099,N_8806);
or U9214 (N_9214,N_8688,N_8869);
xor U9215 (N_9215,N_8248,N_8381);
nor U9216 (N_9216,N_8832,N_8177);
and U9217 (N_9217,N_8005,N_8926);
nand U9218 (N_9218,N_8611,N_8403);
nor U9219 (N_9219,N_8282,N_8391);
nor U9220 (N_9220,N_8124,N_8827);
or U9221 (N_9221,N_8412,N_8214);
or U9222 (N_9222,N_8253,N_8115);
or U9223 (N_9223,N_8985,N_8496);
and U9224 (N_9224,N_8585,N_8969);
nand U9225 (N_9225,N_8347,N_8035);
xor U9226 (N_9226,N_8399,N_8901);
nand U9227 (N_9227,N_8986,N_8660);
or U9228 (N_9228,N_8938,N_8001);
xnor U9229 (N_9229,N_8336,N_8100);
and U9230 (N_9230,N_8054,N_8905);
nand U9231 (N_9231,N_8845,N_8561);
or U9232 (N_9232,N_8516,N_8279);
or U9233 (N_9233,N_8029,N_8424);
nand U9234 (N_9234,N_8724,N_8308);
or U9235 (N_9235,N_8484,N_8536);
xnor U9236 (N_9236,N_8198,N_8095);
nor U9237 (N_9237,N_8786,N_8052);
nor U9238 (N_9238,N_8678,N_8648);
or U9239 (N_9239,N_8898,N_8963);
xnor U9240 (N_9240,N_8004,N_8932);
xnor U9241 (N_9241,N_8971,N_8206);
or U9242 (N_9242,N_8186,N_8470);
and U9243 (N_9243,N_8807,N_8665);
nor U9244 (N_9244,N_8792,N_8132);
nand U9245 (N_9245,N_8880,N_8322);
or U9246 (N_9246,N_8127,N_8473);
or U9247 (N_9247,N_8882,N_8210);
and U9248 (N_9248,N_8086,N_8804);
and U9249 (N_9249,N_8872,N_8928);
or U9250 (N_9250,N_8762,N_8716);
or U9251 (N_9251,N_8576,N_8836);
nand U9252 (N_9252,N_8491,N_8682);
or U9253 (N_9253,N_8478,N_8515);
nor U9254 (N_9254,N_8065,N_8027);
and U9255 (N_9255,N_8553,N_8518);
and U9256 (N_9256,N_8102,N_8778);
xnor U9257 (N_9257,N_8621,N_8506);
nand U9258 (N_9258,N_8771,N_8538);
and U9259 (N_9259,N_8364,N_8128);
nor U9260 (N_9260,N_8043,N_8139);
nand U9261 (N_9261,N_8992,N_8878);
xnor U9262 (N_9262,N_8566,N_8243);
and U9263 (N_9263,N_8732,N_8630);
and U9264 (N_9264,N_8534,N_8736);
nor U9265 (N_9265,N_8080,N_8766);
xnor U9266 (N_9266,N_8526,N_8758);
or U9267 (N_9267,N_8489,N_8924);
or U9268 (N_9268,N_8072,N_8826);
nand U9269 (N_9269,N_8129,N_8929);
xor U9270 (N_9270,N_8382,N_8559);
or U9271 (N_9271,N_8681,N_8371);
xnor U9272 (N_9272,N_8312,N_8982);
and U9273 (N_9273,N_8481,N_8603);
or U9274 (N_9274,N_8150,N_8672);
nor U9275 (N_9275,N_8117,N_8363);
and U9276 (N_9276,N_8613,N_8874);
or U9277 (N_9277,N_8793,N_8749);
nor U9278 (N_9278,N_8638,N_8911);
xor U9279 (N_9279,N_8789,N_8820);
nor U9280 (N_9280,N_8834,N_8021);
nor U9281 (N_9281,N_8469,N_8221);
nand U9282 (N_9282,N_8483,N_8632);
nor U9283 (N_9283,N_8345,N_8423);
or U9284 (N_9284,N_8281,N_8782);
and U9285 (N_9285,N_8401,N_8142);
or U9286 (N_9286,N_8327,N_8189);
nand U9287 (N_9287,N_8452,N_8053);
nor U9288 (N_9288,N_8589,N_8238);
xnor U9289 (N_9289,N_8209,N_8764);
and U9290 (N_9290,N_8298,N_8217);
xnor U9291 (N_9291,N_8317,N_8429);
and U9292 (N_9292,N_8136,N_8964);
xor U9293 (N_9293,N_8635,N_8313);
nand U9294 (N_9294,N_8581,N_8416);
xnor U9295 (N_9295,N_8799,N_8258);
nand U9296 (N_9296,N_8871,N_8722);
nor U9297 (N_9297,N_8242,N_8829);
nor U9298 (N_9298,N_8627,N_8169);
xnor U9299 (N_9299,N_8647,N_8280);
nand U9300 (N_9300,N_8427,N_8479);
xnor U9301 (N_9301,N_8922,N_8628);
and U9302 (N_9302,N_8961,N_8183);
nand U9303 (N_9303,N_8414,N_8463);
or U9304 (N_9304,N_8631,N_8119);
xor U9305 (N_9305,N_8921,N_8979);
or U9306 (N_9306,N_8825,N_8509);
xor U9307 (N_9307,N_8465,N_8112);
nand U9308 (N_9308,N_8870,N_8032);
nand U9309 (N_9309,N_8070,N_8493);
or U9310 (N_9310,N_8187,N_8713);
nand U9311 (N_9311,N_8735,N_8266);
nand U9312 (N_9312,N_8751,N_8495);
or U9313 (N_9313,N_8887,N_8454);
nor U9314 (N_9314,N_8514,N_8517);
xor U9315 (N_9315,N_8519,N_8563);
or U9316 (N_9316,N_8544,N_8074);
xnor U9317 (N_9317,N_8026,N_8287);
nor U9318 (N_9318,N_8577,N_8226);
nor U9319 (N_9319,N_8705,N_8769);
or U9320 (N_9320,N_8618,N_8902);
or U9321 (N_9321,N_8707,N_8350);
nand U9322 (N_9322,N_8157,N_8234);
nor U9323 (N_9323,N_8543,N_8480);
nor U9324 (N_9324,N_8402,N_8138);
xnor U9325 (N_9325,N_8135,N_8942);
xor U9326 (N_9326,N_8375,N_8089);
and U9327 (N_9327,N_8276,N_8564);
and U9328 (N_9328,N_8153,N_8367);
nand U9329 (N_9329,N_8250,N_8050);
and U9330 (N_9330,N_8885,N_8659);
xnor U9331 (N_9331,N_8608,N_8590);
xor U9332 (N_9332,N_8528,N_8014);
nand U9333 (N_9333,N_8354,N_8913);
or U9334 (N_9334,N_8916,N_8339);
and U9335 (N_9335,N_8748,N_8646);
and U9336 (N_9336,N_8975,N_8263);
nor U9337 (N_9337,N_8451,N_8211);
xnor U9338 (N_9338,N_8388,N_8637);
or U9339 (N_9339,N_8854,N_8334);
xor U9340 (N_9340,N_8063,N_8061);
nor U9341 (N_9341,N_8720,N_8330);
or U9342 (N_9342,N_8649,N_8856);
xnor U9343 (N_9343,N_8448,N_8296);
and U9344 (N_9344,N_8984,N_8814);
nor U9345 (N_9345,N_8803,N_8817);
or U9346 (N_9346,N_8653,N_8033);
and U9347 (N_9347,N_8700,N_8775);
and U9348 (N_9348,N_8966,N_8378);
and U9349 (N_9349,N_8383,N_8462);
nand U9350 (N_9350,N_8565,N_8521);
xor U9351 (N_9351,N_8944,N_8106);
nand U9352 (N_9352,N_8741,N_8571);
and U9353 (N_9353,N_8798,N_8443);
or U9354 (N_9354,N_8092,N_8358);
and U9355 (N_9355,N_8192,N_8602);
xor U9356 (N_9356,N_8993,N_8230);
xor U9357 (N_9357,N_8374,N_8864);
nor U9358 (N_9358,N_8851,N_8530);
xor U9359 (N_9359,N_8418,N_8126);
xnor U9360 (N_9360,N_8945,N_8265);
nor U9361 (N_9361,N_8853,N_8831);
nor U9362 (N_9362,N_8241,N_8482);
xor U9363 (N_9363,N_8008,N_8580);
xor U9364 (N_9364,N_8476,N_8025);
nand U9365 (N_9365,N_8828,N_8148);
nand U9366 (N_9366,N_8017,N_8759);
nor U9367 (N_9367,N_8090,N_8216);
xnor U9368 (N_9368,N_8787,N_8256);
and U9369 (N_9369,N_8084,N_8586);
and U9370 (N_9370,N_8160,N_8837);
and U9371 (N_9371,N_8893,N_8351);
nand U9372 (N_9372,N_8858,N_8455);
xor U9373 (N_9373,N_8123,N_8656);
nor U9374 (N_9374,N_8641,N_8406);
xnor U9375 (N_9375,N_8875,N_8889);
and U9376 (N_9376,N_8275,N_8306);
xor U9377 (N_9377,N_8894,N_8068);
nand U9378 (N_9378,N_8320,N_8240);
or U9379 (N_9379,N_8231,N_8812);
xnor U9380 (N_9380,N_8130,N_8745);
nor U9381 (N_9381,N_8233,N_8323);
xnor U9382 (N_9382,N_8051,N_8415);
and U9383 (N_9383,N_8903,N_8002);
and U9384 (N_9384,N_8020,N_8567);
nor U9385 (N_9385,N_8228,N_8122);
nand U9386 (N_9386,N_8988,N_8633);
nand U9387 (N_9387,N_8781,N_8693);
and U9388 (N_9388,N_8434,N_8865);
or U9389 (N_9389,N_8726,N_8556);
xor U9390 (N_9390,N_8562,N_8797);
and U9391 (N_9391,N_8555,N_8023);
and U9392 (N_9392,N_8503,N_8073);
xor U9393 (N_9393,N_8040,N_8795);
and U9394 (N_9394,N_8892,N_8338);
xor U9395 (N_9395,N_8609,N_8162);
nand U9396 (N_9396,N_8428,N_8353);
or U9397 (N_9397,N_8546,N_8307);
and U9398 (N_9398,N_8041,N_8078);
nor U9399 (N_9399,N_8729,N_8419);
nand U9400 (N_9400,N_8395,N_8599);
nand U9401 (N_9401,N_8669,N_8459);
and U9402 (N_9402,N_8349,N_8727);
xnor U9403 (N_9403,N_8857,N_8818);
and U9404 (N_9404,N_8297,N_8695);
or U9405 (N_9405,N_8666,N_8426);
or U9406 (N_9406,N_8055,N_8069);
nand U9407 (N_9407,N_8058,N_8977);
or U9408 (N_9408,N_8291,N_8121);
nor U9409 (N_9409,N_8066,N_8286);
xor U9410 (N_9410,N_8642,N_8624);
and U9411 (N_9411,N_8896,N_8285);
and U9412 (N_9412,N_8490,N_8658);
or U9413 (N_9413,N_8958,N_8674);
nand U9414 (N_9414,N_8540,N_8575);
xor U9415 (N_9415,N_8301,N_8934);
xor U9416 (N_9416,N_8432,N_8765);
or U9417 (N_9417,N_8731,N_8000);
xnor U9418 (N_9418,N_8326,N_8352);
xnor U9419 (N_9419,N_8663,N_8790);
nor U9420 (N_9420,N_8721,N_8018);
xor U9421 (N_9421,N_8315,N_8574);
xor U9422 (N_9422,N_8271,N_8989);
nand U9423 (N_9423,N_8175,N_8968);
nand U9424 (N_9424,N_8098,N_8249);
and U9425 (N_9425,N_8692,N_8433);
nor U9426 (N_9426,N_8146,N_8208);
and U9427 (N_9427,N_8439,N_8059);
and U9428 (N_9428,N_8815,N_8668);
nor U9429 (N_9429,N_8859,N_8103);
nor U9430 (N_9430,N_8557,N_8195);
and U9431 (N_9431,N_8650,N_8219);
nand U9432 (N_9432,N_8441,N_8500);
and U9433 (N_9433,N_8661,N_8809);
or U9434 (N_9434,N_8331,N_8205);
xor U9435 (N_9435,N_8458,N_8548);
xor U9436 (N_9436,N_8377,N_8283);
and U9437 (N_9437,N_8016,N_8318);
and U9438 (N_9438,N_8539,N_8862);
nand U9439 (N_9439,N_8064,N_8821);
or U9440 (N_9440,N_8229,N_8487);
xnor U9441 (N_9441,N_8168,N_8400);
xor U9442 (N_9442,N_8009,N_8421);
xnor U9443 (N_9443,N_8908,N_8430);
and U9444 (N_9444,N_8143,N_8712);
or U9445 (N_9445,N_8839,N_8277);
and U9446 (N_9446,N_8420,N_8846);
nor U9447 (N_9447,N_8883,N_8154);
nand U9448 (N_9448,N_8159,N_8093);
nand U9449 (N_9449,N_8931,N_8447);
or U9450 (N_9450,N_8245,N_8680);
or U9451 (N_9451,N_8730,N_8607);
xor U9452 (N_9452,N_8639,N_8690);
xor U9453 (N_9453,N_8953,N_8990);
and U9454 (N_9454,N_8760,N_8511);
nand U9455 (N_9455,N_8776,N_8167);
or U9456 (N_9456,N_8891,N_8304);
xor U9457 (N_9457,N_8676,N_8504);
xor U9458 (N_9458,N_8134,N_8387);
xnor U9459 (N_9459,N_8223,N_8768);
nor U9460 (N_9460,N_8141,N_8976);
xor U9461 (N_9461,N_8570,N_8031);
nand U9462 (N_9462,N_8604,N_8995);
xnor U9463 (N_9463,N_8773,N_8111);
or U9464 (N_9464,N_8625,N_8791);
xnor U9465 (N_9465,N_8610,N_8409);
nor U9466 (N_9466,N_8461,N_8075);
or U9467 (N_9467,N_8876,N_8513);
or U9468 (N_9468,N_8261,N_8802);
nand U9469 (N_9469,N_8527,N_8919);
and U9470 (N_9470,N_8239,N_8165);
xnor U9471 (N_9471,N_8385,N_8464);
and U9472 (N_9472,N_8843,N_8744);
nand U9473 (N_9473,N_8270,N_8951);
nand U9474 (N_9474,N_8860,N_8444);
or U9475 (N_9475,N_8671,N_8295);
and U9476 (N_9476,N_8244,N_8411);
nor U9477 (N_9477,N_8696,N_8947);
or U9478 (N_9478,N_8288,N_8685);
nor U9479 (N_9479,N_8694,N_8739);
or U9480 (N_9480,N_8498,N_8796);
nor U9481 (N_9481,N_8262,N_8171);
nand U9482 (N_9482,N_8218,N_8772);
nor U9483 (N_9483,N_8194,N_8983);
nor U9484 (N_9484,N_8267,N_8935);
and U9485 (N_9485,N_8113,N_8655);
nor U9486 (N_9486,N_8104,N_8962);
and U9487 (N_9487,N_8956,N_8554);
nand U9488 (N_9488,N_8071,N_8440);
xor U9489 (N_9489,N_8718,N_8199);
or U9490 (N_9490,N_8617,N_8453);
nand U9491 (N_9491,N_8082,N_8202);
or U9492 (N_9492,N_8578,N_8108);
xnor U9493 (N_9493,N_8468,N_8178);
nand U9494 (N_9494,N_8805,N_8107);
nor U9495 (N_9495,N_8212,N_8215);
and U9496 (N_9496,N_8884,N_8835);
nor U9497 (N_9497,N_8524,N_8015);
xor U9498 (N_9498,N_8930,N_8087);
or U9499 (N_9499,N_8684,N_8897);
and U9500 (N_9500,N_8188,N_8078);
nand U9501 (N_9501,N_8194,N_8145);
nor U9502 (N_9502,N_8008,N_8028);
or U9503 (N_9503,N_8712,N_8710);
nor U9504 (N_9504,N_8191,N_8538);
and U9505 (N_9505,N_8763,N_8941);
or U9506 (N_9506,N_8910,N_8941);
and U9507 (N_9507,N_8688,N_8342);
nand U9508 (N_9508,N_8041,N_8612);
and U9509 (N_9509,N_8938,N_8670);
xnor U9510 (N_9510,N_8478,N_8075);
nand U9511 (N_9511,N_8240,N_8290);
nor U9512 (N_9512,N_8633,N_8926);
and U9513 (N_9513,N_8096,N_8757);
or U9514 (N_9514,N_8776,N_8367);
nand U9515 (N_9515,N_8105,N_8066);
nand U9516 (N_9516,N_8760,N_8718);
and U9517 (N_9517,N_8061,N_8806);
nor U9518 (N_9518,N_8911,N_8880);
or U9519 (N_9519,N_8532,N_8919);
and U9520 (N_9520,N_8295,N_8725);
and U9521 (N_9521,N_8677,N_8740);
or U9522 (N_9522,N_8090,N_8823);
nor U9523 (N_9523,N_8411,N_8956);
nand U9524 (N_9524,N_8150,N_8589);
xnor U9525 (N_9525,N_8625,N_8872);
or U9526 (N_9526,N_8401,N_8654);
nand U9527 (N_9527,N_8987,N_8298);
and U9528 (N_9528,N_8372,N_8811);
or U9529 (N_9529,N_8696,N_8484);
or U9530 (N_9530,N_8076,N_8539);
nand U9531 (N_9531,N_8327,N_8029);
and U9532 (N_9532,N_8258,N_8241);
nand U9533 (N_9533,N_8121,N_8631);
nand U9534 (N_9534,N_8544,N_8193);
nand U9535 (N_9535,N_8619,N_8089);
nand U9536 (N_9536,N_8480,N_8386);
nor U9537 (N_9537,N_8227,N_8493);
nor U9538 (N_9538,N_8069,N_8287);
or U9539 (N_9539,N_8702,N_8470);
nor U9540 (N_9540,N_8124,N_8763);
nand U9541 (N_9541,N_8080,N_8932);
nand U9542 (N_9542,N_8811,N_8080);
xnor U9543 (N_9543,N_8827,N_8365);
and U9544 (N_9544,N_8780,N_8943);
and U9545 (N_9545,N_8845,N_8710);
and U9546 (N_9546,N_8205,N_8032);
nor U9547 (N_9547,N_8901,N_8423);
nor U9548 (N_9548,N_8682,N_8552);
and U9549 (N_9549,N_8944,N_8641);
nor U9550 (N_9550,N_8756,N_8444);
xor U9551 (N_9551,N_8074,N_8884);
nor U9552 (N_9552,N_8983,N_8662);
nor U9553 (N_9553,N_8326,N_8251);
xor U9554 (N_9554,N_8940,N_8369);
and U9555 (N_9555,N_8736,N_8016);
and U9556 (N_9556,N_8948,N_8038);
and U9557 (N_9557,N_8567,N_8441);
and U9558 (N_9558,N_8811,N_8825);
and U9559 (N_9559,N_8591,N_8235);
or U9560 (N_9560,N_8389,N_8239);
and U9561 (N_9561,N_8021,N_8941);
nor U9562 (N_9562,N_8911,N_8820);
and U9563 (N_9563,N_8643,N_8435);
or U9564 (N_9564,N_8289,N_8111);
nor U9565 (N_9565,N_8829,N_8284);
or U9566 (N_9566,N_8281,N_8849);
nand U9567 (N_9567,N_8015,N_8395);
or U9568 (N_9568,N_8106,N_8103);
xor U9569 (N_9569,N_8222,N_8752);
nor U9570 (N_9570,N_8806,N_8317);
or U9571 (N_9571,N_8028,N_8750);
or U9572 (N_9572,N_8393,N_8207);
or U9573 (N_9573,N_8341,N_8958);
and U9574 (N_9574,N_8158,N_8274);
or U9575 (N_9575,N_8809,N_8122);
or U9576 (N_9576,N_8479,N_8565);
xnor U9577 (N_9577,N_8676,N_8944);
or U9578 (N_9578,N_8635,N_8955);
nand U9579 (N_9579,N_8300,N_8844);
and U9580 (N_9580,N_8964,N_8140);
xnor U9581 (N_9581,N_8911,N_8096);
xnor U9582 (N_9582,N_8607,N_8188);
and U9583 (N_9583,N_8492,N_8914);
nand U9584 (N_9584,N_8747,N_8418);
nand U9585 (N_9585,N_8571,N_8809);
and U9586 (N_9586,N_8361,N_8977);
and U9587 (N_9587,N_8313,N_8181);
nand U9588 (N_9588,N_8169,N_8781);
or U9589 (N_9589,N_8250,N_8277);
nand U9590 (N_9590,N_8052,N_8971);
nor U9591 (N_9591,N_8465,N_8491);
nor U9592 (N_9592,N_8448,N_8754);
nor U9593 (N_9593,N_8443,N_8049);
xor U9594 (N_9594,N_8880,N_8268);
or U9595 (N_9595,N_8414,N_8882);
xor U9596 (N_9596,N_8941,N_8658);
nand U9597 (N_9597,N_8113,N_8106);
or U9598 (N_9598,N_8274,N_8521);
nor U9599 (N_9599,N_8612,N_8851);
or U9600 (N_9600,N_8642,N_8675);
and U9601 (N_9601,N_8652,N_8887);
nor U9602 (N_9602,N_8063,N_8799);
or U9603 (N_9603,N_8010,N_8101);
xnor U9604 (N_9604,N_8232,N_8218);
or U9605 (N_9605,N_8026,N_8812);
nand U9606 (N_9606,N_8499,N_8035);
xor U9607 (N_9607,N_8251,N_8991);
nor U9608 (N_9608,N_8915,N_8452);
nor U9609 (N_9609,N_8266,N_8721);
nand U9610 (N_9610,N_8624,N_8448);
xnor U9611 (N_9611,N_8380,N_8959);
or U9612 (N_9612,N_8386,N_8928);
nor U9613 (N_9613,N_8676,N_8765);
or U9614 (N_9614,N_8716,N_8234);
and U9615 (N_9615,N_8839,N_8942);
nand U9616 (N_9616,N_8671,N_8501);
and U9617 (N_9617,N_8855,N_8375);
nor U9618 (N_9618,N_8226,N_8158);
nand U9619 (N_9619,N_8207,N_8215);
and U9620 (N_9620,N_8274,N_8566);
xor U9621 (N_9621,N_8970,N_8386);
and U9622 (N_9622,N_8412,N_8024);
xnor U9623 (N_9623,N_8338,N_8861);
or U9624 (N_9624,N_8762,N_8267);
or U9625 (N_9625,N_8509,N_8796);
xor U9626 (N_9626,N_8214,N_8594);
or U9627 (N_9627,N_8027,N_8522);
nor U9628 (N_9628,N_8911,N_8734);
or U9629 (N_9629,N_8913,N_8489);
nand U9630 (N_9630,N_8979,N_8124);
nand U9631 (N_9631,N_8654,N_8305);
or U9632 (N_9632,N_8175,N_8228);
nand U9633 (N_9633,N_8760,N_8568);
nor U9634 (N_9634,N_8116,N_8982);
and U9635 (N_9635,N_8888,N_8765);
or U9636 (N_9636,N_8135,N_8069);
xor U9637 (N_9637,N_8704,N_8971);
and U9638 (N_9638,N_8519,N_8998);
nand U9639 (N_9639,N_8603,N_8228);
xnor U9640 (N_9640,N_8581,N_8502);
xnor U9641 (N_9641,N_8110,N_8807);
nor U9642 (N_9642,N_8833,N_8108);
or U9643 (N_9643,N_8720,N_8323);
nor U9644 (N_9644,N_8096,N_8255);
nor U9645 (N_9645,N_8685,N_8995);
and U9646 (N_9646,N_8270,N_8388);
nand U9647 (N_9647,N_8686,N_8161);
and U9648 (N_9648,N_8255,N_8849);
nand U9649 (N_9649,N_8218,N_8617);
xor U9650 (N_9650,N_8143,N_8088);
nor U9651 (N_9651,N_8423,N_8600);
or U9652 (N_9652,N_8535,N_8513);
nor U9653 (N_9653,N_8598,N_8687);
xnor U9654 (N_9654,N_8404,N_8979);
or U9655 (N_9655,N_8770,N_8725);
and U9656 (N_9656,N_8716,N_8939);
and U9657 (N_9657,N_8120,N_8817);
nand U9658 (N_9658,N_8081,N_8598);
or U9659 (N_9659,N_8176,N_8112);
nor U9660 (N_9660,N_8880,N_8366);
nor U9661 (N_9661,N_8913,N_8171);
xnor U9662 (N_9662,N_8570,N_8503);
nand U9663 (N_9663,N_8617,N_8299);
nand U9664 (N_9664,N_8747,N_8110);
nand U9665 (N_9665,N_8977,N_8031);
xor U9666 (N_9666,N_8721,N_8775);
xor U9667 (N_9667,N_8893,N_8276);
nand U9668 (N_9668,N_8138,N_8267);
and U9669 (N_9669,N_8322,N_8153);
nand U9670 (N_9670,N_8600,N_8750);
nor U9671 (N_9671,N_8294,N_8328);
or U9672 (N_9672,N_8459,N_8478);
nor U9673 (N_9673,N_8785,N_8562);
or U9674 (N_9674,N_8086,N_8039);
nand U9675 (N_9675,N_8786,N_8943);
nand U9676 (N_9676,N_8255,N_8372);
nand U9677 (N_9677,N_8919,N_8893);
or U9678 (N_9678,N_8677,N_8520);
or U9679 (N_9679,N_8698,N_8707);
nand U9680 (N_9680,N_8209,N_8131);
nor U9681 (N_9681,N_8139,N_8652);
nor U9682 (N_9682,N_8598,N_8143);
nor U9683 (N_9683,N_8012,N_8487);
or U9684 (N_9684,N_8660,N_8298);
and U9685 (N_9685,N_8669,N_8038);
nand U9686 (N_9686,N_8657,N_8537);
nand U9687 (N_9687,N_8646,N_8854);
or U9688 (N_9688,N_8036,N_8471);
or U9689 (N_9689,N_8605,N_8296);
nand U9690 (N_9690,N_8217,N_8906);
nor U9691 (N_9691,N_8317,N_8183);
or U9692 (N_9692,N_8143,N_8993);
nand U9693 (N_9693,N_8671,N_8320);
and U9694 (N_9694,N_8425,N_8713);
and U9695 (N_9695,N_8487,N_8582);
nand U9696 (N_9696,N_8497,N_8498);
xor U9697 (N_9697,N_8333,N_8121);
or U9698 (N_9698,N_8267,N_8818);
nand U9699 (N_9699,N_8998,N_8556);
nand U9700 (N_9700,N_8702,N_8292);
and U9701 (N_9701,N_8907,N_8052);
xor U9702 (N_9702,N_8949,N_8924);
nand U9703 (N_9703,N_8817,N_8380);
nor U9704 (N_9704,N_8642,N_8250);
or U9705 (N_9705,N_8837,N_8913);
nand U9706 (N_9706,N_8746,N_8935);
and U9707 (N_9707,N_8782,N_8992);
and U9708 (N_9708,N_8974,N_8033);
and U9709 (N_9709,N_8682,N_8613);
nand U9710 (N_9710,N_8481,N_8208);
xnor U9711 (N_9711,N_8589,N_8392);
nor U9712 (N_9712,N_8766,N_8426);
or U9713 (N_9713,N_8225,N_8603);
or U9714 (N_9714,N_8804,N_8508);
xor U9715 (N_9715,N_8737,N_8901);
or U9716 (N_9716,N_8407,N_8552);
and U9717 (N_9717,N_8759,N_8533);
nor U9718 (N_9718,N_8669,N_8722);
or U9719 (N_9719,N_8774,N_8607);
and U9720 (N_9720,N_8180,N_8961);
and U9721 (N_9721,N_8930,N_8819);
and U9722 (N_9722,N_8461,N_8164);
nand U9723 (N_9723,N_8701,N_8856);
nand U9724 (N_9724,N_8131,N_8588);
nand U9725 (N_9725,N_8727,N_8766);
and U9726 (N_9726,N_8353,N_8352);
nor U9727 (N_9727,N_8845,N_8292);
nor U9728 (N_9728,N_8767,N_8155);
or U9729 (N_9729,N_8756,N_8191);
or U9730 (N_9730,N_8483,N_8924);
and U9731 (N_9731,N_8582,N_8675);
and U9732 (N_9732,N_8186,N_8058);
nand U9733 (N_9733,N_8132,N_8710);
xnor U9734 (N_9734,N_8617,N_8393);
nand U9735 (N_9735,N_8549,N_8011);
xnor U9736 (N_9736,N_8684,N_8827);
or U9737 (N_9737,N_8936,N_8567);
xnor U9738 (N_9738,N_8007,N_8639);
xor U9739 (N_9739,N_8205,N_8459);
or U9740 (N_9740,N_8452,N_8575);
xnor U9741 (N_9741,N_8345,N_8432);
xor U9742 (N_9742,N_8064,N_8908);
and U9743 (N_9743,N_8101,N_8330);
nand U9744 (N_9744,N_8575,N_8743);
xor U9745 (N_9745,N_8895,N_8967);
nor U9746 (N_9746,N_8911,N_8077);
or U9747 (N_9747,N_8869,N_8022);
nand U9748 (N_9748,N_8055,N_8841);
nand U9749 (N_9749,N_8805,N_8097);
nand U9750 (N_9750,N_8170,N_8725);
and U9751 (N_9751,N_8649,N_8713);
and U9752 (N_9752,N_8406,N_8127);
nor U9753 (N_9753,N_8340,N_8859);
xor U9754 (N_9754,N_8204,N_8505);
or U9755 (N_9755,N_8265,N_8317);
and U9756 (N_9756,N_8311,N_8678);
or U9757 (N_9757,N_8350,N_8274);
or U9758 (N_9758,N_8015,N_8618);
nand U9759 (N_9759,N_8954,N_8433);
nor U9760 (N_9760,N_8914,N_8582);
or U9761 (N_9761,N_8856,N_8616);
nand U9762 (N_9762,N_8774,N_8446);
xnor U9763 (N_9763,N_8677,N_8195);
nor U9764 (N_9764,N_8804,N_8029);
xnor U9765 (N_9765,N_8213,N_8005);
and U9766 (N_9766,N_8842,N_8038);
or U9767 (N_9767,N_8586,N_8711);
or U9768 (N_9768,N_8396,N_8088);
and U9769 (N_9769,N_8883,N_8250);
xnor U9770 (N_9770,N_8786,N_8398);
xnor U9771 (N_9771,N_8574,N_8742);
xor U9772 (N_9772,N_8639,N_8256);
xnor U9773 (N_9773,N_8519,N_8277);
and U9774 (N_9774,N_8374,N_8534);
and U9775 (N_9775,N_8033,N_8236);
and U9776 (N_9776,N_8520,N_8675);
nand U9777 (N_9777,N_8651,N_8974);
and U9778 (N_9778,N_8445,N_8408);
nor U9779 (N_9779,N_8771,N_8199);
xnor U9780 (N_9780,N_8908,N_8542);
or U9781 (N_9781,N_8759,N_8961);
and U9782 (N_9782,N_8971,N_8188);
nand U9783 (N_9783,N_8290,N_8186);
xnor U9784 (N_9784,N_8280,N_8551);
and U9785 (N_9785,N_8049,N_8995);
and U9786 (N_9786,N_8717,N_8528);
or U9787 (N_9787,N_8393,N_8328);
nor U9788 (N_9788,N_8723,N_8193);
nand U9789 (N_9789,N_8621,N_8148);
xor U9790 (N_9790,N_8210,N_8266);
and U9791 (N_9791,N_8379,N_8689);
and U9792 (N_9792,N_8097,N_8574);
nor U9793 (N_9793,N_8337,N_8233);
nor U9794 (N_9794,N_8799,N_8903);
or U9795 (N_9795,N_8805,N_8334);
nor U9796 (N_9796,N_8869,N_8648);
nor U9797 (N_9797,N_8644,N_8457);
nor U9798 (N_9798,N_8163,N_8936);
nor U9799 (N_9799,N_8483,N_8063);
and U9800 (N_9800,N_8239,N_8632);
nand U9801 (N_9801,N_8140,N_8623);
xor U9802 (N_9802,N_8594,N_8957);
or U9803 (N_9803,N_8301,N_8368);
nand U9804 (N_9804,N_8756,N_8369);
nor U9805 (N_9805,N_8884,N_8420);
or U9806 (N_9806,N_8183,N_8605);
nand U9807 (N_9807,N_8013,N_8928);
and U9808 (N_9808,N_8982,N_8801);
nand U9809 (N_9809,N_8088,N_8933);
xor U9810 (N_9810,N_8609,N_8021);
nor U9811 (N_9811,N_8683,N_8675);
xnor U9812 (N_9812,N_8319,N_8668);
and U9813 (N_9813,N_8753,N_8687);
nor U9814 (N_9814,N_8052,N_8152);
nor U9815 (N_9815,N_8428,N_8153);
or U9816 (N_9816,N_8260,N_8772);
and U9817 (N_9817,N_8466,N_8642);
and U9818 (N_9818,N_8993,N_8375);
and U9819 (N_9819,N_8478,N_8518);
or U9820 (N_9820,N_8920,N_8921);
or U9821 (N_9821,N_8979,N_8496);
nor U9822 (N_9822,N_8368,N_8438);
and U9823 (N_9823,N_8237,N_8558);
xor U9824 (N_9824,N_8160,N_8667);
xnor U9825 (N_9825,N_8594,N_8806);
xor U9826 (N_9826,N_8567,N_8311);
and U9827 (N_9827,N_8006,N_8173);
and U9828 (N_9828,N_8545,N_8383);
and U9829 (N_9829,N_8547,N_8132);
and U9830 (N_9830,N_8246,N_8985);
nand U9831 (N_9831,N_8242,N_8409);
xnor U9832 (N_9832,N_8118,N_8067);
nand U9833 (N_9833,N_8727,N_8649);
nand U9834 (N_9834,N_8954,N_8221);
xor U9835 (N_9835,N_8778,N_8041);
nor U9836 (N_9836,N_8860,N_8661);
or U9837 (N_9837,N_8766,N_8831);
nand U9838 (N_9838,N_8267,N_8585);
and U9839 (N_9839,N_8275,N_8763);
nand U9840 (N_9840,N_8008,N_8932);
and U9841 (N_9841,N_8102,N_8723);
xor U9842 (N_9842,N_8242,N_8092);
xnor U9843 (N_9843,N_8171,N_8218);
nand U9844 (N_9844,N_8746,N_8572);
nor U9845 (N_9845,N_8456,N_8319);
nand U9846 (N_9846,N_8957,N_8411);
nand U9847 (N_9847,N_8376,N_8351);
nor U9848 (N_9848,N_8189,N_8344);
xor U9849 (N_9849,N_8913,N_8955);
nor U9850 (N_9850,N_8981,N_8089);
nor U9851 (N_9851,N_8911,N_8813);
or U9852 (N_9852,N_8906,N_8241);
xnor U9853 (N_9853,N_8368,N_8065);
and U9854 (N_9854,N_8763,N_8230);
or U9855 (N_9855,N_8398,N_8034);
xor U9856 (N_9856,N_8064,N_8805);
nor U9857 (N_9857,N_8631,N_8003);
xnor U9858 (N_9858,N_8717,N_8081);
or U9859 (N_9859,N_8617,N_8473);
nor U9860 (N_9860,N_8402,N_8730);
nand U9861 (N_9861,N_8026,N_8107);
xnor U9862 (N_9862,N_8710,N_8428);
nand U9863 (N_9863,N_8181,N_8020);
xor U9864 (N_9864,N_8978,N_8900);
nand U9865 (N_9865,N_8151,N_8645);
nor U9866 (N_9866,N_8688,N_8576);
or U9867 (N_9867,N_8022,N_8456);
nor U9868 (N_9868,N_8810,N_8100);
or U9869 (N_9869,N_8891,N_8720);
nor U9870 (N_9870,N_8011,N_8486);
nor U9871 (N_9871,N_8304,N_8461);
nor U9872 (N_9872,N_8362,N_8828);
nand U9873 (N_9873,N_8999,N_8273);
and U9874 (N_9874,N_8695,N_8560);
and U9875 (N_9875,N_8266,N_8246);
or U9876 (N_9876,N_8622,N_8374);
nor U9877 (N_9877,N_8055,N_8540);
nand U9878 (N_9878,N_8033,N_8432);
nand U9879 (N_9879,N_8949,N_8938);
and U9880 (N_9880,N_8971,N_8844);
nor U9881 (N_9881,N_8577,N_8996);
and U9882 (N_9882,N_8780,N_8145);
xnor U9883 (N_9883,N_8135,N_8155);
xor U9884 (N_9884,N_8709,N_8671);
or U9885 (N_9885,N_8062,N_8301);
and U9886 (N_9886,N_8437,N_8577);
xnor U9887 (N_9887,N_8940,N_8899);
nor U9888 (N_9888,N_8636,N_8999);
nand U9889 (N_9889,N_8676,N_8725);
or U9890 (N_9890,N_8135,N_8208);
xor U9891 (N_9891,N_8485,N_8278);
and U9892 (N_9892,N_8423,N_8673);
and U9893 (N_9893,N_8640,N_8509);
nand U9894 (N_9894,N_8568,N_8525);
or U9895 (N_9895,N_8984,N_8435);
xnor U9896 (N_9896,N_8672,N_8048);
xnor U9897 (N_9897,N_8754,N_8112);
nor U9898 (N_9898,N_8026,N_8509);
nor U9899 (N_9899,N_8103,N_8263);
nor U9900 (N_9900,N_8818,N_8678);
nand U9901 (N_9901,N_8961,N_8700);
or U9902 (N_9902,N_8436,N_8248);
nand U9903 (N_9903,N_8423,N_8447);
xor U9904 (N_9904,N_8819,N_8024);
nor U9905 (N_9905,N_8454,N_8778);
nand U9906 (N_9906,N_8116,N_8328);
or U9907 (N_9907,N_8575,N_8591);
or U9908 (N_9908,N_8413,N_8254);
nand U9909 (N_9909,N_8802,N_8502);
or U9910 (N_9910,N_8513,N_8595);
and U9911 (N_9911,N_8654,N_8504);
xnor U9912 (N_9912,N_8263,N_8993);
nor U9913 (N_9913,N_8175,N_8138);
nor U9914 (N_9914,N_8367,N_8444);
or U9915 (N_9915,N_8952,N_8734);
or U9916 (N_9916,N_8436,N_8077);
xor U9917 (N_9917,N_8200,N_8320);
or U9918 (N_9918,N_8534,N_8678);
nand U9919 (N_9919,N_8640,N_8117);
and U9920 (N_9920,N_8548,N_8304);
nor U9921 (N_9921,N_8377,N_8201);
and U9922 (N_9922,N_8047,N_8129);
or U9923 (N_9923,N_8445,N_8647);
xor U9924 (N_9924,N_8445,N_8029);
nand U9925 (N_9925,N_8843,N_8368);
and U9926 (N_9926,N_8726,N_8359);
xor U9927 (N_9927,N_8079,N_8726);
nor U9928 (N_9928,N_8914,N_8613);
or U9929 (N_9929,N_8339,N_8991);
or U9930 (N_9930,N_8839,N_8382);
and U9931 (N_9931,N_8084,N_8499);
or U9932 (N_9932,N_8476,N_8387);
nor U9933 (N_9933,N_8764,N_8487);
and U9934 (N_9934,N_8991,N_8343);
nand U9935 (N_9935,N_8564,N_8335);
xor U9936 (N_9936,N_8349,N_8280);
xor U9937 (N_9937,N_8999,N_8563);
nand U9938 (N_9938,N_8989,N_8847);
xor U9939 (N_9939,N_8698,N_8464);
nor U9940 (N_9940,N_8018,N_8782);
xor U9941 (N_9941,N_8984,N_8024);
nor U9942 (N_9942,N_8072,N_8631);
nand U9943 (N_9943,N_8427,N_8191);
xnor U9944 (N_9944,N_8510,N_8225);
nand U9945 (N_9945,N_8919,N_8607);
xnor U9946 (N_9946,N_8902,N_8468);
and U9947 (N_9947,N_8482,N_8999);
xor U9948 (N_9948,N_8667,N_8241);
nor U9949 (N_9949,N_8721,N_8357);
nor U9950 (N_9950,N_8359,N_8905);
xor U9951 (N_9951,N_8746,N_8905);
or U9952 (N_9952,N_8737,N_8741);
xor U9953 (N_9953,N_8907,N_8422);
or U9954 (N_9954,N_8365,N_8631);
or U9955 (N_9955,N_8267,N_8798);
nand U9956 (N_9956,N_8193,N_8931);
nor U9957 (N_9957,N_8557,N_8154);
nor U9958 (N_9958,N_8228,N_8649);
nand U9959 (N_9959,N_8171,N_8115);
nor U9960 (N_9960,N_8978,N_8120);
nor U9961 (N_9961,N_8317,N_8815);
nor U9962 (N_9962,N_8953,N_8357);
nor U9963 (N_9963,N_8906,N_8717);
xor U9964 (N_9964,N_8791,N_8258);
xnor U9965 (N_9965,N_8512,N_8549);
and U9966 (N_9966,N_8125,N_8228);
nor U9967 (N_9967,N_8971,N_8135);
and U9968 (N_9968,N_8795,N_8339);
nor U9969 (N_9969,N_8619,N_8555);
xor U9970 (N_9970,N_8974,N_8396);
nor U9971 (N_9971,N_8237,N_8743);
xor U9972 (N_9972,N_8156,N_8617);
nor U9973 (N_9973,N_8133,N_8841);
and U9974 (N_9974,N_8127,N_8792);
and U9975 (N_9975,N_8704,N_8116);
or U9976 (N_9976,N_8368,N_8872);
nor U9977 (N_9977,N_8212,N_8189);
xnor U9978 (N_9978,N_8608,N_8680);
nand U9979 (N_9979,N_8048,N_8215);
xnor U9980 (N_9980,N_8494,N_8876);
nand U9981 (N_9981,N_8235,N_8478);
nand U9982 (N_9982,N_8466,N_8056);
or U9983 (N_9983,N_8921,N_8326);
nor U9984 (N_9984,N_8770,N_8781);
and U9985 (N_9985,N_8087,N_8054);
nand U9986 (N_9986,N_8801,N_8456);
xor U9987 (N_9987,N_8831,N_8191);
xor U9988 (N_9988,N_8652,N_8698);
and U9989 (N_9989,N_8997,N_8345);
xor U9990 (N_9990,N_8539,N_8638);
xnor U9991 (N_9991,N_8441,N_8396);
nor U9992 (N_9992,N_8051,N_8668);
and U9993 (N_9993,N_8582,N_8143);
xor U9994 (N_9994,N_8132,N_8716);
xnor U9995 (N_9995,N_8738,N_8697);
nand U9996 (N_9996,N_8162,N_8719);
or U9997 (N_9997,N_8245,N_8074);
nand U9998 (N_9998,N_8145,N_8331);
nand U9999 (N_9999,N_8683,N_8295);
or UO_0 (O_0,N_9849,N_9783);
nand UO_1 (O_1,N_9716,N_9722);
nor UO_2 (O_2,N_9992,N_9087);
and UO_3 (O_3,N_9214,N_9706);
nand UO_4 (O_4,N_9526,N_9175);
nand UO_5 (O_5,N_9945,N_9182);
nand UO_6 (O_6,N_9598,N_9870);
xor UO_7 (O_7,N_9868,N_9865);
nor UO_8 (O_8,N_9724,N_9405);
nand UO_9 (O_9,N_9862,N_9807);
xor UO_10 (O_10,N_9470,N_9277);
xnor UO_11 (O_11,N_9692,N_9154);
or UO_12 (O_12,N_9573,N_9272);
and UO_13 (O_13,N_9645,N_9800);
or UO_14 (O_14,N_9840,N_9274);
nor UO_15 (O_15,N_9981,N_9636);
nor UO_16 (O_16,N_9602,N_9519);
and UO_17 (O_17,N_9371,N_9581);
nor UO_18 (O_18,N_9540,N_9151);
nor UO_19 (O_19,N_9492,N_9975);
nand UO_20 (O_20,N_9253,N_9976);
xor UO_21 (O_21,N_9687,N_9444);
and UO_22 (O_22,N_9583,N_9196);
xor UO_23 (O_23,N_9349,N_9249);
nor UO_24 (O_24,N_9968,N_9856);
or UO_25 (O_25,N_9306,N_9203);
nand UO_26 (O_26,N_9259,N_9717);
nand UO_27 (O_27,N_9209,N_9138);
and UO_28 (O_28,N_9147,N_9913);
nor UO_29 (O_29,N_9971,N_9891);
nand UO_30 (O_30,N_9069,N_9045);
nand UO_31 (O_31,N_9662,N_9163);
nor UO_32 (O_32,N_9502,N_9829);
or UO_33 (O_33,N_9806,N_9431);
and UO_34 (O_34,N_9586,N_9746);
and UO_35 (O_35,N_9097,N_9893);
or UO_36 (O_36,N_9300,N_9179);
or UO_37 (O_37,N_9130,N_9033);
nor UO_38 (O_38,N_9284,N_9419);
nand UO_39 (O_39,N_9879,N_9651);
or UO_40 (O_40,N_9319,N_9226);
xor UO_41 (O_41,N_9423,N_9907);
xnor UO_42 (O_42,N_9858,N_9961);
xor UO_43 (O_43,N_9863,N_9733);
and UO_44 (O_44,N_9506,N_9612);
nand UO_45 (O_45,N_9798,N_9458);
or UO_46 (O_46,N_9321,N_9430);
xnor UO_47 (O_47,N_9940,N_9322);
nor UO_48 (O_48,N_9665,N_9972);
and UO_49 (O_49,N_9185,N_9936);
nor UO_50 (O_50,N_9989,N_9591);
and UO_51 (O_51,N_9691,N_9142);
nand UO_52 (O_52,N_9737,N_9122);
nor UO_53 (O_53,N_9754,N_9592);
and UO_54 (O_54,N_9299,N_9571);
nand UO_55 (O_55,N_9565,N_9049);
nor UO_56 (O_56,N_9118,N_9367);
or UO_57 (O_57,N_9167,N_9370);
nor UO_58 (O_58,N_9345,N_9790);
nor UO_59 (O_59,N_9486,N_9448);
nor UO_60 (O_60,N_9312,N_9273);
xor UO_61 (O_61,N_9315,N_9133);
nand UO_62 (O_62,N_9894,N_9080);
xnor UO_63 (O_63,N_9174,N_9043);
xnor UO_64 (O_64,N_9984,N_9738);
or UO_65 (O_65,N_9445,N_9568);
xor UO_66 (O_66,N_9081,N_9011);
or UO_67 (O_67,N_9648,N_9135);
xor UO_68 (O_68,N_9326,N_9019);
and UO_69 (O_69,N_9335,N_9892);
nand UO_70 (O_70,N_9657,N_9755);
nand UO_71 (O_71,N_9762,N_9295);
nand UO_72 (O_72,N_9451,N_9973);
and UO_73 (O_73,N_9217,N_9885);
xnor UO_74 (O_74,N_9361,N_9333);
nand UO_75 (O_75,N_9603,N_9702);
or UO_76 (O_76,N_9521,N_9801);
and UO_77 (O_77,N_9044,N_9403);
nand UO_78 (O_78,N_9358,N_9567);
nand UO_79 (O_79,N_9629,N_9942);
and UO_80 (O_80,N_9157,N_9394);
nand UO_81 (O_81,N_9908,N_9670);
nand UO_82 (O_82,N_9917,N_9642);
or UO_83 (O_83,N_9794,N_9524);
and UO_84 (O_84,N_9171,N_9079);
xor UO_85 (O_85,N_9343,N_9522);
xor UO_86 (O_86,N_9161,N_9041);
nand UO_87 (O_87,N_9770,N_9632);
xnor UO_88 (O_88,N_9412,N_9239);
xor UO_89 (O_89,N_9169,N_9088);
nand UO_90 (O_90,N_9761,N_9778);
or UO_91 (O_91,N_9339,N_9823);
nand UO_92 (O_92,N_9034,N_9546);
xnor UO_93 (O_93,N_9720,N_9488);
and UO_94 (O_94,N_9771,N_9726);
xor UO_95 (O_95,N_9970,N_9535);
or UO_96 (O_96,N_9094,N_9215);
nor UO_97 (O_97,N_9268,N_9532);
or UO_98 (O_98,N_9186,N_9229);
nand UO_99 (O_99,N_9036,N_9509);
nand UO_100 (O_100,N_9523,N_9918);
nor UO_101 (O_101,N_9897,N_9276);
or UO_102 (O_102,N_9883,N_9510);
nor UO_103 (O_103,N_9597,N_9287);
and UO_104 (O_104,N_9281,N_9734);
xnor UO_105 (O_105,N_9621,N_9388);
xor UO_106 (O_106,N_9495,N_9416);
xnor UO_107 (O_107,N_9980,N_9463);
nand UO_108 (O_108,N_9758,N_9000);
and UO_109 (O_109,N_9666,N_9729);
or UO_110 (O_110,N_9134,N_9541);
nor UO_111 (O_111,N_9813,N_9466);
and UO_112 (O_112,N_9475,N_9835);
or UO_113 (O_113,N_9245,N_9504);
xnor UO_114 (O_114,N_9380,N_9310);
nand UO_115 (O_115,N_9139,N_9655);
or UO_116 (O_116,N_9987,N_9127);
nor UO_117 (O_117,N_9562,N_9904);
nor UO_118 (O_118,N_9355,N_9404);
or UO_119 (O_119,N_9108,N_9331);
nor UO_120 (O_120,N_9450,N_9173);
xnor UO_121 (O_121,N_9517,N_9165);
xor UO_122 (O_122,N_9847,N_9810);
and UO_123 (O_123,N_9503,N_9301);
and UO_124 (O_124,N_9549,N_9967);
xor UO_125 (O_125,N_9838,N_9786);
and UO_126 (O_126,N_9145,N_9525);
nand UO_127 (O_127,N_9620,N_9210);
nor UO_128 (O_128,N_9781,N_9252);
and UO_129 (O_129,N_9415,N_9377);
and UO_130 (O_130,N_9076,N_9035);
xor UO_131 (O_131,N_9283,N_9410);
nor UO_132 (O_132,N_9815,N_9650);
nand UO_133 (O_133,N_9688,N_9797);
or UO_134 (O_134,N_9407,N_9836);
xor UO_135 (O_135,N_9789,N_9796);
and UO_136 (O_136,N_9227,N_9727);
or UO_137 (O_137,N_9582,N_9105);
nand UO_138 (O_138,N_9348,N_9384);
and UO_139 (O_139,N_9042,N_9825);
nand UO_140 (O_140,N_9282,N_9158);
xor UO_141 (O_141,N_9180,N_9378);
xor UO_142 (O_142,N_9822,N_9063);
or UO_143 (O_143,N_9741,N_9457);
and UO_144 (O_144,N_9544,N_9735);
or UO_145 (O_145,N_9515,N_9008);
and UO_146 (O_146,N_9334,N_9327);
and UO_147 (O_147,N_9123,N_9811);
and UO_148 (O_148,N_9429,N_9514);
xor UO_149 (O_149,N_9831,N_9694);
nand UO_150 (O_150,N_9050,N_9777);
xnor UO_151 (O_151,N_9162,N_9854);
nand UO_152 (O_152,N_9278,N_9604);
or UO_153 (O_153,N_9837,N_9479);
nand UO_154 (O_154,N_9064,N_9784);
and UO_155 (O_155,N_9191,N_9255);
nor UO_156 (O_156,N_9022,N_9647);
nand UO_157 (O_157,N_9843,N_9844);
xnor UO_158 (O_158,N_9120,N_9630);
nor UO_159 (O_159,N_9183,N_9285);
nand UO_160 (O_160,N_9817,N_9750);
or UO_161 (O_161,N_9136,N_9164);
xnor UO_162 (O_162,N_9440,N_9491);
nor UO_163 (O_163,N_9328,N_9946);
and UO_164 (O_164,N_9654,N_9235);
or UO_165 (O_165,N_9812,N_9958);
nor UO_166 (O_166,N_9442,N_9697);
and UO_167 (O_167,N_9425,N_9474);
xnor UO_168 (O_168,N_9015,N_9767);
nor UO_169 (O_169,N_9615,N_9112);
nor UO_170 (O_170,N_9082,N_9114);
and UO_171 (O_171,N_9518,N_9258);
xor UO_172 (O_172,N_9159,N_9718);
or UO_173 (O_173,N_9251,N_9799);
or UO_174 (O_174,N_9176,N_9600);
and UO_175 (O_175,N_9024,N_9928);
xnor UO_176 (O_176,N_9710,N_9387);
nor UO_177 (O_177,N_9920,N_9323);
and UO_178 (O_178,N_9626,N_9129);
or UO_179 (O_179,N_9834,N_9414);
nor UO_180 (O_180,N_9742,N_9955);
xor UO_181 (O_181,N_9529,N_9288);
nand UO_182 (O_182,N_9137,N_9638);
xor UO_183 (O_183,N_9668,N_9207);
nor UO_184 (O_184,N_9456,N_9680);
nand UO_185 (O_185,N_9641,N_9508);
and UO_186 (O_186,N_9902,N_9611);
nor UO_187 (O_187,N_9420,N_9505);
nand UO_188 (O_188,N_9585,N_9411);
nand UO_189 (O_189,N_9839,N_9601);
xor UO_190 (O_190,N_9385,N_9313);
nand UO_191 (O_191,N_9267,N_9808);
and UO_192 (O_192,N_9693,N_9464);
or UO_193 (O_193,N_9939,N_9704);
nor UO_194 (O_194,N_9511,N_9441);
and UO_195 (O_195,N_9351,N_9764);
and UO_196 (O_196,N_9469,N_9098);
nand UO_197 (O_197,N_9350,N_9153);
xnor UO_198 (O_198,N_9991,N_9888);
xnor UO_199 (O_199,N_9760,N_9496);
or UO_200 (O_200,N_9279,N_9853);
nor UO_201 (O_201,N_9805,N_9923);
or UO_202 (O_202,N_9951,N_9698);
xor UO_203 (O_203,N_9408,N_9884);
nor UO_204 (O_204,N_9721,N_9305);
and UO_205 (O_205,N_9452,N_9564);
nand UO_206 (O_206,N_9205,N_9520);
or UO_207 (O_207,N_9494,N_9449);
and UO_208 (O_208,N_9117,N_9131);
xnor UO_209 (O_209,N_9409,N_9964);
nand UO_210 (O_210,N_9471,N_9516);
xor UO_211 (O_211,N_9999,N_9934);
nor UO_212 (O_212,N_9330,N_9435);
nand UO_213 (O_213,N_9017,N_9290);
nand UO_214 (O_214,N_9625,N_9937);
nor UO_215 (O_215,N_9149,N_9553);
nand UO_216 (O_216,N_9990,N_9914);
and UO_217 (O_217,N_9714,N_9200);
or UO_218 (O_218,N_9792,N_9874);
xnor UO_219 (O_219,N_9880,N_9211);
or UO_220 (O_220,N_9743,N_9985);
and UO_221 (O_221,N_9896,N_9166);
nor UO_222 (O_222,N_9685,N_9609);
or UO_223 (O_223,N_9085,N_9426);
nor UO_224 (O_224,N_9700,N_9490);
xor UO_225 (O_225,N_9803,N_9690);
nand UO_226 (O_226,N_9298,N_9346);
nor UO_227 (O_227,N_9187,N_9606);
and UO_228 (O_228,N_9393,N_9121);
nor UO_229 (O_229,N_9631,N_9998);
xnor UO_230 (O_230,N_9639,N_9595);
nand UO_231 (O_231,N_9070,N_9878);
and UO_232 (O_232,N_9219,N_9696);
or UO_233 (O_233,N_9857,N_9374);
nand UO_234 (O_234,N_9563,N_9238);
nand UO_235 (O_235,N_9360,N_9247);
nor UO_236 (O_236,N_9204,N_9029);
or UO_237 (O_237,N_9325,N_9689);
or UO_238 (O_238,N_9617,N_9749);
or UO_239 (O_239,N_9341,N_9240);
nand UO_240 (O_240,N_9102,N_9782);
and UO_241 (O_241,N_9744,N_9013);
nor UO_242 (O_242,N_9634,N_9652);
nand UO_243 (O_243,N_9280,N_9254);
or UO_244 (O_244,N_9307,N_9538);
and UO_245 (O_245,N_9552,N_9125);
nor UO_246 (O_246,N_9763,N_9931);
nor UO_247 (O_247,N_9977,N_9925);
and UO_248 (O_248,N_9086,N_9643);
and UO_249 (O_249,N_9318,N_9181);
or UO_250 (O_250,N_9730,N_9140);
nor UO_251 (O_251,N_9910,N_9177);
nand UO_252 (O_252,N_9059,N_9401);
and UO_253 (O_253,N_9788,N_9673);
or UO_254 (O_254,N_9453,N_9842);
nor UO_255 (O_255,N_9398,N_9266);
or UO_256 (O_256,N_9357,N_9188);
or UO_257 (O_257,N_9060,N_9198);
or UO_258 (O_258,N_9093,N_9500);
nor UO_259 (O_259,N_9876,N_9739);
and UO_260 (O_260,N_9293,N_9962);
or UO_261 (O_261,N_9294,N_9633);
xor UO_262 (O_262,N_9004,N_9663);
and UO_263 (O_263,N_9055,N_9170);
and UO_264 (O_264,N_9827,N_9462);
or UO_265 (O_265,N_9804,N_9575);
or UO_266 (O_266,N_9988,N_9912);
or UO_267 (O_267,N_9978,N_9869);
nor UO_268 (O_268,N_9155,N_9588);
xnor UO_269 (O_269,N_9993,N_9664);
xor UO_270 (O_270,N_9428,N_9954);
nand UO_271 (O_271,N_9189,N_9433);
nor UO_272 (O_272,N_9368,N_9481);
and UO_273 (O_273,N_9028,N_9947);
nor UO_274 (O_274,N_9202,N_9460);
nor UO_275 (O_275,N_9895,N_9719);
xnor UO_276 (O_276,N_9422,N_9264);
nor UO_277 (O_277,N_9144,N_9677);
nand UO_278 (O_278,N_9038,N_9675);
or UO_279 (O_279,N_9037,N_9314);
and UO_280 (O_280,N_9396,N_9455);
or UO_281 (O_281,N_9787,N_9051);
nor UO_282 (O_282,N_9774,N_9286);
or UO_283 (O_283,N_9875,N_9821);
and UO_284 (O_284,N_9221,N_9545);
nand UO_285 (O_285,N_9132,N_9311);
nand UO_286 (O_286,N_9480,N_9833);
and UO_287 (O_287,N_9556,N_9201);
nor UO_288 (O_288,N_9048,N_9966);
or UO_289 (O_289,N_9695,N_9848);
xor UO_290 (O_290,N_9599,N_9053);
or UO_291 (O_291,N_9026,N_9745);
nand UO_292 (O_292,N_9194,N_9485);
and UO_293 (O_293,N_9859,N_9501);
nor UO_294 (O_294,N_9828,N_9772);
and UO_295 (O_295,N_9941,N_9230);
nor UO_296 (O_296,N_9418,N_9402);
or UO_297 (O_297,N_9699,N_9372);
nand UO_298 (O_298,N_9536,N_9578);
and UO_299 (O_299,N_9587,N_9785);
or UO_300 (O_300,N_9152,N_9974);
nor UO_301 (O_301,N_9773,N_9555);
and UO_302 (O_302,N_9397,N_9512);
xor UO_303 (O_303,N_9881,N_9559);
nor UO_304 (O_304,N_9107,N_9911);
and UO_305 (O_305,N_9197,N_9062);
and UO_306 (O_306,N_9099,N_9671);
xnor UO_307 (O_307,N_9391,N_9381);
xnor UO_308 (O_308,N_9250,N_9542);
xor UO_309 (O_309,N_9047,N_9101);
and UO_310 (O_310,N_9484,N_9814);
nor UO_311 (O_311,N_9459,N_9231);
nand UO_312 (O_312,N_9950,N_9338);
or UO_313 (O_313,N_9454,N_9543);
and UO_314 (O_314,N_9949,N_9483);
or UO_315 (O_315,N_9432,N_9222);
and UO_316 (O_316,N_9030,N_9924);
nor UO_317 (O_317,N_9447,N_9190);
or UO_318 (O_318,N_9579,N_9329);
and UO_319 (O_319,N_9382,N_9216);
or UO_320 (O_320,N_9659,N_9065);
xor UO_321 (O_321,N_9528,N_9653);
and UO_322 (O_322,N_9906,N_9903);
nor UO_323 (O_323,N_9872,N_9148);
nand UO_324 (O_324,N_9237,N_9003);
nand UO_325 (O_325,N_9243,N_9933);
nand UO_326 (O_326,N_9871,N_9195);
nor UO_327 (O_327,N_9212,N_9270);
nor UO_328 (O_328,N_9084,N_9332);
or UO_329 (O_329,N_9260,N_9867);
nand UO_330 (O_330,N_9531,N_9427);
or UO_331 (O_331,N_9905,N_9354);
nor UO_332 (O_332,N_9852,N_9846);
nor UO_333 (O_333,N_9106,N_9110);
xor UO_334 (O_334,N_9793,N_9759);
or UO_335 (O_335,N_9709,N_9395);
nand UO_336 (O_336,N_9364,N_9256);
xnor UO_337 (O_337,N_9953,N_9607);
nand UO_338 (O_338,N_9056,N_9009);
nor UO_339 (O_339,N_9539,N_9344);
and UO_340 (O_340,N_9554,N_9969);
nor UO_341 (O_341,N_9461,N_9703);
xnor UO_342 (O_342,N_9986,N_9927);
nand UO_343 (O_343,N_9683,N_9873);
nor UO_344 (O_344,N_9021,N_9006);
nor UO_345 (O_345,N_9126,N_9039);
xnor UO_346 (O_346,N_9077,N_9146);
nor UO_347 (O_347,N_9537,N_9948);
nor UO_348 (O_348,N_9096,N_9882);
nor UO_349 (O_349,N_9078,N_9635);
nor UO_350 (O_350,N_9909,N_9889);
nor UO_351 (O_351,N_9845,N_9246);
nor UO_352 (O_352,N_9551,N_9413);
xnor UO_353 (O_353,N_9242,N_9072);
and UO_354 (O_354,N_9437,N_9656);
and UO_355 (O_355,N_9596,N_9627);
and UO_356 (O_356,N_9446,N_9681);
or UO_357 (O_357,N_9373,N_9667);
nand UO_358 (O_358,N_9574,N_9618);
or UO_359 (O_359,N_9715,N_9390);
and UO_360 (O_360,N_9399,N_9468);
or UO_361 (O_361,N_9213,N_9058);
xor UO_362 (O_362,N_9262,N_9225);
nor UO_363 (O_363,N_9802,N_9557);
xnor UO_364 (O_364,N_9850,N_9115);
xor UO_365 (O_365,N_9297,N_9296);
or UO_366 (O_366,N_9956,N_9018);
nand UO_367 (O_367,N_9866,N_9548);
or UO_368 (O_368,N_9851,N_9233);
and UO_369 (O_369,N_9637,N_9753);
nor UO_370 (O_370,N_9886,N_9747);
xor UO_371 (O_371,N_9304,N_9765);
nor UO_372 (O_372,N_9830,N_9944);
nor UO_373 (O_373,N_9560,N_9593);
or UO_374 (O_374,N_9952,N_9473);
nand UO_375 (O_375,N_9111,N_9795);
or UO_376 (O_376,N_9031,N_9590);
xnor UO_377 (O_377,N_9308,N_9569);
and UO_378 (O_378,N_9032,N_9589);
xnor UO_379 (O_379,N_9686,N_9701);
nand UO_380 (O_380,N_9025,N_9089);
and UO_381 (O_381,N_9365,N_9608);
xnor UO_382 (O_382,N_9061,N_9605);
xnor UO_383 (O_383,N_9960,N_9644);
or UO_384 (O_384,N_9369,N_9919);
and UO_385 (O_385,N_9887,N_9820);
nor UO_386 (O_386,N_9580,N_9083);
nor UO_387 (O_387,N_9982,N_9658);
or UO_388 (O_388,N_9731,N_9340);
nand UO_389 (O_389,N_9320,N_9040);
xor UO_390 (O_390,N_9406,N_9100);
and UO_391 (O_391,N_9669,N_9769);
nor UO_392 (O_392,N_9930,N_9316);
and UO_393 (O_393,N_9576,N_9566);
xor UO_394 (O_394,N_9116,N_9624);
nand UO_395 (O_395,N_9071,N_9317);
or UO_396 (O_396,N_9092,N_9926);
xor UO_397 (O_397,N_9275,N_9487);
xnor UO_398 (O_398,N_9932,N_9497);
nand UO_399 (O_399,N_9236,N_9660);
or UO_400 (O_400,N_9899,N_9725);
and UO_401 (O_401,N_9594,N_9527);
nand UO_402 (O_402,N_9066,N_9128);
nand UO_403 (O_403,N_9534,N_9016);
or UO_404 (O_404,N_9223,N_9674);
xor UO_405 (O_405,N_9438,N_9218);
nand UO_406 (O_406,N_9757,N_9054);
nand UO_407 (O_407,N_9756,N_9199);
or UO_408 (O_408,N_9832,N_9498);
nand UO_409 (O_409,N_9610,N_9291);
nor UO_410 (O_410,N_9324,N_9499);
xnor UO_411 (O_411,N_9192,N_9465);
nor UO_412 (O_412,N_9855,N_9678);
or UO_413 (O_413,N_9994,N_9376);
nand UO_414 (O_414,N_9752,N_9616);
and UO_415 (O_415,N_9943,N_9386);
and UO_416 (O_416,N_9068,N_9682);
nor UO_417 (O_417,N_9248,N_9723);
or UO_418 (O_418,N_9861,N_9614);
nor UO_419 (O_419,N_9156,N_9400);
xor UO_420 (O_420,N_9265,N_9020);
or UO_421 (O_421,N_9417,N_9558);
xnor UO_422 (O_422,N_9818,N_9113);
nor UO_423 (O_423,N_9957,N_9860);
and UO_424 (O_424,N_9023,N_9091);
and UO_425 (O_425,N_9561,N_9513);
xor UO_426 (O_426,N_9732,N_9220);
and UO_427 (O_427,N_9168,N_9119);
nand UO_428 (O_428,N_9383,N_9005);
nor UO_429 (O_429,N_9103,N_9915);
nand UO_430 (O_430,N_9073,N_9389);
nand UO_431 (O_431,N_9302,N_9363);
or UO_432 (O_432,N_9996,N_9359);
xnor UO_433 (O_433,N_9779,N_9672);
and UO_434 (O_434,N_9679,N_9232);
and UO_435 (O_435,N_9261,N_9347);
nor UO_436 (O_436,N_9224,N_9929);
or UO_437 (O_437,N_9392,N_9622);
and UO_438 (O_438,N_9027,N_9748);
nor UO_439 (O_439,N_9012,N_9547);
and UO_440 (O_440,N_9963,N_9095);
nand UO_441 (O_441,N_9057,N_9661);
nor UO_442 (O_442,N_9467,N_9751);
nand UO_443 (O_443,N_9356,N_9676);
nor UO_444 (O_444,N_9472,N_9424);
nand UO_445 (O_445,N_9826,N_9309);
xnor UO_446 (O_446,N_9476,N_9206);
and UO_447 (O_447,N_9109,N_9995);
and UO_448 (O_448,N_9143,N_9421);
and UO_449 (O_449,N_9292,N_9877);
nor UO_450 (O_450,N_9184,N_9916);
nand UO_451 (O_451,N_9160,N_9841);
or UO_452 (O_452,N_9478,N_9768);
or UO_453 (O_453,N_9443,N_9684);
and UO_454 (O_454,N_9482,N_9208);
nor UO_455 (O_455,N_9271,N_9628);
nand UO_456 (O_456,N_9646,N_9353);
nand UO_457 (O_457,N_9619,N_9375);
nor UO_458 (O_458,N_9533,N_9766);
xor UO_459 (O_459,N_9439,N_9921);
nor UO_460 (O_460,N_9938,N_9257);
and UO_461 (O_461,N_9613,N_9809);
and UO_462 (O_462,N_9935,N_9014);
xor UO_463 (O_463,N_9705,N_9983);
nand UO_464 (O_464,N_9640,N_9052);
and UO_465 (O_465,N_9959,N_9776);
and UO_466 (O_466,N_9074,N_9922);
or UO_467 (O_467,N_9362,N_9001);
nor UO_468 (O_468,N_9178,N_9493);
nand UO_469 (O_469,N_9342,N_9577);
nor UO_470 (O_470,N_9172,N_9901);
or UO_471 (O_471,N_9104,N_9900);
nor UO_472 (O_472,N_9075,N_9819);
or UO_473 (O_473,N_9864,N_9713);
or UO_474 (O_474,N_9366,N_9244);
xor UO_475 (O_475,N_9150,N_9007);
nor UO_476 (O_476,N_9241,N_9816);
and UO_477 (O_477,N_9728,N_9572);
xnor UO_478 (O_478,N_9067,N_9269);
xor UO_479 (O_479,N_9337,N_9289);
and UO_480 (O_480,N_9550,N_9090);
nand UO_481 (O_481,N_9898,N_9507);
and UO_482 (O_482,N_9434,N_9228);
xnor UO_483 (O_483,N_9708,N_9623);
xor UO_484 (O_484,N_9436,N_9824);
nor UO_485 (O_485,N_9736,N_9570);
nand UO_486 (O_486,N_9775,N_9780);
and UO_487 (O_487,N_9303,N_9979);
nand UO_488 (O_488,N_9336,N_9711);
and UO_489 (O_489,N_9234,N_9352);
nor UO_490 (O_490,N_9707,N_9584);
or UO_491 (O_491,N_9712,N_9740);
or UO_492 (O_492,N_9791,N_9379);
nor UO_493 (O_493,N_9649,N_9530);
nor UO_494 (O_494,N_9489,N_9046);
and UO_495 (O_495,N_9263,N_9124);
nand UO_496 (O_496,N_9965,N_9890);
or UO_497 (O_497,N_9141,N_9002);
nand UO_498 (O_498,N_9010,N_9193);
nor UO_499 (O_499,N_9477,N_9997);
or UO_500 (O_500,N_9143,N_9015);
nor UO_501 (O_501,N_9333,N_9503);
xor UO_502 (O_502,N_9635,N_9383);
nor UO_503 (O_503,N_9513,N_9880);
or UO_504 (O_504,N_9672,N_9620);
or UO_505 (O_505,N_9987,N_9650);
nand UO_506 (O_506,N_9695,N_9046);
and UO_507 (O_507,N_9954,N_9226);
xor UO_508 (O_508,N_9618,N_9171);
or UO_509 (O_509,N_9690,N_9601);
nor UO_510 (O_510,N_9866,N_9636);
and UO_511 (O_511,N_9221,N_9071);
nand UO_512 (O_512,N_9647,N_9956);
xnor UO_513 (O_513,N_9860,N_9759);
nand UO_514 (O_514,N_9451,N_9545);
nor UO_515 (O_515,N_9450,N_9051);
or UO_516 (O_516,N_9361,N_9138);
or UO_517 (O_517,N_9360,N_9219);
and UO_518 (O_518,N_9052,N_9476);
and UO_519 (O_519,N_9888,N_9629);
nor UO_520 (O_520,N_9011,N_9146);
nand UO_521 (O_521,N_9993,N_9630);
or UO_522 (O_522,N_9180,N_9753);
and UO_523 (O_523,N_9628,N_9930);
nor UO_524 (O_524,N_9752,N_9316);
xor UO_525 (O_525,N_9827,N_9318);
nand UO_526 (O_526,N_9804,N_9234);
xor UO_527 (O_527,N_9844,N_9825);
or UO_528 (O_528,N_9988,N_9762);
or UO_529 (O_529,N_9389,N_9687);
and UO_530 (O_530,N_9486,N_9085);
or UO_531 (O_531,N_9933,N_9477);
or UO_532 (O_532,N_9846,N_9060);
and UO_533 (O_533,N_9813,N_9371);
and UO_534 (O_534,N_9451,N_9898);
nor UO_535 (O_535,N_9539,N_9541);
nand UO_536 (O_536,N_9146,N_9259);
nor UO_537 (O_537,N_9394,N_9462);
nor UO_538 (O_538,N_9904,N_9419);
and UO_539 (O_539,N_9469,N_9199);
xnor UO_540 (O_540,N_9754,N_9034);
and UO_541 (O_541,N_9192,N_9418);
xor UO_542 (O_542,N_9731,N_9398);
xor UO_543 (O_543,N_9270,N_9995);
nand UO_544 (O_544,N_9094,N_9291);
xor UO_545 (O_545,N_9320,N_9776);
nand UO_546 (O_546,N_9832,N_9932);
nor UO_547 (O_547,N_9964,N_9798);
nand UO_548 (O_548,N_9975,N_9287);
nand UO_549 (O_549,N_9406,N_9952);
and UO_550 (O_550,N_9606,N_9509);
nand UO_551 (O_551,N_9246,N_9175);
nor UO_552 (O_552,N_9726,N_9257);
and UO_553 (O_553,N_9419,N_9639);
nand UO_554 (O_554,N_9710,N_9276);
nand UO_555 (O_555,N_9937,N_9204);
xor UO_556 (O_556,N_9697,N_9581);
xnor UO_557 (O_557,N_9955,N_9183);
and UO_558 (O_558,N_9030,N_9726);
or UO_559 (O_559,N_9944,N_9104);
nor UO_560 (O_560,N_9861,N_9911);
xnor UO_561 (O_561,N_9911,N_9994);
nor UO_562 (O_562,N_9724,N_9823);
nor UO_563 (O_563,N_9413,N_9052);
xnor UO_564 (O_564,N_9436,N_9384);
xnor UO_565 (O_565,N_9276,N_9443);
or UO_566 (O_566,N_9524,N_9493);
xnor UO_567 (O_567,N_9314,N_9271);
nand UO_568 (O_568,N_9237,N_9743);
nand UO_569 (O_569,N_9471,N_9946);
xnor UO_570 (O_570,N_9920,N_9225);
nand UO_571 (O_571,N_9122,N_9896);
nand UO_572 (O_572,N_9816,N_9732);
nand UO_573 (O_573,N_9147,N_9253);
or UO_574 (O_574,N_9948,N_9080);
xor UO_575 (O_575,N_9149,N_9509);
nor UO_576 (O_576,N_9133,N_9794);
or UO_577 (O_577,N_9960,N_9698);
or UO_578 (O_578,N_9212,N_9731);
nor UO_579 (O_579,N_9690,N_9448);
or UO_580 (O_580,N_9184,N_9018);
xnor UO_581 (O_581,N_9176,N_9142);
nor UO_582 (O_582,N_9873,N_9348);
and UO_583 (O_583,N_9623,N_9751);
or UO_584 (O_584,N_9774,N_9799);
xor UO_585 (O_585,N_9365,N_9197);
nand UO_586 (O_586,N_9357,N_9049);
or UO_587 (O_587,N_9248,N_9265);
or UO_588 (O_588,N_9621,N_9159);
nor UO_589 (O_589,N_9077,N_9450);
and UO_590 (O_590,N_9599,N_9381);
xnor UO_591 (O_591,N_9025,N_9705);
and UO_592 (O_592,N_9058,N_9982);
and UO_593 (O_593,N_9000,N_9776);
and UO_594 (O_594,N_9994,N_9948);
and UO_595 (O_595,N_9644,N_9906);
or UO_596 (O_596,N_9892,N_9020);
and UO_597 (O_597,N_9055,N_9217);
or UO_598 (O_598,N_9450,N_9868);
nor UO_599 (O_599,N_9445,N_9065);
or UO_600 (O_600,N_9491,N_9893);
and UO_601 (O_601,N_9112,N_9553);
nand UO_602 (O_602,N_9831,N_9335);
nand UO_603 (O_603,N_9848,N_9494);
nand UO_604 (O_604,N_9515,N_9172);
or UO_605 (O_605,N_9959,N_9435);
xor UO_606 (O_606,N_9067,N_9790);
xnor UO_607 (O_607,N_9739,N_9560);
nor UO_608 (O_608,N_9323,N_9444);
nand UO_609 (O_609,N_9190,N_9443);
and UO_610 (O_610,N_9884,N_9882);
xnor UO_611 (O_611,N_9025,N_9277);
or UO_612 (O_612,N_9523,N_9522);
or UO_613 (O_613,N_9503,N_9084);
nor UO_614 (O_614,N_9748,N_9755);
nand UO_615 (O_615,N_9796,N_9644);
xor UO_616 (O_616,N_9009,N_9496);
nor UO_617 (O_617,N_9043,N_9200);
and UO_618 (O_618,N_9613,N_9705);
and UO_619 (O_619,N_9748,N_9263);
nor UO_620 (O_620,N_9609,N_9538);
xor UO_621 (O_621,N_9640,N_9400);
xnor UO_622 (O_622,N_9793,N_9384);
or UO_623 (O_623,N_9190,N_9897);
xnor UO_624 (O_624,N_9792,N_9609);
nor UO_625 (O_625,N_9128,N_9528);
nand UO_626 (O_626,N_9152,N_9165);
or UO_627 (O_627,N_9839,N_9866);
or UO_628 (O_628,N_9039,N_9071);
xnor UO_629 (O_629,N_9046,N_9297);
and UO_630 (O_630,N_9375,N_9095);
nor UO_631 (O_631,N_9303,N_9791);
nor UO_632 (O_632,N_9396,N_9410);
nor UO_633 (O_633,N_9366,N_9278);
and UO_634 (O_634,N_9178,N_9192);
nor UO_635 (O_635,N_9492,N_9551);
xnor UO_636 (O_636,N_9284,N_9763);
and UO_637 (O_637,N_9616,N_9596);
nand UO_638 (O_638,N_9590,N_9594);
xnor UO_639 (O_639,N_9746,N_9338);
xor UO_640 (O_640,N_9646,N_9432);
xnor UO_641 (O_641,N_9611,N_9378);
nand UO_642 (O_642,N_9985,N_9569);
and UO_643 (O_643,N_9655,N_9405);
and UO_644 (O_644,N_9606,N_9625);
or UO_645 (O_645,N_9181,N_9107);
xor UO_646 (O_646,N_9738,N_9915);
or UO_647 (O_647,N_9681,N_9055);
and UO_648 (O_648,N_9359,N_9121);
nor UO_649 (O_649,N_9515,N_9560);
nand UO_650 (O_650,N_9220,N_9560);
xnor UO_651 (O_651,N_9973,N_9487);
xnor UO_652 (O_652,N_9245,N_9532);
xnor UO_653 (O_653,N_9604,N_9823);
xor UO_654 (O_654,N_9774,N_9884);
nand UO_655 (O_655,N_9142,N_9805);
or UO_656 (O_656,N_9879,N_9687);
nand UO_657 (O_657,N_9623,N_9922);
and UO_658 (O_658,N_9809,N_9322);
nand UO_659 (O_659,N_9243,N_9173);
and UO_660 (O_660,N_9743,N_9991);
or UO_661 (O_661,N_9910,N_9144);
and UO_662 (O_662,N_9402,N_9007);
or UO_663 (O_663,N_9910,N_9392);
xnor UO_664 (O_664,N_9756,N_9649);
or UO_665 (O_665,N_9868,N_9284);
xnor UO_666 (O_666,N_9044,N_9878);
and UO_667 (O_667,N_9734,N_9448);
or UO_668 (O_668,N_9664,N_9178);
and UO_669 (O_669,N_9949,N_9814);
and UO_670 (O_670,N_9291,N_9423);
xnor UO_671 (O_671,N_9446,N_9462);
nor UO_672 (O_672,N_9285,N_9727);
nor UO_673 (O_673,N_9373,N_9895);
nor UO_674 (O_674,N_9766,N_9993);
or UO_675 (O_675,N_9109,N_9564);
nand UO_676 (O_676,N_9137,N_9640);
and UO_677 (O_677,N_9052,N_9535);
or UO_678 (O_678,N_9129,N_9679);
xor UO_679 (O_679,N_9815,N_9465);
nand UO_680 (O_680,N_9586,N_9082);
nor UO_681 (O_681,N_9809,N_9279);
nand UO_682 (O_682,N_9709,N_9050);
nand UO_683 (O_683,N_9492,N_9547);
xnor UO_684 (O_684,N_9657,N_9766);
or UO_685 (O_685,N_9817,N_9866);
xor UO_686 (O_686,N_9596,N_9756);
and UO_687 (O_687,N_9077,N_9362);
nand UO_688 (O_688,N_9597,N_9443);
and UO_689 (O_689,N_9045,N_9272);
nand UO_690 (O_690,N_9838,N_9263);
nand UO_691 (O_691,N_9409,N_9701);
or UO_692 (O_692,N_9860,N_9677);
xnor UO_693 (O_693,N_9842,N_9930);
or UO_694 (O_694,N_9308,N_9393);
and UO_695 (O_695,N_9287,N_9652);
nor UO_696 (O_696,N_9139,N_9925);
nand UO_697 (O_697,N_9510,N_9670);
or UO_698 (O_698,N_9407,N_9996);
or UO_699 (O_699,N_9158,N_9533);
xnor UO_700 (O_700,N_9677,N_9281);
xnor UO_701 (O_701,N_9113,N_9231);
xor UO_702 (O_702,N_9669,N_9495);
and UO_703 (O_703,N_9798,N_9562);
and UO_704 (O_704,N_9236,N_9643);
xor UO_705 (O_705,N_9292,N_9661);
nand UO_706 (O_706,N_9219,N_9700);
and UO_707 (O_707,N_9598,N_9456);
nand UO_708 (O_708,N_9272,N_9865);
xor UO_709 (O_709,N_9985,N_9976);
or UO_710 (O_710,N_9766,N_9995);
and UO_711 (O_711,N_9380,N_9273);
xnor UO_712 (O_712,N_9128,N_9268);
xnor UO_713 (O_713,N_9165,N_9556);
nor UO_714 (O_714,N_9413,N_9118);
nor UO_715 (O_715,N_9000,N_9469);
nand UO_716 (O_716,N_9471,N_9342);
nand UO_717 (O_717,N_9750,N_9503);
xnor UO_718 (O_718,N_9992,N_9781);
nor UO_719 (O_719,N_9235,N_9801);
xor UO_720 (O_720,N_9642,N_9893);
or UO_721 (O_721,N_9179,N_9019);
nor UO_722 (O_722,N_9541,N_9512);
and UO_723 (O_723,N_9261,N_9276);
and UO_724 (O_724,N_9885,N_9762);
xnor UO_725 (O_725,N_9968,N_9959);
and UO_726 (O_726,N_9089,N_9230);
nand UO_727 (O_727,N_9466,N_9244);
nor UO_728 (O_728,N_9276,N_9591);
and UO_729 (O_729,N_9163,N_9044);
or UO_730 (O_730,N_9627,N_9455);
nand UO_731 (O_731,N_9040,N_9180);
xor UO_732 (O_732,N_9895,N_9348);
and UO_733 (O_733,N_9734,N_9110);
or UO_734 (O_734,N_9067,N_9321);
nand UO_735 (O_735,N_9195,N_9078);
nor UO_736 (O_736,N_9533,N_9311);
nand UO_737 (O_737,N_9194,N_9812);
and UO_738 (O_738,N_9399,N_9883);
nand UO_739 (O_739,N_9403,N_9200);
nor UO_740 (O_740,N_9145,N_9402);
and UO_741 (O_741,N_9855,N_9451);
and UO_742 (O_742,N_9323,N_9657);
nor UO_743 (O_743,N_9934,N_9083);
nand UO_744 (O_744,N_9171,N_9972);
and UO_745 (O_745,N_9554,N_9028);
nand UO_746 (O_746,N_9948,N_9003);
nor UO_747 (O_747,N_9994,N_9175);
and UO_748 (O_748,N_9923,N_9325);
nor UO_749 (O_749,N_9086,N_9636);
xor UO_750 (O_750,N_9289,N_9218);
and UO_751 (O_751,N_9624,N_9587);
xor UO_752 (O_752,N_9096,N_9782);
nor UO_753 (O_753,N_9567,N_9751);
xnor UO_754 (O_754,N_9930,N_9500);
nand UO_755 (O_755,N_9547,N_9485);
nand UO_756 (O_756,N_9441,N_9070);
or UO_757 (O_757,N_9008,N_9428);
nor UO_758 (O_758,N_9849,N_9759);
or UO_759 (O_759,N_9997,N_9682);
nand UO_760 (O_760,N_9490,N_9278);
xor UO_761 (O_761,N_9466,N_9783);
xnor UO_762 (O_762,N_9310,N_9850);
xor UO_763 (O_763,N_9948,N_9313);
nand UO_764 (O_764,N_9565,N_9532);
or UO_765 (O_765,N_9500,N_9124);
nor UO_766 (O_766,N_9121,N_9184);
nor UO_767 (O_767,N_9238,N_9897);
or UO_768 (O_768,N_9806,N_9132);
nand UO_769 (O_769,N_9512,N_9025);
and UO_770 (O_770,N_9685,N_9961);
nand UO_771 (O_771,N_9455,N_9536);
nand UO_772 (O_772,N_9268,N_9800);
xor UO_773 (O_773,N_9357,N_9315);
or UO_774 (O_774,N_9165,N_9187);
or UO_775 (O_775,N_9319,N_9022);
nor UO_776 (O_776,N_9146,N_9868);
or UO_777 (O_777,N_9611,N_9230);
nand UO_778 (O_778,N_9189,N_9102);
nor UO_779 (O_779,N_9828,N_9037);
nor UO_780 (O_780,N_9839,N_9760);
nand UO_781 (O_781,N_9597,N_9063);
xor UO_782 (O_782,N_9378,N_9076);
nand UO_783 (O_783,N_9680,N_9891);
nand UO_784 (O_784,N_9628,N_9088);
nor UO_785 (O_785,N_9930,N_9856);
nor UO_786 (O_786,N_9095,N_9689);
and UO_787 (O_787,N_9127,N_9010);
nor UO_788 (O_788,N_9002,N_9566);
xnor UO_789 (O_789,N_9731,N_9080);
and UO_790 (O_790,N_9372,N_9652);
nor UO_791 (O_791,N_9047,N_9262);
nand UO_792 (O_792,N_9521,N_9347);
nand UO_793 (O_793,N_9916,N_9699);
and UO_794 (O_794,N_9319,N_9868);
nand UO_795 (O_795,N_9233,N_9248);
nand UO_796 (O_796,N_9555,N_9437);
nor UO_797 (O_797,N_9416,N_9486);
xor UO_798 (O_798,N_9586,N_9818);
nand UO_799 (O_799,N_9468,N_9948);
xor UO_800 (O_800,N_9957,N_9758);
nor UO_801 (O_801,N_9577,N_9472);
or UO_802 (O_802,N_9132,N_9992);
nand UO_803 (O_803,N_9189,N_9971);
nor UO_804 (O_804,N_9085,N_9317);
nand UO_805 (O_805,N_9522,N_9866);
or UO_806 (O_806,N_9986,N_9120);
or UO_807 (O_807,N_9523,N_9198);
nor UO_808 (O_808,N_9431,N_9531);
xor UO_809 (O_809,N_9858,N_9173);
nor UO_810 (O_810,N_9851,N_9604);
nor UO_811 (O_811,N_9060,N_9780);
nor UO_812 (O_812,N_9131,N_9589);
xnor UO_813 (O_813,N_9614,N_9227);
nand UO_814 (O_814,N_9497,N_9106);
xnor UO_815 (O_815,N_9263,N_9005);
nor UO_816 (O_816,N_9586,N_9943);
nor UO_817 (O_817,N_9640,N_9087);
or UO_818 (O_818,N_9996,N_9751);
and UO_819 (O_819,N_9148,N_9137);
and UO_820 (O_820,N_9253,N_9729);
and UO_821 (O_821,N_9846,N_9218);
nand UO_822 (O_822,N_9287,N_9396);
or UO_823 (O_823,N_9933,N_9006);
nor UO_824 (O_824,N_9313,N_9459);
or UO_825 (O_825,N_9527,N_9214);
and UO_826 (O_826,N_9156,N_9489);
and UO_827 (O_827,N_9200,N_9977);
and UO_828 (O_828,N_9737,N_9463);
nor UO_829 (O_829,N_9772,N_9680);
nor UO_830 (O_830,N_9824,N_9093);
xnor UO_831 (O_831,N_9565,N_9276);
nand UO_832 (O_832,N_9532,N_9360);
or UO_833 (O_833,N_9074,N_9332);
nor UO_834 (O_834,N_9030,N_9041);
xnor UO_835 (O_835,N_9471,N_9000);
and UO_836 (O_836,N_9958,N_9373);
or UO_837 (O_837,N_9265,N_9343);
or UO_838 (O_838,N_9125,N_9234);
and UO_839 (O_839,N_9679,N_9539);
or UO_840 (O_840,N_9550,N_9600);
xnor UO_841 (O_841,N_9283,N_9626);
or UO_842 (O_842,N_9910,N_9633);
nand UO_843 (O_843,N_9629,N_9190);
and UO_844 (O_844,N_9085,N_9845);
or UO_845 (O_845,N_9967,N_9820);
or UO_846 (O_846,N_9941,N_9172);
xor UO_847 (O_847,N_9619,N_9747);
xnor UO_848 (O_848,N_9118,N_9692);
and UO_849 (O_849,N_9780,N_9421);
nor UO_850 (O_850,N_9899,N_9454);
xnor UO_851 (O_851,N_9300,N_9026);
nor UO_852 (O_852,N_9827,N_9508);
nand UO_853 (O_853,N_9704,N_9410);
and UO_854 (O_854,N_9251,N_9180);
or UO_855 (O_855,N_9277,N_9100);
and UO_856 (O_856,N_9496,N_9748);
xnor UO_857 (O_857,N_9569,N_9123);
nor UO_858 (O_858,N_9662,N_9453);
nand UO_859 (O_859,N_9693,N_9763);
nand UO_860 (O_860,N_9247,N_9195);
nor UO_861 (O_861,N_9237,N_9435);
nor UO_862 (O_862,N_9618,N_9273);
and UO_863 (O_863,N_9432,N_9912);
and UO_864 (O_864,N_9867,N_9248);
and UO_865 (O_865,N_9673,N_9845);
or UO_866 (O_866,N_9030,N_9479);
and UO_867 (O_867,N_9461,N_9521);
and UO_868 (O_868,N_9723,N_9218);
or UO_869 (O_869,N_9995,N_9056);
nand UO_870 (O_870,N_9283,N_9863);
nand UO_871 (O_871,N_9690,N_9008);
or UO_872 (O_872,N_9690,N_9665);
nand UO_873 (O_873,N_9883,N_9817);
and UO_874 (O_874,N_9319,N_9385);
xor UO_875 (O_875,N_9861,N_9910);
nor UO_876 (O_876,N_9234,N_9416);
xor UO_877 (O_877,N_9474,N_9410);
nor UO_878 (O_878,N_9135,N_9617);
nor UO_879 (O_879,N_9312,N_9246);
nor UO_880 (O_880,N_9704,N_9013);
or UO_881 (O_881,N_9968,N_9502);
nor UO_882 (O_882,N_9422,N_9915);
and UO_883 (O_883,N_9699,N_9951);
nand UO_884 (O_884,N_9581,N_9940);
and UO_885 (O_885,N_9141,N_9798);
or UO_886 (O_886,N_9778,N_9872);
nand UO_887 (O_887,N_9644,N_9818);
xnor UO_888 (O_888,N_9941,N_9857);
or UO_889 (O_889,N_9640,N_9037);
xnor UO_890 (O_890,N_9884,N_9594);
nand UO_891 (O_891,N_9001,N_9999);
nand UO_892 (O_892,N_9524,N_9919);
and UO_893 (O_893,N_9452,N_9523);
and UO_894 (O_894,N_9320,N_9927);
nand UO_895 (O_895,N_9290,N_9123);
xnor UO_896 (O_896,N_9922,N_9573);
nor UO_897 (O_897,N_9768,N_9530);
and UO_898 (O_898,N_9376,N_9412);
or UO_899 (O_899,N_9025,N_9004);
and UO_900 (O_900,N_9720,N_9840);
nor UO_901 (O_901,N_9881,N_9958);
nand UO_902 (O_902,N_9891,N_9854);
or UO_903 (O_903,N_9914,N_9033);
nand UO_904 (O_904,N_9147,N_9372);
xnor UO_905 (O_905,N_9869,N_9558);
xor UO_906 (O_906,N_9171,N_9319);
nand UO_907 (O_907,N_9655,N_9751);
and UO_908 (O_908,N_9472,N_9601);
nand UO_909 (O_909,N_9580,N_9714);
and UO_910 (O_910,N_9886,N_9496);
and UO_911 (O_911,N_9652,N_9550);
and UO_912 (O_912,N_9074,N_9480);
or UO_913 (O_913,N_9716,N_9964);
nor UO_914 (O_914,N_9799,N_9483);
or UO_915 (O_915,N_9473,N_9420);
xor UO_916 (O_916,N_9167,N_9863);
nor UO_917 (O_917,N_9057,N_9093);
nor UO_918 (O_918,N_9504,N_9455);
nand UO_919 (O_919,N_9385,N_9960);
nor UO_920 (O_920,N_9736,N_9322);
or UO_921 (O_921,N_9607,N_9082);
nor UO_922 (O_922,N_9960,N_9690);
nor UO_923 (O_923,N_9605,N_9867);
nor UO_924 (O_924,N_9798,N_9076);
nor UO_925 (O_925,N_9472,N_9957);
xor UO_926 (O_926,N_9724,N_9428);
and UO_927 (O_927,N_9802,N_9090);
or UO_928 (O_928,N_9537,N_9425);
nand UO_929 (O_929,N_9015,N_9067);
nand UO_930 (O_930,N_9216,N_9259);
xor UO_931 (O_931,N_9562,N_9323);
nor UO_932 (O_932,N_9066,N_9876);
and UO_933 (O_933,N_9325,N_9562);
nor UO_934 (O_934,N_9222,N_9152);
or UO_935 (O_935,N_9832,N_9550);
nor UO_936 (O_936,N_9082,N_9110);
or UO_937 (O_937,N_9378,N_9374);
nand UO_938 (O_938,N_9391,N_9507);
and UO_939 (O_939,N_9801,N_9955);
or UO_940 (O_940,N_9436,N_9803);
or UO_941 (O_941,N_9750,N_9818);
nand UO_942 (O_942,N_9417,N_9214);
xor UO_943 (O_943,N_9876,N_9826);
or UO_944 (O_944,N_9278,N_9533);
nor UO_945 (O_945,N_9518,N_9689);
and UO_946 (O_946,N_9159,N_9089);
xor UO_947 (O_947,N_9411,N_9876);
xor UO_948 (O_948,N_9763,N_9344);
nand UO_949 (O_949,N_9217,N_9982);
xor UO_950 (O_950,N_9506,N_9337);
or UO_951 (O_951,N_9845,N_9106);
xnor UO_952 (O_952,N_9372,N_9725);
or UO_953 (O_953,N_9020,N_9856);
nor UO_954 (O_954,N_9263,N_9201);
or UO_955 (O_955,N_9973,N_9002);
and UO_956 (O_956,N_9486,N_9916);
xnor UO_957 (O_957,N_9197,N_9795);
and UO_958 (O_958,N_9482,N_9111);
nor UO_959 (O_959,N_9584,N_9084);
and UO_960 (O_960,N_9842,N_9960);
or UO_961 (O_961,N_9121,N_9225);
nor UO_962 (O_962,N_9509,N_9127);
nor UO_963 (O_963,N_9027,N_9650);
nor UO_964 (O_964,N_9666,N_9669);
and UO_965 (O_965,N_9404,N_9822);
and UO_966 (O_966,N_9401,N_9739);
xor UO_967 (O_967,N_9823,N_9152);
or UO_968 (O_968,N_9926,N_9011);
nand UO_969 (O_969,N_9220,N_9227);
xor UO_970 (O_970,N_9099,N_9845);
or UO_971 (O_971,N_9255,N_9435);
and UO_972 (O_972,N_9680,N_9555);
and UO_973 (O_973,N_9931,N_9232);
and UO_974 (O_974,N_9191,N_9975);
nand UO_975 (O_975,N_9583,N_9090);
or UO_976 (O_976,N_9173,N_9594);
or UO_977 (O_977,N_9388,N_9922);
nor UO_978 (O_978,N_9528,N_9553);
xor UO_979 (O_979,N_9173,N_9090);
or UO_980 (O_980,N_9381,N_9847);
xor UO_981 (O_981,N_9685,N_9370);
nand UO_982 (O_982,N_9590,N_9449);
or UO_983 (O_983,N_9931,N_9114);
nor UO_984 (O_984,N_9673,N_9544);
and UO_985 (O_985,N_9769,N_9093);
nand UO_986 (O_986,N_9713,N_9251);
nand UO_987 (O_987,N_9006,N_9012);
or UO_988 (O_988,N_9357,N_9588);
and UO_989 (O_989,N_9933,N_9640);
nand UO_990 (O_990,N_9296,N_9488);
nor UO_991 (O_991,N_9652,N_9605);
xor UO_992 (O_992,N_9558,N_9881);
and UO_993 (O_993,N_9565,N_9822);
nor UO_994 (O_994,N_9139,N_9049);
nand UO_995 (O_995,N_9399,N_9610);
xnor UO_996 (O_996,N_9530,N_9707);
nor UO_997 (O_997,N_9770,N_9964);
and UO_998 (O_998,N_9138,N_9790);
nor UO_999 (O_999,N_9494,N_9162);
and UO_1000 (O_1000,N_9991,N_9577);
xnor UO_1001 (O_1001,N_9962,N_9289);
and UO_1002 (O_1002,N_9570,N_9411);
and UO_1003 (O_1003,N_9983,N_9543);
and UO_1004 (O_1004,N_9646,N_9656);
nand UO_1005 (O_1005,N_9331,N_9303);
xor UO_1006 (O_1006,N_9733,N_9265);
xnor UO_1007 (O_1007,N_9096,N_9177);
xor UO_1008 (O_1008,N_9988,N_9139);
xor UO_1009 (O_1009,N_9418,N_9534);
nor UO_1010 (O_1010,N_9685,N_9930);
or UO_1011 (O_1011,N_9893,N_9169);
nor UO_1012 (O_1012,N_9789,N_9466);
nand UO_1013 (O_1013,N_9259,N_9205);
and UO_1014 (O_1014,N_9963,N_9233);
nor UO_1015 (O_1015,N_9400,N_9938);
or UO_1016 (O_1016,N_9728,N_9839);
nand UO_1017 (O_1017,N_9356,N_9653);
nor UO_1018 (O_1018,N_9029,N_9613);
and UO_1019 (O_1019,N_9030,N_9190);
nand UO_1020 (O_1020,N_9492,N_9114);
nand UO_1021 (O_1021,N_9129,N_9826);
nor UO_1022 (O_1022,N_9211,N_9979);
or UO_1023 (O_1023,N_9326,N_9725);
nand UO_1024 (O_1024,N_9735,N_9766);
nor UO_1025 (O_1025,N_9773,N_9461);
or UO_1026 (O_1026,N_9674,N_9393);
nor UO_1027 (O_1027,N_9767,N_9578);
nand UO_1028 (O_1028,N_9064,N_9455);
nor UO_1029 (O_1029,N_9711,N_9315);
nor UO_1030 (O_1030,N_9434,N_9804);
nor UO_1031 (O_1031,N_9518,N_9486);
nand UO_1032 (O_1032,N_9775,N_9017);
and UO_1033 (O_1033,N_9346,N_9314);
nor UO_1034 (O_1034,N_9290,N_9546);
xnor UO_1035 (O_1035,N_9823,N_9168);
or UO_1036 (O_1036,N_9810,N_9842);
or UO_1037 (O_1037,N_9009,N_9458);
nand UO_1038 (O_1038,N_9741,N_9810);
nand UO_1039 (O_1039,N_9553,N_9029);
nand UO_1040 (O_1040,N_9491,N_9356);
or UO_1041 (O_1041,N_9338,N_9651);
and UO_1042 (O_1042,N_9676,N_9423);
nand UO_1043 (O_1043,N_9592,N_9626);
and UO_1044 (O_1044,N_9703,N_9916);
or UO_1045 (O_1045,N_9686,N_9382);
and UO_1046 (O_1046,N_9491,N_9720);
nand UO_1047 (O_1047,N_9320,N_9536);
or UO_1048 (O_1048,N_9976,N_9045);
nand UO_1049 (O_1049,N_9621,N_9861);
and UO_1050 (O_1050,N_9900,N_9119);
nor UO_1051 (O_1051,N_9758,N_9803);
nand UO_1052 (O_1052,N_9277,N_9353);
nor UO_1053 (O_1053,N_9244,N_9665);
and UO_1054 (O_1054,N_9976,N_9057);
and UO_1055 (O_1055,N_9653,N_9682);
and UO_1056 (O_1056,N_9797,N_9917);
or UO_1057 (O_1057,N_9336,N_9501);
nor UO_1058 (O_1058,N_9582,N_9631);
nor UO_1059 (O_1059,N_9933,N_9236);
and UO_1060 (O_1060,N_9056,N_9973);
nand UO_1061 (O_1061,N_9113,N_9233);
or UO_1062 (O_1062,N_9026,N_9002);
nor UO_1063 (O_1063,N_9122,N_9356);
nand UO_1064 (O_1064,N_9273,N_9105);
or UO_1065 (O_1065,N_9199,N_9453);
nand UO_1066 (O_1066,N_9725,N_9516);
nand UO_1067 (O_1067,N_9832,N_9694);
nor UO_1068 (O_1068,N_9102,N_9302);
or UO_1069 (O_1069,N_9665,N_9722);
nor UO_1070 (O_1070,N_9596,N_9777);
nand UO_1071 (O_1071,N_9314,N_9393);
or UO_1072 (O_1072,N_9814,N_9855);
nor UO_1073 (O_1073,N_9596,N_9854);
nor UO_1074 (O_1074,N_9696,N_9008);
xor UO_1075 (O_1075,N_9144,N_9447);
or UO_1076 (O_1076,N_9027,N_9859);
or UO_1077 (O_1077,N_9378,N_9732);
or UO_1078 (O_1078,N_9465,N_9905);
nand UO_1079 (O_1079,N_9046,N_9487);
or UO_1080 (O_1080,N_9064,N_9617);
nand UO_1081 (O_1081,N_9458,N_9371);
xor UO_1082 (O_1082,N_9979,N_9265);
nand UO_1083 (O_1083,N_9385,N_9559);
nand UO_1084 (O_1084,N_9092,N_9461);
xor UO_1085 (O_1085,N_9950,N_9481);
nand UO_1086 (O_1086,N_9607,N_9002);
xor UO_1087 (O_1087,N_9908,N_9023);
xnor UO_1088 (O_1088,N_9215,N_9275);
xor UO_1089 (O_1089,N_9466,N_9718);
nor UO_1090 (O_1090,N_9130,N_9668);
or UO_1091 (O_1091,N_9999,N_9793);
nor UO_1092 (O_1092,N_9119,N_9662);
xnor UO_1093 (O_1093,N_9604,N_9191);
nor UO_1094 (O_1094,N_9610,N_9249);
nand UO_1095 (O_1095,N_9091,N_9965);
xor UO_1096 (O_1096,N_9216,N_9281);
nand UO_1097 (O_1097,N_9853,N_9704);
nand UO_1098 (O_1098,N_9877,N_9995);
or UO_1099 (O_1099,N_9476,N_9153);
nand UO_1100 (O_1100,N_9977,N_9164);
nand UO_1101 (O_1101,N_9852,N_9094);
nor UO_1102 (O_1102,N_9102,N_9247);
nor UO_1103 (O_1103,N_9264,N_9093);
xor UO_1104 (O_1104,N_9605,N_9387);
xor UO_1105 (O_1105,N_9641,N_9749);
nor UO_1106 (O_1106,N_9211,N_9096);
xnor UO_1107 (O_1107,N_9029,N_9369);
and UO_1108 (O_1108,N_9767,N_9623);
nor UO_1109 (O_1109,N_9167,N_9284);
nor UO_1110 (O_1110,N_9936,N_9475);
and UO_1111 (O_1111,N_9859,N_9601);
nand UO_1112 (O_1112,N_9436,N_9742);
nand UO_1113 (O_1113,N_9666,N_9195);
nand UO_1114 (O_1114,N_9879,N_9539);
or UO_1115 (O_1115,N_9855,N_9243);
nor UO_1116 (O_1116,N_9285,N_9556);
and UO_1117 (O_1117,N_9711,N_9780);
nor UO_1118 (O_1118,N_9991,N_9862);
nor UO_1119 (O_1119,N_9351,N_9159);
nor UO_1120 (O_1120,N_9363,N_9955);
or UO_1121 (O_1121,N_9901,N_9300);
xor UO_1122 (O_1122,N_9053,N_9748);
nor UO_1123 (O_1123,N_9626,N_9930);
nand UO_1124 (O_1124,N_9916,N_9182);
and UO_1125 (O_1125,N_9397,N_9403);
nor UO_1126 (O_1126,N_9890,N_9054);
nand UO_1127 (O_1127,N_9244,N_9504);
nand UO_1128 (O_1128,N_9742,N_9575);
or UO_1129 (O_1129,N_9814,N_9722);
xor UO_1130 (O_1130,N_9434,N_9605);
nor UO_1131 (O_1131,N_9476,N_9813);
nand UO_1132 (O_1132,N_9146,N_9880);
and UO_1133 (O_1133,N_9068,N_9581);
xor UO_1134 (O_1134,N_9161,N_9855);
nand UO_1135 (O_1135,N_9907,N_9203);
and UO_1136 (O_1136,N_9670,N_9011);
xor UO_1137 (O_1137,N_9521,N_9840);
nor UO_1138 (O_1138,N_9466,N_9015);
or UO_1139 (O_1139,N_9519,N_9638);
or UO_1140 (O_1140,N_9665,N_9330);
and UO_1141 (O_1141,N_9948,N_9255);
xnor UO_1142 (O_1142,N_9475,N_9353);
or UO_1143 (O_1143,N_9381,N_9136);
and UO_1144 (O_1144,N_9255,N_9217);
or UO_1145 (O_1145,N_9059,N_9623);
xor UO_1146 (O_1146,N_9295,N_9498);
xnor UO_1147 (O_1147,N_9976,N_9642);
nor UO_1148 (O_1148,N_9569,N_9979);
xnor UO_1149 (O_1149,N_9198,N_9285);
xnor UO_1150 (O_1150,N_9278,N_9774);
and UO_1151 (O_1151,N_9542,N_9855);
or UO_1152 (O_1152,N_9108,N_9270);
and UO_1153 (O_1153,N_9501,N_9888);
nor UO_1154 (O_1154,N_9827,N_9478);
and UO_1155 (O_1155,N_9299,N_9226);
nand UO_1156 (O_1156,N_9625,N_9441);
nor UO_1157 (O_1157,N_9243,N_9422);
nor UO_1158 (O_1158,N_9606,N_9725);
xnor UO_1159 (O_1159,N_9479,N_9140);
nand UO_1160 (O_1160,N_9398,N_9841);
nor UO_1161 (O_1161,N_9556,N_9671);
nor UO_1162 (O_1162,N_9933,N_9003);
nand UO_1163 (O_1163,N_9503,N_9529);
or UO_1164 (O_1164,N_9838,N_9688);
and UO_1165 (O_1165,N_9498,N_9556);
nor UO_1166 (O_1166,N_9556,N_9835);
xor UO_1167 (O_1167,N_9351,N_9222);
and UO_1168 (O_1168,N_9688,N_9516);
nand UO_1169 (O_1169,N_9756,N_9838);
nand UO_1170 (O_1170,N_9848,N_9500);
xnor UO_1171 (O_1171,N_9356,N_9130);
and UO_1172 (O_1172,N_9318,N_9694);
and UO_1173 (O_1173,N_9375,N_9006);
nand UO_1174 (O_1174,N_9536,N_9835);
nand UO_1175 (O_1175,N_9399,N_9680);
xnor UO_1176 (O_1176,N_9802,N_9860);
and UO_1177 (O_1177,N_9793,N_9506);
and UO_1178 (O_1178,N_9216,N_9272);
or UO_1179 (O_1179,N_9133,N_9044);
nor UO_1180 (O_1180,N_9849,N_9184);
or UO_1181 (O_1181,N_9419,N_9584);
nand UO_1182 (O_1182,N_9678,N_9365);
xor UO_1183 (O_1183,N_9040,N_9292);
nor UO_1184 (O_1184,N_9257,N_9790);
xor UO_1185 (O_1185,N_9483,N_9640);
or UO_1186 (O_1186,N_9807,N_9800);
nand UO_1187 (O_1187,N_9396,N_9133);
xnor UO_1188 (O_1188,N_9387,N_9522);
nand UO_1189 (O_1189,N_9767,N_9829);
and UO_1190 (O_1190,N_9662,N_9872);
nor UO_1191 (O_1191,N_9300,N_9406);
xor UO_1192 (O_1192,N_9652,N_9431);
or UO_1193 (O_1193,N_9224,N_9701);
nand UO_1194 (O_1194,N_9772,N_9586);
nand UO_1195 (O_1195,N_9898,N_9348);
xor UO_1196 (O_1196,N_9765,N_9018);
nand UO_1197 (O_1197,N_9428,N_9225);
xnor UO_1198 (O_1198,N_9042,N_9773);
and UO_1199 (O_1199,N_9252,N_9027);
and UO_1200 (O_1200,N_9944,N_9146);
nor UO_1201 (O_1201,N_9633,N_9347);
xnor UO_1202 (O_1202,N_9282,N_9418);
xnor UO_1203 (O_1203,N_9093,N_9767);
xnor UO_1204 (O_1204,N_9818,N_9955);
nand UO_1205 (O_1205,N_9257,N_9086);
and UO_1206 (O_1206,N_9066,N_9456);
and UO_1207 (O_1207,N_9500,N_9982);
nor UO_1208 (O_1208,N_9280,N_9874);
and UO_1209 (O_1209,N_9748,N_9858);
nor UO_1210 (O_1210,N_9884,N_9320);
xor UO_1211 (O_1211,N_9935,N_9900);
xnor UO_1212 (O_1212,N_9520,N_9678);
and UO_1213 (O_1213,N_9526,N_9845);
nor UO_1214 (O_1214,N_9905,N_9913);
or UO_1215 (O_1215,N_9507,N_9099);
nand UO_1216 (O_1216,N_9673,N_9918);
xor UO_1217 (O_1217,N_9142,N_9068);
and UO_1218 (O_1218,N_9796,N_9021);
and UO_1219 (O_1219,N_9802,N_9056);
nand UO_1220 (O_1220,N_9877,N_9924);
or UO_1221 (O_1221,N_9601,N_9598);
or UO_1222 (O_1222,N_9702,N_9175);
nor UO_1223 (O_1223,N_9173,N_9652);
and UO_1224 (O_1224,N_9513,N_9822);
xor UO_1225 (O_1225,N_9962,N_9107);
nor UO_1226 (O_1226,N_9538,N_9456);
nor UO_1227 (O_1227,N_9357,N_9600);
and UO_1228 (O_1228,N_9630,N_9315);
nor UO_1229 (O_1229,N_9634,N_9201);
or UO_1230 (O_1230,N_9030,N_9682);
and UO_1231 (O_1231,N_9095,N_9570);
nor UO_1232 (O_1232,N_9018,N_9290);
nor UO_1233 (O_1233,N_9323,N_9716);
and UO_1234 (O_1234,N_9616,N_9974);
nand UO_1235 (O_1235,N_9014,N_9915);
or UO_1236 (O_1236,N_9717,N_9071);
nor UO_1237 (O_1237,N_9992,N_9013);
and UO_1238 (O_1238,N_9933,N_9338);
or UO_1239 (O_1239,N_9064,N_9171);
or UO_1240 (O_1240,N_9340,N_9989);
xor UO_1241 (O_1241,N_9690,N_9165);
nand UO_1242 (O_1242,N_9936,N_9760);
nand UO_1243 (O_1243,N_9513,N_9814);
xor UO_1244 (O_1244,N_9907,N_9776);
and UO_1245 (O_1245,N_9234,N_9118);
nor UO_1246 (O_1246,N_9511,N_9104);
nand UO_1247 (O_1247,N_9593,N_9335);
nor UO_1248 (O_1248,N_9656,N_9787);
xnor UO_1249 (O_1249,N_9552,N_9556);
xor UO_1250 (O_1250,N_9804,N_9181);
and UO_1251 (O_1251,N_9524,N_9450);
nand UO_1252 (O_1252,N_9898,N_9874);
nand UO_1253 (O_1253,N_9712,N_9148);
or UO_1254 (O_1254,N_9280,N_9345);
and UO_1255 (O_1255,N_9006,N_9740);
nand UO_1256 (O_1256,N_9904,N_9634);
nor UO_1257 (O_1257,N_9227,N_9583);
nand UO_1258 (O_1258,N_9609,N_9766);
and UO_1259 (O_1259,N_9457,N_9543);
nand UO_1260 (O_1260,N_9283,N_9449);
xor UO_1261 (O_1261,N_9121,N_9991);
and UO_1262 (O_1262,N_9055,N_9376);
or UO_1263 (O_1263,N_9367,N_9851);
or UO_1264 (O_1264,N_9347,N_9623);
nand UO_1265 (O_1265,N_9418,N_9434);
nor UO_1266 (O_1266,N_9833,N_9016);
and UO_1267 (O_1267,N_9802,N_9839);
nand UO_1268 (O_1268,N_9723,N_9427);
xnor UO_1269 (O_1269,N_9954,N_9204);
nand UO_1270 (O_1270,N_9749,N_9436);
xor UO_1271 (O_1271,N_9505,N_9533);
xnor UO_1272 (O_1272,N_9717,N_9318);
and UO_1273 (O_1273,N_9496,N_9919);
or UO_1274 (O_1274,N_9016,N_9703);
nor UO_1275 (O_1275,N_9082,N_9182);
and UO_1276 (O_1276,N_9342,N_9448);
nor UO_1277 (O_1277,N_9354,N_9776);
and UO_1278 (O_1278,N_9127,N_9571);
nor UO_1279 (O_1279,N_9707,N_9514);
nor UO_1280 (O_1280,N_9997,N_9100);
and UO_1281 (O_1281,N_9921,N_9183);
and UO_1282 (O_1282,N_9073,N_9659);
xnor UO_1283 (O_1283,N_9103,N_9984);
xnor UO_1284 (O_1284,N_9887,N_9580);
and UO_1285 (O_1285,N_9827,N_9147);
nor UO_1286 (O_1286,N_9113,N_9086);
nor UO_1287 (O_1287,N_9038,N_9016);
or UO_1288 (O_1288,N_9966,N_9295);
or UO_1289 (O_1289,N_9665,N_9580);
or UO_1290 (O_1290,N_9303,N_9143);
nand UO_1291 (O_1291,N_9865,N_9836);
nand UO_1292 (O_1292,N_9806,N_9215);
and UO_1293 (O_1293,N_9676,N_9327);
or UO_1294 (O_1294,N_9560,N_9604);
nand UO_1295 (O_1295,N_9930,N_9713);
xnor UO_1296 (O_1296,N_9810,N_9610);
nor UO_1297 (O_1297,N_9670,N_9320);
or UO_1298 (O_1298,N_9396,N_9463);
nand UO_1299 (O_1299,N_9162,N_9783);
or UO_1300 (O_1300,N_9066,N_9033);
nor UO_1301 (O_1301,N_9524,N_9209);
nand UO_1302 (O_1302,N_9037,N_9207);
or UO_1303 (O_1303,N_9992,N_9479);
nand UO_1304 (O_1304,N_9952,N_9047);
or UO_1305 (O_1305,N_9294,N_9921);
or UO_1306 (O_1306,N_9718,N_9482);
xnor UO_1307 (O_1307,N_9865,N_9266);
nor UO_1308 (O_1308,N_9028,N_9356);
and UO_1309 (O_1309,N_9796,N_9084);
nand UO_1310 (O_1310,N_9286,N_9391);
xor UO_1311 (O_1311,N_9432,N_9066);
nand UO_1312 (O_1312,N_9374,N_9500);
or UO_1313 (O_1313,N_9952,N_9785);
nand UO_1314 (O_1314,N_9723,N_9850);
xnor UO_1315 (O_1315,N_9800,N_9888);
or UO_1316 (O_1316,N_9378,N_9350);
and UO_1317 (O_1317,N_9032,N_9796);
or UO_1318 (O_1318,N_9820,N_9905);
and UO_1319 (O_1319,N_9737,N_9806);
or UO_1320 (O_1320,N_9772,N_9610);
nand UO_1321 (O_1321,N_9345,N_9203);
nand UO_1322 (O_1322,N_9445,N_9037);
or UO_1323 (O_1323,N_9417,N_9850);
nor UO_1324 (O_1324,N_9291,N_9528);
nand UO_1325 (O_1325,N_9582,N_9947);
nor UO_1326 (O_1326,N_9139,N_9300);
and UO_1327 (O_1327,N_9526,N_9639);
xor UO_1328 (O_1328,N_9523,N_9409);
nor UO_1329 (O_1329,N_9174,N_9504);
or UO_1330 (O_1330,N_9852,N_9660);
nor UO_1331 (O_1331,N_9333,N_9700);
nor UO_1332 (O_1332,N_9803,N_9096);
xnor UO_1333 (O_1333,N_9726,N_9723);
nor UO_1334 (O_1334,N_9455,N_9638);
and UO_1335 (O_1335,N_9534,N_9136);
or UO_1336 (O_1336,N_9780,N_9219);
xor UO_1337 (O_1337,N_9469,N_9779);
and UO_1338 (O_1338,N_9520,N_9828);
nor UO_1339 (O_1339,N_9519,N_9488);
nor UO_1340 (O_1340,N_9667,N_9479);
or UO_1341 (O_1341,N_9116,N_9307);
xor UO_1342 (O_1342,N_9231,N_9468);
xor UO_1343 (O_1343,N_9636,N_9478);
and UO_1344 (O_1344,N_9117,N_9529);
nor UO_1345 (O_1345,N_9122,N_9864);
nor UO_1346 (O_1346,N_9189,N_9573);
and UO_1347 (O_1347,N_9976,N_9580);
xor UO_1348 (O_1348,N_9131,N_9850);
nand UO_1349 (O_1349,N_9906,N_9391);
xor UO_1350 (O_1350,N_9730,N_9589);
nor UO_1351 (O_1351,N_9158,N_9256);
nand UO_1352 (O_1352,N_9068,N_9784);
and UO_1353 (O_1353,N_9596,N_9951);
xor UO_1354 (O_1354,N_9864,N_9234);
or UO_1355 (O_1355,N_9988,N_9435);
or UO_1356 (O_1356,N_9582,N_9373);
or UO_1357 (O_1357,N_9240,N_9258);
nand UO_1358 (O_1358,N_9200,N_9873);
nor UO_1359 (O_1359,N_9782,N_9569);
nor UO_1360 (O_1360,N_9579,N_9658);
nand UO_1361 (O_1361,N_9470,N_9710);
or UO_1362 (O_1362,N_9014,N_9882);
nand UO_1363 (O_1363,N_9198,N_9709);
nor UO_1364 (O_1364,N_9888,N_9487);
nor UO_1365 (O_1365,N_9414,N_9935);
or UO_1366 (O_1366,N_9898,N_9326);
xor UO_1367 (O_1367,N_9080,N_9608);
nand UO_1368 (O_1368,N_9011,N_9938);
or UO_1369 (O_1369,N_9429,N_9562);
xor UO_1370 (O_1370,N_9585,N_9237);
nor UO_1371 (O_1371,N_9815,N_9721);
xnor UO_1372 (O_1372,N_9642,N_9476);
and UO_1373 (O_1373,N_9827,N_9999);
nand UO_1374 (O_1374,N_9449,N_9950);
xnor UO_1375 (O_1375,N_9847,N_9336);
or UO_1376 (O_1376,N_9836,N_9254);
and UO_1377 (O_1377,N_9031,N_9734);
and UO_1378 (O_1378,N_9795,N_9555);
nand UO_1379 (O_1379,N_9551,N_9188);
or UO_1380 (O_1380,N_9371,N_9266);
and UO_1381 (O_1381,N_9367,N_9192);
or UO_1382 (O_1382,N_9888,N_9964);
nand UO_1383 (O_1383,N_9955,N_9670);
xor UO_1384 (O_1384,N_9157,N_9514);
or UO_1385 (O_1385,N_9475,N_9372);
nor UO_1386 (O_1386,N_9545,N_9944);
or UO_1387 (O_1387,N_9543,N_9259);
or UO_1388 (O_1388,N_9473,N_9589);
nand UO_1389 (O_1389,N_9440,N_9647);
or UO_1390 (O_1390,N_9456,N_9699);
nand UO_1391 (O_1391,N_9769,N_9612);
or UO_1392 (O_1392,N_9742,N_9961);
or UO_1393 (O_1393,N_9040,N_9779);
nor UO_1394 (O_1394,N_9500,N_9820);
xor UO_1395 (O_1395,N_9149,N_9142);
xnor UO_1396 (O_1396,N_9109,N_9123);
and UO_1397 (O_1397,N_9486,N_9771);
nand UO_1398 (O_1398,N_9811,N_9801);
or UO_1399 (O_1399,N_9414,N_9291);
xor UO_1400 (O_1400,N_9212,N_9606);
and UO_1401 (O_1401,N_9906,N_9886);
and UO_1402 (O_1402,N_9828,N_9018);
nor UO_1403 (O_1403,N_9564,N_9615);
or UO_1404 (O_1404,N_9563,N_9456);
or UO_1405 (O_1405,N_9468,N_9980);
or UO_1406 (O_1406,N_9152,N_9271);
xnor UO_1407 (O_1407,N_9774,N_9837);
or UO_1408 (O_1408,N_9370,N_9747);
nand UO_1409 (O_1409,N_9176,N_9625);
nor UO_1410 (O_1410,N_9720,N_9062);
nor UO_1411 (O_1411,N_9496,N_9924);
and UO_1412 (O_1412,N_9095,N_9373);
nand UO_1413 (O_1413,N_9073,N_9633);
nand UO_1414 (O_1414,N_9522,N_9428);
and UO_1415 (O_1415,N_9267,N_9758);
and UO_1416 (O_1416,N_9425,N_9582);
xnor UO_1417 (O_1417,N_9860,N_9144);
nor UO_1418 (O_1418,N_9625,N_9015);
and UO_1419 (O_1419,N_9113,N_9898);
nand UO_1420 (O_1420,N_9723,N_9522);
and UO_1421 (O_1421,N_9885,N_9578);
or UO_1422 (O_1422,N_9658,N_9614);
nor UO_1423 (O_1423,N_9337,N_9056);
and UO_1424 (O_1424,N_9573,N_9215);
and UO_1425 (O_1425,N_9012,N_9599);
xor UO_1426 (O_1426,N_9999,N_9802);
xor UO_1427 (O_1427,N_9812,N_9937);
and UO_1428 (O_1428,N_9299,N_9621);
xnor UO_1429 (O_1429,N_9340,N_9235);
xor UO_1430 (O_1430,N_9932,N_9955);
nand UO_1431 (O_1431,N_9854,N_9885);
nor UO_1432 (O_1432,N_9378,N_9166);
and UO_1433 (O_1433,N_9716,N_9316);
nand UO_1434 (O_1434,N_9594,N_9927);
nor UO_1435 (O_1435,N_9520,N_9510);
or UO_1436 (O_1436,N_9114,N_9689);
xor UO_1437 (O_1437,N_9494,N_9853);
nor UO_1438 (O_1438,N_9584,N_9048);
nand UO_1439 (O_1439,N_9238,N_9756);
and UO_1440 (O_1440,N_9981,N_9097);
xor UO_1441 (O_1441,N_9127,N_9665);
xnor UO_1442 (O_1442,N_9872,N_9993);
xnor UO_1443 (O_1443,N_9227,N_9431);
xnor UO_1444 (O_1444,N_9499,N_9774);
xnor UO_1445 (O_1445,N_9254,N_9749);
nor UO_1446 (O_1446,N_9100,N_9040);
nand UO_1447 (O_1447,N_9433,N_9860);
nor UO_1448 (O_1448,N_9723,N_9265);
xnor UO_1449 (O_1449,N_9905,N_9923);
nor UO_1450 (O_1450,N_9245,N_9451);
nand UO_1451 (O_1451,N_9127,N_9083);
or UO_1452 (O_1452,N_9029,N_9126);
nand UO_1453 (O_1453,N_9721,N_9635);
or UO_1454 (O_1454,N_9839,N_9751);
nor UO_1455 (O_1455,N_9031,N_9725);
xnor UO_1456 (O_1456,N_9215,N_9757);
nand UO_1457 (O_1457,N_9629,N_9207);
nand UO_1458 (O_1458,N_9552,N_9457);
xor UO_1459 (O_1459,N_9680,N_9039);
xor UO_1460 (O_1460,N_9853,N_9463);
xor UO_1461 (O_1461,N_9351,N_9699);
xor UO_1462 (O_1462,N_9992,N_9971);
nand UO_1463 (O_1463,N_9676,N_9105);
or UO_1464 (O_1464,N_9948,N_9243);
xor UO_1465 (O_1465,N_9732,N_9553);
nand UO_1466 (O_1466,N_9084,N_9394);
and UO_1467 (O_1467,N_9153,N_9806);
xnor UO_1468 (O_1468,N_9209,N_9802);
nand UO_1469 (O_1469,N_9440,N_9922);
nand UO_1470 (O_1470,N_9105,N_9646);
xnor UO_1471 (O_1471,N_9118,N_9420);
nand UO_1472 (O_1472,N_9654,N_9308);
nand UO_1473 (O_1473,N_9750,N_9572);
xnor UO_1474 (O_1474,N_9171,N_9419);
nor UO_1475 (O_1475,N_9750,N_9476);
or UO_1476 (O_1476,N_9093,N_9770);
xnor UO_1477 (O_1477,N_9958,N_9130);
or UO_1478 (O_1478,N_9594,N_9377);
and UO_1479 (O_1479,N_9306,N_9287);
or UO_1480 (O_1480,N_9163,N_9760);
nor UO_1481 (O_1481,N_9180,N_9168);
nor UO_1482 (O_1482,N_9672,N_9247);
nor UO_1483 (O_1483,N_9733,N_9428);
xor UO_1484 (O_1484,N_9359,N_9007);
and UO_1485 (O_1485,N_9746,N_9645);
and UO_1486 (O_1486,N_9472,N_9971);
nand UO_1487 (O_1487,N_9382,N_9240);
or UO_1488 (O_1488,N_9114,N_9618);
xor UO_1489 (O_1489,N_9484,N_9257);
or UO_1490 (O_1490,N_9901,N_9444);
xor UO_1491 (O_1491,N_9745,N_9485);
nand UO_1492 (O_1492,N_9229,N_9234);
nor UO_1493 (O_1493,N_9794,N_9916);
nor UO_1494 (O_1494,N_9273,N_9712);
nand UO_1495 (O_1495,N_9643,N_9874);
nor UO_1496 (O_1496,N_9686,N_9657);
and UO_1497 (O_1497,N_9283,N_9236);
or UO_1498 (O_1498,N_9910,N_9247);
nor UO_1499 (O_1499,N_9776,N_9409);
endmodule